module basic_1500_15000_2000_15_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1280,In_550);
and U1 (N_1,In_395,In_846);
or U2 (N_2,In_303,In_1376);
or U3 (N_3,In_196,In_718);
and U4 (N_4,In_462,In_76);
and U5 (N_5,In_696,In_692);
and U6 (N_6,In_1252,In_991);
and U7 (N_7,In_488,In_664);
or U8 (N_8,In_1258,In_1397);
nand U9 (N_9,In_1103,In_1205);
nor U10 (N_10,In_147,In_563);
nor U11 (N_11,In_1000,In_1112);
nor U12 (N_12,In_1091,In_1354);
and U13 (N_13,In_665,In_561);
and U14 (N_14,In_1032,In_157);
and U15 (N_15,In_785,In_1419);
or U16 (N_16,In_130,In_564);
or U17 (N_17,In_386,In_512);
nor U18 (N_18,In_370,In_210);
or U19 (N_19,In_1242,In_262);
xor U20 (N_20,In_458,In_389);
and U21 (N_21,In_437,In_445);
nand U22 (N_22,In_911,In_783);
nor U23 (N_23,In_1084,In_1158);
or U24 (N_24,In_64,In_493);
nor U25 (N_25,In_1235,In_39);
and U26 (N_26,In_404,In_119);
nand U27 (N_27,In_54,In_484);
or U28 (N_28,In_732,In_578);
xnor U29 (N_29,In_1073,In_1017);
and U30 (N_30,In_1014,In_155);
xnor U31 (N_31,In_1180,In_126);
xor U32 (N_32,In_609,In_1227);
or U33 (N_33,In_2,In_731);
nor U34 (N_34,In_1336,In_951);
or U35 (N_35,In_755,In_858);
nand U36 (N_36,In_1447,In_600);
and U37 (N_37,In_325,In_675);
or U38 (N_38,In_1449,In_554);
nand U39 (N_39,In_222,In_875);
nor U40 (N_40,In_91,In_188);
and U41 (N_41,In_797,In_81);
or U42 (N_42,In_1483,In_1349);
nand U43 (N_43,In_1463,In_1122);
nand U44 (N_44,In_1052,In_737);
nor U45 (N_45,In_624,In_930);
and U46 (N_46,In_888,In_574);
nand U47 (N_47,In_426,In_774);
nor U48 (N_48,In_1229,In_1391);
or U49 (N_49,In_293,In_1348);
nor U50 (N_50,In_219,In_199);
nand U51 (N_51,In_296,In_634);
nor U52 (N_52,In_801,In_656);
and U53 (N_53,In_259,In_655);
nor U54 (N_54,In_270,In_1494);
and U55 (N_55,In_114,In_419);
and U56 (N_56,In_603,In_1490);
nor U57 (N_57,In_322,In_1167);
or U58 (N_58,In_138,In_1257);
and U59 (N_59,In_1302,In_311);
or U60 (N_60,In_289,In_1069);
and U61 (N_61,In_741,In_970);
nand U62 (N_62,In_34,In_695);
nand U63 (N_63,In_337,In_691);
nor U64 (N_64,In_1159,In_1443);
and U65 (N_65,In_316,In_1466);
or U66 (N_66,In_1423,In_1212);
and U67 (N_67,In_763,In_567);
nand U68 (N_68,In_95,In_1094);
nand U69 (N_69,In_341,In_393);
or U70 (N_70,In_509,In_290);
and U71 (N_71,In_661,In_221);
or U72 (N_72,In_559,In_745);
xnor U73 (N_73,In_871,In_100);
xor U74 (N_74,In_1285,In_808);
and U75 (N_75,In_760,In_172);
and U76 (N_76,In_677,In_702);
nand U77 (N_77,In_28,In_127);
nand U78 (N_78,In_848,In_106);
nand U79 (N_79,In_1388,In_708);
nand U80 (N_80,In_1183,In_145);
xnor U81 (N_81,In_709,In_814);
or U82 (N_82,In_403,In_457);
nor U83 (N_83,In_1362,In_979);
and U84 (N_84,In_510,In_189);
or U85 (N_85,In_1221,In_816);
nor U86 (N_86,In_101,In_821);
and U87 (N_87,In_418,In_1291);
nor U88 (N_88,In_1327,In_365);
or U89 (N_89,In_77,In_357);
or U90 (N_90,In_1346,In_998);
or U91 (N_91,In_1199,In_997);
or U92 (N_92,In_1030,In_949);
nand U93 (N_93,In_793,In_1013);
or U94 (N_94,In_534,In_1117);
and U95 (N_95,In_16,In_21);
nor U96 (N_96,In_838,In_1437);
or U97 (N_97,In_1128,In_1131);
nor U98 (N_98,In_1312,In_533);
nor U99 (N_99,In_546,In_562);
nand U100 (N_100,In_133,In_569);
xnor U101 (N_101,In_477,In_608);
nor U102 (N_102,In_233,In_672);
nor U103 (N_103,In_439,In_1427);
nor U104 (N_104,In_1365,In_582);
nor U105 (N_105,In_985,In_809);
or U106 (N_106,In_447,In_1216);
nand U107 (N_107,In_208,In_381);
nor U108 (N_108,In_1109,In_1055);
and U109 (N_109,In_165,In_822);
or U110 (N_110,In_1012,In_1080);
xnor U111 (N_111,In_1224,In_1234);
nor U112 (N_112,In_1297,In_148);
or U113 (N_113,In_944,In_74);
nand U114 (N_114,In_31,In_441);
nor U115 (N_115,In_1037,In_623);
or U116 (N_116,In_383,In_799);
nand U117 (N_117,In_297,In_1428);
and U118 (N_118,In_1123,In_922);
nand U119 (N_119,In_121,In_1150);
nor U120 (N_120,In_110,In_935);
nand U121 (N_121,In_707,In_11);
and U122 (N_122,In_1414,In_1139);
and U123 (N_123,In_1144,In_266);
nand U124 (N_124,In_179,In_1157);
and U125 (N_125,In_1422,In_865);
or U126 (N_126,In_1284,In_32);
nand U127 (N_127,In_849,In_780);
and U128 (N_128,In_693,In_630);
xor U129 (N_129,In_1099,In_628);
and U130 (N_130,In_1175,In_1185);
nor U131 (N_131,In_933,In_787);
or U132 (N_132,In_1200,In_1);
xnor U133 (N_133,In_375,In_195);
xor U134 (N_134,In_859,In_857);
nand U135 (N_135,In_1281,In_1138);
and U136 (N_136,In_648,In_321);
nor U137 (N_137,In_115,In_1236);
xnor U138 (N_138,In_1021,In_1342);
and U139 (N_139,In_1279,In_894);
nor U140 (N_140,In_1344,In_1060);
xor U141 (N_141,In_1196,In_1390);
nor U142 (N_142,In_1385,In_1083);
nor U143 (N_143,In_1398,In_679);
nand U144 (N_144,In_752,In_908);
or U145 (N_145,In_214,In_42);
nor U146 (N_146,In_759,In_831);
and U147 (N_147,In_850,In_962);
xor U148 (N_148,In_1337,In_862);
nor U149 (N_149,In_4,In_876);
or U150 (N_150,In_1309,In_728);
nand U151 (N_151,In_586,In_536);
and U152 (N_152,In_192,In_637);
and U153 (N_153,In_1033,In_256);
nor U154 (N_154,In_1356,In_1201);
nor U155 (N_155,In_1053,In_599);
and U156 (N_156,In_7,In_466);
nor U157 (N_157,In_463,In_1088);
and U158 (N_158,In_873,In_1107);
nor U159 (N_159,In_73,In_1186);
nor U160 (N_160,In_1417,In_1317);
xnor U161 (N_161,In_1481,In_1089);
or U162 (N_162,In_346,In_972);
or U163 (N_163,In_182,In_963);
and U164 (N_164,In_593,In_87);
xor U165 (N_165,In_913,In_1323);
nand U166 (N_166,In_354,In_711);
nand U167 (N_167,In_726,In_482);
nor U168 (N_168,In_680,In_1016);
and U169 (N_169,In_670,In_585);
nor U170 (N_170,In_543,In_532);
and U171 (N_171,In_812,In_722);
and U172 (N_172,In_423,In_584);
and U173 (N_173,In_1334,In_430);
and U174 (N_174,In_1473,In_1497);
nor U175 (N_175,In_1179,In_1009);
and U176 (N_176,In_104,In_248);
xnor U177 (N_177,In_3,In_1047);
nor U178 (N_178,In_832,In_394);
nor U179 (N_179,In_587,In_830);
nand U180 (N_180,In_852,In_274);
nor U181 (N_181,In_24,In_1126);
nand U182 (N_182,In_452,In_471);
xnor U183 (N_183,In_761,In_377);
nor U184 (N_184,In_819,In_1005);
and U185 (N_185,In_1056,In_828);
or U186 (N_186,In_1111,In_253);
nor U187 (N_187,In_892,In_1208);
nor U188 (N_188,In_263,In_5);
or U189 (N_189,In_440,In_897);
or U190 (N_190,In_1164,In_1006);
or U191 (N_191,In_618,In_204);
nand U192 (N_192,In_1194,In_507);
and U193 (N_193,In_132,In_1496);
nor U194 (N_194,In_154,In_1045);
nor U195 (N_195,In_900,In_615);
nand U196 (N_196,In_698,In_88);
and U197 (N_197,In_1108,In_1341);
xnor U198 (N_198,In_372,In_719);
nor U199 (N_199,In_989,In_765);
or U200 (N_200,In_1277,In_235);
or U201 (N_201,In_363,In_1173);
and U202 (N_202,In_746,In_1454);
nand U203 (N_203,In_361,In_44);
and U204 (N_204,In_697,In_1311);
or U205 (N_205,In_246,In_1430);
and U206 (N_206,In_1166,In_72);
or U207 (N_207,In_1322,In_94);
nor U208 (N_208,In_1024,In_893);
and U209 (N_209,In_1036,In_459);
nor U210 (N_210,In_841,In_443);
nor U211 (N_211,In_607,In_1031);
or U212 (N_212,In_1364,In_58);
and U213 (N_213,In_1352,In_59);
nor U214 (N_214,In_583,In_973);
nand U215 (N_215,In_861,In_685);
and U216 (N_216,In_197,In_90);
nor U217 (N_217,In_710,In_1151);
xnor U218 (N_218,In_268,In_521);
or U219 (N_219,In_448,In_653);
nor U220 (N_220,In_1455,In_1161);
nor U221 (N_221,In_391,In_1113);
and U222 (N_222,In_771,In_1412);
or U223 (N_223,In_588,In_1207);
nand U224 (N_224,In_47,In_514);
nor U225 (N_225,In_498,In_735);
and U226 (N_226,In_629,In_261);
nor U227 (N_227,In_1498,In_98);
or U228 (N_228,In_880,In_1004);
nor U229 (N_229,In_264,In_201);
or U230 (N_230,In_1406,In_48);
xor U231 (N_231,In_175,In_1071);
and U232 (N_232,In_597,In_1238);
xor U233 (N_233,In_1254,In_275);
nor U234 (N_234,In_224,In_1253);
or U235 (N_235,In_220,In_1171);
or U236 (N_236,In_1411,In_1424);
nand U237 (N_237,In_1038,In_312);
or U238 (N_238,In_1249,In_314);
nand U239 (N_239,In_715,In_923);
nand U240 (N_240,In_479,In_49);
and U241 (N_241,In_1008,In_557);
and U242 (N_242,In_1270,In_240);
nand U243 (N_243,In_786,In_1410);
nand U244 (N_244,In_990,In_1359);
and U245 (N_245,In_667,In_1141);
and U246 (N_246,In_8,In_886);
nand U247 (N_247,In_284,In_1172);
nor U248 (N_248,In_378,In_117);
or U249 (N_249,In_729,In_125);
nand U250 (N_250,In_171,In_733);
or U251 (N_251,In_662,In_953);
nand U252 (N_252,In_778,In_1153);
nor U253 (N_253,In_1156,In_983);
or U254 (N_254,In_565,In_400);
or U255 (N_255,In_649,In_1335);
nand U256 (N_256,In_1136,In_616);
xnor U257 (N_257,In_1450,In_896);
or U258 (N_258,In_795,In_1146);
nor U259 (N_259,In_734,In_1298);
and U260 (N_260,In_338,In_1445);
nor U261 (N_261,In_1384,In_757);
nand U262 (N_262,In_150,In_412);
and U263 (N_263,In_1010,In_1174);
nor U264 (N_264,In_1070,In_678);
or U265 (N_265,In_85,In_1321);
or U266 (N_266,In_1057,In_183);
nand U267 (N_267,In_1289,In_505);
nand U268 (N_268,In_137,In_553);
and U269 (N_269,In_927,In_347);
xor U270 (N_270,In_1408,In_218);
and U271 (N_271,In_753,In_41);
or U272 (N_272,In_328,In_837);
nand U273 (N_273,In_1195,In_511);
and U274 (N_274,In_449,In_1043);
and U275 (N_275,In_724,In_1461);
and U276 (N_276,In_503,In_800);
nand U277 (N_277,In_823,In_826);
and U278 (N_278,In_551,In_1433);
nor U279 (N_279,In_324,In_176);
or U280 (N_280,In_1370,In_113);
nor U281 (N_281,In_899,In_601);
nor U282 (N_282,In_213,In_1020);
or U283 (N_283,In_727,In_939);
nand U284 (N_284,In_869,In_181);
nor U285 (N_285,In_794,In_272);
nor U286 (N_286,In_1369,In_177);
nand U287 (N_287,In_1066,In_1134);
nor U288 (N_288,In_1377,In_621);
nor U289 (N_289,In_1137,In_15);
or U290 (N_290,In_494,In_669);
nand U291 (N_291,In_1132,In_89);
xor U292 (N_292,In_487,In_681);
and U293 (N_293,In_397,In_173);
and U294 (N_294,In_1246,In_1274);
or U295 (N_295,In_736,In_368);
nor U296 (N_296,In_1239,In_1472);
nor U297 (N_297,In_835,In_834);
xor U298 (N_298,In_1143,In_1343);
nand U299 (N_299,In_388,In_611);
and U300 (N_300,In_604,In_1092);
nor U301 (N_301,In_143,In_942);
nor U302 (N_302,In_647,In_184);
nand U303 (N_303,In_744,In_605);
nor U304 (N_304,In_1404,In_124);
nor U305 (N_305,In_782,In_93);
nand U306 (N_306,In_140,In_13);
or U307 (N_307,In_1162,In_411);
nor U308 (N_308,In_1149,In_1023);
and U309 (N_309,In_19,In_1193);
and U310 (N_310,In_1386,In_287);
and U311 (N_311,In_1303,In_552);
xnor U312 (N_312,In_356,In_1025);
or U313 (N_313,In_544,In_1256);
and U314 (N_314,In_833,In_885);
and U315 (N_315,In_988,In_572);
or U316 (N_316,In_223,In_225);
nand U317 (N_317,In_890,In_827);
nor U318 (N_318,In_1459,In_1295);
and U319 (N_319,In_1368,In_302);
or U320 (N_320,In_410,In_807);
or U321 (N_321,In_1184,In_910);
and U322 (N_322,In_1228,In_491);
nor U323 (N_323,In_1425,In_1154);
nand U324 (N_324,In_1082,In_955);
xor U325 (N_325,In_1396,In_499);
nor U326 (N_326,In_1191,In_1090);
nor U327 (N_327,In_1436,In_0);
or U328 (N_328,In_928,In_234);
nor U329 (N_329,In_163,In_1059);
and U330 (N_330,In_1018,In_977);
nand U331 (N_331,In_690,In_9);
nand U332 (N_332,In_999,In_231);
nand U333 (N_333,In_716,In_118);
nand U334 (N_334,In_1358,In_620);
and U335 (N_335,In_1273,In_829);
nand U336 (N_336,In_339,In_613);
nor U337 (N_337,In_791,In_657);
nand U338 (N_338,In_537,In_160);
xnor U339 (N_339,In_306,In_1288);
nor U340 (N_340,In_929,In_617);
xor U341 (N_341,In_650,In_631);
and U342 (N_342,In_277,In_1313);
or U343 (N_343,In_840,In_1050);
nor U344 (N_344,In_1338,In_641);
and U345 (N_345,In_103,In_269);
nor U346 (N_346,In_1292,In_467);
and U347 (N_347,In_784,In_1268);
and U348 (N_348,In_776,In_1027);
and U349 (N_349,In_326,In_666);
xor U350 (N_350,In_129,In_255);
xor U351 (N_351,In_251,In_1243);
and U352 (N_352,In_185,In_152);
nand U353 (N_353,In_229,In_515);
and U354 (N_354,In_966,In_526);
nand U355 (N_355,In_906,In_1015);
nor U356 (N_356,In_1085,In_1074);
or U357 (N_357,In_815,In_721);
xnor U358 (N_358,In_1275,In_644);
nand U359 (N_359,In_355,In_1395);
or U360 (N_360,In_1003,In_1097);
and U361 (N_361,In_362,In_359);
or U362 (N_362,In_573,In_905);
or U363 (N_363,In_1350,In_348);
xnor U364 (N_364,In_1035,In_43);
nand U365 (N_365,In_1263,In_756);
nor U366 (N_366,In_1394,In_1044);
nor U367 (N_367,In_415,In_79);
nand U368 (N_368,In_465,In_1034);
nand U369 (N_369,In_392,In_1145);
nor U370 (N_370,In_856,In_1409);
or U371 (N_371,In_1147,In_453);
nor U372 (N_372,In_872,In_1345);
and U373 (N_373,In_879,In_689);
or U374 (N_374,In_566,In_1304);
nor U375 (N_375,In_595,In_422);
nor U376 (N_376,In_686,In_946);
and U377 (N_377,In_1392,In_78);
nand U378 (N_378,In_1125,In_625);
or U379 (N_379,In_191,In_406);
or U380 (N_380,In_994,In_1078);
or U381 (N_381,In_788,In_645);
nor U382 (N_382,In_1102,In_854);
nor U383 (N_383,In_1435,In_839);
nor U384 (N_384,In_35,In_434);
nor U385 (N_385,In_1399,In_1096);
or U386 (N_386,In_775,In_947);
nor U387 (N_387,In_14,In_70);
or U388 (N_388,In_502,In_1068);
nand U389 (N_389,In_1488,In_75);
nand U390 (N_390,In_153,In_1452);
and U391 (N_391,In_18,In_1181);
nand U392 (N_392,In_925,In_1415);
nand U393 (N_393,In_740,In_212);
nor U394 (N_394,In_82,In_414);
nand U395 (N_395,In_1306,In_1493);
and U396 (N_396,In_408,In_1451);
or U397 (N_397,In_436,In_340);
nand U398 (N_398,In_640,In_367);
nand U399 (N_399,In_236,In_301);
nor U400 (N_400,In_61,In_902);
nor U401 (N_401,In_450,In_20);
or U402 (N_402,In_258,In_307);
nand U403 (N_403,In_63,In_1098);
or U404 (N_404,In_1499,In_1421);
nand U405 (N_405,In_889,In_398);
nor U406 (N_406,In_190,In_739);
nor U407 (N_407,In_23,In_960);
or U408 (N_408,In_252,In_161);
xnor U409 (N_409,In_674,In_1100);
nand U410 (N_410,In_211,In_717);
and U411 (N_411,In_643,In_142);
xor U412 (N_412,In_1165,In_280);
or U413 (N_413,In_1266,In_198);
and U414 (N_414,In_602,In_571);
nor U415 (N_415,In_1440,In_592);
or U416 (N_416,In_86,In_730);
xnor U417 (N_417,In_1169,In_958);
nor U418 (N_418,In_1314,In_1371);
nand U419 (N_419,In_1290,In_489);
xor U420 (N_420,In_882,In_1357);
or U421 (N_421,In_438,In_1247);
nor U422 (N_422,In_974,In_864);
and U423 (N_423,In_1305,In_1416);
nand U424 (N_424,In_1478,In_399);
xnor U425 (N_425,In_304,In_610);
or U426 (N_426,In_1177,In_842);
or U427 (N_427,In_660,In_762);
xnor U428 (N_428,In_1403,In_1296);
nor U429 (N_429,In_642,In_995);
and U430 (N_430,In_1276,In_528);
and U431 (N_431,In_1299,In_1465);
nand U432 (N_432,In_860,In_1046);
nor U433 (N_433,In_384,In_473);
nor U434 (N_434,In_714,In_1049);
nand U435 (N_435,In_360,In_1294);
and U436 (N_436,In_334,In_435);
nor U437 (N_437,In_446,In_105);
and U438 (N_438,In_904,In_405);
xor U439 (N_439,In_1351,In_1022);
and U440 (N_440,In_817,In_1182);
or U441 (N_441,In_725,In_969);
and U442 (N_442,In_1355,In_174);
and U443 (N_443,In_811,In_144);
nand U444 (N_444,In_244,In_956);
nor U445 (N_445,In_1261,In_1124);
or U446 (N_446,In_1019,In_1468);
or U447 (N_447,In_456,In_1387);
and U448 (N_448,In_1168,In_483);
nand U449 (N_449,In_920,In_149);
nor U450 (N_450,In_1250,In_1366);
nor U451 (N_451,In_790,In_658);
nor U452 (N_452,In_345,In_936);
and U453 (N_453,In_1075,In_1218);
nand U454 (N_454,In_1203,In_92);
xnor U455 (N_455,In_984,In_964);
nor U456 (N_456,In_26,In_194);
or U457 (N_457,In_523,In_996);
nor U458 (N_458,In_60,In_1458);
nand U459 (N_459,In_706,In_506);
nand U460 (N_460,In_1215,In_843);
and U461 (N_461,In_545,In_310);
nor U462 (N_462,In_366,In_878);
nand U463 (N_463,In_684,In_123);
or U464 (N_464,In_769,In_1041);
and U465 (N_465,In_202,In_332);
and U466 (N_466,In_1495,In_429);
nor U467 (N_467,In_273,In_455);
or U468 (N_468,In_464,In_1360);
nand U469 (N_469,In_758,In_668);
nand U470 (N_470,In_1220,In_868);
or U471 (N_471,In_1269,In_283);
nor U472 (N_472,In_288,In_884);
or U473 (N_473,In_1457,In_278);
and U474 (N_474,In_671,In_1367);
and U475 (N_475,In_1347,In_136);
or U476 (N_476,In_1446,In_1120);
xnor U477 (N_477,In_141,In_638);
nor U478 (N_478,In_916,In_1223);
nand U479 (N_479,In_1320,In_333);
nand U480 (N_480,In_558,In_495);
and U481 (N_481,In_1407,In_915);
nor U482 (N_482,In_496,In_30);
nor U483 (N_483,In_1442,In_1192);
and U484 (N_484,In_1469,In_1225);
nand U485 (N_485,In_766,In_329);
nor U486 (N_486,In_317,In_619);
and U487 (N_487,In_486,In_535);
nor U488 (N_488,In_948,In_461);
xor U489 (N_489,In_612,In_1326);
nand U490 (N_490,In_17,In_46);
or U491 (N_491,In_772,In_883);
or U492 (N_492,In_206,In_295);
nand U493 (N_493,In_1431,In_318);
and U494 (N_494,In_27,In_931);
and U495 (N_495,In_1231,In_66);
or U496 (N_496,In_371,In_596);
and U497 (N_497,In_108,In_205);
and U498 (N_498,In_836,In_424);
nand U499 (N_499,In_773,In_187);
nor U500 (N_500,In_178,In_767);
nand U501 (N_501,In_1456,In_1160);
nand U502 (N_502,In_531,In_474);
nand U503 (N_503,In_217,In_961);
xor U504 (N_504,In_941,In_158);
or U505 (N_505,In_1187,In_36);
nand U506 (N_506,In_1106,In_1222);
nor U507 (N_507,In_590,In_1255);
and U508 (N_508,In_813,In_1076);
and U509 (N_509,In_825,In_1418);
or U510 (N_510,In_1011,In_1209);
nor U511 (N_511,In_903,In_1213);
or U512 (N_512,In_500,In_538);
and U513 (N_513,In_245,In_1471);
and U514 (N_514,In_622,In_156);
or U515 (N_515,In_524,In_1340);
nand U516 (N_516,In_548,In_529);
nor U517 (N_517,In_743,In_824);
nor U518 (N_518,In_200,In_1105);
nor U519 (N_519,In_891,In_792);
nor U520 (N_520,In_975,In_460);
nor U521 (N_521,In_38,In_1135);
or U522 (N_522,In_1480,In_313);
or U523 (N_523,In_1389,In_1319);
nor U524 (N_524,In_84,In_789);
xnor U525 (N_525,In_591,In_1127);
or U526 (N_526,In_1214,In_1081);
nor U527 (N_527,In_1307,In_987);
and U528 (N_528,In_1301,In_294);
nor U529 (N_529,In_993,In_128);
and U530 (N_530,In_926,In_798);
xnor U531 (N_531,In_432,In_1474);
xor U532 (N_532,In_682,In_1283);
and U533 (N_533,In_863,In_1248);
or U534 (N_534,In_986,In_750);
nand U535 (N_535,In_575,In_279);
and U536 (N_536,In_497,In_33);
nand U537 (N_537,In_1375,In_917);
or U538 (N_538,In_309,In_282);
and U539 (N_539,In_1267,In_1241);
nor U540 (N_540,In_80,In_818);
and U541 (N_541,In_1133,In_203);
nor U542 (N_542,In_1264,In_1484);
and U543 (N_543,In_687,In_1380);
and U544 (N_544,In_855,In_751);
and U545 (N_545,In_162,In_764);
nor U546 (N_546,In_139,In_877);
or U547 (N_547,In_796,In_1244);
nand U548 (N_548,In_1170,In_851);
nand U549 (N_549,In_779,In_470);
nand U550 (N_550,In_68,In_413);
and U551 (N_551,In_37,In_323);
xnor U552 (N_552,In_626,In_116);
xor U553 (N_553,In_485,In_1325);
nor U554 (N_554,In_895,In_1029);
nor U555 (N_555,In_738,In_1316);
or U556 (N_556,In_847,In_1062);
or U557 (N_557,In_659,In_980);
and U558 (N_558,In_292,In_992);
xnor U559 (N_559,In_257,In_10);
or U560 (N_560,In_382,In_673);
and U561 (N_561,In_699,In_912);
and U562 (N_562,In_1405,In_1489);
nand U563 (N_563,In_1067,In_237);
and U564 (N_564,In_227,In_50);
and U565 (N_565,In_431,In_1492);
and U566 (N_566,In_1237,In_102);
nor U567 (N_567,In_1232,In_454);
nand U568 (N_568,In_965,In_580);
or U569 (N_569,In_380,In_1028);
nand U570 (N_570,In_1233,In_519);
and U571 (N_571,In_207,In_1470);
and U572 (N_572,In_576,In_594);
xnor U573 (N_573,In_238,In_1438);
nand U574 (N_574,In_480,In_954);
and U575 (N_575,In_704,In_1042);
nor U576 (N_576,In_703,In_982);
or U577 (N_577,In_870,In_1373);
nand U578 (N_578,In_651,In_976);
nor U579 (N_579,In_1486,In_241);
nor U580 (N_580,In_409,In_1077);
or U581 (N_581,In_522,In_267);
or U582 (N_582,In_844,In_853);
nand U583 (N_583,In_560,In_1093);
and U584 (N_584,In_805,In_556);
nand U585 (N_585,In_1315,In_1300);
nand U586 (N_586,In_343,In_374);
or U587 (N_587,In_950,In_407);
nand U588 (N_588,In_705,In_376);
nor U589 (N_589,In_476,In_549);
nand U590 (N_590,In_1007,In_396);
or U591 (N_591,In_1383,In_1286);
nand U592 (N_592,In_260,In_1487);
and U593 (N_593,In_134,In_1287);
and U594 (N_594,In_12,In_636);
nor U595 (N_595,In_109,In_806);
nand U596 (N_596,In_120,In_1393);
and U597 (N_597,In_1176,In_99);
and U598 (N_598,In_614,In_901);
or U599 (N_599,In_1188,In_713);
and U600 (N_600,In_25,In_1448);
nor U601 (N_601,In_542,In_1278);
nand U602 (N_602,In_209,In_1063);
nor U603 (N_603,In_1072,In_589);
and U604 (N_604,In_1479,In_451);
or U605 (N_605,In_335,In_62);
and U606 (N_606,In_525,In_417);
and U607 (N_607,In_146,In_1217);
nand U608 (N_608,In_981,In_478);
nand U609 (N_609,In_1190,In_1482);
nand U610 (N_610,In_1485,In_1206);
xor U611 (N_611,In_387,In_701);
xnor U612 (N_612,In_1339,In_934);
nand U613 (N_613,In_1129,In_369);
nor U614 (N_614,In_286,In_444);
or U615 (N_615,In_1372,In_1230);
xor U616 (N_616,In_265,In_820);
or U617 (N_617,In_1282,In_683);
nand U618 (N_618,In_541,In_55);
or U619 (N_619,In_276,In_945);
and U620 (N_620,In_513,In_379);
and U621 (N_621,In_1119,In_6);
or U622 (N_622,In_1272,In_748);
nand U623 (N_623,In_712,In_1402);
nor U624 (N_624,In_938,In_83);
nor U625 (N_625,In_1432,In_350);
or U626 (N_626,In_254,In_1476);
nor U627 (N_627,In_1363,In_1152);
and U628 (N_628,In_579,In_720);
nand U629 (N_629,In_1260,In_1265);
nor U630 (N_630,In_285,In_291);
and U631 (N_631,In_1434,In_1331);
and U632 (N_632,In_469,In_96);
and U633 (N_633,In_508,In_358);
or U634 (N_634,In_1240,In_742);
nand U635 (N_635,In_909,In_754);
or U636 (N_636,In_131,In_349);
nor U637 (N_637,In_330,In_67);
nand U638 (N_638,In_331,In_504);
nor U639 (N_639,In_627,In_688);
or U640 (N_640,In_421,In_694);
xor U641 (N_641,In_1048,In_1401);
or U642 (N_642,In_1475,In_874);
nor U643 (N_643,In_1453,In_940);
and U644 (N_644,In_320,In_249);
nor U645 (N_645,In_40,In_952);
and U646 (N_646,In_352,In_810);
or U647 (N_647,In_887,In_1065);
and U648 (N_648,In_1271,In_45);
and U649 (N_649,In_1245,In_71);
and U650 (N_650,In_428,In_881);
nor U651 (N_651,In_69,In_57);
xnor U652 (N_652,In_232,In_1426);
or U653 (N_653,In_1101,In_420);
and U654 (N_654,In_957,In_654);
and U655 (N_655,In_107,In_1202);
xor U656 (N_656,In_804,In_353);
xor U657 (N_657,In_180,In_768);
nand U658 (N_658,In_803,In_166);
xnor U659 (N_659,In_168,In_1439);
nand U660 (N_660,In_1353,In_1259);
nand U661 (N_661,In_468,In_646);
or U662 (N_662,In_1054,In_319);
nand U663 (N_663,In_425,In_1330);
and U664 (N_664,In_159,In_228);
or U665 (N_665,In_51,In_373);
nor U666 (N_666,In_242,In_1148);
nor U667 (N_667,In_344,In_65);
or U668 (N_668,In_1163,In_170);
or U669 (N_669,In_299,In_364);
nand U670 (N_670,In_971,In_1318);
and U671 (N_671,In_1293,In_520);
nor U672 (N_672,In_781,In_416);
nand U673 (N_673,In_527,In_967);
and U674 (N_674,In_919,In_1464);
nand U675 (N_675,In_635,In_1079);
nor U676 (N_676,In_475,In_112);
and U677 (N_677,In_1142,In_639);
or U678 (N_678,In_530,In_433);
nor U679 (N_679,In_1198,In_1460);
xnor U680 (N_680,In_1333,In_401);
nand U681 (N_681,In_1310,In_151);
nor U682 (N_682,In_1178,In_250);
nand U683 (N_683,In_932,In_1058);
and U684 (N_684,In_1039,In_1491);
or U685 (N_685,In_247,In_1413);
and U686 (N_686,In_1462,In_633);
nand U687 (N_687,In_1118,In_226);
and U688 (N_688,In_652,In_1116);
nor U689 (N_689,In_427,In_492);
or U690 (N_690,In_169,In_1087);
nor U691 (N_691,In_1361,In_186);
and U692 (N_692,In_490,In_336);
or U693 (N_693,In_867,In_898);
nor U694 (N_694,In_918,In_271);
nand U695 (N_695,In_1211,In_676);
nor U696 (N_696,In_1226,In_29);
nor U697 (N_697,In_1189,In_1308);
nand U698 (N_698,In_568,In_481);
or U699 (N_699,In_1382,In_540);
nor U700 (N_700,In_700,In_111);
nand U701 (N_701,In_1026,In_1381);
or U702 (N_702,In_517,In_298);
and U703 (N_703,In_122,In_164);
and U704 (N_704,In_555,In_921);
or U705 (N_705,In_606,In_1002);
nand U706 (N_706,In_663,In_52);
nand U707 (N_707,In_539,In_402);
and U708 (N_708,In_1444,In_351);
nand U709 (N_709,In_749,In_1374);
nand U710 (N_710,In_978,In_723);
or U711 (N_711,In_1477,In_1040);
or U712 (N_712,In_968,In_914);
and U713 (N_713,In_1140,In_1086);
or U714 (N_714,In_937,In_385);
and U715 (N_715,In_1121,In_1104);
nand U716 (N_716,In_547,In_1378);
nand U717 (N_717,In_230,In_1197);
nand U718 (N_718,In_1379,In_1429);
nor U719 (N_719,In_472,In_1219);
nand U720 (N_720,In_216,In_516);
xor U721 (N_721,In_53,In_22);
xnor U722 (N_722,In_1114,In_1329);
and U723 (N_723,In_1441,In_1061);
and U724 (N_724,In_1400,In_215);
and U725 (N_725,In_135,In_1332);
and U726 (N_726,In_1251,In_501);
nor U727 (N_727,In_1110,In_518);
or U728 (N_728,In_581,In_747);
or U729 (N_729,In_1262,In_56);
nand U730 (N_730,In_315,In_1001);
nor U731 (N_731,In_802,In_1064);
and U732 (N_732,In_239,In_442);
nor U733 (N_733,In_305,In_1328);
and U734 (N_734,In_1420,In_598);
nand U735 (N_735,In_845,In_390);
nand U736 (N_736,In_632,In_577);
nand U737 (N_737,In_281,In_1115);
nand U738 (N_738,In_770,In_300);
xnor U739 (N_739,In_97,In_1204);
nor U740 (N_740,In_327,In_907);
nor U741 (N_741,In_1051,In_308);
nor U742 (N_742,In_1155,In_777);
nand U743 (N_743,In_959,In_1467);
nand U744 (N_744,In_342,In_243);
nor U745 (N_745,In_193,In_924);
or U746 (N_746,In_570,In_167);
or U747 (N_747,In_1324,In_866);
nor U748 (N_748,In_1130,In_1095);
nor U749 (N_749,In_1210,In_943);
nor U750 (N_750,In_903,In_320);
or U751 (N_751,In_1185,In_90);
nand U752 (N_752,In_259,In_206);
or U753 (N_753,In_819,In_843);
and U754 (N_754,In_1168,In_1475);
or U755 (N_755,In_1356,In_806);
nor U756 (N_756,In_1162,In_447);
nand U757 (N_757,In_1105,In_1024);
xor U758 (N_758,In_681,In_786);
nor U759 (N_759,In_154,In_586);
nor U760 (N_760,In_929,In_213);
xnor U761 (N_761,In_898,In_1353);
nand U762 (N_762,In_702,In_80);
nand U763 (N_763,In_724,In_21);
and U764 (N_764,In_1278,In_1219);
nand U765 (N_765,In_788,In_565);
xnor U766 (N_766,In_1047,In_211);
xnor U767 (N_767,In_975,In_1012);
nor U768 (N_768,In_1102,In_29);
and U769 (N_769,In_89,In_269);
or U770 (N_770,In_582,In_327);
and U771 (N_771,In_398,In_1418);
nand U772 (N_772,In_1377,In_1140);
nor U773 (N_773,In_1375,In_782);
nand U774 (N_774,In_28,In_226);
nand U775 (N_775,In_1139,In_103);
and U776 (N_776,In_537,In_1476);
nor U777 (N_777,In_1002,In_570);
and U778 (N_778,In_1337,In_1120);
nor U779 (N_779,In_950,In_1273);
and U780 (N_780,In_482,In_1364);
and U781 (N_781,In_634,In_1035);
or U782 (N_782,In_1431,In_61);
nor U783 (N_783,In_1359,In_1198);
and U784 (N_784,In_188,In_15);
nor U785 (N_785,In_1220,In_23);
and U786 (N_786,In_443,In_1063);
nor U787 (N_787,In_611,In_681);
or U788 (N_788,In_822,In_779);
nor U789 (N_789,In_146,In_575);
or U790 (N_790,In_737,In_299);
and U791 (N_791,In_696,In_1045);
or U792 (N_792,In_1415,In_998);
nand U793 (N_793,In_19,In_1200);
or U794 (N_794,In_1333,In_559);
nand U795 (N_795,In_765,In_760);
nor U796 (N_796,In_632,In_464);
and U797 (N_797,In_645,In_1108);
and U798 (N_798,In_1198,In_85);
nor U799 (N_799,In_1340,In_742);
or U800 (N_800,In_568,In_1138);
and U801 (N_801,In_1036,In_1106);
xor U802 (N_802,In_1473,In_751);
and U803 (N_803,In_1072,In_678);
and U804 (N_804,In_631,In_711);
or U805 (N_805,In_1039,In_344);
or U806 (N_806,In_1126,In_1180);
xnor U807 (N_807,In_1324,In_144);
or U808 (N_808,In_502,In_303);
nand U809 (N_809,In_619,In_1355);
or U810 (N_810,In_1070,In_1429);
nor U811 (N_811,In_257,In_1050);
nor U812 (N_812,In_1363,In_541);
xnor U813 (N_813,In_514,In_561);
or U814 (N_814,In_215,In_62);
nand U815 (N_815,In_258,In_1267);
xor U816 (N_816,In_1412,In_617);
or U817 (N_817,In_1293,In_263);
or U818 (N_818,In_1490,In_585);
and U819 (N_819,In_22,In_1497);
nand U820 (N_820,In_446,In_905);
or U821 (N_821,In_338,In_455);
or U822 (N_822,In_348,In_32);
and U823 (N_823,In_550,In_1171);
and U824 (N_824,In_1112,In_479);
nand U825 (N_825,In_339,In_178);
or U826 (N_826,In_1368,In_366);
or U827 (N_827,In_1457,In_586);
or U828 (N_828,In_1414,In_341);
nand U829 (N_829,In_1076,In_1123);
and U830 (N_830,In_1309,In_39);
nand U831 (N_831,In_1219,In_1055);
or U832 (N_832,In_863,In_439);
nand U833 (N_833,In_1084,In_758);
nor U834 (N_834,In_461,In_404);
or U835 (N_835,In_1266,In_99);
nand U836 (N_836,In_196,In_1062);
or U837 (N_837,In_213,In_1076);
nor U838 (N_838,In_405,In_803);
or U839 (N_839,In_719,In_1387);
or U840 (N_840,In_8,In_1014);
nor U841 (N_841,In_1301,In_86);
or U842 (N_842,In_1451,In_161);
or U843 (N_843,In_643,In_811);
nor U844 (N_844,In_1454,In_463);
and U845 (N_845,In_1385,In_435);
nor U846 (N_846,In_339,In_1484);
nor U847 (N_847,In_1459,In_912);
and U848 (N_848,In_870,In_941);
nand U849 (N_849,In_1191,In_422);
nand U850 (N_850,In_1286,In_1394);
nand U851 (N_851,In_1227,In_244);
or U852 (N_852,In_930,In_877);
nor U853 (N_853,In_598,In_708);
or U854 (N_854,In_131,In_947);
or U855 (N_855,In_640,In_668);
xor U856 (N_856,In_1493,In_808);
or U857 (N_857,In_717,In_1272);
and U858 (N_858,In_1221,In_1071);
nand U859 (N_859,In_477,In_257);
nor U860 (N_860,In_163,In_1487);
xnor U861 (N_861,In_0,In_1300);
nor U862 (N_862,In_1227,In_312);
and U863 (N_863,In_1000,In_1048);
nand U864 (N_864,In_746,In_493);
and U865 (N_865,In_1356,In_1050);
and U866 (N_866,In_901,In_352);
and U867 (N_867,In_1084,In_171);
xnor U868 (N_868,In_459,In_178);
or U869 (N_869,In_614,In_154);
or U870 (N_870,In_1010,In_1372);
nor U871 (N_871,In_119,In_187);
xnor U872 (N_872,In_280,In_1206);
xnor U873 (N_873,In_936,In_20);
and U874 (N_874,In_1495,In_163);
nand U875 (N_875,In_574,In_382);
nor U876 (N_876,In_224,In_812);
or U877 (N_877,In_705,In_270);
or U878 (N_878,In_531,In_262);
or U879 (N_879,In_1101,In_368);
and U880 (N_880,In_1027,In_988);
and U881 (N_881,In_1433,In_383);
and U882 (N_882,In_151,In_691);
and U883 (N_883,In_447,In_665);
nand U884 (N_884,In_384,In_954);
xor U885 (N_885,In_536,In_489);
nand U886 (N_886,In_418,In_288);
nand U887 (N_887,In_1171,In_788);
nand U888 (N_888,In_312,In_1288);
or U889 (N_889,In_271,In_940);
and U890 (N_890,In_625,In_295);
or U891 (N_891,In_1265,In_67);
nor U892 (N_892,In_1155,In_77);
nor U893 (N_893,In_1100,In_420);
and U894 (N_894,In_98,In_855);
or U895 (N_895,In_161,In_910);
and U896 (N_896,In_912,In_462);
and U897 (N_897,In_1163,In_1109);
nand U898 (N_898,In_37,In_2);
nand U899 (N_899,In_1167,In_1470);
nand U900 (N_900,In_1188,In_803);
or U901 (N_901,In_243,In_802);
and U902 (N_902,In_899,In_802);
and U903 (N_903,In_1236,In_1127);
nor U904 (N_904,In_554,In_416);
nand U905 (N_905,In_319,In_768);
nor U906 (N_906,In_1228,In_1346);
xor U907 (N_907,In_801,In_557);
xor U908 (N_908,In_188,In_1422);
or U909 (N_909,In_1084,In_1301);
and U910 (N_910,In_295,In_1348);
nor U911 (N_911,In_987,In_849);
nor U912 (N_912,In_718,In_1255);
or U913 (N_913,In_775,In_1042);
or U914 (N_914,In_1449,In_680);
nand U915 (N_915,In_1052,In_271);
nor U916 (N_916,In_1043,In_145);
nor U917 (N_917,In_1377,In_1498);
and U918 (N_918,In_156,In_965);
nand U919 (N_919,In_1333,In_959);
xnor U920 (N_920,In_1317,In_408);
nor U921 (N_921,In_459,In_566);
or U922 (N_922,In_362,In_513);
and U923 (N_923,In_1230,In_163);
xnor U924 (N_924,In_903,In_1163);
and U925 (N_925,In_964,In_630);
xnor U926 (N_926,In_735,In_689);
xnor U927 (N_927,In_632,In_833);
nand U928 (N_928,In_1190,In_702);
xnor U929 (N_929,In_1406,In_455);
or U930 (N_930,In_1477,In_748);
xnor U931 (N_931,In_619,In_617);
nor U932 (N_932,In_1497,In_1140);
nand U933 (N_933,In_1278,In_138);
or U934 (N_934,In_209,In_947);
nor U935 (N_935,In_1292,In_1134);
and U936 (N_936,In_1465,In_916);
and U937 (N_937,In_292,In_1473);
and U938 (N_938,In_97,In_1244);
or U939 (N_939,In_799,In_94);
nor U940 (N_940,In_248,In_666);
xnor U941 (N_941,In_609,In_818);
xor U942 (N_942,In_601,In_39);
xor U943 (N_943,In_453,In_4);
nand U944 (N_944,In_1161,In_678);
and U945 (N_945,In_1379,In_928);
nor U946 (N_946,In_1314,In_386);
or U947 (N_947,In_812,In_622);
xnor U948 (N_948,In_1421,In_313);
and U949 (N_949,In_316,In_949);
and U950 (N_950,In_1360,In_1442);
or U951 (N_951,In_1444,In_1014);
nand U952 (N_952,In_643,In_1265);
or U953 (N_953,In_37,In_1423);
nor U954 (N_954,In_1437,In_1288);
nand U955 (N_955,In_1193,In_1279);
nand U956 (N_956,In_718,In_908);
or U957 (N_957,In_1185,In_556);
or U958 (N_958,In_40,In_451);
nand U959 (N_959,In_21,In_1400);
or U960 (N_960,In_1123,In_186);
and U961 (N_961,In_490,In_974);
or U962 (N_962,In_2,In_491);
or U963 (N_963,In_777,In_1299);
or U964 (N_964,In_804,In_857);
nor U965 (N_965,In_980,In_311);
and U966 (N_966,In_896,In_1124);
and U967 (N_967,In_1066,In_282);
xor U968 (N_968,In_303,In_202);
nand U969 (N_969,In_862,In_1420);
or U970 (N_970,In_1452,In_572);
and U971 (N_971,In_1097,In_115);
nand U972 (N_972,In_325,In_85);
or U973 (N_973,In_612,In_1441);
nor U974 (N_974,In_721,In_195);
nand U975 (N_975,In_1399,In_650);
and U976 (N_976,In_910,In_1071);
nand U977 (N_977,In_748,In_672);
xnor U978 (N_978,In_311,In_288);
or U979 (N_979,In_1282,In_836);
or U980 (N_980,In_1065,In_72);
or U981 (N_981,In_1481,In_1114);
nor U982 (N_982,In_1474,In_1151);
nor U983 (N_983,In_77,In_171);
nand U984 (N_984,In_996,In_194);
nand U985 (N_985,In_1389,In_221);
nor U986 (N_986,In_176,In_1038);
and U987 (N_987,In_879,In_25);
or U988 (N_988,In_1416,In_6);
and U989 (N_989,In_866,In_533);
nand U990 (N_990,In_1084,In_303);
and U991 (N_991,In_588,In_447);
xor U992 (N_992,In_1248,In_860);
nand U993 (N_993,In_1012,In_266);
nor U994 (N_994,In_1289,In_896);
and U995 (N_995,In_960,In_972);
nand U996 (N_996,In_1213,In_295);
or U997 (N_997,In_1187,In_852);
nand U998 (N_998,In_523,In_1099);
xnor U999 (N_999,In_70,In_153);
nand U1000 (N_1000,N_358,N_654);
nor U1001 (N_1001,N_34,N_492);
nor U1002 (N_1002,N_81,N_897);
xnor U1003 (N_1003,N_587,N_984);
or U1004 (N_1004,N_584,N_634);
or U1005 (N_1005,N_330,N_322);
nor U1006 (N_1006,N_732,N_210);
and U1007 (N_1007,N_967,N_51);
and U1008 (N_1008,N_409,N_245);
or U1009 (N_1009,N_78,N_931);
xnor U1010 (N_1010,N_44,N_702);
or U1011 (N_1011,N_518,N_478);
nand U1012 (N_1012,N_577,N_965);
nand U1013 (N_1013,N_3,N_108);
or U1014 (N_1014,N_111,N_972);
or U1015 (N_1015,N_615,N_698);
and U1016 (N_1016,N_817,N_193);
or U1017 (N_1017,N_285,N_214);
and U1018 (N_1018,N_355,N_596);
or U1019 (N_1019,N_802,N_507);
and U1020 (N_1020,N_838,N_862);
or U1021 (N_1021,N_336,N_331);
nor U1022 (N_1022,N_181,N_77);
nor U1023 (N_1023,N_82,N_168);
nand U1024 (N_1024,N_408,N_18);
xnor U1025 (N_1025,N_858,N_808);
nand U1026 (N_1026,N_480,N_717);
nand U1027 (N_1027,N_365,N_554);
nand U1028 (N_1028,N_557,N_341);
xnor U1029 (N_1029,N_672,N_364);
and U1030 (N_1030,N_229,N_957);
and U1031 (N_1031,N_765,N_563);
nand U1032 (N_1032,N_298,N_989);
nor U1033 (N_1033,N_902,N_915);
and U1034 (N_1034,N_286,N_752);
or U1035 (N_1035,N_262,N_651);
and U1036 (N_1036,N_93,N_659);
and U1037 (N_1037,N_2,N_768);
nand U1038 (N_1038,N_813,N_169);
or U1039 (N_1039,N_661,N_421);
nand U1040 (N_1040,N_317,N_595);
nor U1041 (N_1041,N_321,N_469);
and U1042 (N_1042,N_803,N_585);
nand U1043 (N_1043,N_256,N_22);
nor U1044 (N_1044,N_738,N_38);
nor U1045 (N_1045,N_299,N_121);
or U1046 (N_1046,N_98,N_599);
xor U1047 (N_1047,N_558,N_422);
nand U1048 (N_1048,N_849,N_952);
nor U1049 (N_1049,N_104,N_880);
and U1050 (N_1050,N_995,N_243);
nor U1051 (N_1051,N_792,N_109);
and U1052 (N_1052,N_387,N_809);
and U1053 (N_1053,N_474,N_482);
nand U1054 (N_1054,N_707,N_576);
or U1055 (N_1055,N_345,N_427);
nand U1056 (N_1056,N_277,N_945);
and U1057 (N_1057,N_55,N_832);
or U1058 (N_1058,N_176,N_879);
nor U1059 (N_1059,N_332,N_288);
or U1060 (N_1060,N_130,N_338);
nand U1061 (N_1061,N_720,N_65);
and U1062 (N_1062,N_287,N_295);
and U1063 (N_1063,N_124,N_50);
nand U1064 (N_1064,N_757,N_401);
nor U1065 (N_1065,N_515,N_992);
nor U1066 (N_1066,N_419,N_5);
nand U1067 (N_1067,N_57,N_294);
and U1068 (N_1068,N_609,N_59);
and U1069 (N_1069,N_270,N_340);
xor U1070 (N_1070,N_61,N_47);
nor U1071 (N_1071,N_348,N_339);
nand U1072 (N_1072,N_377,N_994);
nand U1073 (N_1073,N_497,N_622);
nor U1074 (N_1074,N_316,N_431);
and U1075 (N_1075,N_356,N_305);
nor U1076 (N_1076,N_208,N_29);
or U1077 (N_1077,N_232,N_561);
and U1078 (N_1078,N_271,N_538);
nor U1079 (N_1079,N_882,N_929);
or U1080 (N_1080,N_451,N_147);
or U1081 (N_1081,N_135,N_905);
nor U1082 (N_1082,N_572,N_385);
nand U1083 (N_1083,N_54,N_102);
and U1084 (N_1084,N_441,N_834);
nor U1085 (N_1085,N_736,N_300);
or U1086 (N_1086,N_11,N_793);
nor U1087 (N_1087,N_63,N_827);
nor U1088 (N_1088,N_8,N_500);
and U1089 (N_1089,N_491,N_910);
nand U1090 (N_1090,N_780,N_264);
and U1091 (N_1091,N_278,N_883);
nor U1092 (N_1092,N_643,N_160);
or U1093 (N_1093,N_559,N_157);
or U1094 (N_1094,N_551,N_600);
nand U1095 (N_1095,N_140,N_904);
or U1096 (N_1096,N_199,N_627);
or U1097 (N_1097,N_112,N_632);
and U1098 (N_1098,N_19,N_620);
or U1099 (N_1099,N_947,N_73);
and U1100 (N_1100,N_32,N_840);
xnor U1101 (N_1101,N_782,N_532);
or U1102 (N_1102,N_520,N_144);
xnor U1103 (N_1103,N_23,N_443);
and U1104 (N_1104,N_624,N_850);
and U1105 (N_1105,N_417,N_280);
xnor U1106 (N_1106,N_835,N_488);
nand U1107 (N_1107,N_655,N_981);
and U1108 (N_1108,N_711,N_586);
and U1109 (N_1109,N_842,N_56);
nand U1110 (N_1110,N_254,N_242);
or U1111 (N_1111,N_787,N_819);
nor U1112 (N_1112,N_693,N_126);
nand U1113 (N_1113,N_115,N_565);
and U1114 (N_1114,N_275,N_416);
nand U1115 (N_1115,N_231,N_760);
and U1116 (N_1116,N_935,N_99);
nor U1117 (N_1117,N_446,N_129);
and U1118 (N_1118,N_454,N_978);
nor U1119 (N_1119,N_663,N_420);
and U1120 (N_1120,N_606,N_297);
or U1121 (N_1121,N_759,N_366);
and U1122 (N_1122,N_202,N_291);
xor U1123 (N_1123,N_699,N_85);
and U1124 (N_1124,N_149,N_916);
and U1125 (N_1125,N_362,N_973);
or U1126 (N_1126,N_145,N_681);
nor U1127 (N_1127,N_908,N_722);
and U1128 (N_1128,N_183,N_762);
or U1129 (N_1129,N_603,N_448);
nor U1130 (N_1130,N_658,N_589);
and U1131 (N_1131,N_456,N_453);
or U1132 (N_1132,N_594,N_150);
and U1133 (N_1133,N_540,N_821);
nand U1134 (N_1134,N_498,N_192);
and U1135 (N_1135,N_493,N_773);
nor U1136 (N_1136,N_296,N_310);
and U1137 (N_1137,N_871,N_975);
nor U1138 (N_1138,N_39,N_865);
or U1139 (N_1139,N_311,N_127);
and U1140 (N_1140,N_686,N_667);
xnor U1141 (N_1141,N_887,N_227);
or U1142 (N_1142,N_696,N_397);
xor U1143 (N_1143,N_204,N_43);
nor U1144 (N_1144,N_412,N_799);
and U1145 (N_1145,N_680,N_465);
and U1146 (N_1146,N_664,N_180);
nor U1147 (N_1147,N_822,N_388);
and U1148 (N_1148,N_928,N_544);
nand U1149 (N_1149,N_796,N_641);
and U1150 (N_1150,N_718,N_354);
or U1151 (N_1151,N_274,N_785);
nor U1152 (N_1152,N_737,N_279);
or U1153 (N_1153,N_92,N_656);
nand U1154 (N_1154,N_79,N_592);
nand U1155 (N_1155,N_900,N_963);
or U1156 (N_1156,N_826,N_607);
and U1157 (N_1157,N_537,N_896);
nor U1158 (N_1158,N_677,N_723);
xnor U1159 (N_1159,N_772,N_598);
or U1160 (N_1160,N_943,N_966);
xnor U1161 (N_1161,N_463,N_933);
and U1162 (N_1162,N_403,N_590);
or U1163 (N_1163,N_120,N_307);
xor U1164 (N_1164,N_174,N_938);
xnor U1165 (N_1165,N_450,N_996);
nor U1166 (N_1166,N_575,N_848);
nand U1167 (N_1167,N_616,N_998);
nand U1168 (N_1168,N_815,N_423);
and U1169 (N_1169,N_650,N_226);
nand U1170 (N_1170,N_314,N_619);
nand U1171 (N_1171,N_376,N_932);
xnor U1172 (N_1172,N_212,N_96);
nand U1173 (N_1173,N_791,N_539);
nand U1174 (N_1174,N_856,N_705);
nand U1175 (N_1175,N_675,N_216);
nor U1176 (N_1176,N_591,N_828);
or U1177 (N_1177,N_660,N_800);
nor U1178 (N_1178,N_178,N_26);
nor U1179 (N_1179,N_766,N_755);
or U1180 (N_1180,N_141,N_712);
xor U1181 (N_1181,N_820,N_874);
nand U1182 (N_1182,N_414,N_251);
or U1183 (N_1183,N_588,N_608);
xor U1184 (N_1184,N_342,N_843);
nor U1185 (N_1185,N_530,N_194);
or U1186 (N_1186,N_186,N_402);
or U1187 (N_1187,N_198,N_770);
or U1188 (N_1188,N_367,N_623);
and U1189 (N_1189,N_552,N_383);
xnor U1190 (N_1190,N_136,N_715);
nand U1191 (N_1191,N_241,N_741);
and U1192 (N_1192,N_349,N_116);
or U1193 (N_1193,N_602,N_425);
xor U1194 (N_1194,N_860,N_976);
nor U1195 (N_1195,N_941,N_618);
and U1196 (N_1196,N_163,N_476);
nand U1197 (N_1197,N_407,N_327);
nand U1198 (N_1198,N_101,N_162);
nor U1199 (N_1199,N_721,N_777);
and U1200 (N_1200,N_206,N_990);
xor U1201 (N_1201,N_223,N_955);
or U1202 (N_1202,N_301,N_158);
or U1203 (N_1203,N_28,N_700);
and U1204 (N_1204,N_642,N_25);
nor U1205 (N_1205,N_977,N_857);
and U1206 (N_1206,N_710,N_579);
or U1207 (N_1207,N_533,N_248);
nand U1208 (N_1208,N_909,N_570);
nor U1209 (N_1209,N_489,N_418);
or U1210 (N_1210,N_228,N_668);
and U1211 (N_1211,N_891,N_62);
and U1212 (N_1212,N_234,N_953);
nor U1213 (N_1213,N_954,N_379);
nor U1214 (N_1214,N_363,N_86);
and U1215 (N_1215,N_683,N_41);
nand U1216 (N_1216,N_939,N_747);
and U1217 (N_1217,N_528,N_119);
or U1218 (N_1218,N_968,N_805);
nor U1219 (N_1219,N_701,N_257);
nand U1220 (N_1220,N_985,N_685);
and U1221 (N_1221,N_133,N_457);
xor U1222 (N_1222,N_312,N_74);
nor U1223 (N_1223,N_714,N_824);
or U1224 (N_1224,N_727,N_903);
nor U1225 (N_1225,N_789,N_283);
and U1226 (N_1226,N_529,N_868);
or U1227 (N_1227,N_368,N_117);
nor U1228 (N_1228,N_325,N_921);
or U1229 (N_1229,N_774,N_906);
or U1230 (N_1230,N_496,N_344);
or U1231 (N_1231,N_613,N_861);
xor U1232 (N_1232,N_343,N_523);
or U1233 (N_1233,N_9,N_697);
or U1234 (N_1234,N_258,N_281);
and U1235 (N_1235,N_823,N_794);
xnor U1236 (N_1236,N_894,N_549);
and U1237 (N_1237,N_167,N_923);
nor U1238 (N_1238,N_514,N_927);
xor U1239 (N_1239,N_611,N_219);
and U1240 (N_1240,N_648,N_499);
or U1241 (N_1241,N_381,N_215);
nand U1242 (N_1242,N_36,N_31);
nor U1243 (N_1243,N_37,N_393);
nand U1244 (N_1244,N_217,N_691);
and U1245 (N_1245,N_640,N_917);
nand U1246 (N_1246,N_353,N_918);
or U1247 (N_1247,N_669,N_494);
or U1248 (N_1248,N_7,N_958);
or U1249 (N_1249,N_581,N_304);
nand U1250 (N_1250,N_201,N_653);
nor U1251 (N_1251,N_58,N_646);
xor U1252 (N_1252,N_797,N_118);
or U1253 (N_1253,N_113,N_839);
nor U1254 (N_1254,N_914,N_814);
nand U1255 (N_1255,N_550,N_52);
nor U1256 (N_1256,N_776,N_830);
and U1257 (N_1257,N_268,N_513);
or U1258 (N_1258,N_378,N_593);
nand U1259 (N_1259,N_847,N_665);
nand U1260 (N_1260,N_106,N_470);
and U1261 (N_1261,N_690,N_128);
nand U1262 (N_1262,N_290,N_266);
nor U1263 (N_1263,N_786,N_795);
xor U1264 (N_1264,N_942,N_30);
nor U1265 (N_1265,N_863,N_913);
nand U1266 (N_1266,N_175,N_153);
xor U1267 (N_1267,N_374,N_255);
nor U1268 (N_1268,N_207,N_380);
nor U1269 (N_1269,N_999,N_458);
or U1270 (N_1270,N_33,N_884);
nor U1271 (N_1271,N_676,N_709);
and U1272 (N_1272,N_761,N_728);
nand U1273 (N_1273,N_524,N_398);
nand U1274 (N_1274,N_806,N_237);
nand U1275 (N_1275,N_439,N_475);
and U1276 (N_1276,N_855,N_637);
nand U1277 (N_1277,N_983,N_224);
nor U1278 (N_1278,N_844,N_788);
or U1279 (N_1279,N_833,N_182);
nand U1280 (N_1280,N_870,N_64);
nor U1281 (N_1281,N_969,N_156);
nor U1282 (N_1282,N_644,N_886);
nor U1283 (N_1283,N_679,N_893);
and U1284 (N_1284,N_404,N_490);
or U1285 (N_1285,N_750,N_148);
or U1286 (N_1286,N_719,N_382);
and U1287 (N_1287,N_812,N_831);
or U1288 (N_1288,N_166,N_936);
nor U1289 (N_1289,N_980,N_185);
or U1290 (N_1290,N_472,N_6);
nor U1291 (N_1291,N_512,N_236);
and U1292 (N_1292,N_413,N_132);
nand U1293 (N_1293,N_437,N_764);
nor U1294 (N_1294,N_508,N_48);
and U1295 (N_1295,N_464,N_763);
xor U1296 (N_1296,N_179,N_371);
nor U1297 (N_1297,N_269,N_481);
nor U1298 (N_1298,N_359,N_926);
nor U1299 (N_1299,N_244,N_892);
and U1300 (N_1300,N_811,N_395);
and U1301 (N_1301,N_221,N_635);
or U1302 (N_1302,N_372,N_673);
nor U1303 (N_1303,N_433,N_756);
nor U1304 (N_1304,N_461,N_484);
xnor U1305 (N_1305,N_347,N_1);
and U1306 (N_1306,N_956,N_249);
or U1307 (N_1307,N_434,N_350);
nor U1308 (N_1308,N_282,N_724);
xor U1309 (N_1309,N_846,N_708);
or U1310 (N_1310,N_267,N_959);
nand U1311 (N_1311,N_265,N_987);
xnor U1312 (N_1312,N_12,N_369);
and U1313 (N_1313,N_222,N_614);
nor U1314 (N_1314,N_467,N_71);
nor U1315 (N_1315,N_922,N_601);
or U1316 (N_1316,N_107,N_293);
and U1317 (N_1317,N_522,N_432);
or U1318 (N_1318,N_466,N_315);
xnor U1319 (N_1319,N_682,N_125);
nor U1320 (N_1320,N_866,N_867);
nor U1321 (N_1321,N_621,N_373);
or U1322 (N_1322,N_20,N_542);
or U1323 (N_1323,N_318,N_829);
xor U1324 (N_1324,N_801,N_666);
nor U1325 (N_1325,N_211,N_907);
or U1326 (N_1326,N_692,N_541);
and U1327 (N_1327,N_726,N_521);
nor U1328 (N_1328,N_778,N_375);
nor U1329 (N_1329,N_754,N_114);
or U1330 (N_1330,N_946,N_562);
and U1331 (N_1331,N_986,N_852);
nor U1332 (N_1332,N_885,N_424);
nor U1333 (N_1333,N_688,N_17);
nor U1334 (N_1334,N_360,N_235);
or U1335 (N_1335,N_390,N_783);
nand U1336 (N_1336,N_810,N_88);
nor U1337 (N_1337,N_394,N_924);
nand U1338 (N_1338,N_191,N_636);
nand U1339 (N_1339,N_462,N_758);
and U1340 (N_1340,N_483,N_993);
or U1341 (N_1341,N_997,N_164);
nand U1342 (N_1342,N_988,N_535);
nor U1343 (N_1343,N_744,N_89);
or U1344 (N_1344,N_610,N_837);
nand U1345 (N_1345,N_303,N_333);
and U1346 (N_1346,N_103,N_652);
nand U1347 (N_1347,N_91,N_543);
or U1348 (N_1348,N_477,N_574);
or U1349 (N_1349,N_745,N_487);
xnor U1350 (N_1350,N_329,N_853);
and U1351 (N_1351,N_742,N_740);
or U1352 (N_1352,N_177,N_888);
nand U1353 (N_1353,N_510,N_137);
or U1354 (N_1354,N_161,N_694);
nand U1355 (N_1355,N_0,N_527);
nand U1356 (N_1356,N_435,N_638);
or U1357 (N_1357,N_818,N_657);
and U1358 (N_1358,N_69,N_964);
or U1359 (N_1359,N_70,N_495);
or U1360 (N_1360,N_190,N_771);
or U1361 (N_1361,N_877,N_152);
or U1362 (N_1362,N_962,N_400);
nor U1363 (N_1363,N_841,N_869);
nand U1364 (N_1364,N_324,N_66);
or U1365 (N_1365,N_873,N_925);
xnor U1366 (N_1366,N_184,N_449);
nor U1367 (N_1367,N_695,N_396);
nand U1368 (N_1368,N_901,N_172);
nor U1369 (N_1369,N_979,N_734);
and U1370 (N_1370,N_361,N_159);
nor U1371 (N_1371,N_671,N_239);
and U1372 (N_1372,N_670,N_511);
nand U1373 (N_1373,N_689,N_898);
nand U1374 (N_1374,N_143,N_459);
and U1375 (N_1375,N_195,N_769);
nor U1376 (N_1376,N_982,N_335);
nand U1377 (N_1377,N_87,N_233);
xnor U1378 (N_1378,N_94,N_951);
nor U1379 (N_1379,N_836,N_949);
nand U1380 (N_1380,N_875,N_426);
or U1381 (N_1381,N_134,N_571);
nand U1382 (N_1382,N_555,N_733);
nand U1383 (N_1383,N_960,N_944);
or U1384 (N_1384,N_320,N_430);
nand U1385 (N_1385,N_580,N_460);
nor U1386 (N_1386,N_674,N_319);
and U1387 (N_1387,N_384,N_974);
nand U1388 (N_1388,N_749,N_784);
xor U1389 (N_1389,N_878,N_60);
or U1390 (N_1390,N_334,N_154);
xnor U1391 (N_1391,N_509,N_735);
and U1392 (N_1392,N_415,N_790);
xnor U1393 (N_1393,N_597,N_564);
and U1394 (N_1394,N_937,N_188);
nor U1395 (N_1395,N_35,N_253);
nor U1396 (N_1396,N_501,N_309);
and U1397 (N_1397,N_452,N_630);
nand U1398 (N_1398,N_713,N_100);
or U1399 (N_1399,N_53,N_238);
nand U1400 (N_1400,N_536,N_816);
nand U1401 (N_1401,N_326,N_546);
nor U1402 (N_1402,N_876,N_105);
nor U1403 (N_1403,N_406,N_247);
xnor U1404 (N_1404,N_779,N_260);
nand U1405 (N_1405,N_547,N_525);
nor U1406 (N_1406,N_131,N_187);
nor U1407 (N_1407,N_170,N_399);
and U1408 (N_1408,N_323,N_583);
or U1409 (N_1409,N_16,N_825);
and U1410 (N_1410,N_246,N_473);
xnor U1411 (N_1411,N_502,N_218);
nor U1412 (N_1412,N_912,N_612);
or U1413 (N_1413,N_24,N_730);
nor U1414 (N_1414,N_519,N_807);
nand U1415 (N_1415,N_503,N_485);
or U1416 (N_1416,N_151,N_639);
or U1417 (N_1417,N_845,N_410);
nand U1418 (N_1418,N_526,N_328);
nand U1419 (N_1419,N_566,N_386);
xnor U1420 (N_1420,N_10,N_438);
nor U1421 (N_1421,N_225,N_436);
and U1422 (N_1422,N_142,N_479);
xnor U1423 (N_1423,N_626,N_948);
xnor U1424 (N_1424,N_569,N_205);
or U1425 (N_1425,N_556,N_370);
or U1426 (N_1426,N_748,N_568);
xnor U1427 (N_1427,N_859,N_289);
and U1428 (N_1428,N_351,N_306);
xor U1429 (N_1429,N_864,N_553);
nor U1430 (N_1430,N_617,N_716);
xnor U1431 (N_1431,N_517,N_919);
nand U1432 (N_1432,N_42,N_687);
or U1433 (N_1433,N_284,N_292);
and U1434 (N_1434,N_961,N_122);
nand U1435 (N_1435,N_46,N_200);
or U1436 (N_1436,N_445,N_171);
xor U1437 (N_1437,N_276,N_15);
nand U1438 (N_1438,N_851,N_471);
nand U1439 (N_1439,N_743,N_872);
nor U1440 (N_1440,N_895,N_313);
and U1441 (N_1441,N_684,N_703);
or U1442 (N_1442,N_911,N_213);
and U1443 (N_1443,N_920,N_173);
and U1444 (N_1444,N_189,N_625);
and U1445 (N_1445,N_560,N_196);
xor U1446 (N_1446,N_725,N_27);
nand U1447 (N_1447,N_678,N_110);
or U1448 (N_1448,N_631,N_890);
nand U1449 (N_1449,N_261,N_971);
or U1450 (N_1450,N_505,N_273);
and U1451 (N_1451,N_259,N_252);
or U1452 (N_1452,N_13,N_854);
nor U1453 (N_1453,N_899,N_352);
nand U1454 (N_1454,N_775,N_950);
and U1455 (N_1455,N_123,N_662);
nor U1456 (N_1456,N_21,N_95);
and U1457 (N_1457,N_67,N_230);
nor U1458 (N_1458,N_930,N_357);
nor U1459 (N_1459,N_83,N_731);
nand U1460 (N_1460,N_76,N_389);
xnor U1461 (N_1461,N_751,N_411);
and U1462 (N_1462,N_14,N_753);
nand U1463 (N_1463,N_506,N_49);
or U1464 (N_1464,N_308,N_991);
and U1465 (N_1465,N_80,N_197);
nand U1466 (N_1466,N_545,N_881);
nand U1467 (N_1467,N_155,N_605);
nor U1468 (N_1468,N_645,N_531);
nand U1469 (N_1469,N_68,N_567);
or U1470 (N_1470,N_767,N_405);
nor U1471 (N_1471,N_604,N_209);
and U1472 (N_1472,N_447,N_392);
nor U1473 (N_1473,N_940,N_746);
or U1474 (N_1474,N_647,N_429);
and U1475 (N_1475,N_40,N_444);
or U1476 (N_1476,N_504,N_428);
and U1477 (N_1477,N_346,N_633);
nor U1478 (N_1478,N_934,N_45);
or U1479 (N_1479,N_302,N_138);
nor U1480 (N_1480,N_146,N_75);
xnor U1481 (N_1481,N_220,N_548);
nor U1482 (N_1482,N_468,N_4);
or U1483 (N_1483,N_729,N_203);
nor U1484 (N_1484,N_649,N_578);
nand U1485 (N_1485,N_706,N_84);
nand U1486 (N_1486,N_440,N_628);
and U1487 (N_1487,N_337,N_391);
nand U1488 (N_1488,N_582,N_970);
nand U1489 (N_1489,N_97,N_455);
and U1490 (N_1490,N_165,N_90);
and U1491 (N_1491,N_263,N_704);
and U1492 (N_1492,N_739,N_573);
nand U1493 (N_1493,N_781,N_534);
nor U1494 (N_1494,N_889,N_516);
and U1495 (N_1495,N_486,N_139);
or U1496 (N_1496,N_804,N_272);
xor U1497 (N_1497,N_442,N_240);
or U1498 (N_1498,N_72,N_629);
nand U1499 (N_1499,N_798,N_250);
and U1500 (N_1500,N_873,N_474);
xnor U1501 (N_1501,N_897,N_71);
nand U1502 (N_1502,N_493,N_823);
nor U1503 (N_1503,N_718,N_664);
nand U1504 (N_1504,N_217,N_900);
nor U1505 (N_1505,N_62,N_895);
nand U1506 (N_1506,N_427,N_860);
and U1507 (N_1507,N_2,N_705);
nand U1508 (N_1508,N_372,N_83);
or U1509 (N_1509,N_402,N_495);
nor U1510 (N_1510,N_119,N_99);
nand U1511 (N_1511,N_72,N_523);
xor U1512 (N_1512,N_938,N_91);
or U1513 (N_1513,N_773,N_293);
or U1514 (N_1514,N_345,N_288);
xor U1515 (N_1515,N_452,N_437);
nor U1516 (N_1516,N_333,N_87);
and U1517 (N_1517,N_156,N_768);
or U1518 (N_1518,N_905,N_890);
nor U1519 (N_1519,N_74,N_260);
or U1520 (N_1520,N_809,N_940);
nor U1521 (N_1521,N_444,N_808);
and U1522 (N_1522,N_392,N_99);
or U1523 (N_1523,N_625,N_349);
or U1524 (N_1524,N_562,N_421);
nand U1525 (N_1525,N_309,N_600);
nor U1526 (N_1526,N_938,N_682);
and U1527 (N_1527,N_686,N_703);
nor U1528 (N_1528,N_831,N_514);
nor U1529 (N_1529,N_301,N_403);
or U1530 (N_1530,N_507,N_764);
nor U1531 (N_1531,N_40,N_331);
nand U1532 (N_1532,N_343,N_925);
or U1533 (N_1533,N_61,N_245);
nor U1534 (N_1534,N_39,N_831);
xnor U1535 (N_1535,N_740,N_695);
and U1536 (N_1536,N_81,N_619);
nor U1537 (N_1537,N_334,N_294);
nand U1538 (N_1538,N_44,N_798);
or U1539 (N_1539,N_263,N_647);
and U1540 (N_1540,N_947,N_633);
nand U1541 (N_1541,N_145,N_817);
and U1542 (N_1542,N_468,N_671);
and U1543 (N_1543,N_640,N_936);
or U1544 (N_1544,N_149,N_753);
or U1545 (N_1545,N_307,N_165);
and U1546 (N_1546,N_917,N_238);
nand U1547 (N_1547,N_906,N_779);
nor U1548 (N_1548,N_543,N_547);
nor U1549 (N_1549,N_234,N_62);
nor U1550 (N_1550,N_24,N_804);
nand U1551 (N_1551,N_724,N_775);
xor U1552 (N_1552,N_132,N_781);
and U1553 (N_1553,N_225,N_797);
or U1554 (N_1554,N_418,N_483);
and U1555 (N_1555,N_228,N_630);
nand U1556 (N_1556,N_75,N_373);
nand U1557 (N_1557,N_63,N_421);
nor U1558 (N_1558,N_644,N_362);
nor U1559 (N_1559,N_23,N_931);
nor U1560 (N_1560,N_774,N_861);
and U1561 (N_1561,N_260,N_813);
nor U1562 (N_1562,N_609,N_441);
and U1563 (N_1563,N_703,N_600);
nor U1564 (N_1564,N_337,N_770);
nand U1565 (N_1565,N_537,N_369);
nand U1566 (N_1566,N_428,N_457);
or U1567 (N_1567,N_936,N_878);
or U1568 (N_1568,N_977,N_403);
nor U1569 (N_1569,N_841,N_397);
and U1570 (N_1570,N_655,N_377);
or U1571 (N_1571,N_776,N_284);
nand U1572 (N_1572,N_107,N_42);
and U1573 (N_1573,N_13,N_23);
nor U1574 (N_1574,N_424,N_262);
nand U1575 (N_1575,N_310,N_308);
nand U1576 (N_1576,N_400,N_387);
xnor U1577 (N_1577,N_60,N_117);
or U1578 (N_1578,N_403,N_300);
nor U1579 (N_1579,N_242,N_13);
or U1580 (N_1580,N_631,N_526);
and U1581 (N_1581,N_329,N_375);
nor U1582 (N_1582,N_516,N_524);
xor U1583 (N_1583,N_40,N_238);
xnor U1584 (N_1584,N_468,N_860);
nand U1585 (N_1585,N_650,N_898);
or U1586 (N_1586,N_675,N_814);
xnor U1587 (N_1587,N_582,N_386);
nor U1588 (N_1588,N_107,N_359);
or U1589 (N_1589,N_400,N_161);
or U1590 (N_1590,N_673,N_739);
and U1591 (N_1591,N_674,N_891);
or U1592 (N_1592,N_359,N_325);
nand U1593 (N_1593,N_825,N_39);
and U1594 (N_1594,N_324,N_979);
nor U1595 (N_1595,N_768,N_755);
and U1596 (N_1596,N_538,N_54);
xnor U1597 (N_1597,N_624,N_544);
nor U1598 (N_1598,N_63,N_810);
nand U1599 (N_1599,N_697,N_495);
nor U1600 (N_1600,N_37,N_953);
xnor U1601 (N_1601,N_767,N_100);
or U1602 (N_1602,N_504,N_740);
nor U1603 (N_1603,N_45,N_407);
nor U1604 (N_1604,N_155,N_871);
or U1605 (N_1605,N_216,N_437);
xor U1606 (N_1606,N_419,N_209);
xnor U1607 (N_1607,N_653,N_406);
nor U1608 (N_1608,N_891,N_945);
or U1609 (N_1609,N_369,N_242);
and U1610 (N_1610,N_382,N_518);
xor U1611 (N_1611,N_780,N_932);
nand U1612 (N_1612,N_310,N_666);
and U1613 (N_1613,N_219,N_727);
nor U1614 (N_1614,N_572,N_515);
and U1615 (N_1615,N_821,N_424);
nand U1616 (N_1616,N_16,N_63);
nand U1617 (N_1617,N_813,N_179);
or U1618 (N_1618,N_712,N_926);
nor U1619 (N_1619,N_320,N_455);
nand U1620 (N_1620,N_163,N_618);
and U1621 (N_1621,N_845,N_797);
nand U1622 (N_1622,N_689,N_425);
or U1623 (N_1623,N_124,N_874);
or U1624 (N_1624,N_13,N_244);
and U1625 (N_1625,N_479,N_444);
nor U1626 (N_1626,N_253,N_693);
or U1627 (N_1627,N_227,N_877);
or U1628 (N_1628,N_316,N_311);
nand U1629 (N_1629,N_561,N_818);
and U1630 (N_1630,N_249,N_894);
nand U1631 (N_1631,N_688,N_777);
and U1632 (N_1632,N_766,N_45);
or U1633 (N_1633,N_931,N_167);
xor U1634 (N_1634,N_847,N_129);
and U1635 (N_1635,N_249,N_80);
or U1636 (N_1636,N_233,N_681);
nand U1637 (N_1637,N_628,N_13);
nor U1638 (N_1638,N_683,N_241);
and U1639 (N_1639,N_925,N_369);
nor U1640 (N_1640,N_231,N_581);
and U1641 (N_1641,N_202,N_780);
nand U1642 (N_1642,N_314,N_865);
or U1643 (N_1643,N_347,N_408);
and U1644 (N_1644,N_614,N_327);
and U1645 (N_1645,N_485,N_876);
nor U1646 (N_1646,N_171,N_272);
or U1647 (N_1647,N_359,N_769);
nor U1648 (N_1648,N_582,N_35);
nor U1649 (N_1649,N_593,N_432);
nor U1650 (N_1650,N_518,N_604);
nand U1651 (N_1651,N_498,N_938);
or U1652 (N_1652,N_812,N_349);
and U1653 (N_1653,N_989,N_606);
nand U1654 (N_1654,N_172,N_547);
nor U1655 (N_1655,N_542,N_630);
and U1656 (N_1656,N_615,N_502);
nand U1657 (N_1657,N_226,N_424);
and U1658 (N_1658,N_249,N_700);
or U1659 (N_1659,N_304,N_607);
nand U1660 (N_1660,N_870,N_338);
nor U1661 (N_1661,N_475,N_344);
and U1662 (N_1662,N_800,N_645);
nand U1663 (N_1663,N_631,N_188);
and U1664 (N_1664,N_588,N_50);
or U1665 (N_1665,N_244,N_86);
and U1666 (N_1666,N_671,N_610);
and U1667 (N_1667,N_488,N_937);
or U1668 (N_1668,N_933,N_756);
nor U1669 (N_1669,N_115,N_597);
xor U1670 (N_1670,N_490,N_711);
xor U1671 (N_1671,N_848,N_303);
or U1672 (N_1672,N_767,N_968);
and U1673 (N_1673,N_162,N_625);
nand U1674 (N_1674,N_690,N_920);
or U1675 (N_1675,N_194,N_6);
nand U1676 (N_1676,N_878,N_914);
and U1677 (N_1677,N_879,N_666);
or U1678 (N_1678,N_688,N_243);
nand U1679 (N_1679,N_684,N_982);
nor U1680 (N_1680,N_986,N_44);
nor U1681 (N_1681,N_239,N_619);
nor U1682 (N_1682,N_186,N_602);
nor U1683 (N_1683,N_729,N_774);
or U1684 (N_1684,N_101,N_418);
nor U1685 (N_1685,N_233,N_127);
and U1686 (N_1686,N_22,N_165);
nor U1687 (N_1687,N_978,N_365);
and U1688 (N_1688,N_363,N_938);
or U1689 (N_1689,N_692,N_101);
nor U1690 (N_1690,N_808,N_933);
nand U1691 (N_1691,N_220,N_490);
and U1692 (N_1692,N_626,N_216);
nand U1693 (N_1693,N_469,N_646);
nor U1694 (N_1694,N_443,N_711);
nand U1695 (N_1695,N_91,N_729);
nand U1696 (N_1696,N_974,N_58);
and U1697 (N_1697,N_446,N_200);
and U1698 (N_1698,N_655,N_708);
and U1699 (N_1699,N_879,N_904);
xor U1700 (N_1700,N_665,N_841);
xnor U1701 (N_1701,N_427,N_3);
and U1702 (N_1702,N_292,N_401);
or U1703 (N_1703,N_381,N_948);
xnor U1704 (N_1704,N_226,N_718);
and U1705 (N_1705,N_368,N_402);
nor U1706 (N_1706,N_25,N_329);
nand U1707 (N_1707,N_260,N_123);
nor U1708 (N_1708,N_998,N_626);
or U1709 (N_1709,N_77,N_665);
or U1710 (N_1710,N_111,N_363);
nand U1711 (N_1711,N_631,N_515);
xnor U1712 (N_1712,N_308,N_360);
nand U1713 (N_1713,N_279,N_136);
nand U1714 (N_1714,N_359,N_868);
nor U1715 (N_1715,N_413,N_92);
and U1716 (N_1716,N_819,N_400);
and U1717 (N_1717,N_558,N_937);
nor U1718 (N_1718,N_545,N_63);
or U1719 (N_1719,N_143,N_356);
xnor U1720 (N_1720,N_773,N_167);
or U1721 (N_1721,N_55,N_907);
nand U1722 (N_1722,N_182,N_304);
nand U1723 (N_1723,N_327,N_326);
nand U1724 (N_1724,N_61,N_355);
and U1725 (N_1725,N_95,N_874);
or U1726 (N_1726,N_264,N_572);
nand U1727 (N_1727,N_687,N_148);
xnor U1728 (N_1728,N_54,N_21);
or U1729 (N_1729,N_997,N_315);
and U1730 (N_1730,N_608,N_786);
nand U1731 (N_1731,N_837,N_241);
and U1732 (N_1732,N_933,N_521);
or U1733 (N_1733,N_629,N_522);
and U1734 (N_1734,N_603,N_731);
nand U1735 (N_1735,N_462,N_568);
xnor U1736 (N_1736,N_825,N_963);
nor U1737 (N_1737,N_37,N_808);
nor U1738 (N_1738,N_556,N_541);
nand U1739 (N_1739,N_878,N_61);
nor U1740 (N_1740,N_888,N_151);
or U1741 (N_1741,N_40,N_578);
nor U1742 (N_1742,N_143,N_306);
or U1743 (N_1743,N_800,N_184);
and U1744 (N_1744,N_639,N_905);
xor U1745 (N_1745,N_903,N_10);
or U1746 (N_1746,N_147,N_413);
and U1747 (N_1747,N_366,N_365);
nor U1748 (N_1748,N_242,N_169);
and U1749 (N_1749,N_611,N_105);
nand U1750 (N_1750,N_434,N_695);
nor U1751 (N_1751,N_417,N_854);
xnor U1752 (N_1752,N_515,N_398);
nand U1753 (N_1753,N_257,N_113);
nor U1754 (N_1754,N_273,N_579);
or U1755 (N_1755,N_743,N_143);
and U1756 (N_1756,N_132,N_481);
nand U1757 (N_1757,N_787,N_210);
and U1758 (N_1758,N_252,N_787);
or U1759 (N_1759,N_83,N_195);
nor U1760 (N_1760,N_976,N_970);
and U1761 (N_1761,N_547,N_353);
or U1762 (N_1762,N_894,N_807);
nand U1763 (N_1763,N_454,N_918);
nor U1764 (N_1764,N_550,N_959);
or U1765 (N_1765,N_526,N_563);
nand U1766 (N_1766,N_471,N_72);
nand U1767 (N_1767,N_842,N_102);
xnor U1768 (N_1768,N_260,N_550);
nand U1769 (N_1769,N_113,N_570);
nand U1770 (N_1770,N_390,N_205);
nor U1771 (N_1771,N_287,N_740);
nor U1772 (N_1772,N_766,N_901);
nand U1773 (N_1773,N_893,N_578);
nand U1774 (N_1774,N_577,N_876);
nand U1775 (N_1775,N_173,N_206);
or U1776 (N_1776,N_170,N_885);
and U1777 (N_1777,N_69,N_870);
xor U1778 (N_1778,N_498,N_852);
or U1779 (N_1779,N_151,N_198);
nor U1780 (N_1780,N_972,N_122);
xor U1781 (N_1781,N_523,N_793);
or U1782 (N_1782,N_804,N_184);
or U1783 (N_1783,N_903,N_367);
or U1784 (N_1784,N_988,N_423);
or U1785 (N_1785,N_582,N_370);
xnor U1786 (N_1786,N_686,N_371);
xor U1787 (N_1787,N_703,N_1);
nand U1788 (N_1788,N_445,N_14);
nand U1789 (N_1789,N_551,N_563);
and U1790 (N_1790,N_215,N_801);
or U1791 (N_1791,N_670,N_977);
and U1792 (N_1792,N_779,N_384);
xor U1793 (N_1793,N_192,N_874);
and U1794 (N_1794,N_839,N_575);
and U1795 (N_1795,N_365,N_699);
nand U1796 (N_1796,N_823,N_668);
and U1797 (N_1797,N_779,N_124);
nand U1798 (N_1798,N_535,N_294);
nor U1799 (N_1799,N_770,N_2);
and U1800 (N_1800,N_441,N_866);
xor U1801 (N_1801,N_806,N_664);
and U1802 (N_1802,N_56,N_173);
and U1803 (N_1803,N_933,N_248);
nor U1804 (N_1804,N_816,N_60);
nand U1805 (N_1805,N_752,N_849);
nor U1806 (N_1806,N_377,N_57);
and U1807 (N_1807,N_200,N_440);
nand U1808 (N_1808,N_165,N_830);
nand U1809 (N_1809,N_109,N_287);
and U1810 (N_1810,N_209,N_938);
and U1811 (N_1811,N_361,N_413);
nor U1812 (N_1812,N_818,N_433);
and U1813 (N_1813,N_580,N_390);
nor U1814 (N_1814,N_72,N_117);
and U1815 (N_1815,N_600,N_132);
nor U1816 (N_1816,N_124,N_734);
or U1817 (N_1817,N_743,N_54);
nor U1818 (N_1818,N_527,N_121);
nand U1819 (N_1819,N_40,N_461);
nor U1820 (N_1820,N_766,N_205);
nor U1821 (N_1821,N_279,N_899);
nand U1822 (N_1822,N_80,N_306);
and U1823 (N_1823,N_801,N_116);
or U1824 (N_1824,N_117,N_292);
or U1825 (N_1825,N_228,N_97);
nor U1826 (N_1826,N_777,N_158);
and U1827 (N_1827,N_479,N_568);
xnor U1828 (N_1828,N_974,N_798);
and U1829 (N_1829,N_364,N_450);
nand U1830 (N_1830,N_535,N_463);
or U1831 (N_1831,N_490,N_586);
nor U1832 (N_1832,N_771,N_779);
or U1833 (N_1833,N_80,N_560);
and U1834 (N_1834,N_286,N_59);
or U1835 (N_1835,N_309,N_997);
nand U1836 (N_1836,N_88,N_157);
and U1837 (N_1837,N_753,N_205);
and U1838 (N_1838,N_794,N_196);
nor U1839 (N_1839,N_90,N_761);
nand U1840 (N_1840,N_876,N_335);
or U1841 (N_1841,N_665,N_144);
nor U1842 (N_1842,N_286,N_334);
or U1843 (N_1843,N_621,N_222);
nand U1844 (N_1844,N_175,N_465);
or U1845 (N_1845,N_10,N_981);
xnor U1846 (N_1846,N_386,N_780);
or U1847 (N_1847,N_931,N_134);
nor U1848 (N_1848,N_673,N_700);
nor U1849 (N_1849,N_36,N_679);
nor U1850 (N_1850,N_155,N_837);
nand U1851 (N_1851,N_232,N_944);
or U1852 (N_1852,N_396,N_20);
or U1853 (N_1853,N_152,N_218);
nor U1854 (N_1854,N_325,N_412);
and U1855 (N_1855,N_477,N_458);
nor U1856 (N_1856,N_417,N_765);
nor U1857 (N_1857,N_56,N_787);
and U1858 (N_1858,N_321,N_729);
nand U1859 (N_1859,N_837,N_962);
and U1860 (N_1860,N_123,N_31);
nor U1861 (N_1861,N_574,N_653);
and U1862 (N_1862,N_524,N_638);
and U1863 (N_1863,N_163,N_44);
xnor U1864 (N_1864,N_210,N_166);
or U1865 (N_1865,N_197,N_622);
or U1866 (N_1866,N_218,N_398);
xor U1867 (N_1867,N_889,N_589);
and U1868 (N_1868,N_393,N_17);
nor U1869 (N_1869,N_567,N_570);
or U1870 (N_1870,N_887,N_341);
nor U1871 (N_1871,N_834,N_649);
or U1872 (N_1872,N_660,N_408);
xor U1873 (N_1873,N_333,N_972);
and U1874 (N_1874,N_395,N_424);
nand U1875 (N_1875,N_712,N_707);
or U1876 (N_1876,N_980,N_212);
or U1877 (N_1877,N_518,N_788);
or U1878 (N_1878,N_965,N_923);
nor U1879 (N_1879,N_18,N_428);
nor U1880 (N_1880,N_996,N_522);
or U1881 (N_1881,N_469,N_344);
nor U1882 (N_1882,N_614,N_645);
nor U1883 (N_1883,N_888,N_259);
and U1884 (N_1884,N_640,N_604);
nor U1885 (N_1885,N_169,N_466);
or U1886 (N_1886,N_749,N_435);
nor U1887 (N_1887,N_635,N_795);
or U1888 (N_1888,N_725,N_979);
and U1889 (N_1889,N_734,N_265);
xnor U1890 (N_1890,N_44,N_193);
nand U1891 (N_1891,N_115,N_673);
xnor U1892 (N_1892,N_118,N_624);
nor U1893 (N_1893,N_199,N_591);
or U1894 (N_1894,N_573,N_680);
nor U1895 (N_1895,N_619,N_674);
nor U1896 (N_1896,N_625,N_136);
nor U1897 (N_1897,N_222,N_957);
nand U1898 (N_1898,N_568,N_886);
and U1899 (N_1899,N_93,N_492);
or U1900 (N_1900,N_375,N_239);
or U1901 (N_1901,N_952,N_196);
or U1902 (N_1902,N_457,N_914);
nor U1903 (N_1903,N_243,N_601);
nor U1904 (N_1904,N_789,N_250);
nor U1905 (N_1905,N_397,N_309);
xnor U1906 (N_1906,N_653,N_440);
xor U1907 (N_1907,N_768,N_868);
nor U1908 (N_1908,N_940,N_661);
or U1909 (N_1909,N_732,N_114);
nand U1910 (N_1910,N_554,N_702);
and U1911 (N_1911,N_328,N_267);
nand U1912 (N_1912,N_491,N_752);
or U1913 (N_1913,N_340,N_938);
nand U1914 (N_1914,N_188,N_101);
or U1915 (N_1915,N_672,N_13);
nand U1916 (N_1916,N_644,N_256);
nor U1917 (N_1917,N_762,N_854);
nor U1918 (N_1918,N_786,N_625);
or U1919 (N_1919,N_442,N_33);
nand U1920 (N_1920,N_34,N_432);
and U1921 (N_1921,N_546,N_131);
or U1922 (N_1922,N_447,N_1);
and U1923 (N_1923,N_492,N_974);
nor U1924 (N_1924,N_540,N_70);
and U1925 (N_1925,N_355,N_300);
or U1926 (N_1926,N_690,N_157);
xor U1927 (N_1927,N_490,N_408);
and U1928 (N_1928,N_185,N_767);
nor U1929 (N_1929,N_116,N_631);
nor U1930 (N_1930,N_276,N_462);
nor U1931 (N_1931,N_661,N_833);
and U1932 (N_1932,N_607,N_956);
or U1933 (N_1933,N_142,N_128);
nor U1934 (N_1934,N_884,N_277);
or U1935 (N_1935,N_38,N_299);
or U1936 (N_1936,N_139,N_733);
and U1937 (N_1937,N_890,N_792);
or U1938 (N_1938,N_20,N_874);
nand U1939 (N_1939,N_836,N_537);
and U1940 (N_1940,N_609,N_483);
nand U1941 (N_1941,N_46,N_23);
and U1942 (N_1942,N_509,N_503);
and U1943 (N_1943,N_577,N_368);
nand U1944 (N_1944,N_229,N_373);
xnor U1945 (N_1945,N_60,N_671);
nand U1946 (N_1946,N_725,N_104);
nor U1947 (N_1947,N_405,N_398);
and U1948 (N_1948,N_281,N_545);
and U1949 (N_1949,N_722,N_346);
and U1950 (N_1950,N_211,N_13);
nor U1951 (N_1951,N_202,N_767);
and U1952 (N_1952,N_308,N_584);
and U1953 (N_1953,N_638,N_154);
or U1954 (N_1954,N_918,N_500);
or U1955 (N_1955,N_876,N_60);
nor U1956 (N_1956,N_263,N_833);
nand U1957 (N_1957,N_971,N_632);
and U1958 (N_1958,N_914,N_26);
or U1959 (N_1959,N_569,N_312);
xnor U1960 (N_1960,N_92,N_525);
or U1961 (N_1961,N_779,N_541);
and U1962 (N_1962,N_116,N_52);
or U1963 (N_1963,N_651,N_772);
or U1964 (N_1964,N_434,N_656);
nand U1965 (N_1965,N_99,N_562);
and U1966 (N_1966,N_613,N_623);
or U1967 (N_1967,N_447,N_948);
xnor U1968 (N_1968,N_535,N_167);
and U1969 (N_1969,N_865,N_754);
and U1970 (N_1970,N_799,N_982);
and U1971 (N_1971,N_205,N_257);
and U1972 (N_1972,N_779,N_531);
nor U1973 (N_1973,N_560,N_447);
xor U1974 (N_1974,N_309,N_492);
and U1975 (N_1975,N_2,N_708);
nor U1976 (N_1976,N_877,N_975);
and U1977 (N_1977,N_916,N_114);
nor U1978 (N_1978,N_490,N_424);
nand U1979 (N_1979,N_3,N_566);
and U1980 (N_1980,N_747,N_655);
and U1981 (N_1981,N_456,N_699);
nand U1982 (N_1982,N_66,N_656);
nor U1983 (N_1983,N_934,N_367);
or U1984 (N_1984,N_671,N_846);
nand U1985 (N_1985,N_833,N_792);
nor U1986 (N_1986,N_447,N_769);
xnor U1987 (N_1987,N_78,N_244);
or U1988 (N_1988,N_926,N_651);
nand U1989 (N_1989,N_185,N_277);
or U1990 (N_1990,N_855,N_817);
nand U1991 (N_1991,N_793,N_159);
xnor U1992 (N_1992,N_222,N_177);
or U1993 (N_1993,N_887,N_337);
xnor U1994 (N_1994,N_516,N_824);
nand U1995 (N_1995,N_519,N_712);
xor U1996 (N_1996,N_43,N_925);
nor U1997 (N_1997,N_301,N_520);
nand U1998 (N_1998,N_393,N_375);
or U1999 (N_1999,N_276,N_2);
xnor U2000 (N_2000,N_1351,N_1434);
nand U2001 (N_2001,N_1643,N_1939);
or U2002 (N_2002,N_1763,N_1052);
and U2003 (N_2003,N_1575,N_1682);
nor U2004 (N_2004,N_1480,N_1704);
xnor U2005 (N_2005,N_1417,N_1166);
nor U2006 (N_2006,N_1927,N_1734);
nand U2007 (N_2007,N_1061,N_1739);
nor U2008 (N_2008,N_1761,N_1104);
or U2009 (N_2009,N_1525,N_1130);
nand U2010 (N_2010,N_1374,N_1644);
xnor U2011 (N_2011,N_1219,N_1147);
and U2012 (N_2012,N_1999,N_1482);
xnor U2013 (N_2013,N_1062,N_1377);
nand U2014 (N_2014,N_1481,N_1199);
or U2015 (N_2015,N_1276,N_1118);
or U2016 (N_2016,N_1093,N_1375);
or U2017 (N_2017,N_1966,N_1212);
nor U2018 (N_2018,N_1263,N_1699);
and U2019 (N_2019,N_1970,N_1047);
xor U2020 (N_2020,N_1688,N_1564);
or U2021 (N_2021,N_1804,N_1720);
or U2022 (N_2022,N_1409,N_1071);
or U2023 (N_2023,N_1940,N_1114);
or U2024 (N_2024,N_1036,N_1043);
and U2025 (N_2025,N_1726,N_1593);
nor U2026 (N_2026,N_1778,N_1233);
nand U2027 (N_2027,N_1509,N_1257);
or U2028 (N_2028,N_1545,N_1703);
nand U2029 (N_2029,N_1444,N_1196);
nor U2030 (N_2030,N_1493,N_1096);
nor U2031 (N_2031,N_1000,N_1568);
and U2032 (N_2032,N_1563,N_1877);
and U2033 (N_2033,N_1412,N_1415);
nor U2034 (N_2034,N_1642,N_1063);
or U2035 (N_2035,N_1401,N_1311);
nor U2036 (N_2036,N_1392,N_1540);
nor U2037 (N_2037,N_1520,N_1458);
nor U2038 (N_2038,N_1471,N_1140);
nor U2039 (N_2039,N_1968,N_1535);
xor U2040 (N_2040,N_1416,N_1156);
or U2041 (N_2041,N_1002,N_1987);
nand U2042 (N_2042,N_1755,N_1078);
and U2043 (N_2043,N_1542,N_1033);
or U2044 (N_2044,N_1132,N_1772);
and U2045 (N_2045,N_1656,N_1406);
or U2046 (N_2046,N_1489,N_1106);
or U2047 (N_2047,N_1089,N_1988);
nor U2048 (N_2048,N_1677,N_1125);
or U2049 (N_2049,N_1760,N_1312);
and U2050 (N_2050,N_1354,N_1991);
or U2051 (N_2051,N_1567,N_1295);
and U2052 (N_2052,N_1165,N_1788);
nand U2053 (N_2053,N_1897,N_1731);
and U2054 (N_2054,N_1916,N_1640);
nand U2055 (N_2055,N_1011,N_1255);
or U2056 (N_2056,N_1866,N_1030);
or U2057 (N_2057,N_1767,N_1967);
xnor U2058 (N_2058,N_1385,N_1997);
xor U2059 (N_2059,N_1014,N_1060);
and U2060 (N_2060,N_1578,N_1422);
and U2061 (N_2061,N_1863,N_1477);
nand U2062 (N_2062,N_1819,N_1019);
xor U2063 (N_2063,N_1608,N_1231);
and U2064 (N_2064,N_1708,N_1474);
or U2065 (N_2065,N_1222,N_1930);
xnor U2066 (N_2066,N_1389,N_1327);
nand U2067 (N_2067,N_1252,N_1102);
nand U2068 (N_2068,N_1020,N_1487);
nand U2069 (N_2069,N_1407,N_1297);
or U2070 (N_2070,N_1645,N_1959);
nor U2071 (N_2071,N_1148,N_1802);
nor U2072 (N_2072,N_1668,N_1712);
nor U2073 (N_2073,N_1825,N_1692);
or U2074 (N_2074,N_1432,N_1789);
nor U2075 (N_2075,N_1037,N_1210);
and U2076 (N_2076,N_1587,N_1594);
and U2077 (N_2077,N_1507,N_1764);
nor U2078 (N_2078,N_1975,N_1439);
or U2079 (N_2079,N_1814,N_1947);
nor U2080 (N_2080,N_1950,N_1485);
and U2081 (N_2081,N_1056,N_1736);
nor U2082 (N_2082,N_1951,N_1119);
nor U2083 (N_2083,N_1003,N_1706);
nand U2084 (N_2084,N_1730,N_1631);
xor U2085 (N_2085,N_1544,N_1678);
nor U2086 (N_2086,N_1470,N_1766);
nand U2087 (N_2087,N_1299,N_1083);
nand U2088 (N_2088,N_1894,N_1486);
xnor U2089 (N_2089,N_1049,N_1710);
nor U2090 (N_2090,N_1261,N_1530);
nor U2091 (N_2091,N_1508,N_1855);
nor U2092 (N_2092,N_1781,N_1356);
and U2093 (N_2093,N_1371,N_1570);
nor U2094 (N_2094,N_1744,N_1289);
nor U2095 (N_2095,N_1346,N_1464);
or U2096 (N_2096,N_1743,N_1473);
and U2097 (N_2097,N_1386,N_1989);
nor U2098 (N_2098,N_1694,N_1634);
and U2099 (N_2099,N_1318,N_1972);
nand U2100 (N_2100,N_1384,N_1438);
nor U2101 (N_2101,N_1903,N_1850);
nor U2102 (N_2102,N_1961,N_1220);
nor U2103 (N_2103,N_1126,N_1752);
and U2104 (N_2104,N_1423,N_1782);
or U2105 (N_2105,N_1807,N_1142);
nor U2106 (N_2106,N_1006,N_1028);
or U2107 (N_2107,N_1316,N_1105);
and U2108 (N_2108,N_1224,N_1902);
nand U2109 (N_2109,N_1214,N_1775);
nor U2110 (N_2110,N_1146,N_1242);
nand U2111 (N_2111,N_1818,N_1057);
and U2112 (N_2112,N_1750,N_1884);
or U2113 (N_2113,N_1552,N_1466);
nand U2114 (N_2114,N_1267,N_1161);
or U2115 (N_2115,N_1264,N_1174);
and U2116 (N_2116,N_1878,N_1762);
or U2117 (N_2117,N_1419,N_1697);
nor U2118 (N_2118,N_1701,N_1141);
nor U2119 (N_2119,N_1094,N_1410);
and U2120 (N_2120,N_1296,N_1601);
and U2121 (N_2121,N_1943,N_1079);
and U2122 (N_2122,N_1537,N_1890);
nor U2123 (N_2123,N_1828,N_1898);
and U2124 (N_2124,N_1483,N_1411);
or U2125 (N_2125,N_1625,N_1728);
and U2126 (N_2126,N_1069,N_1892);
nor U2127 (N_2127,N_1823,N_1149);
or U2128 (N_2128,N_1793,N_1288);
or U2129 (N_2129,N_1499,N_1494);
and U2130 (N_2130,N_1671,N_1247);
nor U2131 (N_2131,N_1433,N_1232);
nor U2132 (N_2132,N_1109,N_1491);
nand U2133 (N_2133,N_1230,N_1662);
or U2134 (N_2134,N_1839,N_1561);
and U2135 (N_2135,N_1176,N_1769);
or U2136 (N_2136,N_1436,N_1500);
nand U2137 (N_2137,N_1050,N_1382);
or U2138 (N_2138,N_1446,N_1364);
and U2139 (N_2139,N_1191,N_1059);
nand U2140 (N_2140,N_1370,N_1867);
nand U2141 (N_2141,N_1541,N_1759);
nand U2142 (N_2142,N_1534,N_1583);
or U2143 (N_2143,N_1580,N_1729);
nand U2144 (N_2144,N_1511,N_1457);
or U2145 (N_2145,N_1572,N_1619);
nor U2146 (N_2146,N_1173,N_1160);
xnor U2147 (N_2147,N_1885,N_1179);
or U2148 (N_2148,N_1463,N_1249);
xnor U2149 (N_2149,N_1691,N_1803);
nand U2150 (N_2150,N_1034,N_1992);
or U2151 (N_2151,N_1503,N_1087);
nor U2152 (N_2152,N_1851,N_1996);
xor U2153 (N_2153,N_1044,N_1323);
nor U2154 (N_2154,N_1963,N_1326);
nand U2155 (N_2155,N_1025,N_1875);
and U2156 (N_2156,N_1531,N_1751);
and U2157 (N_2157,N_1982,N_1287);
nand U2158 (N_2158,N_1195,N_1281);
xnor U2159 (N_2159,N_1426,N_1185);
and U2160 (N_2160,N_1859,N_1820);
nor U2161 (N_2161,N_1824,N_1077);
nor U2162 (N_2162,N_1577,N_1248);
or U2163 (N_2163,N_1722,N_1588);
nand U2164 (N_2164,N_1584,N_1746);
xor U2165 (N_2165,N_1430,N_1971);
or U2166 (N_2166,N_1837,N_1771);
nand U2167 (N_2167,N_1492,N_1277);
and U2168 (N_2168,N_1317,N_1158);
xor U2169 (N_2169,N_1639,N_1742);
or U2170 (N_2170,N_1368,N_1253);
nand U2171 (N_2171,N_1427,N_1053);
or U2172 (N_2172,N_1448,N_1513);
or U2173 (N_2173,N_1424,N_1779);
or U2174 (N_2174,N_1910,N_1546);
and U2175 (N_2175,N_1998,N_1621);
or U2176 (N_2176,N_1893,N_1496);
nor U2177 (N_2177,N_1840,N_1274);
xnor U2178 (N_2178,N_1428,N_1765);
nand U2179 (N_2179,N_1928,N_1139);
nor U2180 (N_2180,N_1238,N_1638);
or U2181 (N_2181,N_1381,N_1361);
or U2182 (N_2182,N_1259,N_1138);
nand U2183 (N_2183,N_1390,N_1012);
nor U2184 (N_2184,N_1957,N_1536);
or U2185 (N_2185,N_1330,N_1573);
and U2186 (N_2186,N_1758,N_1913);
and U2187 (N_2187,N_1075,N_1556);
nand U2188 (N_2188,N_1376,N_1924);
or U2189 (N_2189,N_1889,N_1429);
or U2190 (N_2190,N_1936,N_1243);
nor U2191 (N_2191,N_1021,N_1876);
or U2192 (N_2192,N_1360,N_1908);
nor U2193 (N_2193,N_1955,N_1647);
or U2194 (N_2194,N_1977,N_1123);
or U2195 (N_2195,N_1522,N_1711);
and U2196 (N_2196,N_1891,N_1113);
nor U2197 (N_2197,N_1954,N_1091);
nor U2198 (N_2198,N_1845,N_1282);
xor U2199 (N_2199,N_1945,N_1349);
nand U2200 (N_2200,N_1533,N_1838);
or U2201 (N_2201,N_1651,N_1465);
nand U2202 (N_2202,N_1452,N_1357);
nor U2203 (N_2203,N_1635,N_1134);
xor U2204 (N_2204,N_1286,N_1100);
xnor U2205 (N_2205,N_1843,N_1153);
nand U2206 (N_2206,N_1912,N_1420);
and U2207 (N_2207,N_1168,N_1571);
or U2208 (N_2208,N_1421,N_1298);
nor U2209 (N_2209,N_1596,N_1732);
nand U2210 (N_2210,N_1239,N_1488);
and U2211 (N_2211,N_1240,N_1822);
nor U2212 (N_2212,N_1476,N_1607);
and U2213 (N_2213,N_1154,N_1948);
and U2214 (N_2214,N_1919,N_1344);
nor U2215 (N_2215,N_1209,N_1502);
and U2216 (N_2216,N_1402,N_1292);
nor U2217 (N_2217,N_1099,N_1235);
and U2218 (N_2218,N_1676,N_1151);
and U2219 (N_2219,N_1768,N_1347);
nand U2220 (N_2220,N_1358,N_1633);
or U2221 (N_2221,N_1610,N_1715);
xnor U2222 (N_2222,N_1684,N_1886);
and U2223 (N_2223,N_1952,N_1911);
or U2224 (N_2224,N_1887,N_1440);
and U2225 (N_2225,N_1169,N_1092);
or U2226 (N_2226,N_1953,N_1205);
or U2227 (N_2227,N_1705,N_1674);
xnor U2228 (N_2228,N_1641,N_1042);
nor U2229 (N_2229,N_1110,N_1117);
nand U2230 (N_2230,N_1709,N_1521);
nor U2231 (N_2231,N_1456,N_1009);
or U2232 (N_2232,N_1265,N_1367);
and U2233 (N_2233,N_1505,N_1048);
xnor U2234 (N_2234,N_1504,N_1532);
or U2235 (N_2235,N_1574,N_1909);
and U2236 (N_2236,N_1800,N_1278);
nand U2237 (N_2237,N_1453,N_1150);
or U2238 (N_2238,N_1806,N_1359);
or U2239 (N_2239,N_1801,N_1182);
or U2240 (N_2240,N_1405,N_1455);
nand U2241 (N_2241,N_1717,N_1167);
nand U2242 (N_2242,N_1103,N_1501);
or U2243 (N_2243,N_1241,N_1915);
nor U2244 (N_2244,N_1698,N_1334);
or U2245 (N_2245,N_1589,N_1581);
nand U2246 (N_2246,N_1713,N_1554);
xor U2247 (N_2247,N_1308,N_1721);
and U2248 (N_2248,N_1549,N_1256);
nand U2249 (N_2249,N_1208,N_1171);
and U2250 (N_2250,N_1081,N_1314);
xor U2251 (N_2251,N_1177,N_1135);
nor U2252 (N_2252,N_1462,N_1695);
nand U2253 (N_2253,N_1881,N_1350);
or U2254 (N_2254,N_1780,N_1074);
or U2255 (N_2255,N_1690,N_1181);
or U2256 (N_2256,N_1922,N_1475);
or U2257 (N_2257,N_1551,N_1319);
and U2258 (N_2258,N_1076,N_1321);
nor U2259 (N_2259,N_1686,N_1627);
xor U2260 (N_2260,N_1115,N_1652);
nor U2261 (N_2261,N_1648,N_1526);
and U2262 (N_2262,N_1159,N_1741);
nand U2263 (N_2263,N_1379,N_1022);
xor U2264 (N_2264,N_1260,N_1234);
xor U2265 (N_2265,N_1279,N_1178);
and U2266 (N_2266,N_1335,N_1300);
or U2267 (N_2267,N_1032,N_1495);
nor U2268 (N_2268,N_1904,N_1221);
nor U2269 (N_2269,N_1309,N_1670);
nor U2270 (N_2270,N_1962,N_1320);
nor U2271 (N_2271,N_1155,N_1632);
and U2272 (N_2272,N_1005,N_1403);
nand U2273 (N_2273,N_1776,N_1200);
nor U2274 (N_2274,N_1152,N_1007);
nor U2275 (N_2275,N_1228,N_1796);
and U2276 (N_2276,N_1990,N_1414);
or U2277 (N_2277,N_1849,N_1273);
nand U2278 (N_2278,N_1128,N_1121);
nor U2279 (N_2279,N_1524,N_1258);
and U2280 (N_2280,N_1562,N_1733);
or U2281 (N_2281,N_1122,N_1979);
nand U2282 (N_2282,N_1101,N_1301);
and U2283 (N_2283,N_1934,N_1754);
nand U2284 (N_2284,N_1284,N_1815);
or U2285 (N_2285,N_1027,N_1586);
or U2286 (N_2286,N_1757,N_1856);
nor U2287 (N_2287,N_1935,N_1095);
or U2288 (N_2288,N_1180,N_1696);
nor U2289 (N_2289,N_1517,N_1418);
and U2290 (N_2290,N_1844,N_1058);
nand U2291 (N_2291,N_1790,N_1941);
nor U2292 (N_2292,N_1797,N_1826);
nand U2293 (N_2293,N_1204,N_1745);
nor U2294 (N_2294,N_1938,N_1226);
and U2295 (N_2295,N_1506,N_1127);
nand U2296 (N_2296,N_1097,N_1229);
and U2297 (N_2297,N_1468,N_1748);
nor U2298 (N_2298,N_1557,N_1604);
nand U2299 (N_2299,N_1262,N_1786);
or U2300 (N_2300,N_1834,N_1649);
and U2301 (N_2301,N_1896,N_1207);
xor U2302 (N_2302,N_1770,N_1162);
xor U2303 (N_2303,N_1833,N_1591);
nand U2304 (N_2304,N_1805,N_1969);
nor U2305 (N_2305,N_1777,N_1821);
and U2306 (N_2306,N_1342,N_1792);
or U2307 (N_2307,N_1467,N_1667);
nor U2308 (N_2308,N_1842,N_1917);
nor U2309 (N_2309,N_1340,N_1787);
and U2310 (N_2310,N_1868,N_1206);
nor U2311 (N_2311,N_1082,N_1088);
or U2312 (N_2312,N_1213,N_1313);
nor U2313 (N_2313,N_1628,N_1490);
and U2314 (N_2314,N_1211,N_1548);
or U2315 (N_2315,N_1993,N_1186);
and U2316 (N_2316,N_1227,N_1809);
or U2317 (N_2317,N_1223,N_1447);
xnor U2318 (N_2318,N_1072,N_1599);
or U2319 (N_2319,N_1519,N_1846);
or U2320 (N_2320,N_1035,N_1615);
nor U2321 (N_2321,N_1516,N_1514);
or U2322 (N_2322,N_1654,N_1164);
and U2323 (N_2323,N_1306,N_1873);
nor U2324 (N_2324,N_1983,N_1280);
nor U2325 (N_2325,N_1408,N_1756);
and U2326 (N_2326,N_1921,N_1960);
or U2327 (N_2327,N_1646,N_1973);
nand U2328 (N_2328,N_1184,N_1304);
and U2329 (N_2329,N_1808,N_1858);
nand U2330 (N_2330,N_1799,N_1080);
or U2331 (N_2331,N_1051,N_1600);
and U2332 (N_2332,N_1008,N_1550);
or U2333 (N_2333,N_1847,N_1933);
and U2334 (N_2334,N_1529,N_1920);
or U2335 (N_2335,N_1626,N_1046);
or U2336 (N_2336,N_1145,N_1900);
and U2337 (N_2337,N_1454,N_1813);
and U2338 (N_2338,N_1395,N_1559);
nand U2339 (N_2339,N_1986,N_1425);
xor U2340 (N_2340,N_1740,N_1926);
or U2341 (N_2341,N_1882,N_1435);
and U2342 (N_2342,N_1624,N_1623);
and U2343 (N_2343,N_1795,N_1283);
nor U2344 (N_2344,N_1041,N_1579);
nand U2345 (N_2345,N_1380,N_1747);
nand U2346 (N_2346,N_1985,N_1108);
or U2347 (N_2347,N_1665,N_1391);
or U2348 (N_2348,N_1268,N_1017);
and U2349 (N_2349,N_1333,N_1659);
xor U2350 (N_2350,N_1637,N_1098);
or U2351 (N_2351,N_1461,N_1484);
xor U2352 (N_2352,N_1023,N_1131);
nor U2353 (N_2353,N_1661,N_1669);
xnor U2354 (N_2354,N_1218,N_1291);
or U2355 (N_2355,N_1216,N_1899);
and U2356 (N_2356,N_1653,N_1538);
or U2357 (N_2357,N_1905,N_1609);
and U2358 (N_2358,N_1090,N_1066);
and U2359 (N_2359,N_1879,N_1817);
or U2360 (N_2360,N_1413,N_1613);
nand U2361 (N_2361,N_1681,N_1236);
nor U2362 (N_2362,N_1816,N_1658);
nor U2363 (N_2363,N_1539,N_1266);
xor U2364 (N_2364,N_1459,N_1183);
or U2365 (N_2365,N_1137,N_1718);
and U2366 (N_2366,N_1657,N_1029);
nor U2367 (N_2367,N_1614,N_1666);
or U2368 (N_2368,N_1322,N_1918);
and U2369 (N_2369,N_1112,N_1124);
nor U2370 (N_2370,N_1869,N_1472);
nand U2371 (N_2371,N_1590,N_1272);
and U2372 (N_2372,N_1620,N_1946);
or U2373 (N_2373,N_1172,N_1175);
and U2374 (N_2374,N_1244,N_1315);
nor U2375 (N_2375,N_1965,N_1341);
nor U2376 (N_2376,N_1373,N_1064);
nor U2377 (N_2377,N_1664,N_1864);
xnor U2378 (N_2378,N_1518,N_1016);
or U2379 (N_2379,N_1784,N_1136);
nor U2380 (N_2380,N_1725,N_1964);
nor U2381 (N_2381,N_1498,N_1679);
xor U2382 (N_2382,N_1974,N_1451);
xor U2383 (N_2383,N_1874,N_1566);
or U2384 (N_2384,N_1857,N_1655);
xnor U2385 (N_2385,N_1460,N_1880);
or U2386 (N_2386,N_1618,N_1325);
nand U2387 (N_2387,N_1958,N_1680);
xnor U2388 (N_2388,N_1054,N_1190);
nand U2389 (N_2389,N_1853,N_1835);
and U2390 (N_2390,N_1687,N_1449);
nand U2391 (N_2391,N_1290,N_1307);
nor U2392 (N_2392,N_1442,N_1067);
nand U2393 (N_2393,N_1378,N_1497);
nor U2394 (N_2394,N_1478,N_1724);
and U2395 (N_2395,N_1217,N_1189);
and U2396 (N_2396,N_1170,N_1931);
nor U2397 (N_2397,N_1783,N_1305);
or U2398 (N_2398,N_1038,N_1394);
and U2399 (N_2399,N_1039,N_1883);
and U2400 (N_2400,N_1337,N_1848);
xor U2401 (N_2401,N_1569,N_1716);
xor U2402 (N_2402,N_1107,N_1026);
and U2403 (N_2403,N_1794,N_1942);
and U2404 (N_2404,N_1250,N_1595);
or U2405 (N_2405,N_1749,N_1831);
and U2406 (N_2406,N_1675,N_1443);
xor U2407 (N_2407,N_1558,N_1157);
or U2408 (N_2408,N_1672,N_1854);
or U2409 (N_2409,N_1907,N_1201);
or U2410 (N_2410,N_1302,N_1479);
nor U2411 (N_2411,N_1888,N_1193);
or U2412 (N_2412,N_1348,N_1663);
nor U2413 (N_2413,N_1332,N_1198);
xnor U2414 (N_2414,N_1555,N_1811);
xnor U2415 (N_2415,N_1270,N_1861);
and U2416 (N_2416,N_1396,N_1338);
nor U2417 (N_2417,N_1294,N_1441);
or U2418 (N_2418,N_1871,N_1387);
and U2419 (N_2419,N_1753,N_1031);
nand U2420 (N_2420,N_1133,N_1269);
or U2421 (N_2421,N_1116,N_1660);
nand U2422 (N_2422,N_1310,N_1202);
nor U2423 (N_2423,N_1707,N_1515);
nand U2424 (N_2424,N_1445,N_1245);
and U2425 (N_2425,N_1324,N_1995);
or U2426 (N_2426,N_1120,N_1702);
nor U2427 (N_2427,N_1984,N_1719);
or U2428 (N_2428,N_1275,N_1363);
nor U2429 (N_2429,N_1527,N_1872);
xor U2430 (N_2430,N_1582,N_1832);
and U2431 (N_2431,N_1810,N_1388);
or U2432 (N_2432,N_1215,N_1331);
nand U2433 (N_2433,N_1895,N_1914);
or U2434 (N_2434,N_1812,N_1937);
nor U2435 (N_2435,N_1285,N_1024);
nand U2436 (N_2436,N_1192,N_1689);
or U2437 (N_2437,N_1612,N_1365);
or U2438 (N_2438,N_1978,N_1785);
nor U2439 (N_2439,N_1956,N_1045);
nand U2440 (N_2440,N_1981,N_1700);
and U2441 (N_2441,N_1976,N_1343);
and U2442 (N_2442,N_1798,N_1606);
nand U2443 (N_2443,N_1598,N_1355);
nand U2444 (N_2444,N_1372,N_1870);
or U2445 (N_2445,N_1329,N_1068);
nor U2446 (N_2446,N_1328,N_1018);
or U2447 (N_2447,N_1163,N_1237);
and U2448 (N_2448,N_1723,N_1791);
and U2449 (N_2449,N_1543,N_1271);
and U2450 (N_2450,N_1070,N_1143);
or U2451 (N_2451,N_1949,N_1714);
xnor U2452 (N_2452,N_1013,N_1010);
and U2453 (N_2453,N_1862,N_1188);
xnor U2454 (N_2454,N_1065,N_1592);
nor U2455 (N_2455,N_1576,N_1693);
xnor U2456 (N_2456,N_1437,N_1774);
nand U2457 (N_2457,N_1040,N_1560);
and U2458 (N_2458,N_1523,N_1553);
and U2459 (N_2459,N_1225,N_1830);
or U2460 (N_2460,N_1431,N_1393);
nand U2461 (N_2461,N_1929,N_1510);
nor U2462 (N_2462,N_1398,N_1085);
xor U2463 (N_2463,N_1400,N_1727);
or U2464 (N_2464,N_1293,N_1512);
or U2465 (N_2465,N_1353,N_1547);
and U2466 (N_2466,N_1629,N_1829);
xor U2467 (N_2467,N_1925,N_1111);
xnor U2468 (N_2468,N_1397,N_1383);
nor U2469 (N_2469,N_1683,N_1565);
and U2470 (N_2470,N_1336,N_1673);
nand U2471 (N_2471,N_1611,N_1605);
nand U2472 (N_2472,N_1585,N_1366);
nor U2473 (N_2473,N_1836,N_1622);
nand U2474 (N_2474,N_1251,N_1944);
xnor U2475 (N_2475,N_1203,N_1685);
and U2476 (N_2476,N_1630,N_1015);
and U2477 (N_2477,N_1738,N_1352);
or U2478 (N_2478,N_1339,N_1303);
or U2479 (N_2479,N_1735,N_1650);
nor U2480 (N_2480,N_1450,N_1254);
or U2481 (N_2481,N_1737,N_1345);
nand U2482 (N_2482,N_1194,N_1636);
nor U2483 (N_2483,N_1246,N_1469);
nand U2484 (N_2484,N_1144,N_1932);
nor U2485 (N_2485,N_1086,N_1369);
xnor U2486 (N_2486,N_1980,N_1404);
nor U2487 (N_2487,N_1906,N_1001);
nand U2488 (N_2488,N_1129,N_1865);
nand U2489 (N_2489,N_1860,N_1187);
and U2490 (N_2490,N_1773,N_1004);
and U2491 (N_2491,N_1852,N_1084);
xor U2492 (N_2492,N_1616,N_1827);
nand U2493 (N_2493,N_1841,N_1603);
nand U2494 (N_2494,N_1901,N_1055);
or U2495 (N_2495,N_1923,N_1362);
nor U2496 (N_2496,N_1617,N_1073);
nand U2497 (N_2497,N_1528,N_1602);
and U2498 (N_2498,N_1994,N_1399);
or U2499 (N_2499,N_1597,N_1197);
nand U2500 (N_2500,N_1337,N_1353);
xnor U2501 (N_2501,N_1365,N_1267);
nor U2502 (N_2502,N_1532,N_1077);
nand U2503 (N_2503,N_1276,N_1163);
or U2504 (N_2504,N_1958,N_1686);
or U2505 (N_2505,N_1012,N_1402);
and U2506 (N_2506,N_1448,N_1841);
or U2507 (N_2507,N_1821,N_1325);
xor U2508 (N_2508,N_1010,N_1810);
and U2509 (N_2509,N_1417,N_1256);
or U2510 (N_2510,N_1278,N_1406);
or U2511 (N_2511,N_1544,N_1808);
nor U2512 (N_2512,N_1739,N_1466);
nor U2513 (N_2513,N_1001,N_1871);
or U2514 (N_2514,N_1839,N_1409);
and U2515 (N_2515,N_1865,N_1803);
nor U2516 (N_2516,N_1997,N_1502);
xor U2517 (N_2517,N_1138,N_1217);
or U2518 (N_2518,N_1947,N_1063);
nor U2519 (N_2519,N_1020,N_1262);
or U2520 (N_2520,N_1228,N_1295);
or U2521 (N_2521,N_1818,N_1659);
nor U2522 (N_2522,N_1438,N_1005);
nor U2523 (N_2523,N_1312,N_1904);
xnor U2524 (N_2524,N_1303,N_1201);
nand U2525 (N_2525,N_1564,N_1044);
nand U2526 (N_2526,N_1834,N_1419);
and U2527 (N_2527,N_1866,N_1096);
nor U2528 (N_2528,N_1629,N_1546);
nor U2529 (N_2529,N_1784,N_1231);
nand U2530 (N_2530,N_1173,N_1028);
or U2531 (N_2531,N_1583,N_1268);
or U2532 (N_2532,N_1372,N_1700);
nand U2533 (N_2533,N_1394,N_1549);
nand U2534 (N_2534,N_1759,N_1312);
nand U2535 (N_2535,N_1024,N_1684);
and U2536 (N_2536,N_1643,N_1613);
nor U2537 (N_2537,N_1648,N_1382);
or U2538 (N_2538,N_1864,N_1137);
xnor U2539 (N_2539,N_1349,N_1698);
and U2540 (N_2540,N_1065,N_1633);
and U2541 (N_2541,N_1375,N_1089);
nor U2542 (N_2542,N_1109,N_1811);
xnor U2543 (N_2543,N_1369,N_1634);
nor U2544 (N_2544,N_1228,N_1694);
and U2545 (N_2545,N_1882,N_1599);
and U2546 (N_2546,N_1023,N_1143);
nand U2547 (N_2547,N_1992,N_1763);
xnor U2548 (N_2548,N_1361,N_1139);
nor U2549 (N_2549,N_1812,N_1387);
or U2550 (N_2550,N_1902,N_1663);
nand U2551 (N_2551,N_1729,N_1550);
nor U2552 (N_2552,N_1475,N_1683);
or U2553 (N_2553,N_1429,N_1630);
and U2554 (N_2554,N_1065,N_1366);
or U2555 (N_2555,N_1750,N_1549);
nand U2556 (N_2556,N_1295,N_1866);
or U2557 (N_2557,N_1274,N_1773);
nand U2558 (N_2558,N_1459,N_1538);
or U2559 (N_2559,N_1887,N_1356);
or U2560 (N_2560,N_1269,N_1385);
nor U2561 (N_2561,N_1955,N_1594);
or U2562 (N_2562,N_1949,N_1673);
nand U2563 (N_2563,N_1346,N_1399);
and U2564 (N_2564,N_1914,N_1330);
nor U2565 (N_2565,N_1566,N_1935);
nand U2566 (N_2566,N_1875,N_1739);
nand U2567 (N_2567,N_1730,N_1526);
nor U2568 (N_2568,N_1937,N_1899);
and U2569 (N_2569,N_1290,N_1596);
or U2570 (N_2570,N_1760,N_1766);
or U2571 (N_2571,N_1766,N_1770);
nor U2572 (N_2572,N_1581,N_1845);
nand U2573 (N_2573,N_1389,N_1402);
and U2574 (N_2574,N_1577,N_1735);
nor U2575 (N_2575,N_1248,N_1213);
and U2576 (N_2576,N_1779,N_1097);
and U2577 (N_2577,N_1032,N_1097);
nor U2578 (N_2578,N_1687,N_1074);
nor U2579 (N_2579,N_1960,N_1947);
or U2580 (N_2580,N_1809,N_1549);
nand U2581 (N_2581,N_1393,N_1512);
and U2582 (N_2582,N_1369,N_1884);
and U2583 (N_2583,N_1176,N_1473);
and U2584 (N_2584,N_1550,N_1356);
nand U2585 (N_2585,N_1757,N_1879);
or U2586 (N_2586,N_1320,N_1647);
or U2587 (N_2587,N_1665,N_1498);
and U2588 (N_2588,N_1811,N_1455);
nor U2589 (N_2589,N_1190,N_1604);
nor U2590 (N_2590,N_1383,N_1065);
nor U2591 (N_2591,N_1535,N_1928);
or U2592 (N_2592,N_1323,N_1837);
nand U2593 (N_2593,N_1270,N_1994);
nor U2594 (N_2594,N_1942,N_1725);
or U2595 (N_2595,N_1396,N_1352);
nand U2596 (N_2596,N_1916,N_1917);
or U2597 (N_2597,N_1612,N_1194);
or U2598 (N_2598,N_1351,N_1608);
and U2599 (N_2599,N_1804,N_1769);
nand U2600 (N_2600,N_1356,N_1771);
nand U2601 (N_2601,N_1060,N_1921);
nor U2602 (N_2602,N_1687,N_1407);
nor U2603 (N_2603,N_1775,N_1878);
nor U2604 (N_2604,N_1852,N_1306);
nand U2605 (N_2605,N_1882,N_1369);
nand U2606 (N_2606,N_1394,N_1790);
and U2607 (N_2607,N_1329,N_1793);
and U2608 (N_2608,N_1206,N_1002);
and U2609 (N_2609,N_1652,N_1271);
nand U2610 (N_2610,N_1728,N_1470);
nand U2611 (N_2611,N_1300,N_1001);
and U2612 (N_2612,N_1501,N_1905);
or U2613 (N_2613,N_1591,N_1155);
and U2614 (N_2614,N_1523,N_1583);
nand U2615 (N_2615,N_1820,N_1325);
or U2616 (N_2616,N_1783,N_1428);
and U2617 (N_2617,N_1154,N_1720);
or U2618 (N_2618,N_1809,N_1339);
nor U2619 (N_2619,N_1570,N_1524);
nor U2620 (N_2620,N_1082,N_1735);
and U2621 (N_2621,N_1120,N_1282);
and U2622 (N_2622,N_1295,N_1380);
nand U2623 (N_2623,N_1624,N_1107);
nand U2624 (N_2624,N_1231,N_1631);
nor U2625 (N_2625,N_1210,N_1661);
or U2626 (N_2626,N_1013,N_1592);
or U2627 (N_2627,N_1679,N_1875);
nand U2628 (N_2628,N_1658,N_1019);
and U2629 (N_2629,N_1912,N_1280);
and U2630 (N_2630,N_1054,N_1607);
nor U2631 (N_2631,N_1193,N_1551);
nor U2632 (N_2632,N_1414,N_1885);
xnor U2633 (N_2633,N_1587,N_1449);
or U2634 (N_2634,N_1447,N_1561);
or U2635 (N_2635,N_1365,N_1751);
and U2636 (N_2636,N_1864,N_1855);
and U2637 (N_2637,N_1309,N_1440);
nor U2638 (N_2638,N_1751,N_1781);
nor U2639 (N_2639,N_1254,N_1138);
nor U2640 (N_2640,N_1765,N_1850);
or U2641 (N_2641,N_1629,N_1404);
and U2642 (N_2642,N_1619,N_1017);
or U2643 (N_2643,N_1499,N_1416);
xnor U2644 (N_2644,N_1860,N_1618);
xnor U2645 (N_2645,N_1884,N_1283);
xnor U2646 (N_2646,N_1782,N_1854);
nor U2647 (N_2647,N_1972,N_1223);
nand U2648 (N_2648,N_1587,N_1283);
nor U2649 (N_2649,N_1178,N_1200);
xnor U2650 (N_2650,N_1648,N_1946);
and U2651 (N_2651,N_1366,N_1608);
or U2652 (N_2652,N_1925,N_1943);
nand U2653 (N_2653,N_1966,N_1078);
or U2654 (N_2654,N_1195,N_1425);
and U2655 (N_2655,N_1143,N_1898);
and U2656 (N_2656,N_1901,N_1758);
and U2657 (N_2657,N_1959,N_1614);
and U2658 (N_2658,N_1660,N_1622);
or U2659 (N_2659,N_1643,N_1029);
or U2660 (N_2660,N_1666,N_1770);
nand U2661 (N_2661,N_1666,N_1305);
and U2662 (N_2662,N_1825,N_1497);
nor U2663 (N_2663,N_1896,N_1254);
nand U2664 (N_2664,N_1944,N_1903);
nor U2665 (N_2665,N_1845,N_1922);
and U2666 (N_2666,N_1574,N_1845);
xnor U2667 (N_2667,N_1771,N_1479);
xnor U2668 (N_2668,N_1598,N_1132);
nor U2669 (N_2669,N_1494,N_1448);
xor U2670 (N_2670,N_1204,N_1991);
nand U2671 (N_2671,N_1706,N_1046);
xor U2672 (N_2672,N_1565,N_1413);
or U2673 (N_2673,N_1492,N_1642);
xnor U2674 (N_2674,N_1881,N_1647);
nor U2675 (N_2675,N_1107,N_1717);
and U2676 (N_2676,N_1693,N_1294);
nor U2677 (N_2677,N_1045,N_1649);
xnor U2678 (N_2678,N_1363,N_1572);
nand U2679 (N_2679,N_1781,N_1230);
and U2680 (N_2680,N_1759,N_1470);
and U2681 (N_2681,N_1445,N_1076);
and U2682 (N_2682,N_1723,N_1838);
or U2683 (N_2683,N_1699,N_1032);
nor U2684 (N_2684,N_1794,N_1584);
or U2685 (N_2685,N_1914,N_1277);
and U2686 (N_2686,N_1500,N_1208);
nand U2687 (N_2687,N_1947,N_1363);
xor U2688 (N_2688,N_1731,N_1368);
and U2689 (N_2689,N_1778,N_1090);
nor U2690 (N_2690,N_1882,N_1571);
or U2691 (N_2691,N_1552,N_1835);
and U2692 (N_2692,N_1124,N_1839);
nand U2693 (N_2693,N_1163,N_1288);
nor U2694 (N_2694,N_1538,N_1991);
xnor U2695 (N_2695,N_1274,N_1813);
nor U2696 (N_2696,N_1450,N_1617);
nor U2697 (N_2697,N_1091,N_1785);
xnor U2698 (N_2698,N_1896,N_1579);
nor U2699 (N_2699,N_1851,N_1292);
nand U2700 (N_2700,N_1668,N_1293);
nand U2701 (N_2701,N_1894,N_1572);
nor U2702 (N_2702,N_1810,N_1950);
nand U2703 (N_2703,N_1963,N_1405);
nand U2704 (N_2704,N_1138,N_1040);
nand U2705 (N_2705,N_1435,N_1520);
nor U2706 (N_2706,N_1759,N_1136);
or U2707 (N_2707,N_1173,N_1753);
or U2708 (N_2708,N_1160,N_1075);
or U2709 (N_2709,N_1483,N_1351);
or U2710 (N_2710,N_1132,N_1749);
or U2711 (N_2711,N_1234,N_1663);
or U2712 (N_2712,N_1152,N_1333);
or U2713 (N_2713,N_1051,N_1127);
or U2714 (N_2714,N_1823,N_1566);
and U2715 (N_2715,N_1405,N_1793);
nor U2716 (N_2716,N_1042,N_1446);
nor U2717 (N_2717,N_1952,N_1565);
nor U2718 (N_2718,N_1714,N_1195);
nand U2719 (N_2719,N_1906,N_1654);
or U2720 (N_2720,N_1255,N_1472);
nand U2721 (N_2721,N_1078,N_1371);
nor U2722 (N_2722,N_1711,N_1692);
xor U2723 (N_2723,N_1497,N_1437);
or U2724 (N_2724,N_1841,N_1611);
nand U2725 (N_2725,N_1709,N_1253);
or U2726 (N_2726,N_1962,N_1398);
or U2727 (N_2727,N_1464,N_1393);
xor U2728 (N_2728,N_1468,N_1178);
xnor U2729 (N_2729,N_1529,N_1030);
and U2730 (N_2730,N_1227,N_1703);
or U2731 (N_2731,N_1444,N_1796);
nand U2732 (N_2732,N_1579,N_1455);
nor U2733 (N_2733,N_1225,N_1368);
and U2734 (N_2734,N_1755,N_1838);
nor U2735 (N_2735,N_1839,N_1958);
or U2736 (N_2736,N_1428,N_1940);
or U2737 (N_2737,N_1953,N_1891);
nand U2738 (N_2738,N_1735,N_1818);
nor U2739 (N_2739,N_1680,N_1506);
and U2740 (N_2740,N_1332,N_1666);
and U2741 (N_2741,N_1495,N_1672);
nand U2742 (N_2742,N_1315,N_1418);
nand U2743 (N_2743,N_1012,N_1510);
xor U2744 (N_2744,N_1722,N_1939);
xor U2745 (N_2745,N_1216,N_1496);
nand U2746 (N_2746,N_1541,N_1192);
or U2747 (N_2747,N_1460,N_1629);
xnor U2748 (N_2748,N_1116,N_1065);
and U2749 (N_2749,N_1760,N_1389);
and U2750 (N_2750,N_1078,N_1181);
nor U2751 (N_2751,N_1843,N_1128);
and U2752 (N_2752,N_1632,N_1174);
nor U2753 (N_2753,N_1811,N_1882);
and U2754 (N_2754,N_1458,N_1350);
nor U2755 (N_2755,N_1064,N_1843);
xnor U2756 (N_2756,N_1011,N_1097);
nor U2757 (N_2757,N_1009,N_1938);
and U2758 (N_2758,N_1466,N_1647);
and U2759 (N_2759,N_1619,N_1604);
nor U2760 (N_2760,N_1772,N_1636);
and U2761 (N_2761,N_1547,N_1845);
nor U2762 (N_2762,N_1279,N_1469);
or U2763 (N_2763,N_1000,N_1751);
or U2764 (N_2764,N_1503,N_1133);
nor U2765 (N_2765,N_1497,N_1984);
or U2766 (N_2766,N_1052,N_1271);
xnor U2767 (N_2767,N_1207,N_1046);
nor U2768 (N_2768,N_1408,N_1751);
nand U2769 (N_2769,N_1595,N_1266);
and U2770 (N_2770,N_1578,N_1055);
nand U2771 (N_2771,N_1259,N_1847);
or U2772 (N_2772,N_1254,N_1194);
nand U2773 (N_2773,N_1297,N_1483);
nor U2774 (N_2774,N_1889,N_1709);
nor U2775 (N_2775,N_1150,N_1128);
nor U2776 (N_2776,N_1881,N_1905);
nor U2777 (N_2777,N_1581,N_1202);
nor U2778 (N_2778,N_1164,N_1336);
or U2779 (N_2779,N_1990,N_1808);
nand U2780 (N_2780,N_1098,N_1977);
nand U2781 (N_2781,N_1234,N_1150);
nand U2782 (N_2782,N_1534,N_1489);
nand U2783 (N_2783,N_1909,N_1885);
nand U2784 (N_2784,N_1733,N_1096);
xor U2785 (N_2785,N_1615,N_1387);
or U2786 (N_2786,N_1532,N_1146);
nand U2787 (N_2787,N_1653,N_1119);
nand U2788 (N_2788,N_1774,N_1724);
nor U2789 (N_2789,N_1142,N_1853);
xor U2790 (N_2790,N_1198,N_1564);
and U2791 (N_2791,N_1366,N_1171);
nor U2792 (N_2792,N_1064,N_1975);
or U2793 (N_2793,N_1920,N_1351);
nand U2794 (N_2794,N_1962,N_1637);
nand U2795 (N_2795,N_1841,N_1139);
nor U2796 (N_2796,N_1388,N_1175);
nand U2797 (N_2797,N_1007,N_1445);
and U2798 (N_2798,N_1366,N_1637);
and U2799 (N_2799,N_1830,N_1260);
nand U2800 (N_2800,N_1542,N_1652);
nor U2801 (N_2801,N_1607,N_1783);
nand U2802 (N_2802,N_1568,N_1265);
nand U2803 (N_2803,N_1478,N_1562);
nor U2804 (N_2804,N_1112,N_1184);
nand U2805 (N_2805,N_1110,N_1071);
xor U2806 (N_2806,N_1999,N_1017);
or U2807 (N_2807,N_1741,N_1639);
nand U2808 (N_2808,N_1749,N_1641);
or U2809 (N_2809,N_1021,N_1119);
nor U2810 (N_2810,N_1988,N_1299);
and U2811 (N_2811,N_1814,N_1247);
or U2812 (N_2812,N_1034,N_1293);
and U2813 (N_2813,N_1732,N_1953);
and U2814 (N_2814,N_1093,N_1457);
and U2815 (N_2815,N_1412,N_1555);
or U2816 (N_2816,N_1613,N_1009);
xor U2817 (N_2817,N_1971,N_1676);
nor U2818 (N_2818,N_1578,N_1127);
nand U2819 (N_2819,N_1374,N_1632);
nor U2820 (N_2820,N_1580,N_1397);
or U2821 (N_2821,N_1629,N_1262);
nand U2822 (N_2822,N_1554,N_1724);
or U2823 (N_2823,N_1070,N_1013);
nand U2824 (N_2824,N_1629,N_1470);
or U2825 (N_2825,N_1417,N_1013);
or U2826 (N_2826,N_1031,N_1737);
and U2827 (N_2827,N_1823,N_1435);
xnor U2828 (N_2828,N_1090,N_1509);
nand U2829 (N_2829,N_1380,N_1767);
nand U2830 (N_2830,N_1610,N_1862);
xor U2831 (N_2831,N_1754,N_1376);
or U2832 (N_2832,N_1908,N_1203);
nor U2833 (N_2833,N_1040,N_1132);
or U2834 (N_2834,N_1751,N_1312);
nor U2835 (N_2835,N_1614,N_1258);
or U2836 (N_2836,N_1589,N_1893);
nor U2837 (N_2837,N_1695,N_1598);
and U2838 (N_2838,N_1851,N_1863);
and U2839 (N_2839,N_1148,N_1650);
nor U2840 (N_2840,N_1042,N_1583);
xor U2841 (N_2841,N_1648,N_1576);
nor U2842 (N_2842,N_1142,N_1255);
nor U2843 (N_2843,N_1087,N_1068);
nand U2844 (N_2844,N_1216,N_1053);
and U2845 (N_2845,N_1240,N_1285);
or U2846 (N_2846,N_1739,N_1740);
and U2847 (N_2847,N_1190,N_1669);
or U2848 (N_2848,N_1543,N_1612);
nand U2849 (N_2849,N_1673,N_1388);
xor U2850 (N_2850,N_1556,N_1238);
xor U2851 (N_2851,N_1511,N_1736);
and U2852 (N_2852,N_1077,N_1827);
nand U2853 (N_2853,N_1695,N_1071);
and U2854 (N_2854,N_1125,N_1958);
and U2855 (N_2855,N_1892,N_1765);
or U2856 (N_2856,N_1374,N_1194);
nor U2857 (N_2857,N_1750,N_1031);
nand U2858 (N_2858,N_1558,N_1110);
xor U2859 (N_2859,N_1367,N_1644);
nor U2860 (N_2860,N_1657,N_1638);
nor U2861 (N_2861,N_1786,N_1057);
and U2862 (N_2862,N_1319,N_1288);
nor U2863 (N_2863,N_1534,N_1956);
nor U2864 (N_2864,N_1305,N_1887);
and U2865 (N_2865,N_1475,N_1148);
and U2866 (N_2866,N_1129,N_1692);
nor U2867 (N_2867,N_1115,N_1714);
nand U2868 (N_2868,N_1399,N_1591);
nor U2869 (N_2869,N_1314,N_1527);
or U2870 (N_2870,N_1829,N_1999);
and U2871 (N_2871,N_1766,N_1208);
and U2872 (N_2872,N_1086,N_1955);
and U2873 (N_2873,N_1625,N_1155);
or U2874 (N_2874,N_1326,N_1864);
and U2875 (N_2875,N_1244,N_1220);
and U2876 (N_2876,N_1171,N_1548);
nor U2877 (N_2877,N_1683,N_1939);
nor U2878 (N_2878,N_1019,N_1916);
and U2879 (N_2879,N_1259,N_1079);
xnor U2880 (N_2880,N_1081,N_1473);
nand U2881 (N_2881,N_1462,N_1860);
or U2882 (N_2882,N_1899,N_1687);
and U2883 (N_2883,N_1769,N_1342);
nand U2884 (N_2884,N_1509,N_1961);
nor U2885 (N_2885,N_1894,N_1472);
nor U2886 (N_2886,N_1853,N_1862);
nand U2887 (N_2887,N_1942,N_1807);
and U2888 (N_2888,N_1388,N_1946);
nand U2889 (N_2889,N_1554,N_1534);
nand U2890 (N_2890,N_1305,N_1385);
nand U2891 (N_2891,N_1057,N_1310);
or U2892 (N_2892,N_1568,N_1484);
nand U2893 (N_2893,N_1850,N_1333);
xor U2894 (N_2894,N_1917,N_1374);
or U2895 (N_2895,N_1283,N_1531);
or U2896 (N_2896,N_1960,N_1840);
and U2897 (N_2897,N_1156,N_1781);
xor U2898 (N_2898,N_1452,N_1790);
nand U2899 (N_2899,N_1006,N_1149);
nand U2900 (N_2900,N_1157,N_1427);
nand U2901 (N_2901,N_1623,N_1703);
xor U2902 (N_2902,N_1646,N_1698);
or U2903 (N_2903,N_1363,N_1375);
or U2904 (N_2904,N_1985,N_1497);
nor U2905 (N_2905,N_1803,N_1714);
and U2906 (N_2906,N_1560,N_1728);
nor U2907 (N_2907,N_1044,N_1999);
nand U2908 (N_2908,N_1770,N_1278);
or U2909 (N_2909,N_1465,N_1355);
and U2910 (N_2910,N_1515,N_1712);
nand U2911 (N_2911,N_1101,N_1404);
nor U2912 (N_2912,N_1431,N_1703);
or U2913 (N_2913,N_1844,N_1617);
or U2914 (N_2914,N_1973,N_1918);
or U2915 (N_2915,N_1997,N_1518);
nor U2916 (N_2916,N_1349,N_1439);
and U2917 (N_2917,N_1719,N_1419);
or U2918 (N_2918,N_1972,N_1463);
and U2919 (N_2919,N_1124,N_1620);
and U2920 (N_2920,N_1316,N_1848);
nor U2921 (N_2921,N_1826,N_1001);
nand U2922 (N_2922,N_1895,N_1058);
nand U2923 (N_2923,N_1010,N_1956);
xor U2924 (N_2924,N_1607,N_1938);
nand U2925 (N_2925,N_1577,N_1675);
nand U2926 (N_2926,N_1991,N_1875);
and U2927 (N_2927,N_1107,N_1287);
and U2928 (N_2928,N_1391,N_1972);
and U2929 (N_2929,N_1026,N_1416);
xnor U2930 (N_2930,N_1608,N_1218);
and U2931 (N_2931,N_1502,N_1568);
xor U2932 (N_2932,N_1879,N_1727);
xnor U2933 (N_2933,N_1079,N_1963);
and U2934 (N_2934,N_1313,N_1822);
or U2935 (N_2935,N_1663,N_1777);
or U2936 (N_2936,N_1294,N_1058);
nor U2937 (N_2937,N_1681,N_1922);
nor U2938 (N_2938,N_1432,N_1108);
nor U2939 (N_2939,N_1236,N_1277);
nor U2940 (N_2940,N_1257,N_1060);
or U2941 (N_2941,N_1048,N_1466);
and U2942 (N_2942,N_1136,N_1740);
and U2943 (N_2943,N_1033,N_1392);
and U2944 (N_2944,N_1706,N_1071);
nand U2945 (N_2945,N_1686,N_1290);
or U2946 (N_2946,N_1361,N_1690);
nand U2947 (N_2947,N_1507,N_1625);
nor U2948 (N_2948,N_1235,N_1097);
and U2949 (N_2949,N_1141,N_1792);
or U2950 (N_2950,N_1846,N_1347);
nand U2951 (N_2951,N_1744,N_1981);
nor U2952 (N_2952,N_1854,N_1690);
or U2953 (N_2953,N_1581,N_1490);
xor U2954 (N_2954,N_1676,N_1474);
or U2955 (N_2955,N_1190,N_1673);
and U2956 (N_2956,N_1629,N_1369);
nor U2957 (N_2957,N_1765,N_1046);
nand U2958 (N_2958,N_1666,N_1497);
xor U2959 (N_2959,N_1261,N_1351);
and U2960 (N_2960,N_1971,N_1841);
nor U2961 (N_2961,N_1999,N_1281);
or U2962 (N_2962,N_1482,N_1763);
nor U2963 (N_2963,N_1680,N_1339);
nor U2964 (N_2964,N_1267,N_1861);
and U2965 (N_2965,N_1011,N_1899);
or U2966 (N_2966,N_1851,N_1639);
or U2967 (N_2967,N_1291,N_1485);
nor U2968 (N_2968,N_1607,N_1920);
and U2969 (N_2969,N_1865,N_1839);
nor U2970 (N_2970,N_1417,N_1435);
or U2971 (N_2971,N_1045,N_1655);
or U2972 (N_2972,N_1597,N_1868);
or U2973 (N_2973,N_1147,N_1513);
nor U2974 (N_2974,N_1488,N_1332);
nor U2975 (N_2975,N_1260,N_1361);
nand U2976 (N_2976,N_1013,N_1859);
nand U2977 (N_2977,N_1664,N_1538);
nor U2978 (N_2978,N_1342,N_1173);
or U2979 (N_2979,N_1503,N_1864);
nand U2980 (N_2980,N_1534,N_1537);
or U2981 (N_2981,N_1397,N_1820);
xnor U2982 (N_2982,N_1987,N_1590);
xor U2983 (N_2983,N_1030,N_1042);
nor U2984 (N_2984,N_1209,N_1489);
nor U2985 (N_2985,N_1237,N_1426);
or U2986 (N_2986,N_1213,N_1880);
and U2987 (N_2987,N_1797,N_1915);
or U2988 (N_2988,N_1255,N_1927);
nand U2989 (N_2989,N_1996,N_1183);
xnor U2990 (N_2990,N_1638,N_1902);
or U2991 (N_2991,N_1690,N_1962);
nor U2992 (N_2992,N_1764,N_1099);
nand U2993 (N_2993,N_1674,N_1928);
nand U2994 (N_2994,N_1282,N_1140);
nor U2995 (N_2995,N_1984,N_1559);
and U2996 (N_2996,N_1306,N_1111);
or U2997 (N_2997,N_1393,N_1768);
nor U2998 (N_2998,N_1951,N_1476);
or U2999 (N_2999,N_1188,N_1934);
and U3000 (N_3000,N_2674,N_2550);
and U3001 (N_3001,N_2486,N_2769);
nor U3002 (N_3002,N_2371,N_2372);
or U3003 (N_3003,N_2730,N_2879);
nor U3004 (N_3004,N_2300,N_2154);
nand U3005 (N_3005,N_2388,N_2793);
nand U3006 (N_3006,N_2766,N_2788);
and U3007 (N_3007,N_2814,N_2297);
nand U3008 (N_3008,N_2619,N_2250);
nand U3009 (N_3009,N_2682,N_2050);
nand U3010 (N_3010,N_2129,N_2200);
or U3011 (N_3011,N_2685,N_2346);
nand U3012 (N_3012,N_2936,N_2626);
nand U3013 (N_3013,N_2510,N_2440);
or U3014 (N_3014,N_2437,N_2610);
nor U3015 (N_3015,N_2954,N_2729);
or U3016 (N_3016,N_2181,N_2801);
nor U3017 (N_3017,N_2798,N_2597);
nor U3018 (N_3018,N_2985,N_2697);
xor U3019 (N_3019,N_2802,N_2772);
nand U3020 (N_3020,N_2901,N_2148);
nor U3021 (N_3021,N_2781,N_2774);
and U3022 (N_3022,N_2585,N_2829);
nor U3023 (N_3023,N_2376,N_2184);
xor U3024 (N_3024,N_2976,N_2330);
and U3025 (N_3025,N_2928,N_2574);
nor U3026 (N_3026,N_2828,N_2799);
nand U3027 (N_3027,N_2321,N_2957);
and U3028 (N_3028,N_2015,N_2858);
nor U3029 (N_3029,N_2439,N_2961);
or U3030 (N_3030,N_2199,N_2964);
nor U3031 (N_3031,N_2659,N_2020);
and U3032 (N_3032,N_2123,N_2998);
and U3033 (N_3033,N_2456,N_2640);
or U3034 (N_3034,N_2091,N_2977);
nand U3035 (N_3035,N_2933,N_2172);
or U3036 (N_3036,N_2892,N_2744);
nor U3037 (N_3037,N_2229,N_2355);
nor U3038 (N_3038,N_2546,N_2377);
nand U3039 (N_3039,N_2225,N_2874);
nor U3040 (N_3040,N_2228,N_2883);
nand U3041 (N_3041,N_2571,N_2813);
nor U3042 (N_3042,N_2131,N_2278);
nand U3043 (N_3043,N_2084,N_2064);
xnor U3044 (N_3044,N_2467,N_2276);
nand U3045 (N_3045,N_2203,N_2182);
nand U3046 (N_3046,N_2838,N_2273);
xor U3047 (N_3047,N_2383,N_2863);
nor U3048 (N_3048,N_2833,N_2119);
and U3049 (N_3049,N_2653,N_2245);
or U3050 (N_3050,N_2533,N_2785);
and U3051 (N_3051,N_2545,N_2749);
nor U3052 (N_3052,N_2378,N_2304);
or U3053 (N_3053,N_2004,N_2623);
nand U3054 (N_3054,N_2541,N_2677);
nor U3055 (N_3055,N_2318,N_2975);
xnor U3056 (N_3056,N_2434,N_2444);
xor U3057 (N_3057,N_2691,N_2726);
or U3058 (N_3058,N_2501,N_2153);
or U3059 (N_3059,N_2221,N_2483);
nor U3060 (N_3060,N_2582,N_2641);
or U3061 (N_3061,N_2668,N_2758);
nor U3062 (N_3062,N_2683,N_2692);
nor U3063 (N_3063,N_2480,N_2116);
and U3064 (N_3064,N_2516,N_2452);
and U3065 (N_3065,N_2776,N_2227);
xor U3066 (N_3066,N_2851,N_2634);
or U3067 (N_3067,N_2596,N_2676);
nor U3068 (N_3068,N_2824,N_2521);
or U3069 (N_3069,N_2025,N_2605);
nand U3070 (N_3070,N_2435,N_2098);
and U3071 (N_3071,N_2494,N_2312);
or U3072 (N_3072,N_2862,N_2016);
and U3073 (N_3073,N_2800,N_2466);
and U3074 (N_3074,N_2359,N_2348);
and U3075 (N_3075,N_2587,N_2738);
xor U3076 (N_3076,N_2028,N_2576);
nand U3077 (N_3077,N_2812,N_2681);
nand U3078 (N_3078,N_2805,N_2556);
nand U3079 (N_3079,N_2219,N_2027);
nor U3080 (N_3080,N_2673,N_2384);
xnor U3081 (N_3081,N_2732,N_2398);
or U3082 (N_3082,N_2899,N_2941);
nor U3083 (N_3083,N_2558,N_2128);
and U3084 (N_3084,N_2872,N_2826);
nor U3085 (N_3085,N_2926,N_2881);
xnor U3086 (N_3086,N_2846,N_2115);
or U3087 (N_3087,N_2670,N_2743);
nor U3088 (N_3088,N_2657,N_2731);
or U3089 (N_3089,N_2678,N_2529);
nand U3090 (N_3090,N_2239,N_2174);
nand U3091 (N_3091,N_2306,N_2402);
nor U3092 (N_3092,N_2725,N_2260);
xor U3093 (N_3093,N_2931,N_2443);
and U3094 (N_3094,N_2827,N_2006);
xnor U3095 (N_3095,N_2996,N_2328);
xnor U3096 (N_3096,N_2196,N_2918);
nor U3097 (N_3097,N_2431,N_2042);
or U3098 (N_3098,N_2621,N_2762);
and U3099 (N_3099,N_2555,N_2269);
nor U3100 (N_3100,N_2099,N_2488);
xnor U3101 (N_3101,N_2989,N_2352);
nand U3102 (N_3102,N_2625,N_2544);
nand U3103 (N_3103,N_2473,N_2157);
xnor U3104 (N_3104,N_2747,N_2009);
xor U3105 (N_3105,N_2173,N_2547);
nor U3106 (N_3106,N_2924,N_2051);
and U3107 (N_3107,N_2295,N_2403);
or U3108 (N_3108,N_2675,N_2719);
xor U3109 (N_3109,N_2686,N_2667);
nand U3110 (N_3110,N_2096,N_2999);
nor U3111 (N_3111,N_2615,N_2748);
xnor U3112 (N_3112,N_2241,N_2648);
nand U3113 (N_3113,N_2320,N_2938);
or U3114 (N_3114,N_2255,N_2669);
nor U3115 (N_3115,N_2700,N_2343);
xnor U3116 (N_3116,N_2534,N_2518);
nand U3117 (N_3117,N_2904,N_2281);
and U3118 (N_3118,N_2303,N_2284);
or U3119 (N_3119,N_2840,N_2316);
nand U3120 (N_3120,N_2179,N_2037);
nor U3121 (N_3121,N_2289,N_2259);
or U3122 (N_3122,N_2045,N_2804);
or U3123 (N_3123,N_2076,N_2591);
and U3124 (N_3124,N_2958,N_2689);
and U3125 (N_3125,N_2716,N_2995);
nor U3126 (N_3126,N_2854,N_2424);
xnor U3127 (N_3127,N_2072,N_2275);
and U3128 (N_3128,N_2438,N_2392);
or U3129 (N_3129,N_2755,N_2986);
and U3130 (N_3130,N_2885,N_2206);
and U3131 (N_3131,N_2238,N_2540);
or U3132 (N_3132,N_2651,N_2902);
or U3133 (N_3133,N_2859,N_2167);
xor U3134 (N_3134,N_2337,N_2927);
or U3135 (N_3135,N_2477,N_2142);
nor U3136 (N_3136,N_2818,N_2039);
or U3137 (N_3137,N_2145,N_2637);
xor U3138 (N_3138,N_2213,N_2363);
or U3139 (N_3139,N_2432,N_2877);
nand U3140 (N_3140,N_2427,N_2498);
nand U3141 (N_3141,N_2897,N_2898);
or U3142 (N_3142,N_2194,N_2308);
nor U3143 (N_3143,N_2083,N_2723);
nor U3144 (N_3144,N_2500,N_2970);
and U3145 (N_3145,N_2379,N_2391);
or U3146 (N_3146,N_2387,N_2264);
or U3147 (N_3147,N_2768,N_2095);
nand U3148 (N_3148,N_2717,N_2470);
and U3149 (N_3149,N_2044,N_2141);
and U3150 (N_3150,N_2412,N_2205);
or U3151 (N_3151,N_2487,N_2207);
or U3152 (N_3152,N_2335,N_2595);
and U3153 (N_3153,N_2929,N_2548);
nor U3154 (N_3154,N_2475,N_2257);
and U3155 (N_3155,N_2442,N_2414);
nand U3156 (N_3156,N_2823,N_2132);
nor U3157 (N_3157,N_2984,N_2056);
nor U3158 (N_3158,N_2616,N_2169);
nor U3159 (N_3159,N_2422,N_2162);
xnor U3160 (N_3160,N_2476,N_2664);
and U3161 (N_3161,N_2436,N_2244);
or U3162 (N_3162,N_2048,N_2404);
and U3163 (N_3163,N_2508,N_2588);
nand U3164 (N_3164,N_2535,N_2581);
nand U3165 (N_3165,N_2043,N_2794);
and U3166 (N_3166,N_2347,N_2103);
nor U3167 (N_3167,N_2644,N_2334);
nand U3168 (N_3168,N_2313,N_2302);
nor U3169 (N_3169,N_2951,N_2850);
or U3170 (N_3170,N_2628,N_2538);
and U3171 (N_3171,N_2513,N_2127);
nand U3172 (N_3172,N_2137,N_2080);
nor U3173 (N_3173,N_2635,N_2570);
nand U3174 (N_3174,N_2703,N_2658);
nor U3175 (N_3175,N_2013,N_2565);
and U3176 (N_3176,N_2912,N_2191);
nand U3177 (N_3177,N_2698,N_2505);
nand U3178 (N_3178,N_2362,N_2557);
and U3179 (N_3179,N_2580,N_2982);
or U3180 (N_3180,N_2138,N_2638);
nor U3181 (N_3181,N_2948,N_2839);
nor U3182 (N_3182,N_2617,N_2707);
or U3183 (N_3183,N_2710,N_2946);
or U3184 (N_3184,N_2711,N_2869);
xor U3185 (N_3185,N_2240,N_2397);
nor U3186 (N_3186,N_2867,N_2599);
nand U3187 (N_3187,N_2968,N_2151);
or U3188 (N_3188,N_2413,N_2601);
nor U3189 (N_3189,N_2552,N_2822);
nor U3190 (N_3190,N_2370,N_2893);
or U3191 (N_3191,N_2003,N_2071);
and U3192 (N_3192,N_2357,N_2987);
nand U3193 (N_3193,N_2536,N_2531);
nor U3194 (N_3194,N_2290,N_2114);
nand U3195 (N_3195,N_2592,N_2147);
xor U3196 (N_3196,N_2578,N_2267);
or U3197 (N_3197,N_2124,N_2249);
or U3198 (N_3198,N_2602,N_2382);
nand U3199 (N_3199,N_2509,N_2107);
nand U3200 (N_3200,N_2230,N_2190);
or U3201 (N_3201,N_2243,N_2779);
nand U3202 (N_3202,N_2909,N_2889);
or U3203 (N_3203,N_2624,N_2469);
nand U3204 (N_3204,N_2612,N_2932);
nor U3205 (N_3205,N_2293,N_2569);
and U3206 (N_3206,N_2121,N_2282);
nand U3207 (N_3207,N_2288,N_2176);
nand U3208 (N_3208,N_2062,N_2980);
or U3209 (N_3209,N_2694,N_2763);
and U3210 (N_3210,N_2923,N_2136);
xor U3211 (N_3211,N_2420,N_2490);
and U3212 (N_3212,N_2113,N_2900);
nand U3213 (N_3213,N_2279,N_2465);
or U3214 (N_3214,N_2296,N_2507);
nor U3215 (N_3215,N_2908,N_2075);
xor U3216 (N_3216,N_2369,N_2277);
nor U3217 (N_3217,N_2706,N_2482);
or U3218 (N_3218,N_2461,N_2633);
nor U3219 (N_3219,N_2187,N_2024);
or U3220 (N_3220,N_2198,N_2563);
or U3221 (N_3221,N_2821,N_2515);
nor U3222 (N_3222,N_2778,N_2093);
or U3223 (N_3223,N_2708,N_2226);
nand U3224 (N_3224,N_2220,N_2709);
or U3225 (N_3225,N_2981,N_2770);
or U3226 (N_3226,N_2344,N_2861);
xnor U3227 (N_3227,N_2234,N_2943);
or U3228 (N_3228,N_2089,N_2242);
nor U3229 (N_3229,N_2525,N_2223);
nand U3230 (N_3230,N_2584,N_2061);
or U3231 (N_3231,N_2643,N_2849);
nand U3232 (N_3232,N_2325,N_2193);
or U3233 (N_3233,N_2600,N_2149);
nor U3234 (N_3234,N_2807,N_2265);
or U3235 (N_3235,N_2993,N_2607);
or U3236 (N_3236,N_2082,N_2971);
nor U3237 (N_3237,N_2543,N_2672);
nand U3238 (N_3238,N_2752,N_2735);
xnor U3239 (N_3239,N_2395,N_2524);
nand U3240 (N_3240,N_2088,N_2636);
nor U3241 (N_3241,N_2002,N_2474);
and U3242 (N_3242,N_2497,N_2365);
and U3243 (N_3243,N_2905,N_2063);
nor U3244 (N_3244,N_2216,N_2988);
nor U3245 (N_3245,N_2102,N_2385);
nand U3246 (N_3246,N_2029,N_2163);
or U3247 (N_3247,N_2101,N_2426);
or U3248 (N_3248,N_2125,N_2451);
nor U3249 (N_3249,N_2930,N_2155);
nor U3250 (N_3250,N_2661,N_2967);
and U3251 (N_3251,N_2159,N_2736);
nand U3252 (N_3252,N_2007,N_2140);
nor U3253 (N_3253,N_2577,N_2008);
and U3254 (N_3254,N_2342,N_2322);
nand U3255 (N_3255,N_2445,N_2459);
nor U3256 (N_3256,N_2301,N_2329);
or U3257 (N_3257,N_2575,N_2554);
or U3258 (N_3258,N_2333,N_2287);
and U3259 (N_3259,N_2396,N_2252);
or U3260 (N_3260,N_2262,N_2417);
xnor U3261 (N_3261,N_2268,N_2110);
nor U3262 (N_3262,N_2134,N_2983);
nand U3263 (N_3263,N_2573,N_2419);
nand U3264 (N_3264,N_2236,N_2105);
or U3265 (N_3265,N_2690,N_2937);
or U3266 (N_3266,N_2614,N_2094);
nor U3267 (N_3267,N_2254,N_2418);
nor U3268 (N_3268,N_2068,N_2598);
nand U3269 (N_3269,N_2796,N_2210);
nor U3270 (N_3270,N_2258,N_2608);
and U3271 (N_3271,N_2997,N_2882);
and U3272 (N_3272,N_2057,N_2049);
and U3273 (N_3273,N_2085,N_2724);
xnor U3274 (N_3274,N_2895,N_2504);
nor U3275 (N_3275,N_2652,N_2760);
and U3276 (N_3276,N_2055,N_2327);
nor U3277 (N_3277,N_2323,N_2784);
nand U3278 (N_3278,N_2311,N_2843);
nor U3279 (N_3279,N_2046,N_2665);
nand U3280 (N_3280,N_2503,N_2903);
nor U3281 (N_3281,N_2109,N_2035);
or U3282 (N_3282,N_2942,N_2916);
nor U3283 (N_3283,N_2345,N_2122);
or U3284 (N_3284,N_2884,N_2857);
nor U3285 (N_3285,N_2449,N_2914);
nor U3286 (N_3286,N_2773,N_2701);
or U3287 (N_3287,N_2520,N_2012);
nand U3288 (N_3288,N_2782,N_2713);
and U3289 (N_3289,N_2407,N_2654);
or U3290 (N_3290,N_2041,N_2000);
nand U3291 (N_3291,N_2266,N_2896);
xor U3292 (N_3292,N_2201,N_2087);
and U3293 (N_3293,N_2662,N_2058);
nor U3294 (N_3294,N_2023,N_2684);
nor U3295 (N_3295,N_2143,N_2647);
or U3296 (N_3296,N_2888,N_2511);
nor U3297 (N_3297,N_2542,N_2687);
nand U3298 (N_3298,N_2375,N_2847);
and U3299 (N_3299,N_2400,N_2561);
xor U3300 (N_3300,N_2512,N_2705);
nor U3301 (N_3301,N_2386,N_2150);
and U3302 (N_3302,N_2564,N_2650);
xor U3303 (N_3303,N_2235,N_2695);
or U3304 (N_3304,N_2714,N_2354);
or U3305 (N_3305,N_2324,N_2906);
xor U3306 (N_3306,N_2522,N_2464);
nor U3307 (N_3307,N_2118,N_2825);
and U3308 (N_3308,N_2253,N_2990);
and U3309 (N_3309,N_2117,N_2120);
nand U3310 (N_3310,N_2204,N_2646);
and U3311 (N_3311,N_2960,N_2660);
nor U3312 (N_3312,N_2441,N_2820);
or U3313 (N_3313,N_2609,N_2485);
xnor U3314 (N_3314,N_2539,N_2666);
and U3315 (N_3315,N_2034,N_2326);
and U3316 (N_3316,N_2183,N_2920);
nand U3317 (N_3317,N_2401,N_2492);
nor U3318 (N_3318,N_2972,N_2361);
nand U3319 (N_3319,N_2368,N_2491);
nand U3320 (N_3320,N_2560,N_2005);
nor U3321 (N_3321,N_2356,N_2780);
nor U3322 (N_3322,N_2146,N_2935);
or U3323 (N_3323,N_2462,N_2745);
nand U3324 (N_3324,N_2627,N_2910);
nand U3325 (N_3325,N_2759,N_2166);
nand U3326 (N_3326,N_2186,N_2502);
nor U3327 (N_3327,N_2994,N_2270);
and U3328 (N_3328,N_2519,N_2022);
or U3329 (N_3329,N_2263,N_2815);
and U3330 (N_3330,N_2848,N_2283);
nand U3331 (N_3331,N_2010,N_2215);
nor U3332 (N_3332,N_2133,N_2314);
nor U3333 (N_3333,N_2992,N_2246);
and U3334 (N_3334,N_2448,N_2594);
and U3335 (N_3335,N_2059,N_2750);
and U3336 (N_3336,N_2733,N_2453);
nand U3337 (N_3337,N_2939,N_2680);
and U3338 (N_3338,N_2630,N_2679);
or U3339 (N_3339,N_2632,N_2158);
or U3340 (N_3340,N_2712,N_2338);
nor U3341 (N_3341,N_2517,N_2272);
and U3342 (N_3342,N_2613,N_2164);
nor U3343 (N_3343,N_2819,N_2170);
nand U3344 (N_3344,N_2070,N_2471);
nor U3345 (N_3345,N_2073,N_2878);
xnor U3346 (N_3346,N_2484,N_2298);
xnor U3347 (N_3347,N_2830,N_2030);
nand U3348 (N_3348,N_2952,N_2969);
nor U3349 (N_3349,N_2855,N_2197);
xnor U3350 (N_3350,N_2891,N_2792);
nor U3351 (N_3351,N_2727,N_2887);
nor U3352 (N_3352,N_2721,N_2754);
and U3353 (N_3353,N_2523,N_2699);
and U3354 (N_3354,N_2751,N_2195);
or U3355 (N_3355,N_2702,N_2175);
nor U3356 (N_3356,N_2532,N_2100);
and U3357 (N_3357,N_2069,N_2880);
and U3358 (N_3358,N_2618,N_2551);
nor U3359 (N_3359,N_2086,N_2693);
and U3360 (N_3360,N_2586,N_2890);
nand U3361 (N_3361,N_2374,N_2081);
or U3362 (N_3362,N_2292,N_2139);
nand U3363 (N_3363,N_2966,N_2108);
nor U3364 (N_3364,N_2688,N_2649);
or U3365 (N_3365,N_2496,N_2017);
and U3366 (N_3366,N_2457,N_2911);
nand U3367 (N_3367,N_2790,N_2033);
nor U3368 (N_3368,N_2373,N_2870);
nor U3369 (N_3369,N_2310,N_2789);
and U3370 (N_3370,N_2366,N_2405);
and U3371 (N_3371,N_2589,N_2741);
or U3372 (N_3372,N_2737,N_2720);
and U3373 (N_3373,N_2715,N_2415);
nand U3374 (N_3374,N_2349,N_2604);
xor U3375 (N_3375,N_2481,N_2499);
nor U3376 (N_3376,N_2844,N_2963);
or U3377 (N_3377,N_2468,N_2130);
and U3378 (N_3378,N_2810,N_2358);
and U3379 (N_3379,N_2251,N_2168);
nand U3380 (N_3380,N_2797,N_2078);
xor U3381 (N_3381,N_2014,N_2180);
nor U3382 (N_3382,N_2332,N_2307);
and U3383 (N_3383,N_2959,N_2286);
xor U3384 (N_3384,N_2568,N_2777);
or U3385 (N_3385,N_2757,N_2962);
nand U3386 (N_3386,N_2052,N_2066);
nor U3387 (N_3387,N_2026,N_2663);
nor U3388 (N_3388,N_2450,N_2340);
xnor U3389 (N_3389,N_2171,N_2309);
xnor U3390 (N_3390,N_2562,N_2416);
and U3391 (N_3391,N_2074,N_2917);
nor U3392 (N_3392,N_2144,N_2177);
and U3393 (N_3393,N_2156,N_2873);
and U3394 (N_3394,N_2831,N_2161);
or U3395 (N_3395,N_2835,N_2606);
or U3396 (N_3396,N_2746,N_2421);
nand U3397 (N_3397,N_2603,N_2836);
and U3398 (N_3398,N_2925,N_2274);
nor U3399 (N_3399,N_2202,N_2054);
nand U3400 (N_3400,N_2528,N_2280);
nor U3401 (N_3401,N_2866,N_2423);
nor U3402 (N_3402,N_2019,N_2549);
and U3403 (N_3403,N_2940,N_2237);
xor U3404 (N_3404,N_2360,N_2655);
or U3405 (N_3405,N_2742,N_2077);
nor U3406 (N_3406,N_2631,N_2092);
nand U3407 (N_3407,N_2067,N_2408);
nor U3408 (N_3408,N_2865,N_2734);
or U3409 (N_3409,N_2559,N_2430);
nor U3410 (N_3410,N_2811,N_2806);
and U3411 (N_3411,N_2222,N_2217);
nand U3412 (N_3412,N_2740,N_2090);
and U3413 (N_3413,N_2152,N_2611);
nand U3414 (N_3414,N_2947,N_2231);
xor U3415 (N_3415,N_2868,N_2214);
and U3416 (N_3416,N_2786,N_2319);
nor U3417 (N_3417,N_2261,N_2852);
nor U3418 (N_3418,N_2506,N_2425);
nor U3419 (N_3419,N_2915,N_2886);
nor U3420 (N_3420,N_2209,N_2871);
xnor U3421 (N_3421,N_2919,N_2514);
and U3422 (N_3422,N_2192,N_2285);
nor U3423 (N_3423,N_2950,N_2864);
nor U3424 (N_3424,N_2922,N_2718);
nor U3425 (N_3425,N_2189,N_2894);
and U3426 (N_3426,N_2350,N_2956);
nand U3427 (N_3427,N_2876,N_2394);
or U3428 (N_3428,N_2765,N_2639);
xnor U3429 (N_3429,N_2188,N_2527);
nand U3430 (N_3430,N_2271,N_2097);
or U3431 (N_3431,N_2429,N_2853);
nand U3432 (N_3432,N_2803,N_2447);
and U3433 (N_3433,N_2208,N_2001);
and U3434 (N_3434,N_2949,N_2489);
nor U3435 (N_3435,N_2978,N_2381);
or U3436 (N_3436,N_2291,N_2671);
and U3437 (N_3437,N_2339,N_2390);
and U3438 (N_3438,N_2460,N_2380);
or U3439 (N_3439,N_2256,N_2106);
and U3440 (N_3440,N_2944,N_2248);
and U3441 (N_3441,N_2856,N_2126);
and U3442 (N_3442,N_2218,N_2934);
or U3443 (N_3443,N_2053,N_2472);
nor U3444 (N_3444,N_2845,N_2620);
nand U3445 (N_3445,N_2341,N_2247);
nor U3446 (N_3446,N_2065,N_2040);
nand U3447 (N_3447,N_2353,N_2526);
nand U3448 (N_3448,N_2454,N_2572);
and U3449 (N_3449,N_2060,N_2364);
and U3450 (N_3450,N_2767,N_2583);
and U3451 (N_3451,N_2367,N_2795);
nand U3452 (N_3452,N_2233,N_2808);
nor U3453 (N_3453,N_2458,N_2047);
nand U3454 (N_3454,N_2530,N_2955);
or U3455 (N_3455,N_2656,N_2590);
nor U3456 (N_3456,N_2428,N_2409);
or U3457 (N_3457,N_2593,N_2834);
nand U3458 (N_3458,N_2135,N_2816);
or U3459 (N_3459,N_2455,N_2704);
xnor U3460 (N_3460,N_2493,N_2479);
and U3461 (N_3461,N_2974,N_2739);
and U3462 (N_3462,N_2771,N_2495);
nor U3463 (N_3463,N_2446,N_2224);
or U3464 (N_3464,N_2764,N_2178);
and U3465 (N_3465,N_2331,N_2953);
nor U3466 (N_3466,N_2406,N_2791);
nor U3467 (N_3467,N_2478,N_2579);
or U3468 (N_3468,N_2991,N_2299);
and U3469 (N_3469,N_2775,N_2553);
or U3470 (N_3470,N_2079,N_2032);
or U3471 (N_3471,N_2111,N_2756);
or U3472 (N_3472,N_2160,N_2393);
or U3473 (N_3473,N_2761,N_2753);
xor U3474 (N_3474,N_2038,N_2317);
nand U3475 (N_3475,N_2165,N_2629);
nor U3476 (N_3476,N_2294,N_2832);
or U3477 (N_3477,N_2907,N_2973);
or U3478 (N_3478,N_2315,N_2809);
or U3479 (N_3479,N_2021,N_2945);
and U3480 (N_3480,N_2913,N_2837);
xnor U3481 (N_3481,N_2567,N_2566);
or U3482 (N_3482,N_2433,N_2232);
and U3483 (N_3483,N_2842,N_2211);
nand U3484 (N_3484,N_2875,N_2696);
or U3485 (N_3485,N_2860,N_2411);
nand U3486 (N_3486,N_2011,N_2305);
nor U3487 (N_3487,N_2645,N_2537);
or U3488 (N_3488,N_2410,N_2787);
and U3489 (N_3489,N_2841,N_2185);
or U3490 (N_3490,N_2399,N_2018);
and U3491 (N_3491,N_2722,N_2728);
and U3492 (N_3492,N_2965,N_2921);
nor U3493 (N_3493,N_2817,N_2112);
nor U3494 (N_3494,N_2783,N_2622);
or U3495 (N_3495,N_2642,N_2031);
or U3496 (N_3496,N_2351,N_2336);
nand U3497 (N_3497,N_2979,N_2212);
nand U3498 (N_3498,N_2104,N_2389);
nand U3499 (N_3499,N_2036,N_2463);
nand U3500 (N_3500,N_2334,N_2679);
nand U3501 (N_3501,N_2332,N_2384);
or U3502 (N_3502,N_2726,N_2856);
nor U3503 (N_3503,N_2387,N_2574);
or U3504 (N_3504,N_2984,N_2033);
nand U3505 (N_3505,N_2569,N_2128);
and U3506 (N_3506,N_2986,N_2762);
nand U3507 (N_3507,N_2142,N_2552);
nand U3508 (N_3508,N_2658,N_2085);
and U3509 (N_3509,N_2567,N_2368);
nor U3510 (N_3510,N_2430,N_2528);
or U3511 (N_3511,N_2417,N_2996);
xor U3512 (N_3512,N_2380,N_2271);
or U3513 (N_3513,N_2125,N_2485);
nor U3514 (N_3514,N_2175,N_2615);
nor U3515 (N_3515,N_2888,N_2584);
and U3516 (N_3516,N_2172,N_2287);
or U3517 (N_3517,N_2822,N_2614);
nor U3518 (N_3518,N_2519,N_2990);
xnor U3519 (N_3519,N_2373,N_2025);
or U3520 (N_3520,N_2569,N_2337);
xor U3521 (N_3521,N_2937,N_2198);
and U3522 (N_3522,N_2384,N_2568);
and U3523 (N_3523,N_2727,N_2421);
nor U3524 (N_3524,N_2955,N_2294);
nor U3525 (N_3525,N_2785,N_2165);
and U3526 (N_3526,N_2051,N_2503);
xnor U3527 (N_3527,N_2683,N_2431);
or U3528 (N_3528,N_2203,N_2882);
nor U3529 (N_3529,N_2705,N_2212);
nor U3530 (N_3530,N_2606,N_2336);
or U3531 (N_3531,N_2300,N_2945);
nand U3532 (N_3532,N_2724,N_2189);
and U3533 (N_3533,N_2350,N_2085);
nor U3534 (N_3534,N_2572,N_2910);
and U3535 (N_3535,N_2912,N_2146);
nand U3536 (N_3536,N_2766,N_2849);
or U3537 (N_3537,N_2410,N_2926);
nand U3538 (N_3538,N_2281,N_2031);
nand U3539 (N_3539,N_2841,N_2683);
and U3540 (N_3540,N_2118,N_2586);
nand U3541 (N_3541,N_2730,N_2225);
and U3542 (N_3542,N_2743,N_2415);
nand U3543 (N_3543,N_2656,N_2579);
nand U3544 (N_3544,N_2924,N_2543);
or U3545 (N_3545,N_2180,N_2940);
and U3546 (N_3546,N_2573,N_2899);
nand U3547 (N_3547,N_2127,N_2105);
or U3548 (N_3548,N_2471,N_2424);
or U3549 (N_3549,N_2446,N_2209);
nand U3550 (N_3550,N_2482,N_2596);
nor U3551 (N_3551,N_2132,N_2762);
nand U3552 (N_3552,N_2903,N_2260);
or U3553 (N_3553,N_2703,N_2366);
and U3554 (N_3554,N_2240,N_2955);
xnor U3555 (N_3555,N_2950,N_2115);
nor U3556 (N_3556,N_2945,N_2652);
or U3557 (N_3557,N_2238,N_2052);
nand U3558 (N_3558,N_2277,N_2721);
xor U3559 (N_3559,N_2726,N_2947);
and U3560 (N_3560,N_2123,N_2928);
and U3561 (N_3561,N_2397,N_2176);
nor U3562 (N_3562,N_2299,N_2362);
or U3563 (N_3563,N_2262,N_2092);
or U3564 (N_3564,N_2430,N_2263);
or U3565 (N_3565,N_2986,N_2975);
nor U3566 (N_3566,N_2149,N_2596);
nand U3567 (N_3567,N_2569,N_2452);
nand U3568 (N_3568,N_2825,N_2589);
nand U3569 (N_3569,N_2363,N_2105);
nor U3570 (N_3570,N_2142,N_2113);
or U3571 (N_3571,N_2820,N_2782);
nor U3572 (N_3572,N_2699,N_2121);
nand U3573 (N_3573,N_2048,N_2007);
xor U3574 (N_3574,N_2829,N_2158);
xnor U3575 (N_3575,N_2225,N_2628);
or U3576 (N_3576,N_2434,N_2155);
nor U3577 (N_3577,N_2928,N_2556);
or U3578 (N_3578,N_2872,N_2080);
or U3579 (N_3579,N_2207,N_2273);
and U3580 (N_3580,N_2884,N_2870);
and U3581 (N_3581,N_2987,N_2544);
xor U3582 (N_3582,N_2584,N_2665);
nand U3583 (N_3583,N_2057,N_2773);
xnor U3584 (N_3584,N_2151,N_2429);
and U3585 (N_3585,N_2482,N_2049);
nor U3586 (N_3586,N_2256,N_2473);
nand U3587 (N_3587,N_2831,N_2481);
nor U3588 (N_3588,N_2556,N_2576);
nor U3589 (N_3589,N_2076,N_2375);
nand U3590 (N_3590,N_2992,N_2805);
nand U3591 (N_3591,N_2383,N_2988);
nor U3592 (N_3592,N_2098,N_2300);
nor U3593 (N_3593,N_2485,N_2237);
nor U3594 (N_3594,N_2076,N_2426);
and U3595 (N_3595,N_2795,N_2183);
and U3596 (N_3596,N_2380,N_2442);
nand U3597 (N_3597,N_2549,N_2619);
and U3598 (N_3598,N_2435,N_2243);
nand U3599 (N_3599,N_2811,N_2539);
nor U3600 (N_3600,N_2898,N_2657);
nand U3601 (N_3601,N_2909,N_2578);
and U3602 (N_3602,N_2221,N_2028);
nand U3603 (N_3603,N_2479,N_2997);
nand U3604 (N_3604,N_2300,N_2183);
and U3605 (N_3605,N_2413,N_2829);
nand U3606 (N_3606,N_2144,N_2297);
and U3607 (N_3607,N_2230,N_2053);
and U3608 (N_3608,N_2111,N_2799);
or U3609 (N_3609,N_2261,N_2759);
or U3610 (N_3610,N_2742,N_2937);
and U3611 (N_3611,N_2461,N_2562);
and U3612 (N_3612,N_2772,N_2773);
and U3613 (N_3613,N_2573,N_2094);
nor U3614 (N_3614,N_2806,N_2891);
and U3615 (N_3615,N_2562,N_2124);
and U3616 (N_3616,N_2191,N_2941);
and U3617 (N_3617,N_2631,N_2220);
nand U3618 (N_3618,N_2654,N_2933);
or U3619 (N_3619,N_2723,N_2681);
nor U3620 (N_3620,N_2215,N_2563);
or U3621 (N_3621,N_2253,N_2222);
and U3622 (N_3622,N_2415,N_2238);
or U3623 (N_3623,N_2152,N_2918);
xor U3624 (N_3624,N_2883,N_2974);
or U3625 (N_3625,N_2798,N_2372);
nand U3626 (N_3626,N_2751,N_2595);
or U3627 (N_3627,N_2068,N_2808);
nor U3628 (N_3628,N_2954,N_2629);
and U3629 (N_3629,N_2566,N_2134);
nor U3630 (N_3630,N_2713,N_2461);
nand U3631 (N_3631,N_2938,N_2067);
or U3632 (N_3632,N_2571,N_2913);
xnor U3633 (N_3633,N_2350,N_2584);
nand U3634 (N_3634,N_2705,N_2726);
nand U3635 (N_3635,N_2725,N_2747);
and U3636 (N_3636,N_2511,N_2375);
xor U3637 (N_3637,N_2826,N_2521);
nor U3638 (N_3638,N_2512,N_2876);
nor U3639 (N_3639,N_2588,N_2029);
and U3640 (N_3640,N_2880,N_2006);
nand U3641 (N_3641,N_2645,N_2860);
nor U3642 (N_3642,N_2453,N_2110);
and U3643 (N_3643,N_2458,N_2459);
nand U3644 (N_3644,N_2966,N_2747);
nand U3645 (N_3645,N_2756,N_2914);
nand U3646 (N_3646,N_2608,N_2714);
nor U3647 (N_3647,N_2627,N_2458);
or U3648 (N_3648,N_2777,N_2165);
nand U3649 (N_3649,N_2935,N_2967);
or U3650 (N_3650,N_2254,N_2561);
nor U3651 (N_3651,N_2590,N_2681);
or U3652 (N_3652,N_2285,N_2855);
and U3653 (N_3653,N_2419,N_2369);
and U3654 (N_3654,N_2581,N_2995);
and U3655 (N_3655,N_2276,N_2146);
nor U3656 (N_3656,N_2978,N_2061);
nor U3657 (N_3657,N_2430,N_2153);
nor U3658 (N_3658,N_2157,N_2740);
and U3659 (N_3659,N_2718,N_2897);
nor U3660 (N_3660,N_2384,N_2297);
and U3661 (N_3661,N_2310,N_2686);
or U3662 (N_3662,N_2026,N_2734);
or U3663 (N_3663,N_2035,N_2983);
xnor U3664 (N_3664,N_2852,N_2916);
nand U3665 (N_3665,N_2096,N_2437);
or U3666 (N_3666,N_2908,N_2247);
or U3667 (N_3667,N_2521,N_2963);
nand U3668 (N_3668,N_2478,N_2717);
and U3669 (N_3669,N_2856,N_2884);
and U3670 (N_3670,N_2927,N_2583);
and U3671 (N_3671,N_2214,N_2073);
and U3672 (N_3672,N_2048,N_2649);
and U3673 (N_3673,N_2658,N_2962);
or U3674 (N_3674,N_2022,N_2591);
nor U3675 (N_3675,N_2818,N_2257);
and U3676 (N_3676,N_2205,N_2017);
nand U3677 (N_3677,N_2539,N_2979);
nor U3678 (N_3678,N_2545,N_2372);
nand U3679 (N_3679,N_2853,N_2893);
nand U3680 (N_3680,N_2618,N_2318);
nand U3681 (N_3681,N_2418,N_2238);
nand U3682 (N_3682,N_2841,N_2242);
xnor U3683 (N_3683,N_2540,N_2067);
nor U3684 (N_3684,N_2684,N_2683);
or U3685 (N_3685,N_2484,N_2872);
nand U3686 (N_3686,N_2709,N_2593);
and U3687 (N_3687,N_2996,N_2529);
nand U3688 (N_3688,N_2736,N_2203);
or U3689 (N_3689,N_2924,N_2456);
and U3690 (N_3690,N_2811,N_2808);
and U3691 (N_3691,N_2066,N_2743);
xor U3692 (N_3692,N_2884,N_2638);
nor U3693 (N_3693,N_2711,N_2071);
or U3694 (N_3694,N_2556,N_2199);
or U3695 (N_3695,N_2618,N_2039);
or U3696 (N_3696,N_2310,N_2135);
nor U3697 (N_3697,N_2694,N_2318);
and U3698 (N_3698,N_2600,N_2871);
nor U3699 (N_3699,N_2039,N_2855);
nor U3700 (N_3700,N_2154,N_2551);
or U3701 (N_3701,N_2096,N_2787);
and U3702 (N_3702,N_2951,N_2993);
xnor U3703 (N_3703,N_2572,N_2737);
or U3704 (N_3704,N_2463,N_2167);
nor U3705 (N_3705,N_2994,N_2381);
nor U3706 (N_3706,N_2339,N_2723);
nand U3707 (N_3707,N_2959,N_2006);
nor U3708 (N_3708,N_2788,N_2514);
nand U3709 (N_3709,N_2480,N_2354);
nand U3710 (N_3710,N_2715,N_2887);
and U3711 (N_3711,N_2636,N_2285);
nand U3712 (N_3712,N_2675,N_2134);
nand U3713 (N_3713,N_2879,N_2434);
and U3714 (N_3714,N_2592,N_2196);
nand U3715 (N_3715,N_2964,N_2229);
or U3716 (N_3716,N_2715,N_2702);
nand U3717 (N_3717,N_2626,N_2854);
or U3718 (N_3718,N_2222,N_2483);
and U3719 (N_3719,N_2310,N_2711);
nand U3720 (N_3720,N_2000,N_2326);
and U3721 (N_3721,N_2171,N_2941);
or U3722 (N_3722,N_2925,N_2386);
nor U3723 (N_3723,N_2042,N_2727);
and U3724 (N_3724,N_2467,N_2129);
and U3725 (N_3725,N_2850,N_2811);
xor U3726 (N_3726,N_2078,N_2681);
or U3727 (N_3727,N_2239,N_2828);
and U3728 (N_3728,N_2767,N_2162);
xnor U3729 (N_3729,N_2315,N_2334);
and U3730 (N_3730,N_2879,N_2703);
xnor U3731 (N_3731,N_2716,N_2259);
nand U3732 (N_3732,N_2196,N_2515);
nand U3733 (N_3733,N_2493,N_2341);
nand U3734 (N_3734,N_2039,N_2644);
nor U3735 (N_3735,N_2921,N_2973);
nand U3736 (N_3736,N_2031,N_2152);
nor U3737 (N_3737,N_2413,N_2111);
and U3738 (N_3738,N_2380,N_2550);
or U3739 (N_3739,N_2933,N_2456);
and U3740 (N_3740,N_2740,N_2176);
nand U3741 (N_3741,N_2480,N_2709);
nand U3742 (N_3742,N_2805,N_2347);
nand U3743 (N_3743,N_2776,N_2816);
or U3744 (N_3744,N_2366,N_2458);
or U3745 (N_3745,N_2239,N_2883);
and U3746 (N_3746,N_2514,N_2548);
or U3747 (N_3747,N_2541,N_2738);
nand U3748 (N_3748,N_2394,N_2599);
nor U3749 (N_3749,N_2659,N_2954);
xor U3750 (N_3750,N_2128,N_2483);
and U3751 (N_3751,N_2993,N_2723);
or U3752 (N_3752,N_2466,N_2865);
nand U3753 (N_3753,N_2931,N_2870);
nand U3754 (N_3754,N_2515,N_2779);
nor U3755 (N_3755,N_2391,N_2390);
and U3756 (N_3756,N_2081,N_2604);
nor U3757 (N_3757,N_2465,N_2980);
xor U3758 (N_3758,N_2788,N_2389);
and U3759 (N_3759,N_2681,N_2093);
xor U3760 (N_3760,N_2726,N_2659);
nor U3761 (N_3761,N_2510,N_2186);
nor U3762 (N_3762,N_2665,N_2450);
nand U3763 (N_3763,N_2950,N_2623);
and U3764 (N_3764,N_2658,N_2298);
nand U3765 (N_3765,N_2041,N_2281);
nor U3766 (N_3766,N_2144,N_2373);
and U3767 (N_3767,N_2606,N_2196);
nor U3768 (N_3768,N_2536,N_2177);
and U3769 (N_3769,N_2220,N_2276);
or U3770 (N_3770,N_2122,N_2287);
and U3771 (N_3771,N_2051,N_2557);
xnor U3772 (N_3772,N_2600,N_2096);
and U3773 (N_3773,N_2907,N_2596);
and U3774 (N_3774,N_2807,N_2142);
xor U3775 (N_3775,N_2265,N_2566);
xor U3776 (N_3776,N_2772,N_2309);
nand U3777 (N_3777,N_2288,N_2106);
nor U3778 (N_3778,N_2662,N_2340);
nand U3779 (N_3779,N_2948,N_2355);
and U3780 (N_3780,N_2289,N_2162);
nand U3781 (N_3781,N_2547,N_2767);
and U3782 (N_3782,N_2314,N_2253);
or U3783 (N_3783,N_2311,N_2477);
and U3784 (N_3784,N_2879,N_2633);
or U3785 (N_3785,N_2209,N_2954);
nand U3786 (N_3786,N_2036,N_2501);
and U3787 (N_3787,N_2119,N_2992);
and U3788 (N_3788,N_2577,N_2892);
nor U3789 (N_3789,N_2144,N_2403);
nor U3790 (N_3790,N_2552,N_2681);
or U3791 (N_3791,N_2553,N_2019);
and U3792 (N_3792,N_2469,N_2895);
nand U3793 (N_3793,N_2778,N_2651);
xnor U3794 (N_3794,N_2507,N_2523);
or U3795 (N_3795,N_2020,N_2701);
or U3796 (N_3796,N_2721,N_2894);
nand U3797 (N_3797,N_2679,N_2107);
nand U3798 (N_3798,N_2700,N_2470);
nand U3799 (N_3799,N_2500,N_2342);
and U3800 (N_3800,N_2720,N_2194);
or U3801 (N_3801,N_2170,N_2296);
nor U3802 (N_3802,N_2370,N_2529);
xor U3803 (N_3803,N_2661,N_2963);
and U3804 (N_3804,N_2628,N_2873);
or U3805 (N_3805,N_2709,N_2590);
nor U3806 (N_3806,N_2736,N_2315);
or U3807 (N_3807,N_2633,N_2837);
and U3808 (N_3808,N_2371,N_2718);
and U3809 (N_3809,N_2823,N_2970);
nand U3810 (N_3810,N_2585,N_2681);
nor U3811 (N_3811,N_2775,N_2340);
or U3812 (N_3812,N_2010,N_2665);
nand U3813 (N_3813,N_2102,N_2565);
nor U3814 (N_3814,N_2564,N_2000);
nand U3815 (N_3815,N_2034,N_2363);
nand U3816 (N_3816,N_2265,N_2183);
nor U3817 (N_3817,N_2673,N_2483);
xnor U3818 (N_3818,N_2780,N_2244);
nor U3819 (N_3819,N_2595,N_2217);
nand U3820 (N_3820,N_2006,N_2633);
nor U3821 (N_3821,N_2573,N_2013);
xnor U3822 (N_3822,N_2451,N_2565);
xnor U3823 (N_3823,N_2570,N_2243);
or U3824 (N_3824,N_2859,N_2758);
nand U3825 (N_3825,N_2741,N_2460);
nor U3826 (N_3826,N_2366,N_2634);
nand U3827 (N_3827,N_2486,N_2309);
nor U3828 (N_3828,N_2992,N_2138);
or U3829 (N_3829,N_2984,N_2851);
and U3830 (N_3830,N_2343,N_2919);
nand U3831 (N_3831,N_2720,N_2722);
nand U3832 (N_3832,N_2970,N_2524);
and U3833 (N_3833,N_2985,N_2986);
xnor U3834 (N_3834,N_2888,N_2925);
or U3835 (N_3835,N_2370,N_2270);
xnor U3836 (N_3836,N_2298,N_2621);
nor U3837 (N_3837,N_2013,N_2399);
nor U3838 (N_3838,N_2139,N_2544);
nor U3839 (N_3839,N_2487,N_2728);
or U3840 (N_3840,N_2848,N_2521);
and U3841 (N_3841,N_2746,N_2159);
or U3842 (N_3842,N_2577,N_2494);
or U3843 (N_3843,N_2455,N_2819);
nand U3844 (N_3844,N_2722,N_2496);
and U3845 (N_3845,N_2120,N_2935);
nand U3846 (N_3846,N_2478,N_2903);
nor U3847 (N_3847,N_2196,N_2816);
nor U3848 (N_3848,N_2075,N_2380);
and U3849 (N_3849,N_2127,N_2236);
xnor U3850 (N_3850,N_2574,N_2370);
xnor U3851 (N_3851,N_2984,N_2263);
or U3852 (N_3852,N_2239,N_2909);
nor U3853 (N_3853,N_2965,N_2113);
and U3854 (N_3854,N_2358,N_2671);
and U3855 (N_3855,N_2703,N_2840);
or U3856 (N_3856,N_2333,N_2370);
or U3857 (N_3857,N_2566,N_2126);
nor U3858 (N_3858,N_2699,N_2376);
or U3859 (N_3859,N_2597,N_2660);
or U3860 (N_3860,N_2861,N_2548);
or U3861 (N_3861,N_2637,N_2635);
and U3862 (N_3862,N_2368,N_2904);
and U3863 (N_3863,N_2132,N_2924);
nand U3864 (N_3864,N_2695,N_2973);
xor U3865 (N_3865,N_2084,N_2942);
or U3866 (N_3866,N_2463,N_2406);
and U3867 (N_3867,N_2163,N_2544);
or U3868 (N_3868,N_2019,N_2061);
nand U3869 (N_3869,N_2177,N_2538);
nor U3870 (N_3870,N_2247,N_2777);
and U3871 (N_3871,N_2448,N_2443);
and U3872 (N_3872,N_2054,N_2526);
nor U3873 (N_3873,N_2571,N_2831);
and U3874 (N_3874,N_2992,N_2023);
nand U3875 (N_3875,N_2505,N_2656);
nand U3876 (N_3876,N_2804,N_2613);
nor U3877 (N_3877,N_2683,N_2727);
nand U3878 (N_3878,N_2330,N_2318);
nor U3879 (N_3879,N_2870,N_2874);
or U3880 (N_3880,N_2022,N_2307);
nor U3881 (N_3881,N_2223,N_2553);
or U3882 (N_3882,N_2340,N_2272);
and U3883 (N_3883,N_2599,N_2127);
and U3884 (N_3884,N_2561,N_2592);
xor U3885 (N_3885,N_2789,N_2473);
nand U3886 (N_3886,N_2037,N_2452);
nor U3887 (N_3887,N_2563,N_2357);
xnor U3888 (N_3888,N_2840,N_2873);
and U3889 (N_3889,N_2699,N_2434);
and U3890 (N_3890,N_2498,N_2745);
or U3891 (N_3891,N_2471,N_2788);
or U3892 (N_3892,N_2772,N_2341);
or U3893 (N_3893,N_2272,N_2192);
nand U3894 (N_3894,N_2660,N_2889);
xor U3895 (N_3895,N_2105,N_2647);
and U3896 (N_3896,N_2537,N_2883);
nor U3897 (N_3897,N_2485,N_2835);
nand U3898 (N_3898,N_2887,N_2521);
and U3899 (N_3899,N_2752,N_2517);
and U3900 (N_3900,N_2968,N_2286);
or U3901 (N_3901,N_2050,N_2456);
or U3902 (N_3902,N_2311,N_2333);
nand U3903 (N_3903,N_2202,N_2457);
and U3904 (N_3904,N_2329,N_2697);
or U3905 (N_3905,N_2764,N_2467);
nor U3906 (N_3906,N_2557,N_2372);
xnor U3907 (N_3907,N_2371,N_2018);
and U3908 (N_3908,N_2664,N_2712);
nand U3909 (N_3909,N_2650,N_2409);
and U3910 (N_3910,N_2787,N_2933);
nand U3911 (N_3911,N_2861,N_2723);
and U3912 (N_3912,N_2792,N_2348);
or U3913 (N_3913,N_2498,N_2208);
nand U3914 (N_3914,N_2379,N_2222);
nor U3915 (N_3915,N_2346,N_2147);
or U3916 (N_3916,N_2140,N_2857);
and U3917 (N_3917,N_2062,N_2288);
and U3918 (N_3918,N_2035,N_2422);
or U3919 (N_3919,N_2125,N_2274);
nand U3920 (N_3920,N_2803,N_2727);
nand U3921 (N_3921,N_2481,N_2525);
nand U3922 (N_3922,N_2190,N_2497);
nand U3923 (N_3923,N_2599,N_2036);
nor U3924 (N_3924,N_2428,N_2009);
xnor U3925 (N_3925,N_2529,N_2413);
nor U3926 (N_3926,N_2507,N_2964);
or U3927 (N_3927,N_2005,N_2569);
and U3928 (N_3928,N_2262,N_2611);
or U3929 (N_3929,N_2860,N_2518);
nor U3930 (N_3930,N_2824,N_2525);
nand U3931 (N_3931,N_2883,N_2671);
nand U3932 (N_3932,N_2438,N_2282);
nor U3933 (N_3933,N_2640,N_2651);
nor U3934 (N_3934,N_2801,N_2745);
or U3935 (N_3935,N_2705,N_2993);
xnor U3936 (N_3936,N_2824,N_2752);
and U3937 (N_3937,N_2874,N_2130);
or U3938 (N_3938,N_2829,N_2438);
nand U3939 (N_3939,N_2757,N_2961);
and U3940 (N_3940,N_2081,N_2649);
xnor U3941 (N_3941,N_2256,N_2429);
nand U3942 (N_3942,N_2698,N_2048);
nor U3943 (N_3943,N_2780,N_2097);
and U3944 (N_3944,N_2034,N_2239);
or U3945 (N_3945,N_2079,N_2100);
or U3946 (N_3946,N_2692,N_2320);
and U3947 (N_3947,N_2035,N_2658);
xor U3948 (N_3948,N_2283,N_2813);
or U3949 (N_3949,N_2845,N_2078);
xnor U3950 (N_3950,N_2682,N_2839);
and U3951 (N_3951,N_2801,N_2438);
and U3952 (N_3952,N_2579,N_2675);
nand U3953 (N_3953,N_2713,N_2215);
or U3954 (N_3954,N_2688,N_2568);
nor U3955 (N_3955,N_2442,N_2281);
nand U3956 (N_3956,N_2007,N_2364);
and U3957 (N_3957,N_2064,N_2650);
and U3958 (N_3958,N_2169,N_2883);
or U3959 (N_3959,N_2033,N_2699);
nand U3960 (N_3960,N_2088,N_2639);
or U3961 (N_3961,N_2271,N_2546);
nand U3962 (N_3962,N_2846,N_2507);
nor U3963 (N_3963,N_2486,N_2982);
and U3964 (N_3964,N_2305,N_2702);
or U3965 (N_3965,N_2046,N_2894);
or U3966 (N_3966,N_2115,N_2391);
nand U3967 (N_3967,N_2254,N_2606);
nand U3968 (N_3968,N_2332,N_2871);
and U3969 (N_3969,N_2015,N_2515);
xor U3970 (N_3970,N_2171,N_2670);
and U3971 (N_3971,N_2112,N_2972);
nor U3972 (N_3972,N_2656,N_2991);
and U3973 (N_3973,N_2286,N_2389);
nor U3974 (N_3974,N_2718,N_2674);
xnor U3975 (N_3975,N_2891,N_2027);
xor U3976 (N_3976,N_2865,N_2226);
nor U3977 (N_3977,N_2837,N_2159);
and U3978 (N_3978,N_2521,N_2737);
or U3979 (N_3979,N_2357,N_2484);
xnor U3980 (N_3980,N_2568,N_2919);
nor U3981 (N_3981,N_2995,N_2914);
xnor U3982 (N_3982,N_2677,N_2077);
nor U3983 (N_3983,N_2736,N_2638);
nand U3984 (N_3984,N_2352,N_2502);
or U3985 (N_3985,N_2741,N_2882);
nand U3986 (N_3986,N_2312,N_2558);
xnor U3987 (N_3987,N_2736,N_2039);
nand U3988 (N_3988,N_2790,N_2022);
or U3989 (N_3989,N_2470,N_2755);
or U3990 (N_3990,N_2288,N_2629);
nand U3991 (N_3991,N_2435,N_2856);
xnor U3992 (N_3992,N_2400,N_2818);
nand U3993 (N_3993,N_2166,N_2363);
nor U3994 (N_3994,N_2126,N_2049);
nor U3995 (N_3995,N_2566,N_2792);
or U3996 (N_3996,N_2336,N_2034);
nand U3997 (N_3997,N_2629,N_2999);
nor U3998 (N_3998,N_2820,N_2726);
nor U3999 (N_3999,N_2346,N_2652);
or U4000 (N_4000,N_3169,N_3499);
nand U4001 (N_4001,N_3543,N_3170);
or U4002 (N_4002,N_3295,N_3808);
nor U4003 (N_4003,N_3761,N_3740);
and U4004 (N_4004,N_3519,N_3141);
nand U4005 (N_4005,N_3276,N_3282);
nand U4006 (N_4006,N_3721,N_3887);
or U4007 (N_4007,N_3696,N_3552);
nand U4008 (N_4008,N_3832,N_3949);
and U4009 (N_4009,N_3825,N_3620);
and U4010 (N_4010,N_3258,N_3707);
and U4011 (N_4011,N_3588,N_3171);
and U4012 (N_4012,N_3708,N_3946);
or U4013 (N_4013,N_3792,N_3078);
nor U4014 (N_4014,N_3383,N_3524);
or U4015 (N_4015,N_3624,N_3550);
and U4016 (N_4016,N_3851,N_3812);
and U4017 (N_4017,N_3065,N_3712);
and U4018 (N_4018,N_3862,N_3309);
nor U4019 (N_4019,N_3021,N_3965);
xor U4020 (N_4020,N_3109,N_3474);
nor U4021 (N_4021,N_3354,N_3496);
and U4022 (N_4022,N_3268,N_3894);
nand U4023 (N_4023,N_3113,N_3000);
and U4024 (N_4024,N_3444,N_3306);
xor U4025 (N_4025,N_3183,N_3586);
and U4026 (N_4026,N_3424,N_3771);
xor U4027 (N_4027,N_3015,N_3039);
nor U4028 (N_4028,N_3980,N_3538);
or U4029 (N_4029,N_3226,N_3540);
and U4030 (N_4030,N_3714,N_3323);
xnor U4031 (N_4031,N_3618,N_3683);
or U4032 (N_4032,N_3345,N_3180);
or U4033 (N_4033,N_3558,N_3725);
nor U4034 (N_4034,N_3191,N_3446);
nor U4035 (N_4035,N_3824,N_3728);
nor U4036 (N_4036,N_3619,N_3351);
and U4037 (N_4037,N_3574,N_3206);
or U4038 (N_4038,N_3755,N_3794);
nor U4039 (N_4039,N_3119,N_3998);
and U4040 (N_4040,N_3938,N_3184);
nor U4041 (N_4041,N_3421,N_3981);
or U4042 (N_4042,N_3944,N_3898);
nor U4043 (N_4043,N_3148,N_3733);
and U4044 (N_4044,N_3880,N_3147);
xor U4045 (N_4045,N_3986,N_3906);
nor U4046 (N_4046,N_3172,N_3259);
nor U4047 (N_4047,N_3304,N_3360);
and U4048 (N_4048,N_3572,N_3263);
and U4049 (N_4049,N_3956,N_3156);
or U4050 (N_4050,N_3705,N_3407);
or U4051 (N_4051,N_3387,N_3372);
nor U4052 (N_4052,N_3168,N_3318);
or U4053 (N_4053,N_3530,N_3943);
or U4054 (N_4054,N_3891,N_3215);
and U4055 (N_4055,N_3048,N_3094);
nor U4056 (N_4056,N_3577,N_3012);
or U4057 (N_4057,N_3357,N_3283);
and U4058 (N_4058,N_3365,N_3265);
nor U4059 (N_4059,N_3589,N_3816);
or U4060 (N_4060,N_3062,N_3117);
nor U4061 (N_4061,N_3413,N_3320);
nand U4062 (N_4062,N_3236,N_3801);
and U4063 (N_4063,N_3674,N_3487);
and U4064 (N_4064,N_3715,N_3079);
or U4065 (N_4065,N_3930,N_3899);
nand U4066 (N_4066,N_3381,N_3256);
or U4067 (N_4067,N_3702,N_3827);
nand U4068 (N_4068,N_3692,N_3270);
or U4069 (N_4069,N_3132,N_3479);
nor U4070 (N_4070,N_3770,N_3881);
nor U4071 (N_4071,N_3330,N_3607);
nor U4072 (N_4072,N_3778,N_3626);
or U4073 (N_4073,N_3272,N_3598);
or U4074 (N_4074,N_3888,N_3672);
nand U4075 (N_4075,N_3326,N_3368);
or U4076 (N_4076,N_3815,N_3573);
nand U4077 (N_4077,N_3562,N_3810);
xor U4078 (N_4078,N_3690,N_3918);
nor U4079 (N_4079,N_3511,N_3685);
nand U4080 (N_4080,N_3393,N_3566);
nor U4081 (N_4081,N_3190,N_3466);
nor U4082 (N_4082,N_3652,N_3205);
and U4083 (N_4083,N_3961,N_3353);
nor U4084 (N_4084,N_3146,N_3252);
and U4085 (N_4085,N_3197,N_3092);
nand U4086 (N_4086,N_3045,N_3260);
or U4087 (N_4087,N_3996,N_3068);
nand U4088 (N_4088,N_3214,N_3303);
and U4089 (N_4089,N_3704,N_3369);
and U4090 (N_4090,N_3315,N_3143);
or U4091 (N_4091,N_3570,N_3599);
and U4092 (N_4092,N_3322,N_3130);
nor U4093 (N_4093,N_3697,N_3941);
nand U4094 (N_4094,N_3793,N_3426);
and U4095 (N_4095,N_3483,N_3419);
and U4096 (N_4096,N_3207,N_3164);
xor U4097 (N_4097,N_3001,N_3642);
or U4098 (N_4098,N_3166,N_3768);
nor U4099 (N_4099,N_3105,N_3789);
xnor U4100 (N_4100,N_3405,N_3352);
or U4101 (N_4101,N_3913,N_3960);
nor U4102 (N_4102,N_3547,N_3036);
and U4103 (N_4103,N_3748,N_3211);
or U4104 (N_4104,N_3641,N_3947);
or U4105 (N_4105,N_3507,N_3933);
xnor U4106 (N_4106,N_3379,N_3654);
nand U4107 (N_4107,N_3010,N_3890);
and U4108 (N_4108,N_3449,N_3083);
nor U4109 (N_4109,N_3706,N_3845);
nor U4110 (N_4110,N_3163,N_3992);
and U4111 (N_4111,N_3797,N_3134);
or U4112 (N_4112,N_3514,N_3679);
nor U4113 (N_4113,N_3003,N_3592);
nand U4114 (N_4114,N_3433,N_3610);
or U4115 (N_4115,N_3394,N_3814);
or U4116 (N_4116,N_3836,N_3729);
nand U4117 (N_4117,N_3803,N_3374);
or U4118 (N_4118,N_3942,N_3159);
or U4119 (N_4119,N_3210,N_3773);
nand U4120 (N_4120,N_3600,N_3666);
and U4121 (N_4121,N_3209,N_3907);
and U4122 (N_4122,N_3527,N_3532);
xor U4123 (N_4123,N_3288,N_3711);
nand U4124 (N_4124,N_3084,N_3482);
or U4125 (N_4125,N_3217,N_3175);
xor U4126 (N_4126,N_3723,N_3865);
or U4127 (N_4127,N_3945,N_3468);
and U4128 (N_4128,N_3126,N_3248);
or U4129 (N_4129,N_3990,N_3766);
or U4130 (N_4130,N_3489,N_3905);
or U4131 (N_4131,N_3024,N_3388);
or U4132 (N_4132,N_3877,N_3979);
or U4133 (N_4133,N_3718,N_3492);
and U4134 (N_4134,N_3673,N_3809);
or U4135 (N_4135,N_3587,N_3701);
nor U4136 (N_4136,N_3621,N_3634);
or U4137 (N_4137,N_3627,N_3680);
nor U4138 (N_4138,N_3615,N_3359);
nor U4139 (N_4139,N_3834,N_3929);
xor U4140 (N_4140,N_3380,N_3462);
or U4141 (N_4141,N_3328,N_3194);
nand U4142 (N_4142,N_3515,N_3070);
or U4143 (N_4143,N_3958,N_3135);
and U4144 (N_4144,N_3555,N_3075);
or U4145 (N_4145,N_3281,N_3237);
or U4146 (N_4146,N_3266,N_3417);
xor U4147 (N_4147,N_3640,N_3886);
and U4148 (N_4148,N_3123,N_3089);
or U4149 (N_4149,N_3734,N_3107);
nor U4150 (N_4150,N_3777,N_3046);
and U4151 (N_4151,N_3860,N_3554);
xnor U4152 (N_4152,N_3428,N_3301);
and U4153 (N_4153,N_3875,N_3931);
nand U4154 (N_4154,N_3285,N_3686);
nor U4155 (N_4155,N_3534,N_3099);
or U4156 (N_4156,N_3578,N_3670);
nand U4157 (N_4157,N_3081,N_3478);
nor U4158 (N_4158,N_3085,N_3840);
xnor U4159 (N_4159,N_3804,N_3435);
nor U4160 (N_4160,N_3613,N_3967);
nor U4161 (N_4161,N_3067,N_3193);
nand U4162 (N_4162,N_3361,N_3103);
and U4163 (N_4163,N_3727,N_3456);
nand U4164 (N_4164,N_3779,N_3106);
nor U4165 (N_4165,N_3392,N_3593);
and U4166 (N_4166,N_3461,N_3739);
xnor U4167 (N_4167,N_3402,N_3453);
xor U4168 (N_4168,N_3014,N_3495);
nor U4169 (N_4169,N_3290,N_3513);
nand U4170 (N_4170,N_3490,N_3756);
nand U4171 (N_4171,N_3985,N_3999);
nand U4172 (N_4172,N_3028,N_3275);
and U4173 (N_4173,N_3822,N_3335);
nand U4174 (N_4174,N_3420,N_3316);
and U4175 (N_4175,N_3830,N_3299);
and U4176 (N_4176,N_3920,N_3235);
nor U4177 (N_4177,N_3498,N_3378);
nand U4178 (N_4178,N_3348,N_3994);
nand U4179 (N_4179,N_3198,N_3294);
and U4180 (N_4180,N_3928,N_3878);
and U4181 (N_4181,N_3535,N_3160);
and U4182 (N_4182,N_3430,N_3019);
and U4183 (N_4183,N_3581,N_3464);
nor U4184 (N_4184,N_3518,N_3017);
nor U4185 (N_4185,N_3800,N_3289);
and U4186 (N_4186,N_3682,N_3227);
or U4187 (N_4187,N_3653,N_3597);
and U4188 (N_4188,N_3576,N_3189);
nand U4189 (N_4189,N_3662,N_3337);
and U4190 (N_4190,N_3895,N_3410);
xnor U4191 (N_4191,N_3854,N_3525);
nor U4192 (N_4192,N_3583,N_3937);
and U4193 (N_4193,N_3041,N_3422);
nor U4194 (N_4194,N_3762,N_3063);
or U4195 (N_4195,N_3149,N_3187);
nand U4196 (N_4196,N_3745,N_3950);
and U4197 (N_4197,N_3788,N_3011);
nand U4198 (N_4198,N_3245,N_3321);
or U4199 (N_4199,N_3018,N_3279);
nand U4200 (N_4200,N_3616,N_3988);
nor U4201 (N_4201,N_3232,N_3839);
nor U4202 (N_4202,N_3628,N_3883);
nor U4203 (N_4203,N_3546,N_3885);
xor U4204 (N_4204,N_3549,N_3658);
and U4205 (N_4205,N_3909,N_3327);
or U4206 (N_4206,N_3564,N_3848);
and U4207 (N_4207,N_3060,N_3781);
nand U4208 (N_4208,N_3310,N_3921);
and U4209 (N_4209,N_3638,N_3399);
and U4210 (N_4210,N_3450,N_3404);
nand U4211 (N_4211,N_3473,N_3516);
or U4212 (N_4212,N_3675,N_3469);
nand U4213 (N_4213,N_3142,N_3477);
nand U4214 (N_4214,N_3884,N_3689);
and U4215 (N_4215,N_3026,N_3855);
xnor U4216 (N_4216,N_3811,N_3350);
and U4217 (N_4217,N_3298,N_3648);
nand U4218 (N_4218,N_3108,N_3726);
and U4219 (N_4219,N_3805,N_3751);
or U4220 (N_4220,N_3138,N_3040);
or U4221 (N_4221,N_3951,N_3594);
nand U4222 (N_4222,N_3660,N_3425);
nand U4223 (N_4223,N_3241,N_3749);
or U4224 (N_4224,N_3630,N_3497);
nand U4225 (N_4225,N_3936,N_3287);
or U4226 (N_4226,N_3765,N_3255);
or U4227 (N_4227,N_3565,N_3661);
and U4228 (N_4228,N_3750,N_3776);
nand U4229 (N_4229,N_3769,N_3072);
or U4230 (N_4230,N_3847,N_3086);
or U4231 (N_4231,N_3485,N_3976);
or U4232 (N_4232,N_3284,N_3844);
nor U4233 (N_4233,N_3505,N_3528);
nand U4234 (N_4234,N_3775,N_3118);
nor U4235 (N_4235,N_3759,N_3784);
nor U4236 (N_4236,N_3452,N_3914);
xor U4237 (N_4237,N_3398,N_3182);
nand U4238 (N_4238,N_3694,N_3561);
or U4239 (N_4239,N_3059,N_3720);
nand U4240 (N_4240,N_3545,N_3440);
nand U4241 (N_4241,N_3858,N_3897);
and U4242 (N_4242,N_3445,N_3336);
nand U4243 (N_4243,N_3560,N_3731);
and U4244 (N_4244,N_3502,N_3659);
nor U4245 (N_4245,N_3324,N_3385);
nand U4246 (N_4246,N_3396,N_3764);
xor U4247 (N_4247,N_3719,N_3722);
nor U4248 (N_4248,N_3423,N_3828);
xor U4249 (N_4249,N_3278,N_3982);
or U4250 (N_4250,N_3475,N_3331);
nand U4251 (N_4251,N_3125,N_3140);
nand U4252 (N_4252,N_3962,N_3225);
nand U4253 (N_4253,N_3606,N_3977);
or U4254 (N_4254,N_3127,N_3850);
nand U4255 (N_4255,N_3051,N_3370);
and U4256 (N_4256,N_3458,N_3199);
nand U4257 (N_4257,N_3639,N_3054);
nor U4258 (N_4258,N_3604,N_3151);
or U4259 (N_4259,N_3438,N_3512);
nand U4260 (N_4260,N_3747,N_3664);
and U4261 (N_4261,N_3500,N_3030);
and U4262 (N_4262,N_3088,N_3744);
nor U4263 (N_4263,N_3693,N_3843);
nand U4264 (N_4264,N_3667,N_3195);
xnor U4265 (N_4265,N_3467,N_3539);
and U4266 (N_4266,N_3200,N_3742);
xnor U4267 (N_4267,N_3178,N_3677);
nand U4268 (N_4268,N_3602,N_3264);
nand U4269 (N_4269,N_3313,N_3454);
or U4270 (N_4270,N_3434,N_3614);
nand U4271 (N_4271,N_3096,N_3339);
nand U4272 (N_4272,N_3415,N_3669);
nand U4273 (N_4273,N_3073,N_3665);
and U4274 (N_4274,N_3964,N_3411);
and U4275 (N_4275,N_3635,N_3363);
and U4276 (N_4276,N_3743,N_3364);
nand U4277 (N_4277,N_3991,N_3154);
or U4278 (N_4278,N_3384,N_3754);
nor U4279 (N_4279,N_3471,N_3786);
nor U4280 (N_4280,N_3432,N_3904);
or U4281 (N_4281,N_3043,N_3857);
and U4282 (N_4282,N_3213,N_3568);
or U4283 (N_4283,N_3416,N_3317);
or U4284 (N_4284,N_3212,N_3481);
or U4285 (N_4285,N_3520,N_3542);
nor U4286 (N_4286,N_3332,N_3239);
or U4287 (N_4287,N_3185,N_3536);
nand U4288 (N_4288,N_3849,N_3655);
xor U4289 (N_4289,N_3813,N_3603);
nor U4290 (N_4290,N_3102,N_3133);
nand U4291 (N_4291,N_3716,N_3873);
nand U4292 (N_4292,N_3111,N_3228);
and U4293 (N_4293,N_3173,N_3219);
or U4294 (N_4294,N_3181,N_3650);
xor U4295 (N_4295,N_3098,N_3314);
or U4296 (N_4296,N_3293,N_3091);
nor U4297 (N_4297,N_3758,N_3344);
and U4298 (N_4298,N_3772,N_3861);
nand U4299 (N_4299,N_3736,N_3867);
nor U4300 (N_4300,N_3058,N_3637);
nor U4301 (N_4301,N_3681,N_3975);
or U4302 (N_4302,N_3596,N_3939);
xnor U4303 (N_4303,N_3934,N_3397);
nor U4304 (N_4304,N_3963,N_3161);
xnor U4305 (N_4305,N_3557,N_3767);
nor U4306 (N_4306,N_3548,N_3969);
and U4307 (N_4307,N_3129,N_3333);
and U4308 (N_4308,N_3699,N_3459);
or U4309 (N_4309,N_3870,N_3376);
xor U4310 (N_4310,N_3177,N_3732);
or U4311 (N_4311,N_3013,N_3342);
nor U4312 (N_4312,N_3863,N_3571);
or U4313 (N_4313,N_3122,N_3978);
and U4314 (N_4314,N_3935,N_3343);
nand U4315 (N_4315,N_3186,N_3710);
nand U4316 (N_4316,N_3752,N_3157);
nor U4317 (N_4317,N_3308,N_3842);
xnor U4318 (N_4318,N_3403,N_3643);
or U4319 (N_4319,N_3837,N_3373);
or U4320 (N_4320,N_3448,N_3806);
nor U4321 (N_4321,N_3508,N_3647);
or U4322 (N_4322,N_3261,N_3480);
and U4323 (N_4323,N_3790,N_3254);
nand U4324 (N_4324,N_3463,N_3908);
xnor U4325 (N_4325,N_3267,N_3005);
and U4326 (N_4326,N_3970,N_3608);
nor U4327 (N_4327,N_3429,N_3002);
nor U4328 (N_4328,N_3911,N_3957);
xor U4329 (N_4329,N_3889,N_3247);
nand U4330 (N_4330,N_3510,N_3644);
xor U4331 (N_4331,N_3069,N_3631);
and U4332 (N_4332,N_3853,N_3609);
nor U4333 (N_4333,N_3044,N_3575);
nor U4334 (N_4334,N_3037,N_3738);
or U4335 (N_4335,N_3691,N_3128);
or U4336 (N_4336,N_3240,N_3023);
nor U4337 (N_4337,N_3932,N_3819);
or U4338 (N_4338,N_3176,N_3250);
and U4339 (N_4339,N_3912,N_3919);
xor U4340 (N_4340,N_3223,N_3544);
and U4341 (N_4341,N_3179,N_3038);
and U4342 (N_4342,N_3782,N_3605);
and U4343 (N_4343,N_3846,N_3273);
and U4344 (N_4344,N_3229,N_3537);
nor U4345 (N_4345,N_3533,N_3076);
and U4346 (N_4346,N_3307,N_3503);
or U4347 (N_4347,N_3050,N_3645);
and U4348 (N_4348,N_3636,N_3869);
and U4349 (N_4349,N_3162,N_3188);
nor U4350 (N_4350,N_3506,N_3153);
xor U4351 (N_4351,N_3874,N_3136);
nor U4352 (N_4352,N_3795,N_3852);
or U4353 (N_4353,N_3968,N_3902);
nand U4354 (N_4354,N_3901,N_3823);
nor U4355 (N_4355,N_3917,N_3053);
and U4356 (N_4356,N_3406,N_3915);
nand U4357 (N_4357,N_3006,N_3451);
or U4358 (N_4358,N_3676,N_3066);
nor U4359 (N_4359,N_3280,N_3218);
and U4360 (N_4360,N_3238,N_3349);
nand U4361 (N_4361,N_3055,N_3971);
nand U4362 (N_4362,N_3972,N_3983);
and U4363 (N_4363,N_3052,N_3391);
nor U4364 (N_4364,N_3818,N_3152);
nand U4365 (N_4365,N_3703,N_3080);
nand U4366 (N_4366,N_3955,N_3663);
xor U4367 (N_4367,N_3753,N_3892);
nand U4368 (N_4368,N_3022,N_3780);
nor U4369 (N_4369,N_3174,N_3923);
and U4370 (N_4370,N_3879,N_3296);
and U4371 (N_4371,N_3717,N_3526);
or U4372 (N_4372,N_3437,N_3995);
xnor U4373 (N_4373,N_3925,N_3121);
or U4374 (N_4374,N_3124,N_3243);
nor U4375 (N_4375,N_3087,N_3559);
nor U4376 (N_4376,N_3684,N_3027);
and U4377 (N_4377,N_3484,N_3807);
or U4378 (N_4378,N_3047,N_3042);
and U4379 (N_4379,N_3334,N_3427);
and U4380 (N_4380,N_3251,N_3418);
or U4381 (N_4381,N_3612,N_3799);
nand U4382 (N_4382,N_3035,N_3580);
and U4383 (N_4383,N_3071,N_3305);
nor U4384 (N_4384,N_3622,N_3004);
or U4385 (N_4385,N_3355,N_3927);
nor U4386 (N_4386,N_3460,N_3436);
xnor U4387 (N_4387,N_3486,N_3472);
nor U4388 (N_4388,N_3760,N_3838);
nand U4389 (N_4389,N_3651,N_3476);
nand U4390 (N_4390,N_3953,N_3131);
nand U4391 (N_4391,N_3220,N_3896);
xor U4392 (N_4392,N_3903,N_3112);
or U4393 (N_4393,N_3367,N_3292);
or U4394 (N_4394,N_3582,N_3698);
and U4395 (N_4395,N_3590,N_3442);
and U4396 (N_4396,N_3623,N_3144);
and U4397 (N_4397,N_3034,N_3922);
nor U4398 (N_4398,N_3443,N_3077);
xnor U4399 (N_4399,N_3488,N_3257);
nor U4400 (N_4400,N_3989,N_3277);
or U4401 (N_4401,N_3090,N_3517);
nand U4402 (N_4402,N_3671,N_3431);
nand U4403 (N_4403,N_3414,N_3329);
nand U4404 (N_4404,N_3649,N_3493);
and U4405 (N_4405,N_3954,N_3893);
nand U4406 (N_4406,N_3774,N_3796);
or U4407 (N_4407,N_3523,N_3678);
nor U4408 (N_4408,N_3216,N_3959);
nor U4409 (N_4409,N_3763,N_3591);
and U4410 (N_4410,N_3082,N_3286);
or U4411 (N_4411,N_3504,N_3139);
nor U4412 (N_4412,N_3868,N_3700);
or U4413 (N_4413,N_3377,N_3032);
xnor U4414 (N_4414,N_3730,N_3491);
nor U4415 (N_4415,N_3916,N_3551);
xor U4416 (N_4416,N_3595,N_3300);
nand U4417 (N_4417,N_3031,N_3409);
or U4418 (N_4418,N_3116,N_3926);
or U4419 (N_4419,N_3356,N_3390);
nand U4420 (N_4420,N_3470,N_3695);
nor U4421 (N_4421,N_3829,N_3375);
nand U4422 (N_4422,N_3632,N_3882);
nor U4423 (N_4423,N_3033,N_3231);
xnor U4424 (N_4424,N_3900,N_3521);
nand U4425 (N_4425,N_3340,N_3871);
and U4426 (N_4426,N_3371,N_3110);
and U4427 (N_4427,N_3668,N_3093);
and U4428 (N_4428,N_3522,N_3100);
and U4429 (N_4429,N_3095,N_3222);
xor U4430 (N_4430,N_3584,N_3757);
nand U4431 (N_4431,N_3579,N_3441);
and U4432 (N_4432,N_3529,N_3319);
nor U4433 (N_4433,N_3246,N_3097);
and U4434 (N_4434,N_3791,N_3202);
or U4435 (N_4435,N_3952,N_3611);
or U4436 (N_4436,N_3233,N_3074);
and U4437 (N_4437,N_3984,N_3563);
nand U4438 (N_4438,N_3509,N_3987);
and U4439 (N_4439,N_3709,N_3966);
nor U4440 (N_4440,N_3338,N_3876);
or U4441 (N_4441,N_3687,N_3291);
or U4442 (N_4442,N_3221,N_3688);
xor U4443 (N_4443,N_3553,N_3234);
nand U4444 (N_4444,N_3457,N_3785);
nor U4445 (N_4445,N_3724,N_3826);
or U4446 (N_4446,N_3556,N_3020);
xnor U4447 (N_4447,N_3325,N_3646);
or U4448 (N_4448,N_3585,N_3856);
or U4449 (N_4449,N_3016,N_3567);
or U4450 (N_4450,N_3269,N_3569);
nand U4451 (N_4451,N_3401,N_3008);
or U4452 (N_4452,N_3201,N_3347);
nand U4453 (N_4453,N_3833,N_3137);
and U4454 (N_4454,N_3057,N_3993);
nor U4455 (N_4455,N_3866,N_3798);
or U4456 (N_4456,N_3341,N_3271);
and U4457 (N_4457,N_3737,N_3311);
and U4458 (N_4458,N_3244,N_3049);
and U4459 (N_4459,N_3948,N_3872);
and U4460 (N_4460,N_3297,N_3841);
nand U4461 (N_4461,N_3115,N_3910);
or U4462 (N_4462,N_3165,N_3974);
or U4463 (N_4463,N_3859,N_3312);
nand U4464 (N_4464,N_3713,N_3625);
and U4465 (N_4465,N_3224,N_3657);
nor U4466 (N_4466,N_3362,N_3346);
nand U4467 (N_4467,N_3208,N_3787);
and U4468 (N_4468,N_3382,N_3120);
nand U4469 (N_4469,N_3007,N_3064);
nor U4470 (N_4470,N_3009,N_3358);
and U4471 (N_4471,N_3395,N_3104);
and U4472 (N_4472,N_3465,N_3746);
xnor U4473 (N_4473,N_3501,N_3389);
nand U4474 (N_4474,N_3101,N_3302);
nor U4475 (N_4475,N_3203,N_3997);
nand U4476 (N_4476,N_3262,N_3817);
nand U4477 (N_4477,N_3835,N_3155);
and U4478 (N_4478,N_3494,N_3366);
and U4479 (N_4479,N_3242,N_3455);
nor U4480 (N_4480,N_3820,N_3629);
nor U4481 (N_4481,N_3802,N_3025);
nand U4482 (N_4482,N_3617,N_3656);
nor U4483 (N_4483,N_3940,N_3735);
nor U4484 (N_4484,N_3447,N_3114);
xor U4485 (N_4485,N_3150,N_3167);
nor U4486 (N_4486,N_3633,N_3531);
nand U4487 (N_4487,N_3783,N_3821);
nand U4488 (N_4488,N_3249,N_3924);
and U4489 (N_4489,N_3158,N_3408);
nand U4490 (N_4490,N_3230,N_3439);
and U4491 (N_4491,N_3864,N_3831);
xnor U4492 (N_4492,N_3741,N_3145);
and U4493 (N_4493,N_3204,N_3541);
nor U4494 (N_4494,N_3253,N_3973);
and U4495 (N_4495,N_3029,N_3274);
xor U4496 (N_4496,N_3412,N_3601);
and U4497 (N_4497,N_3400,N_3192);
and U4498 (N_4498,N_3061,N_3386);
xor U4499 (N_4499,N_3056,N_3196);
nand U4500 (N_4500,N_3710,N_3501);
nand U4501 (N_4501,N_3268,N_3014);
nor U4502 (N_4502,N_3952,N_3994);
and U4503 (N_4503,N_3038,N_3261);
xor U4504 (N_4504,N_3615,N_3632);
or U4505 (N_4505,N_3580,N_3710);
nand U4506 (N_4506,N_3991,N_3107);
nand U4507 (N_4507,N_3296,N_3642);
nand U4508 (N_4508,N_3251,N_3683);
or U4509 (N_4509,N_3307,N_3460);
and U4510 (N_4510,N_3023,N_3074);
and U4511 (N_4511,N_3152,N_3714);
nor U4512 (N_4512,N_3143,N_3155);
and U4513 (N_4513,N_3699,N_3975);
and U4514 (N_4514,N_3854,N_3114);
or U4515 (N_4515,N_3679,N_3663);
or U4516 (N_4516,N_3447,N_3660);
xor U4517 (N_4517,N_3650,N_3276);
nor U4518 (N_4518,N_3628,N_3178);
and U4519 (N_4519,N_3088,N_3644);
nand U4520 (N_4520,N_3519,N_3681);
nand U4521 (N_4521,N_3625,N_3975);
nand U4522 (N_4522,N_3591,N_3852);
nand U4523 (N_4523,N_3154,N_3838);
or U4524 (N_4524,N_3748,N_3164);
nor U4525 (N_4525,N_3546,N_3990);
or U4526 (N_4526,N_3273,N_3286);
xor U4527 (N_4527,N_3593,N_3365);
nand U4528 (N_4528,N_3238,N_3572);
and U4529 (N_4529,N_3743,N_3137);
and U4530 (N_4530,N_3126,N_3808);
nor U4531 (N_4531,N_3893,N_3041);
or U4532 (N_4532,N_3994,N_3310);
nor U4533 (N_4533,N_3140,N_3487);
nor U4534 (N_4534,N_3715,N_3034);
xor U4535 (N_4535,N_3255,N_3510);
or U4536 (N_4536,N_3925,N_3654);
nor U4537 (N_4537,N_3315,N_3016);
nor U4538 (N_4538,N_3155,N_3900);
or U4539 (N_4539,N_3803,N_3989);
and U4540 (N_4540,N_3911,N_3604);
or U4541 (N_4541,N_3685,N_3634);
xor U4542 (N_4542,N_3484,N_3242);
nand U4543 (N_4543,N_3467,N_3643);
and U4544 (N_4544,N_3779,N_3508);
nand U4545 (N_4545,N_3876,N_3366);
or U4546 (N_4546,N_3767,N_3912);
nand U4547 (N_4547,N_3777,N_3766);
nor U4548 (N_4548,N_3198,N_3533);
or U4549 (N_4549,N_3765,N_3514);
and U4550 (N_4550,N_3155,N_3130);
and U4551 (N_4551,N_3181,N_3686);
nor U4552 (N_4552,N_3746,N_3299);
and U4553 (N_4553,N_3941,N_3168);
nor U4554 (N_4554,N_3541,N_3960);
nor U4555 (N_4555,N_3099,N_3778);
nand U4556 (N_4556,N_3389,N_3585);
nor U4557 (N_4557,N_3039,N_3636);
nor U4558 (N_4558,N_3193,N_3664);
and U4559 (N_4559,N_3702,N_3606);
or U4560 (N_4560,N_3715,N_3754);
or U4561 (N_4561,N_3521,N_3174);
nor U4562 (N_4562,N_3035,N_3115);
and U4563 (N_4563,N_3341,N_3447);
nand U4564 (N_4564,N_3878,N_3626);
nor U4565 (N_4565,N_3025,N_3203);
and U4566 (N_4566,N_3168,N_3749);
nor U4567 (N_4567,N_3702,N_3749);
and U4568 (N_4568,N_3095,N_3614);
nor U4569 (N_4569,N_3468,N_3239);
nand U4570 (N_4570,N_3852,N_3136);
or U4571 (N_4571,N_3461,N_3229);
nor U4572 (N_4572,N_3238,N_3256);
or U4573 (N_4573,N_3355,N_3567);
and U4574 (N_4574,N_3870,N_3556);
or U4575 (N_4575,N_3097,N_3440);
or U4576 (N_4576,N_3888,N_3574);
and U4577 (N_4577,N_3073,N_3187);
and U4578 (N_4578,N_3016,N_3509);
xnor U4579 (N_4579,N_3374,N_3213);
nand U4580 (N_4580,N_3164,N_3769);
and U4581 (N_4581,N_3525,N_3393);
xor U4582 (N_4582,N_3462,N_3492);
nand U4583 (N_4583,N_3588,N_3809);
or U4584 (N_4584,N_3460,N_3376);
and U4585 (N_4585,N_3126,N_3774);
or U4586 (N_4586,N_3675,N_3511);
nand U4587 (N_4587,N_3213,N_3602);
nand U4588 (N_4588,N_3202,N_3928);
nand U4589 (N_4589,N_3416,N_3725);
nor U4590 (N_4590,N_3103,N_3437);
nand U4591 (N_4591,N_3541,N_3337);
nand U4592 (N_4592,N_3325,N_3850);
or U4593 (N_4593,N_3769,N_3624);
xnor U4594 (N_4594,N_3673,N_3050);
nand U4595 (N_4595,N_3314,N_3807);
nor U4596 (N_4596,N_3612,N_3141);
and U4597 (N_4597,N_3163,N_3108);
nor U4598 (N_4598,N_3974,N_3903);
xnor U4599 (N_4599,N_3156,N_3597);
or U4600 (N_4600,N_3347,N_3364);
xnor U4601 (N_4601,N_3527,N_3574);
and U4602 (N_4602,N_3708,N_3199);
or U4603 (N_4603,N_3989,N_3901);
nand U4604 (N_4604,N_3073,N_3940);
or U4605 (N_4605,N_3374,N_3517);
and U4606 (N_4606,N_3388,N_3688);
nor U4607 (N_4607,N_3194,N_3676);
xnor U4608 (N_4608,N_3536,N_3218);
nand U4609 (N_4609,N_3313,N_3466);
and U4610 (N_4610,N_3816,N_3029);
or U4611 (N_4611,N_3251,N_3808);
nor U4612 (N_4612,N_3873,N_3349);
and U4613 (N_4613,N_3964,N_3120);
nor U4614 (N_4614,N_3571,N_3649);
nand U4615 (N_4615,N_3970,N_3304);
nor U4616 (N_4616,N_3315,N_3967);
or U4617 (N_4617,N_3231,N_3929);
and U4618 (N_4618,N_3353,N_3178);
nand U4619 (N_4619,N_3899,N_3509);
nor U4620 (N_4620,N_3273,N_3968);
xor U4621 (N_4621,N_3706,N_3617);
nor U4622 (N_4622,N_3386,N_3478);
nor U4623 (N_4623,N_3402,N_3858);
and U4624 (N_4624,N_3316,N_3984);
nor U4625 (N_4625,N_3987,N_3297);
or U4626 (N_4626,N_3864,N_3127);
or U4627 (N_4627,N_3097,N_3120);
or U4628 (N_4628,N_3044,N_3732);
nor U4629 (N_4629,N_3139,N_3816);
xor U4630 (N_4630,N_3147,N_3976);
and U4631 (N_4631,N_3822,N_3127);
nor U4632 (N_4632,N_3120,N_3310);
or U4633 (N_4633,N_3839,N_3604);
and U4634 (N_4634,N_3979,N_3726);
or U4635 (N_4635,N_3395,N_3387);
or U4636 (N_4636,N_3282,N_3368);
nand U4637 (N_4637,N_3809,N_3213);
or U4638 (N_4638,N_3053,N_3785);
or U4639 (N_4639,N_3394,N_3162);
nor U4640 (N_4640,N_3152,N_3078);
and U4641 (N_4641,N_3438,N_3996);
nor U4642 (N_4642,N_3077,N_3938);
nand U4643 (N_4643,N_3827,N_3429);
nand U4644 (N_4644,N_3604,N_3610);
nor U4645 (N_4645,N_3668,N_3291);
and U4646 (N_4646,N_3780,N_3973);
and U4647 (N_4647,N_3380,N_3426);
xor U4648 (N_4648,N_3963,N_3518);
nand U4649 (N_4649,N_3269,N_3156);
nor U4650 (N_4650,N_3747,N_3880);
nand U4651 (N_4651,N_3476,N_3189);
or U4652 (N_4652,N_3589,N_3245);
nor U4653 (N_4653,N_3536,N_3814);
nand U4654 (N_4654,N_3111,N_3498);
or U4655 (N_4655,N_3698,N_3670);
nand U4656 (N_4656,N_3277,N_3833);
and U4657 (N_4657,N_3276,N_3835);
nand U4658 (N_4658,N_3500,N_3579);
or U4659 (N_4659,N_3199,N_3418);
xor U4660 (N_4660,N_3804,N_3838);
xnor U4661 (N_4661,N_3830,N_3079);
xor U4662 (N_4662,N_3632,N_3023);
and U4663 (N_4663,N_3469,N_3245);
nor U4664 (N_4664,N_3183,N_3465);
nor U4665 (N_4665,N_3672,N_3887);
nor U4666 (N_4666,N_3364,N_3778);
nand U4667 (N_4667,N_3720,N_3037);
nor U4668 (N_4668,N_3543,N_3943);
nand U4669 (N_4669,N_3414,N_3779);
nand U4670 (N_4670,N_3140,N_3142);
xnor U4671 (N_4671,N_3881,N_3838);
and U4672 (N_4672,N_3760,N_3511);
or U4673 (N_4673,N_3341,N_3675);
nor U4674 (N_4674,N_3605,N_3178);
nor U4675 (N_4675,N_3217,N_3706);
xor U4676 (N_4676,N_3084,N_3353);
or U4677 (N_4677,N_3946,N_3159);
and U4678 (N_4678,N_3312,N_3797);
or U4679 (N_4679,N_3209,N_3731);
nand U4680 (N_4680,N_3008,N_3873);
or U4681 (N_4681,N_3880,N_3573);
nand U4682 (N_4682,N_3162,N_3802);
nor U4683 (N_4683,N_3124,N_3980);
or U4684 (N_4684,N_3470,N_3144);
or U4685 (N_4685,N_3620,N_3411);
nand U4686 (N_4686,N_3367,N_3366);
and U4687 (N_4687,N_3473,N_3709);
or U4688 (N_4688,N_3712,N_3705);
nand U4689 (N_4689,N_3852,N_3130);
or U4690 (N_4690,N_3247,N_3391);
and U4691 (N_4691,N_3730,N_3876);
nor U4692 (N_4692,N_3242,N_3032);
and U4693 (N_4693,N_3308,N_3990);
or U4694 (N_4694,N_3248,N_3774);
or U4695 (N_4695,N_3820,N_3603);
nand U4696 (N_4696,N_3645,N_3741);
and U4697 (N_4697,N_3227,N_3140);
nand U4698 (N_4698,N_3410,N_3269);
or U4699 (N_4699,N_3061,N_3555);
xnor U4700 (N_4700,N_3340,N_3936);
or U4701 (N_4701,N_3781,N_3036);
and U4702 (N_4702,N_3783,N_3762);
xnor U4703 (N_4703,N_3451,N_3255);
nor U4704 (N_4704,N_3793,N_3078);
nor U4705 (N_4705,N_3891,N_3428);
nor U4706 (N_4706,N_3012,N_3943);
or U4707 (N_4707,N_3392,N_3468);
nor U4708 (N_4708,N_3388,N_3400);
nor U4709 (N_4709,N_3556,N_3925);
and U4710 (N_4710,N_3991,N_3425);
nand U4711 (N_4711,N_3702,N_3104);
or U4712 (N_4712,N_3834,N_3612);
and U4713 (N_4713,N_3306,N_3798);
nand U4714 (N_4714,N_3860,N_3200);
or U4715 (N_4715,N_3034,N_3050);
xnor U4716 (N_4716,N_3904,N_3149);
nor U4717 (N_4717,N_3689,N_3988);
nor U4718 (N_4718,N_3899,N_3891);
nor U4719 (N_4719,N_3218,N_3499);
or U4720 (N_4720,N_3028,N_3600);
xor U4721 (N_4721,N_3258,N_3363);
xnor U4722 (N_4722,N_3088,N_3035);
xor U4723 (N_4723,N_3233,N_3399);
and U4724 (N_4724,N_3394,N_3894);
nand U4725 (N_4725,N_3346,N_3308);
or U4726 (N_4726,N_3218,N_3543);
or U4727 (N_4727,N_3347,N_3066);
or U4728 (N_4728,N_3496,N_3210);
and U4729 (N_4729,N_3285,N_3727);
and U4730 (N_4730,N_3406,N_3158);
or U4731 (N_4731,N_3517,N_3945);
nand U4732 (N_4732,N_3498,N_3271);
or U4733 (N_4733,N_3151,N_3743);
or U4734 (N_4734,N_3196,N_3606);
or U4735 (N_4735,N_3060,N_3902);
xnor U4736 (N_4736,N_3174,N_3699);
and U4737 (N_4737,N_3545,N_3857);
and U4738 (N_4738,N_3301,N_3711);
nor U4739 (N_4739,N_3890,N_3606);
nand U4740 (N_4740,N_3811,N_3632);
xor U4741 (N_4741,N_3144,N_3392);
or U4742 (N_4742,N_3297,N_3502);
or U4743 (N_4743,N_3649,N_3103);
nand U4744 (N_4744,N_3124,N_3820);
nor U4745 (N_4745,N_3442,N_3104);
or U4746 (N_4746,N_3084,N_3126);
nor U4747 (N_4747,N_3775,N_3802);
nand U4748 (N_4748,N_3920,N_3184);
nand U4749 (N_4749,N_3557,N_3580);
or U4750 (N_4750,N_3295,N_3932);
and U4751 (N_4751,N_3104,N_3171);
nand U4752 (N_4752,N_3458,N_3810);
or U4753 (N_4753,N_3459,N_3210);
nor U4754 (N_4754,N_3781,N_3893);
and U4755 (N_4755,N_3778,N_3343);
and U4756 (N_4756,N_3282,N_3606);
and U4757 (N_4757,N_3598,N_3060);
and U4758 (N_4758,N_3721,N_3022);
nor U4759 (N_4759,N_3239,N_3322);
nand U4760 (N_4760,N_3406,N_3217);
and U4761 (N_4761,N_3463,N_3114);
or U4762 (N_4762,N_3332,N_3544);
or U4763 (N_4763,N_3442,N_3671);
nor U4764 (N_4764,N_3067,N_3151);
and U4765 (N_4765,N_3352,N_3032);
and U4766 (N_4766,N_3204,N_3946);
and U4767 (N_4767,N_3369,N_3841);
xnor U4768 (N_4768,N_3846,N_3136);
or U4769 (N_4769,N_3423,N_3720);
nand U4770 (N_4770,N_3772,N_3418);
nor U4771 (N_4771,N_3583,N_3840);
or U4772 (N_4772,N_3957,N_3582);
nand U4773 (N_4773,N_3436,N_3386);
nor U4774 (N_4774,N_3678,N_3920);
or U4775 (N_4775,N_3623,N_3311);
nor U4776 (N_4776,N_3755,N_3254);
or U4777 (N_4777,N_3149,N_3633);
or U4778 (N_4778,N_3496,N_3929);
nor U4779 (N_4779,N_3759,N_3453);
or U4780 (N_4780,N_3700,N_3671);
nand U4781 (N_4781,N_3611,N_3127);
nor U4782 (N_4782,N_3385,N_3614);
nand U4783 (N_4783,N_3214,N_3057);
nor U4784 (N_4784,N_3937,N_3291);
nand U4785 (N_4785,N_3454,N_3720);
or U4786 (N_4786,N_3803,N_3610);
nor U4787 (N_4787,N_3981,N_3193);
and U4788 (N_4788,N_3938,N_3357);
nand U4789 (N_4789,N_3995,N_3309);
or U4790 (N_4790,N_3690,N_3506);
xor U4791 (N_4791,N_3521,N_3902);
and U4792 (N_4792,N_3577,N_3721);
and U4793 (N_4793,N_3925,N_3282);
nand U4794 (N_4794,N_3596,N_3896);
nand U4795 (N_4795,N_3476,N_3821);
or U4796 (N_4796,N_3475,N_3517);
and U4797 (N_4797,N_3098,N_3940);
nor U4798 (N_4798,N_3688,N_3397);
nor U4799 (N_4799,N_3986,N_3983);
and U4800 (N_4800,N_3592,N_3990);
nor U4801 (N_4801,N_3187,N_3529);
and U4802 (N_4802,N_3733,N_3025);
or U4803 (N_4803,N_3186,N_3361);
nand U4804 (N_4804,N_3667,N_3896);
and U4805 (N_4805,N_3726,N_3128);
and U4806 (N_4806,N_3256,N_3850);
nor U4807 (N_4807,N_3806,N_3572);
nor U4808 (N_4808,N_3893,N_3841);
nor U4809 (N_4809,N_3948,N_3593);
or U4810 (N_4810,N_3878,N_3399);
nand U4811 (N_4811,N_3073,N_3183);
or U4812 (N_4812,N_3009,N_3241);
or U4813 (N_4813,N_3698,N_3692);
nand U4814 (N_4814,N_3199,N_3069);
and U4815 (N_4815,N_3617,N_3289);
or U4816 (N_4816,N_3343,N_3184);
and U4817 (N_4817,N_3973,N_3776);
and U4818 (N_4818,N_3706,N_3128);
nor U4819 (N_4819,N_3919,N_3590);
nor U4820 (N_4820,N_3492,N_3926);
or U4821 (N_4821,N_3233,N_3281);
nor U4822 (N_4822,N_3220,N_3576);
or U4823 (N_4823,N_3893,N_3455);
nor U4824 (N_4824,N_3766,N_3039);
or U4825 (N_4825,N_3112,N_3837);
nand U4826 (N_4826,N_3892,N_3717);
nor U4827 (N_4827,N_3912,N_3635);
or U4828 (N_4828,N_3462,N_3562);
or U4829 (N_4829,N_3811,N_3342);
or U4830 (N_4830,N_3759,N_3671);
and U4831 (N_4831,N_3170,N_3154);
and U4832 (N_4832,N_3408,N_3286);
nor U4833 (N_4833,N_3552,N_3551);
nor U4834 (N_4834,N_3767,N_3653);
or U4835 (N_4835,N_3684,N_3676);
or U4836 (N_4836,N_3465,N_3870);
nand U4837 (N_4837,N_3441,N_3477);
and U4838 (N_4838,N_3959,N_3272);
and U4839 (N_4839,N_3520,N_3168);
and U4840 (N_4840,N_3053,N_3214);
or U4841 (N_4841,N_3735,N_3763);
nor U4842 (N_4842,N_3249,N_3316);
or U4843 (N_4843,N_3461,N_3545);
or U4844 (N_4844,N_3446,N_3409);
nand U4845 (N_4845,N_3940,N_3865);
nor U4846 (N_4846,N_3801,N_3391);
or U4847 (N_4847,N_3419,N_3094);
nor U4848 (N_4848,N_3628,N_3598);
nand U4849 (N_4849,N_3153,N_3683);
xor U4850 (N_4850,N_3872,N_3199);
or U4851 (N_4851,N_3485,N_3780);
and U4852 (N_4852,N_3234,N_3990);
nand U4853 (N_4853,N_3521,N_3469);
nor U4854 (N_4854,N_3686,N_3306);
nor U4855 (N_4855,N_3448,N_3164);
xor U4856 (N_4856,N_3716,N_3840);
and U4857 (N_4857,N_3081,N_3523);
nor U4858 (N_4858,N_3722,N_3416);
and U4859 (N_4859,N_3372,N_3780);
nand U4860 (N_4860,N_3738,N_3193);
and U4861 (N_4861,N_3555,N_3354);
or U4862 (N_4862,N_3120,N_3296);
nor U4863 (N_4863,N_3304,N_3180);
nand U4864 (N_4864,N_3490,N_3322);
nand U4865 (N_4865,N_3102,N_3294);
and U4866 (N_4866,N_3533,N_3247);
or U4867 (N_4867,N_3654,N_3990);
or U4868 (N_4868,N_3562,N_3058);
xor U4869 (N_4869,N_3823,N_3561);
nor U4870 (N_4870,N_3112,N_3574);
and U4871 (N_4871,N_3167,N_3004);
and U4872 (N_4872,N_3056,N_3178);
nor U4873 (N_4873,N_3110,N_3784);
nand U4874 (N_4874,N_3920,N_3162);
or U4875 (N_4875,N_3163,N_3619);
and U4876 (N_4876,N_3239,N_3382);
nor U4877 (N_4877,N_3684,N_3183);
and U4878 (N_4878,N_3180,N_3526);
nor U4879 (N_4879,N_3914,N_3430);
or U4880 (N_4880,N_3138,N_3042);
xor U4881 (N_4881,N_3248,N_3587);
nor U4882 (N_4882,N_3093,N_3752);
or U4883 (N_4883,N_3509,N_3197);
and U4884 (N_4884,N_3242,N_3864);
and U4885 (N_4885,N_3629,N_3893);
nand U4886 (N_4886,N_3672,N_3406);
and U4887 (N_4887,N_3454,N_3942);
and U4888 (N_4888,N_3265,N_3191);
nand U4889 (N_4889,N_3415,N_3075);
nand U4890 (N_4890,N_3859,N_3116);
xnor U4891 (N_4891,N_3055,N_3788);
nand U4892 (N_4892,N_3055,N_3075);
and U4893 (N_4893,N_3736,N_3200);
nor U4894 (N_4894,N_3844,N_3724);
and U4895 (N_4895,N_3103,N_3665);
and U4896 (N_4896,N_3787,N_3081);
nand U4897 (N_4897,N_3223,N_3285);
xor U4898 (N_4898,N_3997,N_3006);
or U4899 (N_4899,N_3694,N_3293);
nand U4900 (N_4900,N_3118,N_3249);
and U4901 (N_4901,N_3670,N_3076);
or U4902 (N_4902,N_3393,N_3997);
nand U4903 (N_4903,N_3723,N_3785);
nand U4904 (N_4904,N_3450,N_3222);
nand U4905 (N_4905,N_3644,N_3240);
or U4906 (N_4906,N_3700,N_3116);
nand U4907 (N_4907,N_3077,N_3178);
or U4908 (N_4908,N_3393,N_3779);
nor U4909 (N_4909,N_3569,N_3781);
nor U4910 (N_4910,N_3599,N_3344);
or U4911 (N_4911,N_3980,N_3013);
and U4912 (N_4912,N_3611,N_3722);
nor U4913 (N_4913,N_3697,N_3642);
nor U4914 (N_4914,N_3819,N_3140);
or U4915 (N_4915,N_3178,N_3461);
nor U4916 (N_4916,N_3628,N_3965);
and U4917 (N_4917,N_3703,N_3406);
nor U4918 (N_4918,N_3265,N_3225);
and U4919 (N_4919,N_3854,N_3614);
or U4920 (N_4920,N_3314,N_3449);
nor U4921 (N_4921,N_3769,N_3250);
nor U4922 (N_4922,N_3928,N_3218);
and U4923 (N_4923,N_3158,N_3063);
nor U4924 (N_4924,N_3616,N_3060);
nor U4925 (N_4925,N_3354,N_3528);
nand U4926 (N_4926,N_3150,N_3479);
nand U4927 (N_4927,N_3264,N_3745);
or U4928 (N_4928,N_3723,N_3533);
xor U4929 (N_4929,N_3736,N_3136);
nand U4930 (N_4930,N_3336,N_3486);
nor U4931 (N_4931,N_3954,N_3580);
nand U4932 (N_4932,N_3903,N_3904);
and U4933 (N_4933,N_3119,N_3918);
nand U4934 (N_4934,N_3420,N_3349);
nand U4935 (N_4935,N_3180,N_3518);
nor U4936 (N_4936,N_3701,N_3533);
nand U4937 (N_4937,N_3631,N_3242);
nand U4938 (N_4938,N_3401,N_3420);
xor U4939 (N_4939,N_3157,N_3502);
and U4940 (N_4940,N_3508,N_3268);
or U4941 (N_4941,N_3296,N_3363);
nor U4942 (N_4942,N_3227,N_3909);
nor U4943 (N_4943,N_3757,N_3408);
nor U4944 (N_4944,N_3539,N_3888);
xnor U4945 (N_4945,N_3400,N_3286);
and U4946 (N_4946,N_3540,N_3824);
or U4947 (N_4947,N_3719,N_3322);
or U4948 (N_4948,N_3227,N_3517);
nand U4949 (N_4949,N_3316,N_3376);
nor U4950 (N_4950,N_3754,N_3361);
or U4951 (N_4951,N_3608,N_3535);
and U4952 (N_4952,N_3055,N_3539);
nand U4953 (N_4953,N_3823,N_3176);
or U4954 (N_4954,N_3055,N_3210);
nor U4955 (N_4955,N_3781,N_3455);
and U4956 (N_4956,N_3247,N_3677);
or U4957 (N_4957,N_3185,N_3438);
and U4958 (N_4958,N_3413,N_3343);
and U4959 (N_4959,N_3585,N_3300);
or U4960 (N_4960,N_3928,N_3358);
xnor U4961 (N_4961,N_3809,N_3159);
and U4962 (N_4962,N_3432,N_3303);
nand U4963 (N_4963,N_3136,N_3279);
nor U4964 (N_4964,N_3858,N_3234);
nor U4965 (N_4965,N_3985,N_3908);
or U4966 (N_4966,N_3439,N_3057);
and U4967 (N_4967,N_3897,N_3198);
nor U4968 (N_4968,N_3910,N_3377);
or U4969 (N_4969,N_3898,N_3931);
or U4970 (N_4970,N_3773,N_3902);
or U4971 (N_4971,N_3879,N_3391);
and U4972 (N_4972,N_3697,N_3820);
and U4973 (N_4973,N_3412,N_3747);
and U4974 (N_4974,N_3096,N_3381);
nor U4975 (N_4975,N_3414,N_3930);
nand U4976 (N_4976,N_3374,N_3234);
nand U4977 (N_4977,N_3379,N_3729);
or U4978 (N_4978,N_3265,N_3458);
nand U4979 (N_4979,N_3114,N_3176);
nor U4980 (N_4980,N_3795,N_3421);
nor U4981 (N_4981,N_3511,N_3323);
nor U4982 (N_4982,N_3292,N_3673);
nand U4983 (N_4983,N_3416,N_3040);
nand U4984 (N_4984,N_3298,N_3294);
nor U4985 (N_4985,N_3409,N_3546);
nand U4986 (N_4986,N_3328,N_3473);
and U4987 (N_4987,N_3895,N_3935);
nand U4988 (N_4988,N_3552,N_3752);
xor U4989 (N_4989,N_3780,N_3297);
or U4990 (N_4990,N_3818,N_3533);
or U4991 (N_4991,N_3570,N_3656);
nor U4992 (N_4992,N_3734,N_3018);
nor U4993 (N_4993,N_3480,N_3699);
xnor U4994 (N_4994,N_3009,N_3571);
and U4995 (N_4995,N_3005,N_3456);
or U4996 (N_4996,N_3467,N_3103);
nor U4997 (N_4997,N_3663,N_3611);
nand U4998 (N_4998,N_3093,N_3332);
nand U4999 (N_4999,N_3519,N_3662);
or U5000 (N_5000,N_4659,N_4353);
nor U5001 (N_5001,N_4280,N_4493);
nor U5002 (N_5002,N_4996,N_4157);
nand U5003 (N_5003,N_4494,N_4861);
and U5004 (N_5004,N_4173,N_4385);
or U5005 (N_5005,N_4428,N_4835);
nor U5006 (N_5006,N_4994,N_4595);
and U5007 (N_5007,N_4958,N_4352);
and U5008 (N_5008,N_4350,N_4827);
nor U5009 (N_5009,N_4452,N_4236);
and U5010 (N_5010,N_4924,N_4468);
nor U5011 (N_5011,N_4764,N_4439);
nand U5012 (N_5012,N_4107,N_4311);
or U5013 (N_5013,N_4873,N_4331);
or U5014 (N_5014,N_4471,N_4437);
nand U5015 (N_5015,N_4046,N_4127);
or U5016 (N_5016,N_4825,N_4907);
nor U5017 (N_5017,N_4482,N_4248);
and U5018 (N_5018,N_4158,N_4799);
or U5019 (N_5019,N_4866,N_4684);
nand U5020 (N_5020,N_4070,N_4637);
nand U5021 (N_5021,N_4681,N_4536);
and U5022 (N_5022,N_4770,N_4259);
and U5023 (N_5023,N_4583,N_4612);
and U5024 (N_5024,N_4765,N_4189);
nand U5025 (N_5025,N_4038,N_4445);
and U5026 (N_5026,N_4746,N_4450);
and U5027 (N_5027,N_4402,N_4997);
or U5028 (N_5028,N_4050,N_4376);
nand U5029 (N_5029,N_4335,N_4992);
nand U5030 (N_5030,N_4059,N_4601);
or U5031 (N_5031,N_4089,N_4670);
or U5032 (N_5032,N_4544,N_4296);
and U5033 (N_5033,N_4140,N_4962);
or U5034 (N_5034,N_4074,N_4118);
and U5035 (N_5035,N_4863,N_4581);
nor U5036 (N_5036,N_4441,N_4174);
xor U5037 (N_5037,N_4606,N_4965);
xnor U5038 (N_5038,N_4033,N_4704);
or U5039 (N_5039,N_4413,N_4087);
xor U5040 (N_5040,N_4200,N_4278);
nand U5041 (N_5041,N_4508,N_4917);
and U5042 (N_5042,N_4291,N_4776);
nor U5043 (N_5043,N_4198,N_4082);
and U5044 (N_5044,N_4910,N_4184);
nor U5045 (N_5045,N_4381,N_4330);
nand U5046 (N_5046,N_4404,N_4021);
nor U5047 (N_5047,N_4150,N_4665);
or U5048 (N_5048,N_4027,N_4339);
and U5049 (N_5049,N_4640,N_4206);
and U5050 (N_5050,N_4430,N_4769);
nor U5051 (N_5051,N_4516,N_4461);
nor U5052 (N_5052,N_4549,N_4496);
nor U5053 (N_5053,N_4579,N_4239);
or U5054 (N_5054,N_4946,N_4750);
or U5055 (N_5055,N_4796,N_4973);
or U5056 (N_5056,N_4609,N_4442);
nor U5057 (N_5057,N_4253,N_4929);
or U5058 (N_5058,N_4165,N_4023);
or U5059 (N_5059,N_4272,N_4409);
nor U5060 (N_5060,N_4029,N_4918);
and U5061 (N_5061,N_4592,N_4304);
or U5062 (N_5062,N_4787,N_4136);
and U5063 (N_5063,N_4137,N_4534);
nor U5064 (N_5064,N_4889,N_4963);
and U5065 (N_5065,N_4773,N_4752);
nand U5066 (N_5066,N_4618,N_4242);
nand U5067 (N_5067,N_4995,N_4129);
nand U5068 (N_5068,N_4176,N_4099);
and U5069 (N_5069,N_4346,N_4322);
nor U5070 (N_5070,N_4552,N_4328);
and U5071 (N_5071,N_4072,N_4794);
nand U5072 (N_5072,N_4811,N_4641);
and U5073 (N_5073,N_4748,N_4371);
and U5074 (N_5074,N_4833,N_4486);
and U5075 (N_5075,N_4630,N_4839);
and U5076 (N_5076,N_4542,N_4388);
nor U5077 (N_5077,N_4203,N_4451);
nor U5078 (N_5078,N_4120,N_4101);
nor U5079 (N_5079,N_4596,N_4210);
and U5080 (N_5080,N_4489,N_4897);
nand U5081 (N_5081,N_4777,N_4806);
and U5082 (N_5082,N_4491,N_4130);
and U5083 (N_5083,N_4957,N_4745);
nor U5084 (N_5084,N_4467,N_4421);
nand U5085 (N_5085,N_4423,N_4650);
or U5086 (N_5086,N_4938,N_4585);
and U5087 (N_5087,N_4808,N_4740);
and U5088 (N_5088,N_4512,N_4531);
or U5089 (N_5089,N_4832,N_4999);
nand U5090 (N_5090,N_4290,N_4816);
and U5091 (N_5091,N_4546,N_4805);
xor U5092 (N_5092,N_4978,N_4394);
xnor U5093 (N_5093,N_4204,N_4801);
nand U5094 (N_5094,N_4310,N_4324);
or U5095 (N_5095,N_4890,N_4022);
nor U5096 (N_5096,N_4678,N_4077);
nand U5097 (N_5097,N_4626,N_4905);
and U5098 (N_5098,N_4913,N_4378);
nor U5099 (N_5099,N_4343,N_4395);
nand U5100 (N_5100,N_4824,N_4446);
nand U5101 (N_5101,N_4367,N_4718);
nor U5102 (N_5102,N_4791,N_4538);
or U5103 (N_5103,N_4901,N_4669);
nor U5104 (N_5104,N_4587,N_4109);
or U5105 (N_5105,N_4187,N_4840);
or U5106 (N_5106,N_4406,N_4666);
nand U5107 (N_5107,N_4274,N_4519);
and U5108 (N_5108,N_4916,N_4939);
nand U5109 (N_5109,N_4528,N_4876);
or U5110 (N_5110,N_4984,N_4266);
nand U5111 (N_5111,N_4810,N_4543);
nand U5112 (N_5112,N_4822,N_4273);
nand U5113 (N_5113,N_4244,N_4193);
nand U5114 (N_5114,N_4893,N_4517);
nor U5115 (N_5115,N_4084,N_4553);
and U5116 (N_5116,N_4106,N_4642);
and U5117 (N_5117,N_4636,N_4032);
and U5118 (N_5118,N_4644,N_4447);
nand U5119 (N_5119,N_4102,N_4742);
or U5120 (N_5120,N_4171,N_4075);
xnor U5121 (N_5121,N_4284,N_4500);
or U5122 (N_5122,N_4753,N_4725);
nor U5123 (N_5123,N_4041,N_4898);
and U5124 (N_5124,N_4231,N_4622);
xnor U5125 (N_5125,N_4037,N_4312);
xor U5126 (N_5126,N_4686,N_4586);
nor U5127 (N_5127,N_4031,N_4474);
nand U5128 (N_5128,N_4007,N_4279);
nor U5129 (N_5129,N_4663,N_4424);
nor U5130 (N_5130,N_4572,N_4188);
nor U5131 (N_5131,N_4035,N_4366);
or U5132 (N_5132,N_4535,N_4108);
or U5133 (N_5133,N_4830,N_4823);
or U5134 (N_5134,N_4900,N_4359);
nor U5135 (N_5135,N_4507,N_4444);
xor U5136 (N_5136,N_4604,N_4116);
nand U5137 (N_5137,N_4611,N_4817);
or U5138 (N_5138,N_4610,N_4357);
and U5139 (N_5139,N_4195,N_4317);
xor U5140 (N_5140,N_4779,N_4230);
or U5141 (N_5141,N_4761,N_4219);
xor U5142 (N_5142,N_4731,N_4710);
and U5143 (N_5143,N_4192,N_4044);
nor U5144 (N_5144,N_4540,N_4522);
nand U5145 (N_5145,N_4813,N_4695);
nor U5146 (N_5146,N_4372,N_4379);
nand U5147 (N_5147,N_4687,N_4785);
and U5148 (N_5148,N_4976,N_4697);
nor U5149 (N_5149,N_4139,N_4202);
and U5150 (N_5150,N_4243,N_4480);
and U5151 (N_5151,N_4975,N_4078);
nand U5152 (N_5152,N_4256,N_4656);
nor U5153 (N_5153,N_4292,N_4302);
or U5154 (N_5154,N_4968,N_4054);
or U5155 (N_5155,N_4019,N_4289);
and U5156 (N_5156,N_4092,N_4162);
or U5157 (N_5157,N_4793,N_4240);
or U5158 (N_5158,N_4392,N_4503);
or U5159 (N_5159,N_4927,N_4739);
nor U5160 (N_5160,N_4479,N_4705);
or U5161 (N_5161,N_4340,N_4555);
nor U5162 (N_5162,N_4375,N_4030);
nor U5163 (N_5163,N_4719,N_4712);
nand U5164 (N_5164,N_4980,N_4218);
and U5165 (N_5165,N_4868,N_4170);
and U5166 (N_5166,N_4886,N_4514);
and U5167 (N_5167,N_4629,N_4143);
and U5168 (N_5168,N_4217,N_4238);
nand U5169 (N_5169,N_4869,N_4034);
or U5170 (N_5170,N_4495,N_4919);
or U5171 (N_5171,N_4621,N_4246);
or U5172 (N_5172,N_4386,N_4028);
and U5173 (N_5173,N_4743,N_4627);
nand U5174 (N_5174,N_4055,N_4631);
nand U5175 (N_5175,N_4578,N_4234);
or U5176 (N_5176,N_4433,N_4607);
nand U5177 (N_5177,N_4233,N_4168);
nand U5178 (N_5178,N_4842,N_4247);
or U5179 (N_5179,N_4369,N_4417);
or U5180 (N_5180,N_4967,N_4123);
nand U5181 (N_5181,N_4255,N_4914);
xnor U5182 (N_5182,N_4945,N_4398);
nor U5183 (N_5183,N_4690,N_4648);
or U5184 (N_5184,N_4175,N_4305);
or U5185 (N_5185,N_4185,N_4316);
nand U5186 (N_5186,N_4181,N_4095);
nand U5187 (N_5187,N_4481,N_4262);
and U5188 (N_5188,N_4459,N_4591);
nor U5189 (N_5189,N_4228,N_4241);
xor U5190 (N_5190,N_4497,N_4879);
and U5191 (N_5191,N_4133,N_4577);
or U5192 (N_5192,N_4201,N_4724);
and U5193 (N_5193,N_4458,N_4942);
or U5194 (N_5194,N_4936,N_4048);
nand U5195 (N_5195,N_4727,N_4649);
nor U5196 (N_5196,N_4025,N_4981);
and U5197 (N_5197,N_4672,N_4111);
and U5198 (N_5198,N_4925,N_4196);
nor U5199 (N_5199,N_4790,N_4923);
or U5200 (N_5200,N_4220,N_4935);
nand U5201 (N_5201,N_4216,N_4571);
or U5202 (N_5202,N_4707,N_4537);
and U5203 (N_5203,N_4397,N_4252);
nor U5204 (N_5204,N_4530,N_4608);
nand U5205 (N_5205,N_4026,N_4662);
xor U5206 (N_5206,N_4294,N_4485);
nor U5207 (N_5207,N_4576,N_4036);
or U5208 (N_5208,N_4269,N_4558);
nor U5209 (N_5209,N_4756,N_4411);
and U5210 (N_5210,N_4420,N_4042);
and U5211 (N_5211,N_4634,N_4061);
xor U5212 (N_5212,N_4426,N_4852);
nor U5213 (N_5213,N_4664,N_4545);
or U5214 (N_5214,N_4431,N_4723);
nand U5215 (N_5215,N_4891,N_4877);
and U5216 (N_5216,N_4757,N_4655);
nor U5217 (N_5217,N_4425,N_4836);
or U5218 (N_5218,N_4342,N_4870);
nand U5219 (N_5219,N_4899,N_4320);
and U5220 (N_5220,N_4564,N_4632);
nor U5221 (N_5221,N_4906,N_4131);
or U5222 (N_5222,N_4097,N_4152);
xnor U5223 (N_5223,N_4344,N_4829);
nor U5224 (N_5224,N_4915,N_4271);
or U5225 (N_5225,N_4871,N_4122);
and U5226 (N_5226,N_4982,N_4850);
xor U5227 (N_5227,N_4419,N_4937);
nor U5228 (N_5228,N_4683,N_4675);
or U5229 (N_5229,N_4760,N_4892);
nand U5230 (N_5230,N_4229,N_4800);
and U5231 (N_5231,N_4977,N_4205);
xnor U5232 (N_5232,N_4254,N_4265);
nand U5233 (N_5233,N_4768,N_4334);
or U5234 (N_5234,N_4853,N_4073);
and U5235 (N_5235,N_4066,N_4178);
and U5236 (N_5236,N_4146,N_4454);
nand U5237 (N_5237,N_4887,N_4554);
nand U5238 (N_5238,N_4293,N_4338);
nand U5239 (N_5239,N_4685,N_4039);
nand U5240 (N_5240,N_4548,N_4812);
or U5241 (N_5241,N_4755,N_4270);
nand U5242 (N_5242,N_4509,N_4221);
nand U5243 (N_5243,N_4014,N_4191);
nor U5244 (N_5244,N_4933,N_4858);
and U5245 (N_5245,N_4227,N_4064);
and U5246 (N_5246,N_4551,N_4733);
nor U5247 (N_5247,N_4318,N_4734);
or U5248 (N_5248,N_4797,N_4510);
or U5249 (N_5249,N_4478,N_4332);
or U5250 (N_5250,N_4401,N_4315);
nand U5251 (N_5251,N_4974,N_4065);
xor U5252 (N_5252,N_4597,N_4301);
and U5253 (N_5253,N_4156,N_4865);
nor U5254 (N_5254,N_4160,N_4380);
or U5255 (N_5255,N_4053,N_4348);
nor U5256 (N_5256,N_4396,N_4645);
and U5257 (N_5257,N_4285,N_4383);
xor U5258 (N_5258,N_4443,N_4619);
and U5259 (N_5259,N_4215,N_4506);
nand U5260 (N_5260,N_4658,N_4856);
nand U5261 (N_5261,N_4488,N_4747);
or U5262 (N_5262,N_4602,N_4169);
nand U5263 (N_5263,N_4166,N_4434);
nor U5264 (N_5264,N_4857,N_4953);
nand U5265 (N_5265,N_4282,N_4691);
or U5266 (N_5266,N_4814,N_4058);
and U5267 (N_5267,N_4911,N_4298);
nand U5268 (N_5268,N_4638,N_4941);
or U5269 (N_5269,N_4275,N_4407);
or U5270 (N_5270,N_4002,N_4934);
nand U5271 (N_5271,N_4703,N_4722);
nand U5272 (N_5272,N_4943,N_4260);
nand U5273 (N_5273,N_4455,N_4567);
and U5274 (N_5274,N_4605,N_4009);
or U5275 (N_5275,N_4056,N_4438);
and U5276 (N_5276,N_4737,N_4713);
and U5277 (N_5277,N_4501,N_4709);
nand U5278 (N_5278,N_4490,N_4151);
nor U5279 (N_5279,N_4786,N_4142);
nand U5280 (N_5280,N_4860,N_4399);
nand U5281 (N_5281,N_4112,N_4847);
nor U5282 (N_5282,N_4121,N_4671);
xor U5283 (N_5283,N_4998,N_4373);
nand U5284 (N_5284,N_4159,N_4700);
and U5285 (N_5285,N_4067,N_4594);
and U5286 (N_5286,N_4083,N_4613);
nand U5287 (N_5287,N_4759,N_4211);
nand U5288 (N_5288,N_4345,N_4382);
and U5289 (N_5289,N_4989,N_4556);
nand U5290 (N_5290,N_4831,N_4483);
nand U5291 (N_5291,N_4696,N_4932);
nor U5292 (N_5292,N_4321,N_4926);
or U5293 (N_5293,N_4237,N_4872);
nand U5294 (N_5294,N_4895,N_4336);
and U5295 (N_5295,N_4826,N_4792);
or U5296 (N_5296,N_4069,N_4726);
nand U5297 (N_5297,N_4281,N_4529);
nor U5298 (N_5298,N_4303,N_4498);
nor U5299 (N_5299,N_4706,N_4708);
nand U5300 (N_5300,N_4308,N_4190);
or U5301 (N_5301,N_4086,N_4432);
nor U5302 (N_5302,N_4052,N_4565);
and U5303 (N_5303,N_4620,N_4969);
or U5304 (N_5304,N_4807,N_4960);
nand U5305 (N_5305,N_4377,N_4463);
nand U5306 (N_5306,N_4570,N_4896);
or U5307 (N_5307,N_4803,N_4145);
nand U5308 (N_5308,N_4880,N_4261);
or U5309 (N_5309,N_4124,N_4593);
nand U5310 (N_5310,N_4063,N_4333);
nand U5311 (N_5311,N_4716,N_4149);
xor U5312 (N_5312,N_4527,N_4874);
or U5313 (N_5313,N_4466,N_4940);
nor U5314 (N_5314,N_4511,N_4469);
nor U5315 (N_5315,N_4214,N_4828);
nor U5316 (N_5316,N_4100,N_4337);
and U5317 (N_5317,N_4701,N_4885);
or U5318 (N_5318,N_4134,N_4389);
or U5319 (N_5319,N_4584,N_4125);
nand U5320 (N_5320,N_4862,N_4795);
or U5321 (N_5321,N_4226,N_4286);
or U5322 (N_5322,N_4020,N_4138);
and U5323 (N_5323,N_4117,N_4513);
xnor U5324 (N_5324,N_4005,N_4153);
or U5325 (N_5325,N_4904,N_4643);
and U5326 (N_5326,N_4177,N_4264);
nand U5327 (N_5327,N_4624,N_4251);
nand U5328 (N_5328,N_4728,N_4400);
nor U5329 (N_5329,N_4949,N_4616);
nor U5330 (N_5330,N_4987,N_4952);
or U5331 (N_5331,N_4016,N_4405);
or U5332 (N_5332,N_4574,N_4566);
and U5333 (N_5333,N_4183,N_4403);
xnor U5334 (N_5334,N_4347,N_4688);
and U5335 (N_5335,N_4472,N_4329);
nor U5336 (N_5336,N_4000,N_4654);
nor U5337 (N_5337,N_4928,N_4135);
and U5338 (N_5338,N_4588,N_4798);
nand U5339 (N_5339,N_4010,N_4881);
and U5340 (N_5340,N_4043,N_4435);
nor U5341 (N_5341,N_4429,N_4802);
xnor U5342 (N_5342,N_4921,N_4922);
nor U5343 (N_5343,N_4300,N_4128);
nand U5344 (N_5344,N_4299,N_4250);
and U5345 (N_5345,N_4361,N_4351);
nor U5346 (N_5346,N_4418,N_4520);
nor U5347 (N_5347,N_4991,N_4615);
or U5348 (N_5348,N_4094,N_4068);
nand U5349 (N_5349,N_4288,N_4222);
and U5350 (N_5350,N_4954,N_4635);
and U5351 (N_5351,N_4387,N_4679);
and U5352 (N_5352,N_4208,N_4462);
nor U5353 (N_5353,N_4148,N_4582);
nor U5354 (N_5354,N_4956,N_4057);
or U5355 (N_5355,N_4465,N_4809);
or U5356 (N_5356,N_4071,N_4573);
and U5357 (N_5357,N_4360,N_4197);
and U5358 (N_5358,N_4667,N_4464);
and U5359 (N_5359,N_4778,N_4550);
nand U5360 (N_5360,N_4096,N_4781);
nor U5361 (N_5361,N_4818,N_4851);
nand U5362 (N_5362,N_4179,N_4533);
or U5363 (N_5363,N_4017,N_4875);
nand U5364 (N_5364,N_4855,N_4557);
and U5365 (N_5365,N_4754,N_4721);
and U5366 (N_5366,N_4349,N_4090);
nand U5367 (N_5367,N_4163,N_4883);
nor U5368 (N_5368,N_4848,N_4410);
nand U5369 (N_5369,N_4625,N_4931);
or U5370 (N_5370,N_4306,N_4408);
or U5371 (N_5371,N_4951,N_4325);
nor U5372 (N_5372,N_4689,N_4319);
nor U5373 (N_5373,N_4103,N_4841);
nor U5374 (N_5374,N_4126,N_4456);
nand U5375 (N_5375,N_4682,N_4788);
nand U5376 (N_5376,N_4199,N_4532);
and U5377 (N_5377,N_4979,N_4001);
and U5378 (N_5378,N_4313,N_4844);
and U5379 (N_5379,N_4356,N_4674);
and U5380 (N_5380,N_4213,N_4846);
or U5381 (N_5381,N_4692,N_4948);
nand U5382 (N_5382,N_4235,N_4427);
nor U5383 (N_5383,N_4207,N_4964);
or U5384 (N_5384,N_4088,N_4820);
or U5385 (N_5385,N_4575,N_4355);
nand U5386 (N_5386,N_4966,N_4539);
nor U5387 (N_5387,N_4390,N_4223);
and U5388 (N_5388,N_4180,N_4012);
and U5389 (N_5389,N_4815,N_4487);
nor U5390 (N_5390,N_4113,N_4772);
or U5391 (N_5391,N_4694,N_4849);
nand U5392 (N_5392,N_4104,N_4295);
nand U5393 (N_5393,N_4603,N_4172);
xnor U5394 (N_5394,N_4568,N_4060);
nor U5395 (N_5395,N_4714,N_4477);
and U5396 (N_5396,N_4698,N_4661);
xor U5397 (N_5397,N_4085,N_4049);
nand U5398 (N_5398,N_4751,N_4309);
nor U5399 (N_5399,N_4393,N_4720);
nor U5400 (N_5400,N_4307,N_4590);
and U5401 (N_5401,N_4523,N_4526);
nand U5402 (N_5402,N_4354,N_4651);
and U5403 (N_5403,N_4422,N_4453);
or U5404 (N_5404,N_4115,N_4011);
nor U5405 (N_5405,N_4182,N_4944);
nand U5406 (N_5406,N_4374,N_4614);
nand U5407 (N_5407,N_4888,N_4364);
nor U5408 (N_5408,N_4062,N_4878);
nor U5409 (N_5409,N_4867,N_4147);
nand U5410 (N_5410,N_4673,N_4580);
and U5411 (N_5411,N_4782,N_4837);
and U5412 (N_5412,N_4961,N_4741);
xor U5413 (N_5413,N_4093,N_4653);
and U5414 (N_5414,N_4047,N_4947);
nor U5415 (N_5415,N_4633,N_4677);
xor U5416 (N_5416,N_4283,N_4245);
and U5417 (N_5417,N_4783,N_4297);
or U5418 (N_5418,N_4515,N_4448);
nand U5419 (N_5419,N_4484,N_4473);
nand U5420 (N_5420,N_4144,N_4562);
nor U5421 (N_5421,N_4263,N_4209);
nor U5422 (N_5422,N_4859,N_4368);
and U5423 (N_5423,N_4589,N_4657);
xor U5424 (N_5424,N_4647,N_4224);
and U5425 (N_5425,N_4560,N_4541);
or U5426 (N_5426,N_4729,N_4323);
nand U5427 (N_5427,N_4518,N_4110);
or U5428 (N_5428,N_4930,N_4091);
or U5429 (N_5429,N_4008,N_4780);
or U5430 (N_5430,N_4971,N_4164);
nor U5431 (N_5431,N_4983,N_4882);
or U5432 (N_5432,N_4476,N_4789);
nand U5433 (N_5433,N_4819,N_4771);
xor U5434 (N_5434,N_4652,N_4521);
nor U5435 (N_5435,N_4416,N_4105);
nor U5436 (N_5436,N_4717,N_4440);
nor U5437 (N_5437,N_4492,N_4970);
nand U5438 (N_5438,N_4460,N_4762);
nor U5439 (N_5439,N_4076,N_4327);
nand U5440 (N_5440,N_4711,N_4628);
nor U5441 (N_5441,N_4155,N_4412);
xnor U5442 (N_5442,N_4024,N_4775);
or U5443 (N_5443,N_4972,N_4912);
and U5444 (N_5444,N_4598,N_4051);
or U5445 (N_5445,N_4370,N_4212);
nor U5446 (N_5446,N_4045,N_4600);
xnor U5447 (N_5447,N_4003,N_4524);
nor U5448 (N_5448,N_4660,N_4838);
nand U5449 (N_5449,N_4902,N_4766);
and U5450 (N_5450,N_4081,N_4268);
nor U5451 (N_5451,N_4732,N_4693);
xnor U5452 (N_5452,N_4079,N_4362);
and U5453 (N_5453,N_4470,N_4436);
nand U5454 (N_5454,N_4391,N_4141);
and U5455 (N_5455,N_4276,N_4950);
and U5456 (N_5456,N_4225,N_4617);
or U5457 (N_5457,N_4004,N_4015);
or U5458 (N_5458,N_4730,N_4985);
nand U5459 (N_5459,N_4843,N_4744);
or U5460 (N_5460,N_4563,N_4821);
nor U5461 (N_5461,N_4884,N_4326);
nand U5462 (N_5462,N_4763,N_4988);
and U5463 (N_5463,N_4845,N_4749);
or U5464 (N_5464,N_4363,N_4894);
or U5465 (N_5465,N_4167,N_4006);
nand U5466 (N_5466,N_4475,N_4161);
and U5467 (N_5467,N_4559,N_4499);
nor U5468 (N_5468,N_4358,N_4646);
and U5469 (N_5469,N_4702,N_4314);
nor U5470 (N_5470,N_4132,N_4715);
nand U5471 (N_5471,N_4384,N_4735);
or U5472 (N_5472,N_4993,N_4258);
nor U5473 (N_5473,N_4561,N_4232);
or U5474 (N_5474,N_4676,N_4699);
nand U5475 (N_5475,N_4018,N_4986);
xor U5476 (N_5476,N_4864,N_4277);
xor U5477 (N_5477,N_4119,N_4908);
or U5478 (N_5478,N_4639,N_4040);
nor U5479 (N_5479,N_4013,N_4547);
nand U5480 (N_5480,N_4920,N_4623);
and U5481 (N_5481,N_4154,N_4955);
nand U5482 (N_5482,N_4186,N_4415);
and U5483 (N_5483,N_4903,N_4599);
nand U5484 (N_5484,N_4114,N_4257);
nand U5485 (N_5485,N_4505,N_4668);
and U5486 (N_5486,N_4502,N_4784);
or U5487 (N_5487,N_4959,N_4767);
and U5488 (N_5488,N_4569,N_4774);
or U5489 (N_5489,N_4080,N_4834);
or U5490 (N_5490,N_4909,N_4365);
and U5491 (N_5491,N_4758,N_4804);
or U5492 (N_5492,N_4525,N_4854);
nand U5493 (N_5493,N_4457,N_4736);
xnor U5494 (N_5494,N_4249,N_4738);
and U5495 (N_5495,N_4267,N_4194);
or U5496 (N_5496,N_4990,N_4098);
nor U5497 (N_5497,N_4341,N_4449);
nor U5498 (N_5498,N_4414,N_4287);
xnor U5499 (N_5499,N_4680,N_4504);
and U5500 (N_5500,N_4536,N_4680);
and U5501 (N_5501,N_4957,N_4777);
nand U5502 (N_5502,N_4552,N_4081);
nand U5503 (N_5503,N_4713,N_4196);
or U5504 (N_5504,N_4982,N_4666);
or U5505 (N_5505,N_4715,N_4278);
or U5506 (N_5506,N_4240,N_4179);
and U5507 (N_5507,N_4177,N_4978);
or U5508 (N_5508,N_4990,N_4507);
nor U5509 (N_5509,N_4630,N_4031);
nand U5510 (N_5510,N_4365,N_4402);
or U5511 (N_5511,N_4205,N_4057);
xor U5512 (N_5512,N_4050,N_4059);
xnor U5513 (N_5513,N_4474,N_4550);
nor U5514 (N_5514,N_4952,N_4440);
nand U5515 (N_5515,N_4664,N_4295);
xnor U5516 (N_5516,N_4280,N_4370);
xor U5517 (N_5517,N_4876,N_4764);
nor U5518 (N_5518,N_4670,N_4796);
nor U5519 (N_5519,N_4488,N_4258);
or U5520 (N_5520,N_4894,N_4102);
and U5521 (N_5521,N_4833,N_4432);
and U5522 (N_5522,N_4234,N_4989);
nand U5523 (N_5523,N_4522,N_4670);
and U5524 (N_5524,N_4104,N_4692);
nand U5525 (N_5525,N_4770,N_4863);
nand U5526 (N_5526,N_4715,N_4382);
and U5527 (N_5527,N_4260,N_4163);
or U5528 (N_5528,N_4375,N_4239);
or U5529 (N_5529,N_4220,N_4197);
or U5530 (N_5530,N_4916,N_4001);
or U5531 (N_5531,N_4376,N_4519);
xnor U5532 (N_5532,N_4130,N_4999);
xor U5533 (N_5533,N_4923,N_4753);
xor U5534 (N_5534,N_4879,N_4301);
nor U5535 (N_5535,N_4815,N_4461);
and U5536 (N_5536,N_4067,N_4342);
nor U5537 (N_5537,N_4940,N_4430);
and U5538 (N_5538,N_4618,N_4696);
nor U5539 (N_5539,N_4781,N_4195);
xor U5540 (N_5540,N_4030,N_4352);
nand U5541 (N_5541,N_4050,N_4721);
nor U5542 (N_5542,N_4991,N_4403);
nor U5543 (N_5543,N_4807,N_4338);
nor U5544 (N_5544,N_4120,N_4364);
and U5545 (N_5545,N_4324,N_4297);
and U5546 (N_5546,N_4641,N_4336);
or U5547 (N_5547,N_4837,N_4279);
or U5548 (N_5548,N_4747,N_4304);
nor U5549 (N_5549,N_4179,N_4616);
or U5550 (N_5550,N_4114,N_4825);
nand U5551 (N_5551,N_4180,N_4218);
nand U5552 (N_5552,N_4129,N_4058);
and U5553 (N_5553,N_4846,N_4318);
and U5554 (N_5554,N_4952,N_4692);
or U5555 (N_5555,N_4539,N_4887);
nand U5556 (N_5556,N_4792,N_4693);
xnor U5557 (N_5557,N_4619,N_4400);
nand U5558 (N_5558,N_4283,N_4681);
nor U5559 (N_5559,N_4848,N_4078);
nand U5560 (N_5560,N_4326,N_4285);
nand U5561 (N_5561,N_4988,N_4802);
and U5562 (N_5562,N_4709,N_4685);
or U5563 (N_5563,N_4101,N_4822);
and U5564 (N_5564,N_4566,N_4981);
nor U5565 (N_5565,N_4363,N_4777);
or U5566 (N_5566,N_4896,N_4200);
nand U5567 (N_5567,N_4010,N_4128);
and U5568 (N_5568,N_4342,N_4422);
or U5569 (N_5569,N_4630,N_4909);
and U5570 (N_5570,N_4561,N_4343);
and U5571 (N_5571,N_4340,N_4852);
nor U5572 (N_5572,N_4253,N_4417);
or U5573 (N_5573,N_4937,N_4753);
nor U5574 (N_5574,N_4526,N_4689);
or U5575 (N_5575,N_4439,N_4159);
nor U5576 (N_5576,N_4600,N_4340);
nor U5577 (N_5577,N_4770,N_4432);
nand U5578 (N_5578,N_4199,N_4978);
nor U5579 (N_5579,N_4173,N_4485);
and U5580 (N_5580,N_4466,N_4507);
or U5581 (N_5581,N_4931,N_4048);
or U5582 (N_5582,N_4694,N_4860);
or U5583 (N_5583,N_4834,N_4214);
nand U5584 (N_5584,N_4519,N_4241);
or U5585 (N_5585,N_4396,N_4687);
and U5586 (N_5586,N_4271,N_4725);
or U5587 (N_5587,N_4678,N_4469);
nand U5588 (N_5588,N_4968,N_4371);
nand U5589 (N_5589,N_4854,N_4006);
or U5590 (N_5590,N_4896,N_4907);
and U5591 (N_5591,N_4406,N_4427);
nand U5592 (N_5592,N_4985,N_4071);
nor U5593 (N_5593,N_4342,N_4186);
and U5594 (N_5594,N_4369,N_4148);
nor U5595 (N_5595,N_4972,N_4890);
xor U5596 (N_5596,N_4889,N_4496);
nand U5597 (N_5597,N_4427,N_4740);
nand U5598 (N_5598,N_4238,N_4519);
and U5599 (N_5599,N_4856,N_4144);
nand U5600 (N_5600,N_4257,N_4031);
nor U5601 (N_5601,N_4928,N_4132);
and U5602 (N_5602,N_4428,N_4945);
nor U5603 (N_5603,N_4756,N_4581);
nor U5604 (N_5604,N_4559,N_4183);
nor U5605 (N_5605,N_4275,N_4342);
nor U5606 (N_5606,N_4384,N_4993);
or U5607 (N_5607,N_4471,N_4938);
nor U5608 (N_5608,N_4966,N_4737);
nor U5609 (N_5609,N_4637,N_4044);
nor U5610 (N_5610,N_4732,N_4267);
and U5611 (N_5611,N_4390,N_4277);
or U5612 (N_5612,N_4611,N_4099);
and U5613 (N_5613,N_4252,N_4912);
or U5614 (N_5614,N_4937,N_4246);
nand U5615 (N_5615,N_4540,N_4223);
or U5616 (N_5616,N_4508,N_4641);
nor U5617 (N_5617,N_4538,N_4524);
nand U5618 (N_5618,N_4592,N_4146);
nand U5619 (N_5619,N_4522,N_4074);
nand U5620 (N_5620,N_4189,N_4193);
nor U5621 (N_5621,N_4926,N_4985);
nor U5622 (N_5622,N_4946,N_4085);
and U5623 (N_5623,N_4831,N_4999);
xor U5624 (N_5624,N_4623,N_4098);
or U5625 (N_5625,N_4634,N_4773);
nand U5626 (N_5626,N_4907,N_4117);
and U5627 (N_5627,N_4770,N_4608);
nor U5628 (N_5628,N_4645,N_4844);
and U5629 (N_5629,N_4768,N_4806);
and U5630 (N_5630,N_4514,N_4263);
nand U5631 (N_5631,N_4565,N_4385);
and U5632 (N_5632,N_4541,N_4334);
and U5633 (N_5633,N_4782,N_4723);
and U5634 (N_5634,N_4362,N_4599);
nor U5635 (N_5635,N_4049,N_4280);
nor U5636 (N_5636,N_4525,N_4129);
nor U5637 (N_5637,N_4638,N_4242);
nand U5638 (N_5638,N_4826,N_4262);
and U5639 (N_5639,N_4245,N_4661);
and U5640 (N_5640,N_4983,N_4803);
and U5641 (N_5641,N_4026,N_4086);
or U5642 (N_5642,N_4260,N_4876);
nor U5643 (N_5643,N_4042,N_4637);
or U5644 (N_5644,N_4646,N_4170);
and U5645 (N_5645,N_4695,N_4749);
or U5646 (N_5646,N_4590,N_4165);
and U5647 (N_5647,N_4631,N_4141);
and U5648 (N_5648,N_4262,N_4603);
nand U5649 (N_5649,N_4052,N_4875);
or U5650 (N_5650,N_4055,N_4649);
and U5651 (N_5651,N_4023,N_4408);
or U5652 (N_5652,N_4111,N_4142);
nand U5653 (N_5653,N_4463,N_4054);
or U5654 (N_5654,N_4623,N_4460);
xnor U5655 (N_5655,N_4215,N_4796);
and U5656 (N_5656,N_4677,N_4355);
nor U5657 (N_5657,N_4823,N_4377);
nand U5658 (N_5658,N_4167,N_4526);
and U5659 (N_5659,N_4846,N_4756);
nand U5660 (N_5660,N_4316,N_4799);
nor U5661 (N_5661,N_4394,N_4824);
nand U5662 (N_5662,N_4866,N_4947);
or U5663 (N_5663,N_4657,N_4348);
and U5664 (N_5664,N_4240,N_4455);
or U5665 (N_5665,N_4634,N_4606);
nor U5666 (N_5666,N_4418,N_4901);
or U5667 (N_5667,N_4348,N_4007);
or U5668 (N_5668,N_4278,N_4787);
xor U5669 (N_5669,N_4045,N_4261);
or U5670 (N_5670,N_4837,N_4230);
nand U5671 (N_5671,N_4492,N_4500);
nand U5672 (N_5672,N_4016,N_4645);
nand U5673 (N_5673,N_4880,N_4492);
or U5674 (N_5674,N_4556,N_4652);
nor U5675 (N_5675,N_4128,N_4353);
nor U5676 (N_5676,N_4816,N_4139);
nand U5677 (N_5677,N_4438,N_4370);
nor U5678 (N_5678,N_4282,N_4374);
nand U5679 (N_5679,N_4734,N_4024);
and U5680 (N_5680,N_4633,N_4386);
nor U5681 (N_5681,N_4512,N_4532);
nor U5682 (N_5682,N_4152,N_4612);
nor U5683 (N_5683,N_4307,N_4214);
nand U5684 (N_5684,N_4098,N_4000);
and U5685 (N_5685,N_4159,N_4135);
or U5686 (N_5686,N_4198,N_4727);
and U5687 (N_5687,N_4885,N_4175);
nor U5688 (N_5688,N_4708,N_4577);
xnor U5689 (N_5689,N_4752,N_4374);
nor U5690 (N_5690,N_4836,N_4937);
nor U5691 (N_5691,N_4957,N_4881);
and U5692 (N_5692,N_4105,N_4898);
and U5693 (N_5693,N_4336,N_4593);
nor U5694 (N_5694,N_4259,N_4784);
nand U5695 (N_5695,N_4791,N_4421);
nor U5696 (N_5696,N_4289,N_4618);
nor U5697 (N_5697,N_4464,N_4200);
xor U5698 (N_5698,N_4145,N_4250);
and U5699 (N_5699,N_4106,N_4977);
nand U5700 (N_5700,N_4477,N_4448);
nor U5701 (N_5701,N_4065,N_4943);
xor U5702 (N_5702,N_4914,N_4101);
and U5703 (N_5703,N_4329,N_4450);
or U5704 (N_5704,N_4809,N_4078);
nand U5705 (N_5705,N_4427,N_4187);
nor U5706 (N_5706,N_4086,N_4846);
nor U5707 (N_5707,N_4563,N_4170);
nand U5708 (N_5708,N_4702,N_4746);
nand U5709 (N_5709,N_4093,N_4955);
nor U5710 (N_5710,N_4401,N_4430);
xor U5711 (N_5711,N_4750,N_4531);
or U5712 (N_5712,N_4538,N_4999);
and U5713 (N_5713,N_4332,N_4119);
or U5714 (N_5714,N_4400,N_4343);
nor U5715 (N_5715,N_4548,N_4409);
nor U5716 (N_5716,N_4831,N_4707);
nand U5717 (N_5717,N_4311,N_4009);
nand U5718 (N_5718,N_4839,N_4667);
nor U5719 (N_5719,N_4654,N_4987);
nand U5720 (N_5720,N_4827,N_4935);
and U5721 (N_5721,N_4959,N_4500);
and U5722 (N_5722,N_4086,N_4214);
or U5723 (N_5723,N_4707,N_4337);
nor U5724 (N_5724,N_4470,N_4489);
or U5725 (N_5725,N_4433,N_4421);
nand U5726 (N_5726,N_4312,N_4024);
or U5727 (N_5727,N_4490,N_4441);
nor U5728 (N_5728,N_4721,N_4140);
nor U5729 (N_5729,N_4081,N_4784);
or U5730 (N_5730,N_4946,N_4001);
xor U5731 (N_5731,N_4099,N_4955);
xor U5732 (N_5732,N_4060,N_4553);
and U5733 (N_5733,N_4399,N_4854);
nand U5734 (N_5734,N_4872,N_4232);
xnor U5735 (N_5735,N_4500,N_4152);
xor U5736 (N_5736,N_4693,N_4703);
nand U5737 (N_5737,N_4557,N_4587);
or U5738 (N_5738,N_4529,N_4981);
nand U5739 (N_5739,N_4067,N_4249);
nand U5740 (N_5740,N_4241,N_4293);
or U5741 (N_5741,N_4993,N_4171);
or U5742 (N_5742,N_4251,N_4968);
nand U5743 (N_5743,N_4917,N_4306);
and U5744 (N_5744,N_4342,N_4136);
and U5745 (N_5745,N_4453,N_4654);
nor U5746 (N_5746,N_4096,N_4329);
or U5747 (N_5747,N_4734,N_4468);
or U5748 (N_5748,N_4795,N_4455);
and U5749 (N_5749,N_4162,N_4852);
nand U5750 (N_5750,N_4033,N_4098);
and U5751 (N_5751,N_4485,N_4033);
nand U5752 (N_5752,N_4839,N_4550);
nor U5753 (N_5753,N_4089,N_4055);
and U5754 (N_5754,N_4222,N_4321);
and U5755 (N_5755,N_4993,N_4992);
nand U5756 (N_5756,N_4125,N_4497);
and U5757 (N_5757,N_4876,N_4620);
nor U5758 (N_5758,N_4776,N_4053);
xnor U5759 (N_5759,N_4777,N_4287);
or U5760 (N_5760,N_4881,N_4268);
nand U5761 (N_5761,N_4394,N_4973);
nor U5762 (N_5762,N_4484,N_4614);
nor U5763 (N_5763,N_4250,N_4846);
and U5764 (N_5764,N_4773,N_4260);
and U5765 (N_5765,N_4408,N_4045);
and U5766 (N_5766,N_4719,N_4206);
or U5767 (N_5767,N_4730,N_4254);
and U5768 (N_5768,N_4354,N_4014);
xnor U5769 (N_5769,N_4571,N_4247);
xor U5770 (N_5770,N_4654,N_4328);
or U5771 (N_5771,N_4986,N_4758);
or U5772 (N_5772,N_4916,N_4507);
or U5773 (N_5773,N_4133,N_4118);
or U5774 (N_5774,N_4349,N_4884);
nand U5775 (N_5775,N_4442,N_4910);
nor U5776 (N_5776,N_4506,N_4764);
nand U5777 (N_5777,N_4601,N_4559);
xor U5778 (N_5778,N_4496,N_4562);
nor U5779 (N_5779,N_4113,N_4366);
nand U5780 (N_5780,N_4312,N_4109);
nand U5781 (N_5781,N_4402,N_4048);
or U5782 (N_5782,N_4641,N_4117);
xor U5783 (N_5783,N_4322,N_4741);
nand U5784 (N_5784,N_4217,N_4017);
or U5785 (N_5785,N_4182,N_4489);
and U5786 (N_5786,N_4825,N_4623);
or U5787 (N_5787,N_4617,N_4571);
and U5788 (N_5788,N_4115,N_4164);
nand U5789 (N_5789,N_4619,N_4644);
or U5790 (N_5790,N_4437,N_4882);
nand U5791 (N_5791,N_4413,N_4960);
and U5792 (N_5792,N_4205,N_4559);
and U5793 (N_5793,N_4806,N_4740);
nor U5794 (N_5794,N_4146,N_4043);
nand U5795 (N_5795,N_4433,N_4617);
and U5796 (N_5796,N_4379,N_4775);
nand U5797 (N_5797,N_4001,N_4282);
and U5798 (N_5798,N_4218,N_4596);
nor U5799 (N_5799,N_4263,N_4240);
and U5800 (N_5800,N_4815,N_4625);
or U5801 (N_5801,N_4581,N_4397);
nand U5802 (N_5802,N_4565,N_4006);
nand U5803 (N_5803,N_4487,N_4792);
or U5804 (N_5804,N_4496,N_4125);
and U5805 (N_5805,N_4173,N_4448);
nor U5806 (N_5806,N_4075,N_4553);
nand U5807 (N_5807,N_4735,N_4389);
or U5808 (N_5808,N_4998,N_4718);
and U5809 (N_5809,N_4440,N_4213);
and U5810 (N_5810,N_4201,N_4004);
and U5811 (N_5811,N_4252,N_4029);
nand U5812 (N_5812,N_4384,N_4876);
and U5813 (N_5813,N_4952,N_4616);
or U5814 (N_5814,N_4860,N_4466);
xnor U5815 (N_5815,N_4807,N_4378);
nor U5816 (N_5816,N_4951,N_4392);
or U5817 (N_5817,N_4929,N_4393);
nand U5818 (N_5818,N_4638,N_4682);
nor U5819 (N_5819,N_4172,N_4865);
nand U5820 (N_5820,N_4718,N_4324);
xnor U5821 (N_5821,N_4660,N_4692);
xnor U5822 (N_5822,N_4597,N_4321);
nand U5823 (N_5823,N_4569,N_4241);
or U5824 (N_5824,N_4608,N_4749);
nor U5825 (N_5825,N_4628,N_4663);
or U5826 (N_5826,N_4895,N_4053);
xor U5827 (N_5827,N_4518,N_4351);
nor U5828 (N_5828,N_4397,N_4341);
nand U5829 (N_5829,N_4725,N_4324);
or U5830 (N_5830,N_4170,N_4884);
and U5831 (N_5831,N_4440,N_4311);
or U5832 (N_5832,N_4962,N_4878);
and U5833 (N_5833,N_4077,N_4960);
xnor U5834 (N_5834,N_4142,N_4780);
and U5835 (N_5835,N_4327,N_4340);
nor U5836 (N_5836,N_4111,N_4691);
and U5837 (N_5837,N_4999,N_4151);
and U5838 (N_5838,N_4772,N_4741);
and U5839 (N_5839,N_4541,N_4227);
and U5840 (N_5840,N_4312,N_4540);
nor U5841 (N_5841,N_4755,N_4126);
and U5842 (N_5842,N_4157,N_4815);
nand U5843 (N_5843,N_4046,N_4852);
and U5844 (N_5844,N_4435,N_4458);
and U5845 (N_5845,N_4143,N_4625);
or U5846 (N_5846,N_4785,N_4066);
nor U5847 (N_5847,N_4620,N_4007);
or U5848 (N_5848,N_4468,N_4852);
and U5849 (N_5849,N_4174,N_4331);
nor U5850 (N_5850,N_4459,N_4297);
nor U5851 (N_5851,N_4315,N_4112);
or U5852 (N_5852,N_4469,N_4155);
and U5853 (N_5853,N_4127,N_4535);
nand U5854 (N_5854,N_4129,N_4895);
or U5855 (N_5855,N_4930,N_4842);
and U5856 (N_5856,N_4244,N_4191);
nor U5857 (N_5857,N_4372,N_4536);
xnor U5858 (N_5858,N_4298,N_4408);
and U5859 (N_5859,N_4342,N_4492);
or U5860 (N_5860,N_4903,N_4317);
xnor U5861 (N_5861,N_4754,N_4681);
nand U5862 (N_5862,N_4223,N_4535);
or U5863 (N_5863,N_4636,N_4493);
nor U5864 (N_5864,N_4732,N_4271);
nand U5865 (N_5865,N_4559,N_4843);
nand U5866 (N_5866,N_4074,N_4117);
xor U5867 (N_5867,N_4349,N_4380);
xor U5868 (N_5868,N_4453,N_4822);
nand U5869 (N_5869,N_4093,N_4550);
nand U5870 (N_5870,N_4227,N_4568);
and U5871 (N_5871,N_4674,N_4727);
nor U5872 (N_5872,N_4672,N_4927);
nand U5873 (N_5873,N_4024,N_4055);
nand U5874 (N_5874,N_4604,N_4628);
and U5875 (N_5875,N_4815,N_4041);
or U5876 (N_5876,N_4011,N_4683);
nand U5877 (N_5877,N_4138,N_4754);
nand U5878 (N_5878,N_4933,N_4478);
or U5879 (N_5879,N_4002,N_4904);
xnor U5880 (N_5880,N_4350,N_4949);
nor U5881 (N_5881,N_4874,N_4677);
xor U5882 (N_5882,N_4875,N_4502);
nand U5883 (N_5883,N_4032,N_4299);
and U5884 (N_5884,N_4608,N_4321);
and U5885 (N_5885,N_4965,N_4517);
or U5886 (N_5886,N_4455,N_4297);
or U5887 (N_5887,N_4227,N_4052);
or U5888 (N_5888,N_4487,N_4188);
or U5889 (N_5889,N_4001,N_4063);
or U5890 (N_5890,N_4847,N_4546);
and U5891 (N_5891,N_4426,N_4274);
or U5892 (N_5892,N_4963,N_4143);
nand U5893 (N_5893,N_4858,N_4413);
xor U5894 (N_5894,N_4414,N_4590);
xnor U5895 (N_5895,N_4883,N_4946);
and U5896 (N_5896,N_4222,N_4514);
or U5897 (N_5897,N_4965,N_4888);
xor U5898 (N_5898,N_4319,N_4171);
nand U5899 (N_5899,N_4715,N_4554);
or U5900 (N_5900,N_4384,N_4581);
nor U5901 (N_5901,N_4942,N_4596);
or U5902 (N_5902,N_4905,N_4162);
nor U5903 (N_5903,N_4934,N_4359);
nand U5904 (N_5904,N_4487,N_4100);
and U5905 (N_5905,N_4285,N_4651);
xor U5906 (N_5906,N_4595,N_4360);
or U5907 (N_5907,N_4691,N_4893);
nand U5908 (N_5908,N_4469,N_4744);
nor U5909 (N_5909,N_4452,N_4415);
or U5910 (N_5910,N_4825,N_4642);
or U5911 (N_5911,N_4091,N_4266);
or U5912 (N_5912,N_4432,N_4868);
and U5913 (N_5913,N_4831,N_4196);
or U5914 (N_5914,N_4283,N_4984);
nand U5915 (N_5915,N_4517,N_4662);
or U5916 (N_5916,N_4969,N_4520);
nor U5917 (N_5917,N_4886,N_4538);
nand U5918 (N_5918,N_4986,N_4405);
nor U5919 (N_5919,N_4893,N_4037);
or U5920 (N_5920,N_4597,N_4837);
nand U5921 (N_5921,N_4637,N_4879);
nand U5922 (N_5922,N_4398,N_4925);
and U5923 (N_5923,N_4484,N_4727);
and U5924 (N_5924,N_4293,N_4968);
xnor U5925 (N_5925,N_4161,N_4063);
and U5926 (N_5926,N_4427,N_4364);
or U5927 (N_5927,N_4043,N_4625);
or U5928 (N_5928,N_4593,N_4076);
and U5929 (N_5929,N_4535,N_4675);
or U5930 (N_5930,N_4330,N_4003);
nand U5931 (N_5931,N_4439,N_4711);
nand U5932 (N_5932,N_4959,N_4659);
or U5933 (N_5933,N_4836,N_4944);
nand U5934 (N_5934,N_4766,N_4778);
nand U5935 (N_5935,N_4631,N_4166);
or U5936 (N_5936,N_4420,N_4894);
or U5937 (N_5937,N_4994,N_4130);
nand U5938 (N_5938,N_4481,N_4905);
and U5939 (N_5939,N_4862,N_4081);
and U5940 (N_5940,N_4619,N_4034);
and U5941 (N_5941,N_4897,N_4624);
nand U5942 (N_5942,N_4030,N_4978);
xor U5943 (N_5943,N_4876,N_4828);
nor U5944 (N_5944,N_4994,N_4029);
nor U5945 (N_5945,N_4195,N_4089);
nor U5946 (N_5946,N_4860,N_4287);
xnor U5947 (N_5947,N_4240,N_4848);
nand U5948 (N_5948,N_4607,N_4373);
nor U5949 (N_5949,N_4959,N_4183);
or U5950 (N_5950,N_4796,N_4084);
nand U5951 (N_5951,N_4725,N_4819);
or U5952 (N_5952,N_4725,N_4210);
nor U5953 (N_5953,N_4256,N_4977);
and U5954 (N_5954,N_4575,N_4191);
and U5955 (N_5955,N_4762,N_4375);
xnor U5956 (N_5956,N_4640,N_4354);
or U5957 (N_5957,N_4590,N_4043);
nand U5958 (N_5958,N_4386,N_4734);
or U5959 (N_5959,N_4713,N_4008);
and U5960 (N_5960,N_4217,N_4549);
or U5961 (N_5961,N_4331,N_4081);
nand U5962 (N_5962,N_4730,N_4032);
or U5963 (N_5963,N_4873,N_4942);
or U5964 (N_5964,N_4933,N_4837);
and U5965 (N_5965,N_4565,N_4891);
nor U5966 (N_5966,N_4390,N_4944);
or U5967 (N_5967,N_4270,N_4981);
or U5968 (N_5968,N_4336,N_4603);
nor U5969 (N_5969,N_4088,N_4262);
nand U5970 (N_5970,N_4808,N_4576);
xor U5971 (N_5971,N_4589,N_4272);
and U5972 (N_5972,N_4008,N_4874);
nand U5973 (N_5973,N_4839,N_4094);
nor U5974 (N_5974,N_4939,N_4235);
nand U5975 (N_5975,N_4332,N_4429);
and U5976 (N_5976,N_4794,N_4015);
nand U5977 (N_5977,N_4877,N_4627);
nand U5978 (N_5978,N_4236,N_4606);
nor U5979 (N_5979,N_4960,N_4196);
nand U5980 (N_5980,N_4163,N_4633);
or U5981 (N_5981,N_4103,N_4851);
nand U5982 (N_5982,N_4621,N_4910);
nand U5983 (N_5983,N_4897,N_4028);
nand U5984 (N_5984,N_4215,N_4570);
nor U5985 (N_5985,N_4442,N_4870);
xnor U5986 (N_5986,N_4843,N_4747);
xnor U5987 (N_5987,N_4981,N_4850);
or U5988 (N_5988,N_4734,N_4032);
and U5989 (N_5989,N_4062,N_4600);
nand U5990 (N_5990,N_4755,N_4780);
nor U5991 (N_5991,N_4834,N_4536);
nand U5992 (N_5992,N_4273,N_4351);
nor U5993 (N_5993,N_4183,N_4274);
and U5994 (N_5994,N_4509,N_4413);
nor U5995 (N_5995,N_4291,N_4227);
or U5996 (N_5996,N_4399,N_4809);
nand U5997 (N_5997,N_4062,N_4924);
or U5998 (N_5998,N_4523,N_4966);
nor U5999 (N_5999,N_4713,N_4866);
or U6000 (N_6000,N_5084,N_5099);
and U6001 (N_6001,N_5219,N_5089);
nor U6002 (N_6002,N_5845,N_5326);
nand U6003 (N_6003,N_5036,N_5346);
and U6004 (N_6004,N_5037,N_5543);
and U6005 (N_6005,N_5976,N_5888);
nor U6006 (N_6006,N_5924,N_5134);
nand U6007 (N_6007,N_5832,N_5760);
or U6008 (N_6008,N_5006,N_5053);
and U6009 (N_6009,N_5223,N_5176);
or U6010 (N_6010,N_5467,N_5491);
nor U6011 (N_6011,N_5727,N_5653);
or U6012 (N_6012,N_5501,N_5698);
and U6013 (N_6013,N_5095,N_5007);
nand U6014 (N_6014,N_5933,N_5798);
nand U6015 (N_6015,N_5387,N_5474);
nand U6016 (N_6016,N_5351,N_5286);
nor U6017 (N_6017,N_5447,N_5364);
nor U6018 (N_6018,N_5334,N_5399);
and U6019 (N_6019,N_5138,N_5785);
nor U6020 (N_6020,N_5621,N_5405);
or U6021 (N_6021,N_5449,N_5208);
or U6022 (N_6022,N_5726,N_5265);
nor U6023 (N_6023,N_5600,N_5633);
or U6024 (N_6024,N_5397,N_5817);
nor U6025 (N_6025,N_5964,N_5586);
and U6026 (N_6026,N_5630,N_5946);
nand U6027 (N_6027,N_5807,N_5808);
and U6028 (N_6028,N_5854,N_5603);
nand U6029 (N_6029,N_5379,N_5041);
nand U6030 (N_6030,N_5672,N_5228);
or U6031 (N_6031,N_5169,N_5662);
nand U6032 (N_6032,N_5076,N_5980);
or U6033 (N_6033,N_5168,N_5377);
and U6034 (N_6034,N_5165,N_5713);
nand U6035 (N_6035,N_5678,N_5688);
xor U6036 (N_6036,N_5156,N_5434);
nor U6037 (N_6037,N_5482,N_5602);
or U6038 (N_6038,N_5802,N_5240);
nand U6039 (N_6039,N_5712,N_5120);
nand U6040 (N_6040,N_5526,N_5161);
nor U6041 (N_6041,N_5073,N_5948);
nand U6042 (N_6042,N_5883,N_5093);
or U6043 (N_6043,N_5551,N_5699);
nand U6044 (N_6044,N_5097,N_5042);
or U6045 (N_6045,N_5711,N_5507);
and U6046 (N_6046,N_5730,N_5233);
nand U6047 (N_6047,N_5339,N_5429);
and U6048 (N_6048,N_5287,N_5347);
or U6049 (N_6049,N_5128,N_5503);
and U6050 (N_6050,N_5506,N_5859);
nand U6051 (N_6051,N_5516,N_5654);
and U6052 (N_6052,N_5135,N_5673);
or U6053 (N_6053,N_5126,N_5444);
nor U6054 (N_6054,N_5562,N_5674);
nand U6055 (N_6055,N_5754,N_5663);
or U6056 (N_6056,N_5133,N_5763);
and U6057 (N_6057,N_5220,N_5009);
nor U6058 (N_6058,N_5060,N_5306);
nand U6059 (N_6059,N_5361,N_5159);
nor U6060 (N_6060,N_5715,N_5432);
or U6061 (N_6061,N_5427,N_5408);
nor U6062 (N_6062,N_5105,N_5871);
nand U6063 (N_6063,N_5034,N_5840);
and U6064 (N_6064,N_5420,N_5823);
nand U6065 (N_6065,N_5256,N_5075);
or U6066 (N_6066,N_5174,N_5568);
xor U6067 (N_6067,N_5343,N_5544);
xor U6068 (N_6068,N_5033,N_5731);
nor U6069 (N_6069,N_5224,N_5625);
or U6070 (N_6070,N_5511,N_5775);
nand U6071 (N_6071,N_5709,N_5786);
nand U6072 (N_6072,N_5862,N_5787);
and U6073 (N_6073,N_5446,N_5490);
or U6074 (N_6074,N_5864,N_5940);
xnor U6075 (N_6075,N_5484,N_5649);
and U6076 (N_6076,N_5899,N_5701);
nor U6077 (N_6077,N_5062,N_5358);
nand U6078 (N_6078,N_5183,N_5173);
and U6079 (N_6079,N_5067,N_5355);
nor U6080 (N_6080,N_5282,N_5904);
nor U6081 (N_6081,N_5370,N_5676);
nand U6082 (N_6082,N_5349,N_5741);
nand U6083 (N_6083,N_5695,N_5929);
or U6084 (N_6084,N_5026,N_5172);
nand U6085 (N_6085,N_5154,N_5396);
nand U6086 (N_6086,N_5632,N_5315);
nand U6087 (N_6087,N_5108,N_5212);
nor U6088 (N_6088,N_5542,N_5270);
and U6089 (N_6089,N_5866,N_5372);
or U6090 (N_6090,N_5495,N_5189);
nor U6091 (N_6091,N_5556,N_5739);
and U6092 (N_6092,N_5456,N_5327);
and U6093 (N_6093,N_5644,N_5365);
and U6094 (N_6094,N_5818,N_5710);
and U6095 (N_6095,N_5241,N_5734);
nand U6096 (N_6096,N_5191,N_5525);
nor U6097 (N_6097,N_5504,N_5769);
or U6098 (N_6098,N_5912,N_5117);
and U6099 (N_6099,N_5069,N_5416);
and U6100 (N_6100,N_5837,N_5519);
nor U6101 (N_6101,N_5198,N_5719);
and U6102 (N_6102,N_5475,N_5557);
nor U6103 (N_6103,N_5524,N_5570);
nand U6104 (N_6104,N_5949,N_5577);
nor U6105 (N_6105,N_5629,N_5951);
nor U6106 (N_6106,N_5990,N_5881);
nor U6107 (N_6107,N_5812,N_5402);
nor U6108 (N_6108,N_5266,N_5297);
nand U6109 (N_6109,N_5004,N_5911);
and U6110 (N_6110,N_5445,N_5826);
nor U6111 (N_6111,N_5532,N_5038);
nor U6112 (N_6112,N_5943,N_5560);
nor U6113 (N_6113,N_5927,N_5129);
or U6114 (N_6114,N_5919,N_5874);
or U6115 (N_6115,N_5764,N_5584);
nor U6116 (N_6116,N_5002,N_5112);
and U6117 (N_6117,N_5045,N_5522);
nor U6118 (N_6118,N_5248,N_5805);
xor U6119 (N_6119,N_5103,N_5916);
and U6120 (N_6120,N_5635,N_5657);
or U6121 (N_6121,N_5955,N_5063);
nor U6122 (N_6122,N_5953,N_5576);
nand U6123 (N_6123,N_5246,N_5459);
or U6124 (N_6124,N_5891,N_5815);
nor U6125 (N_6125,N_5656,N_5296);
and U6126 (N_6126,N_5765,N_5043);
or U6127 (N_6127,N_5025,N_5055);
and U6128 (N_6128,N_5332,N_5243);
nand U6129 (N_6129,N_5460,N_5974);
or U6130 (N_6130,N_5483,N_5792);
xor U6131 (N_6131,N_5380,N_5061);
nor U6132 (N_6132,N_5131,N_5909);
or U6133 (N_6133,N_5594,N_5969);
nor U6134 (N_6134,N_5356,N_5797);
nand U6135 (N_6135,N_5274,N_5162);
or U6136 (N_6136,N_5618,N_5637);
or U6137 (N_6137,N_5563,N_5439);
nand U6138 (N_6138,N_5641,N_5958);
nand U6139 (N_6139,N_5796,N_5921);
xnor U6140 (N_6140,N_5886,N_5622);
nor U6141 (N_6141,N_5294,N_5206);
or U6142 (N_6142,N_5923,N_5342);
or U6143 (N_6143,N_5552,N_5694);
nand U6144 (N_6144,N_5421,N_5195);
xor U6145 (N_6145,N_5825,N_5122);
nand U6146 (N_6146,N_5669,N_5596);
or U6147 (N_6147,N_5777,N_5824);
nand U6148 (N_6148,N_5424,N_5636);
or U6149 (N_6149,N_5702,N_5993);
nor U6150 (N_6150,N_5264,N_5865);
and U6151 (N_6151,N_5070,N_5468);
nand U6152 (N_6152,N_5589,N_5583);
nor U6153 (N_6153,N_5896,N_5058);
xnor U6154 (N_6154,N_5203,N_5956);
and U6155 (N_6155,N_5268,N_5123);
or U6156 (N_6156,N_5647,N_5113);
nor U6157 (N_6157,N_5328,N_5231);
and U6158 (N_6158,N_5217,N_5163);
and U6159 (N_6159,N_5436,N_5150);
or U6160 (N_6160,N_5360,N_5366);
and U6161 (N_6161,N_5788,N_5455);
and U6162 (N_6162,N_5018,N_5121);
nand U6163 (N_6163,N_5151,N_5391);
and U6164 (N_6164,N_5350,N_5857);
or U6165 (N_6165,N_5975,N_5487);
or U6166 (N_6166,N_5118,N_5218);
and U6167 (N_6167,N_5932,N_5747);
xnor U6168 (N_6168,N_5376,N_5239);
and U6169 (N_6169,N_5806,N_5317);
xor U6170 (N_6170,N_5308,N_5035);
or U6171 (N_6171,N_5677,N_5898);
nor U6172 (N_6172,N_5180,N_5795);
or U6173 (N_6173,N_5092,N_5530);
nor U6174 (N_6174,N_5601,N_5738);
nor U6175 (N_6175,N_5406,N_5938);
nand U6176 (N_6176,N_5152,N_5725);
or U6177 (N_6177,N_5723,N_5690);
nand U6178 (N_6178,N_5083,N_5140);
nand U6179 (N_6179,N_5804,N_5272);
or U6180 (N_6180,N_5080,N_5861);
or U6181 (N_6181,N_5531,N_5598);
nand U6182 (N_6182,N_5894,N_5100);
nand U6183 (N_6183,N_5448,N_5793);
nor U6184 (N_6184,N_5454,N_5931);
and U6185 (N_6185,N_5970,N_5384);
or U6186 (N_6186,N_5010,N_5978);
nand U6187 (N_6187,N_5079,N_5915);
nand U6188 (N_6188,N_5196,N_5890);
and U6189 (N_6189,N_5028,N_5984);
and U6190 (N_6190,N_5450,N_5994);
nor U6191 (N_6191,N_5561,N_5031);
xor U6192 (N_6192,N_5481,N_5211);
nor U6193 (N_6193,N_5573,N_5882);
and U6194 (N_6194,N_5820,N_5245);
or U6195 (N_6195,N_5517,N_5145);
nand U6196 (N_6196,N_5816,N_5950);
or U6197 (N_6197,N_5609,N_5383);
nand U6198 (N_6198,N_5341,N_5452);
nor U6199 (N_6199,N_5616,N_5494);
nor U6200 (N_6200,N_5528,N_5071);
nor U6201 (N_6201,N_5143,N_5740);
nand U6202 (N_6202,N_5569,N_5205);
nand U6203 (N_6203,N_5628,N_5375);
nor U6204 (N_6204,N_5799,N_5720);
or U6205 (N_6205,N_5177,N_5939);
and U6206 (N_6206,N_5226,N_5510);
xnor U6207 (N_6207,N_5546,N_5645);
nor U6208 (N_6208,N_5558,N_5348);
nand U6209 (N_6209,N_5304,N_5473);
nor U6210 (N_6210,N_5064,N_5838);
and U6211 (N_6211,N_5367,N_5767);
nor U6212 (N_6212,N_5389,N_5110);
and U6213 (N_6213,N_5513,N_5409);
nor U6214 (N_6214,N_5724,N_5257);
nand U6215 (N_6215,N_5395,N_5300);
and U6216 (N_6216,N_5703,N_5972);
nor U6217 (N_6217,N_5537,N_5914);
nand U6218 (N_6218,N_5534,N_5860);
nand U6219 (N_6219,N_5499,N_5566);
nand U6220 (N_6220,N_5784,N_5571);
or U6221 (N_6221,N_5288,N_5608);
nor U6222 (N_6222,N_5142,N_5518);
and U6223 (N_6223,N_5498,N_5390);
nor U6224 (N_6224,N_5147,N_5856);
or U6225 (N_6225,N_5853,N_5340);
and U6226 (N_6226,N_5433,N_5858);
or U6227 (N_6227,N_5954,N_5839);
nor U6228 (N_6228,N_5170,N_5307);
nor U6229 (N_6229,N_5612,N_5054);
or U6230 (N_6230,N_5471,N_5193);
nor U6231 (N_6231,N_5761,N_5316);
nand U6232 (N_6232,N_5947,N_5381);
and U6233 (N_6233,N_5352,N_5019);
or U6234 (N_6234,N_5579,N_5422);
nor U6235 (N_6235,N_5250,N_5281);
nand U6236 (N_6236,N_5235,N_5329);
or U6237 (N_6237,N_5512,N_5209);
nand U6238 (N_6238,N_5850,N_5291);
or U6239 (N_6239,N_5213,N_5425);
xor U6240 (N_6240,N_5884,N_5305);
or U6241 (N_6241,N_5144,N_5486);
nand U6242 (N_6242,N_5800,N_5574);
nand U6243 (N_6243,N_5782,N_5988);
nand U6244 (N_6244,N_5908,N_5944);
and U6245 (N_6245,N_5697,N_5252);
or U6246 (N_6246,N_5283,N_5021);
nand U6247 (N_6247,N_5175,N_5101);
nor U6248 (N_6248,N_5776,N_5892);
nand U6249 (N_6249,N_5930,N_5968);
nor U6250 (N_6250,N_5215,N_5046);
or U6251 (N_6251,N_5199,N_5385);
nand U6252 (N_6252,N_5648,N_5852);
and U6253 (N_6253,N_5290,N_5922);
xnor U6254 (N_6254,N_5736,N_5158);
nand U6255 (N_6255,N_5016,N_5462);
and U6256 (N_6256,N_5696,N_5412);
or U6257 (N_6257,N_5849,N_5995);
and U6258 (N_6258,N_5124,N_5827);
and U6259 (N_6259,N_5575,N_5335);
nor U6260 (N_6260,N_5255,N_5115);
nand U6261 (N_6261,N_5497,N_5684);
and U6262 (N_6262,N_5072,N_5087);
and U6263 (N_6263,N_5074,N_5756);
or U6264 (N_6264,N_5878,N_5961);
nand U6265 (N_6265,N_5781,N_5936);
xor U6266 (N_6266,N_5435,N_5547);
xnor U6267 (N_6267,N_5626,N_5210);
nor U6268 (N_6268,N_5311,N_5664);
nand U6269 (N_6269,N_5357,N_5130);
xor U6270 (N_6270,N_5572,N_5545);
or U6271 (N_6271,N_5178,N_5284);
nand U6272 (N_6272,N_5721,N_5689);
or U6273 (N_6273,N_5363,N_5027);
xnor U6274 (N_6274,N_5771,N_5125);
and U6275 (N_6275,N_5989,N_5431);
or U6276 (N_6276,N_5834,N_5309);
nand U6277 (N_6277,N_5591,N_5935);
nor U6278 (N_6278,N_5164,N_5607);
nand U6279 (N_6279,N_5515,N_5292);
nor U6280 (N_6280,N_5666,N_5998);
nor U6281 (N_6281,N_5863,N_5821);
nand U6282 (N_6282,N_5533,N_5017);
and U6283 (N_6283,N_5643,N_5407);
or U6284 (N_6284,N_5870,N_5267);
nand U6285 (N_6285,N_5285,N_5289);
nand U6286 (N_6286,N_5751,N_5373);
xnor U6287 (N_6287,N_5873,N_5453);
and U6288 (N_6288,N_5634,N_5214);
or U6289 (N_6289,N_5905,N_5780);
nand U6290 (N_6290,N_5082,N_5279);
and U6291 (N_6291,N_5691,N_5755);
and U6292 (N_6292,N_5249,N_5437);
or U6293 (N_6293,N_5928,N_5655);
xnor U6294 (N_6294,N_5386,N_5813);
nor U6295 (N_6295,N_5417,N_5809);
and U6296 (N_6296,N_5614,N_5020);
nand U6297 (N_6297,N_5259,N_5867);
nand U6298 (N_6298,N_5015,N_5477);
nor U6299 (N_6299,N_5090,N_5234);
nand U6300 (N_6300,N_5750,N_5597);
nor U6301 (N_6301,N_5963,N_5104);
or U6302 (N_6302,N_5423,N_5508);
nand U6303 (N_6303,N_5605,N_5997);
nor U6304 (N_6304,N_5393,N_5564);
xnor U6305 (N_6305,N_5842,N_5746);
and U6306 (N_6306,N_5299,N_5548);
nor U6307 (N_6307,N_5369,N_5094);
and U6308 (N_6308,N_5620,N_5277);
nand U6309 (N_6309,N_5496,N_5464);
or U6310 (N_6310,N_5085,N_5611);
nand U6311 (N_6311,N_5059,N_5962);
nand U6312 (N_6312,N_5977,N_5116);
nor U6313 (N_6313,N_5012,N_5879);
nand U6314 (N_6314,N_5841,N_5242);
xnor U6315 (N_6315,N_5378,N_5952);
nand U6316 (N_6316,N_5253,N_5661);
nand U6317 (N_6317,N_5639,N_5368);
or U6318 (N_6318,N_5302,N_5470);
nor U6319 (N_6319,N_5638,N_5658);
nor U6320 (N_6320,N_5077,N_5830);
nand U6321 (N_6321,N_5735,N_5003);
nor U6322 (N_6322,N_5204,N_5237);
xnor U6323 (N_6323,N_5032,N_5748);
xor U6324 (N_6324,N_5013,N_5523);
or U6325 (N_6325,N_5303,N_5500);
xnor U6326 (N_6326,N_5157,N_5682);
and U6327 (N_6327,N_5791,N_5251);
nor U6328 (N_6328,N_5008,N_5565);
or U6329 (N_6329,N_5106,N_5766);
nand U6330 (N_6330,N_5489,N_5918);
or U6331 (N_6331,N_5029,N_5700);
or U6332 (N_6332,N_5388,N_5414);
or U6333 (N_6333,N_5039,N_5986);
and U6334 (N_6334,N_5665,N_5221);
and U6335 (N_6335,N_5187,N_5065);
nor U6336 (N_6336,N_5410,N_5493);
nand U6337 (N_6337,N_5107,N_5167);
and U6338 (N_6338,N_5318,N_5650);
nand U6339 (N_6339,N_5707,N_5778);
nor U6340 (N_6340,N_5109,N_5717);
or U6341 (N_6341,N_5520,N_5394);
or U6342 (N_6342,N_5835,N_5617);
nand U6343 (N_6343,N_5441,N_5418);
xnor U6344 (N_6344,N_5298,N_5553);
nand U6345 (N_6345,N_5040,N_5836);
and U6346 (N_6346,N_5202,N_5322);
nor U6347 (N_6347,N_5023,N_5773);
and U6348 (N_6348,N_5230,N_5426);
or U6349 (N_6349,N_5153,N_5048);
nand U6350 (N_6350,N_5232,N_5774);
and U6351 (N_6351,N_5743,N_5509);
xnor U6352 (N_6352,N_5991,N_5957);
and U6353 (N_6353,N_5768,N_5492);
or U6354 (N_6354,N_5996,N_5679);
nand U6355 (N_6355,N_5275,N_5675);
nand U6356 (N_6356,N_5758,N_5502);
nand U6357 (N_6357,N_5238,N_5555);
or U6358 (N_6358,N_5960,N_5190);
nor U6359 (N_6359,N_5262,N_5068);
nand U6360 (N_6360,N_5590,N_5102);
xor U6361 (N_6361,N_5000,N_5344);
nor U6362 (N_6362,N_5521,N_5320);
nor U6363 (N_6363,N_5578,N_5877);
nand U6364 (N_6364,N_5732,N_5581);
nand U6365 (N_6365,N_5716,N_5801);
nor U6366 (N_6366,N_5201,N_5185);
nand U6367 (N_6367,N_5457,N_5024);
or U6368 (N_6368,N_5312,N_5917);
nor U6369 (N_6369,N_5959,N_5889);
nor U6370 (N_6370,N_5744,N_5683);
and U6371 (N_6371,N_5066,N_5982);
xor U6372 (N_6372,N_5926,N_5398);
nand U6373 (N_6373,N_5868,N_5321);
nor U6374 (N_6374,N_5985,N_5681);
nor U6375 (N_6375,N_5472,N_5651);
nor U6376 (N_6376,N_5295,N_5538);
nand U6377 (N_6377,N_5148,N_5992);
nand U6378 (N_6378,N_5880,N_5869);
xnor U6379 (N_6379,N_5280,N_5722);
nor U6380 (N_6380,N_5708,N_5411);
nor U6381 (N_6381,N_5667,N_5906);
and U6382 (N_6382,N_5687,N_5599);
or U6383 (N_6383,N_5078,N_5330);
or U6384 (N_6384,N_5942,N_5907);
or U6385 (N_6385,N_5338,N_5983);
or U6386 (N_6386,N_5987,N_5671);
nor U6387 (N_6387,N_5336,N_5966);
and U6388 (N_6388,N_5188,N_5604);
or U6389 (N_6389,N_5981,N_5704);
and U6390 (N_6390,N_5415,N_5670);
nand U6391 (N_6391,N_5624,N_5762);
nand U6392 (N_6392,N_5337,N_5937);
or U6393 (N_6393,N_5718,N_5011);
and U6394 (N_6394,N_5155,N_5705);
nor U6395 (N_6395,N_5759,N_5465);
and U6396 (N_6396,N_5149,N_5001);
or U6397 (N_6397,N_5132,N_5770);
and U6398 (N_6398,N_5831,N_5114);
xor U6399 (N_6399,N_5680,N_5476);
nor U6400 (N_6400,N_5333,N_5222);
xor U6401 (N_6401,N_5052,N_5595);
or U6402 (N_6402,N_5463,N_5371);
nor U6403 (N_6403,N_5772,N_5325);
nand U6404 (N_6404,N_5419,N_5278);
and U6405 (N_6405,N_5592,N_5005);
nand U6406 (N_6406,N_5692,N_5354);
nand U6407 (N_6407,N_5737,N_5428);
nor U6408 (N_6408,N_5529,N_5194);
nor U6409 (N_6409,N_5324,N_5086);
nor U6410 (N_6410,N_5401,N_5686);
or U6411 (N_6411,N_5783,N_5876);
and U6412 (N_6412,N_5779,N_5096);
and U6413 (N_6413,N_5269,N_5119);
nand U6414 (N_6414,N_5659,N_5631);
and U6415 (N_6415,N_5895,N_5875);
and U6416 (N_6416,N_5200,N_5893);
nor U6417 (N_6417,N_5945,N_5789);
nand U6418 (N_6418,N_5244,N_5541);
nor U6419 (N_6419,N_5646,N_5192);
or U6420 (N_6420,N_5685,N_5313);
or U6421 (N_6421,N_5851,N_5137);
or U6422 (N_6422,N_5623,N_5403);
nor U6423 (N_6423,N_5822,N_5934);
nor U6424 (N_6424,N_5182,N_5803);
and U6425 (N_6425,N_5833,N_5706);
nand U6426 (N_6426,N_5088,N_5745);
and U6427 (N_6427,N_5098,N_5536);
and U6428 (N_6428,N_5941,N_5461);
nor U6429 (N_6429,N_5897,N_5642);
or U6430 (N_6430,N_5810,N_5728);
nand U6431 (N_6431,N_5829,N_5901);
and U6432 (N_6432,N_5846,N_5127);
and U6433 (N_6433,N_5451,N_5790);
nand U6434 (N_6434,N_5049,N_5549);
or U6435 (N_6435,N_5606,N_5965);
or U6436 (N_6436,N_5971,N_5587);
nand U6437 (N_6437,N_5458,N_5184);
nand U6438 (N_6438,N_5273,N_5828);
xor U6439 (N_6439,N_5111,N_5050);
nor U6440 (N_6440,N_5580,N_5353);
and U6441 (N_6441,N_5627,N_5051);
nor U6442 (N_6442,N_5443,N_5258);
nand U6443 (N_6443,N_5582,N_5903);
nand U6444 (N_6444,N_5550,N_5216);
nand U6445 (N_6445,N_5967,N_5181);
or U6446 (N_6446,N_5749,N_5478);
or U6447 (N_6447,N_5593,N_5814);
nor U6448 (N_6448,N_5392,N_5413);
xor U6449 (N_6449,N_5247,N_5872);
or U6450 (N_6450,N_5136,N_5640);
or U6451 (N_6451,N_5714,N_5166);
and U6452 (N_6452,N_5374,N_5973);
or U6453 (N_6453,N_5811,N_5081);
or U6454 (N_6454,N_5588,N_5619);
or U6455 (N_6455,N_5479,N_5847);
nor U6456 (N_6456,N_5261,N_5197);
nor U6457 (N_6457,N_5310,N_5920);
or U6458 (N_6458,N_5615,N_5733);
or U6459 (N_6459,N_5260,N_5382);
xor U6460 (N_6460,N_5505,N_5056);
and U6461 (N_6461,N_5047,N_5276);
or U6462 (N_6462,N_5146,N_5913);
xor U6463 (N_6463,N_5225,N_5539);
nor U6464 (N_6464,N_5999,N_5668);
and U6465 (N_6465,N_5660,N_5902);
nand U6466 (N_6466,N_5844,N_5752);
or U6467 (N_6467,N_5900,N_5331);
nand U6468 (N_6468,N_5171,N_5613);
or U6469 (N_6469,N_5263,N_5585);
or U6470 (N_6470,N_5044,N_5757);
and U6471 (N_6471,N_5141,N_5438);
nor U6472 (N_6472,N_5554,N_5430);
nor U6473 (N_6473,N_5540,N_5139);
xor U6474 (N_6474,N_5314,N_5319);
and U6475 (N_6475,N_5179,N_5794);
and U6476 (N_6476,N_5819,N_5729);
nor U6477 (N_6477,N_5485,N_5271);
xor U6478 (N_6478,N_5488,N_5014);
nand U6479 (N_6479,N_5925,N_5843);
xor U6480 (N_6480,N_5610,N_5559);
or U6481 (N_6481,N_5753,N_5440);
nand U6482 (N_6482,N_5466,N_5855);
and U6483 (N_6483,N_5848,N_5091);
xor U6484 (N_6484,N_5567,N_5910);
and U6485 (N_6485,N_5293,N_5514);
nand U6486 (N_6486,N_5469,N_5979);
and U6487 (N_6487,N_5742,N_5400);
and U6488 (N_6488,N_5207,N_5885);
or U6489 (N_6489,N_5535,N_5345);
nand U6490 (N_6490,N_5323,N_5186);
and U6491 (N_6491,N_5359,N_5227);
nor U6492 (N_6492,N_5229,N_5254);
nand U6493 (N_6493,N_5057,N_5301);
nand U6494 (N_6494,N_5480,N_5404);
or U6495 (N_6495,N_5693,N_5652);
and U6496 (N_6496,N_5160,N_5442);
nor U6497 (N_6497,N_5236,N_5022);
nor U6498 (N_6498,N_5887,N_5362);
nand U6499 (N_6499,N_5527,N_5030);
nand U6500 (N_6500,N_5848,N_5853);
and U6501 (N_6501,N_5838,N_5421);
nand U6502 (N_6502,N_5304,N_5140);
and U6503 (N_6503,N_5426,N_5674);
nor U6504 (N_6504,N_5914,N_5974);
or U6505 (N_6505,N_5446,N_5616);
nor U6506 (N_6506,N_5774,N_5002);
and U6507 (N_6507,N_5295,N_5826);
and U6508 (N_6508,N_5271,N_5555);
or U6509 (N_6509,N_5323,N_5462);
nand U6510 (N_6510,N_5146,N_5227);
nand U6511 (N_6511,N_5861,N_5049);
and U6512 (N_6512,N_5323,N_5070);
nor U6513 (N_6513,N_5646,N_5082);
and U6514 (N_6514,N_5988,N_5462);
and U6515 (N_6515,N_5104,N_5922);
nor U6516 (N_6516,N_5860,N_5300);
and U6517 (N_6517,N_5138,N_5239);
or U6518 (N_6518,N_5780,N_5653);
or U6519 (N_6519,N_5313,N_5225);
and U6520 (N_6520,N_5653,N_5604);
and U6521 (N_6521,N_5811,N_5388);
or U6522 (N_6522,N_5745,N_5441);
or U6523 (N_6523,N_5383,N_5919);
nand U6524 (N_6524,N_5718,N_5181);
xor U6525 (N_6525,N_5182,N_5711);
or U6526 (N_6526,N_5392,N_5276);
or U6527 (N_6527,N_5588,N_5130);
nand U6528 (N_6528,N_5586,N_5906);
nand U6529 (N_6529,N_5512,N_5742);
nor U6530 (N_6530,N_5426,N_5236);
nand U6531 (N_6531,N_5094,N_5701);
nor U6532 (N_6532,N_5532,N_5870);
and U6533 (N_6533,N_5165,N_5753);
or U6534 (N_6534,N_5798,N_5723);
nor U6535 (N_6535,N_5800,N_5710);
nand U6536 (N_6536,N_5944,N_5108);
and U6537 (N_6537,N_5249,N_5592);
nand U6538 (N_6538,N_5117,N_5814);
or U6539 (N_6539,N_5452,N_5391);
nand U6540 (N_6540,N_5546,N_5905);
and U6541 (N_6541,N_5764,N_5811);
or U6542 (N_6542,N_5131,N_5683);
nand U6543 (N_6543,N_5105,N_5712);
nor U6544 (N_6544,N_5870,N_5926);
or U6545 (N_6545,N_5674,N_5670);
nor U6546 (N_6546,N_5449,N_5356);
nand U6547 (N_6547,N_5168,N_5942);
or U6548 (N_6548,N_5000,N_5027);
and U6549 (N_6549,N_5693,N_5324);
and U6550 (N_6550,N_5008,N_5455);
nor U6551 (N_6551,N_5148,N_5683);
xor U6552 (N_6552,N_5873,N_5479);
nand U6553 (N_6553,N_5175,N_5657);
or U6554 (N_6554,N_5250,N_5082);
or U6555 (N_6555,N_5599,N_5506);
or U6556 (N_6556,N_5931,N_5647);
and U6557 (N_6557,N_5603,N_5330);
nor U6558 (N_6558,N_5277,N_5363);
and U6559 (N_6559,N_5765,N_5679);
and U6560 (N_6560,N_5322,N_5874);
and U6561 (N_6561,N_5586,N_5771);
or U6562 (N_6562,N_5429,N_5888);
nand U6563 (N_6563,N_5777,N_5119);
nand U6564 (N_6564,N_5002,N_5069);
nand U6565 (N_6565,N_5287,N_5001);
and U6566 (N_6566,N_5635,N_5866);
nor U6567 (N_6567,N_5894,N_5664);
nand U6568 (N_6568,N_5598,N_5237);
nand U6569 (N_6569,N_5441,N_5679);
nand U6570 (N_6570,N_5896,N_5455);
xor U6571 (N_6571,N_5924,N_5121);
or U6572 (N_6572,N_5764,N_5745);
nor U6573 (N_6573,N_5138,N_5475);
nand U6574 (N_6574,N_5814,N_5802);
nand U6575 (N_6575,N_5988,N_5990);
or U6576 (N_6576,N_5235,N_5232);
nor U6577 (N_6577,N_5601,N_5466);
nor U6578 (N_6578,N_5684,N_5287);
nor U6579 (N_6579,N_5666,N_5662);
nor U6580 (N_6580,N_5989,N_5826);
nand U6581 (N_6581,N_5677,N_5849);
or U6582 (N_6582,N_5257,N_5828);
and U6583 (N_6583,N_5546,N_5334);
nor U6584 (N_6584,N_5702,N_5469);
nand U6585 (N_6585,N_5611,N_5658);
or U6586 (N_6586,N_5793,N_5256);
and U6587 (N_6587,N_5392,N_5240);
or U6588 (N_6588,N_5571,N_5102);
nor U6589 (N_6589,N_5058,N_5118);
and U6590 (N_6590,N_5136,N_5765);
or U6591 (N_6591,N_5407,N_5673);
nor U6592 (N_6592,N_5812,N_5271);
nand U6593 (N_6593,N_5526,N_5372);
or U6594 (N_6594,N_5944,N_5075);
nand U6595 (N_6595,N_5165,N_5665);
nand U6596 (N_6596,N_5891,N_5896);
nor U6597 (N_6597,N_5853,N_5771);
nor U6598 (N_6598,N_5178,N_5048);
nand U6599 (N_6599,N_5928,N_5277);
nand U6600 (N_6600,N_5308,N_5380);
nand U6601 (N_6601,N_5978,N_5993);
xor U6602 (N_6602,N_5707,N_5772);
nor U6603 (N_6603,N_5574,N_5545);
and U6604 (N_6604,N_5147,N_5815);
nor U6605 (N_6605,N_5716,N_5151);
nand U6606 (N_6606,N_5200,N_5393);
and U6607 (N_6607,N_5385,N_5667);
nand U6608 (N_6608,N_5034,N_5699);
or U6609 (N_6609,N_5471,N_5961);
nor U6610 (N_6610,N_5120,N_5001);
nand U6611 (N_6611,N_5133,N_5639);
and U6612 (N_6612,N_5477,N_5330);
and U6613 (N_6613,N_5949,N_5625);
or U6614 (N_6614,N_5550,N_5955);
and U6615 (N_6615,N_5118,N_5878);
nor U6616 (N_6616,N_5924,N_5428);
nand U6617 (N_6617,N_5148,N_5864);
or U6618 (N_6618,N_5558,N_5777);
xnor U6619 (N_6619,N_5678,N_5590);
or U6620 (N_6620,N_5691,N_5758);
nor U6621 (N_6621,N_5189,N_5284);
xor U6622 (N_6622,N_5857,N_5114);
nand U6623 (N_6623,N_5299,N_5979);
and U6624 (N_6624,N_5141,N_5677);
nor U6625 (N_6625,N_5116,N_5017);
nor U6626 (N_6626,N_5687,N_5596);
nand U6627 (N_6627,N_5209,N_5999);
or U6628 (N_6628,N_5527,N_5308);
nand U6629 (N_6629,N_5533,N_5950);
or U6630 (N_6630,N_5900,N_5188);
or U6631 (N_6631,N_5877,N_5067);
nand U6632 (N_6632,N_5598,N_5524);
nor U6633 (N_6633,N_5705,N_5273);
nor U6634 (N_6634,N_5303,N_5746);
and U6635 (N_6635,N_5296,N_5741);
and U6636 (N_6636,N_5494,N_5568);
and U6637 (N_6637,N_5168,N_5789);
nand U6638 (N_6638,N_5001,N_5903);
or U6639 (N_6639,N_5959,N_5775);
nand U6640 (N_6640,N_5110,N_5753);
nand U6641 (N_6641,N_5742,N_5579);
nand U6642 (N_6642,N_5971,N_5647);
nand U6643 (N_6643,N_5795,N_5744);
nand U6644 (N_6644,N_5214,N_5748);
and U6645 (N_6645,N_5881,N_5236);
or U6646 (N_6646,N_5894,N_5113);
or U6647 (N_6647,N_5783,N_5551);
or U6648 (N_6648,N_5633,N_5563);
and U6649 (N_6649,N_5434,N_5734);
nor U6650 (N_6650,N_5994,N_5011);
and U6651 (N_6651,N_5075,N_5063);
or U6652 (N_6652,N_5859,N_5997);
or U6653 (N_6653,N_5377,N_5388);
nor U6654 (N_6654,N_5296,N_5375);
nor U6655 (N_6655,N_5343,N_5192);
nor U6656 (N_6656,N_5477,N_5279);
and U6657 (N_6657,N_5200,N_5696);
and U6658 (N_6658,N_5073,N_5599);
or U6659 (N_6659,N_5410,N_5136);
nor U6660 (N_6660,N_5386,N_5455);
xor U6661 (N_6661,N_5977,N_5956);
and U6662 (N_6662,N_5769,N_5398);
or U6663 (N_6663,N_5134,N_5047);
and U6664 (N_6664,N_5406,N_5059);
xor U6665 (N_6665,N_5146,N_5448);
nand U6666 (N_6666,N_5919,N_5373);
nand U6667 (N_6667,N_5548,N_5838);
nor U6668 (N_6668,N_5038,N_5491);
nand U6669 (N_6669,N_5192,N_5812);
nor U6670 (N_6670,N_5299,N_5025);
xor U6671 (N_6671,N_5350,N_5472);
xor U6672 (N_6672,N_5033,N_5001);
nor U6673 (N_6673,N_5498,N_5546);
xnor U6674 (N_6674,N_5371,N_5752);
nor U6675 (N_6675,N_5560,N_5500);
nor U6676 (N_6676,N_5025,N_5494);
or U6677 (N_6677,N_5244,N_5578);
nand U6678 (N_6678,N_5954,N_5706);
nand U6679 (N_6679,N_5976,N_5754);
or U6680 (N_6680,N_5612,N_5392);
nand U6681 (N_6681,N_5857,N_5356);
nand U6682 (N_6682,N_5376,N_5430);
and U6683 (N_6683,N_5013,N_5041);
xnor U6684 (N_6684,N_5264,N_5610);
and U6685 (N_6685,N_5724,N_5552);
nand U6686 (N_6686,N_5891,N_5778);
nor U6687 (N_6687,N_5079,N_5616);
nor U6688 (N_6688,N_5219,N_5589);
xnor U6689 (N_6689,N_5858,N_5265);
nand U6690 (N_6690,N_5090,N_5650);
or U6691 (N_6691,N_5614,N_5737);
nand U6692 (N_6692,N_5758,N_5481);
nor U6693 (N_6693,N_5875,N_5563);
or U6694 (N_6694,N_5294,N_5843);
or U6695 (N_6695,N_5638,N_5275);
and U6696 (N_6696,N_5950,N_5467);
or U6697 (N_6697,N_5972,N_5818);
nor U6698 (N_6698,N_5438,N_5814);
nand U6699 (N_6699,N_5930,N_5599);
and U6700 (N_6700,N_5273,N_5908);
or U6701 (N_6701,N_5855,N_5351);
nor U6702 (N_6702,N_5581,N_5201);
nand U6703 (N_6703,N_5840,N_5223);
nand U6704 (N_6704,N_5933,N_5499);
or U6705 (N_6705,N_5896,N_5756);
nand U6706 (N_6706,N_5389,N_5695);
or U6707 (N_6707,N_5900,N_5742);
and U6708 (N_6708,N_5348,N_5718);
and U6709 (N_6709,N_5884,N_5148);
nand U6710 (N_6710,N_5492,N_5629);
or U6711 (N_6711,N_5055,N_5306);
nand U6712 (N_6712,N_5472,N_5875);
nor U6713 (N_6713,N_5300,N_5038);
nor U6714 (N_6714,N_5748,N_5775);
xor U6715 (N_6715,N_5621,N_5826);
and U6716 (N_6716,N_5982,N_5235);
and U6717 (N_6717,N_5796,N_5186);
xor U6718 (N_6718,N_5993,N_5920);
nand U6719 (N_6719,N_5240,N_5403);
and U6720 (N_6720,N_5331,N_5270);
and U6721 (N_6721,N_5733,N_5357);
and U6722 (N_6722,N_5793,N_5501);
nor U6723 (N_6723,N_5884,N_5302);
nor U6724 (N_6724,N_5985,N_5653);
or U6725 (N_6725,N_5605,N_5949);
or U6726 (N_6726,N_5808,N_5149);
nand U6727 (N_6727,N_5479,N_5795);
nand U6728 (N_6728,N_5553,N_5489);
or U6729 (N_6729,N_5848,N_5976);
or U6730 (N_6730,N_5557,N_5547);
and U6731 (N_6731,N_5595,N_5951);
nor U6732 (N_6732,N_5851,N_5067);
nand U6733 (N_6733,N_5452,N_5189);
or U6734 (N_6734,N_5931,N_5477);
nand U6735 (N_6735,N_5292,N_5147);
or U6736 (N_6736,N_5871,N_5817);
nor U6737 (N_6737,N_5016,N_5625);
nor U6738 (N_6738,N_5634,N_5500);
nor U6739 (N_6739,N_5643,N_5186);
nor U6740 (N_6740,N_5146,N_5346);
or U6741 (N_6741,N_5603,N_5702);
nor U6742 (N_6742,N_5720,N_5728);
nand U6743 (N_6743,N_5691,N_5095);
or U6744 (N_6744,N_5671,N_5829);
and U6745 (N_6745,N_5952,N_5905);
and U6746 (N_6746,N_5177,N_5620);
nand U6747 (N_6747,N_5022,N_5007);
nor U6748 (N_6748,N_5460,N_5286);
or U6749 (N_6749,N_5783,N_5044);
nor U6750 (N_6750,N_5373,N_5356);
and U6751 (N_6751,N_5078,N_5250);
xnor U6752 (N_6752,N_5561,N_5725);
xnor U6753 (N_6753,N_5776,N_5538);
nand U6754 (N_6754,N_5156,N_5932);
nand U6755 (N_6755,N_5411,N_5787);
or U6756 (N_6756,N_5710,N_5359);
nor U6757 (N_6757,N_5231,N_5281);
nand U6758 (N_6758,N_5002,N_5031);
or U6759 (N_6759,N_5118,N_5665);
and U6760 (N_6760,N_5382,N_5017);
nand U6761 (N_6761,N_5493,N_5069);
xor U6762 (N_6762,N_5549,N_5373);
and U6763 (N_6763,N_5293,N_5446);
nor U6764 (N_6764,N_5001,N_5463);
nor U6765 (N_6765,N_5925,N_5884);
nor U6766 (N_6766,N_5132,N_5520);
nor U6767 (N_6767,N_5615,N_5796);
and U6768 (N_6768,N_5955,N_5091);
nand U6769 (N_6769,N_5124,N_5040);
or U6770 (N_6770,N_5485,N_5344);
xnor U6771 (N_6771,N_5386,N_5835);
or U6772 (N_6772,N_5113,N_5171);
and U6773 (N_6773,N_5314,N_5461);
or U6774 (N_6774,N_5321,N_5201);
nor U6775 (N_6775,N_5606,N_5603);
and U6776 (N_6776,N_5254,N_5217);
and U6777 (N_6777,N_5381,N_5542);
and U6778 (N_6778,N_5574,N_5260);
xnor U6779 (N_6779,N_5195,N_5317);
and U6780 (N_6780,N_5940,N_5472);
nor U6781 (N_6781,N_5843,N_5345);
and U6782 (N_6782,N_5569,N_5773);
and U6783 (N_6783,N_5673,N_5740);
nand U6784 (N_6784,N_5821,N_5128);
nor U6785 (N_6785,N_5509,N_5694);
and U6786 (N_6786,N_5646,N_5808);
nor U6787 (N_6787,N_5628,N_5976);
or U6788 (N_6788,N_5352,N_5573);
nand U6789 (N_6789,N_5955,N_5162);
nor U6790 (N_6790,N_5456,N_5094);
or U6791 (N_6791,N_5825,N_5326);
nand U6792 (N_6792,N_5089,N_5863);
and U6793 (N_6793,N_5137,N_5669);
and U6794 (N_6794,N_5258,N_5322);
or U6795 (N_6795,N_5114,N_5615);
or U6796 (N_6796,N_5917,N_5459);
and U6797 (N_6797,N_5844,N_5021);
and U6798 (N_6798,N_5920,N_5566);
or U6799 (N_6799,N_5140,N_5822);
or U6800 (N_6800,N_5010,N_5993);
xnor U6801 (N_6801,N_5732,N_5402);
or U6802 (N_6802,N_5164,N_5436);
nand U6803 (N_6803,N_5830,N_5941);
or U6804 (N_6804,N_5923,N_5858);
nor U6805 (N_6805,N_5687,N_5767);
nand U6806 (N_6806,N_5290,N_5720);
nand U6807 (N_6807,N_5207,N_5893);
and U6808 (N_6808,N_5112,N_5510);
nor U6809 (N_6809,N_5804,N_5113);
and U6810 (N_6810,N_5439,N_5696);
and U6811 (N_6811,N_5749,N_5499);
or U6812 (N_6812,N_5218,N_5913);
xor U6813 (N_6813,N_5314,N_5205);
nand U6814 (N_6814,N_5688,N_5137);
and U6815 (N_6815,N_5700,N_5414);
and U6816 (N_6816,N_5458,N_5078);
or U6817 (N_6817,N_5711,N_5681);
or U6818 (N_6818,N_5417,N_5705);
and U6819 (N_6819,N_5895,N_5166);
nand U6820 (N_6820,N_5716,N_5356);
nand U6821 (N_6821,N_5365,N_5109);
and U6822 (N_6822,N_5299,N_5087);
xor U6823 (N_6823,N_5064,N_5285);
or U6824 (N_6824,N_5407,N_5035);
nand U6825 (N_6825,N_5955,N_5625);
or U6826 (N_6826,N_5433,N_5098);
nand U6827 (N_6827,N_5431,N_5020);
and U6828 (N_6828,N_5463,N_5416);
or U6829 (N_6829,N_5540,N_5533);
and U6830 (N_6830,N_5738,N_5951);
and U6831 (N_6831,N_5142,N_5164);
nand U6832 (N_6832,N_5955,N_5009);
or U6833 (N_6833,N_5871,N_5303);
and U6834 (N_6834,N_5547,N_5489);
or U6835 (N_6835,N_5394,N_5086);
or U6836 (N_6836,N_5433,N_5548);
nor U6837 (N_6837,N_5634,N_5482);
nor U6838 (N_6838,N_5521,N_5089);
xor U6839 (N_6839,N_5496,N_5659);
or U6840 (N_6840,N_5308,N_5561);
xnor U6841 (N_6841,N_5966,N_5917);
nor U6842 (N_6842,N_5284,N_5293);
and U6843 (N_6843,N_5004,N_5386);
nor U6844 (N_6844,N_5972,N_5037);
or U6845 (N_6845,N_5223,N_5806);
nor U6846 (N_6846,N_5405,N_5210);
nor U6847 (N_6847,N_5286,N_5323);
and U6848 (N_6848,N_5442,N_5408);
nor U6849 (N_6849,N_5655,N_5822);
nor U6850 (N_6850,N_5755,N_5911);
and U6851 (N_6851,N_5041,N_5087);
nor U6852 (N_6852,N_5889,N_5046);
and U6853 (N_6853,N_5194,N_5391);
and U6854 (N_6854,N_5875,N_5179);
nor U6855 (N_6855,N_5175,N_5698);
nand U6856 (N_6856,N_5273,N_5017);
nor U6857 (N_6857,N_5649,N_5105);
or U6858 (N_6858,N_5785,N_5592);
or U6859 (N_6859,N_5160,N_5918);
xor U6860 (N_6860,N_5160,N_5688);
nand U6861 (N_6861,N_5858,N_5469);
nand U6862 (N_6862,N_5924,N_5467);
nand U6863 (N_6863,N_5851,N_5022);
and U6864 (N_6864,N_5052,N_5539);
and U6865 (N_6865,N_5746,N_5517);
nor U6866 (N_6866,N_5297,N_5083);
nand U6867 (N_6867,N_5583,N_5734);
or U6868 (N_6868,N_5068,N_5805);
or U6869 (N_6869,N_5200,N_5575);
or U6870 (N_6870,N_5570,N_5412);
nand U6871 (N_6871,N_5205,N_5867);
or U6872 (N_6872,N_5408,N_5506);
or U6873 (N_6873,N_5442,N_5434);
and U6874 (N_6874,N_5980,N_5615);
or U6875 (N_6875,N_5356,N_5503);
nand U6876 (N_6876,N_5964,N_5999);
nor U6877 (N_6877,N_5654,N_5957);
or U6878 (N_6878,N_5966,N_5192);
or U6879 (N_6879,N_5204,N_5494);
xor U6880 (N_6880,N_5601,N_5004);
nor U6881 (N_6881,N_5010,N_5752);
xor U6882 (N_6882,N_5242,N_5594);
and U6883 (N_6883,N_5751,N_5141);
nand U6884 (N_6884,N_5101,N_5924);
or U6885 (N_6885,N_5887,N_5666);
nand U6886 (N_6886,N_5253,N_5020);
nor U6887 (N_6887,N_5658,N_5989);
or U6888 (N_6888,N_5385,N_5305);
or U6889 (N_6889,N_5770,N_5690);
or U6890 (N_6890,N_5668,N_5147);
or U6891 (N_6891,N_5696,N_5763);
nor U6892 (N_6892,N_5525,N_5862);
and U6893 (N_6893,N_5561,N_5379);
nor U6894 (N_6894,N_5290,N_5382);
or U6895 (N_6895,N_5915,N_5289);
and U6896 (N_6896,N_5268,N_5391);
nand U6897 (N_6897,N_5133,N_5757);
nor U6898 (N_6898,N_5389,N_5376);
nor U6899 (N_6899,N_5999,N_5775);
nand U6900 (N_6900,N_5222,N_5879);
nor U6901 (N_6901,N_5377,N_5715);
nor U6902 (N_6902,N_5522,N_5537);
nor U6903 (N_6903,N_5834,N_5201);
and U6904 (N_6904,N_5983,N_5859);
nand U6905 (N_6905,N_5603,N_5070);
and U6906 (N_6906,N_5476,N_5138);
and U6907 (N_6907,N_5167,N_5573);
nor U6908 (N_6908,N_5959,N_5583);
nor U6909 (N_6909,N_5698,N_5255);
or U6910 (N_6910,N_5771,N_5635);
xnor U6911 (N_6911,N_5653,N_5869);
or U6912 (N_6912,N_5722,N_5519);
and U6913 (N_6913,N_5966,N_5027);
and U6914 (N_6914,N_5324,N_5368);
or U6915 (N_6915,N_5502,N_5450);
nand U6916 (N_6916,N_5905,N_5817);
and U6917 (N_6917,N_5750,N_5905);
or U6918 (N_6918,N_5701,N_5015);
and U6919 (N_6919,N_5858,N_5562);
nor U6920 (N_6920,N_5944,N_5458);
or U6921 (N_6921,N_5534,N_5831);
and U6922 (N_6922,N_5551,N_5838);
or U6923 (N_6923,N_5415,N_5085);
nand U6924 (N_6924,N_5449,N_5344);
nand U6925 (N_6925,N_5346,N_5726);
nand U6926 (N_6926,N_5482,N_5601);
nand U6927 (N_6927,N_5773,N_5491);
xor U6928 (N_6928,N_5917,N_5184);
and U6929 (N_6929,N_5603,N_5880);
or U6930 (N_6930,N_5575,N_5919);
or U6931 (N_6931,N_5372,N_5417);
and U6932 (N_6932,N_5321,N_5568);
or U6933 (N_6933,N_5421,N_5669);
nand U6934 (N_6934,N_5564,N_5425);
and U6935 (N_6935,N_5918,N_5976);
and U6936 (N_6936,N_5127,N_5246);
and U6937 (N_6937,N_5144,N_5476);
and U6938 (N_6938,N_5653,N_5269);
nand U6939 (N_6939,N_5455,N_5683);
nand U6940 (N_6940,N_5904,N_5873);
xor U6941 (N_6941,N_5655,N_5594);
or U6942 (N_6942,N_5127,N_5105);
xnor U6943 (N_6943,N_5481,N_5416);
nand U6944 (N_6944,N_5618,N_5440);
nand U6945 (N_6945,N_5507,N_5011);
or U6946 (N_6946,N_5136,N_5255);
or U6947 (N_6947,N_5046,N_5098);
nand U6948 (N_6948,N_5430,N_5259);
and U6949 (N_6949,N_5615,N_5392);
or U6950 (N_6950,N_5851,N_5316);
and U6951 (N_6951,N_5591,N_5110);
xor U6952 (N_6952,N_5190,N_5831);
nand U6953 (N_6953,N_5145,N_5044);
nand U6954 (N_6954,N_5836,N_5822);
nor U6955 (N_6955,N_5113,N_5478);
nand U6956 (N_6956,N_5154,N_5041);
nor U6957 (N_6957,N_5680,N_5523);
nand U6958 (N_6958,N_5417,N_5938);
nor U6959 (N_6959,N_5212,N_5041);
xor U6960 (N_6960,N_5481,N_5288);
or U6961 (N_6961,N_5300,N_5608);
and U6962 (N_6962,N_5970,N_5560);
and U6963 (N_6963,N_5165,N_5972);
and U6964 (N_6964,N_5996,N_5733);
nand U6965 (N_6965,N_5609,N_5856);
or U6966 (N_6966,N_5216,N_5834);
or U6967 (N_6967,N_5106,N_5308);
xnor U6968 (N_6968,N_5850,N_5878);
and U6969 (N_6969,N_5246,N_5341);
and U6970 (N_6970,N_5702,N_5023);
nor U6971 (N_6971,N_5311,N_5078);
and U6972 (N_6972,N_5038,N_5793);
nor U6973 (N_6973,N_5817,N_5250);
or U6974 (N_6974,N_5126,N_5496);
nand U6975 (N_6975,N_5347,N_5035);
nor U6976 (N_6976,N_5709,N_5214);
nand U6977 (N_6977,N_5967,N_5307);
or U6978 (N_6978,N_5682,N_5855);
nor U6979 (N_6979,N_5128,N_5299);
nand U6980 (N_6980,N_5804,N_5144);
xnor U6981 (N_6981,N_5418,N_5845);
nand U6982 (N_6982,N_5812,N_5059);
nor U6983 (N_6983,N_5990,N_5345);
nor U6984 (N_6984,N_5317,N_5022);
xnor U6985 (N_6985,N_5468,N_5422);
and U6986 (N_6986,N_5604,N_5474);
and U6987 (N_6987,N_5391,N_5239);
or U6988 (N_6988,N_5144,N_5670);
and U6989 (N_6989,N_5968,N_5939);
and U6990 (N_6990,N_5577,N_5898);
and U6991 (N_6991,N_5478,N_5754);
and U6992 (N_6992,N_5211,N_5645);
or U6993 (N_6993,N_5724,N_5097);
xor U6994 (N_6994,N_5366,N_5258);
nand U6995 (N_6995,N_5865,N_5848);
or U6996 (N_6996,N_5454,N_5499);
or U6997 (N_6997,N_5098,N_5847);
nand U6998 (N_6998,N_5732,N_5688);
or U6999 (N_6999,N_5833,N_5867);
nand U7000 (N_7000,N_6677,N_6119);
nand U7001 (N_7001,N_6564,N_6583);
xnor U7002 (N_7002,N_6504,N_6651);
xnor U7003 (N_7003,N_6082,N_6446);
nand U7004 (N_7004,N_6840,N_6562);
or U7005 (N_7005,N_6491,N_6739);
and U7006 (N_7006,N_6737,N_6422);
or U7007 (N_7007,N_6543,N_6786);
xor U7008 (N_7008,N_6993,N_6406);
or U7009 (N_7009,N_6022,N_6478);
nand U7010 (N_7010,N_6402,N_6557);
and U7011 (N_7011,N_6820,N_6096);
and U7012 (N_7012,N_6963,N_6713);
or U7013 (N_7013,N_6642,N_6295);
nor U7014 (N_7014,N_6456,N_6091);
nor U7015 (N_7015,N_6577,N_6912);
or U7016 (N_7016,N_6596,N_6163);
nor U7017 (N_7017,N_6021,N_6113);
nand U7018 (N_7018,N_6072,N_6383);
nand U7019 (N_7019,N_6452,N_6080);
and U7020 (N_7020,N_6899,N_6857);
nor U7021 (N_7021,N_6217,N_6716);
nand U7022 (N_7022,N_6995,N_6484);
or U7023 (N_7023,N_6821,N_6767);
and U7024 (N_7024,N_6126,N_6712);
or U7025 (N_7025,N_6334,N_6549);
nand U7026 (N_7026,N_6646,N_6848);
and U7027 (N_7027,N_6950,N_6715);
and U7028 (N_7028,N_6747,N_6469);
or U7029 (N_7029,N_6523,N_6885);
nand U7030 (N_7030,N_6490,N_6903);
xnor U7031 (N_7031,N_6429,N_6224);
or U7032 (N_7032,N_6678,N_6059);
xor U7033 (N_7033,N_6172,N_6173);
nor U7034 (N_7034,N_6438,N_6033);
xor U7035 (N_7035,N_6386,N_6315);
nand U7036 (N_7036,N_6166,N_6443);
nand U7037 (N_7037,N_6893,N_6971);
or U7038 (N_7038,N_6408,N_6180);
nand U7039 (N_7039,N_6801,N_6179);
and U7040 (N_7040,N_6928,N_6140);
xor U7041 (N_7041,N_6590,N_6621);
nor U7042 (N_7042,N_6351,N_6304);
nor U7043 (N_7043,N_6322,N_6299);
nand U7044 (N_7044,N_6707,N_6718);
nand U7045 (N_7045,N_6150,N_6477);
and U7046 (N_7046,N_6637,N_6421);
nor U7047 (N_7047,N_6956,N_6155);
nand U7048 (N_7048,N_6598,N_6203);
or U7049 (N_7049,N_6953,N_6571);
and U7050 (N_7050,N_6510,N_6708);
or U7051 (N_7051,N_6145,N_6182);
nand U7052 (N_7052,N_6246,N_6257);
nor U7053 (N_7053,N_6358,N_6136);
nor U7054 (N_7054,N_6917,N_6360);
nand U7055 (N_7055,N_6281,N_6068);
nand U7056 (N_7056,N_6333,N_6536);
or U7057 (N_7057,N_6615,N_6066);
xor U7058 (N_7058,N_6003,N_6415);
nor U7059 (N_7059,N_6313,N_6768);
nand U7060 (N_7060,N_6775,N_6541);
nor U7061 (N_7061,N_6134,N_6781);
xnor U7062 (N_7062,N_6785,N_6254);
and U7063 (N_7063,N_6240,N_6178);
nor U7064 (N_7064,N_6740,N_6690);
or U7065 (N_7065,N_6978,N_6280);
and U7066 (N_7066,N_6401,N_6440);
and U7067 (N_7067,N_6326,N_6200);
nand U7068 (N_7068,N_6814,N_6578);
and U7069 (N_7069,N_6496,N_6964);
and U7070 (N_7070,N_6221,N_6389);
or U7071 (N_7071,N_6585,N_6473);
nand U7072 (N_7072,N_6976,N_6819);
or U7073 (N_7073,N_6435,N_6472);
nor U7074 (N_7074,N_6143,N_6765);
nor U7075 (N_7075,N_6808,N_6805);
or U7076 (N_7076,N_6465,N_6984);
nand U7077 (N_7077,N_6509,N_6309);
xnor U7078 (N_7078,N_6142,N_6448);
nand U7079 (N_7079,N_6584,N_6455);
nor U7080 (N_7080,N_6266,N_6243);
nor U7081 (N_7081,N_6194,N_6551);
nor U7082 (N_7082,N_6752,N_6568);
nand U7083 (N_7083,N_6366,N_6769);
nand U7084 (N_7084,N_6714,N_6486);
nor U7085 (N_7085,N_6701,N_6032);
nand U7086 (N_7086,N_6339,N_6601);
nand U7087 (N_7087,N_6547,N_6359);
xor U7088 (N_7088,N_6904,N_6973);
nor U7089 (N_7089,N_6692,N_6579);
and U7090 (N_7090,N_6555,N_6700);
nand U7091 (N_7091,N_6195,N_6397);
and U7092 (N_7092,N_6248,N_6132);
or U7093 (N_7093,N_6005,N_6336);
nand U7094 (N_7094,N_6253,N_6225);
nor U7095 (N_7095,N_6955,N_6090);
or U7096 (N_7096,N_6889,N_6611);
xor U7097 (N_7097,N_6105,N_6285);
nand U7098 (N_7098,N_6250,N_6494);
nor U7099 (N_7099,N_6234,N_6563);
nand U7100 (N_7100,N_6756,N_6791);
or U7101 (N_7101,N_6652,N_6365);
and U7102 (N_7102,N_6839,N_6325);
or U7103 (N_7103,N_6294,N_6233);
xnor U7104 (N_7104,N_6108,N_6574);
nand U7105 (N_7105,N_6048,N_6267);
nor U7106 (N_7106,N_6567,N_6927);
xnor U7107 (N_7107,N_6232,N_6444);
nand U7108 (N_7108,N_6362,N_6817);
and U7109 (N_7109,N_6260,N_6139);
and U7110 (N_7110,N_6460,N_6850);
and U7111 (N_7111,N_6025,N_6544);
and U7112 (N_7112,N_6515,N_6778);
nor U7113 (N_7113,N_6211,N_6831);
or U7114 (N_7114,N_6619,N_6844);
nand U7115 (N_7115,N_6418,N_6107);
nand U7116 (N_7116,N_6069,N_6414);
and U7117 (N_7117,N_6356,N_6898);
nor U7118 (N_7118,N_6158,N_6580);
xor U7119 (N_7119,N_6201,N_6731);
nor U7120 (N_7120,N_6487,N_6131);
and U7121 (N_7121,N_6900,N_6772);
nor U7122 (N_7122,N_6863,N_6499);
nor U7123 (N_7123,N_6968,N_6192);
and U7124 (N_7124,N_6999,N_6639);
or U7125 (N_7125,N_6015,N_6717);
or U7126 (N_7126,N_6230,N_6931);
or U7127 (N_7127,N_6057,N_6252);
xnor U7128 (N_7128,N_6582,N_6297);
or U7129 (N_7129,N_6554,N_6560);
nor U7130 (N_7130,N_6908,N_6783);
and U7131 (N_7131,N_6942,N_6007);
nand U7132 (N_7132,N_6761,N_6753);
nand U7133 (N_7133,N_6895,N_6745);
nand U7134 (N_7134,N_6332,N_6502);
or U7135 (N_7135,N_6390,N_6017);
xnor U7136 (N_7136,N_6676,N_6771);
or U7137 (N_7137,N_6559,N_6860);
or U7138 (N_7138,N_6065,N_6018);
nor U7139 (N_7139,N_6102,N_6667);
and U7140 (N_7140,N_6736,N_6866);
nand U7141 (N_7141,N_6097,N_6937);
or U7142 (N_7142,N_6875,N_6788);
xor U7143 (N_7143,N_6608,N_6321);
and U7144 (N_7144,N_6529,N_6770);
nor U7145 (N_7145,N_6933,N_6540);
and U7146 (N_7146,N_6877,N_6610);
nor U7147 (N_7147,N_6659,N_6123);
and U7148 (N_7148,N_6011,N_6990);
nand U7149 (N_7149,N_6935,N_6640);
xor U7150 (N_7150,N_6573,N_6614);
xor U7151 (N_7151,N_6241,N_6884);
and U7152 (N_7152,N_6095,N_6666);
nor U7153 (N_7153,N_6330,N_6498);
and U7154 (N_7154,N_6974,N_6532);
nand U7155 (N_7155,N_6635,N_6067);
nand U7156 (N_7156,N_6843,N_6597);
xnor U7157 (N_7157,N_6255,N_6062);
nand U7158 (N_7158,N_6570,N_6115);
nand U7159 (N_7159,N_6865,N_6023);
xnor U7160 (N_7160,N_6988,N_6682);
nand U7161 (N_7161,N_6897,N_6288);
and U7162 (N_7162,N_6355,N_6924);
nand U7163 (N_7163,N_6689,N_6374);
or U7164 (N_7164,N_6835,N_6849);
nor U7165 (N_7165,N_6156,N_6874);
xnor U7166 (N_7166,N_6101,N_6871);
or U7167 (N_7167,N_6471,N_6319);
nand U7168 (N_7168,N_6705,N_6109);
nor U7169 (N_7169,N_6467,N_6436);
or U7170 (N_7170,N_6760,N_6349);
nor U7171 (N_7171,N_6409,N_6357);
nor U7172 (N_7172,N_6363,N_6275);
or U7173 (N_7173,N_6980,N_6873);
nor U7174 (N_7174,N_6000,N_6581);
or U7175 (N_7175,N_6946,N_6034);
and U7176 (N_7176,N_6479,N_6671);
nand U7177 (N_7177,N_6214,N_6948);
and U7178 (N_7178,N_6149,N_6704);
nand U7179 (N_7179,N_6348,N_6957);
nor U7180 (N_7180,N_6012,N_6633);
or U7181 (N_7181,N_6038,N_6774);
or U7182 (N_7182,N_6982,N_6437);
and U7183 (N_7183,N_6604,N_6388);
nand U7184 (N_7184,N_6238,N_6392);
nor U7185 (N_7185,N_6511,N_6047);
and U7186 (N_7186,N_6181,N_6077);
nand U7187 (N_7187,N_6493,N_6036);
nor U7188 (N_7188,N_6335,N_6694);
nor U7189 (N_7189,N_6991,N_6174);
and U7190 (N_7190,N_6894,N_6412);
nor U7191 (N_7191,N_6237,N_6273);
or U7192 (N_7192,N_6169,N_6847);
nor U7193 (N_7193,N_6395,N_6272);
nor U7194 (N_7194,N_6447,N_6699);
and U7195 (N_7195,N_6430,N_6734);
nor U7196 (N_7196,N_6074,N_6996);
nand U7197 (N_7197,N_6328,N_6782);
nand U7198 (N_7198,N_6944,N_6079);
nor U7199 (N_7199,N_6528,N_6787);
or U7200 (N_7200,N_6997,N_6475);
and U7201 (N_7201,N_6028,N_6235);
nor U7202 (N_7202,N_6063,N_6223);
and U7203 (N_7203,N_6723,N_6265);
xnor U7204 (N_7204,N_6852,N_6810);
and U7205 (N_7205,N_6277,N_6725);
nand U7206 (N_7206,N_6104,N_6656);
nand U7207 (N_7207,N_6915,N_6624);
nor U7208 (N_7208,N_6279,N_6816);
nand U7209 (N_7209,N_6492,N_6306);
and U7210 (N_7210,N_6052,N_6367);
or U7211 (N_7211,N_6416,N_6683);
nor U7212 (N_7212,N_6301,N_6433);
nor U7213 (N_7213,N_6684,N_6364);
nor U7214 (N_7214,N_6981,N_6879);
xnor U7215 (N_7215,N_6797,N_6673);
nand U7216 (N_7216,N_6858,N_6014);
nor U7217 (N_7217,N_6445,N_6645);
nor U7218 (N_7218,N_6337,N_6545);
and U7219 (N_7219,N_6868,N_6943);
and U7220 (N_7220,N_6229,N_6722);
nand U7221 (N_7221,N_6594,N_6586);
and U7222 (N_7222,N_6258,N_6076);
or U7223 (N_7223,N_6878,N_6343);
xnor U7224 (N_7224,N_6081,N_6271);
nor U7225 (N_7225,N_6249,N_6176);
nand U7226 (N_7226,N_6561,N_6861);
xor U7227 (N_7227,N_6970,N_6087);
nor U7228 (N_7228,N_6110,N_6815);
or U7229 (N_7229,N_6071,N_6576);
nand U7230 (N_7230,N_6552,N_6311);
nor U7231 (N_7231,N_6754,N_6727);
and U7232 (N_7232,N_6481,N_6051);
xor U7233 (N_7233,N_6157,N_6009);
nor U7234 (N_7234,N_6757,N_6830);
nor U7235 (N_7235,N_6167,N_6353);
and U7236 (N_7236,N_6983,N_6887);
xnor U7237 (N_7237,N_6381,N_6043);
or U7238 (N_7238,N_6135,N_6083);
nand U7239 (N_7239,N_6199,N_6368);
xnor U7240 (N_7240,N_6114,N_6521);
nand U7241 (N_7241,N_6064,N_6451);
xnor U7242 (N_7242,N_6245,N_6985);
nand U7243 (N_7243,N_6269,N_6688);
nor U7244 (N_7244,N_6729,N_6662);
nand U7245 (N_7245,N_6175,N_6599);
xor U7246 (N_7246,N_6385,N_6869);
and U7247 (N_7247,N_6376,N_6546);
nor U7248 (N_7248,N_6159,N_6453);
xnor U7249 (N_7249,N_6605,N_6751);
nor U7250 (N_7250,N_6346,N_6458);
nor U7251 (N_7251,N_6949,N_6958);
and U7252 (N_7252,N_6724,N_6361);
and U7253 (N_7253,N_6539,N_6161);
and U7254 (N_7254,N_6212,N_6035);
and U7255 (N_7255,N_6213,N_6439);
nand U7256 (N_7256,N_6204,N_6932);
or U7257 (N_7257,N_6384,N_6296);
or U7258 (N_7258,N_6117,N_6653);
and U7259 (N_7259,N_6634,N_6118);
and U7260 (N_7260,N_6314,N_6403);
xnor U7261 (N_7261,N_6764,N_6324);
and U7262 (N_7262,N_6647,N_6426);
nand U7263 (N_7263,N_6218,N_6587);
nand U7264 (N_7264,N_6901,N_6709);
nor U7265 (N_7265,N_6058,N_6298);
xnor U7266 (N_7266,N_6940,N_6482);
or U7267 (N_7267,N_6607,N_6987);
and U7268 (N_7268,N_6922,N_6603);
or U7269 (N_7269,N_6489,N_6525);
nor U7270 (N_7270,N_6538,N_6806);
and U7271 (N_7271,N_6641,N_6872);
or U7272 (N_7272,N_6530,N_6404);
xnor U7273 (N_7273,N_6124,N_6372);
or U7274 (N_7274,N_6154,N_6189);
nand U7275 (N_7275,N_6312,N_6193);
nand U7276 (N_7276,N_6111,N_6289);
nand U7277 (N_7277,N_6292,N_6670);
nand U7278 (N_7278,N_6784,N_6503);
nand U7279 (N_7279,N_6303,N_6907);
or U7280 (N_7280,N_6674,N_6405);
nand U7281 (N_7281,N_6242,N_6088);
nor U7282 (N_7282,N_6146,N_6205);
and U7283 (N_7283,N_6345,N_6799);
nand U7284 (N_7284,N_6986,N_6016);
nand U7285 (N_7285,N_6160,N_6413);
and U7286 (N_7286,N_6720,N_6672);
xor U7287 (N_7287,N_6829,N_6954);
and U7288 (N_7288,N_6120,N_6896);
nor U7289 (N_7289,N_6291,N_6410);
nand U7290 (N_7290,N_6377,N_6263);
or U7291 (N_7291,N_6270,N_6780);
or U7292 (N_7292,N_6612,N_6951);
nor U7293 (N_7293,N_6268,N_6735);
and U7294 (N_7294,N_6627,N_6459);
and U7295 (N_7295,N_6046,N_6882);
nor U7296 (N_7296,N_6206,N_6902);
and U7297 (N_7297,N_6053,N_6251);
nand U7298 (N_7298,N_6183,N_6909);
nor U7299 (N_7299,N_6941,N_6750);
or U7300 (N_7300,N_6329,N_6137);
or U7301 (N_7301,N_6049,N_6476);
xor U7302 (N_7302,N_6696,N_6247);
and U7303 (N_7303,N_6441,N_6827);
or U7304 (N_7304,N_6870,N_6282);
nand U7305 (N_7305,N_6450,N_6106);
and U7306 (N_7306,N_6828,N_6762);
and U7307 (N_7307,N_6026,N_6226);
or U7308 (N_7308,N_6196,N_6024);
or U7309 (N_7309,N_6616,N_6084);
nand U7310 (N_7310,N_6618,N_6029);
nor U7311 (N_7311,N_6379,N_6045);
nand U7312 (N_7312,N_6170,N_6638);
and U7313 (N_7313,N_6338,N_6862);
or U7314 (N_7314,N_6595,N_6613);
or U7315 (N_7315,N_6936,N_6202);
xor U7316 (N_7316,N_6396,N_6151);
and U7317 (N_7317,N_6055,N_6207);
and U7318 (N_7318,N_6125,N_6112);
and U7319 (N_7319,N_6864,N_6210);
or U7320 (N_7320,N_6042,N_6308);
and U7321 (N_7321,N_6141,N_6350);
nor U7322 (N_7322,N_6556,N_6620);
and U7323 (N_7323,N_6378,N_6320);
and U7324 (N_7324,N_6663,N_6960);
nand U7325 (N_7325,N_6470,N_6811);
nor U7326 (N_7326,N_6209,N_6906);
nand U7327 (N_7327,N_6758,N_6913);
and U7328 (N_7328,N_6888,N_6220);
or U7329 (N_7329,N_6128,N_6431);
nand U7330 (N_7330,N_6041,N_6890);
nor U7331 (N_7331,N_6919,N_6305);
and U7332 (N_7332,N_6462,N_6256);
or U7333 (N_7333,N_6457,N_6732);
xnor U7334 (N_7334,N_6216,N_6449);
nand U7335 (N_7335,N_6741,N_6380);
nor U7336 (N_7336,N_6733,N_6524);
and U7337 (N_7337,N_6773,N_6880);
nand U7338 (N_7338,N_6500,N_6191);
xor U7339 (N_7339,N_6698,N_6188);
nand U7340 (N_7340,N_6798,N_6507);
nand U7341 (N_7341,N_6693,N_6979);
or U7342 (N_7342,N_6075,N_6914);
nor U7343 (N_7343,N_6592,N_6755);
and U7344 (N_7344,N_6061,N_6854);
nor U7345 (N_7345,N_6373,N_6420);
and U7346 (N_7346,N_6628,N_6056);
nor U7347 (N_7347,N_6144,N_6794);
and U7348 (N_7348,N_6691,N_6466);
and U7349 (N_7349,N_6636,N_6961);
and U7350 (N_7350,N_6534,N_6920);
xnor U7351 (N_7351,N_6276,N_6040);
xnor U7352 (N_7352,N_6905,N_6965);
and U7353 (N_7353,N_6442,N_6197);
nor U7354 (N_7354,N_6514,N_6759);
or U7355 (N_7355,N_6044,N_6650);
and U7356 (N_7356,N_6148,N_6630);
and U7357 (N_7357,N_6967,N_6800);
and U7358 (N_7358,N_6654,N_6632);
nand U7359 (N_7359,N_6369,N_6742);
or U7360 (N_7360,N_6186,N_6929);
nor U7361 (N_7361,N_6548,N_6501);
or U7362 (N_7362,N_6975,N_6341);
and U7363 (N_7363,N_6461,N_6394);
nand U7364 (N_7364,N_6177,N_6851);
nor U7365 (N_7365,N_6994,N_6842);
and U7366 (N_7366,N_6803,N_6208);
or U7367 (N_7367,N_6558,N_6001);
and U7368 (N_7368,N_6911,N_6977);
nor U7369 (N_7369,N_6721,N_6290);
or U7370 (N_7370,N_6841,N_6728);
or U7371 (N_7371,N_6886,N_6531);
or U7372 (N_7372,N_6591,N_6286);
nor U7373 (N_7373,N_6030,N_6938);
and U7374 (N_7374,N_6726,N_6744);
nand U7375 (N_7375,N_6138,N_6262);
and U7376 (N_7376,N_6317,N_6520);
or U7377 (N_7377,N_6427,N_6657);
or U7378 (N_7378,N_6488,N_6644);
and U7379 (N_7379,N_6008,N_6130);
nor U7380 (N_7380,N_6164,N_6660);
nand U7381 (N_7381,N_6278,N_6763);
nor U7382 (N_7382,N_6400,N_6483);
nand U7383 (N_7383,N_6832,N_6078);
and U7384 (N_7384,N_6687,N_6428);
or U7385 (N_7385,N_6089,N_6506);
nor U7386 (N_7386,N_6399,N_6809);
nand U7387 (N_7387,N_6347,N_6789);
and U7388 (N_7388,N_6398,N_6454);
or U7389 (N_7389,N_6575,N_6103);
xnor U7390 (N_7390,N_6122,N_6992);
or U7391 (N_7391,N_6092,N_6617);
nand U7392 (N_7392,N_6855,N_6921);
nor U7393 (N_7393,N_6287,N_6463);
nand U7394 (N_7394,N_6050,N_6846);
nor U7395 (N_7395,N_6190,N_6316);
nand U7396 (N_7396,N_6681,N_6474);
nand U7397 (N_7397,N_6926,N_6686);
and U7398 (N_7398,N_6464,N_6411);
or U7399 (N_7399,N_6836,N_6168);
nor U7400 (N_7400,N_6962,N_6790);
or U7401 (N_7401,N_6031,N_6318);
or U7402 (N_7402,N_6236,N_6925);
xor U7403 (N_7403,N_6039,N_6609);
nor U7404 (N_7404,N_6152,N_6432);
nand U7405 (N_7405,N_6845,N_6572);
and U7406 (N_7406,N_6323,N_6658);
or U7407 (N_7407,N_6513,N_6093);
and U7408 (N_7408,N_6434,N_6833);
nor U7409 (N_7409,N_6812,N_6244);
or U7410 (N_7410,N_6792,N_6505);
and U7411 (N_7411,N_6824,N_6382);
xnor U7412 (N_7412,N_6934,N_6661);
and U7413 (N_7413,N_6517,N_6004);
and U7414 (N_7414,N_6300,N_6099);
nor U7415 (N_7415,N_6054,N_6537);
xnor U7416 (N_7416,N_6825,N_6804);
and U7417 (N_7417,N_6606,N_6533);
or U7418 (N_7418,N_6593,N_6129);
nand U7419 (N_7419,N_6837,N_6668);
nor U7420 (N_7420,N_6675,N_6302);
and U7421 (N_7421,N_6649,N_6730);
xnor U7422 (N_7422,N_6834,N_6133);
nor U7423 (N_7423,N_6340,N_6629);
nand U7424 (N_7424,N_6966,N_6655);
nand U7425 (N_7425,N_6264,N_6766);
or U7426 (N_7426,N_6969,N_6147);
and U7427 (N_7427,N_6085,N_6697);
or U7428 (N_7428,N_6749,N_6779);
nand U7429 (N_7429,N_6187,N_6989);
and U7430 (N_7430,N_6519,N_6823);
nand U7431 (N_7431,N_6738,N_6526);
or U7432 (N_7432,N_6518,N_6227);
nor U7433 (N_7433,N_6910,N_6952);
nor U7434 (N_7434,N_6284,N_6086);
and U7435 (N_7435,N_6480,N_6883);
xor U7436 (N_7436,N_6945,N_6622);
nand U7437 (N_7437,N_6859,N_6522);
and U7438 (N_7438,N_6121,N_6795);
or U7439 (N_7439,N_6665,N_6527);
nand U7440 (N_7440,N_6391,N_6261);
or U7441 (N_7441,N_6239,N_6019);
nand U7442 (N_7442,N_6198,N_6070);
nand U7443 (N_7443,N_6274,N_6485);
and U7444 (N_7444,N_6838,N_6094);
or U7445 (N_7445,N_6807,N_6387);
and U7446 (N_7446,N_6425,N_6939);
and U7447 (N_7447,N_6959,N_6853);
and U7448 (N_7448,N_6802,N_6695);
nand U7449 (N_7449,N_6370,N_6891);
nor U7450 (N_7450,N_6664,N_6669);
xor U7451 (N_7451,N_6231,N_6535);
and U7452 (N_7452,N_6947,N_6037);
nor U7453 (N_7453,N_6127,N_6998);
or U7454 (N_7454,N_6916,N_6293);
nor U7455 (N_7455,N_6215,N_6424);
nor U7456 (N_7456,N_6569,N_6685);
nand U7457 (N_7457,N_6027,N_6116);
and U7458 (N_7458,N_6352,N_6495);
nand U7459 (N_7459,N_6918,N_6793);
or U7460 (N_7460,N_6002,N_6098);
nand U7461 (N_7461,N_6972,N_6228);
and U7462 (N_7462,N_6867,N_6375);
or U7463 (N_7463,N_6648,N_6776);
nor U7464 (N_7464,N_6344,N_6856);
or U7465 (N_7465,N_6566,N_6826);
nand U7466 (N_7466,N_6219,N_6719);
nand U7467 (N_7467,N_6407,N_6073);
nand U7468 (N_7468,N_6743,N_6354);
and U7469 (N_7469,N_6010,N_6625);
or U7470 (N_7470,N_6818,N_6060);
or U7471 (N_7471,N_6331,N_6393);
nor U7472 (N_7472,N_6813,N_6680);
and U7473 (N_7473,N_6006,N_6165);
or U7474 (N_7474,N_6930,N_6923);
nand U7475 (N_7475,N_6542,N_6748);
xnor U7476 (N_7476,N_6553,N_6631);
nor U7477 (N_7477,N_6876,N_6777);
and U7478 (N_7478,N_6679,N_6600);
or U7479 (N_7479,N_6419,N_6565);
nand U7480 (N_7480,N_6259,N_6307);
or U7481 (N_7481,N_6283,N_6643);
nand U7482 (N_7482,N_6162,N_6417);
xnor U7483 (N_7483,N_6100,N_6710);
nor U7484 (N_7484,N_6516,N_6746);
and U7485 (N_7485,N_6822,N_6508);
and U7486 (N_7486,N_6706,N_6703);
nor U7487 (N_7487,N_6153,N_6892);
and U7488 (N_7488,N_6310,N_6184);
and U7489 (N_7489,N_6512,N_6588);
nor U7490 (N_7490,N_6423,N_6013);
nand U7491 (N_7491,N_6623,N_6626);
xnor U7492 (N_7492,N_6327,N_6602);
and U7493 (N_7493,N_6185,N_6711);
nor U7494 (N_7494,N_6796,N_6371);
nor U7495 (N_7495,N_6468,N_6497);
xor U7496 (N_7496,N_6171,N_6222);
nand U7497 (N_7497,N_6702,N_6589);
and U7498 (N_7498,N_6550,N_6020);
nand U7499 (N_7499,N_6881,N_6342);
xnor U7500 (N_7500,N_6183,N_6410);
nand U7501 (N_7501,N_6256,N_6411);
nor U7502 (N_7502,N_6092,N_6087);
nand U7503 (N_7503,N_6901,N_6928);
nand U7504 (N_7504,N_6490,N_6296);
and U7505 (N_7505,N_6821,N_6063);
and U7506 (N_7506,N_6518,N_6008);
nor U7507 (N_7507,N_6470,N_6681);
nand U7508 (N_7508,N_6558,N_6533);
or U7509 (N_7509,N_6284,N_6714);
or U7510 (N_7510,N_6984,N_6278);
or U7511 (N_7511,N_6545,N_6050);
or U7512 (N_7512,N_6576,N_6783);
xnor U7513 (N_7513,N_6458,N_6812);
nand U7514 (N_7514,N_6221,N_6023);
nand U7515 (N_7515,N_6904,N_6649);
xnor U7516 (N_7516,N_6479,N_6621);
or U7517 (N_7517,N_6462,N_6000);
and U7518 (N_7518,N_6858,N_6873);
nor U7519 (N_7519,N_6119,N_6024);
xnor U7520 (N_7520,N_6644,N_6348);
xnor U7521 (N_7521,N_6302,N_6075);
nor U7522 (N_7522,N_6447,N_6920);
nor U7523 (N_7523,N_6813,N_6580);
and U7524 (N_7524,N_6211,N_6828);
nor U7525 (N_7525,N_6192,N_6049);
and U7526 (N_7526,N_6918,N_6939);
nand U7527 (N_7527,N_6966,N_6545);
and U7528 (N_7528,N_6544,N_6867);
and U7529 (N_7529,N_6060,N_6382);
or U7530 (N_7530,N_6215,N_6792);
and U7531 (N_7531,N_6164,N_6736);
and U7532 (N_7532,N_6475,N_6577);
and U7533 (N_7533,N_6860,N_6996);
nand U7534 (N_7534,N_6837,N_6486);
nand U7535 (N_7535,N_6750,N_6967);
nor U7536 (N_7536,N_6492,N_6159);
nor U7537 (N_7537,N_6580,N_6824);
nand U7538 (N_7538,N_6692,N_6928);
nand U7539 (N_7539,N_6081,N_6334);
or U7540 (N_7540,N_6888,N_6897);
xnor U7541 (N_7541,N_6324,N_6371);
and U7542 (N_7542,N_6304,N_6449);
nor U7543 (N_7543,N_6166,N_6044);
or U7544 (N_7544,N_6327,N_6733);
and U7545 (N_7545,N_6873,N_6386);
nor U7546 (N_7546,N_6073,N_6673);
nand U7547 (N_7547,N_6827,N_6783);
or U7548 (N_7548,N_6380,N_6198);
nor U7549 (N_7549,N_6935,N_6081);
nor U7550 (N_7550,N_6526,N_6996);
xor U7551 (N_7551,N_6292,N_6924);
or U7552 (N_7552,N_6944,N_6156);
nor U7553 (N_7553,N_6606,N_6484);
or U7554 (N_7554,N_6226,N_6884);
nand U7555 (N_7555,N_6322,N_6872);
and U7556 (N_7556,N_6217,N_6422);
nor U7557 (N_7557,N_6732,N_6100);
xnor U7558 (N_7558,N_6411,N_6796);
or U7559 (N_7559,N_6615,N_6792);
nor U7560 (N_7560,N_6848,N_6952);
or U7561 (N_7561,N_6067,N_6455);
or U7562 (N_7562,N_6388,N_6772);
and U7563 (N_7563,N_6076,N_6750);
and U7564 (N_7564,N_6136,N_6083);
and U7565 (N_7565,N_6392,N_6947);
nor U7566 (N_7566,N_6431,N_6163);
or U7567 (N_7567,N_6587,N_6188);
xor U7568 (N_7568,N_6449,N_6477);
nor U7569 (N_7569,N_6547,N_6966);
or U7570 (N_7570,N_6275,N_6547);
nor U7571 (N_7571,N_6924,N_6162);
xor U7572 (N_7572,N_6967,N_6415);
and U7573 (N_7573,N_6973,N_6029);
nand U7574 (N_7574,N_6708,N_6418);
nor U7575 (N_7575,N_6011,N_6069);
nand U7576 (N_7576,N_6723,N_6198);
or U7577 (N_7577,N_6119,N_6352);
nand U7578 (N_7578,N_6553,N_6224);
nand U7579 (N_7579,N_6753,N_6408);
nand U7580 (N_7580,N_6474,N_6680);
xnor U7581 (N_7581,N_6622,N_6978);
or U7582 (N_7582,N_6845,N_6574);
nor U7583 (N_7583,N_6980,N_6567);
nor U7584 (N_7584,N_6612,N_6953);
nand U7585 (N_7585,N_6111,N_6744);
or U7586 (N_7586,N_6126,N_6721);
nor U7587 (N_7587,N_6362,N_6155);
nand U7588 (N_7588,N_6807,N_6332);
nor U7589 (N_7589,N_6631,N_6346);
and U7590 (N_7590,N_6460,N_6680);
nor U7591 (N_7591,N_6931,N_6294);
or U7592 (N_7592,N_6605,N_6824);
or U7593 (N_7593,N_6913,N_6011);
nand U7594 (N_7594,N_6330,N_6980);
nor U7595 (N_7595,N_6758,N_6384);
or U7596 (N_7596,N_6771,N_6526);
or U7597 (N_7597,N_6774,N_6878);
or U7598 (N_7598,N_6532,N_6947);
and U7599 (N_7599,N_6555,N_6946);
or U7600 (N_7600,N_6754,N_6423);
nor U7601 (N_7601,N_6224,N_6351);
or U7602 (N_7602,N_6464,N_6804);
nand U7603 (N_7603,N_6189,N_6551);
or U7604 (N_7604,N_6752,N_6334);
nand U7605 (N_7605,N_6596,N_6055);
or U7606 (N_7606,N_6864,N_6193);
and U7607 (N_7607,N_6833,N_6056);
and U7608 (N_7608,N_6066,N_6993);
nand U7609 (N_7609,N_6429,N_6422);
xnor U7610 (N_7610,N_6737,N_6319);
xor U7611 (N_7611,N_6790,N_6606);
nor U7612 (N_7612,N_6613,N_6978);
nand U7613 (N_7613,N_6349,N_6121);
nand U7614 (N_7614,N_6908,N_6421);
xnor U7615 (N_7615,N_6948,N_6731);
and U7616 (N_7616,N_6172,N_6164);
or U7617 (N_7617,N_6489,N_6869);
nand U7618 (N_7618,N_6690,N_6426);
or U7619 (N_7619,N_6553,N_6668);
or U7620 (N_7620,N_6088,N_6263);
or U7621 (N_7621,N_6955,N_6323);
nand U7622 (N_7622,N_6788,N_6445);
and U7623 (N_7623,N_6925,N_6660);
or U7624 (N_7624,N_6761,N_6790);
nor U7625 (N_7625,N_6330,N_6236);
nor U7626 (N_7626,N_6151,N_6353);
or U7627 (N_7627,N_6077,N_6180);
xor U7628 (N_7628,N_6022,N_6593);
nand U7629 (N_7629,N_6767,N_6029);
and U7630 (N_7630,N_6960,N_6345);
or U7631 (N_7631,N_6159,N_6389);
or U7632 (N_7632,N_6273,N_6101);
nand U7633 (N_7633,N_6921,N_6025);
nand U7634 (N_7634,N_6046,N_6023);
and U7635 (N_7635,N_6812,N_6560);
and U7636 (N_7636,N_6891,N_6246);
and U7637 (N_7637,N_6898,N_6127);
nor U7638 (N_7638,N_6472,N_6256);
nand U7639 (N_7639,N_6244,N_6519);
nand U7640 (N_7640,N_6126,N_6768);
nor U7641 (N_7641,N_6865,N_6348);
and U7642 (N_7642,N_6308,N_6136);
nand U7643 (N_7643,N_6007,N_6734);
xor U7644 (N_7644,N_6559,N_6654);
xor U7645 (N_7645,N_6249,N_6788);
nor U7646 (N_7646,N_6907,N_6838);
nand U7647 (N_7647,N_6458,N_6374);
and U7648 (N_7648,N_6000,N_6611);
nand U7649 (N_7649,N_6642,N_6241);
or U7650 (N_7650,N_6761,N_6663);
and U7651 (N_7651,N_6659,N_6183);
nand U7652 (N_7652,N_6579,N_6277);
nor U7653 (N_7653,N_6811,N_6115);
xor U7654 (N_7654,N_6755,N_6214);
and U7655 (N_7655,N_6932,N_6924);
nand U7656 (N_7656,N_6685,N_6236);
or U7657 (N_7657,N_6450,N_6519);
xor U7658 (N_7658,N_6274,N_6555);
and U7659 (N_7659,N_6780,N_6310);
and U7660 (N_7660,N_6499,N_6814);
xnor U7661 (N_7661,N_6969,N_6093);
or U7662 (N_7662,N_6107,N_6161);
xnor U7663 (N_7663,N_6529,N_6440);
xor U7664 (N_7664,N_6133,N_6830);
and U7665 (N_7665,N_6856,N_6205);
xor U7666 (N_7666,N_6849,N_6334);
nand U7667 (N_7667,N_6017,N_6666);
or U7668 (N_7668,N_6389,N_6225);
nand U7669 (N_7669,N_6459,N_6747);
and U7670 (N_7670,N_6380,N_6121);
nand U7671 (N_7671,N_6434,N_6804);
or U7672 (N_7672,N_6978,N_6802);
or U7673 (N_7673,N_6594,N_6578);
or U7674 (N_7674,N_6403,N_6346);
and U7675 (N_7675,N_6915,N_6850);
xnor U7676 (N_7676,N_6511,N_6584);
and U7677 (N_7677,N_6034,N_6361);
xor U7678 (N_7678,N_6503,N_6650);
or U7679 (N_7679,N_6641,N_6436);
and U7680 (N_7680,N_6102,N_6197);
xor U7681 (N_7681,N_6306,N_6830);
and U7682 (N_7682,N_6656,N_6484);
or U7683 (N_7683,N_6549,N_6792);
nand U7684 (N_7684,N_6720,N_6423);
and U7685 (N_7685,N_6141,N_6532);
nor U7686 (N_7686,N_6314,N_6777);
and U7687 (N_7687,N_6054,N_6913);
and U7688 (N_7688,N_6730,N_6936);
nand U7689 (N_7689,N_6145,N_6011);
nor U7690 (N_7690,N_6208,N_6312);
nand U7691 (N_7691,N_6384,N_6025);
nand U7692 (N_7692,N_6405,N_6418);
nor U7693 (N_7693,N_6160,N_6767);
nand U7694 (N_7694,N_6989,N_6024);
nand U7695 (N_7695,N_6851,N_6576);
or U7696 (N_7696,N_6928,N_6358);
and U7697 (N_7697,N_6306,N_6486);
nor U7698 (N_7698,N_6345,N_6668);
and U7699 (N_7699,N_6973,N_6448);
nor U7700 (N_7700,N_6757,N_6173);
or U7701 (N_7701,N_6700,N_6444);
nor U7702 (N_7702,N_6090,N_6081);
or U7703 (N_7703,N_6229,N_6633);
nor U7704 (N_7704,N_6345,N_6544);
and U7705 (N_7705,N_6606,N_6122);
and U7706 (N_7706,N_6845,N_6982);
nand U7707 (N_7707,N_6008,N_6167);
or U7708 (N_7708,N_6324,N_6339);
nand U7709 (N_7709,N_6847,N_6500);
or U7710 (N_7710,N_6600,N_6336);
or U7711 (N_7711,N_6565,N_6740);
nor U7712 (N_7712,N_6421,N_6589);
nand U7713 (N_7713,N_6209,N_6439);
xor U7714 (N_7714,N_6410,N_6598);
or U7715 (N_7715,N_6113,N_6199);
and U7716 (N_7716,N_6268,N_6561);
nor U7717 (N_7717,N_6240,N_6292);
nand U7718 (N_7718,N_6610,N_6457);
or U7719 (N_7719,N_6003,N_6900);
and U7720 (N_7720,N_6202,N_6303);
nand U7721 (N_7721,N_6198,N_6460);
nor U7722 (N_7722,N_6818,N_6470);
nand U7723 (N_7723,N_6486,N_6516);
or U7724 (N_7724,N_6098,N_6198);
xor U7725 (N_7725,N_6776,N_6553);
xor U7726 (N_7726,N_6967,N_6949);
or U7727 (N_7727,N_6419,N_6112);
nor U7728 (N_7728,N_6651,N_6999);
nor U7729 (N_7729,N_6768,N_6273);
nand U7730 (N_7730,N_6446,N_6743);
or U7731 (N_7731,N_6723,N_6029);
nor U7732 (N_7732,N_6868,N_6769);
nor U7733 (N_7733,N_6094,N_6968);
nand U7734 (N_7734,N_6810,N_6591);
and U7735 (N_7735,N_6915,N_6845);
and U7736 (N_7736,N_6962,N_6240);
or U7737 (N_7737,N_6222,N_6218);
and U7738 (N_7738,N_6622,N_6348);
or U7739 (N_7739,N_6856,N_6365);
or U7740 (N_7740,N_6812,N_6815);
nand U7741 (N_7741,N_6882,N_6947);
or U7742 (N_7742,N_6899,N_6284);
nor U7743 (N_7743,N_6273,N_6295);
and U7744 (N_7744,N_6966,N_6199);
xor U7745 (N_7745,N_6851,N_6662);
or U7746 (N_7746,N_6780,N_6508);
nor U7747 (N_7747,N_6931,N_6343);
xnor U7748 (N_7748,N_6055,N_6759);
and U7749 (N_7749,N_6026,N_6211);
nor U7750 (N_7750,N_6158,N_6592);
or U7751 (N_7751,N_6955,N_6695);
and U7752 (N_7752,N_6266,N_6185);
or U7753 (N_7753,N_6330,N_6141);
or U7754 (N_7754,N_6880,N_6886);
nor U7755 (N_7755,N_6830,N_6829);
nand U7756 (N_7756,N_6528,N_6517);
or U7757 (N_7757,N_6895,N_6188);
nand U7758 (N_7758,N_6880,N_6482);
nor U7759 (N_7759,N_6336,N_6311);
and U7760 (N_7760,N_6774,N_6081);
nand U7761 (N_7761,N_6529,N_6684);
nand U7762 (N_7762,N_6239,N_6202);
or U7763 (N_7763,N_6126,N_6865);
xnor U7764 (N_7764,N_6043,N_6036);
xor U7765 (N_7765,N_6396,N_6572);
or U7766 (N_7766,N_6045,N_6155);
xnor U7767 (N_7767,N_6839,N_6930);
nand U7768 (N_7768,N_6196,N_6794);
nor U7769 (N_7769,N_6547,N_6180);
nand U7770 (N_7770,N_6260,N_6537);
or U7771 (N_7771,N_6531,N_6092);
and U7772 (N_7772,N_6448,N_6324);
xnor U7773 (N_7773,N_6748,N_6089);
nor U7774 (N_7774,N_6272,N_6099);
nor U7775 (N_7775,N_6101,N_6473);
nor U7776 (N_7776,N_6448,N_6905);
or U7777 (N_7777,N_6578,N_6972);
and U7778 (N_7778,N_6374,N_6788);
and U7779 (N_7779,N_6605,N_6322);
nand U7780 (N_7780,N_6385,N_6411);
nand U7781 (N_7781,N_6210,N_6823);
or U7782 (N_7782,N_6805,N_6963);
and U7783 (N_7783,N_6649,N_6384);
and U7784 (N_7784,N_6957,N_6571);
or U7785 (N_7785,N_6474,N_6289);
nor U7786 (N_7786,N_6032,N_6290);
xnor U7787 (N_7787,N_6224,N_6576);
nand U7788 (N_7788,N_6555,N_6575);
and U7789 (N_7789,N_6921,N_6572);
or U7790 (N_7790,N_6350,N_6311);
xnor U7791 (N_7791,N_6776,N_6108);
nor U7792 (N_7792,N_6461,N_6381);
xnor U7793 (N_7793,N_6487,N_6684);
and U7794 (N_7794,N_6607,N_6837);
nor U7795 (N_7795,N_6689,N_6917);
nor U7796 (N_7796,N_6172,N_6890);
xnor U7797 (N_7797,N_6071,N_6284);
nor U7798 (N_7798,N_6483,N_6741);
nor U7799 (N_7799,N_6326,N_6441);
xnor U7800 (N_7800,N_6402,N_6731);
xnor U7801 (N_7801,N_6463,N_6802);
nand U7802 (N_7802,N_6798,N_6257);
or U7803 (N_7803,N_6938,N_6546);
nand U7804 (N_7804,N_6214,N_6709);
nand U7805 (N_7805,N_6832,N_6027);
nor U7806 (N_7806,N_6406,N_6245);
or U7807 (N_7807,N_6833,N_6604);
nand U7808 (N_7808,N_6311,N_6764);
nor U7809 (N_7809,N_6775,N_6003);
xor U7810 (N_7810,N_6994,N_6645);
or U7811 (N_7811,N_6190,N_6443);
xnor U7812 (N_7812,N_6296,N_6658);
nor U7813 (N_7813,N_6512,N_6327);
xnor U7814 (N_7814,N_6792,N_6702);
or U7815 (N_7815,N_6450,N_6714);
or U7816 (N_7816,N_6151,N_6193);
nor U7817 (N_7817,N_6164,N_6268);
nand U7818 (N_7818,N_6342,N_6781);
and U7819 (N_7819,N_6051,N_6505);
nor U7820 (N_7820,N_6571,N_6820);
nand U7821 (N_7821,N_6148,N_6428);
and U7822 (N_7822,N_6914,N_6481);
and U7823 (N_7823,N_6621,N_6181);
nor U7824 (N_7824,N_6764,N_6251);
nor U7825 (N_7825,N_6380,N_6786);
and U7826 (N_7826,N_6513,N_6224);
and U7827 (N_7827,N_6639,N_6418);
nor U7828 (N_7828,N_6828,N_6414);
or U7829 (N_7829,N_6128,N_6597);
and U7830 (N_7830,N_6412,N_6311);
or U7831 (N_7831,N_6124,N_6208);
xor U7832 (N_7832,N_6252,N_6808);
nor U7833 (N_7833,N_6480,N_6384);
or U7834 (N_7834,N_6934,N_6641);
xor U7835 (N_7835,N_6050,N_6914);
nor U7836 (N_7836,N_6412,N_6584);
and U7837 (N_7837,N_6625,N_6369);
and U7838 (N_7838,N_6366,N_6122);
and U7839 (N_7839,N_6006,N_6008);
and U7840 (N_7840,N_6715,N_6966);
and U7841 (N_7841,N_6976,N_6991);
or U7842 (N_7842,N_6529,N_6294);
nand U7843 (N_7843,N_6187,N_6784);
and U7844 (N_7844,N_6029,N_6971);
nand U7845 (N_7845,N_6252,N_6631);
or U7846 (N_7846,N_6473,N_6905);
xnor U7847 (N_7847,N_6849,N_6047);
nand U7848 (N_7848,N_6490,N_6053);
nor U7849 (N_7849,N_6446,N_6241);
and U7850 (N_7850,N_6578,N_6836);
xor U7851 (N_7851,N_6593,N_6368);
nor U7852 (N_7852,N_6769,N_6562);
or U7853 (N_7853,N_6271,N_6946);
xor U7854 (N_7854,N_6618,N_6832);
xnor U7855 (N_7855,N_6191,N_6852);
nor U7856 (N_7856,N_6541,N_6582);
xor U7857 (N_7857,N_6147,N_6112);
or U7858 (N_7858,N_6741,N_6577);
nand U7859 (N_7859,N_6770,N_6852);
or U7860 (N_7860,N_6112,N_6701);
xor U7861 (N_7861,N_6216,N_6804);
and U7862 (N_7862,N_6989,N_6860);
nor U7863 (N_7863,N_6653,N_6654);
or U7864 (N_7864,N_6794,N_6699);
nor U7865 (N_7865,N_6936,N_6832);
nand U7866 (N_7866,N_6228,N_6335);
xor U7867 (N_7867,N_6722,N_6067);
and U7868 (N_7868,N_6353,N_6712);
nand U7869 (N_7869,N_6417,N_6442);
nand U7870 (N_7870,N_6772,N_6024);
and U7871 (N_7871,N_6564,N_6075);
nor U7872 (N_7872,N_6854,N_6433);
nand U7873 (N_7873,N_6208,N_6739);
or U7874 (N_7874,N_6117,N_6284);
nor U7875 (N_7875,N_6398,N_6356);
nor U7876 (N_7876,N_6611,N_6641);
or U7877 (N_7877,N_6600,N_6704);
xnor U7878 (N_7878,N_6274,N_6495);
and U7879 (N_7879,N_6538,N_6675);
nand U7880 (N_7880,N_6552,N_6103);
nand U7881 (N_7881,N_6251,N_6117);
nand U7882 (N_7882,N_6399,N_6266);
nor U7883 (N_7883,N_6873,N_6716);
xnor U7884 (N_7884,N_6958,N_6488);
nand U7885 (N_7885,N_6578,N_6975);
nand U7886 (N_7886,N_6767,N_6938);
nor U7887 (N_7887,N_6618,N_6412);
and U7888 (N_7888,N_6707,N_6418);
or U7889 (N_7889,N_6266,N_6479);
or U7890 (N_7890,N_6676,N_6581);
and U7891 (N_7891,N_6683,N_6948);
nand U7892 (N_7892,N_6157,N_6014);
xor U7893 (N_7893,N_6284,N_6479);
and U7894 (N_7894,N_6380,N_6128);
nor U7895 (N_7895,N_6631,N_6054);
nand U7896 (N_7896,N_6286,N_6757);
nor U7897 (N_7897,N_6799,N_6466);
xor U7898 (N_7898,N_6843,N_6515);
and U7899 (N_7899,N_6989,N_6889);
or U7900 (N_7900,N_6839,N_6183);
nand U7901 (N_7901,N_6237,N_6836);
or U7902 (N_7902,N_6349,N_6264);
nand U7903 (N_7903,N_6785,N_6924);
nor U7904 (N_7904,N_6775,N_6260);
and U7905 (N_7905,N_6316,N_6015);
xnor U7906 (N_7906,N_6471,N_6628);
nand U7907 (N_7907,N_6039,N_6561);
and U7908 (N_7908,N_6310,N_6097);
and U7909 (N_7909,N_6951,N_6062);
and U7910 (N_7910,N_6158,N_6693);
xnor U7911 (N_7911,N_6723,N_6677);
nor U7912 (N_7912,N_6053,N_6319);
or U7913 (N_7913,N_6574,N_6223);
and U7914 (N_7914,N_6720,N_6733);
nand U7915 (N_7915,N_6185,N_6187);
xor U7916 (N_7916,N_6841,N_6946);
and U7917 (N_7917,N_6379,N_6708);
nand U7918 (N_7918,N_6200,N_6238);
or U7919 (N_7919,N_6919,N_6538);
nor U7920 (N_7920,N_6940,N_6005);
nor U7921 (N_7921,N_6014,N_6908);
and U7922 (N_7922,N_6685,N_6917);
nor U7923 (N_7923,N_6680,N_6214);
nand U7924 (N_7924,N_6223,N_6005);
and U7925 (N_7925,N_6510,N_6593);
or U7926 (N_7926,N_6811,N_6226);
or U7927 (N_7927,N_6435,N_6017);
and U7928 (N_7928,N_6791,N_6960);
and U7929 (N_7929,N_6416,N_6122);
and U7930 (N_7930,N_6356,N_6505);
and U7931 (N_7931,N_6330,N_6328);
and U7932 (N_7932,N_6486,N_6498);
nand U7933 (N_7933,N_6778,N_6491);
xnor U7934 (N_7934,N_6097,N_6205);
xnor U7935 (N_7935,N_6767,N_6961);
nor U7936 (N_7936,N_6689,N_6071);
or U7937 (N_7937,N_6913,N_6114);
or U7938 (N_7938,N_6473,N_6647);
and U7939 (N_7939,N_6548,N_6320);
nand U7940 (N_7940,N_6949,N_6282);
and U7941 (N_7941,N_6832,N_6722);
nand U7942 (N_7942,N_6987,N_6270);
and U7943 (N_7943,N_6504,N_6106);
or U7944 (N_7944,N_6533,N_6742);
or U7945 (N_7945,N_6275,N_6677);
nor U7946 (N_7946,N_6673,N_6248);
or U7947 (N_7947,N_6898,N_6644);
xnor U7948 (N_7948,N_6072,N_6733);
or U7949 (N_7949,N_6079,N_6487);
and U7950 (N_7950,N_6336,N_6844);
and U7951 (N_7951,N_6651,N_6711);
nand U7952 (N_7952,N_6048,N_6631);
nand U7953 (N_7953,N_6823,N_6071);
nor U7954 (N_7954,N_6253,N_6015);
nor U7955 (N_7955,N_6203,N_6202);
nor U7956 (N_7956,N_6454,N_6791);
and U7957 (N_7957,N_6903,N_6212);
nor U7958 (N_7958,N_6840,N_6801);
nand U7959 (N_7959,N_6474,N_6786);
xor U7960 (N_7960,N_6632,N_6696);
nand U7961 (N_7961,N_6228,N_6677);
nand U7962 (N_7962,N_6825,N_6071);
xor U7963 (N_7963,N_6800,N_6434);
and U7964 (N_7964,N_6293,N_6459);
or U7965 (N_7965,N_6096,N_6755);
nor U7966 (N_7966,N_6620,N_6134);
nor U7967 (N_7967,N_6515,N_6900);
or U7968 (N_7968,N_6463,N_6272);
and U7969 (N_7969,N_6819,N_6679);
and U7970 (N_7970,N_6317,N_6647);
nand U7971 (N_7971,N_6740,N_6829);
or U7972 (N_7972,N_6119,N_6326);
nand U7973 (N_7973,N_6077,N_6450);
or U7974 (N_7974,N_6403,N_6152);
nor U7975 (N_7975,N_6691,N_6562);
or U7976 (N_7976,N_6743,N_6851);
nand U7977 (N_7977,N_6379,N_6825);
and U7978 (N_7978,N_6265,N_6479);
or U7979 (N_7979,N_6988,N_6756);
and U7980 (N_7980,N_6053,N_6002);
nor U7981 (N_7981,N_6384,N_6881);
nand U7982 (N_7982,N_6421,N_6461);
nand U7983 (N_7983,N_6987,N_6505);
nand U7984 (N_7984,N_6943,N_6026);
nor U7985 (N_7985,N_6658,N_6423);
nand U7986 (N_7986,N_6574,N_6243);
nand U7987 (N_7987,N_6920,N_6516);
and U7988 (N_7988,N_6645,N_6014);
or U7989 (N_7989,N_6898,N_6866);
or U7990 (N_7990,N_6076,N_6025);
or U7991 (N_7991,N_6583,N_6035);
nand U7992 (N_7992,N_6557,N_6274);
and U7993 (N_7993,N_6215,N_6284);
xnor U7994 (N_7994,N_6720,N_6899);
or U7995 (N_7995,N_6609,N_6362);
nor U7996 (N_7996,N_6627,N_6200);
nor U7997 (N_7997,N_6209,N_6821);
or U7998 (N_7998,N_6738,N_6598);
or U7999 (N_7999,N_6278,N_6769);
or U8000 (N_8000,N_7501,N_7572);
nand U8001 (N_8001,N_7405,N_7265);
nand U8002 (N_8002,N_7578,N_7616);
nor U8003 (N_8003,N_7907,N_7036);
and U8004 (N_8004,N_7493,N_7612);
nor U8005 (N_8005,N_7762,N_7797);
or U8006 (N_8006,N_7415,N_7239);
or U8007 (N_8007,N_7842,N_7108);
nand U8008 (N_8008,N_7173,N_7002);
or U8009 (N_8009,N_7961,N_7628);
or U8010 (N_8010,N_7291,N_7970);
nor U8011 (N_8011,N_7644,N_7109);
and U8012 (N_8012,N_7465,N_7581);
and U8013 (N_8013,N_7323,N_7783);
nand U8014 (N_8014,N_7049,N_7969);
xnor U8015 (N_8015,N_7330,N_7182);
xnor U8016 (N_8016,N_7351,N_7694);
or U8017 (N_8017,N_7867,N_7993);
and U8018 (N_8018,N_7498,N_7152);
or U8019 (N_8019,N_7463,N_7116);
nor U8020 (N_8020,N_7489,N_7930);
nand U8021 (N_8021,N_7104,N_7278);
or U8022 (N_8022,N_7853,N_7926);
xor U8023 (N_8023,N_7507,N_7425);
or U8024 (N_8024,N_7600,N_7359);
or U8025 (N_8025,N_7187,N_7376);
nor U8026 (N_8026,N_7076,N_7032);
and U8027 (N_8027,N_7928,N_7657);
xnor U8028 (N_8028,N_7666,N_7039);
nor U8029 (N_8029,N_7114,N_7886);
nand U8030 (N_8030,N_7509,N_7846);
nand U8031 (N_8031,N_7322,N_7096);
and U8032 (N_8032,N_7219,N_7899);
xnor U8033 (N_8033,N_7448,N_7488);
or U8034 (N_8034,N_7284,N_7902);
nor U8035 (N_8035,N_7643,N_7472);
and U8036 (N_8036,N_7226,N_7776);
nor U8037 (N_8037,N_7453,N_7045);
nand U8038 (N_8038,N_7834,N_7151);
or U8039 (N_8039,N_7863,N_7872);
nor U8040 (N_8040,N_7954,N_7388);
nor U8041 (N_8041,N_7431,N_7378);
nor U8042 (N_8042,N_7306,N_7195);
or U8043 (N_8043,N_7174,N_7619);
and U8044 (N_8044,N_7720,N_7709);
nor U8045 (N_8045,N_7295,N_7972);
nor U8046 (N_8046,N_7528,N_7952);
and U8047 (N_8047,N_7656,N_7212);
xnor U8048 (N_8048,N_7981,N_7208);
xor U8049 (N_8049,N_7023,N_7156);
or U8050 (N_8050,N_7565,N_7125);
nor U8051 (N_8051,N_7971,N_7980);
nand U8052 (N_8052,N_7221,N_7826);
nor U8053 (N_8053,N_7966,N_7796);
xnor U8054 (N_8054,N_7582,N_7963);
nor U8055 (N_8055,N_7638,N_7369);
and U8056 (N_8056,N_7247,N_7682);
or U8057 (N_8057,N_7311,N_7426);
nor U8058 (N_8058,N_7160,N_7207);
and U8059 (N_8059,N_7874,N_7767);
and U8060 (N_8060,N_7601,N_7445);
and U8061 (N_8061,N_7135,N_7920);
or U8062 (N_8062,N_7040,N_7546);
nand U8063 (N_8063,N_7833,N_7234);
or U8064 (N_8064,N_7486,N_7804);
nand U8065 (N_8065,N_7761,N_7436);
nor U8066 (N_8066,N_7115,N_7811);
or U8067 (N_8067,N_7778,N_7715);
or U8068 (N_8068,N_7157,N_7771);
nand U8069 (N_8069,N_7932,N_7461);
or U8070 (N_8070,N_7175,N_7676);
xor U8071 (N_8071,N_7766,N_7785);
or U8072 (N_8072,N_7557,N_7944);
nand U8073 (N_8073,N_7809,N_7094);
nor U8074 (N_8074,N_7814,N_7051);
xnor U8075 (N_8075,N_7377,N_7285);
nand U8076 (N_8076,N_7007,N_7325);
and U8077 (N_8077,N_7894,N_7865);
nand U8078 (N_8078,N_7693,N_7646);
or U8079 (N_8079,N_7113,N_7434);
or U8080 (N_8080,N_7397,N_7086);
and U8081 (N_8081,N_7494,N_7988);
nor U8082 (N_8082,N_7244,N_7908);
or U8083 (N_8083,N_7667,N_7428);
nand U8084 (N_8084,N_7120,N_7898);
and U8085 (N_8085,N_7877,N_7091);
nand U8086 (N_8086,N_7592,N_7671);
or U8087 (N_8087,N_7340,N_7299);
nand U8088 (N_8088,N_7844,N_7320);
nand U8089 (N_8089,N_7913,N_7413);
and U8090 (N_8090,N_7469,N_7731);
xor U8091 (N_8091,N_7301,N_7257);
nor U8092 (N_8092,N_7589,N_7866);
and U8093 (N_8093,N_7089,N_7995);
xor U8094 (N_8094,N_7362,N_7895);
nor U8095 (N_8095,N_7951,N_7348);
nand U8096 (N_8096,N_7477,N_7610);
and U8097 (N_8097,N_7206,N_7645);
or U8098 (N_8098,N_7707,N_7310);
nor U8099 (N_8099,N_7381,N_7941);
xnor U8100 (N_8100,N_7637,N_7881);
or U8101 (N_8101,N_7407,N_7060);
nor U8102 (N_8102,N_7847,N_7746);
or U8103 (N_8103,N_7396,N_7129);
and U8104 (N_8104,N_7101,N_7551);
nand U8105 (N_8105,N_7389,N_7805);
and U8106 (N_8106,N_7550,N_7105);
and U8107 (N_8107,N_7634,N_7909);
nor U8108 (N_8108,N_7754,N_7631);
nor U8109 (N_8109,N_7673,N_7356);
or U8110 (N_8110,N_7836,N_7368);
nor U8111 (N_8111,N_7992,N_7680);
nor U8112 (N_8112,N_7700,N_7430);
nor U8113 (N_8113,N_7497,N_7364);
nand U8114 (N_8114,N_7548,N_7132);
xor U8115 (N_8115,N_7879,N_7912);
and U8116 (N_8116,N_7256,N_7942);
or U8117 (N_8117,N_7547,N_7033);
nand U8118 (N_8118,N_7190,N_7529);
or U8119 (N_8119,N_7292,N_7649);
and U8120 (N_8120,N_7177,N_7495);
and U8121 (N_8121,N_7655,N_7755);
and U8122 (N_8122,N_7417,N_7901);
xor U8123 (N_8123,N_7375,N_7537);
nor U8124 (N_8124,N_7579,N_7663);
and U8125 (N_8125,N_7499,N_7411);
nor U8126 (N_8126,N_7556,N_7987);
and U8127 (N_8127,N_7456,N_7274);
nand U8128 (N_8128,N_7354,N_7080);
or U8129 (N_8129,N_7316,N_7815);
nand U8130 (N_8130,N_7964,N_7337);
or U8131 (N_8131,N_7611,N_7245);
or U8132 (N_8132,N_7399,N_7530);
xnor U8133 (N_8133,N_7103,N_7324);
nor U8134 (N_8134,N_7722,N_7636);
nand U8135 (N_8135,N_7986,N_7522);
and U8136 (N_8136,N_7989,N_7480);
nor U8137 (N_8137,N_7946,N_7880);
or U8138 (N_8138,N_7701,N_7213);
or U8139 (N_8139,N_7353,N_7163);
xor U8140 (N_8140,N_7735,N_7542);
and U8141 (N_8141,N_7845,N_7384);
nor U8142 (N_8142,N_7838,N_7022);
or U8143 (N_8143,N_7167,N_7892);
and U8144 (N_8144,N_7552,N_7008);
and U8145 (N_8145,N_7059,N_7027);
and U8146 (N_8146,N_7905,N_7317);
nor U8147 (N_8147,N_7728,N_7669);
and U8148 (N_8148,N_7539,N_7736);
nor U8149 (N_8149,N_7540,N_7336);
and U8150 (N_8150,N_7147,N_7593);
and U8151 (N_8151,N_7651,N_7824);
and U8152 (N_8152,N_7272,N_7164);
nand U8153 (N_8153,N_7690,N_7191);
nand U8154 (N_8154,N_7297,N_7181);
nor U8155 (N_8155,N_7748,N_7615);
nand U8156 (N_8156,N_7617,N_7281);
nand U8157 (N_8157,N_7535,N_7686);
xnor U8158 (N_8158,N_7897,N_7000);
or U8159 (N_8159,N_7092,N_7596);
xor U8160 (N_8160,N_7883,N_7140);
nand U8161 (N_8161,N_7392,N_7314);
nand U8162 (N_8162,N_7126,N_7280);
nand U8163 (N_8163,N_7705,N_7440);
or U8164 (N_8164,N_7267,N_7119);
nand U8165 (N_8165,N_7774,N_7678);
nor U8166 (N_8166,N_7861,N_7420);
or U8167 (N_8167,N_7192,N_7800);
nand U8168 (N_8168,N_7222,N_7238);
nor U8169 (N_8169,N_7478,N_7878);
and U8170 (N_8170,N_7347,N_7924);
or U8171 (N_8171,N_7958,N_7575);
nor U8172 (N_8172,N_7211,N_7034);
nand U8173 (N_8173,N_7081,N_7464);
or U8174 (N_8174,N_7732,N_7597);
or U8175 (N_8175,N_7888,N_7217);
xnor U8176 (N_8176,N_7470,N_7335);
nor U8177 (N_8177,N_7777,N_7041);
and U8178 (N_8178,N_7711,N_7155);
and U8179 (N_8179,N_7672,N_7569);
nand U8180 (N_8180,N_7432,N_7231);
and U8181 (N_8181,N_7401,N_7520);
nand U8182 (N_8182,N_7885,N_7111);
and U8183 (N_8183,N_7982,N_7015);
nand U8184 (N_8184,N_7232,N_7973);
nor U8185 (N_8185,N_7810,N_7994);
and U8186 (N_8186,N_7409,N_7268);
nor U8187 (N_8187,N_7048,N_7717);
nand U8188 (N_8188,N_7275,N_7055);
nand U8189 (N_8189,N_7661,N_7840);
and U8190 (N_8190,N_7806,N_7654);
nor U8191 (N_8191,N_7756,N_7940);
and U8192 (N_8192,N_7228,N_7516);
and U8193 (N_8193,N_7817,N_7443);
or U8194 (N_8194,N_7254,N_7025);
xor U8195 (N_8195,N_7412,N_7985);
nand U8196 (N_8196,N_7090,N_7568);
nand U8197 (N_8197,N_7220,N_7248);
and U8198 (N_8198,N_7020,N_7884);
or U8199 (N_8199,N_7296,N_7553);
xnor U8200 (N_8200,N_7189,N_7227);
xor U8201 (N_8201,N_7503,N_7067);
and U8202 (N_8202,N_7283,N_7176);
or U8203 (N_8203,N_7276,N_7074);
xnor U8204 (N_8204,N_7702,N_7005);
and U8205 (N_8205,N_7492,N_7695);
xnor U8206 (N_8206,N_7851,N_7670);
nand U8207 (N_8207,N_7936,N_7962);
or U8208 (N_8208,N_7146,N_7757);
nand U8209 (N_8209,N_7483,N_7889);
nand U8210 (N_8210,N_7640,N_7893);
xnor U8211 (N_8211,N_7554,N_7279);
nand U8212 (N_8212,N_7361,N_7047);
nand U8213 (N_8213,N_7315,N_7689);
or U8214 (N_8214,N_7787,N_7763);
and U8215 (N_8215,N_7910,N_7142);
nand U8216 (N_8216,N_7410,N_7618);
and U8217 (N_8217,N_7143,N_7939);
nand U8218 (N_8218,N_7696,N_7016);
and U8219 (N_8219,N_7068,N_7466);
or U8220 (N_8220,N_7996,N_7960);
or U8221 (N_8221,N_7747,N_7035);
nand U8222 (N_8222,N_7014,N_7261);
or U8223 (N_8223,N_7843,N_7848);
nand U8224 (N_8224,N_7798,N_7538);
and U8225 (N_8225,N_7684,N_7950);
nor U8226 (N_8226,N_7215,N_7876);
nand U8227 (N_8227,N_7668,N_7243);
nand U8228 (N_8228,N_7590,N_7949);
nor U8229 (N_8229,N_7224,N_7468);
nor U8230 (N_8230,N_7527,N_7745);
or U8231 (N_8231,N_7482,N_7312);
nand U8232 (N_8232,N_7473,N_7009);
or U8233 (N_8233,N_7263,N_7740);
and U8234 (N_8234,N_7795,N_7319);
nand U8235 (N_8235,N_7052,N_7093);
or U8236 (N_8236,N_7769,N_7571);
nand U8237 (N_8237,N_7917,N_7737);
or U8238 (N_8238,N_7629,N_7003);
or U8239 (N_8239,N_7688,N_7246);
and U8240 (N_8240,N_7588,N_7402);
nor U8241 (N_8241,N_7698,N_7511);
or U8242 (N_8242,N_7161,N_7458);
and U8243 (N_8243,N_7484,N_7726);
nand U8244 (N_8244,N_7967,N_7760);
nand U8245 (N_8245,N_7948,N_7223);
nor U8246 (N_8246,N_7580,N_7945);
or U8247 (N_8247,N_7641,N_7828);
and U8248 (N_8248,N_7262,N_7692);
nand U8249 (N_8249,N_7270,N_7773);
and U8250 (N_8250,N_7998,N_7652);
nand U8251 (N_8251,N_7915,N_7414);
nor U8252 (N_8252,N_7438,N_7199);
or U8253 (N_8253,N_7435,N_7504);
xnor U8254 (N_8254,N_7380,N_7162);
and U8255 (N_8255,N_7321,N_7475);
nand U8256 (N_8256,N_7338,N_7070);
nand U8257 (N_8257,N_7869,N_7308);
and U8258 (N_8258,N_7991,N_7518);
or U8259 (N_8259,N_7400,N_7794);
nor U8260 (N_8260,N_7719,N_7044);
nand U8261 (N_8261,N_7429,N_7549);
nand U8262 (N_8262,N_7237,N_7046);
nand U8263 (N_8263,N_7632,N_7439);
and U8264 (N_8264,N_7563,N_7521);
or U8265 (N_8265,N_7896,N_7724);
and U8266 (N_8266,N_7976,N_7862);
xor U8267 (N_8267,N_7573,N_7449);
xor U8268 (N_8268,N_7054,N_7071);
and U8269 (N_8269,N_7753,N_7560);
or U8270 (N_8270,N_7534,N_7779);
or U8271 (N_8271,N_7789,N_7562);
or U8272 (N_8272,N_7128,N_7733);
nand U8273 (N_8273,N_7374,N_7857);
nor U8274 (N_8274,N_7710,N_7006);
or U8275 (N_8275,N_7259,N_7305);
or U8276 (N_8276,N_7555,N_7024);
or U8277 (N_8277,N_7699,N_7452);
nor U8278 (N_8278,N_7603,N_7558);
and U8279 (N_8279,N_7532,N_7122);
or U8280 (N_8280,N_7250,N_7937);
nor U8281 (N_8281,N_7180,N_7136);
nor U8282 (N_8282,N_7594,N_7765);
or U8283 (N_8283,N_7525,N_7772);
nor U8284 (N_8284,N_7997,N_7346);
or U8285 (N_8285,N_7209,N_7999);
and U8286 (N_8286,N_7660,N_7764);
or U8287 (N_8287,N_7864,N_7855);
nand U8288 (N_8288,N_7077,N_7916);
nand U8289 (N_8289,N_7607,N_7602);
xnor U8290 (N_8290,N_7391,N_7185);
and U8291 (N_8291,N_7138,N_7309);
or U8292 (N_8292,N_7169,N_7752);
nand U8293 (N_8293,N_7642,N_7481);
nor U8294 (N_8294,N_7729,N_7403);
and U8295 (N_8295,N_7471,N_7802);
nor U8296 (N_8296,N_7371,N_7255);
or U8297 (N_8297,N_7127,N_7433);
and U8298 (N_8298,N_7923,N_7240);
and U8299 (N_8299,N_7822,N_7703);
and U8300 (N_8300,N_7394,N_7541);
or U8301 (N_8301,N_7379,N_7825);
nand U8302 (N_8302,N_7069,N_7957);
nand U8303 (N_8303,N_7854,N_7447);
nand U8304 (N_8304,N_7821,N_7770);
nand U8305 (N_8305,N_7282,N_7056);
and U8306 (N_8306,N_7066,N_7358);
or U8307 (N_8307,N_7633,N_7918);
nand U8308 (N_8308,N_7955,N_7061);
nand U8309 (N_8309,N_7647,N_7137);
or U8310 (N_8310,N_7013,N_7965);
and U8311 (N_8311,N_7620,N_7029);
nand U8312 (N_8312,N_7734,N_7978);
or U8313 (N_8313,N_7406,N_7159);
xor U8314 (N_8314,N_7437,N_7210);
and U8315 (N_8315,N_7390,N_7216);
and U8316 (N_8316,N_7419,N_7591);
and U8317 (N_8317,N_7900,N_7459);
nand U8318 (N_8318,N_7627,N_7253);
and U8319 (N_8319,N_7201,N_7112);
nand U8320 (N_8320,N_7635,N_7318);
and U8321 (N_8321,N_7614,N_7574);
nor U8322 (N_8322,N_7808,N_7818);
xor U8323 (N_8323,N_7730,N_7031);
or U8324 (N_8324,N_7623,N_7704);
and U8325 (N_8325,N_7807,N_7084);
nor U8326 (N_8326,N_7107,N_7333);
nor U8327 (N_8327,N_7172,N_7057);
nand U8328 (N_8328,N_7085,N_7011);
and U8329 (N_8329,N_7837,N_7196);
nand U8330 (N_8330,N_7890,N_7373);
and U8331 (N_8331,N_7365,N_7968);
nand U8332 (N_8332,N_7799,N_7083);
xor U8333 (N_8333,N_7904,N_7801);
and U8334 (N_8334,N_7567,N_7868);
nand U8335 (N_8335,N_7313,N_7218);
nor U8336 (N_8336,N_7037,N_7050);
nor U8337 (N_8337,N_7441,N_7271);
or U8338 (N_8338,N_7630,N_7302);
or U8339 (N_8339,N_7708,N_7536);
nand U8340 (N_8340,N_7454,N_7508);
and U8341 (N_8341,N_7249,N_7653);
and U8342 (N_8342,N_7513,N_7519);
and U8343 (N_8343,N_7974,N_7154);
and U8344 (N_8344,N_7858,N_7131);
or U8345 (N_8345,N_7514,N_7713);
and U8346 (N_8346,N_7922,N_7398);
nand U8347 (N_8347,N_7307,N_7664);
nor U8348 (N_8348,N_7017,N_7533);
or U8349 (N_8349,N_7150,N_7018);
xor U8350 (N_8350,N_7831,N_7674);
nor U8351 (N_8351,N_7442,N_7485);
or U8352 (N_8352,N_7788,N_7675);
or U8353 (N_8353,N_7121,N_7194);
nor U8354 (N_8354,N_7576,N_7813);
nor U8355 (N_8355,N_7938,N_7933);
or U8356 (N_8356,N_7241,N_7658);
and U8357 (N_8357,N_7205,N_7339);
and U8358 (N_8358,N_7564,N_7827);
nand U8359 (N_8359,N_7184,N_7875);
nand U8360 (N_8360,N_7124,N_7683);
nand U8361 (N_8361,N_7178,N_7098);
or U8362 (N_8362,N_7500,N_7506);
nand U8363 (N_8363,N_7697,N_7123);
nand U8364 (N_8364,N_7515,N_7490);
nand U8365 (N_8365,N_7079,N_7739);
xnor U8366 (N_8366,N_7030,N_7832);
nor U8367 (N_8367,N_7395,N_7100);
or U8368 (N_8368,N_7749,N_7782);
nor U8369 (N_8369,N_7523,N_7286);
nand U8370 (N_8370,N_7956,N_7665);
or U8371 (N_8371,N_7983,N_7133);
nand U8372 (N_8372,N_7775,N_7784);
nor U8373 (N_8373,N_7058,N_7606);
nor U8374 (N_8374,N_7609,N_7106);
and U8375 (N_8375,N_7288,N_7839);
and U8376 (N_8376,N_7148,N_7570);
and U8377 (N_8377,N_7332,N_7608);
nand U8378 (N_8378,N_7510,N_7416);
or U8379 (N_8379,N_7063,N_7812);
nor U8380 (N_8380,N_7613,N_7345);
or U8381 (N_8381,N_7975,N_7427);
and U8382 (N_8382,N_7158,N_7650);
nor U8383 (N_8383,N_7360,N_7457);
and U8384 (N_8384,N_7648,N_7242);
and U8385 (N_8385,N_7010,N_7850);
nor U8386 (N_8386,N_7326,N_7873);
xor U8387 (N_8387,N_7743,N_7460);
nand U8388 (N_8388,N_7141,N_7450);
nand U8389 (N_8389,N_7871,N_7758);
nor U8390 (N_8390,N_7204,N_7544);
xnor U8391 (N_8391,N_7906,N_7977);
xnor U8392 (N_8392,N_7639,N_7605);
nand U8393 (N_8393,N_7197,N_7424);
nand U8394 (N_8394,N_7496,N_7543);
or U8395 (N_8395,N_7229,N_7294);
nand U8396 (N_8396,N_7153,N_7768);
nor U8397 (N_8397,N_7479,N_7200);
or U8398 (N_8398,N_7064,N_7203);
nand U8399 (N_8399,N_7383,N_7363);
and U8400 (N_8400,N_7681,N_7919);
nand U8401 (N_8401,N_7742,N_7677);
or U8402 (N_8402,N_7979,N_7598);
nor U8403 (N_8403,N_7266,N_7087);
or U8404 (N_8404,N_7943,N_7984);
nand U8405 (N_8405,N_7474,N_7595);
or U8406 (N_8406,N_7102,N_7342);
nand U8407 (N_8407,N_7531,N_7790);
nor U8408 (N_8408,N_7110,N_7097);
xnor U8409 (N_8409,N_7235,N_7685);
or U8410 (N_8410,N_7829,N_7366);
nor U8411 (N_8411,N_7935,N_7078);
nor U8412 (N_8412,N_7251,N_7451);
and U8413 (N_8413,N_7718,N_7830);
nand U8414 (N_8414,N_7387,N_7277);
xnor U8415 (N_8415,N_7082,N_7751);
and U8416 (N_8416,N_7852,N_7331);
xor U8417 (N_8417,N_7927,N_7487);
or U8418 (N_8418,N_7502,N_7233);
or U8419 (N_8419,N_7856,N_7870);
and U8420 (N_8420,N_7328,N_7264);
xnor U8421 (N_8421,N_7293,N_7491);
nand U8422 (N_8422,N_7462,N_7584);
and U8423 (N_8423,N_7791,N_7624);
xor U8424 (N_8424,N_7179,N_7021);
nand U8425 (N_8425,N_7372,N_7750);
nor U8426 (N_8426,N_7171,N_7139);
nand U8427 (N_8427,N_7088,N_7236);
nor U8428 (N_8428,N_7370,N_7914);
or U8429 (N_8429,N_7042,N_7382);
nor U8430 (N_8430,N_7599,N_7386);
nor U8431 (N_8431,N_7823,N_7170);
nor U8432 (N_8432,N_7467,N_7921);
and U8433 (N_8433,N_7408,N_7026);
nor U8434 (N_8434,N_7260,N_7099);
nand U8435 (N_8435,N_7476,N_7947);
nor U8436 (N_8436,N_7446,N_7214);
and U8437 (N_8437,N_7300,N_7625);
or U8438 (N_8438,N_7367,N_7357);
or U8439 (N_8439,N_7741,N_7849);
nand U8440 (N_8440,N_7355,N_7911);
or U8441 (N_8441,N_7759,N_7421);
xnor U8442 (N_8442,N_7118,N_7882);
and U8443 (N_8443,N_7891,N_7352);
or U8444 (N_8444,N_7166,N_7327);
xor U8445 (N_8445,N_7792,N_7714);
or U8446 (N_8446,N_7723,N_7038);
nand U8447 (N_8447,N_7577,N_7781);
or U8448 (N_8448,N_7202,N_7816);
or U8449 (N_8449,N_7290,N_7586);
nand U8450 (N_8450,N_7786,N_7903);
or U8451 (N_8451,N_7188,N_7225);
nand U8452 (N_8452,N_7193,N_7780);
and U8453 (N_8453,N_7258,N_7043);
xnor U8454 (N_8454,N_7925,N_7621);
or U8455 (N_8455,N_7350,N_7820);
and U8456 (N_8456,N_7727,N_7004);
nor U8457 (N_8457,N_7168,N_7418);
nor U8458 (N_8458,N_7343,N_7344);
and U8459 (N_8459,N_7404,N_7073);
and U8460 (N_8460,N_7422,N_7072);
and U8461 (N_8461,N_7329,N_7583);
nand U8462 (N_8462,N_7545,N_7298);
nor U8463 (N_8463,N_7725,N_7959);
xnor U8464 (N_8464,N_7183,N_7931);
and U8465 (N_8465,N_7444,N_7062);
or U8466 (N_8466,N_7393,N_7165);
nand U8467 (N_8467,N_7028,N_7887);
and U8468 (N_8468,N_7334,N_7385);
and U8469 (N_8469,N_7053,N_7001);
nor U8470 (N_8470,N_7585,N_7679);
and U8471 (N_8471,N_7145,N_7012);
nand U8472 (N_8472,N_7716,N_7198);
and U8473 (N_8473,N_7587,N_7144);
nand U8474 (N_8474,N_7341,N_7512);
and U8475 (N_8475,N_7721,N_7687);
nor U8476 (N_8476,N_7793,N_7075);
or U8477 (N_8477,N_7859,N_7691);
and U8478 (N_8478,N_7289,N_7738);
and U8479 (N_8479,N_7803,N_7134);
nand U8480 (N_8480,N_7524,N_7130);
nor U8481 (N_8481,N_7841,N_7304);
and U8482 (N_8482,N_7517,N_7953);
nand U8483 (N_8483,N_7819,N_7835);
nand U8484 (N_8484,N_7934,N_7626);
nor U8485 (N_8485,N_7526,N_7065);
and U8486 (N_8486,N_7561,N_7149);
nand U8487 (N_8487,N_7659,N_7303);
nor U8488 (N_8488,N_7423,N_7455);
nand U8489 (N_8489,N_7252,N_7505);
nand U8490 (N_8490,N_7604,N_7117);
and U8491 (N_8491,N_7662,N_7269);
and U8492 (N_8492,N_7230,N_7622);
or U8493 (N_8493,N_7712,N_7929);
nand U8494 (N_8494,N_7287,N_7990);
nor U8495 (N_8495,N_7349,N_7019);
nand U8496 (N_8496,N_7559,N_7706);
or U8497 (N_8497,N_7744,N_7273);
and U8498 (N_8498,N_7186,N_7095);
and U8499 (N_8499,N_7860,N_7566);
and U8500 (N_8500,N_7320,N_7222);
and U8501 (N_8501,N_7408,N_7205);
nor U8502 (N_8502,N_7165,N_7582);
nand U8503 (N_8503,N_7914,N_7725);
xnor U8504 (N_8504,N_7060,N_7096);
nor U8505 (N_8505,N_7921,N_7979);
nand U8506 (N_8506,N_7949,N_7859);
or U8507 (N_8507,N_7986,N_7453);
or U8508 (N_8508,N_7629,N_7758);
nand U8509 (N_8509,N_7220,N_7034);
xor U8510 (N_8510,N_7420,N_7606);
and U8511 (N_8511,N_7919,N_7761);
or U8512 (N_8512,N_7173,N_7577);
nand U8513 (N_8513,N_7598,N_7189);
and U8514 (N_8514,N_7584,N_7074);
nor U8515 (N_8515,N_7879,N_7347);
nand U8516 (N_8516,N_7239,N_7374);
or U8517 (N_8517,N_7743,N_7047);
or U8518 (N_8518,N_7041,N_7820);
and U8519 (N_8519,N_7164,N_7392);
nor U8520 (N_8520,N_7573,N_7015);
nand U8521 (N_8521,N_7443,N_7549);
nor U8522 (N_8522,N_7894,N_7313);
and U8523 (N_8523,N_7663,N_7931);
nor U8524 (N_8524,N_7891,N_7715);
nand U8525 (N_8525,N_7167,N_7855);
and U8526 (N_8526,N_7427,N_7521);
xnor U8527 (N_8527,N_7742,N_7029);
nand U8528 (N_8528,N_7609,N_7501);
and U8529 (N_8529,N_7872,N_7604);
nand U8530 (N_8530,N_7907,N_7712);
nand U8531 (N_8531,N_7948,N_7874);
xor U8532 (N_8532,N_7002,N_7784);
and U8533 (N_8533,N_7293,N_7489);
and U8534 (N_8534,N_7097,N_7042);
nor U8535 (N_8535,N_7294,N_7224);
nand U8536 (N_8536,N_7820,N_7518);
and U8537 (N_8537,N_7197,N_7614);
nor U8538 (N_8538,N_7286,N_7108);
nor U8539 (N_8539,N_7065,N_7974);
or U8540 (N_8540,N_7295,N_7118);
xor U8541 (N_8541,N_7924,N_7237);
or U8542 (N_8542,N_7532,N_7953);
nand U8543 (N_8543,N_7400,N_7931);
or U8544 (N_8544,N_7697,N_7863);
nand U8545 (N_8545,N_7924,N_7938);
nand U8546 (N_8546,N_7698,N_7598);
nor U8547 (N_8547,N_7061,N_7700);
or U8548 (N_8548,N_7712,N_7974);
nand U8549 (N_8549,N_7897,N_7190);
nor U8550 (N_8550,N_7019,N_7093);
or U8551 (N_8551,N_7242,N_7512);
nor U8552 (N_8552,N_7696,N_7046);
and U8553 (N_8553,N_7709,N_7520);
nand U8554 (N_8554,N_7285,N_7959);
nand U8555 (N_8555,N_7048,N_7927);
nor U8556 (N_8556,N_7135,N_7235);
and U8557 (N_8557,N_7966,N_7312);
or U8558 (N_8558,N_7324,N_7251);
nor U8559 (N_8559,N_7171,N_7643);
nand U8560 (N_8560,N_7175,N_7020);
nor U8561 (N_8561,N_7072,N_7310);
nand U8562 (N_8562,N_7412,N_7346);
and U8563 (N_8563,N_7697,N_7553);
nand U8564 (N_8564,N_7746,N_7491);
xor U8565 (N_8565,N_7603,N_7449);
nand U8566 (N_8566,N_7013,N_7029);
nor U8567 (N_8567,N_7820,N_7860);
or U8568 (N_8568,N_7067,N_7150);
nor U8569 (N_8569,N_7695,N_7227);
nor U8570 (N_8570,N_7171,N_7201);
and U8571 (N_8571,N_7028,N_7892);
nor U8572 (N_8572,N_7832,N_7178);
nor U8573 (N_8573,N_7740,N_7909);
and U8574 (N_8574,N_7910,N_7196);
or U8575 (N_8575,N_7268,N_7108);
or U8576 (N_8576,N_7808,N_7471);
or U8577 (N_8577,N_7194,N_7167);
nor U8578 (N_8578,N_7279,N_7367);
nand U8579 (N_8579,N_7014,N_7854);
nand U8580 (N_8580,N_7476,N_7314);
xnor U8581 (N_8581,N_7191,N_7460);
and U8582 (N_8582,N_7993,N_7494);
and U8583 (N_8583,N_7706,N_7471);
nand U8584 (N_8584,N_7023,N_7456);
and U8585 (N_8585,N_7905,N_7083);
or U8586 (N_8586,N_7996,N_7898);
xnor U8587 (N_8587,N_7539,N_7231);
and U8588 (N_8588,N_7320,N_7719);
or U8589 (N_8589,N_7167,N_7701);
and U8590 (N_8590,N_7378,N_7915);
or U8591 (N_8591,N_7033,N_7661);
xor U8592 (N_8592,N_7312,N_7575);
nor U8593 (N_8593,N_7842,N_7866);
nand U8594 (N_8594,N_7935,N_7949);
or U8595 (N_8595,N_7816,N_7219);
and U8596 (N_8596,N_7521,N_7879);
xor U8597 (N_8597,N_7110,N_7292);
nand U8598 (N_8598,N_7629,N_7080);
nor U8599 (N_8599,N_7599,N_7821);
or U8600 (N_8600,N_7444,N_7245);
nor U8601 (N_8601,N_7499,N_7678);
or U8602 (N_8602,N_7584,N_7716);
and U8603 (N_8603,N_7401,N_7307);
nand U8604 (N_8604,N_7969,N_7356);
or U8605 (N_8605,N_7409,N_7341);
and U8606 (N_8606,N_7709,N_7525);
nor U8607 (N_8607,N_7299,N_7078);
nor U8608 (N_8608,N_7726,N_7722);
nor U8609 (N_8609,N_7142,N_7421);
or U8610 (N_8610,N_7324,N_7963);
or U8611 (N_8611,N_7581,N_7745);
nor U8612 (N_8612,N_7287,N_7852);
and U8613 (N_8613,N_7620,N_7454);
nand U8614 (N_8614,N_7089,N_7937);
nand U8615 (N_8615,N_7484,N_7180);
and U8616 (N_8616,N_7137,N_7799);
nand U8617 (N_8617,N_7469,N_7255);
nand U8618 (N_8618,N_7554,N_7906);
or U8619 (N_8619,N_7881,N_7239);
xor U8620 (N_8620,N_7541,N_7084);
and U8621 (N_8621,N_7525,N_7902);
or U8622 (N_8622,N_7944,N_7284);
and U8623 (N_8623,N_7704,N_7908);
and U8624 (N_8624,N_7733,N_7915);
nand U8625 (N_8625,N_7433,N_7777);
nor U8626 (N_8626,N_7115,N_7688);
xor U8627 (N_8627,N_7443,N_7230);
and U8628 (N_8628,N_7384,N_7951);
nand U8629 (N_8629,N_7933,N_7481);
and U8630 (N_8630,N_7306,N_7347);
nor U8631 (N_8631,N_7180,N_7160);
xor U8632 (N_8632,N_7536,N_7635);
nand U8633 (N_8633,N_7243,N_7154);
nand U8634 (N_8634,N_7729,N_7389);
or U8635 (N_8635,N_7037,N_7063);
xor U8636 (N_8636,N_7929,N_7452);
nand U8637 (N_8637,N_7941,N_7915);
and U8638 (N_8638,N_7891,N_7349);
or U8639 (N_8639,N_7842,N_7445);
and U8640 (N_8640,N_7189,N_7115);
and U8641 (N_8641,N_7625,N_7669);
or U8642 (N_8642,N_7434,N_7732);
nor U8643 (N_8643,N_7597,N_7128);
or U8644 (N_8644,N_7710,N_7934);
xor U8645 (N_8645,N_7821,N_7501);
or U8646 (N_8646,N_7509,N_7099);
and U8647 (N_8647,N_7700,N_7706);
and U8648 (N_8648,N_7876,N_7289);
or U8649 (N_8649,N_7918,N_7192);
nand U8650 (N_8650,N_7902,N_7200);
xor U8651 (N_8651,N_7729,N_7073);
nand U8652 (N_8652,N_7539,N_7969);
nor U8653 (N_8653,N_7923,N_7039);
and U8654 (N_8654,N_7059,N_7369);
and U8655 (N_8655,N_7069,N_7732);
or U8656 (N_8656,N_7976,N_7469);
or U8657 (N_8657,N_7321,N_7173);
nand U8658 (N_8658,N_7566,N_7347);
and U8659 (N_8659,N_7508,N_7689);
or U8660 (N_8660,N_7189,N_7292);
nand U8661 (N_8661,N_7833,N_7105);
nand U8662 (N_8662,N_7407,N_7938);
xnor U8663 (N_8663,N_7068,N_7715);
nand U8664 (N_8664,N_7213,N_7054);
or U8665 (N_8665,N_7247,N_7787);
or U8666 (N_8666,N_7428,N_7088);
and U8667 (N_8667,N_7010,N_7393);
nand U8668 (N_8668,N_7476,N_7017);
and U8669 (N_8669,N_7198,N_7680);
and U8670 (N_8670,N_7878,N_7892);
nand U8671 (N_8671,N_7914,N_7633);
nor U8672 (N_8672,N_7548,N_7683);
nand U8673 (N_8673,N_7199,N_7231);
or U8674 (N_8674,N_7311,N_7559);
and U8675 (N_8675,N_7101,N_7387);
nor U8676 (N_8676,N_7418,N_7688);
nand U8677 (N_8677,N_7841,N_7621);
and U8678 (N_8678,N_7975,N_7080);
and U8679 (N_8679,N_7738,N_7118);
nand U8680 (N_8680,N_7206,N_7030);
or U8681 (N_8681,N_7829,N_7584);
or U8682 (N_8682,N_7166,N_7661);
nor U8683 (N_8683,N_7645,N_7067);
and U8684 (N_8684,N_7259,N_7127);
nand U8685 (N_8685,N_7102,N_7807);
nand U8686 (N_8686,N_7046,N_7531);
or U8687 (N_8687,N_7984,N_7353);
or U8688 (N_8688,N_7657,N_7893);
and U8689 (N_8689,N_7608,N_7627);
or U8690 (N_8690,N_7857,N_7881);
nand U8691 (N_8691,N_7867,N_7361);
or U8692 (N_8692,N_7141,N_7833);
nor U8693 (N_8693,N_7404,N_7716);
and U8694 (N_8694,N_7396,N_7764);
or U8695 (N_8695,N_7969,N_7293);
nand U8696 (N_8696,N_7875,N_7809);
nor U8697 (N_8697,N_7548,N_7202);
and U8698 (N_8698,N_7621,N_7940);
nor U8699 (N_8699,N_7614,N_7015);
or U8700 (N_8700,N_7928,N_7061);
and U8701 (N_8701,N_7814,N_7155);
nand U8702 (N_8702,N_7975,N_7139);
and U8703 (N_8703,N_7250,N_7598);
nor U8704 (N_8704,N_7685,N_7764);
nor U8705 (N_8705,N_7068,N_7873);
nor U8706 (N_8706,N_7781,N_7509);
nand U8707 (N_8707,N_7613,N_7644);
nor U8708 (N_8708,N_7458,N_7956);
nor U8709 (N_8709,N_7994,N_7655);
nand U8710 (N_8710,N_7959,N_7241);
and U8711 (N_8711,N_7889,N_7466);
or U8712 (N_8712,N_7529,N_7278);
xor U8713 (N_8713,N_7473,N_7157);
nand U8714 (N_8714,N_7864,N_7861);
nor U8715 (N_8715,N_7774,N_7569);
nand U8716 (N_8716,N_7533,N_7712);
or U8717 (N_8717,N_7448,N_7119);
nand U8718 (N_8718,N_7686,N_7586);
nand U8719 (N_8719,N_7800,N_7525);
nor U8720 (N_8720,N_7182,N_7589);
nor U8721 (N_8721,N_7380,N_7714);
and U8722 (N_8722,N_7615,N_7125);
or U8723 (N_8723,N_7635,N_7399);
nand U8724 (N_8724,N_7171,N_7157);
xor U8725 (N_8725,N_7988,N_7798);
or U8726 (N_8726,N_7290,N_7845);
nor U8727 (N_8727,N_7244,N_7710);
nor U8728 (N_8728,N_7127,N_7247);
or U8729 (N_8729,N_7289,N_7089);
or U8730 (N_8730,N_7416,N_7602);
and U8731 (N_8731,N_7326,N_7555);
or U8732 (N_8732,N_7861,N_7176);
nand U8733 (N_8733,N_7940,N_7368);
nor U8734 (N_8734,N_7365,N_7177);
or U8735 (N_8735,N_7237,N_7784);
or U8736 (N_8736,N_7758,N_7952);
nand U8737 (N_8737,N_7787,N_7760);
nor U8738 (N_8738,N_7737,N_7967);
and U8739 (N_8739,N_7842,N_7064);
nand U8740 (N_8740,N_7144,N_7343);
nor U8741 (N_8741,N_7397,N_7509);
nand U8742 (N_8742,N_7406,N_7668);
and U8743 (N_8743,N_7285,N_7791);
or U8744 (N_8744,N_7385,N_7619);
nand U8745 (N_8745,N_7739,N_7766);
nand U8746 (N_8746,N_7847,N_7237);
or U8747 (N_8747,N_7147,N_7026);
or U8748 (N_8748,N_7386,N_7526);
or U8749 (N_8749,N_7988,N_7451);
nand U8750 (N_8750,N_7805,N_7623);
nand U8751 (N_8751,N_7919,N_7467);
and U8752 (N_8752,N_7887,N_7675);
nor U8753 (N_8753,N_7533,N_7399);
nor U8754 (N_8754,N_7107,N_7385);
nor U8755 (N_8755,N_7473,N_7610);
and U8756 (N_8756,N_7858,N_7021);
nand U8757 (N_8757,N_7064,N_7004);
nor U8758 (N_8758,N_7893,N_7512);
nand U8759 (N_8759,N_7248,N_7686);
or U8760 (N_8760,N_7412,N_7549);
xnor U8761 (N_8761,N_7774,N_7358);
nand U8762 (N_8762,N_7160,N_7931);
nand U8763 (N_8763,N_7610,N_7341);
nor U8764 (N_8764,N_7732,N_7943);
or U8765 (N_8765,N_7081,N_7729);
nor U8766 (N_8766,N_7695,N_7238);
and U8767 (N_8767,N_7692,N_7718);
nand U8768 (N_8768,N_7708,N_7861);
or U8769 (N_8769,N_7890,N_7712);
nor U8770 (N_8770,N_7592,N_7019);
nor U8771 (N_8771,N_7316,N_7881);
nor U8772 (N_8772,N_7058,N_7125);
or U8773 (N_8773,N_7163,N_7830);
xor U8774 (N_8774,N_7843,N_7849);
nand U8775 (N_8775,N_7125,N_7966);
xnor U8776 (N_8776,N_7574,N_7398);
nor U8777 (N_8777,N_7606,N_7961);
or U8778 (N_8778,N_7515,N_7418);
nor U8779 (N_8779,N_7475,N_7451);
nand U8780 (N_8780,N_7197,N_7466);
and U8781 (N_8781,N_7669,N_7180);
nor U8782 (N_8782,N_7413,N_7154);
nand U8783 (N_8783,N_7181,N_7416);
nand U8784 (N_8784,N_7909,N_7669);
or U8785 (N_8785,N_7551,N_7784);
or U8786 (N_8786,N_7530,N_7101);
or U8787 (N_8787,N_7129,N_7829);
nor U8788 (N_8788,N_7160,N_7918);
or U8789 (N_8789,N_7168,N_7190);
or U8790 (N_8790,N_7202,N_7568);
or U8791 (N_8791,N_7320,N_7186);
or U8792 (N_8792,N_7287,N_7143);
nor U8793 (N_8793,N_7343,N_7538);
and U8794 (N_8794,N_7439,N_7455);
and U8795 (N_8795,N_7509,N_7862);
and U8796 (N_8796,N_7652,N_7655);
or U8797 (N_8797,N_7710,N_7301);
nand U8798 (N_8798,N_7724,N_7457);
and U8799 (N_8799,N_7676,N_7444);
or U8800 (N_8800,N_7555,N_7783);
nor U8801 (N_8801,N_7980,N_7801);
nand U8802 (N_8802,N_7915,N_7044);
nand U8803 (N_8803,N_7925,N_7480);
or U8804 (N_8804,N_7218,N_7837);
and U8805 (N_8805,N_7784,N_7408);
nor U8806 (N_8806,N_7224,N_7731);
and U8807 (N_8807,N_7020,N_7914);
nor U8808 (N_8808,N_7174,N_7956);
or U8809 (N_8809,N_7099,N_7586);
nand U8810 (N_8810,N_7183,N_7269);
nand U8811 (N_8811,N_7433,N_7864);
nor U8812 (N_8812,N_7840,N_7205);
nand U8813 (N_8813,N_7031,N_7708);
xor U8814 (N_8814,N_7043,N_7580);
or U8815 (N_8815,N_7317,N_7169);
nand U8816 (N_8816,N_7377,N_7761);
xnor U8817 (N_8817,N_7770,N_7798);
xnor U8818 (N_8818,N_7031,N_7369);
xnor U8819 (N_8819,N_7517,N_7403);
nor U8820 (N_8820,N_7799,N_7148);
or U8821 (N_8821,N_7129,N_7772);
nor U8822 (N_8822,N_7231,N_7436);
or U8823 (N_8823,N_7653,N_7161);
nand U8824 (N_8824,N_7433,N_7114);
nor U8825 (N_8825,N_7590,N_7730);
and U8826 (N_8826,N_7309,N_7273);
nand U8827 (N_8827,N_7227,N_7778);
and U8828 (N_8828,N_7859,N_7864);
nor U8829 (N_8829,N_7251,N_7156);
nor U8830 (N_8830,N_7935,N_7692);
nor U8831 (N_8831,N_7719,N_7643);
nor U8832 (N_8832,N_7763,N_7470);
xor U8833 (N_8833,N_7645,N_7798);
and U8834 (N_8834,N_7726,N_7760);
nand U8835 (N_8835,N_7540,N_7010);
nor U8836 (N_8836,N_7364,N_7088);
nor U8837 (N_8837,N_7375,N_7464);
nand U8838 (N_8838,N_7549,N_7189);
and U8839 (N_8839,N_7872,N_7722);
and U8840 (N_8840,N_7789,N_7509);
or U8841 (N_8841,N_7054,N_7801);
nand U8842 (N_8842,N_7188,N_7341);
xor U8843 (N_8843,N_7916,N_7430);
or U8844 (N_8844,N_7215,N_7684);
or U8845 (N_8845,N_7222,N_7686);
nand U8846 (N_8846,N_7672,N_7517);
and U8847 (N_8847,N_7087,N_7163);
nand U8848 (N_8848,N_7249,N_7713);
or U8849 (N_8849,N_7336,N_7564);
and U8850 (N_8850,N_7152,N_7077);
nand U8851 (N_8851,N_7469,N_7137);
nor U8852 (N_8852,N_7511,N_7798);
nor U8853 (N_8853,N_7456,N_7526);
xnor U8854 (N_8854,N_7803,N_7991);
nor U8855 (N_8855,N_7231,N_7412);
nand U8856 (N_8856,N_7534,N_7546);
or U8857 (N_8857,N_7127,N_7107);
xnor U8858 (N_8858,N_7753,N_7582);
or U8859 (N_8859,N_7314,N_7662);
and U8860 (N_8860,N_7209,N_7538);
nor U8861 (N_8861,N_7260,N_7496);
nor U8862 (N_8862,N_7558,N_7372);
nor U8863 (N_8863,N_7505,N_7488);
and U8864 (N_8864,N_7750,N_7667);
or U8865 (N_8865,N_7834,N_7156);
xor U8866 (N_8866,N_7669,N_7419);
nor U8867 (N_8867,N_7055,N_7063);
nand U8868 (N_8868,N_7668,N_7757);
nand U8869 (N_8869,N_7205,N_7995);
or U8870 (N_8870,N_7855,N_7327);
nor U8871 (N_8871,N_7410,N_7017);
nor U8872 (N_8872,N_7765,N_7863);
and U8873 (N_8873,N_7816,N_7140);
or U8874 (N_8874,N_7326,N_7695);
and U8875 (N_8875,N_7923,N_7626);
and U8876 (N_8876,N_7920,N_7137);
and U8877 (N_8877,N_7403,N_7544);
nand U8878 (N_8878,N_7265,N_7716);
or U8879 (N_8879,N_7027,N_7196);
or U8880 (N_8880,N_7829,N_7223);
and U8881 (N_8881,N_7207,N_7384);
xor U8882 (N_8882,N_7642,N_7944);
nand U8883 (N_8883,N_7970,N_7810);
xnor U8884 (N_8884,N_7991,N_7293);
or U8885 (N_8885,N_7050,N_7323);
nor U8886 (N_8886,N_7609,N_7834);
and U8887 (N_8887,N_7080,N_7369);
and U8888 (N_8888,N_7969,N_7823);
or U8889 (N_8889,N_7548,N_7920);
and U8890 (N_8890,N_7956,N_7115);
or U8891 (N_8891,N_7497,N_7347);
nor U8892 (N_8892,N_7572,N_7978);
or U8893 (N_8893,N_7959,N_7404);
or U8894 (N_8894,N_7986,N_7215);
xnor U8895 (N_8895,N_7156,N_7857);
or U8896 (N_8896,N_7239,N_7946);
and U8897 (N_8897,N_7610,N_7210);
and U8898 (N_8898,N_7312,N_7225);
nor U8899 (N_8899,N_7856,N_7599);
and U8900 (N_8900,N_7451,N_7690);
or U8901 (N_8901,N_7169,N_7281);
and U8902 (N_8902,N_7861,N_7513);
or U8903 (N_8903,N_7286,N_7359);
xor U8904 (N_8904,N_7801,N_7545);
nor U8905 (N_8905,N_7797,N_7272);
xor U8906 (N_8906,N_7982,N_7428);
xnor U8907 (N_8907,N_7235,N_7992);
nor U8908 (N_8908,N_7185,N_7863);
nor U8909 (N_8909,N_7326,N_7260);
xnor U8910 (N_8910,N_7097,N_7490);
nor U8911 (N_8911,N_7987,N_7533);
nand U8912 (N_8912,N_7237,N_7689);
nand U8913 (N_8913,N_7153,N_7749);
nand U8914 (N_8914,N_7624,N_7310);
and U8915 (N_8915,N_7439,N_7792);
nand U8916 (N_8916,N_7914,N_7695);
nand U8917 (N_8917,N_7315,N_7197);
nor U8918 (N_8918,N_7503,N_7226);
or U8919 (N_8919,N_7659,N_7614);
nand U8920 (N_8920,N_7603,N_7543);
nand U8921 (N_8921,N_7148,N_7713);
or U8922 (N_8922,N_7723,N_7176);
and U8923 (N_8923,N_7419,N_7655);
nand U8924 (N_8924,N_7624,N_7094);
and U8925 (N_8925,N_7502,N_7014);
and U8926 (N_8926,N_7871,N_7235);
nand U8927 (N_8927,N_7881,N_7591);
nor U8928 (N_8928,N_7836,N_7640);
nand U8929 (N_8929,N_7132,N_7251);
nor U8930 (N_8930,N_7112,N_7158);
nor U8931 (N_8931,N_7609,N_7290);
xnor U8932 (N_8932,N_7023,N_7932);
or U8933 (N_8933,N_7432,N_7991);
nand U8934 (N_8934,N_7052,N_7424);
and U8935 (N_8935,N_7954,N_7669);
nand U8936 (N_8936,N_7813,N_7785);
nor U8937 (N_8937,N_7343,N_7566);
and U8938 (N_8938,N_7885,N_7839);
xnor U8939 (N_8939,N_7212,N_7034);
nand U8940 (N_8940,N_7363,N_7650);
nand U8941 (N_8941,N_7202,N_7056);
or U8942 (N_8942,N_7967,N_7040);
nand U8943 (N_8943,N_7308,N_7566);
or U8944 (N_8944,N_7308,N_7137);
nand U8945 (N_8945,N_7097,N_7900);
nand U8946 (N_8946,N_7339,N_7449);
or U8947 (N_8947,N_7454,N_7496);
nor U8948 (N_8948,N_7446,N_7270);
or U8949 (N_8949,N_7720,N_7310);
or U8950 (N_8950,N_7389,N_7873);
and U8951 (N_8951,N_7952,N_7183);
nor U8952 (N_8952,N_7243,N_7475);
nand U8953 (N_8953,N_7940,N_7229);
nand U8954 (N_8954,N_7438,N_7054);
nor U8955 (N_8955,N_7693,N_7746);
or U8956 (N_8956,N_7970,N_7114);
xor U8957 (N_8957,N_7657,N_7089);
nor U8958 (N_8958,N_7643,N_7689);
nor U8959 (N_8959,N_7331,N_7231);
nand U8960 (N_8960,N_7289,N_7935);
nor U8961 (N_8961,N_7171,N_7471);
and U8962 (N_8962,N_7431,N_7317);
nand U8963 (N_8963,N_7565,N_7189);
or U8964 (N_8964,N_7845,N_7427);
nand U8965 (N_8965,N_7888,N_7914);
xor U8966 (N_8966,N_7961,N_7147);
or U8967 (N_8967,N_7590,N_7221);
xor U8968 (N_8968,N_7717,N_7441);
nand U8969 (N_8969,N_7221,N_7186);
nand U8970 (N_8970,N_7742,N_7353);
nand U8971 (N_8971,N_7613,N_7597);
or U8972 (N_8972,N_7891,N_7397);
nor U8973 (N_8973,N_7510,N_7924);
nor U8974 (N_8974,N_7676,N_7055);
nor U8975 (N_8975,N_7048,N_7611);
xnor U8976 (N_8976,N_7667,N_7107);
nand U8977 (N_8977,N_7061,N_7735);
nand U8978 (N_8978,N_7987,N_7527);
nor U8979 (N_8979,N_7957,N_7960);
or U8980 (N_8980,N_7936,N_7008);
and U8981 (N_8981,N_7406,N_7360);
nor U8982 (N_8982,N_7969,N_7847);
and U8983 (N_8983,N_7487,N_7723);
or U8984 (N_8984,N_7735,N_7643);
nand U8985 (N_8985,N_7744,N_7613);
nand U8986 (N_8986,N_7187,N_7028);
and U8987 (N_8987,N_7454,N_7686);
and U8988 (N_8988,N_7269,N_7723);
or U8989 (N_8989,N_7953,N_7429);
nor U8990 (N_8990,N_7189,N_7708);
nor U8991 (N_8991,N_7799,N_7200);
nand U8992 (N_8992,N_7961,N_7045);
nor U8993 (N_8993,N_7090,N_7057);
and U8994 (N_8994,N_7079,N_7188);
and U8995 (N_8995,N_7986,N_7323);
and U8996 (N_8996,N_7514,N_7138);
and U8997 (N_8997,N_7866,N_7840);
nand U8998 (N_8998,N_7967,N_7635);
or U8999 (N_8999,N_7947,N_7838);
nand U9000 (N_9000,N_8794,N_8922);
nor U9001 (N_9001,N_8321,N_8024);
and U9002 (N_9002,N_8222,N_8564);
or U9003 (N_9003,N_8701,N_8925);
nand U9004 (N_9004,N_8475,N_8692);
or U9005 (N_9005,N_8995,N_8967);
or U9006 (N_9006,N_8089,N_8803);
nor U9007 (N_9007,N_8631,N_8651);
and U9008 (N_9008,N_8713,N_8663);
or U9009 (N_9009,N_8776,N_8882);
nand U9010 (N_9010,N_8593,N_8239);
nand U9011 (N_9011,N_8290,N_8691);
or U9012 (N_9012,N_8318,N_8777);
or U9013 (N_9013,N_8848,N_8044);
and U9014 (N_9014,N_8204,N_8231);
nor U9015 (N_9015,N_8910,N_8994);
or U9016 (N_9016,N_8850,N_8530);
nand U9017 (N_9017,N_8829,N_8235);
nor U9018 (N_9018,N_8033,N_8953);
nor U9019 (N_9019,N_8924,N_8462);
nand U9020 (N_9020,N_8283,N_8774);
nor U9021 (N_9021,N_8048,N_8039);
xnor U9022 (N_9022,N_8810,N_8801);
xor U9023 (N_9023,N_8413,N_8862);
nor U9024 (N_9024,N_8589,N_8758);
and U9025 (N_9025,N_8330,N_8843);
nor U9026 (N_9026,N_8301,N_8468);
xnor U9027 (N_9027,N_8399,N_8835);
nor U9028 (N_9028,N_8073,N_8415);
nand U9029 (N_9029,N_8133,N_8920);
nand U9030 (N_9030,N_8090,N_8366);
nor U9031 (N_9031,N_8597,N_8212);
or U9032 (N_9032,N_8601,N_8488);
or U9033 (N_9033,N_8045,N_8122);
nor U9034 (N_9034,N_8097,N_8310);
nor U9035 (N_9035,N_8965,N_8229);
or U9036 (N_9036,N_8729,N_8359);
nor U9037 (N_9037,N_8508,N_8317);
nand U9038 (N_9038,N_8240,N_8904);
and U9039 (N_9039,N_8436,N_8827);
nor U9040 (N_9040,N_8215,N_8060);
nor U9041 (N_9041,N_8938,N_8258);
nor U9042 (N_9042,N_8677,N_8149);
xnor U9043 (N_9043,N_8199,N_8875);
or U9044 (N_9044,N_8216,N_8539);
xor U9045 (N_9045,N_8951,N_8182);
nor U9046 (N_9046,N_8770,N_8277);
nand U9047 (N_9047,N_8087,N_8251);
nor U9048 (N_9048,N_8689,N_8630);
xor U9049 (N_9049,N_8380,N_8489);
or U9050 (N_9050,N_8561,N_8647);
or U9051 (N_9051,N_8656,N_8595);
and U9052 (N_9052,N_8983,N_8858);
xor U9053 (N_9053,N_8932,N_8568);
nor U9054 (N_9054,N_8238,N_8752);
nor U9055 (N_9055,N_8658,N_8471);
nor U9056 (N_9056,N_8476,N_8790);
or U9057 (N_9057,N_8515,N_8009);
or U9058 (N_9058,N_8613,N_8887);
nand U9059 (N_9059,N_8678,N_8985);
nor U9060 (N_9060,N_8012,N_8406);
nor U9061 (N_9061,N_8464,N_8357);
nand U9062 (N_9062,N_8335,N_8859);
and U9063 (N_9063,N_8410,N_8679);
or U9064 (N_9064,N_8587,N_8351);
xor U9065 (N_9065,N_8531,N_8401);
or U9066 (N_9066,N_8662,N_8879);
nor U9067 (N_9067,N_8372,N_8798);
or U9068 (N_9068,N_8154,N_8778);
or U9069 (N_9069,N_8138,N_8062);
and U9070 (N_9070,N_8362,N_8896);
or U9071 (N_9071,N_8316,N_8292);
nor U9072 (N_9072,N_8522,N_8263);
or U9073 (N_9073,N_8479,N_8830);
and U9074 (N_9074,N_8693,N_8501);
nor U9075 (N_9075,N_8421,N_8017);
and U9076 (N_9076,N_8453,N_8035);
nand U9077 (N_9077,N_8695,N_8754);
or U9078 (N_9078,N_8140,N_8383);
nor U9079 (N_9079,N_8234,N_8818);
or U9080 (N_9080,N_8846,N_8120);
or U9081 (N_9081,N_8634,N_8387);
nand U9082 (N_9082,N_8513,N_8712);
nand U9083 (N_9083,N_8057,N_8353);
xnor U9084 (N_9084,N_8864,N_8937);
and U9085 (N_9085,N_8562,N_8586);
or U9086 (N_9086,N_8596,N_8000);
nand U9087 (N_9087,N_8825,N_8303);
and U9088 (N_9088,N_8096,N_8946);
nor U9089 (N_9089,N_8749,N_8168);
nor U9090 (N_9090,N_8757,N_8854);
xnor U9091 (N_9091,N_8111,N_8123);
and U9092 (N_9092,N_8177,N_8378);
or U9093 (N_9093,N_8502,N_8247);
nor U9094 (N_9094,N_8999,N_8124);
nand U9095 (N_9095,N_8414,N_8346);
and U9096 (N_9096,N_8931,N_8333);
and U9097 (N_9097,N_8645,N_8698);
or U9098 (N_9098,N_8541,N_8193);
xor U9099 (N_9099,N_8305,N_8127);
and U9100 (N_9100,N_8217,N_8973);
nor U9101 (N_9101,N_8425,N_8746);
or U9102 (N_9102,N_8671,N_8886);
and U9103 (N_9103,N_8724,N_8164);
nor U9104 (N_9104,N_8473,N_8437);
and U9105 (N_9105,N_8962,N_8440);
nor U9106 (N_9106,N_8288,N_8264);
nor U9107 (N_9107,N_8812,N_8328);
and U9108 (N_9108,N_8141,N_8960);
nor U9109 (N_9109,N_8675,N_8510);
nand U9110 (N_9110,N_8390,N_8573);
and U9111 (N_9111,N_8876,N_8025);
or U9112 (N_9112,N_8143,N_8914);
nor U9113 (N_9113,N_8386,N_8314);
nor U9114 (N_9114,N_8398,N_8908);
nand U9115 (N_9115,N_8132,N_8441);
and U9116 (N_9116,N_8418,N_8323);
or U9117 (N_9117,N_8061,N_8972);
or U9118 (N_9118,N_8772,N_8916);
and U9119 (N_9119,N_8736,N_8320);
nor U9120 (N_9120,N_8884,N_8889);
and U9121 (N_9121,N_8828,N_8431);
nor U9122 (N_9122,N_8881,N_8873);
nand U9123 (N_9123,N_8557,N_8579);
or U9124 (N_9124,N_8744,N_8104);
nor U9125 (N_9125,N_8709,N_8863);
nor U9126 (N_9126,N_8481,N_8241);
nand U9127 (N_9127,N_8661,N_8270);
or U9128 (N_9128,N_8535,N_8610);
or U9129 (N_9129,N_8350,N_8367);
nor U9130 (N_9130,N_8918,N_8052);
or U9131 (N_9131,N_8230,N_8358);
and U9132 (N_9132,N_8186,N_8957);
xnor U9133 (N_9133,N_8620,N_8851);
nand U9134 (N_9134,N_8200,N_8540);
or U9135 (N_9135,N_8393,N_8456);
or U9136 (N_9136,N_8871,N_8484);
xnor U9137 (N_9137,N_8706,N_8611);
and U9138 (N_9138,N_8625,N_8069);
nand U9139 (N_9139,N_8838,N_8542);
or U9140 (N_9140,N_8732,N_8548);
nand U9141 (N_9141,N_8948,N_8385);
nor U9142 (N_9142,N_8519,N_8092);
or U9143 (N_9143,N_8255,N_8796);
nand U9144 (N_9144,N_8298,N_8091);
nor U9145 (N_9145,N_8402,N_8767);
and U9146 (N_9146,N_8416,N_8114);
and U9147 (N_9147,N_8460,N_8486);
nor U9148 (N_9148,N_8849,N_8162);
nor U9149 (N_9149,N_8644,N_8322);
xnor U9150 (N_9150,N_8345,N_8629);
nand U9151 (N_9151,N_8733,N_8756);
and U9152 (N_9152,N_8616,N_8831);
or U9153 (N_9153,N_8979,N_8528);
or U9154 (N_9154,N_8341,N_8008);
nand U9155 (N_9155,N_8529,N_8660);
nand U9156 (N_9156,N_8071,N_8198);
nand U9157 (N_9157,N_8116,N_8265);
xor U9158 (N_9158,N_8655,N_8961);
and U9159 (N_9159,N_8452,N_8254);
or U9160 (N_9160,N_8536,N_8411);
nor U9161 (N_9161,N_8434,N_8930);
or U9162 (N_9162,N_8901,N_8727);
and U9163 (N_9163,N_8715,N_8594);
nand U9164 (N_9164,N_8259,N_8964);
xor U9165 (N_9165,N_8201,N_8694);
nor U9166 (N_9166,N_8424,N_8417);
xnor U9167 (N_9167,N_8093,N_8989);
nor U9168 (N_9168,N_8897,N_8438);
and U9169 (N_9169,N_8105,N_8667);
xnor U9170 (N_9170,N_8274,N_8505);
or U9171 (N_9171,N_8720,N_8252);
nor U9172 (N_9172,N_8731,N_8600);
and U9173 (N_9173,N_8928,N_8286);
or U9174 (N_9174,N_8276,N_8623);
nor U9175 (N_9175,N_8545,N_8684);
or U9176 (N_9176,N_8329,N_8364);
or U9177 (N_9177,N_8512,N_8294);
and U9178 (N_9178,N_8764,N_8100);
nand U9179 (N_9179,N_8567,N_8172);
and U9180 (N_9180,N_8996,N_8054);
or U9181 (N_9181,N_8449,N_8152);
nand U9182 (N_9182,N_8118,N_8950);
and U9183 (N_9183,N_8477,N_8907);
nand U9184 (N_9184,N_8407,N_8883);
and U9185 (N_9185,N_8181,N_8246);
and U9186 (N_9186,N_8993,N_8195);
or U9187 (N_9187,N_8253,N_8793);
or U9188 (N_9188,N_8942,N_8894);
nor U9189 (N_9189,N_8606,N_8430);
and U9190 (N_9190,N_8446,N_8670);
nand U9191 (N_9191,N_8779,N_8211);
or U9192 (N_9192,N_8547,N_8725);
and U9193 (N_9193,N_8668,N_8112);
nand U9194 (N_9194,N_8833,N_8377);
nor U9195 (N_9195,N_8046,N_8635);
or U9196 (N_9196,N_8454,N_8992);
nor U9197 (N_9197,N_8227,N_8943);
or U9198 (N_9198,N_8360,N_8011);
and U9199 (N_9199,N_8299,N_8409);
or U9200 (N_9200,N_8459,N_8248);
nor U9201 (N_9201,N_8839,N_8273);
and U9202 (N_9202,N_8337,N_8603);
and U9203 (N_9203,N_8743,N_8053);
nand U9204 (N_9204,N_8750,N_8503);
xnor U9205 (N_9205,N_8990,N_8837);
nor U9206 (N_9206,N_8748,N_8768);
and U9207 (N_9207,N_8817,N_8624);
nor U9208 (N_9208,N_8870,N_8432);
nand U9209 (N_9209,N_8309,N_8400);
and U9210 (N_9210,N_8082,N_8506);
nor U9211 (N_9211,N_8051,N_8444);
nor U9212 (N_9212,N_8860,N_8947);
or U9213 (N_9213,N_8982,N_8130);
xor U9214 (N_9214,N_8391,N_8065);
nor U9215 (N_9215,N_8042,N_8428);
nand U9216 (N_9216,N_8064,N_8147);
xor U9217 (N_9217,N_8912,N_8184);
and U9218 (N_9218,N_8565,N_8968);
nor U9219 (N_9219,N_8110,N_8218);
nand U9220 (N_9220,N_8180,N_8448);
nor U9221 (N_9221,N_8190,N_8232);
and U9222 (N_9222,N_8574,N_8716);
nor U9223 (N_9223,N_8028,N_8919);
xor U9224 (N_9224,N_8869,N_8971);
nor U9225 (N_9225,N_8394,N_8038);
nand U9226 (N_9226,N_8269,N_8178);
or U9227 (N_9227,N_8722,N_8219);
or U9228 (N_9228,N_8034,N_8702);
and U9229 (N_9229,N_8496,N_8699);
or U9230 (N_9230,N_8179,N_8555);
nand U9231 (N_9231,N_8155,N_8893);
and U9232 (N_9232,N_8639,N_8572);
nor U9233 (N_9233,N_8580,N_8319);
and U9234 (N_9234,N_8207,N_8049);
or U9235 (N_9235,N_8392,N_8643);
or U9236 (N_9236,N_8868,N_8905);
and U9237 (N_9237,N_8700,N_8681);
and U9238 (N_9238,N_8002,N_8030);
or U9239 (N_9239,N_8707,N_8537);
nand U9240 (N_9240,N_8084,N_8569);
xnor U9241 (N_9241,N_8435,N_8867);
or U9242 (N_9242,N_8786,N_8344);
xnor U9243 (N_9243,N_8811,N_8591);
or U9244 (N_9244,N_8202,N_8783);
and U9245 (N_9245,N_8327,N_8945);
or U9246 (N_9246,N_8369,N_8036);
nor U9247 (N_9247,N_8673,N_8244);
nor U9248 (N_9248,N_8281,N_8293);
or U9249 (N_9249,N_8497,N_8741);
xnor U9250 (N_9250,N_8792,N_8003);
nor U9251 (N_9251,N_8214,N_8261);
xor U9252 (N_9252,N_8526,N_8885);
nand U9253 (N_9253,N_8495,N_8368);
nor U9254 (N_9254,N_8855,N_8823);
nor U9255 (N_9255,N_8721,N_8389);
nor U9256 (N_9256,N_8083,N_8153);
and U9257 (N_9257,N_8952,N_8010);
xnor U9258 (N_9258,N_8142,N_8760);
nand U9259 (N_9259,N_8395,N_8755);
nor U9260 (N_9260,N_8081,N_8223);
and U9261 (N_9261,N_8483,N_8331);
xnor U9262 (N_9262,N_8272,N_8534);
xnor U9263 (N_9263,N_8791,N_8680);
or U9264 (N_9264,N_8816,N_8742);
and U9265 (N_9265,N_8005,N_8516);
nand U9266 (N_9266,N_8077,N_8278);
or U9267 (N_9267,N_8189,N_8987);
nor U9268 (N_9268,N_8326,N_8325);
and U9269 (N_9269,N_8955,N_8730);
or U9270 (N_9270,N_8514,N_8095);
nor U9271 (N_9271,N_8878,N_8847);
or U9272 (N_9272,N_8422,N_8094);
nor U9273 (N_9273,N_8146,N_8307);
nand U9274 (N_9274,N_8923,N_8031);
nand U9275 (N_9275,N_8852,N_8191);
nand U9276 (N_9276,N_8139,N_8205);
and U9277 (N_9277,N_8279,N_8027);
nand U9278 (N_9278,N_8233,N_8880);
xnor U9279 (N_9279,N_8004,N_8020);
or U9280 (N_9280,N_8121,N_8221);
nor U9281 (N_9281,N_8072,N_8311);
nor U9282 (N_9282,N_8160,N_8935);
nand U9283 (N_9283,N_8324,N_8958);
and U9284 (N_9284,N_8704,N_8926);
nand U9285 (N_9285,N_8384,N_8349);
and U9286 (N_9286,N_8210,N_8174);
nor U9287 (N_9287,N_8058,N_8915);
nand U9288 (N_9288,N_8976,N_8717);
nor U9289 (N_9289,N_8666,N_8078);
or U9290 (N_9290,N_8490,N_8352);
and U9291 (N_9291,N_8936,N_8066);
or U9292 (N_9292,N_8396,N_8397);
and U9293 (N_9293,N_8738,N_8841);
nand U9294 (N_9294,N_8379,N_8795);
and U9295 (N_9295,N_8762,N_8780);
and U9296 (N_9296,N_8621,N_8373);
nor U9297 (N_9297,N_8861,N_8682);
xor U9298 (N_9298,N_8605,N_8740);
and U9299 (N_9299,N_8457,N_8461);
nor U9300 (N_9300,N_8023,N_8509);
and U9301 (N_9301,N_8988,N_8518);
nor U9302 (N_9302,N_8819,N_8649);
and U9303 (N_9303,N_8636,N_8726);
or U9304 (N_9304,N_8775,N_8899);
and U9305 (N_9305,N_8225,N_8041);
nor U9306 (N_9306,N_8998,N_8617);
and U9307 (N_9307,N_8271,N_8131);
and U9308 (N_9308,N_8055,N_8267);
nand U9309 (N_9309,N_8109,N_8037);
nor U9310 (N_9310,N_8332,N_8342);
and U9311 (N_9311,N_8719,N_8170);
nand U9312 (N_9312,N_8429,N_8315);
or U9313 (N_9313,N_8642,N_8525);
or U9314 (N_9314,N_8013,N_8161);
nand U9315 (N_9315,N_8898,N_8646);
nand U9316 (N_9316,N_8063,N_8659);
or U9317 (N_9317,N_8275,N_8708);
and U9318 (N_9318,N_8059,N_8627);
xnor U9319 (N_9319,N_8821,N_8494);
nor U9320 (N_9320,N_8807,N_8842);
and U9321 (N_9321,N_8256,N_8280);
and U9322 (N_9322,N_8888,N_8136);
nand U9323 (N_9323,N_8085,N_8697);
and U9324 (N_9324,N_8633,N_8511);
xor U9325 (N_9325,N_8466,N_8356);
and U9326 (N_9326,N_8365,N_8618);
or U9327 (N_9327,N_8577,N_8169);
nand U9328 (N_9328,N_8439,N_8137);
and U9329 (N_9329,N_8236,N_8799);
and U9330 (N_9330,N_8944,N_8759);
or U9331 (N_9331,N_8284,N_8266);
or U9332 (N_9332,N_8813,N_8304);
nand U9333 (N_9333,N_8463,N_8785);
nor U9334 (N_9334,N_8688,N_8374);
nand U9335 (N_9335,N_8674,N_8187);
and U9336 (N_9336,N_8451,N_8076);
xnor U9337 (N_9337,N_8237,N_8956);
and U9338 (N_9338,N_8080,N_8480);
xor U9339 (N_9339,N_8206,N_8844);
or U9340 (N_9340,N_8302,N_8891);
or U9341 (N_9341,N_8075,N_8086);
nor U9342 (N_9342,N_8376,N_8019);
nand U9343 (N_9343,N_8523,N_8067);
or U9344 (N_9344,N_8134,N_8683);
nor U9345 (N_9345,N_8581,N_8228);
or U9346 (N_9346,N_8194,N_8203);
nand U9347 (N_9347,N_8933,N_8619);
nor U9348 (N_9348,N_8576,N_8363);
nand U9349 (N_9349,N_8427,N_8705);
nor U9350 (N_9350,N_8737,N_8442);
nand U9351 (N_9351,N_8500,N_8544);
and U9352 (N_9352,N_8157,N_8125);
nand U9353 (N_9353,N_8895,N_8289);
nor U9354 (N_9354,N_8312,N_8099);
nand U9355 (N_9355,N_8917,N_8609);
or U9356 (N_9356,N_8723,N_8443);
nor U9357 (N_9357,N_8485,N_8308);
nand U9358 (N_9358,N_8563,N_8626);
and U9359 (N_9359,N_8602,N_8478);
or U9360 (N_9360,N_8354,N_8450);
nand U9361 (N_9361,N_8690,N_8467);
nand U9362 (N_9362,N_8001,N_8213);
and U9363 (N_9363,N_8614,N_8188);
or U9364 (N_9364,N_8787,N_8173);
or U9365 (N_9365,N_8107,N_8804);
and U9366 (N_9366,N_8499,N_8527);
xor U9367 (N_9367,N_8520,N_8521);
or U9368 (N_9368,N_8102,N_8966);
nor U9369 (N_9369,N_8026,N_8834);
or U9370 (N_9370,N_8382,N_8734);
nor U9371 (N_9371,N_8208,N_8159);
nand U9372 (N_9372,N_8487,N_8648);
or U9373 (N_9373,N_8445,N_8088);
nand U9374 (N_9374,N_8672,N_8313);
nand U9375 (N_9375,N_8113,N_8021);
or U9376 (N_9376,N_8814,N_8117);
nor U9377 (N_9377,N_8771,N_8650);
and U9378 (N_9378,N_8652,N_8306);
nor U9379 (N_9379,N_8970,N_8297);
nand U9380 (N_9380,N_8608,N_8242);
or U9381 (N_9381,N_8664,N_8653);
xnor U9382 (N_9382,N_8669,N_8615);
nand U9383 (N_9383,N_8420,N_8538);
and U9384 (N_9384,N_8781,N_8815);
nand U9385 (N_9385,N_8158,N_8582);
nor U9386 (N_9386,N_8032,N_8892);
and U9387 (N_9387,N_8981,N_8176);
or U9388 (N_9388,N_8151,N_8939);
and U9389 (N_9389,N_8543,N_8654);
and U9390 (N_9390,N_8043,N_8739);
or U9391 (N_9391,N_8556,N_8447);
and U9392 (N_9392,N_8296,N_8334);
and U9393 (N_9393,N_8552,N_8590);
xor U9394 (N_9394,N_8108,N_8056);
nand U9395 (N_9395,N_8832,N_8098);
or U9396 (N_9396,N_8566,N_8282);
nor U9397 (N_9397,N_8361,N_8977);
xnor U9398 (N_9398,N_8978,N_8533);
and U9399 (N_9399,N_8984,N_8578);
and U9400 (N_9400,N_8163,N_8622);
nand U9401 (N_9401,N_8766,N_8986);
or U9402 (N_9402,N_8607,N_8913);
nand U9403 (N_9403,N_8560,N_8115);
or U9404 (N_9404,N_8765,N_8347);
or U9405 (N_9405,N_8103,N_8865);
or U9406 (N_9406,N_8802,N_8465);
nand U9407 (N_9407,N_8997,N_8941);
or U9408 (N_9408,N_8262,N_8974);
xnor U9409 (N_9409,N_8388,N_8047);
nor U9410 (N_9410,N_8339,N_8549);
nor U9411 (N_9411,N_8903,N_8735);
or U9412 (N_9412,N_8183,N_8638);
xnor U9413 (N_9413,N_8632,N_8800);
and U9414 (N_9414,N_8185,N_8482);
or U9415 (N_9415,N_8890,N_8822);
or U9416 (N_9416,N_8135,N_8074);
or U9417 (N_9417,N_8469,N_8806);
and U9418 (N_9418,N_8797,N_8585);
nand U9419 (N_9419,N_8007,N_8954);
and U9420 (N_9420,N_8474,N_8599);
and U9421 (N_9421,N_8584,N_8657);
nand U9422 (N_9422,N_8050,N_8840);
xnor U9423 (N_9423,N_8665,N_8551);
or U9424 (N_9424,N_8458,N_8745);
nor U9425 (N_9425,N_8826,N_8145);
nor U9426 (N_9426,N_8921,N_8929);
or U9427 (N_9427,N_8343,N_8604);
or U9428 (N_9428,N_8433,N_8524);
or U9429 (N_9429,N_8166,N_8773);
nor U9430 (N_9430,N_8018,N_8370);
nor U9431 (N_9431,N_8403,N_8348);
and U9432 (N_9432,N_8196,N_8686);
and U9433 (N_9433,N_8676,N_8789);
or U9434 (N_9434,N_8969,N_8249);
and U9435 (N_9435,N_8703,N_8751);
xnor U9436 (N_9436,N_8836,N_8769);
or U9437 (N_9437,N_8148,N_8150);
or U9438 (N_9438,N_8761,N_8507);
nor U9439 (N_9439,N_8492,N_8220);
nor U9440 (N_9440,N_8014,N_8763);
or U9441 (N_9441,N_8612,N_8546);
nor U9442 (N_9442,N_8029,N_8696);
or U9443 (N_9443,N_8845,N_8728);
nand U9444 (N_9444,N_8070,N_8902);
nor U9445 (N_9445,N_8588,N_8250);
and U9446 (N_9446,N_8245,N_8872);
xnor U9447 (N_9447,N_8820,N_8338);
nand U9448 (N_9448,N_8171,N_8711);
nor U9449 (N_9449,N_8909,N_8853);
nand U9450 (N_9450,N_8144,N_8975);
or U9451 (N_9451,N_8718,N_8423);
nand U9452 (N_9452,N_8295,N_8558);
or U9453 (N_9453,N_8300,N_8857);
and U9454 (N_9454,N_8934,N_8226);
and U9455 (N_9455,N_8106,N_8980);
and U9456 (N_9456,N_8570,N_8470);
or U9457 (N_9457,N_8687,N_8371);
and U9458 (N_9458,N_8156,N_8128);
or U9459 (N_9459,N_8498,N_8165);
or U9460 (N_9460,N_8016,N_8167);
nand U9461 (N_9461,N_8068,N_8532);
and U9462 (N_9462,N_8553,N_8710);
or U9463 (N_9463,N_8405,N_8554);
nand U9464 (N_9464,N_8243,N_8285);
and U9465 (N_9465,N_8598,N_8963);
and U9466 (N_9466,N_8808,N_8504);
or U9467 (N_9467,N_8375,N_8784);
nand U9468 (N_9468,N_8455,N_8788);
or U9469 (N_9469,N_8355,N_8906);
nand U9470 (N_9470,N_8753,N_8824);
nor U9471 (N_9471,N_8640,N_8419);
or U9472 (N_9472,N_8404,N_8129);
nor U9473 (N_9473,N_8022,N_8927);
xor U9474 (N_9474,N_8583,N_8412);
or U9475 (N_9475,N_8224,N_8101);
nor U9476 (N_9476,N_8805,N_8197);
and U9477 (N_9477,N_8381,N_8336);
nand U9478 (N_9478,N_8192,N_8015);
or U9479 (N_9479,N_8268,N_8714);
or U9480 (N_9480,N_8991,N_8571);
xnor U9481 (N_9481,N_8940,N_8291);
or U9482 (N_9482,N_8517,N_8900);
or U9483 (N_9483,N_8628,N_8408);
nand U9484 (N_9484,N_8126,N_8856);
nand U9485 (N_9485,N_8866,N_8877);
or U9486 (N_9486,N_8175,N_8959);
xnor U9487 (N_9487,N_8685,N_8209);
nand U9488 (N_9488,N_8911,N_8006);
or U9489 (N_9489,N_8637,N_8257);
nor U9490 (N_9490,N_8809,N_8874);
nor U9491 (N_9491,N_8472,N_8287);
and U9492 (N_9492,N_8426,N_8592);
nand U9493 (N_9493,N_8559,N_8340);
xor U9494 (N_9494,N_8493,N_8550);
or U9495 (N_9495,N_8491,N_8747);
xor U9496 (N_9496,N_8949,N_8260);
xor U9497 (N_9497,N_8641,N_8079);
nand U9498 (N_9498,N_8040,N_8575);
or U9499 (N_9499,N_8119,N_8782);
nor U9500 (N_9500,N_8967,N_8477);
nor U9501 (N_9501,N_8557,N_8559);
nand U9502 (N_9502,N_8938,N_8862);
or U9503 (N_9503,N_8595,N_8435);
nand U9504 (N_9504,N_8312,N_8739);
and U9505 (N_9505,N_8188,N_8007);
nand U9506 (N_9506,N_8103,N_8734);
nand U9507 (N_9507,N_8096,N_8065);
nand U9508 (N_9508,N_8054,N_8108);
or U9509 (N_9509,N_8483,N_8419);
nand U9510 (N_9510,N_8609,N_8437);
nand U9511 (N_9511,N_8911,N_8917);
or U9512 (N_9512,N_8650,N_8428);
or U9513 (N_9513,N_8409,N_8574);
and U9514 (N_9514,N_8586,N_8227);
and U9515 (N_9515,N_8246,N_8042);
xor U9516 (N_9516,N_8875,N_8333);
nor U9517 (N_9517,N_8745,N_8675);
nor U9518 (N_9518,N_8995,N_8673);
nor U9519 (N_9519,N_8326,N_8453);
or U9520 (N_9520,N_8960,N_8029);
nor U9521 (N_9521,N_8860,N_8532);
nand U9522 (N_9522,N_8454,N_8013);
or U9523 (N_9523,N_8828,N_8091);
or U9524 (N_9524,N_8518,N_8571);
nand U9525 (N_9525,N_8555,N_8561);
and U9526 (N_9526,N_8744,N_8202);
and U9527 (N_9527,N_8657,N_8049);
nor U9528 (N_9528,N_8969,N_8893);
nor U9529 (N_9529,N_8050,N_8519);
xor U9530 (N_9530,N_8724,N_8818);
and U9531 (N_9531,N_8986,N_8949);
nand U9532 (N_9532,N_8055,N_8725);
nor U9533 (N_9533,N_8610,N_8064);
and U9534 (N_9534,N_8468,N_8127);
nor U9535 (N_9535,N_8750,N_8891);
nand U9536 (N_9536,N_8194,N_8510);
nand U9537 (N_9537,N_8793,N_8260);
nor U9538 (N_9538,N_8136,N_8023);
and U9539 (N_9539,N_8882,N_8913);
and U9540 (N_9540,N_8866,N_8172);
nand U9541 (N_9541,N_8678,N_8247);
or U9542 (N_9542,N_8206,N_8833);
or U9543 (N_9543,N_8242,N_8805);
xnor U9544 (N_9544,N_8487,N_8314);
nand U9545 (N_9545,N_8527,N_8619);
nor U9546 (N_9546,N_8259,N_8023);
and U9547 (N_9547,N_8412,N_8707);
nor U9548 (N_9548,N_8237,N_8733);
nor U9549 (N_9549,N_8761,N_8571);
or U9550 (N_9550,N_8354,N_8444);
and U9551 (N_9551,N_8914,N_8464);
or U9552 (N_9552,N_8641,N_8500);
nor U9553 (N_9553,N_8764,N_8120);
xnor U9554 (N_9554,N_8177,N_8922);
and U9555 (N_9555,N_8441,N_8262);
and U9556 (N_9556,N_8096,N_8730);
or U9557 (N_9557,N_8613,N_8963);
nor U9558 (N_9558,N_8492,N_8674);
nor U9559 (N_9559,N_8713,N_8507);
or U9560 (N_9560,N_8747,N_8711);
nand U9561 (N_9561,N_8860,N_8309);
and U9562 (N_9562,N_8278,N_8485);
or U9563 (N_9563,N_8633,N_8037);
and U9564 (N_9564,N_8492,N_8993);
or U9565 (N_9565,N_8889,N_8584);
and U9566 (N_9566,N_8911,N_8794);
and U9567 (N_9567,N_8208,N_8317);
nand U9568 (N_9568,N_8607,N_8071);
xnor U9569 (N_9569,N_8867,N_8146);
nand U9570 (N_9570,N_8810,N_8736);
xnor U9571 (N_9571,N_8706,N_8413);
and U9572 (N_9572,N_8576,N_8795);
nor U9573 (N_9573,N_8935,N_8022);
nor U9574 (N_9574,N_8373,N_8832);
or U9575 (N_9575,N_8653,N_8457);
xnor U9576 (N_9576,N_8078,N_8084);
nor U9577 (N_9577,N_8557,N_8734);
and U9578 (N_9578,N_8834,N_8361);
xnor U9579 (N_9579,N_8092,N_8666);
and U9580 (N_9580,N_8840,N_8857);
nor U9581 (N_9581,N_8176,N_8811);
nand U9582 (N_9582,N_8089,N_8054);
and U9583 (N_9583,N_8504,N_8520);
or U9584 (N_9584,N_8053,N_8932);
nand U9585 (N_9585,N_8662,N_8458);
xor U9586 (N_9586,N_8180,N_8745);
and U9587 (N_9587,N_8187,N_8314);
nand U9588 (N_9588,N_8366,N_8385);
xor U9589 (N_9589,N_8054,N_8656);
nand U9590 (N_9590,N_8404,N_8604);
or U9591 (N_9591,N_8463,N_8670);
xnor U9592 (N_9592,N_8575,N_8951);
nand U9593 (N_9593,N_8049,N_8103);
or U9594 (N_9594,N_8185,N_8993);
nor U9595 (N_9595,N_8117,N_8312);
or U9596 (N_9596,N_8647,N_8431);
nor U9597 (N_9597,N_8693,N_8377);
and U9598 (N_9598,N_8394,N_8455);
nor U9599 (N_9599,N_8627,N_8713);
nor U9600 (N_9600,N_8718,N_8567);
or U9601 (N_9601,N_8264,N_8777);
and U9602 (N_9602,N_8866,N_8966);
or U9603 (N_9603,N_8603,N_8755);
and U9604 (N_9604,N_8603,N_8079);
nor U9605 (N_9605,N_8400,N_8766);
and U9606 (N_9606,N_8151,N_8631);
and U9607 (N_9607,N_8664,N_8270);
or U9608 (N_9608,N_8674,N_8981);
nor U9609 (N_9609,N_8642,N_8437);
or U9610 (N_9610,N_8327,N_8932);
nand U9611 (N_9611,N_8008,N_8970);
nor U9612 (N_9612,N_8097,N_8970);
nor U9613 (N_9613,N_8648,N_8969);
and U9614 (N_9614,N_8249,N_8640);
nor U9615 (N_9615,N_8610,N_8301);
nor U9616 (N_9616,N_8652,N_8799);
or U9617 (N_9617,N_8351,N_8311);
nor U9618 (N_9618,N_8362,N_8516);
or U9619 (N_9619,N_8531,N_8758);
nand U9620 (N_9620,N_8168,N_8080);
nor U9621 (N_9621,N_8255,N_8423);
xnor U9622 (N_9622,N_8287,N_8493);
nand U9623 (N_9623,N_8467,N_8381);
and U9624 (N_9624,N_8053,N_8313);
nand U9625 (N_9625,N_8087,N_8505);
and U9626 (N_9626,N_8638,N_8433);
and U9627 (N_9627,N_8757,N_8737);
or U9628 (N_9628,N_8216,N_8088);
nand U9629 (N_9629,N_8791,N_8483);
or U9630 (N_9630,N_8210,N_8937);
and U9631 (N_9631,N_8573,N_8629);
xnor U9632 (N_9632,N_8540,N_8206);
nand U9633 (N_9633,N_8675,N_8917);
nor U9634 (N_9634,N_8909,N_8824);
and U9635 (N_9635,N_8571,N_8365);
and U9636 (N_9636,N_8881,N_8353);
nand U9637 (N_9637,N_8943,N_8877);
xnor U9638 (N_9638,N_8846,N_8203);
nand U9639 (N_9639,N_8822,N_8194);
nand U9640 (N_9640,N_8107,N_8270);
nand U9641 (N_9641,N_8677,N_8463);
or U9642 (N_9642,N_8544,N_8042);
nand U9643 (N_9643,N_8461,N_8234);
and U9644 (N_9644,N_8045,N_8829);
or U9645 (N_9645,N_8248,N_8278);
nand U9646 (N_9646,N_8801,N_8742);
nand U9647 (N_9647,N_8913,N_8856);
nand U9648 (N_9648,N_8692,N_8456);
nand U9649 (N_9649,N_8260,N_8927);
or U9650 (N_9650,N_8846,N_8319);
nand U9651 (N_9651,N_8033,N_8505);
and U9652 (N_9652,N_8892,N_8445);
nand U9653 (N_9653,N_8610,N_8459);
and U9654 (N_9654,N_8371,N_8349);
nor U9655 (N_9655,N_8734,N_8866);
and U9656 (N_9656,N_8495,N_8581);
nor U9657 (N_9657,N_8263,N_8737);
or U9658 (N_9658,N_8294,N_8255);
nand U9659 (N_9659,N_8762,N_8246);
xnor U9660 (N_9660,N_8162,N_8750);
nand U9661 (N_9661,N_8721,N_8168);
xor U9662 (N_9662,N_8040,N_8955);
nand U9663 (N_9663,N_8927,N_8328);
xor U9664 (N_9664,N_8302,N_8335);
and U9665 (N_9665,N_8458,N_8259);
nor U9666 (N_9666,N_8467,N_8669);
or U9667 (N_9667,N_8371,N_8341);
nor U9668 (N_9668,N_8257,N_8830);
nand U9669 (N_9669,N_8408,N_8480);
nand U9670 (N_9670,N_8436,N_8663);
and U9671 (N_9671,N_8272,N_8425);
and U9672 (N_9672,N_8065,N_8668);
or U9673 (N_9673,N_8792,N_8250);
nor U9674 (N_9674,N_8303,N_8405);
and U9675 (N_9675,N_8719,N_8890);
nor U9676 (N_9676,N_8533,N_8332);
or U9677 (N_9677,N_8578,N_8468);
nand U9678 (N_9678,N_8182,N_8982);
or U9679 (N_9679,N_8628,N_8751);
or U9680 (N_9680,N_8817,N_8421);
and U9681 (N_9681,N_8405,N_8922);
and U9682 (N_9682,N_8832,N_8717);
nand U9683 (N_9683,N_8205,N_8871);
nor U9684 (N_9684,N_8965,N_8850);
nand U9685 (N_9685,N_8678,N_8750);
and U9686 (N_9686,N_8151,N_8805);
or U9687 (N_9687,N_8782,N_8509);
and U9688 (N_9688,N_8706,N_8079);
or U9689 (N_9689,N_8026,N_8547);
nor U9690 (N_9690,N_8057,N_8584);
or U9691 (N_9691,N_8000,N_8359);
nand U9692 (N_9692,N_8442,N_8201);
nand U9693 (N_9693,N_8080,N_8695);
or U9694 (N_9694,N_8043,N_8310);
or U9695 (N_9695,N_8956,N_8172);
and U9696 (N_9696,N_8914,N_8736);
nand U9697 (N_9697,N_8939,N_8041);
and U9698 (N_9698,N_8175,N_8431);
or U9699 (N_9699,N_8587,N_8052);
and U9700 (N_9700,N_8992,N_8392);
and U9701 (N_9701,N_8948,N_8101);
nand U9702 (N_9702,N_8076,N_8436);
or U9703 (N_9703,N_8898,N_8738);
or U9704 (N_9704,N_8272,N_8945);
and U9705 (N_9705,N_8133,N_8294);
nor U9706 (N_9706,N_8642,N_8728);
and U9707 (N_9707,N_8577,N_8440);
and U9708 (N_9708,N_8239,N_8443);
nand U9709 (N_9709,N_8021,N_8203);
nor U9710 (N_9710,N_8271,N_8290);
or U9711 (N_9711,N_8589,N_8940);
nand U9712 (N_9712,N_8282,N_8778);
and U9713 (N_9713,N_8102,N_8155);
nand U9714 (N_9714,N_8935,N_8903);
or U9715 (N_9715,N_8160,N_8025);
or U9716 (N_9716,N_8475,N_8081);
nor U9717 (N_9717,N_8898,N_8394);
nand U9718 (N_9718,N_8693,N_8987);
nand U9719 (N_9719,N_8832,N_8495);
and U9720 (N_9720,N_8479,N_8837);
or U9721 (N_9721,N_8323,N_8082);
nor U9722 (N_9722,N_8275,N_8257);
or U9723 (N_9723,N_8943,N_8349);
nand U9724 (N_9724,N_8487,N_8501);
and U9725 (N_9725,N_8532,N_8614);
nand U9726 (N_9726,N_8425,N_8183);
nor U9727 (N_9727,N_8459,N_8206);
nor U9728 (N_9728,N_8339,N_8699);
or U9729 (N_9729,N_8697,N_8806);
or U9730 (N_9730,N_8529,N_8217);
xor U9731 (N_9731,N_8047,N_8097);
nor U9732 (N_9732,N_8405,N_8178);
nand U9733 (N_9733,N_8258,N_8914);
or U9734 (N_9734,N_8811,N_8253);
nor U9735 (N_9735,N_8628,N_8339);
nor U9736 (N_9736,N_8067,N_8101);
nand U9737 (N_9737,N_8520,N_8975);
nand U9738 (N_9738,N_8914,N_8627);
or U9739 (N_9739,N_8015,N_8752);
nor U9740 (N_9740,N_8550,N_8337);
nand U9741 (N_9741,N_8126,N_8397);
and U9742 (N_9742,N_8096,N_8568);
and U9743 (N_9743,N_8153,N_8324);
xor U9744 (N_9744,N_8264,N_8138);
nand U9745 (N_9745,N_8783,N_8678);
nand U9746 (N_9746,N_8556,N_8830);
xor U9747 (N_9747,N_8987,N_8279);
nand U9748 (N_9748,N_8943,N_8625);
nor U9749 (N_9749,N_8150,N_8024);
or U9750 (N_9750,N_8298,N_8435);
and U9751 (N_9751,N_8827,N_8525);
and U9752 (N_9752,N_8084,N_8440);
or U9753 (N_9753,N_8619,N_8988);
or U9754 (N_9754,N_8691,N_8991);
or U9755 (N_9755,N_8706,N_8682);
or U9756 (N_9756,N_8906,N_8758);
or U9757 (N_9757,N_8097,N_8857);
and U9758 (N_9758,N_8862,N_8837);
and U9759 (N_9759,N_8079,N_8271);
nor U9760 (N_9760,N_8181,N_8862);
nor U9761 (N_9761,N_8424,N_8034);
or U9762 (N_9762,N_8329,N_8523);
nor U9763 (N_9763,N_8296,N_8752);
nor U9764 (N_9764,N_8626,N_8121);
and U9765 (N_9765,N_8301,N_8281);
and U9766 (N_9766,N_8770,N_8493);
nor U9767 (N_9767,N_8749,N_8720);
nor U9768 (N_9768,N_8365,N_8075);
nor U9769 (N_9769,N_8747,N_8901);
and U9770 (N_9770,N_8275,N_8562);
and U9771 (N_9771,N_8338,N_8020);
nor U9772 (N_9772,N_8755,N_8830);
or U9773 (N_9773,N_8835,N_8396);
or U9774 (N_9774,N_8088,N_8403);
and U9775 (N_9775,N_8282,N_8919);
and U9776 (N_9776,N_8663,N_8324);
and U9777 (N_9777,N_8276,N_8041);
nand U9778 (N_9778,N_8567,N_8975);
nor U9779 (N_9779,N_8763,N_8806);
or U9780 (N_9780,N_8594,N_8259);
nand U9781 (N_9781,N_8614,N_8601);
and U9782 (N_9782,N_8491,N_8574);
nor U9783 (N_9783,N_8133,N_8233);
and U9784 (N_9784,N_8819,N_8231);
and U9785 (N_9785,N_8730,N_8712);
and U9786 (N_9786,N_8422,N_8315);
nand U9787 (N_9787,N_8758,N_8108);
nor U9788 (N_9788,N_8891,N_8728);
nand U9789 (N_9789,N_8058,N_8381);
xor U9790 (N_9790,N_8430,N_8053);
or U9791 (N_9791,N_8043,N_8166);
nor U9792 (N_9792,N_8610,N_8181);
and U9793 (N_9793,N_8522,N_8205);
xnor U9794 (N_9794,N_8833,N_8909);
or U9795 (N_9795,N_8748,N_8782);
or U9796 (N_9796,N_8785,N_8301);
and U9797 (N_9797,N_8930,N_8482);
nand U9798 (N_9798,N_8753,N_8261);
xnor U9799 (N_9799,N_8819,N_8378);
xor U9800 (N_9800,N_8541,N_8415);
and U9801 (N_9801,N_8825,N_8302);
nor U9802 (N_9802,N_8019,N_8168);
or U9803 (N_9803,N_8820,N_8168);
nand U9804 (N_9804,N_8963,N_8214);
nor U9805 (N_9805,N_8447,N_8658);
and U9806 (N_9806,N_8749,N_8754);
xor U9807 (N_9807,N_8185,N_8724);
nand U9808 (N_9808,N_8632,N_8520);
or U9809 (N_9809,N_8431,N_8630);
and U9810 (N_9810,N_8428,N_8987);
nor U9811 (N_9811,N_8086,N_8995);
nor U9812 (N_9812,N_8967,N_8607);
nor U9813 (N_9813,N_8800,N_8833);
nor U9814 (N_9814,N_8809,N_8097);
nor U9815 (N_9815,N_8326,N_8850);
nand U9816 (N_9816,N_8757,N_8985);
nand U9817 (N_9817,N_8123,N_8649);
nand U9818 (N_9818,N_8083,N_8470);
and U9819 (N_9819,N_8136,N_8054);
nor U9820 (N_9820,N_8013,N_8284);
nor U9821 (N_9821,N_8088,N_8454);
nor U9822 (N_9822,N_8976,N_8467);
nand U9823 (N_9823,N_8143,N_8810);
nor U9824 (N_9824,N_8078,N_8873);
and U9825 (N_9825,N_8810,N_8350);
xnor U9826 (N_9826,N_8895,N_8492);
nor U9827 (N_9827,N_8064,N_8877);
nor U9828 (N_9828,N_8515,N_8441);
nor U9829 (N_9829,N_8413,N_8318);
and U9830 (N_9830,N_8141,N_8208);
nor U9831 (N_9831,N_8724,N_8548);
nor U9832 (N_9832,N_8487,N_8444);
and U9833 (N_9833,N_8575,N_8327);
and U9834 (N_9834,N_8860,N_8976);
and U9835 (N_9835,N_8777,N_8349);
or U9836 (N_9836,N_8477,N_8264);
nor U9837 (N_9837,N_8413,N_8068);
nand U9838 (N_9838,N_8232,N_8856);
nor U9839 (N_9839,N_8787,N_8432);
nor U9840 (N_9840,N_8601,N_8042);
nand U9841 (N_9841,N_8097,N_8627);
or U9842 (N_9842,N_8730,N_8888);
nor U9843 (N_9843,N_8639,N_8014);
or U9844 (N_9844,N_8246,N_8740);
xnor U9845 (N_9845,N_8737,N_8101);
nand U9846 (N_9846,N_8023,N_8002);
and U9847 (N_9847,N_8167,N_8477);
and U9848 (N_9848,N_8332,N_8359);
nor U9849 (N_9849,N_8829,N_8726);
or U9850 (N_9850,N_8484,N_8284);
nand U9851 (N_9851,N_8784,N_8585);
nor U9852 (N_9852,N_8200,N_8775);
nor U9853 (N_9853,N_8436,N_8928);
or U9854 (N_9854,N_8708,N_8462);
and U9855 (N_9855,N_8006,N_8461);
and U9856 (N_9856,N_8163,N_8802);
and U9857 (N_9857,N_8419,N_8804);
nand U9858 (N_9858,N_8035,N_8438);
nand U9859 (N_9859,N_8988,N_8732);
nor U9860 (N_9860,N_8589,N_8522);
and U9861 (N_9861,N_8420,N_8914);
and U9862 (N_9862,N_8809,N_8055);
nor U9863 (N_9863,N_8297,N_8177);
nand U9864 (N_9864,N_8646,N_8693);
or U9865 (N_9865,N_8259,N_8410);
and U9866 (N_9866,N_8816,N_8374);
and U9867 (N_9867,N_8528,N_8017);
nand U9868 (N_9868,N_8472,N_8869);
nand U9869 (N_9869,N_8815,N_8647);
or U9870 (N_9870,N_8135,N_8904);
nor U9871 (N_9871,N_8245,N_8932);
or U9872 (N_9872,N_8597,N_8203);
or U9873 (N_9873,N_8168,N_8445);
nand U9874 (N_9874,N_8464,N_8698);
nor U9875 (N_9875,N_8806,N_8917);
nand U9876 (N_9876,N_8991,N_8169);
or U9877 (N_9877,N_8079,N_8366);
nor U9878 (N_9878,N_8627,N_8244);
xor U9879 (N_9879,N_8536,N_8190);
or U9880 (N_9880,N_8081,N_8875);
or U9881 (N_9881,N_8922,N_8426);
and U9882 (N_9882,N_8462,N_8714);
xor U9883 (N_9883,N_8591,N_8395);
or U9884 (N_9884,N_8888,N_8015);
nand U9885 (N_9885,N_8385,N_8625);
or U9886 (N_9886,N_8995,N_8444);
nand U9887 (N_9887,N_8508,N_8935);
nor U9888 (N_9888,N_8940,N_8093);
or U9889 (N_9889,N_8211,N_8429);
nor U9890 (N_9890,N_8235,N_8131);
nor U9891 (N_9891,N_8991,N_8558);
nor U9892 (N_9892,N_8945,N_8439);
nand U9893 (N_9893,N_8122,N_8549);
and U9894 (N_9894,N_8685,N_8007);
and U9895 (N_9895,N_8650,N_8781);
and U9896 (N_9896,N_8907,N_8414);
xor U9897 (N_9897,N_8823,N_8665);
nand U9898 (N_9898,N_8880,N_8303);
xor U9899 (N_9899,N_8259,N_8821);
nand U9900 (N_9900,N_8557,N_8452);
xnor U9901 (N_9901,N_8660,N_8650);
nand U9902 (N_9902,N_8086,N_8958);
nand U9903 (N_9903,N_8699,N_8175);
xor U9904 (N_9904,N_8693,N_8101);
and U9905 (N_9905,N_8747,N_8118);
and U9906 (N_9906,N_8015,N_8560);
nand U9907 (N_9907,N_8274,N_8036);
xnor U9908 (N_9908,N_8897,N_8068);
and U9909 (N_9909,N_8564,N_8454);
nor U9910 (N_9910,N_8681,N_8414);
nand U9911 (N_9911,N_8953,N_8511);
nor U9912 (N_9912,N_8796,N_8939);
nor U9913 (N_9913,N_8126,N_8223);
or U9914 (N_9914,N_8901,N_8663);
and U9915 (N_9915,N_8491,N_8611);
nand U9916 (N_9916,N_8004,N_8985);
nor U9917 (N_9917,N_8552,N_8521);
and U9918 (N_9918,N_8748,N_8952);
or U9919 (N_9919,N_8291,N_8506);
and U9920 (N_9920,N_8506,N_8081);
or U9921 (N_9921,N_8272,N_8305);
nand U9922 (N_9922,N_8518,N_8909);
or U9923 (N_9923,N_8642,N_8636);
and U9924 (N_9924,N_8083,N_8779);
or U9925 (N_9925,N_8961,N_8857);
xor U9926 (N_9926,N_8292,N_8280);
or U9927 (N_9927,N_8248,N_8112);
and U9928 (N_9928,N_8086,N_8601);
nor U9929 (N_9929,N_8742,N_8154);
nand U9930 (N_9930,N_8589,N_8224);
nand U9931 (N_9931,N_8574,N_8015);
nor U9932 (N_9932,N_8709,N_8549);
nor U9933 (N_9933,N_8930,N_8555);
xnor U9934 (N_9934,N_8564,N_8367);
nor U9935 (N_9935,N_8329,N_8607);
and U9936 (N_9936,N_8593,N_8030);
and U9937 (N_9937,N_8930,N_8074);
nor U9938 (N_9938,N_8779,N_8100);
and U9939 (N_9939,N_8462,N_8272);
and U9940 (N_9940,N_8493,N_8039);
and U9941 (N_9941,N_8685,N_8982);
nor U9942 (N_9942,N_8737,N_8594);
and U9943 (N_9943,N_8788,N_8507);
nand U9944 (N_9944,N_8071,N_8323);
and U9945 (N_9945,N_8379,N_8744);
xnor U9946 (N_9946,N_8202,N_8829);
nand U9947 (N_9947,N_8788,N_8756);
xor U9948 (N_9948,N_8201,N_8655);
and U9949 (N_9949,N_8870,N_8836);
and U9950 (N_9950,N_8776,N_8402);
nand U9951 (N_9951,N_8569,N_8711);
nor U9952 (N_9952,N_8662,N_8369);
or U9953 (N_9953,N_8137,N_8482);
nand U9954 (N_9954,N_8041,N_8391);
nor U9955 (N_9955,N_8452,N_8732);
and U9956 (N_9956,N_8539,N_8339);
and U9957 (N_9957,N_8100,N_8810);
nand U9958 (N_9958,N_8924,N_8191);
nor U9959 (N_9959,N_8810,N_8897);
nand U9960 (N_9960,N_8841,N_8960);
xnor U9961 (N_9961,N_8377,N_8047);
and U9962 (N_9962,N_8925,N_8426);
xnor U9963 (N_9963,N_8902,N_8588);
and U9964 (N_9964,N_8939,N_8181);
nand U9965 (N_9965,N_8139,N_8500);
nand U9966 (N_9966,N_8859,N_8645);
nor U9967 (N_9967,N_8140,N_8438);
or U9968 (N_9968,N_8806,N_8171);
nand U9969 (N_9969,N_8094,N_8263);
nor U9970 (N_9970,N_8543,N_8948);
or U9971 (N_9971,N_8459,N_8061);
and U9972 (N_9972,N_8497,N_8577);
or U9973 (N_9973,N_8236,N_8879);
or U9974 (N_9974,N_8628,N_8671);
and U9975 (N_9975,N_8360,N_8931);
and U9976 (N_9976,N_8753,N_8692);
nor U9977 (N_9977,N_8027,N_8642);
nand U9978 (N_9978,N_8576,N_8134);
and U9979 (N_9979,N_8322,N_8989);
or U9980 (N_9980,N_8388,N_8376);
nand U9981 (N_9981,N_8888,N_8724);
nor U9982 (N_9982,N_8990,N_8521);
nand U9983 (N_9983,N_8594,N_8089);
nor U9984 (N_9984,N_8839,N_8424);
and U9985 (N_9985,N_8012,N_8875);
nor U9986 (N_9986,N_8558,N_8767);
nor U9987 (N_9987,N_8203,N_8982);
or U9988 (N_9988,N_8542,N_8217);
nand U9989 (N_9989,N_8850,N_8284);
nor U9990 (N_9990,N_8630,N_8998);
nor U9991 (N_9991,N_8535,N_8317);
nand U9992 (N_9992,N_8187,N_8205);
or U9993 (N_9993,N_8785,N_8655);
nand U9994 (N_9994,N_8947,N_8913);
or U9995 (N_9995,N_8887,N_8255);
nand U9996 (N_9996,N_8896,N_8130);
nor U9997 (N_9997,N_8375,N_8437);
or U9998 (N_9998,N_8585,N_8299);
or U9999 (N_9999,N_8833,N_8343);
xnor U10000 (N_10000,N_9877,N_9874);
nor U10001 (N_10001,N_9083,N_9880);
and U10002 (N_10002,N_9522,N_9887);
or U10003 (N_10003,N_9638,N_9329);
and U10004 (N_10004,N_9573,N_9983);
or U10005 (N_10005,N_9871,N_9389);
nand U10006 (N_10006,N_9636,N_9507);
and U10007 (N_10007,N_9323,N_9563);
or U10008 (N_10008,N_9431,N_9778);
nand U10009 (N_10009,N_9729,N_9174);
and U10010 (N_10010,N_9049,N_9524);
nand U10011 (N_10011,N_9761,N_9833);
nor U10012 (N_10012,N_9053,N_9666);
or U10013 (N_10013,N_9660,N_9190);
nor U10014 (N_10014,N_9099,N_9231);
nor U10015 (N_10015,N_9500,N_9537);
and U10016 (N_10016,N_9753,N_9069);
and U10017 (N_10017,N_9107,N_9813);
nand U10018 (N_10018,N_9001,N_9037);
and U10019 (N_10019,N_9978,N_9162);
and U10020 (N_10020,N_9979,N_9624);
and U10021 (N_10021,N_9044,N_9501);
xnor U10022 (N_10022,N_9139,N_9548);
nor U10023 (N_10023,N_9203,N_9909);
or U10024 (N_10024,N_9294,N_9234);
nor U10025 (N_10025,N_9052,N_9726);
nand U10026 (N_10026,N_9351,N_9590);
nor U10027 (N_10027,N_9187,N_9773);
nor U10028 (N_10028,N_9487,N_9169);
nand U10029 (N_10029,N_9132,N_9095);
nand U10030 (N_10030,N_9968,N_9568);
nand U10031 (N_10031,N_9752,N_9505);
xnor U10032 (N_10032,N_9683,N_9807);
or U10033 (N_10033,N_9796,N_9863);
nand U10034 (N_10034,N_9045,N_9461);
nor U10035 (N_10035,N_9677,N_9919);
or U10036 (N_10036,N_9885,N_9027);
nor U10037 (N_10037,N_9712,N_9376);
and U10038 (N_10038,N_9895,N_9738);
nand U10039 (N_10039,N_9516,N_9763);
nand U10040 (N_10040,N_9101,N_9743);
and U10041 (N_10041,N_9504,N_9082);
nand U10042 (N_10042,N_9582,N_9064);
nor U10043 (N_10043,N_9239,N_9583);
or U10044 (N_10044,N_9612,N_9555);
and U10045 (N_10045,N_9702,N_9920);
or U10046 (N_10046,N_9433,N_9759);
nor U10047 (N_10047,N_9365,N_9302);
and U10048 (N_10048,N_9454,N_9350);
and U10049 (N_10049,N_9549,N_9198);
nand U10050 (N_10050,N_9685,N_9426);
or U10051 (N_10051,N_9337,N_9087);
nand U10052 (N_10052,N_9896,N_9934);
and U10053 (N_10053,N_9442,N_9315);
xnor U10054 (N_10054,N_9314,N_9894);
and U10055 (N_10055,N_9085,N_9318);
nand U10056 (N_10056,N_9875,N_9274);
xnor U10057 (N_10057,N_9219,N_9960);
nand U10058 (N_10058,N_9710,N_9646);
xor U10059 (N_10059,N_9211,N_9301);
nand U10060 (N_10060,N_9236,N_9765);
nor U10061 (N_10061,N_9860,N_9286);
nor U10062 (N_10062,N_9688,N_9912);
nand U10063 (N_10063,N_9380,N_9950);
nor U10064 (N_10064,N_9445,N_9385);
and U10065 (N_10065,N_9453,N_9496);
and U10066 (N_10066,N_9072,N_9040);
or U10067 (N_10067,N_9870,N_9892);
nand U10068 (N_10068,N_9249,N_9526);
or U10069 (N_10069,N_9299,N_9093);
xnor U10070 (N_10070,N_9075,N_9260);
nor U10071 (N_10071,N_9071,N_9471);
xnor U10072 (N_10072,N_9525,N_9626);
xor U10073 (N_10073,N_9556,N_9593);
or U10074 (N_10074,N_9475,N_9921);
and U10075 (N_10075,N_9576,N_9747);
nand U10076 (N_10076,N_9366,N_9240);
or U10077 (N_10077,N_9937,N_9956);
or U10078 (N_10078,N_9775,N_9109);
nand U10079 (N_10079,N_9756,N_9316);
or U10080 (N_10080,N_9066,N_9022);
xor U10081 (N_10081,N_9403,N_9485);
nand U10082 (N_10082,N_9742,N_9119);
nor U10083 (N_10083,N_9489,N_9985);
xor U10084 (N_10084,N_9558,N_9336);
and U10085 (N_10085,N_9657,N_9283);
nand U10086 (N_10086,N_9208,N_9760);
or U10087 (N_10087,N_9347,N_9546);
nor U10088 (N_10088,N_9217,N_9514);
or U10089 (N_10089,N_9331,N_9220);
and U10090 (N_10090,N_9594,N_9922);
or U10091 (N_10091,N_9459,N_9758);
nor U10092 (N_10092,N_9928,N_9395);
and U10093 (N_10093,N_9751,N_9907);
or U10094 (N_10094,N_9958,N_9357);
and U10095 (N_10095,N_9797,N_9477);
nand U10096 (N_10096,N_9000,N_9084);
nor U10097 (N_10097,N_9488,N_9021);
or U10098 (N_10098,N_9237,N_9016);
or U10099 (N_10099,N_9003,N_9635);
nand U10100 (N_10100,N_9447,N_9961);
or U10101 (N_10101,N_9716,N_9312);
and U10102 (N_10102,N_9559,N_9964);
nor U10103 (N_10103,N_9076,N_9035);
and U10104 (N_10104,N_9725,N_9023);
and U10105 (N_10105,N_9146,N_9223);
or U10106 (N_10106,N_9161,N_9578);
nor U10107 (N_10107,N_9906,N_9104);
nand U10108 (N_10108,N_9838,N_9543);
and U10109 (N_10109,N_9705,N_9882);
or U10110 (N_10110,N_9618,N_9793);
or U10111 (N_10111,N_9070,N_9349);
nor U10112 (N_10112,N_9888,N_9814);
or U10113 (N_10113,N_9566,N_9293);
or U10114 (N_10114,N_9135,N_9984);
nor U10115 (N_10115,N_9105,N_9630);
nand U10116 (N_10116,N_9383,N_9017);
nor U10117 (N_10117,N_9057,N_9143);
nor U10118 (N_10118,N_9943,N_9258);
nor U10119 (N_10119,N_9899,N_9295);
nor U10120 (N_10120,N_9289,N_9317);
and U10121 (N_10121,N_9408,N_9930);
nand U10122 (N_10122,N_9762,N_9873);
xnor U10123 (N_10123,N_9340,N_9739);
or U10124 (N_10124,N_9569,N_9042);
and U10125 (N_10125,N_9659,N_9149);
and U10126 (N_10126,N_9328,N_9263);
and U10127 (N_10127,N_9798,N_9370);
and U10128 (N_10128,N_9415,N_9966);
and U10129 (N_10129,N_9640,N_9138);
xor U10130 (N_10130,N_9118,N_9128);
or U10131 (N_10131,N_9100,N_9163);
nor U10132 (N_10132,N_9772,N_9451);
or U10133 (N_10133,N_9073,N_9839);
nor U10134 (N_10134,N_9939,N_9734);
nor U10135 (N_10135,N_9290,N_9338);
nor U10136 (N_10136,N_9440,N_9605);
nor U10137 (N_10137,N_9430,N_9777);
nor U10138 (N_10138,N_9722,N_9086);
and U10139 (N_10139,N_9131,N_9846);
nand U10140 (N_10140,N_9615,N_9717);
or U10141 (N_10141,N_9450,N_9058);
or U10142 (N_10142,N_9924,N_9697);
or U10143 (N_10143,N_9932,N_9209);
and U10144 (N_10144,N_9266,N_9221);
nor U10145 (N_10145,N_9868,N_9804);
or U10146 (N_10146,N_9390,N_9836);
or U10147 (N_10147,N_9092,N_9661);
and U10148 (N_10148,N_9378,N_9973);
and U10149 (N_10149,N_9495,N_9650);
and U10150 (N_10150,N_9394,N_9009);
nor U10151 (N_10151,N_9754,N_9173);
and U10152 (N_10152,N_9359,N_9330);
xor U10153 (N_10153,N_9832,N_9847);
or U10154 (N_10154,N_9438,N_9554);
nor U10155 (N_10155,N_9464,N_9157);
nand U10156 (N_10156,N_9801,N_9474);
nor U10157 (N_10157,N_9925,N_9553);
xor U10158 (N_10158,N_9421,N_9781);
and U10159 (N_10159,N_9903,N_9625);
nor U10160 (N_10160,N_9872,N_9610);
nand U10161 (N_10161,N_9935,N_9959);
and U10162 (N_10162,N_9602,N_9397);
nand U10163 (N_10163,N_9156,N_9680);
nand U10164 (N_10164,N_9986,N_9372);
or U10165 (N_10165,N_9195,N_9965);
nor U10166 (N_10166,N_9998,N_9831);
xnor U10167 (N_10167,N_9923,N_9186);
and U10168 (N_10168,N_9669,N_9641);
nand U10169 (N_10169,N_9435,N_9374);
nor U10170 (N_10170,N_9769,N_9377);
nand U10171 (N_10171,N_9013,N_9422);
or U10172 (N_10172,N_9326,N_9288);
nand U10173 (N_10173,N_9898,N_9499);
and U10174 (N_10174,N_9929,N_9355);
or U10175 (N_10175,N_9110,N_9437);
nand U10176 (N_10176,N_9207,N_9183);
or U10177 (N_10177,N_9160,N_9028);
nand U10178 (N_10178,N_9749,N_9396);
and U10179 (N_10179,N_9571,N_9165);
nand U10180 (N_10180,N_9424,N_9992);
or U10181 (N_10181,N_9147,N_9835);
and U10182 (N_10182,N_9539,N_9155);
xor U10183 (N_10183,N_9029,N_9024);
nor U10184 (N_10184,N_9348,N_9989);
xnor U10185 (N_10185,N_9994,N_9371);
nor U10186 (N_10186,N_9402,N_9213);
xor U10187 (N_10187,N_9393,N_9202);
xnor U10188 (N_10188,N_9088,N_9609);
nor U10189 (N_10189,N_9369,N_9731);
and U10190 (N_10190,N_9681,N_9812);
nand U10191 (N_10191,N_9164,N_9060);
nand U10192 (N_10192,N_9809,N_9458);
and U10193 (N_10193,N_9200,N_9787);
and U10194 (N_10194,N_9551,N_9764);
and U10195 (N_10195,N_9611,N_9810);
xor U10196 (N_10196,N_9354,N_9206);
or U10197 (N_10197,N_9952,N_9056);
nand U10198 (N_10198,N_9015,N_9830);
nand U10199 (N_10199,N_9005,N_9840);
xnor U10200 (N_10200,N_9512,N_9168);
and U10201 (N_10201,N_9025,N_9278);
or U10202 (N_10202,N_9770,N_9837);
or U10203 (N_10203,N_9261,N_9419);
xor U10204 (N_10204,N_9910,N_9343);
or U10205 (N_10205,N_9276,N_9470);
nor U10206 (N_10206,N_9478,N_9598);
and U10207 (N_10207,N_9241,N_9905);
nor U10208 (N_10208,N_9736,N_9308);
nor U10209 (N_10209,N_9434,N_9783);
or U10210 (N_10210,N_9311,N_9363);
or U10211 (N_10211,N_9901,N_9439);
nand U10212 (N_10212,N_9412,N_9648);
nand U10213 (N_10213,N_9281,N_9197);
nand U10214 (N_10214,N_9825,N_9916);
xor U10215 (N_10215,N_9955,N_9230);
nor U10216 (N_10216,N_9802,N_9843);
or U10217 (N_10217,N_9006,N_9720);
xor U10218 (N_10218,N_9800,N_9382);
nor U10219 (N_10219,N_9491,N_9120);
or U10220 (N_10220,N_9864,N_9745);
nor U10221 (N_10221,N_9228,N_9628);
nor U10222 (N_10222,N_9352,N_9446);
or U10223 (N_10223,N_9255,N_9560);
nor U10224 (N_10224,N_9869,N_9970);
or U10225 (N_10225,N_9719,N_9038);
nand U10226 (N_10226,N_9094,N_9841);
nor U10227 (N_10227,N_9490,N_9307);
nand U10228 (N_10228,N_9699,N_9353);
nor U10229 (N_10229,N_9232,N_9178);
or U10230 (N_10230,N_9790,N_9091);
nor U10231 (N_10231,N_9805,N_9806);
xnor U10232 (N_10232,N_9121,N_9601);
xor U10233 (N_10233,N_9185,N_9816);
and U10234 (N_10234,N_9361,N_9218);
nor U10235 (N_10235,N_9243,N_9711);
xor U10236 (N_10236,N_9997,N_9401);
nand U10237 (N_10237,N_9740,N_9862);
nand U10238 (N_10238,N_9297,N_9849);
nor U10239 (N_10239,N_9616,N_9649);
xor U10240 (N_10240,N_9858,N_9492);
or U10241 (N_10241,N_9768,N_9730);
xnor U10242 (N_10242,N_9327,N_9528);
and U10243 (N_10243,N_9346,N_9002);
and U10244 (N_10244,N_9980,N_9334);
and U10245 (N_10245,N_9713,N_9684);
or U10246 (N_10246,N_9991,N_9233);
nand U10247 (N_10247,N_9589,N_9229);
and U10248 (N_10248,N_9866,N_9196);
nand U10249 (N_10249,N_9667,N_9245);
nor U10250 (N_10250,N_9090,N_9031);
nor U10251 (N_10251,N_9951,N_9420);
or U10252 (N_10252,N_9269,N_9767);
or U10253 (N_10253,N_9159,N_9853);
nor U10254 (N_10254,N_9786,N_9384);
or U10255 (N_10255,N_9913,N_9134);
xor U10256 (N_10256,N_9172,N_9788);
or U10257 (N_10257,N_9803,N_9727);
nor U10258 (N_10258,N_9857,N_9513);
nand U10259 (N_10259,N_9141,N_9116);
and U10260 (N_10260,N_9409,N_9339);
or U10261 (N_10261,N_9448,N_9126);
nor U10262 (N_10262,N_9476,N_9606);
nor U10263 (N_10263,N_9158,N_9686);
nor U10264 (N_10264,N_9123,N_9672);
or U10265 (N_10265,N_9530,N_9881);
nor U10266 (N_10266,N_9962,N_9285);
and U10267 (N_10267,N_9482,N_9463);
and U10268 (N_10268,N_9242,N_9981);
and U10269 (N_10269,N_9519,N_9815);
and U10270 (N_10270,N_9527,N_9580);
or U10271 (N_10271,N_9272,N_9262);
nor U10272 (N_10272,N_9851,N_9122);
xor U10273 (N_10273,N_9404,N_9254);
and U10274 (N_10274,N_9826,N_9642);
or U10275 (N_10275,N_9971,N_9591);
and U10276 (N_10276,N_9055,N_9577);
nor U10277 (N_10277,N_9063,N_9225);
or U10278 (N_10278,N_9226,N_9368);
nor U10279 (N_10279,N_9545,N_9400);
nor U10280 (N_10280,N_9189,N_9631);
or U10281 (N_10281,N_9235,N_9171);
nor U10282 (N_10282,N_9204,N_9808);
nor U10283 (N_10283,N_9144,N_9309);
nand U10284 (N_10284,N_9750,N_9671);
nor U10285 (N_10285,N_9452,N_9608);
nand U10286 (N_10286,N_9222,N_9124);
and U10287 (N_10287,N_9647,N_9416);
nand U10288 (N_10288,N_9637,N_9665);
or U10289 (N_10289,N_9592,N_9969);
xor U10290 (N_10290,N_9304,N_9678);
nor U10291 (N_10291,N_9982,N_9322);
or U10292 (N_10292,N_9506,N_9620);
nand U10293 (N_10293,N_9707,N_9547);
nor U10294 (N_10294,N_9523,N_9142);
xor U10295 (N_10295,N_9305,N_9561);
nand U10296 (N_10296,N_9709,N_9466);
or U10297 (N_10297,N_9014,N_9785);
nand U10298 (N_10298,N_9046,N_9565);
xnor U10299 (N_10299,N_9509,N_9067);
nor U10300 (N_10300,N_9534,N_9824);
nand U10301 (N_10301,N_9460,N_9388);
and U10302 (N_10302,N_9867,N_9427);
nor U10303 (N_10303,N_9472,N_9776);
nand U10304 (N_10304,N_9948,N_9940);
xnor U10305 (N_10305,N_9270,N_9728);
nand U10306 (N_10306,N_9498,N_9247);
nand U10307 (N_10307,N_9655,N_9303);
xor U10308 (N_10308,N_9879,N_9536);
nand U10309 (N_10309,N_9782,N_9850);
or U10310 (N_10310,N_9938,N_9700);
or U10311 (N_10311,N_9273,N_9191);
xnor U10312 (N_10312,N_9941,N_9737);
nand U10313 (N_10313,N_9148,N_9170);
or U10314 (N_10314,N_9199,N_9856);
and U10315 (N_10315,N_9947,N_9227);
and U10316 (N_10316,N_9428,N_9517);
nand U10317 (N_10317,N_9999,N_9410);
xnor U10318 (N_10318,N_9033,N_9600);
and U10319 (N_10319,N_9391,N_9257);
or U10320 (N_10320,N_9387,N_9845);
xnor U10321 (N_10321,N_9581,N_9486);
and U10322 (N_10322,N_9531,N_9967);
or U10323 (N_10323,N_9429,N_9244);
and U10324 (N_10324,N_9570,N_9030);
nand U10325 (N_10325,N_9818,N_9819);
nor U10326 (N_10326,N_9585,N_9399);
and U10327 (N_10327,N_9047,N_9356);
or U10328 (N_10328,N_9579,N_9541);
nand U10329 (N_10329,N_9633,N_9051);
nor U10330 (N_10330,N_9724,N_9639);
and U10331 (N_10331,N_9976,N_9306);
and U10332 (N_10332,N_9518,N_9521);
nand U10333 (N_10333,N_9990,N_9617);
and U10334 (N_10334,N_9298,N_9904);
nand U10335 (N_10335,N_9953,N_9893);
and U10336 (N_10336,N_9876,N_9908);
nor U10337 (N_10337,N_9567,N_9820);
or U10338 (N_10338,N_9004,N_9714);
or U10339 (N_10339,N_9373,N_9996);
or U10340 (N_10340,N_9766,N_9644);
and U10341 (N_10341,N_9654,N_9103);
xnor U10342 (N_10342,N_9693,N_9535);
and U10343 (N_10343,N_9332,N_9175);
nor U10344 (N_10344,N_9732,N_9279);
or U10345 (N_10345,N_9643,N_9861);
and U10346 (N_10346,N_9687,N_9020);
nand U10347 (N_10347,N_9675,N_9417);
or U10348 (N_10348,N_9811,N_9081);
or U10349 (N_10349,N_9629,N_9918);
nand U10350 (N_10350,N_9375,N_9153);
nand U10351 (N_10351,N_9603,N_9268);
nand U10352 (N_10352,N_9596,N_9529);
and U10353 (N_10353,N_9455,N_9562);
nand U10354 (N_10354,N_9413,N_9167);
or U10355 (N_10355,N_9250,N_9050);
or U10356 (N_10356,N_9265,N_9089);
and U10357 (N_10357,N_9456,N_9133);
nor U10358 (N_10358,N_9480,N_9721);
nor U10359 (N_10359,N_9689,N_9313);
and U10360 (N_10360,N_9411,N_9036);
xor U10361 (N_10361,N_9886,N_9744);
and U10362 (N_10362,N_9193,N_9364);
xnor U10363 (N_10363,N_9607,N_9587);
or U10364 (N_10364,N_9271,N_9102);
nand U10365 (N_10365,N_9310,N_9564);
nand U10366 (N_10366,N_9280,N_9398);
and U10367 (N_10367,N_9344,N_9188);
and U10368 (N_10368,N_9345,N_9884);
and U10369 (N_10369,N_9321,N_9622);
nand U10370 (N_10370,N_9708,N_9771);
or U10371 (N_10371,N_9414,N_9897);
nor U10372 (N_10372,N_9077,N_9432);
nor U10373 (N_10373,N_9902,N_9360);
or U10374 (N_10374,N_9041,N_9696);
nor U10375 (N_10375,N_9214,N_9748);
nand U10376 (N_10376,N_9854,N_9406);
nor U10377 (N_10377,N_9484,N_9865);
or U10378 (N_10378,N_9113,N_9248);
nor U10379 (N_10379,N_9179,N_9098);
nand U10380 (N_10380,N_9386,N_9392);
or U10381 (N_10381,N_9441,N_9292);
nand U10382 (N_10382,N_9176,N_9205);
and U10383 (N_10383,N_9829,N_9619);
xor U10384 (N_10384,N_9074,N_9467);
or U10385 (N_10385,N_9933,N_9718);
nor U10386 (N_10386,N_9936,N_9468);
or U10387 (N_10387,N_9817,N_9859);
nand U10388 (N_10388,N_9652,N_9510);
and U10389 (N_10389,N_9735,N_9481);
and U10390 (N_10390,N_9828,N_9151);
and U10391 (N_10391,N_9575,N_9963);
or U10392 (N_10392,N_9140,N_9694);
and U10393 (N_10393,N_9341,N_9927);
nor U10394 (N_10394,N_9878,N_9502);
nand U10395 (N_10395,N_9026,N_9129);
or U10396 (N_10396,N_9515,N_9827);
nor U10397 (N_10397,N_9325,N_9425);
and U10398 (N_10398,N_9212,N_9457);
nand U10399 (N_10399,N_9795,N_9698);
or U10400 (N_10400,N_9112,N_9848);
xnor U10401 (N_10401,N_9673,N_9703);
and U10402 (N_10402,N_9931,N_9111);
or U10403 (N_10403,N_9018,N_9078);
or U10404 (N_10404,N_9706,N_9127);
nand U10405 (N_10405,N_9469,N_9358);
or U10406 (N_10406,N_9957,N_9613);
and U10407 (N_10407,N_9946,N_9949);
xor U10408 (N_10408,N_9224,N_9494);
nor U10409 (N_10409,N_9043,N_9993);
nor U10410 (N_10410,N_9789,N_9079);
xnor U10411 (N_10411,N_9180,N_9096);
or U10412 (N_10412,N_9125,N_9267);
xnor U10413 (N_10413,N_9059,N_9690);
nand U10414 (N_10414,N_9479,N_9658);
nand U10415 (N_10415,N_9300,N_9599);
nand U10416 (N_10416,N_9890,N_9115);
xor U10417 (N_10417,N_9588,N_9114);
nand U10418 (N_10418,N_9215,N_9503);
nor U10419 (N_10419,N_9852,N_9799);
nor U10420 (N_10420,N_9319,N_9842);
or U10421 (N_10421,N_9627,N_9520);
and U10422 (N_10422,N_9911,N_9032);
nand U10423 (N_10423,N_9844,N_9900);
nor U10424 (N_10424,N_9855,N_9011);
or U10425 (N_10425,N_9915,N_9574);
xor U10426 (N_10426,N_9423,N_9282);
and U10427 (N_10427,N_9823,N_9645);
nor U10428 (N_10428,N_9715,N_9988);
nand U10429 (N_10429,N_9741,N_9791);
nor U10430 (N_10430,N_9792,N_9152);
or U10431 (N_10431,N_9259,N_9550);
nor U10432 (N_10432,N_9584,N_9597);
nand U10433 (N_10433,N_9511,N_9977);
xnor U10434 (N_10434,N_9508,N_9604);
or U10435 (N_10435,N_9651,N_9670);
nand U10436 (N_10436,N_9062,N_9061);
nor U10437 (N_10437,N_9614,N_9108);
or U10438 (N_10438,N_9662,N_9019);
and U10439 (N_10439,N_9664,N_9883);
nand U10440 (N_10440,N_9342,N_9945);
and U10441 (N_10441,N_9238,N_9917);
nand U10442 (N_10442,N_9540,N_9595);
and U10443 (N_10443,N_9251,N_9889);
nor U10444 (N_10444,N_9333,N_9277);
and U10445 (N_10445,N_9891,N_9632);
nor U10446 (N_10446,N_9780,N_9733);
nand U10447 (N_10447,N_9834,N_9944);
xnor U10448 (N_10448,N_9533,N_9379);
or U10449 (N_10449,N_9012,N_9975);
xnor U10450 (N_10450,N_9544,N_9253);
or U10451 (N_10451,N_9822,N_9821);
and U10452 (N_10452,N_9972,N_9008);
nand U10453 (N_10453,N_9668,N_9291);
and U10454 (N_10454,N_9065,N_9926);
or U10455 (N_10455,N_9210,N_9653);
nand U10456 (N_10456,N_9942,N_9246);
nor U10457 (N_10457,N_9177,N_9695);
xnor U10458 (N_10458,N_9462,N_9723);
nor U10459 (N_10459,N_9405,N_9381);
and U10460 (N_10460,N_9691,N_9995);
nand U10461 (N_10461,N_9154,N_9552);
nor U10462 (N_10462,N_9444,N_9572);
and U10463 (N_10463,N_9007,N_9256);
nand U10464 (N_10464,N_9623,N_9166);
and U10465 (N_10465,N_9068,N_9216);
or U10466 (N_10466,N_9048,N_9784);
nand U10467 (N_10467,N_9682,N_9150);
nor U10468 (N_10468,N_9034,N_9145);
and U10469 (N_10469,N_9182,N_9701);
and U10470 (N_10470,N_9252,N_9586);
or U10471 (N_10471,N_9974,N_9264);
nand U10472 (N_10472,N_9914,N_9275);
and U10473 (N_10473,N_9181,N_9954);
xnor U10474 (N_10474,N_9296,N_9493);
xor U10475 (N_10475,N_9130,N_9757);
xor U10476 (N_10476,N_9497,N_9755);
xor U10477 (N_10477,N_9676,N_9794);
nand U10478 (N_10478,N_9054,N_9746);
or U10479 (N_10479,N_9692,N_9407);
nand U10480 (N_10480,N_9449,N_9184);
nand U10481 (N_10481,N_9418,N_9774);
nor U10482 (N_10482,N_9137,N_9483);
nor U10483 (N_10483,N_9542,N_9324);
nand U10484 (N_10484,N_9679,N_9538);
nand U10485 (N_10485,N_9287,N_9656);
nand U10486 (N_10486,N_9080,N_9201);
nor U10487 (N_10487,N_9634,N_9443);
and U10488 (N_10488,N_9136,N_9367);
nor U10489 (N_10489,N_9532,N_9704);
and U10490 (N_10490,N_9557,N_9779);
nor U10491 (N_10491,N_9010,N_9663);
nor U10492 (N_10492,N_9320,N_9194);
xnor U10493 (N_10493,N_9465,N_9039);
and U10494 (N_10494,N_9117,N_9362);
nor U10495 (N_10495,N_9106,N_9436);
or U10496 (N_10496,N_9284,N_9473);
xnor U10497 (N_10497,N_9097,N_9674);
xor U10498 (N_10498,N_9621,N_9987);
xnor U10499 (N_10499,N_9192,N_9335);
nand U10500 (N_10500,N_9052,N_9555);
and U10501 (N_10501,N_9800,N_9770);
or U10502 (N_10502,N_9991,N_9955);
or U10503 (N_10503,N_9797,N_9182);
and U10504 (N_10504,N_9689,N_9371);
and U10505 (N_10505,N_9114,N_9826);
nand U10506 (N_10506,N_9464,N_9178);
xor U10507 (N_10507,N_9527,N_9635);
and U10508 (N_10508,N_9781,N_9554);
and U10509 (N_10509,N_9444,N_9560);
or U10510 (N_10510,N_9945,N_9198);
nand U10511 (N_10511,N_9577,N_9502);
nand U10512 (N_10512,N_9916,N_9740);
and U10513 (N_10513,N_9823,N_9489);
nand U10514 (N_10514,N_9947,N_9976);
or U10515 (N_10515,N_9641,N_9550);
nor U10516 (N_10516,N_9687,N_9234);
or U10517 (N_10517,N_9434,N_9951);
or U10518 (N_10518,N_9737,N_9570);
nor U10519 (N_10519,N_9049,N_9412);
or U10520 (N_10520,N_9817,N_9508);
or U10521 (N_10521,N_9233,N_9270);
and U10522 (N_10522,N_9190,N_9694);
nor U10523 (N_10523,N_9902,N_9681);
or U10524 (N_10524,N_9831,N_9130);
nor U10525 (N_10525,N_9363,N_9429);
and U10526 (N_10526,N_9564,N_9568);
or U10527 (N_10527,N_9855,N_9972);
or U10528 (N_10528,N_9287,N_9240);
and U10529 (N_10529,N_9160,N_9971);
nand U10530 (N_10530,N_9402,N_9181);
or U10531 (N_10531,N_9792,N_9397);
nor U10532 (N_10532,N_9377,N_9664);
or U10533 (N_10533,N_9363,N_9017);
and U10534 (N_10534,N_9107,N_9956);
xnor U10535 (N_10535,N_9758,N_9142);
nand U10536 (N_10536,N_9068,N_9683);
and U10537 (N_10537,N_9535,N_9314);
nor U10538 (N_10538,N_9495,N_9668);
nand U10539 (N_10539,N_9786,N_9268);
and U10540 (N_10540,N_9276,N_9221);
or U10541 (N_10541,N_9326,N_9085);
xor U10542 (N_10542,N_9516,N_9266);
nor U10543 (N_10543,N_9039,N_9774);
or U10544 (N_10544,N_9923,N_9385);
and U10545 (N_10545,N_9192,N_9722);
and U10546 (N_10546,N_9157,N_9737);
or U10547 (N_10547,N_9736,N_9657);
or U10548 (N_10548,N_9830,N_9543);
and U10549 (N_10549,N_9465,N_9638);
and U10550 (N_10550,N_9117,N_9700);
or U10551 (N_10551,N_9593,N_9436);
or U10552 (N_10552,N_9726,N_9201);
nor U10553 (N_10553,N_9119,N_9758);
and U10554 (N_10554,N_9926,N_9624);
or U10555 (N_10555,N_9082,N_9960);
or U10556 (N_10556,N_9016,N_9889);
or U10557 (N_10557,N_9786,N_9037);
or U10558 (N_10558,N_9498,N_9240);
or U10559 (N_10559,N_9958,N_9234);
xor U10560 (N_10560,N_9561,N_9949);
nor U10561 (N_10561,N_9854,N_9830);
nor U10562 (N_10562,N_9692,N_9116);
nor U10563 (N_10563,N_9815,N_9438);
nor U10564 (N_10564,N_9294,N_9707);
and U10565 (N_10565,N_9278,N_9376);
or U10566 (N_10566,N_9085,N_9182);
nor U10567 (N_10567,N_9899,N_9507);
and U10568 (N_10568,N_9433,N_9649);
nand U10569 (N_10569,N_9615,N_9754);
nor U10570 (N_10570,N_9044,N_9836);
and U10571 (N_10571,N_9460,N_9845);
and U10572 (N_10572,N_9306,N_9931);
or U10573 (N_10573,N_9358,N_9939);
nor U10574 (N_10574,N_9937,N_9240);
nor U10575 (N_10575,N_9361,N_9950);
nand U10576 (N_10576,N_9056,N_9783);
and U10577 (N_10577,N_9654,N_9843);
nand U10578 (N_10578,N_9208,N_9792);
or U10579 (N_10579,N_9830,N_9351);
nand U10580 (N_10580,N_9324,N_9529);
nor U10581 (N_10581,N_9616,N_9307);
nor U10582 (N_10582,N_9878,N_9432);
or U10583 (N_10583,N_9485,N_9673);
nand U10584 (N_10584,N_9678,N_9811);
and U10585 (N_10585,N_9149,N_9476);
nand U10586 (N_10586,N_9691,N_9353);
nor U10587 (N_10587,N_9915,N_9816);
and U10588 (N_10588,N_9381,N_9800);
and U10589 (N_10589,N_9781,N_9954);
xnor U10590 (N_10590,N_9521,N_9543);
and U10591 (N_10591,N_9521,N_9504);
nor U10592 (N_10592,N_9922,N_9627);
nor U10593 (N_10593,N_9490,N_9669);
and U10594 (N_10594,N_9824,N_9933);
nand U10595 (N_10595,N_9681,N_9408);
and U10596 (N_10596,N_9232,N_9650);
or U10597 (N_10597,N_9245,N_9679);
nor U10598 (N_10598,N_9744,N_9860);
or U10599 (N_10599,N_9387,N_9712);
nand U10600 (N_10600,N_9540,N_9770);
nor U10601 (N_10601,N_9212,N_9247);
and U10602 (N_10602,N_9720,N_9197);
or U10603 (N_10603,N_9000,N_9151);
nor U10604 (N_10604,N_9726,N_9429);
and U10605 (N_10605,N_9355,N_9419);
xnor U10606 (N_10606,N_9636,N_9663);
nor U10607 (N_10607,N_9221,N_9943);
xor U10608 (N_10608,N_9767,N_9417);
and U10609 (N_10609,N_9754,N_9061);
or U10610 (N_10610,N_9870,N_9255);
and U10611 (N_10611,N_9925,N_9657);
nor U10612 (N_10612,N_9428,N_9814);
nand U10613 (N_10613,N_9638,N_9573);
nor U10614 (N_10614,N_9808,N_9365);
or U10615 (N_10615,N_9509,N_9925);
nor U10616 (N_10616,N_9656,N_9709);
or U10617 (N_10617,N_9758,N_9290);
or U10618 (N_10618,N_9833,N_9668);
nor U10619 (N_10619,N_9248,N_9281);
xnor U10620 (N_10620,N_9296,N_9490);
and U10621 (N_10621,N_9694,N_9856);
nand U10622 (N_10622,N_9031,N_9468);
and U10623 (N_10623,N_9753,N_9569);
nand U10624 (N_10624,N_9108,N_9093);
or U10625 (N_10625,N_9597,N_9279);
and U10626 (N_10626,N_9040,N_9819);
nand U10627 (N_10627,N_9831,N_9825);
and U10628 (N_10628,N_9310,N_9024);
xnor U10629 (N_10629,N_9843,N_9554);
nand U10630 (N_10630,N_9166,N_9133);
nand U10631 (N_10631,N_9736,N_9379);
and U10632 (N_10632,N_9281,N_9101);
or U10633 (N_10633,N_9612,N_9542);
and U10634 (N_10634,N_9170,N_9918);
or U10635 (N_10635,N_9641,N_9092);
nor U10636 (N_10636,N_9901,N_9366);
nand U10637 (N_10637,N_9402,N_9428);
nand U10638 (N_10638,N_9574,N_9482);
nor U10639 (N_10639,N_9218,N_9579);
nor U10640 (N_10640,N_9497,N_9048);
nand U10641 (N_10641,N_9666,N_9969);
or U10642 (N_10642,N_9167,N_9608);
nor U10643 (N_10643,N_9826,N_9270);
or U10644 (N_10644,N_9591,N_9063);
nand U10645 (N_10645,N_9211,N_9623);
nor U10646 (N_10646,N_9002,N_9387);
nor U10647 (N_10647,N_9241,N_9184);
and U10648 (N_10648,N_9920,N_9670);
or U10649 (N_10649,N_9831,N_9083);
nor U10650 (N_10650,N_9140,N_9742);
nand U10651 (N_10651,N_9403,N_9117);
nand U10652 (N_10652,N_9166,N_9400);
or U10653 (N_10653,N_9624,N_9606);
and U10654 (N_10654,N_9762,N_9894);
or U10655 (N_10655,N_9042,N_9695);
nand U10656 (N_10656,N_9659,N_9769);
xor U10657 (N_10657,N_9357,N_9209);
nor U10658 (N_10658,N_9176,N_9471);
and U10659 (N_10659,N_9152,N_9728);
nand U10660 (N_10660,N_9716,N_9659);
xnor U10661 (N_10661,N_9105,N_9492);
nand U10662 (N_10662,N_9792,N_9521);
and U10663 (N_10663,N_9165,N_9884);
and U10664 (N_10664,N_9934,N_9425);
or U10665 (N_10665,N_9021,N_9712);
and U10666 (N_10666,N_9319,N_9709);
nand U10667 (N_10667,N_9653,N_9580);
nand U10668 (N_10668,N_9627,N_9900);
nor U10669 (N_10669,N_9939,N_9889);
and U10670 (N_10670,N_9683,N_9325);
and U10671 (N_10671,N_9583,N_9912);
nand U10672 (N_10672,N_9379,N_9722);
nand U10673 (N_10673,N_9014,N_9997);
and U10674 (N_10674,N_9588,N_9210);
and U10675 (N_10675,N_9915,N_9584);
nand U10676 (N_10676,N_9604,N_9246);
nand U10677 (N_10677,N_9180,N_9683);
nand U10678 (N_10678,N_9333,N_9550);
nor U10679 (N_10679,N_9286,N_9129);
nor U10680 (N_10680,N_9652,N_9434);
nand U10681 (N_10681,N_9429,N_9150);
and U10682 (N_10682,N_9604,N_9268);
nor U10683 (N_10683,N_9535,N_9575);
nand U10684 (N_10684,N_9898,N_9821);
or U10685 (N_10685,N_9883,N_9223);
nor U10686 (N_10686,N_9837,N_9700);
nand U10687 (N_10687,N_9246,N_9071);
nor U10688 (N_10688,N_9451,N_9088);
nor U10689 (N_10689,N_9801,N_9982);
and U10690 (N_10690,N_9455,N_9830);
and U10691 (N_10691,N_9372,N_9701);
nand U10692 (N_10692,N_9785,N_9489);
or U10693 (N_10693,N_9585,N_9352);
nor U10694 (N_10694,N_9051,N_9993);
xor U10695 (N_10695,N_9264,N_9607);
or U10696 (N_10696,N_9218,N_9740);
nand U10697 (N_10697,N_9107,N_9309);
nand U10698 (N_10698,N_9078,N_9413);
nand U10699 (N_10699,N_9624,N_9167);
and U10700 (N_10700,N_9557,N_9275);
and U10701 (N_10701,N_9659,N_9672);
or U10702 (N_10702,N_9915,N_9585);
xnor U10703 (N_10703,N_9002,N_9050);
nor U10704 (N_10704,N_9349,N_9544);
and U10705 (N_10705,N_9283,N_9681);
nor U10706 (N_10706,N_9835,N_9135);
and U10707 (N_10707,N_9384,N_9074);
nand U10708 (N_10708,N_9869,N_9904);
or U10709 (N_10709,N_9383,N_9480);
nand U10710 (N_10710,N_9774,N_9018);
nor U10711 (N_10711,N_9650,N_9561);
and U10712 (N_10712,N_9260,N_9252);
and U10713 (N_10713,N_9260,N_9026);
nand U10714 (N_10714,N_9052,N_9992);
and U10715 (N_10715,N_9702,N_9385);
xor U10716 (N_10716,N_9694,N_9781);
and U10717 (N_10717,N_9709,N_9126);
nand U10718 (N_10718,N_9235,N_9392);
nand U10719 (N_10719,N_9193,N_9254);
nand U10720 (N_10720,N_9493,N_9691);
nor U10721 (N_10721,N_9144,N_9947);
xor U10722 (N_10722,N_9556,N_9170);
nand U10723 (N_10723,N_9702,N_9780);
nor U10724 (N_10724,N_9783,N_9576);
nor U10725 (N_10725,N_9674,N_9128);
and U10726 (N_10726,N_9870,N_9869);
nand U10727 (N_10727,N_9851,N_9229);
or U10728 (N_10728,N_9968,N_9574);
nor U10729 (N_10729,N_9752,N_9316);
nand U10730 (N_10730,N_9503,N_9937);
or U10731 (N_10731,N_9661,N_9495);
and U10732 (N_10732,N_9872,N_9803);
nand U10733 (N_10733,N_9400,N_9070);
and U10734 (N_10734,N_9935,N_9478);
and U10735 (N_10735,N_9658,N_9060);
nand U10736 (N_10736,N_9095,N_9298);
or U10737 (N_10737,N_9372,N_9868);
nor U10738 (N_10738,N_9625,N_9365);
and U10739 (N_10739,N_9017,N_9145);
or U10740 (N_10740,N_9510,N_9856);
nor U10741 (N_10741,N_9000,N_9408);
nand U10742 (N_10742,N_9077,N_9992);
nor U10743 (N_10743,N_9930,N_9557);
nor U10744 (N_10744,N_9125,N_9726);
nor U10745 (N_10745,N_9014,N_9618);
nand U10746 (N_10746,N_9381,N_9758);
or U10747 (N_10747,N_9814,N_9121);
and U10748 (N_10748,N_9992,N_9347);
or U10749 (N_10749,N_9053,N_9925);
xor U10750 (N_10750,N_9562,N_9078);
nor U10751 (N_10751,N_9203,N_9947);
nor U10752 (N_10752,N_9253,N_9387);
and U10753 (N_10753,N_9252,N_9223);
nor U10754 (N_10754,N_9726,N_9910);
nand U10755 (N_10755,N_9601,N_9537);
and U10756 (N_10756,N_9908,N_9958);
or U10757 (N_10757,N_9695,N_9648);
nor U10758 (N_10758,N_9250,N_9116);
or U10759 (N_10759,N_9391,N_9162);
and U10760 (N_10760,N_9762,N_9501);
nor U10761 (N_10761,N_9880,N_9957);
nor U10762 (N_10762,N_9902,N_9656);
and U10763 (N_10763,N_9384,N_9856);
or U10764 (N_10764,N_9318,N_9404);
nand U10765 (N_10765,N_9027,N_9075);
nand U10766 (N_10766,N_9646,N_9612);
nor U10767 (N_10767,N_9383,N_9223);
or U10768 (N_10768,N_9549,N_9257);
and U10769 (N_10769,N_9260,N_9553);
nand U10770 (N_10770,N_9448,N_9125);
nand U10771 (N_10771,N_9437,N_9810);
nand U10772 (N_10772,N_9429,N_9194);
nor U10773 (N_10773,N_9875,N_9793);
nor U10774 (N_10774,N_9446,N_9843);
and U10775 (N_10775,N_9422,N_9412);
and U10776 (N_10776,N_9365,N_9363);
xor U10777 (N_10777,N_9758,N_9692);
or U10778 (N_10778,N_9354,N_9236);
or U10779 (N_10779,N_9985,N_9551);
and U10780 (N_10780,N_9139,N_9702);
nor U10781 (N_10781,N_9302,N_9008);
or U10782 (N_10782,N_9079,N_9478);
nand U10783 (N_10783,N_9657,N_9208);
nor U10784 (N_10784,N_9467,N_9649);
xor U10785 (N_10785,N_9610,N_9280);
nor U10786 (N_10786,N_9746,N_9203);
or U10787 (N_10787,N_9107,N_9923);
nor U10788 (N_10788,N_9777,N_9872);
and U10789 (N_10789,N_9781,N_9208);
nor U10790 (N_10790,N_9697,N_9602);
or U10791 (N_10791,N_9991,N_9674);
and U10792 (N_10792,N_9702,N_9029);
or U10793 (N_10793,N_9482,N_9102);
or U10794 (N_10794,N_9253,N_9478);
and U10795 (N_10795,N_9011,N_9546);
nor U10796 (N_10796,N_9894,N_9489);
or U10797 (N_10797,N_9696,N_9875);
nor U10798 (N_10798,N_9005,N_9575);
nor U10799 (N_10799,N_9968,N_9666);
and U10800 (N_10800,N_9644,N_9672);
and U10801 (N_10801,N_9490,N_9505);
or U10802 (N_10802,N_9379,N_9601);
or U10803 (N_10803,N_9380,N_9454);
and U10804 (N_10804,N_9583,N_9687);
nand U10805 (N_10805,N_9865,N_9197);
xnor U10806 (N_10806,N_9592,N_9310);
nor U10807 (N_10807,N_9858,N_9615);
nand U10808 (N_10808,N_9659,N_9597);
or U10809 (N_10809,N_9373,N_9372);
nand U10810 (N_10810,N_9097,N_9901);
or U10811 (N_10811,N_9740,N_9275);
nor U10812 (N_10812,N_9911,N_9153);
nand U10813 (N_10813,N_9268,N_9046);
xnor U10814 (N_10814,N_9147,N_9117);
or U10815 (N_10815,N_9310,N_9121);
or U10816 (N_10816,N_9910,N_9237);
nand U10817 (N_10817,N_9120,N_9684);
nor U10818 (N_10818,N_9638,N_9016);
nand U10819 (N_10819,N_9681,N_9719);
and U10820 (N_10820,N_9582,N_9021);
nor U10821 (N_10821,N_9522,N_9015);
nor U10822 (N_10822,N_9726,N_9192);
and U10823 (N_10823,N_9783,N_9543);
or U10824 (N_10824,N_9084,N_9191);
xnor U10825 (N_10825,N_9415,N_9958);
nor U10826 (N_10826,N_9907,N_9580);
nand U10827 (N_10827,N_9089,N_9968);
and U10828 (N_10828,N_9842,N_9403);
or U10829 (N_10829,N_9103,N_9380);
or U10830 (N_10830,N_9797,N_9153);
nand U10831 (N_10831,N_9149,N_9064);
xor U10832 (N_10832,N_9802,N_9498);
and U10833 (N_10833,N_9950,N_9219);
xnor U10834 (N_10834,N_9399,N_9117);
and U10835 (N_10835,N_9941,N_9310);
nand U10836 (N_10836,N_9604,N_9135);
and U10837 (N_10837,N_9875,N_9857);
or U10838 (N_10838,N_9382,N_9092);
and U10839 (N_10839,N_9866,N_9089);
nor U10840 (N_10840,N_9310,N_9042);
nor U10841 (N_10841,N_9563,N_9669);
nand U10842 (N_10842,N_9267,N_9493);
and U10843 (N_10843,N_9087,N_9604);
and U10844 (N_10844,N_9325,N_9546);
nor U10845 (N_10845,N_9525,N_9843);
nand U10846 (N_10846,N_9659,N_9777);
xnor U10847 (N_10847,N_9715,N_9243);
and U10848 (N_10848,N_9155,N_9622);
nor U10849 (N_10849,N_9442,N_9633);
nor U10850 (N_10850,N_9217,N_9564);
or U10851 (N_10851,N_9616,N_9407);
and U10852 (N_10852,N_9347,N_9650);
or U10853 (N_10853,N_9493,N_9879);
nand U10854 (N_10854,N_9370,N_9621);
nand U10855 (N_10855,N_9160,N_9821);
nand U10856 (N_10856,N_9440,N_9560);
nor U10857 (N_10857,N_9346,N_9568);
or U10858 (N_10858,N_9399,N_9261);
nand U10859 (N_10859,N_9144,N_9911);
nand U10860 (N_10860,N_9493,N_9211);
and U10861 (N_10861,N_9122,N_9073);
nor U10862 (N_10862,N_9918,N_9115);
nand U10863 (N_10863,N_9933,N_9235);
nand U10864 (N_10864,N_9519,N_9289);
or U10865 (N_10865,N_9350,N_9732);
or U10866 (N_10866,N_9535,N_9810);
nand U10867 (N_10867,N_9433,N_9948);
and U10868 (N_10868,N_9575,N_9063);
nand U10869 (N_10869,N_9054,N_9076);
xor U10870 (N_10870,N_9783,N_9615);
or U10871 (N_10871,N_9699,N_9149);
nor U10872 (N_10872,N_9133,N_9117);
nor U10873 (N_10873,N_9278,N_9511);
and U10874 (N_10874,N_9909,N_9361);
xnor U10875 (N_10875,N_9884,N_9480);
and U10876 (N_10876,N_9991,N_9744);
or U10877 (N_10877,N_9081,N_9141);
nand U10878 (N_10878,N_9953,N_9261);
and U10879 (N_10879,N_9139,N_9203);
and U10880 (N_10880,N_9395,N_9847);
nor U10881 (N_10881,N_9554,N_9703);
and U10882 (N_10882,N_9056,N_9122);
or U10883 (N_10883,N_9120,N_9499);
nor U10884 (N_10884,N_9903,N_9316);
and U10885 (N_10885,N_9162,N_9479);
nand U10886 (N_10886,N_9150,N_9342);
nor U10887 (N_10887,N_9647,N_9680);
and U10888 (N_10888,N_9076,N_9929);
or U10889 (N_10889,N_9564,N_9097);
nand U10890 (N_10890,N_9151,N_9784);
and U10891 (N_10891,N_9746,N_9971);
xor U10892 (N_10892,N_9851,N_9679);
nor U10893 (N_10893,N_9554,N_9923);
or U10894 (N_10894,N_9094,N_9630);
xor U10895 (N_10895,N_9958,N_9023);
nand U10896 (N_10896,N_9716,N_9830);
or U10897 (N_10897,N_9170,N_9466);
or U10898 (N_10898,N_9486,N_9609);
or U10899 (N_10899,N_9870,N_9300);
nor U10900 (N_10900,N_9481,N_9713);
and U10901 (N_10901,N_9070,N_9149);
nor U10902 (N_10902,N_9465,N_9600);
or U10903 (N_10903,N_9329,N_9100);
and U10904 (N_10904,N_9825,N_9031);
and U10905 (N_10905,N_9042,N_9485);
and U10906 (N_10906,N_9101,N_9431);
and U10907 (N_10907,N_9467,N_9958);
or U10908 (N_10908,N_9225,N_9530);
nand U10909 (N_10909,N_9704,N_9215);
or U10910 (N_10910,N_9958,N_9954);
nor U10911 (N_10911,N_9889,N_9066);
or U10912 (N_10912,N_9767,N_9321);
or U10913 (N_10913,N_9361,N_9118);
and U10914 (N_10914,N_9106,N_9396);
and U10915 (N_10915,N_9219,N_9235);
nand U10916 (N_10916,N_9092,N_9625);
nor U10917 (N_10917,N_9303,N_9978);
or U10918 (N_10918,N_9919,N_9641);
nand U10919 (N_10919,N_9606,N_9029);
nand U10920 (N_10920,N_9280,N_9713);
nand U10921 (N_10921,N_9849,N_9314);
nand U10922 (N_10922,N_9120,N_9384);
nand U10923 (N_10923,N_9850,N_9138);
or U10924 (N_10924,N_9012,N_9323);
and U10925 (N_10925,N_9605,N_9826);
and U10926 (N_10926,N_9498,N_9609);
nand U10927 (N_10927,N_9076,N_9042);
nand U10928 (N_10928,N_9269,N_9296);
nand U10929 (N_10929,N_9236,N_9152);
and U10930 (N_10930,N_9769,N_9513);
nand U10931 (N_10931,N_9525,N_9106);
nand U10932 (N_10932,N_9536,N_9112);
xor U10933 (N_10933,N_9105,N_9973);
nand U10934 (N_10934,N_9093,N_9246);
nand U10935 (N_10935,N_9045,N_9731);
or U10936 (N_10936,N_9427,N_9636);
xnor U10937 (N_10937,N_9745,N_9914);
and U10938 (N_10938,N_9573,N_9021);
nand U10939 (N_10939,N_9224,N_9473);
nor U10940 (N_10940,N_9087,N_9575);
nor U10941 (N_10941,N_9697,N_9123);
or U10942 (N_10942,N_9044,N_9496);
or U10943 (N_10943,N_9038,N_9094);
or U10944 (N_10944,N_9293,N_9848);
or U10945 (N_10945,N_9306,N_9398);
nor U10946 (N_10946,N_9292,N_9102);
nand U10947 (N_10947,N_9062,N_9087);
xnor U10948 (N_10948,N_9373,N_9483);
nor U10949 (N_10949,N_9459,N_9980);
and U10950 (N_10950,N_9559,N_9265);
nand U10951 (N_10951,N_9104,N_9545);
or U10952 (N_10952,N_9990,N_9862);
or U10953 (N_10953,N_9454,N_9398);
nand U10954 (N_10954,N_9288,N_9882);
nor U10955 (N_10955,N_9849,N_9239);
and U10956 (N_10956,N_9137,N_9139);
nand U10957 (N_10957,N_9950,N_9747);
nand U10958 (N_10958,N_9475,N_9649);
nor U10959 (N_10959,N_9378,N_9342);
or U10960 (N_10960,N_9471,N_9862);
xnor U10961 (N_10961,N_9116,N_9375);
or U10962 (N_10962,N_9720,N_9858);
or U10963 (N_10963,N_9119,N_9574);
nand U10964 (N_10964,N_9477,N_9706);
nor U10965 (N_10965,N_9489,N_9779);
nand U10966 (N_10966,N_9142,N_9348);
xor U10967 (N_10967,N_9593,N_9988);
and U10968 (N_10968,N_9830,N_9194);
nand U10969 (N_10969,N_9705,N_9816);
nand U10970 (N_10970,N_9510,N_9017);
xnor U10971 (N_10971,N_9194,N_9708);
nand U10972 (N_10972,N_9478,N_9522);
nor U10973 (N_10973,N_9385,N_9072);
and U10974 (N_10974,N_9729,N_9746);
and U10975 (N_10975,N_9972,N_9847);
or U10976 (N_10976,N_9933,N_9741);
nor U10977 (N_10977,N_9158,N_9824);
or U10978 (N_10978,N_9238,N_9778);
or U10979 (N_10979,N_9894,N_9585);
nand U10980 (N_10980,N_9828,N_9224);
or U10981 (N_10981,N_9298,N_9213);
and U10982 (N_10982,N_9140,N_9514);
nand U10983 (N_10983,N_9512,N_9436);
or U10984 (N_10984,N_9778,N_9941);
nand U10985 (N_10985,N_9425,N_9587);
nor U10986 (N_10986,N_9442,N_9573);
nand U10987 (N_10987,N_9923,N_9523);
and U10988 (N_10988,N_9939,N_9092);
and U10989 (N_10989,N_9992,N_9815);
nand U10990 (N_10990,N_9754,N_9448);
nand U10991 (N_10991,N_9367,N_9228);
nand U10992 (N_10992,N_9116,N_9050);
xnor U10993 (N_10993,N_9240,N_9244);
or U10994 (N_10994,N_9409,N_9045);
or U10995 (N_10995,N_9226,N_9821);
nand U10996 (N_10996,N_9697,N_9945);
nor U10997 (N_10997,N_9579,N_9429);
nand U10998 (N_10998,N_9201,N_9848);
or U10999 (N_10999,N_9849,N_9548);
or U11000 (N_11000,N_10571,N_10783);
nor U11001 (N_11001,N_10090,N_10251);
nor U11002 (N_11002,N_10607,N_10905);
nand U11003 (N_11003,N_10636,N_10020);
nand U11004 (N_11004,N_10363,N_10511);
and U11005 (N_11005,N_10445,N_10823);
nand U11006 (N_11006,N_10854,N_10214);
xor U11007 (N_11007,N_10052,N_10894);
and U11008 (N_11008,N_10631,N_10004);
and U11009 (N_11009,N_10129,N_10520);
nor U11010 (N_11010,N_10717,N_10486);
nand U11011 (N_11011,N_10911,N_10827);
and U11012 (N_11012,N_10016,N_10040);
nand U11013 (N_11013,N_10076,N_10992);
xor U11014 (N_11014,N_10710,N_10546);
xnor U11015 (N_11015,N_10628,N_10950);
and U11016 (N_11016,N_10712,N_10061);
nand U11017 (N_11017,N_10149,N_10860);
or U11018 (N_11018,N_10741,N_10617);
nor U11019 (N_11019,N_10037,N_10064);
xor U11020 (N_11020,N_10472,N_10421);
or U11021 (N_11021,N_10752,N_10643);
or U11022 (N_11022,N_10248,N_10570);
nand U11023 (N_11023,N_10838,N_10082);
nand U11024 (N_11024,N_10857,N_10085);
xor U11025 (N_11025,N_10097,N_10024);
xnor U11026 (N_11026,N_10612,N_10260);
nand U11027 (N_11027,N_10518,N_10945);
or U11028 (N_11028,N_10389,N_10941);
nand U11029 (N_11029,N_10733,N_10918);
or U11030 (N_11030,N_10545,N_10808);
nor U11031 (N_11031,N_10556,N_10604);
and U11032 (N_11032,N_10044,N_10409);
nand U11033 (N_11033,N_10953,N_10167);
and U11034 (N_11034,N_10596,N_10405);
nor U11035 (N_11035,N_10746,N_10831);
or U11036 (N_11036,N_10873,N_10909);
nor U11037 (N_11037,N_10448,N_10530);
xnor U11038 (N_11038,N_10263,N_10947);
and U11039 (N_11039,N_10275,N_10753);
xnor U11040 (N_11040,N_10849,N_10364);
nand U11041 (N_11041,N_10858,N_10328);
and U11042 (N_11042,N_10122,N_10246);
nand U11043 (N_11043,N_10458,N_10975);
nand U11044 (N_11044,N_10738,N_10960);
nand U11045 (N_11045,N_10152,N_10428);
or U11046 (N_11046,N_10406,N_10946);
xnor U11047 (N_11047,N_10295,N_10692);
nand U11048 (N_11048,N_10681,N_10308);
xnor U11049 (N_11049,N_10540,N_10666);
or U11050 (N_11050,N_10079,N_10142);
nor U11051 (N_11051,N_10730,N_10893);
nor U11052 (N_11052,N_10469,N_10983);
nand U11053 (N_11053,N_10656,N_10749);
and U11054 (N_11054,N_10886,N_10713);
xor U11055 (N_11055,N_10492,N_10525);
nand U11056 (N_11056,N_10991,N_10771);
and U11057 (N_11057,N_10460,N_10514);
xor U11058 (N_11058,N_10550,N_10025);
nand U11059 (N_11059,N_10735,N_10228);
nor U11060 (N_11060,N_10819,N_10537);
nor U11061 (N_11061,N_10900,N_10826);
nand U11062 (N_11062,N_10270,N_10553);
nand U11063 (N_11063,N_10673,N_10637);
nor U11064 (N_11064,N_10668,N_10578);
nor U11065 (N_11065,N_10046,N_10990);
and U11066 (N_11066,N_10128,N_10772);
and U11067 (N_11067,N_10199,N_10386);
or U11068 (N_11068,N_10255,N_10832);
or U11069 (N_11069,N_10362,N_10528);
nand U11070 (N_11070,N_10923,N_10850);
and U11071 (N_11071,N_10474,N_10473);
xor U11072 (N_11072,N_10567,N_10848);
nor U11073 (N_11073,N_10249,N_10341);
nand U11074 (N_11074,N_10307,N_10536);
nand U11075 (N_11075,N_10592,N_10906);
or U11076 (N_11076,N_10840,N_10930);
or U11077 (N_11077,N_10573,N_10459);
nand U11078 (N_11078,N_10433,N_10060);
or U11079 (N_11079,N_10081,N_10172);
xnor U11080 (N_11080,N_10332,N_10695);
and U11081 (N_11081,N_10729,N_10069);
nand U11082 (N_11082,N_10683,N_10679);
nand U11083 (N_11083,N_10271,N_10449);
and U11084 (N_11084,N_10215,N_10714);
nor U11085 (N_11085,N_10324,N_10676);
or U11086 (N_11086,N_10359,N_10117);
or U11087 (N_11087,N_10088,N_10696);
and U11088 (N_11088,N_10303,N_10345);
nor U11089 (N_11089,N_10429,N_10340);
nor U11090 (N_11090,N_10030,N_10611);
nor U11091 (N_11091,N_10635,N_10851);
nor U11092 (N_11092,N_10613,N_10532);
nand U11093 (N_11093,N_10670,N_10555);
nor U11094 (N_11094,N_10739,N_10073);
and U11095 (N_11095,N_10132,N_10552);
nor U11096 (N_11096,N_10484,N_10391);
nor U11097 (N_11097,N_10407,N_10410);
nor U11098 (N_11098,N_10927,N_10560);
and U11099 (N_11099,N_10885,N_10856);
xnor U11100 (N_11100,N_10426,N_10551);
nand U11101 (N_11101,N_10820,N_10365);
xor U11102 (N_11102,N_10222,N_10865);
xnor U11103 (N_11103,N_10863,N_10963);
and U11104 (N_11104,N_10059,N_10720);
nor U11105 (N_11105,N_10579,N_10043);
nor U11106 (N_11106,N_10479,N_10456);
or U11107 (N_11107,N_10284,N_10057);
or U11108 (N_11108,N_10661,N_10910);
or U11109 (N_11109,N_10745,N_10161);
nand U11110 (N_11110,N_10427,N_10357);
nor U11111 (N_11111,N_10504,N_10987);
nand U11112 (N_11112,N_10701,N_10381);
and U11113 (N_11113,N_10166,N_10790);
nor U11114 (N_11114,N_10541,N_10399);
and U11115 (N_11115,N_10119,N_10707);
nand U11116 (N_11116,N_10675,N_10318);
nand U11117 (N_11117,N_10182,N_10881);
and U11118 (N_11118,N_10224,N_10903);
or U11119 (N_11119,N_10134,N_10033);
or U11120 (N_11120,N_10976,N_10217);
nor U11121 (N_11121,N_10252,N_10022);
nand U11122 (N_11122,N_10743,N_10339);
nand U11123 (N_11123,N_10141,N_10056);
xnor U11124 (N_11124,N_10915,N_10159);
nand U11125 (N_11125,N_10188,N_10121);
nor U11126 (N_11126,N_10765,N_10958);
and U11127 (N_11127,N_10093,N_10964);
nand U11128 (N_11128,N_10192,N_10795);
nor U11129 (N_11129,N_10277,N_10967);
nor U11130 (N_11130,N_10653,N_10180);
or U11131 (N_11131,N_10503,N_10736);
nand U11132 (N_11132,N_10115,N_10299);
and U11133 (N_11133,N_10387,N_10205);
nand U11134 (N_11134,N_10400,N_10603);
or U11135 (N_11135,N_10273,N_10286);
and U11136 (N_11136,N_10379,N_10652);
or U11137 (N_11137,N_10118,N_10092);
or U11138 (N_11138,N_10225,N_10558);
nand U11139 (N_11139,N_10747,N_10276);
xnor U11140 (N_11140,N_10825,N_10583);
and U11141 (N_11141,N_10241,N_10305);
nand U11142 (N_11142,N_10651,N_10414);
xnor U11143 (N_11143,N_10220,N_10727);
nand U11144 (N_11144,N_10574,N_10706);
and U11145 (N_11145,N_10780,N_10822);
xnor U11146 (N_11146,N_10042,N_10138);
and U11147 (N_11147,N_10306,N_10094);
nor U11148 (N_11148,N_10023,N_10366);
nor U11149 (N_11149,N_10351,N_10053);
nand U11150 (N_11150,N_10792,N_10902);
or U11151 (N_11151,N_10105,N_10360);
nor U11152 (N_11152,N_10791,N_10066);
nor U11153 (N_11153,N_10853,N_10144);
nor U11154 (N_11154,N_10561,N_10794);
or U11155 (N_11155,N_10098,N_10843);
and U11156 (N_11156,N_10658,N_10928);
xor U11157 (N_11157,N_10678,N_10181);
or U11158 (N_11158,N_10354,N_10232);
xor U11159 (N_11159,N_10793,N_10424);
and U11160 (N_11160,N_10936,N_10281);
nor U11161 (N_11161,N_10431,N_10810);
or U11162 (N_11162,N_10507,N_10148);
nand U11163 (N_11163,N_10493,N_10078);
or U11164 (N_11164,N_10187,N_10879);
or U11165 (N_11165,N_10471,N_10883);
nor U11166 (N_11166,N_10803,N_10644);
and U11167 (N_11167,N_10750,N_10002);
or U11168 (N_11168,N_10123,N_10602);
nand U11169 (N_11169,N_10801,N_10837);
nor U11170 (N_11170,N_10971,N_10029);
or U11171 (N_11171,N_10719,N_10355);
nor U11172 (N_11172,N_10347,N_10087);
nand U11173 (N_11173,N_10660,N_10589);
and U11174 (N_11174,N_10338,N_10477);
and U11175 (N_11175,N_10145,N_10380);
or U11176 (N_11176,N_10096,N_10461);
and U11177 (N_11177,N_10333,N_10648);
nand U11178 (N_11178,N_10895,N_10403);
nor U11179 (N_11179,N_10777,N_10268);
or U11180 (N_11180,N_10995,N_10012);
nor U11181 (N_11181,N_10321,N_10642);
and U11182 (N_11182,N_10049,N_10799);
nor U11183 (N_11183,N_10715,N_10375);
nand U11184 (N_11184,N_10422,N_10845);
nor U11185 (N_11185,N_10210,N_10008);
nand U11186 (N_11186,N_10147,N_10665);
or U11187 (N_11187,N_10256,N_10349);
xnor U11188 (N_11188,N_10155,N_10979);
or U11189 (N_11189,N_10265,N_10898);
xor U11190 (N_11190,N_10314,N_10104);
nor U11191 (N_11191,N_10266,N_10582);
nor U11192 (N_11192,N_10892,N_10154);
and U11193 (N_11193,N_10075,N_10973);
or U11194 (N_11194,N_10954,N_10417);
nor U11195 (N_11195,N_10113,N_10526);
nor U11196 (N_11196,N_10758,N_10505);
and U11197 (N_11197,N_10168,N_10356);
xor U11198 (N_11198,N_10133,N_10430);
and U11199 (N_11199,N_10291,N_10319);
nand U11200 (N_11200,N_10352,N_10289);
nor U11201 (N_11201,N_10705,N_10773);
or U11202 (N_11202,N_10208,N_10213);
and U11203 (N_11203,N_10184,N_10462);
nand U11204 (N_11204,N_10005,N_10419);
and U11205 (N_11205,N_10544,N_10183);
or U11206 (N_11206,N_10259,N_10331);
nand U11207 (N_11207,N_10988,N_10709);
xnor U11208 (N_11208,N_10982,N_10301);
nand U11209 (N_11209,N_10382,N_10968);
xnor U11210 (N_11210,N_10444,N_10640);
xnor U11211 (N_11211,N_10869,N_10485);
nor U11212 (N_11212,N_10564,N_10438);
nand U11213 (N_11213,N_10841,N_10726);
and U11214 (N_11214,N_10922,N_10302);
nand U11215 (N_11215,N_10818,N_10487);
or U11216 (N_11216,N_10209,N_10369);
and U11217 (N_11217,N_10500,N_10674);
nand U11218 (N_11218,N_10948,N_10805);
and U11219 (N_11219,N_10370,N_10377);
nor U11220 (N_11220,N_10938,N_10102);
xnor U11221 (N_11221,N_10616,N_10998);
or U11222 (N_11222,N_10871,N_10385);
or U11223 (N_11223,N_10236,N_10813);
nor U11224 (N_11224,N_10164,N_10027);
nand U11225 (N_11225,N_10880,N_10189);
nand U11226 (N_11226,N_10659,N_10390);
nand U11227 (N_11227,N_10839,N_10916);
xor U11228 (N_11228,N_10939,N_10358);
and U11229 (N_11229,N_10348,N_10921);
and U11230 (N_11230,N_10581,N_10663);
or U11231 (N_11231,N_10908,N_10283);
xnor U11232 (N_11232,N_10623,N_10598);
nor U11233 (N_11233,N_10562,N_10684);
nor U11234 (N_11234,N_10874,N_10760);
or U11235 (N_11235,N_10396,N_10697);
nor U11236 (N_11236,N_10501,N_10408);
nand U11237 (N_11237,N_10196,N_10535);
nor U11238 (N_11238,N_10383,N_10548);
xor U11239 (N_11239,N_10935,N_10566);
or U11240 (N_11240,N_10021,N_10453);
nand U11241 (N_11241,N_10048,N_10436);
nand U11242 (N_11242,N_10542,N_10361);
nand U11243 (N_11243,N_10957,N_10420);
xnor U11244 (N_11244,N_10388,N_10326);
xor U11245 (N_11245,N_10577,N_10650);
nand U11246 (N_11246,N_10211,N_10816);
nor U11247 (N_11247,N_10914,N_10212);
or U11248 (N_11248,N_10036,N_10506);
or U11249 (N_11249,N_10242,N_10517);
and U11250 (N_11250,N_10101,N_10330);
and U11251 (N_11251,N_10404,N_10169);
and U11252 (N_11252,N_10455,N_10051);
nor U11253 (N_11253,N_10722,N_10143);
xor U11254 (N_11254,N_10931,N_10494);
xor U11255 (N_11255,N_10654,N_10480);
nor U11256 (N_11256,N_10015,N_10071);
nand U11257 (N_11257,N_10074,N_10335);
nand U11258 (N_11258,N_10748,N_10063);
nor U11259 (N_11259,N_10787,N_10201);
and U11260 (N_11260,N_10605,N_10907);
xnor U11261 (N_11261,N_10185,N_10533);
nand U11262 (N_11262,N_10139,N_10467);
xor U11263 (N_11263,N_10757,N_10929);
nor U11264 (N_11264,N_10434,N_10543);
and U11265 (N_11265,N_10206,N_10751);
nand U11266 (N_11266,N_10110,N_10243);
or U11267 (N_11267,N_10646,N_10944);
nor U11268 (N_11268,N_10776,N_10350);
and U11269 (N_11269,N_10600,N_10084);
nor U11270 (N_11270,N_10759,N_10667);
nand U11271 (N_11271,N_10797,N_10267);
nor U11272 (N_11272,N_10465,N_10896);
and U11273 (N_11273,N_10413,N_10647);
or U11274 (N_11274,N_10013,N_10688);
or U11275 (N_11275,N_10497,N_10884);
and U11276 (N_11276,N_10786,N_10219);
xnor U11277 (N_11277,N_10834,N_10320);
nor U11278 (N_11278,N_10498,N_10997);
nor U11279 (N_11279,N_10584,N_10641);
nor U11280 (N_11280,N_10913,N_10398);
and U11281 (N_11281,N_10112,N_10077);
or U11282 (N_11282,N_10293,N_10107);
or U11283 (N_11283,N_10828,N_10124);
or U11284 (N_11284,N_10942,N_10146);
and U11285 (N_11285,N_10933,N_10313);
nand U11286 (N_11286,N_10346,N_10014);
nor U11287 (N_11287,N_10239,N_10156);
or U11288 (N_11288,N_10952,N_10620);
nand U11289 (N_11289,N_10502,N_10711);
nor U11290 (N_11290,N_10019,N_10416);
nor U11291 (N_11291,N_10626,N_10523);
nand U11292 (N_11292,N_10315,N_10230);
or U11293 (N_11293,N_10890,N_10833);
or U11294 (N_11294,N_10778,N_10280);
or U11295 (N_11295,N_10200,N_10068);
or U11296 (N_11296,N_10519,N_10153);
or U11297 (N_11297,N_10585,N_10789);
xor U11298 (N_11298,N_10130,N_10703);
nor U11299 (N_11299,N_10179,N_10374);
or U11300 (N_11300,N_10039,N_10586);
nand U11301 (N_11301,N_10859,N_10924);
or U11302 (N_11302,N_10755,N_10258);
and U11303 (N_11303,N_10993,N_10394);
or U11304 (N_11304,N_10026,N_10980);
xor U11305 (N_11305,N_10999,N_10830);
and U11306 (N_11306,N_10116,N_10547);
or U11307 (N_11307,N_10452,N_10691);
nor U11308 (N_11308,N_10767,N_10136);
nor U11309 (N_11309,N_10238,N_10468);
nor U11310 (N_11310,N_10708,N_10806);
nor U11311 (N_11311,N_10297,N_10089);
nand U11312 (N_11312,N_10889,N_10619);
and U11313 (N_11313,N_10296,N_10870);
nand U11314 (N_11314,N_10186,N_10244);
and U11315 (N_11315,N_10887,N_10601);
nand U11316 (N_11316,N_10300,N_10231);
xnor U11317 (N_11317,N_10698,N_10512);
nor U11318 (N_11318,N_10058,N_10510);
or U11319 (N_11319,N_10001,N_10899);
and U11320 (N_11320,N_10981,N_10978);
or U11321 (N_11321,N_10229,N_10111);
nand U11322 (N_11322,N_10234,N_10091);
nor U11323 (N_11323,N_10011,N_10557);
or U11324 (N_11324,N_10443,N_10513);
or U11325 (N_11325,N_10731,N_10784);
nor U11326 (N_11326,N_10316,N_10233);
and U11327 (N_11327,N_10996,N_10344);
or U11328 (N_11328,N_10203,N_10534);
nor U11329 (N_11329,N_10974,N_10694);
and U11330 (N_11330,N_10262,N_10815);
or U11331 (N_11331,N_10618,N_10312);
or U11332 (N_11332,N_10401,N_10744);
nor U11333 (N_11333,N_10614,N_10590);
and U11334 (N_11334,N_10861,N_10934);
or U11335 (N_11335,N_10687,N_10835);
nand U11336 (N_11336,N_10041,N_10131);
nand U11337 (N_11337,N_10264,N_10664);
nor U11338 (N_11338,N_10086,N_10272);
and U11339 (N_11339,N_10446,N_10812);
and U11340 (N_11340,N_10395,N_10309);
nor U11341 (N_11341,N_10955,N_10050);
nand U11342 (N_11342,N_10864,N_10926);
nand U11343 (N_11343,N_10877,N_10202);
or U11344 (N_11344,N_10904,N_10699);
nand U11345 (N_11345,N_10028,N_10633);
nand U11346 (N_11346,N_10095,N_10689);
xnor U11347 (N_11347,N_10031,N_10768);
xnor U11348 (N_11348,N_10221,N_10782);
and U11349 (N_11349,N_10677,N_10829);
nand U11350 (N_11350,N_10919,N_10163);
or U11351 (N_11351,N_10476,N_10655);
nor U11352 (N_11352,N_10972,N_10207);
and U11353 (N_11353,N_10065,N_10943);
and U11354 (N_11354,N_10000,N_10754);
nand U11355 (N_11355,N_10171,N_10007);
nand U11356 (N_11356,N_10178,N_10055);
or U11357 (N_11357,N_10017,N_10606);
nand U11358 (N_11358,N_10304,N_10742);
xor U11359 (N_11359,N_10464,N_10126);
nand U11360 (N_11360,N_10878,N_10559);
xor U11361 (N_11361,N_10191,N_10716);
or U11362 (N_11362,N_10959,N_10287);
and U11363 (N_11363,N_10488,N_10317);
or U11364 (N_11364,N_10470,N_10624);
and U11365 (N_11365,N_10940,N_10531);
or U11366 (N_11366,N_10872,N_10140);
or U11367 (N_11367,N_10593,N_10175);
or U11368 (N_11368,N_10568,N_10588);
or U11369 (N_11369,N_10282,N_10176);
and U11370 (N_11370,N_10437,N_10435);
nor U11371 (N_11371,N_10956,N_10006);
nand U11372 (N_11372,N_10100,N_10466);
and U11373 (N_11373,N_10587,N_10327);
nand U11374 (N_11374,N_10932,N_10725);
nor U11375 (N_11375,N_10965,N_10595);
or U11376 (N_11376,N_10285,N_10591);
and U11377 (N_11377,N_10962,N_10227);
and U11378 (N_11378,N_10240,N_10250);
or U11379 (N_11379,N_10322,N_10852);
or U11380 (N_11380,N_10693,N_10257);
nor U11381 (N_11381,N_10925,N_10127);
nor U11382 (N_11382,N_10197,N_10496);
and U11383 (N_11383,N_10190,N_10237);
nand U11384 (N_11384,N_10384,N_10412);
and U11385 (N_11385,N_10682,N_10451);
nand U11386 (N_11386,N_10969,N_10554);
nand U11387 (N_11387,N_10868,N_10245);
or U11388 (N_11388,N_10376,N_10432);
nand U11389 (N_11389,N_10495,N_10261);
and U11390 (N_11390,N_10855,N_10732);
nand U11391 (N_11391,N_10441,N_10294);
nor U11392 (N_11392,N_10195,N_10522);
and U11393 (N_11393,N_10690,N_10108);
nand U11394 (N_11394,N_10610,N_10080);
or U11395 (N_11395,N_10157,N_10003);
or U11396 (N_11396,N_10378,N_10576);
nand U11397 (N_11397,N_10740,N_10521);
nand U11398 (N_11398,N_10489,N_10756);
nor U11399 (N_11399,N_10937,N_10762);
nor U11400 (N_11400,N_10173,N_10622);
nand U11401 (N_11401,N_10804,N_10516);
nor U11402 (N_11402,N_10917,N_10809);
nor U11403 (N_11403,N_10103,N_10846);
nor U11404 (N_11404,N_10125,N_10862);
xnor U11405 (N_11405,N_10970,N_10704);
xnor U11406 (N_11406,N_10483,N_10985);
nand U11407 (N_11407,N_10204,N_10254);
nor U11408 (N_11408,N_10669,N_10608);
or U11409 (N_11409,N_10775,N_10475);
and U11410 (N_11410,N_10572,N_10977);
and U11411 (N_11411,N_10323,N_10769);
or U11412 (N_11412,N_10625,N_10070);
nand U11413 (N_11413,N_10193,N_10034);
xnor U11414 (N_11414,N_10888,N_10515);
nand U11415 (N_11415,N_10671,N_10411);
xor U11416 (N_11416,N_10170,N_10106);
or U11417 (N_11417,N_10174,N_10649);
nand U11418 (N_11418,N_10876,N_10353);
xor U11419 (N_11419,N_10842,N_10882);
xor U11420 (N_11420,N_10539,N_10800);
nor U11421 (N_11421,N_10439,N_10529);
or U11422 (N_11422,N_10788,N_10425);
nor U11423 (N_11423,N_10770,N_10311);
and U11424 (N_11424,N_10450,N_10083);
or U11425 (N_11425,N_10912,N_10580);
nor U11426 (N_11426,N_10440,N_10866);
nor U11427 (N_11427,N_10491,N_10062);
or U11428 (N_11428,N_10986,N_10198);
nand U11429 (N_11429,N_10632,N_10290);
and U11430 (N_11430,N_10150,N_10621);
xor U11431 (N_11431,N_10627,N_10045);
and U11432 (N_11432,N_10067,N_10798);
and U11433 (N_11433,N_10645,N_10599);
nor U11434 (N_11434,N_10524,N_10018);
nand U11435 (N_11435,N_10702,N_10811);
and U11436 (N_11436,N_10718,N_10032);
or U11437 (N_11437,N_10072,N_10994);
nor U11438 (N_11438,N_10372,N_10099);
or U11439 (N_11439,N_10951,N_10274);
or U11440 (N_11440,N_10686,N_10490);
nand U11441 (N_11441,N_10035,N_10235);
nor U11442 (N_11442,N_10336,N_10672);
nand U11443 (N_11443,N_10734,N_10630);
nor U11444 (N_11444,N_10844,N_10565);
or U11445 (N_11445,N_10194,N_10785);
nand U11446 (N_11446,N_10549,N_10817);
nor U11447 (N_11447,N_10781,N_10223);
nor U11448 (N_11448,N_10278,N_10447);
or U11449 (N_11449,N_10920,N_10766);
and U11450 (N_11450,N_10310,N_10392);
xor U11451 (N_11451,N_10814,N_10764);
nand U11452 (N_11452,N_10463,N_10891);
and U11453 (N_11453,N_10478,N_10160);
and U11454 (N_11454,N_10538,N_10499);
and U11455 (N_11455,N_10508,N_10325);
or U11456 (N_11456,N_10680,N_10629);
and U11457 (N_11457,N_10373,N_10796);
nand U11458 (N_11458,N_10721,N_10454);
xor U11459 (N_11459,N_10685,N_10054);
nand U11460 (N_11460,N_10802,N_10824);
and U11461 (N_11461,N_10120,N_10821);
and U11462 (N_11462,N_10609,N_10269);
or U11463 (N_11463,N_10038,N_10763);
or U11464 (N_11464,N_10638,N_10594);
xnor U11465 (N_11465,N_10226,N_10867);
nand U11466 (N_11466,N_10009,N_10662);
nand U11467 (N_11467,N_10615,N_10457);
nand U11468 (N_11468,N_10216,N_10151);
nor U11469 (N_11469,N_10700,N_10010);
xnor U11470 (N_11470,N_10761,N_10984);
nor U11471 (N_11471,N_10334,N_10177);
and U11472 (N_11472,N_10397,N_10901);
and U11473 (N_11473,N_10897,N_10563);
xnor U11474 (N_11474,N_10288,N_10569);
and U11475 (N_11475,N_10135,N_10253);
or U11476 (N_11476,N_10218,N_10836);
xor U11477 (N_11477,N_10989,N_10137);
and U11478 (N_11478,N_10114,N_10415);
or U11479 (N_11479,N_10343,N_10737);
or U11480 (N_11480,N_10949,N_10724);
nand U11481 (N_11481,N_10527,N_10875);
nand U11482 (N_11482,N_10639,N_10442);
xor U11483 (N_11483,N_10847,N_10966);
xnor U11484 (N_11484,N_10393,N_10728);
xor U11485 (N_11485,N_10423,N_10657);
and U11486 (N_11486,N_10961,N_10402);
nor U11487 (N_11487,N_10329,N_10575);
and U11488 (N_11488,N_10158,N_10162);
nand U11489 (N_11489,N_10774,N_10279);
and U11490 (N_11490,N_10292,N_10482);
nand U11491 (N_11491,N_10509,N_10337);
or U11492 (N_11492,N_10597,N_10247);
or U11493 (N_11493,N_10807,N_10368);
or U11494 (N_11494,N_10367,N_10298);
or U11495 (N_11495,N_10109,N_10723);
nor U11496 (N_11496,N_10371,N_10418);
nand U11497 (N_11497,N_10779,N_10165);
nor U11498 (N_11498,N_10481,N_10342);
nand U11499 (N_11499,N_10047,N_10634);
or U11500 (N_11500,N_10497,N_10810);
nor U11501 (N_11501,N_10894,N_10677);
xnor U11502 (N_11502,N_10280,N_10292);
or U11503 (N_11503,N_10849,N_10089);
or U11504 (N_11504,N_10416,N_10913);
and U11505 (N_11505,N_10141,N_10038);
or U11506 (N_11506,N_10068,N_10087);
and U11507 (N_11507,N_10534,N_10303);
or U11508 (N_11508,N_10576,N_10474);
or U11509 (N_11509,N_10382,N_10405);
nand U11510 (N_11510,N_10210,N_10242);
xnor U11511 (N_11511,N_10859,N_10094);
or U11512 (N_11512,N_10951,N_10966);
nor U11513 (N_11513,N_10977,N_10266);
nand U11514 (N_11514,N_10018,N_10663);
nor U11515 (N_11515,N_10792,N_10615);
xor U11516 (N_11516,N_10686,N_10722);
nand U11517 (N_11517,N_10862,N_10847);
and U11518 (N_11518,N_10430,N_10784);
or U11519 (N_11519,N_10955,N_10627);
nand U11520 (N_11520,N_10113,N_10698);
or U11521 (N_11521,N_10674,N_10654);
xor U11522 (N_11522,N_10974,N_10221);
nor U11523 (N_11523,N_10712,N_10936);
nor U11524 (N_11524,N_10833,N_10900);
nor U11525 (N_11525,N_10041,N_10016);
nor U11526 (N_11526,N_10827,N_10627);
nand U11527 (N_11527,N_10636,N_10431);
nand U11528 (N_11528,N_10991,N_10634);
nand U11529 (N_11529,N_10465,N_10112);
nand U11530 (N_11530,N_10045,N_10461);
and U11531 (N_11531,N_10146,N_10274);
xnor U11532 (N_11532,N_10428,N_10699);
nand U11533 (N_11533,N_10849,N_10343);
nand U11534 (N_11534,N_10263,N_10514);
xor U11535 (N_11535,N_10227,N_10176);
and U11536 (N_11536,N_10008,N_10193);
nor U11537 (N_11537,N_10467,N_10208);
nor U11538 (N_11538,N_10948,N_10725);
or U11539 (N_11539,N_10514,N_10822);
and U11540 (N_11540,N_10104,N_10940);
or U11541 (N_11541,N_10214,N_10002);
and U11542 (N_11542,N_10100,N_10967);
or U11543 (N_11543,N_10503,N_10800);
and U11544 (N_11544,N_10410,N_10257);
nor U11545 (N_11545,N_10966,N_10003);
or U11546 (N_11546,N_10712,N_10607);
nor U11547 (N_11547,N_10711,N_10501);
nand U11548 (N_11548,N_10803,N_10099);
or U11549 (N_11549,N_10235,N_10620);
nand U11550 (N_11550,N_10865,N_10182);
nand U11551 (N_11551,N_10779,N_10573);
and U11552 (N_11552,N_10235,N_10086);
nor U11553 (N_11553,N_10797,N_10662);
and U11554 (N_11554,N_10392,N_10197);
xor U11555 (N_11555,N_10834,N_10152);
and U11556 (N_11556,N_10461,N_10854);
nand U11557 (N_11557,N_10958,N_10255);
or U11558 (N_11558,N_10914,N_10957);
or U11559 (N_11559,N_10960,N_10238);
and U11560 (N_11560,N_10417,N_10492);
nand U11561 (N_11561,N_10606,N_10843);
or U11562 (N_11562,N_10508,N_10835);
nand U11563 (N_11563,N_10127,N_10207);
xor U11564 (N_11564,N_10050,N_10889);
xnor U11565 (N_11565,N_10045,N_10476);
nor U11566 (N_11566,N_10616,N_10817);
or U11567 (N_11567,N_10545,N_10446);
or U11568 (N_11568,N_10390,N_10363);
nand U11569 (N_11569,N_10746,N_10335);
nor U11570 (N_11570,N_10573,N_10396);
or U11571 (N_11571,N_10834,N_10805);
nor U11572 (N_11572,N_10130,N_10085);
or U11573 (N_11573,N_10440,N_10544);
nand U11574 (N_11574,N_10399,N_10141);
nor U11575 (N_11575,N_10947,N_10780);
xnor U11576 (N_11576,N_10271,N_10771);
xor U11577 (N_11577,N_10958,N_10959);
nand U11578 (N_11578,N_10721,N_10931);
and U11579 (N_11579,N_10420,N_10687);
nand U11580 (N_11580,N_10103,N_10195);
and U11581 (N_11581,N_10693,N_10888);
nor U11582 (N_11582,N_10792,N_10562);
or U11583 (N_11583,N_10669,N_10158);
or U11584 (N_11584,N_10614,N_10837);
or U11585 (N_11585,N_10408,N_10515);
or U11586 (N_11586,N_10001,N_10240);
xnor U11587 (N_11587,N_10638,N_10465);
or U11588 (N_11588,N_10693,N_10433);
nor U11589 (N_11589,N_10893,N_10981);
and U11590 (N_11590,N_10381,N_10014);
nor U11591 (N_11591,N_10392,N_10563);
nand U11592 (N_11592,N_10214,N_10245);
and U11593 (N_11593,N_10839,N_10306);
nand U11594 (N_11594,N_10107,N_10254);
nor U11595 (N_11595,N_10105,N_10656);
nor U11596 (N_11596,N_10368,N_10766);
and U11597 (N_11597,N_10279,N_10714);
or U11598 (N_11598,N_10317,N_10919);
or U11599 (N_11599,N_10794,N_10464);
and U11600 (N_11600,N_10258,N_10118);
nor U11601 (N_11601,N_10080,N_10469);
nor U11602 (N_11602,N_10382,N_10688);
or U11603 (N_11603,N_10637,N_10854);
xor U11604 (N_11604,N_10995,N_10551);
nor U11605 (N_11605,N_10620,N_10974);
nand U11606 (N_11606,N_10068,N_10588);
nor U11607 (N_11607,N_10474,N_10396);
nor U11608 (N_11608,N_10835,N_10474);
nor U11609 (N_11609,N_10929,N_10628);
or U11610 (N_11610,N_10645,N_10590);
nand U11611 (N_11611,N_10576,N_10182);
nand U11612 (N_11612,N_10733,N_10707);
and U11613 (N_11613,N_10495,N_10225);
and U11614 (N_11614,N_10703,N_10458);
nand U11615 (N_11615,N_10548,N_10412);
or U11616 (N_11616,N_10802,N_10520);
xor U11617 (N_11617,N_10598,N_10467);
and U11618 (N_11618,N_10066,N_10830);
xnor U11619 (N_11619,N_10842,N_10256);
or U11620 (N_11620,N_10825,N_10516);
nand U11621 (N_11621,N_10628,N_10579);
nor U11622 (N_11622,N_10501,N_10780);
and U11623 (N_11623,N_10223,N_10653);
or U11624 (N_11624,N_10398,N_10493);
nor U11625 (N_11625,N_10331,N_10999);
nor U11626 (N_11626,N_10707,N_10817);
or U11627 (N_11627,N_10141,N_10446);
nand U11628 (N_11628,N_10122,N_10117);
nor U11629 (N_11629,N_10839,N_10979);
nand U11630 (N_11630,N_10233,N_10559);
xor U11631 (N_11631,N_10485,N_10038);
nor U11632 (N_11632,N_10044,N_10163);
or U11633 (N_11633,N_10110,N_10852);
xor U11634 (N_11634,N_10543,N_10020);
or U11635 (N_11635,N_10050,N_10528);
and U11636 (N_11636,N_10273,N_10195);
and U11637 (N_11637,N_10817,N_10571);
nand U11638 (N_11638,N_10521,N_10639);
nand U11639 (N_11639,N_10496,N_10678);
xor U11640 (N_11640,N_10552,N_10337);
and U11641 (N_11641,N_10585,N_10372);
nor U11642 (N_11642,N_10671,N_10549);
nor U11643 (N_11643,N_10378,N_10284);
or U11644 (N_11644,N_10780,N_10591);
xnor U11645 (N_11645,N_10347,N_10368);
nor U11646 (N_11646,N_10451,N_10019);
nand U11647 (N_11647,N_10407,N_10497);
nor U11648 (N_11648,N_10036,N_10549);
nand U11649 (N_11649,N_10099,N_10422);
nand U11650 (N_11650,N_10017,N_10752);
nand U11651 (N_11651,N_10865,N_10696);
or U11652 (N_11652,N_10486,N_10463);
and U11653 (N_11653,N_10779,N_10001);
nor U11654 (N_11654,N_10946,N_10680);
nand U11655 (N_11655,N_10483,N_10284);
and U11656 (N_11656,N_10662,N_10710);
and U11657 (N_11657,N_10121,N_10162);
and U11658 (N_11658,N_10088,N_10422);
and U11659 (N_11659,N_10194,N_10316);
and U11660 (N_11660,N_10632,N_10918);
nand U11661 (N_11661,N_10559,N_10067);
nand U11662 (N_11662,N_10990,N_10838);
or U11663 (N_11663,N_10508,N_10690);
nand U11664 (N_11664,N_10254,N_10559);
or U11665 (N_11665,N_10992,N_10557);
xor U11666 (N_11666,N_10945,N_10769);
nor U11667 (N_11667,N_10209,N_10582);
or U11668 (N_11668,N_10316,N_10454);
or U11669 (N_11669,N_10117,N_10676);
or U11670 (N_11670,N_10249,N_10314);
nand U11671 (N_11671,N_10341,N_10492);
or U11672 (N_11672,N_10329,N_10708);
nor U11673 (N_11673,N_10958,N_10242);
or U11674 (N_11674,N_10373,N_10252);
or U11675 (N_11675,N_10783,N_10066);
or U11676 (N_11676,N_10672,N_10746);
and U11677 (N_11677,N_10278,N_10449);
xor U11678 (N_11678,N_10600,N_10482);
xnor U11679 (N_11679,N_10959,N_10229);
or U11680 (N_11680,N_10819,N_10678);
xor U11681 (N_11681,N_10972,N_10587);
nand U11682 (N_11682,N_10010,N_10041);
or U11683 (N_11683,N_10760,N_10093);
or U11684 (N_11684,N_10957,N_10822);
nor U11685 (N_11685,N_10805,N_10112);
and U11686 (N_11686,N_10175,N_10975);
nor U11687 (N_11687,N_10370,N_10031);
xnor U11688 (N_11688,N_10736,N_10033);
nor U11689 (N_11689,N_10997,N_10389);
nor U11690 (N_11690,N_10545,N_10395);
and U11691 (N_11691,N_10781,N_10832);
nor U11692 (N_11692,N_10936,N_10242);
nor U11693 (N_11693,N_10771,N_10172);
nand U11694 (N_11694,N_10910,N_10078);
or U11695 (N_11695,N_10286,N_10440);
or U11696 (N_11696,N_10932,N_10784);
nor U11697 (N_11697,N_10170,N_10364);
nor U11698 (N_11698,N_10538,N_10386);
xor U11699 (N_11699,N_10487,N_10599);
xnor U11700 (N_11700,N_10575,N_10611);
nor U11701 (N_11701,N_10028,N_10658);
nand U11702 (N_11702,N_10468,N_10741);
and U11703 (N_11703,N_10237,N_10442);
xor U11704 (N_11704,N_10074,N_10985);
and U11705 (N_11705,N_10778,N_10215);
and U11706 (N_11706,N_10171,N_10676);
nor U11707 (N_11707,N_10527,N_10072);
and U11708 (N_11708,N_10775,N_10205);
or U11709 (N_11709,N_10574,N_10648);
nor U11710 (N_11710,N_10899,N_10972);
or U11711 (N_11711,N_10181,N_10974);
nor U11712 (N_11712,N_10786,N_10251);
nor U11713 (N_11713,N_10945,N_10646);
nor U11714 (N_11714,N_10251,N_10962);
xor U11715 (N_11715,N_10683,N_10819);
and U11716 (N_11716,N_10844,N_10036);
nand U11717 (N_11717,N_10539,N_10934);
nand U11718 (N_11718,N_10384,N_10294);
or U11719 (N_11719,N_10153,N_10792);
and U11720 (N_11720,N_10709,N_10319);
or U11721 (N_11721,N_10403,N_10279);
xor U11722 (N_11722,N_10162,N_10605);
nor U11723 (N_11723,N_10771,N_10760);
and U11724 (N_11724,N_10253,N_10376);
and U11725 (N_11725,N_10496,N_10280);
and U11726 (N_11726,N_10539,N_10212);
nor U11727 (N_11727,N_10363,N_10027);
and U11728 (N_11728,N_10448,N_10413);
nor U11729 (N_11729,N_10840,N_10830);
nand U11730 (N_11730,N_10850,N_10711);
xor U11731 (N_11731,N_10768,N_10292);
nand U11732 (N_11732,N_10356,N_10092);
and U11733 (N_11733,N_10345,N_10739);
nand U11734 (N_11734,N_10935,N_10312);
and U11735 (N_11735,N_10041,N_10665);
xnor U11736 (N_11736,N_10518,N_10496);
or U11737 (N_11737,N_10480,N_10998);
nor U11738 (N_11738,N_10941,N_10865);
nor U11739 (N_11739,N_10270,N_10041);
and U11740 (N_11740,N_10939,N_10687);
xor U11741 (N_11741,N_10805,N_10829);
nor U11742 (N_11742,N_10260,N_10484);
or U11743 (N_11743,N_10704,N_10407);
and U11744 (N_11744,N_10956,N_10923);
nand U11745 (N_11745,N_10804,N_10894);
xnor U11746 (N_11746,N_10158,N_10827);
nand U11747 (N_11747,N_10596,N_10537);
or U11748 (N_11748,N_10890,N_10119);
or U11749 (N_11749,N_10157,N_10209);
or U11750 (N_11750,N_10018,N_10034);
and U11751 (N_11751,N_10876,N_10079);
nand U11752 (N_11752,N_10695,N_10009);
nor U11753 (N_11753,N_10501,N_10875);
and U11754 (N_11754,N_10640,N_10883);
and U11755 (N_11755,N_10262,N_10878);
nand U11756 (N_11756,N_10848,N_10738);
nor U11757 (N_11757,N_10953,N_10877);
nand U11758 (N_11758,N_10620,N_10204);
nor U11759 (N_11759,N_10138,N_10968);
or U11760 (N_11760,N_10422,N_10138);
nand U11761 (N_11761,N_10435,N_10210);
or U11762 (N_11762,N_10149,N_10139);
and U11763 (N_11763,N_10277,N_10638);
or U11764 (N_11764,N_10235,N_10300);
nand U11765 (N_11765,N_10070,N_10251);
nand U11766 (N_11766,N_10898,N_10202);
nor U11767 (N_11767,N_10631,N_10043);
and U11768 (N_11768,N_10074,N_10807);
or U11769 (N_11769,N_10844,N_10216);
nand U11770 (N_11770,N_10452,N_10838);
nor U11771 (N_11771,N_10569,N_10270);
or U11772 (N_11772,N_10194,N_10566);
or U11773 (N_11773,N_10052,N_10714);
and U11774 (N_11774,N_10849,N_10725);
and U11775 (N_11775,N_10338,N_10113);
or U11776 (N_11776,N_10348,N_10012);
and U11777 (N_11777,N_10074,N_10284);
and U11778 (N_11778,N_10826,N_10241);
nor U11779 (N_11779,N_10475,N_10911);
nor U11780 (N_11780,N_10489,N_10801);
nor U11781 (N_11781,N_10388,N_10054);
or U11782 (N_11782,N_10556,N_10033);
nand U11783 (N_11783,N_10666,N_10079);
or U11784 (N_11784,N_10505,N_10017);
and U11785 (N_11785,N_10288,N_10327);
and U11786 (N_11786,N_10965,N_10024);
nand U11787 (N_11787,N_10328,N_10405);
nand U11788 (N_11788,N_10553,N_10807);
xnor U11789 (N_11789,N_10807,N_10315);
xnor U11790 (N_11790,N_10239,N_10184);
and U11791 (N_11791,N_10755,N_10088);
nor U11792 (N_11792,N_10266,N_10746);
nand U11793 (N_11793,N_10540,N_10709);
and U11794 (N_11794,N_10835,N_10919);
or U11795 (N_11795,N_10743,N_10076);
and U11796 (N_11796,N_10483,N_10164);
and U11797 (N_11797,N_10355,N_10466);
and U11798 (N_11798,N_10604,N_10429);
nor U11799 (N_11799,N_10243,N_10731);
nor U11800 (N_11800,N_10100,N_10197);
nor U11801 (N_11801,N_10788,N_10486);
or U11802 (N_11802,N_10717,N_10700);
nor U11803 (N_11803,N_10492,N_10798);
and U11804 (N_11804,N_10130,N_10735);
and U11805 (N_11805,N_10414,N_10114);
and U11806 (N_11806,N_10455,N_10388);
nand U11807 (N_11807,N_10254,N_10989);
and U11808 (N_11808,N_10453,N_10121);
nand U11809 (N_11809,N_10757,N_10492);
nor U11810 (N_11810,N_10381,N_10389);
and U11811 (N_11811,N_10890,N_10759);
nand U11812 (N_11812,N_10833,N_10498);
and U11813 (N_11813,N_10508,N_10665);
and U11814 (N_11814,N_10545,N_10478);
and U11815 (N_11815,N_10435,N_10639);
nand U11816 (N_11816,N_10617,N_10683);
and U11817 (N_11817,N_10758,N_10860);
and U11818 (N_11818,N_10470,N_10814);
and U11819 (N_11819,N_10019,N_10233);
nand U11820 (N_11820,N_10396,N_10670);
nand U11821 (N_11821,N_10584,N_10163);
xnor U11822 (N_11822,N_10034,N_10748);
nand U11823 (N_11823,N_10841,N_10189);
nand U11824 (N_11824,N_10951,N_10008);
and U11825 (N_11825,N_10759,N_10000);
xnor U11826 (N_11826,N_10437,N_10431);
nor U11827 (N_11827,N_10492,N_10960);
nor U11828 (N_11828,N_10620,N_10097);
or U11829 (N_11829,N_10264,N_10396);
and U11830 (N_11830,N_10363,N_10830);
nand U11831 (N_11831,N_10167,N_10166);
nor U11832 (N_11832,N_10695,N_10788);
nand U11833 (N_11833,N_10074,N_10401);
and U11834 (N_11834,N_10821,N_10708);
nand U11835 (N_11835,N_10775,N_10416);
xor U11836 (N_11836,N_10124,N_10633);
and U11837 (N_11837,N_10209,N_10447);
nand U11838 (N_11838,N_10942,N_10817);
nand U11839 (N_11839,N_10959,N_10012);
nand U11840 (N_11840,N_10989,N_10099);
and U11841 (N_11841,N_10865,N_10085);
nor U11842 (N_11842,N_10594,N_10932);
or U11843 (N_11843,N_10260,N_10289);
and U11844 (N_11844,N_10586,N_10003);
nand U11845 (N_11845,N_10171,N_10400);
nor U11846 (N_11846,N_10687,N_10739);
or U11847 (N_11847,N_10468,N_10226);
or U11848 (N_11848,N_10519,N_10037);
and U11849 (N_11849,N_10323,N_10953);
nor U11850 (N_11850,N_10520,N_10394);
nor U11851 (N_11851,N_10122,N_10635);
nor U11852 (N_11852,N_10035,N_10515);
xnor U11853 (N_11853,N_10961,N_10230);
and U11854 (N_11854,N_10186,N_10509);
or U11855 (N_11855,N_10507,N_10629);
or U11856 (N_11856,N_10404,N_10947);
nand U11857 (N_11857,N_10808,N_10976);
nand U11858 (N_11858,N_10167,N_10668);
or U11859 (N_11859,N_10657,N_10799);
nor U11860 (N_11860,N_10087,N_10393);
or U11861 (N_11861,N_10033,N_10763);
and U11862 (N_11862,N_10941,N_10641);
xnor U11863 (N_11863,N_10034,N_10740);
nand U11864 (N_11864,N_10163,N_10142);
and U11865 (N_11865,N_10917,N_10949);
or U11866 (N_11866,N_10095,N_10624);
and U11867 (N_11867,N_10985,N_10608);
or U11868 (N_11868,N_10691,N_10190);
nand U11869 (N_11869,N_10018,N_10200);
nor U11870 (N_11870,N_10187,N_10906);
nor U11871 (N_11871,N_10479,N_10906);
and U11872 (N_11872,N_10845,N_10561);
xnor U11873 (N_11873,N_10986,N_10719);
nor U11874 (N_11874,N_10398,N_10482);
and U11875 (N_11875,N_10288,N_10581);
xnor U11876 (N_11876,N_10164,N_10526);
or U11877 (N_11877,N_10868,N_10787);
or U11878 (N_11878,N_10204,N_10723);
or U11879 (N_11879,N_10428,N_10582);
and U11880 (N_11880,N_10785,N_10187);
and U11881 (N_11881,N_10729,N_10416);
nand U11882 (N_11882,N_10504,N_10295);
xor U11883 (N_11883,N_10902,N_10864);
or U11884 (N_11884,N_10796,N_10942);
nand U11885 (N_11885,N_10318,N_10602);
and U11886 (N_11886,N_10994,N_10241);
nor U11887 (N_11887,N_10791,N_10502);
nor U11888 (N_11888,N_10952,N_10031);
or U11889 (N_11889,N_10765,N_10266);
or U11890 (N_11890,N_10123,N_10390);
and U11891 (N_11891,N_10027,N_10993);
or U11892 (N_11892,N_10693,N_10281);
nor U11893 (N_11893,N_10071,N_10628);
nand U11894 (N_11894,N_10859,N_10651);
or U11895 (N_11895,N_10645,N_10691);
xnor U11896 (N_11896,N_10831,N_10059);
nand U11897 (N_11897,N_10900,N_10760);
or U11898 (N_11898,N_10189,N_10905);
or U11899 (N_11899,N_10442,N_10541);
or U11900 (N_11900,N_10416,N_10888);
nor U11901 (N_11901,N_10283,N_10672);
or U11902 (N_11902,N_10272,N_10970);
xnor U11903 (N_11903,N_10750,N_10846);
nor U11904 (N_11904,N_10614,N_10061);
or U11905 (N_11905,N_10344,N_10822);
and U11906 (N_11906,N_10966,N_10721);
and U11907 (N_11907,N_10876,N_10698);
xnor U11908 (N_11908,N_10323,N_10988);
and U11909 (N_11909,N_10573,N_10911);
nor U11910 (N_11910,N_10706,N_10595);
and U11911 (N_11911,N_10200,N_10623);
and U11912 (N_11912,N_10509,N_10654);
or U11913 (N_11913,N_10048,N_10944);
nand U11914 (N_11914,N_10562,N_10768);
nor U11915 (N_11915,N_10176,N_10817);
or U11916 (N_11916,N_10504,N_10635);
nor U11917 (N_11917,N_10677,N_10234);
or U11918 (N_11918,N_10770,N_10967);
nor U11919 (N_11919,N_10311,N_10122);
nor U11920 (N_11920,N_10474,N_10429);
and U11921 (N_11921,N_10277,N_10570);
and U11922 (N_11922,N_10892,N_10282);
nand U11923 (N_11923,N_10427,N_10120);
nand U11924 (N_11924,N_10767,N_10573);
nand U11925 (N_11925,N_10015,N_10841);
nor U11926 (N_11926,N_10847,N_10364);
nand U11927 (N_11927,N_10292,N_10388);
nor U11928 (N_11928,N_10344,N_10452);
nor U11929 (N_11929,N_10119,N_10917);
nor U11930 (N_11930,N_10987,N_10703);
or U11931 (N_11931,N_10917,N_10815);
and U11932 (N_11932,N_10999,N_10935);
or U11933 (N_11933,N_10412,N_10263);
or U11934 (N_11934,N_10971,N_10989);
xnor U11935 (N_11935,N_10331,N_10228);
or U11936 (N_11936,N_10754,N_10492);
or U11937 (N_11937,N_10390,N_10244);
nor U11938 (N_11938,N_10894,N_10769);
xnor U11939 (N_11939,N_10222,N_10363);
or U11940 (N_11940,N_10060,N_10393);
and U11941 (N_11941,N_10395,N_10059);
xnor U11942 (N_11942,N_10306,N_10798);
and U11943 (N_11943,N_10953,N_10907);
nor U11944 (N_11944,N_10124,N_10594);
or U11945 (N_11945,N_10216,N_10815);
or U11946 (N_11946,N_10323,N_10697);
xor U11947 (N_11947,N_10058,N_10776);
nor U11948 (N_11948,N_10796,N_10383);
nor U11949 (N_11949,N_10066,N_10091);
and U11950 (N_11950,N_10752,N_10527);
nand U11951 (N_11951,N_10737,N_10098);
nor U11952 (N_11952,N_10358,N_10771);
nand U11953 (N_11953,N_10090,N_10526);
nor U11954 (N_11954,N_10687,N_10163);
and U11955 (N_11955,N_10197,N_10345);
and U11956 (N_11956,N_10365,N_10461);
and U11957 (N_11957,N_10511,N_10548);
nand U11958 (N_11958,N_10420,N_10553);
nand U11959 (N_11959,N_10233,N_10368);
nor U11960 (N_11960,N_10183,N_10572);
nor U11961 (N_11961,N_10381,N_10041);
nand U11962 (N_11962,N_10288,N_10090);
or U11963 (N_11963,N_10434,N_10521);
nor U11964 (N_11964,N_10862,N_10596);
nand U11965 (N_11965,N_10337,N_10881);
nand U11966 (N_11966,N_10234,N_10189);
or U11967 (N_11967,N_10847,N_10970);
xor U11968 (N_11968,N_10514,N_10912);
xnor U11969 (N_11969,N_10877,N_10755);
nor U11970 (N_11970,N_10604,N_10632);
or U11971 (N_11971,N_10614,N_10826);
or U11972 (N_11972,N_10444,N_10045);
nor U11973 (N_11973,N_10973,N_10287);
or U11974 (N_11974,N_10489,N_10949);
xor U11975 (N_11975,N_10719,N_10690);
nor U11976 (N_11976,N_10995,N_10119);
or U11977 (N_11977,N_10721,N_10527);
xor U11978 (N_11978,N_10635,N_10676);
or U11979 (N_11979,N_10834,N_10738);
nor U11980 (N_11980,N_10392,N_10638);
nand U11981 (N_11981,N_10348,N_10204);
nor U11982 (N_11982,N_10259,N_10628);
or U11983 (N_11983,N_10840,N_10324);
nor U11984 (N_11984,N_10772,N_10752);
xor U11985 (N_11985,N_10968,N_10061);
nor U11986 (N_11986,N_10995,N_10515);
nor U11987 (N_11987,N_10350,N_10488);
nor U11988 (N_11988,N_10232,N_10533);
nand U11989 (N_11989,N_10366,N_10841);
nor U11990 (N_11990,N_10757,N_10223);
or U11991 (N_11991,N_10361,N_10543);
or U11992 (N_11992,N_10269,N_10282);
xor U11993 (N_11993,N_10278,N_10797);
and U11994 (N_11994,N_10312,N_10358);
or U11995 (N_11995,N_10529,N_10715);
or U11996 (N_11996,N_10858,N_10193);
and U11997 (N_11997,N_10238,N_10262);
or U11998 (N_11998,N_10719,N_10679);
or U11999 (N_11999,N_10767,N_10577);
nand U12000 (N_12000,N_11077,N_11877);
or U12001 (N_12001,N_11871,N_11254);
nand U12002 (N_12002,N_11236,N_11846);
nand U12003 (N_12003,N_11943,N_11243);
xnor U12004 (N_12004,N_11592,N_11750);
or U12005 (N_12005,N_11714,N_11476);
or U12006 (N_12006,N_11951,N_11845);
and U12007 (N_12007,N_11699,N_11352);
or U12008 (N_12008,N_11582,N_11895);
nor U12009 (N_12009,N_11210,N_11090);
and U12010 (N_12010,N_11291,N_11333);
nor U12011 (N_12011,N_11514,N_11079);
and U12012 (N_12012,N_11506,N_11889);
or U12013 (N_12013,N_11121,N_11744);
or U12014 (N_12014,N_11452,N_11302);
nor U12015 (N_12015,N_11171,N_11158);
or U12016 (N_12016,N_11635,N_11983);
and U12017 (N_12017,N_11162,N_11349);
nor U12018 (N_12018,N_11838,N_11773);
nand U12019 (N_12019,N_11651,N_11567);
nand U12020 (N_12020,N_11425,N_11284);
nor U12021 (N_12021,N_11030,N_11135);
and U12022 (N_12022,N_11029,N_11998);
or U12023 (N_12023,N_11320,N_11404);
nor U12024 (N_12024,N_11874,N_11763);
xnor U12025 (N_12025,N_11016,N_11550);
and U12026 (N_12026,N_11536,N_11681);
and U12027 (N_12027,N_11769,N_11534);
nor U12028 (N_12028,N_11081,N_11814);
nor U12029 (N_12029,N_11644,N_11042);
and U12030 (N_12030,N_11579,N_11001);
nand U12031 (N_12031,N_11310,N_11208);
xnor U12032 (N_12032,N_11419,N_11387);
and U12033 (N_12033,N_11562,N_11321);
nor U12034 (N_12034,N_11554,N_11545);
and U12035 (N_12035,N_11264,N_11782);
and U12036 (N_12036,N_11199,N_11695);
nand U12037 (N_12037,N_11609,N_11747);
and U12038 (N_12038,N_11612,N_11606);
or U12039 (N_12039,N_11849,N_11745);
and U12040 (N_12040,N_11794,N_11500);
or U12041 (N_12041,N_11881,N_11867);
or U12042 (N_12042,N_11980,N_11361);
nor U12043 (N_12043,N_11702,N_11484);
and U12044 (N_12044,N_11356,N_11667);
and U12045 (N_12045,N_11824,N_11385);
or U12046 (N_12046,N_11143,N_11442);
and U12047 (N_12047,N_11923,N_11422);
or U12048 (N_12048,N_11429,N_11522);
and U12049 (N_12049,N_11239,N_11383);
nor U12050 (N_12050,N_11549,N_11212);
and U12051 (N_12051,N_11891,N_11656);
and U12052 (N_12052,N_11602,N_11682);
nor U12053 (N_12053,N_11398,N_11839);
nand U12054 (N_12054,N_11053,N_11069);
or U12055 (N_12055,N_11386,N_11965);
nor U12056 (N_12056,N_11961,N_11289);
and U12057 (N_12057,N_11257,N_11924);
nand U12058 (N_12058,N_11293,N_11049);
or U12059 (N_12059,N_11156,N_11481);
xor U12060 (N_12060,N_11104,N_11395);
or U12061 (N_12061,N_11409,N_11338);
nand U12062 (N_12062,N_11604,N_11066);
nor U12063 (N_12063,N_11344,N_11672);
nand U12064 (N_12064,N_11444,N_11477);
or U12065 (N_12065,N_11724,N_11987);
nor U12066 (N_12066,N_11250,N_11326);
nand U12067 (N_12067,N_11125,N_11453);
nand U12068 (N_12068,N_11022,N_11648);
and U12069 (N_12069,N_11560,N_11973);
nand U12070 (N_12070,N_11529,N_11054);
or U12071 (N_12071,N_11775,N_11365);
nor U12072 (N_12072,N_11428,N_11229);
nor U12073 (N_12073,N_11465,N_11979);
nand U12074 (N_12074,N_11211,N_11064);
and U12075 (N_12075,N_11013,N_11581);
nor U12076 (N_12076,N_11274,N_11245);
nand U12077 (N_12077,N_11155,N_11524);
and U12078 (N_12078,N_11263,N_11863);
nor U12079 (N_12079,N_11508,N_11046);
or U12080 (N_12080,N_11886,N_11176);
nor U12081 (N_12081,N_11780,N_11128);
nand U12082 (N_12082,N_11455,N_11901);
nand U12083 (N_12083,N_11905,N_11397);
and U12084 (N_12084,N_11706,N_11220);
xnor U12085 (N_12085,N_11255,N_11677);
nor U12086 (N_12086,N_11828,N_11177);
nor U12087 (N_12087,N_11134,N_11223);
nor U12088 (N_12088,N_11768,N_11730);
and U12089 (N_12089,N_11840,N_11527);
and U12090 (N_12090,N_11723,N_11811);
and U12091 (N_12091,N_11370,N_11312);
xor U12092 (N_12092,N_11778,N_11486);
or U12093 (N_12093,N_11993,N_11201);
or U12094 (N_12094,N_11096,N_11258);
xor U12095 (N_12095,N_11078,N_11160);
or U12096 (N_12096,N_11072,N_11627);
or U12097 (N_12097,N_11411,N_11140);
nand U12098 (N_12098,N_11615,N_11842);
and U12099 (N_12099,N_11926,N_11329);
xor U12100 (N_12100,N_11178,N_11466);
nor U12101 (N_12101,N_11721,N_11770);
or U12102 (N_12102,N_11503,N_11463);
or U12103 (N_12103,N_11447,N_11292);
nand U12104 (N_12104,N_11711,N_11087);
and U12105 (N_12105,N_11108,N_11678);
or U12106 (N_12106,N_11456,N_11316);
nand U12107 (N_12107,N_11671,N_11313);
nor U12108 (N_12108,N_11643,N_11531);
and U12109 (N_12109,N_11153,N_11192);
or U12110 (N_12110,N_11832,N_11005);
nor U12111 (N_12111,N_11319,N_11185);
nor U12112 (N_12112,N_11417,N_11253);
or U12113 (N_12113,N_11556,N_11434);
and U12114 (N_12114,N_11114,N_11573);
xnor U12115 (N_12115,N_11939,N_11958);
nand U12116 (N_12116,N_11804,N_11431);
and U12117 (N_12117,N_11106,N_11538);
or U12118 (N_12118,N_11198,N_11897);
or U12119 (N_12119,N_11646,N_11517);
nor U12120 (N_12120,N_11812,N_11376);
nor U12121 (N_12121,N_11869,N_11642);
and U12122 (N_12122,N_11179,N_11729);
or U12123 (N_12123,N_11019,N_11371);
and U12124 (N_12124,N_11577,N_11414);
nor U12125 (N_12125,N_11184,N_11661);
nor U12126 (N_12126,N_11787,N_11304);
nand U12127 (N_12127,N_11910,N_11918);
and U12128 (N_12128,N_11995,N_11323);
nor U12129 (N_12129,N_11488,N_11962);
nor U12130 (N_12130,N_11970,N_11570);
nand U12131 (N_12131,N_11168,N_11443);
and U12132 (N_12132,N_11265,N_11836);
nand U12133 (N_12133,N_11260,N_11172);
nor U12134 (N_12134,N_11107,N_11413);
and U12135 (N_12135,N_11240,N_11718);
nand U12136 (N_12136,N_11753,N_11922);
xor U12137 (N_12137,N_11144,N_11194);
nand U12138 (N_12138,N_11530,N_11613);
nand U12139 (N_12139,N_11969,N_11098);
or U12140 (N_12140,N_11080,N_11708);
or U12141 (N_12141,N_11318,N_11688);
nand U12142 (N_12142,N_11767,N_11189);
nand U12143 (N_12143,N_11410,N_11354);
nand U12144 (N_12144,N_11296,N_11197);
nand U12145 (N_12145,N_11544,N_11948);
and U12146 (N_12146,N_11468,N_11335);
nor U12147 (N_12147,N_11216,N_11345);
nor U12148 (N_12148,N_11805,N_11990);
and U12149 (N_12149,N_11563,N_11626);
and U12150 (N_12150,N_11213,N_11774);
xor U12151 (N_12151,N_11328,N_11136);
or U12152 (N_12152,N_11362,N_11101);
and U12153 (N_12153,N_11006,N_11887);
and U12154 (N_12154,N_11650,N_11813);
nand U12155 (N_12155,N_11149,N_11132);
nor U12156 (N_12156,N_11789,N_11252);
nor U12157 (N_12157,N_11587,N_11683);
nand U12158 (N_12158,N_11050,N_11408);
nor U12159 (N_12159,N_11788,N_11139);
or U12160 (N_12160,N_11940,N_11652);
and U12161 (N_12161,N_11148,N_11935);
nand U12162 (N_12162,N_11623,N_11464);
and U12163 (N_12163,N_11966,N_11272);
nand U12164 (N_12164,N_11917,N_11955);
or U12165 (N_12165,N_11416,N_11232);
nor U12166 (N_12166,N_11543,N_11694);
nor U12167 (N_12167,N_11301,N_11366);
nor U12168 (N_12168,N_11390,N_11621);
xnor U12169 (N_12169,N_11857,N_11781);
and U12170 (N_12170,N_11707,N_11834);
or U12171 (N_12171,N_11147,N_11214);
nand U12172 (N_12172,N_11424,N_11637);
xor U12173 (N_12173,N_11692,N_11916);
xor U12174 (N_12174,N_11401,N_11547);
nor U12175 (N_12175,N_11262,N_11472);
and U12176 (N_12176,N_11848,N_11566);
nor U12177 (N_12177,N_11430,N_11827);
xor U12178 (N_12178,N_11009,N_11535);
nor U12179 (N_12179,N_11892,N_11188);
nand U12180 (N_12180,N_11141,N_11756);
and U12181 (N_12181,N_11331,N_11608);
or U12182 (N_12182,N_11084,N_11498);
nand U12183 (N_12183,N_11382,N_11883);
nor U12184 (N_12184,N_11475,N_11680);
nand U12185 (N_12185,N_11640,N_11010);
and U12186 (N_12186,N_11421,N_11467);
nor U12187 (N_12187,N_11752,N_11696);
and U12188 (N_12188,N_11297,N_11954);
nor U12189 (N_12189,N_11012,N_11673);
and U12190 (N_12190,N_11283,N_11499);
nand U12191 (N_12191,N_11890,N_11186);
and U12192 (N_12192,N_11266,N_11818);
nor U12193 (N_12193,N_11028,N_11523);
nand U12194 (N_12194,N_11574,N_11632);
xor U12195 (N_12195,N_11526,N_11070);
nand U12196 (N_12196,N_11594,N_11116);
nand U12197 (N_12197,N_11516,N_11306);
nand U12198 (N_12198,N_11357,N_11256);
nor U12199 (N_12199,N_11525,N_11518);
nor U12200 (N_12200,N_11393,N_11580);
nand U12201 (N_12201,N_11837,N_11088);
and U12202 (N_12202,N_11728,N_11949);
nand U12203 (N_12203,N_11299,N_11553);
or U12204 (N_12204,N_11348,N_11657);
and U12205 (N_12205,N_11666,N_11164);
nor U12206 (N_12206,N_11600,N_11909);
or U12207 (N_12207,N_11709,N_11377);
nor U12208 (N_12208,N_11616,N_11669);
or U12209 (N_12209,N_11737,N_11654);
and U12210 (N_12210,N_11440,N_11548);
and U12211 (N_12211,N_11882,N_11865);
and U12212 (N_12212,N_11461,N_11884);
nor U12213 (N_12213,N_11533,N_11094);
nand U12214 (N_12214,N_11539,N_11187);
or U12215 (N_12215,N_11795,N_11858);
or U12216 (N_12216,N_11624,N_11802);
nor U12217 (N_12217,N_11457,N_11927);
nor U12218 (N_12218,N_11492,N_11639);
nor U12219 (N_12219,N_11697,N_11485);
xor U12220 (N_12220,N_11900,N_11375);
and U12221 (N_12221,N_11314,N_11379);
xor U12222 (N_12222,N_11057,N_11938);
or U12223 (N_12223,N_11269,N_11131);
nand U12224 (N_12224,N_11885,N_11843);
nand U12225 (N_12225,N_11315,N_11145);
xnor U12226 (N_12226,N_11427,N_11816);
or U12227 (N_12227,N_11165,N_11378);
xor U12228 (N_12228,N_11278,N_11967);
and U12229 (N_12229,N_11809,N_11275);
and U12230 (N_12230,N_11436,N_11908);
xnor U12231 (N_12231,N_11031,N_11311);
and U12232 (N_12232,N_11290,N_11180);
and U12233 (N_12233,N_11037,N_11268);
nand U12234 (N_12234,N_11700,N_11203);
and U12235 (N_12235,N_11822,N_11929);
nand U12236 (N_12236,N_11879,N_11873);
and U12237 (N_12237,N_11451,N_11551);
xnor U12238 (N_12238,N_11294,N_11823);
nor U12239 (N_12239,N_11614,N_11607);
or U12240 (N_12240,N_11835,N_11668);
nand U12241 (N_12241,N_11693,N_11618);
nand U12242 (N_12242,N_11964,N_11373);
nor U12243 (N_12243,N_11280,N_11925);
nor U12244 (N_12244,N_11052,N_11074);
and U12245 (N_12245,N_11282,N_11799);
or U12246 (N_12246,N_11633,N_11117);
nand U12247 (N_12247,N_11450,N_11821);
nor U12248 (N_12248,N_11032,N_11023);
or U12249 (N_12249,N_11512,N_11025);
and U12250 (N_12250,N_11933,N_11771);
nor U12251 (N_12251,N_11137,N_11638);
xor U12252 (N_12252,N_11439,N_11986);
xor U12253 (N_12253,N_11241,N_11270);
and U12254 (N_12254,N_11586,N_11803);
xor U12255 (N_12255,N_11852,N_11124);
nand U12256 (N_12256,N_11878,N_11462);
or U12257 (N_12257,N_11020,N_11097);
nor U12258 (N_12258,N_11303,N_11433);
xor U12259 (N_12259,N_11758,N_11636);
xnor U12260 (N_12260,N_11571,N_11739);
nor U12261 (N_12261,N_11120,N_11992);
nor U12262 (N_12262,N_11941,N_11276);
nor U12263 (N_12263,N_11994,N_11620);
nor U12264 (N_12264,N_11670,N_11797);
nand U12265 (N_12265,N_11285,N_11267);
nor U12266 (N_12266,N_11710,N_11853);
and U12267 (N_12267,N_11991,N_11764);
nor U12268 (N_12268,N_11118,N_11099);
nand U12269 (N_12269,N_11222,N_11662);
xor U12270 (N_12270,N_11972,N_11641);
nand U12271 (N_12271,N_11625,N_11899);
nand U12272 (N_12272,N_11279,N_11287);
or U12273 (N_12273,N_11261,N_11095);
nor U12274 (N_12274,N_11784,N_11583);
nand U12275 (N_12275,N_11062,N_11575);
and U12276 (N_12276,N_11438,N_11202);
nand U12277 (N_12277,N_11847,N_11528);
nor U12278 (N_12278,N_11045,N_11235);
or U12279 (N_12279,N_11934,N_11217);
nand U12280 (N_12280,N_11898,N_11996);
nor U12281 (N_12281,N_11322,N_11051);
nand U12282 (N_12282,N_11561,N_11113);
nor U12283 (N_12283,N_11205,N_11532);
or U12284 (N_12284,N_11792,N_11734);
and U12285 (N_12285,N_11068,N_11937);
or U12286 (N_12286,N_11237,N_11815);
nand U12287 (N_12287,N_11478,N_11719);
and U12288 (N_12288,N_11585,N_11684);
or U12289 (N_12289,N_11565,N_11740);
or U12290 (N_12290,N_11244,N_11482);
nor U12291 (N_12291,N_11687,N_11448);
and U12292 (N_12292,N_11412,N_11127);
xor U12293 (N_12293,N_11913,N_11112);
nand U12294 (N_12294,N_11957,N_11590);
or U12295 (N_12295,N_11988,N_11449);
or U12296 (N_12296,N_11645,N_11494);
and U12297 (N_12297,N_11277,N_11713);
nor U12298 (N_12298,N_11369,N_11219);
nand U12299 (N_12299,N_11601,N_11100);
nand U12300 (N_12300,N_11743,N_11946);
and U12301 (N_12301,N_11800,N_11295);
nor U12302 (N_12302,N_11435,N_11950);
xor U12303 (N_12303,N_11520,N_11251);
or U12304 (N_12304,N_11327,N_11055);
nor U12305 (N_12305,N_11975,N_11493);
nand U12306 (N_12306,N_11474,N_11381);
xor U12307 (N_12307,N_11231,N_11437);
or U12308 (N_12308,N_11584,N_11405);
nand U12309 (N_12309,N_11402,N_11190);
nand U12310 (N_12310,N_11854,N_11446);
and U12311 (N_12311,N_11930,N_11655);
nand U12312 (N_12312,N_11021,N_11904);
nand U12313 (N_12313,N_11083,N_11002);
xor U12314 (N_12314,N_11163,N_11350);
and U12315 (N_12315,N_11082,N_11597);
nand U12316 (N_12316,N_11552,N_11521);
and U12317 (N_12317,N_11757,N_11830);
and U12318 (N_12318,N_11075,N_11035);
or U12319 (N_12319,N_11558,N_11833);
nor U12320 (N_12320,N_11173,N_11353);
nand U12321 (N_12321,N_11974,N_11791);
nor U12322 (N_12322,N_11872,N_11036);
or U12323 (N_12323,N_11167,N_11856);
nor U12324 (N_12324,N_11230,N_11859);
nand U12325 (N_12325,N_11762,N_11591);
or U12326 (N_12326,N_11460,N_11491);
or U12327 (N_12327,N_11047,N_11346);
or U12328 (N_12328,N_11919,N_11091);
nor U12329 (N_12329,N_11110,N_11902);
or U12330 (N_12330,N_11426,N_11007);
or U12331 (N_12331,N_11751,N_11334);
or U12332 (N_12332,N_11109,N_11479);
and U12333 (N_12333,N_11086,N_11720);
xnor U12334 (N_12334,N_11589,N_11779);
nor U12335 (N_12335,N_11542,N_11564);
or U12336 (N_12336,N_11674,N_11454);
nand U12337 (N_12337,N_11071,N_11073);
and U12338 (N_12338,N_11505,N_11206);
and U12339 (N_12339,N_11698,N_11896);
nor U12340 (N_12340,N_11459,N_11391);
nand U12341 (N_12341,N_11907,N_11701);
or U12342 (N_12342,N_11796,N_11207);
or U12343 (N_12343,N_11027,N_11741);
or U12344 (N_12344,N_11105,N_11004);
and U12345 (N_12345,N_11906,N_11942);
and U12346 (N_12346,N_11248,N_11415);
nor U12347 (N_12347,N_11717,N_11689);
nand U12348 (N_12348,N_11649,N_11634);
or U12349 (N_12349,N_11611,N_11420);
or U12350 (N_12350,N_11396,N_11510);
xnor U12351 (N_12351,N_11765,N_11281);
nand U12352 (N_12352,N_11738,N_11242);
nor U12353 (N_12353,N_11932,N_11166);
or U12354 (N_12354,N_11195,N_11324);
and U12355 (N_12355,N_11722,N_11894);
or U12356 (N_12356,N_11507,N_11509);
nor U12357 (N_12357,N_11806,N_11473);
or U12358 (N_12358,N_11159,N_11018);
and U12359 (N_12359,N_11471,N_11928);
or U12360 (N_12360,N_11039,N_11384);
or U12361 (N_12361,N_11617,N_11102);
nand U12362 (N_12362,N_11766,N_11749);
and U12363 (N_12363,N_11423,N_11130);
nand U12364 (N_12364,N_11759,N_11691);
or U12365 (N_12365,N_11952,N_11048);
nand U12366 (N_12366,N_11685,N_11920);
nand U12367 (N_12367,N_11196,N_11487);
nand U12368 (N_12368,N_11540,N_11150);
xnor U12369 (N_12369,N_11690,N_11546);
xnor U12370 (N_12370,N_11191,N_11953);
nor U12371 (N_12371,N_11981,N_11663);
nor U12372 (N_12372,N_11568,N_11271);
and U12373 (N_12373,N_11968,N_11676);
nor U12374 (N_12374,N_11831,N_11161);
nand U12375 (N_12375,N_11142,N_11569);
nor U12376 (N_12376,N_11619,N_11407);
nand U12377 (N_12377,N_11664,N_11059);
nor U12378 (N_12378,N_11228,N_11599);
and U12379 (N_12379,N_11793,N_11754);
or U12380 (N_12380,N_11576,N_11122);
xor U12381 (N_12381,N_11458,N_11497);
nor U12382 (N_12382,N_11880,N_11798);
and U12383 (N_12383,N_11736,N_11971);
and U12384 (N_12384,N_11989,N_11513);
or U12385 (N_12385,N_11945,N_11033);
xor U12386 (N_12386,N_11286,N_11174);
nor U12387 (N_12387,N_11870,N_11469);
nor U12388 (N_12388,N_11123,N_11598);
xor U12389 (N_12389,N_11999,N_11735);
nor U12390 (N_12390,N_11658,N_11596);
or U12391 (N_12391,N_11157,N_11665);
xor U12392 (N_12392,N_11403,N_11786);
and U12393 (N_12393,N_11193,N_11183);
nor U12394 (N_12394,N_11043,N_11629);
or U12395 (N_12395,N_11686,N_11067);
and U12396 (N_12396,N_11209,N_11234);
or U12397 (N_12397,N_11982,N_11238);
xnor U12398 (N_12398,N_11772,N_11363);
nor U12399 (N_12399,N_11703,N_11912);
nor U12400 (N_12400,N_11496,N_11034);
nor U12401 (N_12401,N_11914,N_11631);
and U12402 (N_12402,N_11725,N_11727);
nor U12403 (N_12403,N_11038,N_11519);
nor U12404 (N_12404,N_11227,N_11876);
or U12405 (N_12405,N_11888,N_11182);
and U12406 (N_12406,N_11380,N_11247);
and U12407 (N_12407,N_11841,N_11483);
and U12408 (N_12408,N_11810,N_11445);
nand U12409 (N_12409,N_11400,N_11441);
nand U12410 (N_12410,N_11317,N_11515);
or U12411 (N_12411,N_11808,N_11399);
and U12412 (N_12412,N_11392,N_11578);
xnor U12413 (N_12413,N_11151,N_11976);
xnor U12414 (N_12414,N_11480,N_11011);
and U12415 (N_12415,N_11092,N_11221);
and U12416 (N_12416,N_11470,N_11343);
or U12417 (N_12417,N_11200,N_11820);
or U12418 (N_12418,N_11921,N_11175);
or U12419 (N_12419,N_11777,N_11489);
or U12420 (N_12420,N_11298,N_11418);
or U12421 (N_12421,N_11307,N_11790);
nor U12422 (N_12422,N_11305,N_11588);
and U12423 (N_12423,N_11374,N_11855);
and U12424 (N_12424,N_11978,N_11732);
nor U12425 (N_12425,N_11541,N_11259);
nor U12426 (N_12426,N_11504,N_11061);
or U12427 (N_12427,N_11893,N_11060);
nand U12428 (N_12428,N_11785,N_11911);
nor U12429 (N_12429,N_11659,N_11861);
and U12430 (N_12430,N_11537,N_11603);
nor U12431 (N_12431,N_11406,N_11358);
and U12432 (N_12432,N_11224,N_11014);
and U12433 (N_12433,N_11860,N_11605);
nor U12434 (N_12434,N_11628,N_11829);
or U12435 (N_12435,N_11704,N_11040);
and U12436 (N_12436,N_11817,N_11063);
or U12437 (N_12437,N_11129,N_11003);
or U12438 (N_12438,N_11760,N_11862);
nand U12439 (N_12439,N_11931,N_11355);
nand U12440 (N_12440,N_11093,N_11807);
nor U12441 (N_12441,N_11501,N_11984);
nand U12442 (N_12442,N_11360,N_11715);
or U12443 (N_12443,N_11000,N_11875);
or U12444 (N_12444,N_11015,N_11115);
and U12445 (N_12445,N_11850,N_11226);
nand U12446 (N_12446,N_11065,N_11742);
or U12447 (N_12447,N_11325,N_11056);
and U12448 (N_12448,N_11716,N_11364);
nor U12449 (N_12449,N_11026,N_11776);
or U12450 (N_12450,N_11336,N_11339);
nor U12451 (N_12451,N_11170,N_11731);
or U12452 (N_12452,N_11660,N_11308);
nor U12453 (N_12453,N_11089,N_11273);
or U12454 (N_12454,N_11630,N_11300);
and U12455 (N_12455,N_11342,N_11783);
nor U12456 (N_12456,N_11389,N_11372);
nor U12457 (N_12457,N_11755,N_11246);
or U12458 (N_12458,N_11309,N_11748);
and U12459 (N_12459,N_11337,N_11705);
nand U12460 (N_12460,N_11915,N_11733);
nand U12461 (N_12461,N_11559,N_11490);
and U12462 (N_12462,N_11152,N_11225);
and U12463 (N_12463,N_11944,N_11368);
or U12464 (N_12464,N_11555,N_11249);
nor U12465 (N_12465,N_11181,N_11947);
and U12466 (N_12466,N_11218,N_11595);
or U12467 (N_12467,N_11985,N_11233);
and U12468 (N_12468,N_11864,N_11367);
nor U12469 (N_12469,N_11432,N_11959);
or U12470 (N_12470,N_11977,N_11936);
nor U12471 (N_12471,N_11746,N_11044);
and U12472 (N_12472,N_11557,N_11511);
and U12473 (N_12473,N_11085,N_11351);
nand U12474 (N_12474,N_11963,N_11801);
xor U12475 (N_12475,N_11572,N_11204);
xnor U12476 (N_12476,N_11997,N_11712);
or U12477 (N_12477,N_11154,N_11647);
and U12478 (N_12478,N_11126,N_11146);
or U12479 (N_12479,N_11388,N_11119);
and U12480 (N_12480,N_11495,N_11169);
and U12481 (N_12481,N_11076,N_11394);
or U12482 (N_12482,N_11347,N_11851);
nor U12483 (N_12483,N_11041,N_11960);
nand U12484 (N_12484,N_11866,N_11868);
nor U12485 (N_12485,N_11138,N_11215);
xnor U12486 (N_12486,N_11330,N_11826);
xor U12487 (N_12487,N_11761,N_11726);
nor U12488 (N_12488,N_11111,N_11653);
and U12489 (N_12489,N_11008,N_11956);
nor U12490 (N_12490,N_11024,N_11825);
and U12491 (N_12491,N_11288,N_11340);
and U12492 (N_12492,N_11133,N_11332);
or U12493 (N_12493,N_11610,N_11844);
or U12494 (N_12494,N_11341,N_11058);
xor U12495 (N_12495,N_11622,N_11593);
nor U12496 (N_12496,N_11103,N_11017);
and U12497 (N_12497,N_11359,N_11502);
nand U12498 (N_12498,N_11819,N_11903);
or U12499 (N_12499,N_11679,N_11675);
or U12500 (N_12500,N_11587,N_11552);
nand U12501 (N_12501,N_11238,N_11795);
nand U12502 (N_12502,N_11368,N_11009);
nand U12503 (N_12503,N_11785,N_11446);
nor U12504 (N_12504,N_11484,N_11563);
or U12505 (N_12505,N_11017,N_11829);
nor U12506 (N_12506,N_11027,N_11627);
or U12507 (N_12507,N_11109,N_11606);
nand U12508 (N_12508,N_11530,N_11151);
or U12509 (N_12509,N_11751,N_11436);
nor U12510 (N_12510,N_11679,N_11687);
or U12511 (N_12511,N_11842,N_11707);
nand U12512 (N_12512,N_11536,N_11714);
and U12513 (N_12513,N_11848,N_11772);
or U12514 (N_12514,N_11977,N_11746);
nand U12515 (N_12515,N_11868,N_11005);
or U12516 (N_12516,N_11310,N_11542);
or U12517 (N_12517,N_11602,N_11356);
and U12518 (N_12518,N_11291,N_11098);
nor U12519 (N_12519,N_11444,N_11426);
xnor U12520 (N_12520,N_11090,N_11140);
nand U12521 (N_12521,N_11240,N_11708);
nand U12522 (N_12522,N_11436,N_11753);
and U12523 (N_12523,N_11535,N_11388);
or U12524 (N_12524,N_11242,N_11867);
nand U12525 (N_12525,N_11722,N_11857);
nand U12526 (N_12526,N_11017,N_11105);
nor U12527 (N_12527,N_11548,N_11727);
and U12528 (N_12528,N_11905,N_11157);
xnor U12529 (N_12529,N_11177,N_11183);
xor U12530 (N_12530,N_11875,N_11294);
nor U12531 (N_12531,N_11436,N_11115);
nor U12532 (N_12532,N_11516,N_11583);
nand U12533 (N_12533,N_11659,N_11859);
and U12534 (N_12534,N_11455,N_11917);
nand U12535 (N_12535,N_11188,N_11388);
and U12536 (N_12536,N_11993,N_11829);
nand U12537 (N_12537,N_11887,N_11294);
nor U12538 (N_12538,N_11826,N_11913);
nand U12539 (N_12539,N_11349,N_11036);
or U12540 (N_12540,N_11439,N_11316);
and U12541 (N_12541,N_11253,N_11178);
nor U12542 (N_12542,N_11380,N_11744);
and U12543 (N_12543,N_11204,N_11773);
nor U12544 (N_12544,N_11823,N_11986);
nor U12545 (N_12545,N_11376,N_11106);
nor U12546 (N_12546,N_11080,N_11896);
or U12547 (N_12547,N_11636,N_11990);
nand U12548 (N_12548,N_11605,N_11103);
or U12549 (N_12549,N_11502,N_11829);
or U12550 (N_12550,N_11895,N_11445);
nor U12551 (N_12551,N_11141,N_11014);
or U12552 (N_12552,N_11299,N_11480);
and U12553 (N_12553,N_11483,N_11964);
nor U12554 (N_12554,N_11092,N_11248);
nand U12555 (N_12555,N_11808,N_11918);
nor U12556 (N_12556,N_11262,N_11033);
nor U12557 (N_12557,N_11578,N_11916);
and U12558 (N_12558,N_11587,N_11412);
or U12559 (N_12559,N_11580,N_11292);
or U12560 (N_12560,N_11101,N_11038);
or U12561 (N_12561,N_11445,N_11323);
nor U12562 (N_12562,N_11662,N_11407);
nor U12563 (N_12563,N_11413,N_11865);
and U12564 (N_12564,N_11131,N_11117);
xor U12565 (N_12565,N_11552,N_11762);
nand U12566 (N_12566,N_11450,N_11545);
xor U12567 (N_12567,N_11047,N_11222);
and U12568 (N_12568,N_11081,N_11101);
xor U12569 (N_12569,N_11313,N_11725);
and U12570 (N_12570,N_11363,N_11723);
or U12571 (N_12571,N_11809,N_11499);
nor U12572 (N_12572,N_11935,N_11221);
nor U12573 (N_12573,N_11249,N_11608);
nand U12574 (N_12574,N_11418,N_11875);
and U12575 (N_12575,N_11372,N_11493);
and U12576 (N_12576,N_11582,N_11642);
or U12577 (N_12577,N_11639,N_11250);
and U12578 (N_12578,N_11089,N_11216);
nor U12579 (N_12579,N_11368,N_11442);
nor U12580 (N_12580,N_11991,N_11063);
nor U12581 (N_12581,N_11510,N_11829);
or U12582 (N_12582,N_11233,N_11055);
and U12583 (N_12583,N_11619,N_11870);
and U12584 (N_12584,N_11187,N_11443);
nand U12585 (N_12585,N_11828,N_11125);
and U12586 (N_12586,N_11690,N_11229);
nor U12587 (N_12587,N_11582,N_11781);
nor U12588 (N_12588,N_11012,N_11951);
nor U12589 (N_12589,N_11827,N_11968);
xnor U12590 (N_12590,N_11991,N_11163);
xor U12591 (N_12591,N_11959,N_11618);
or U12592 (N_12592,N_11336,N_11207);
nand U12593 (N_12593,N_11735,N_11113);
nor U12594 (N_12594,N_11101,N_11393);
xor U12595 (N_12595,N_11792,N_11762);
nor U12596 (N_12596,N_11686,N_11872);
or U12597 (N_12597,N_11905,N_11692);
nor U12598 (N_12598,N_11858,N_11178);
and U12599 (N_12599,N_11761,N_11251);
nand U12600 (N_12600,N_11561,N_11864);
or U12601 (N_12601,N_11682,N_11107);
nand U12602 (N_12602,N_11475,N_11652);
and U12603 (N_12603,N_11436,N_11250);
or U12604 (N_12604,N_11621,N_11097);
nor U12605 (N_12605,N_11112,N_11764);
and U12606 (N_12606,N_11691,N_11025);
nand U12607 (N_12607,N_11131,N_11863);
or U12608 (N_12608,N_11972,N_11843);
nand U12609 (N_12609,N_11480,N_11354);
nand U12610 (N_12610,N_11135,N_11181);
nand U12611 (N_12611,N_11433,N_11383);
xnor U12612 (N_12612,N_11257,N_11865);
nand U12613 (N_12613,N_11840,N_11979);
nor U12614 (N_12614,N_11389,N_11625);
or U12615 (N_12615,N_11544,N_11899);
and U12616 (N_12616,N_11952,N_11046);
and U12617 (N_12617,N_11773,N_11597);
nor U12618 (N_12618,N_11307,N_11394);
nor U12619 (N_12619,N_11863,N_11653);
xor U12620 (N_12620,N_11427,N_11316);
and U12621 (N_12621,N_11792,N_11217);
nor U12622 (N_12622,N_11919,N_11721);
nor U12623 (N_12623,N_11859,N_11484);
and U12624 (N_12624,N_11037,N_11756);
and U12625 (N_12625,N_11062,N_11045);
nor U12626 (N_12626,N_11914,N_11940);
and U12627 (N_12627,N_11920,N_11908);
and U12628 (N_12628,N_11174,N_11307);
nand U12629 (N_12629,N_11038,N_11871);
and U12630 (N_12630,N_11208,N_11185);
nor U12631 (N_12631,N_11379,N_11492);
nand U12632 (N_12632,N_11103,N_11482);
nand U12633 (N_12633,N_11453,N_11105);
nor U12634 (N_12634,N_11051,N_11160);
or U12635 (N_12635,N_11480,N_11594);
nor U12636 (N_12636,N_11235,N_11189);
nand U12637 (N_12637,N_11962,N_11436);
nor U12638 (N_12638,N_11287,N_11794);
or U12639 (N_12639,N_11773,N_11719);
and U12640 (N_12640,N_11633,N_11569);
and U12641 (N_12641,N_11680,N_11265);
nor U12642 (N_12642,N_11315,N_11978);
nand U12643 (N_12643,N_11442,N_11372);
nor U12644 (N_12644,N_11800,N_11042);
and U12645 (N_12645,N_11534,N_11207);
nor U12646 (N_12646,N_11797,N_11046);
or U12647 (N_12647,N_11768,N_11076);
and U12648 (N_12648,N_11817,N_11905);
nand U12649 (N_12649,N_11718,N_11852);
and U12650 (N_12650,N_11552,N_11938);
and U12651 (N_12651,N_11269,N_11246);
and U12652 (N_12652,N_11194,N_11488);
and U12653 (N_12653,N_11752,N_11693);
nand U12654 (N_12654,N_11451,N_11745);
xnor U12655 (N_12655,N_11990,N_11064);
nor U12656 (N_12656,N_11319,N_11621);
and U12657 (N_12657,N_11663,N_11591);
and U12658 (N_12658,N_11782,N_11545);
nand U12659 (N_12659,N_11871,N_11821);
xor U12660 (N_12660,N_11838,N_11699);
nand U12661 (N_12661,N_11163,N_11024);
nor U12662 (N_12662,N_11762,N_11682);
and U12663 (N_12663,N_11584,N_11847);
nor U12664 (N_12664,N_11551,N_11005);
nor U12665 (N_12665,N_11051,N_11433);
or U12666 (N_12666,N_11852,N_11812);
nor U12667 (N_12667,N_11214,N_11291);
or U12668 (N_12668,N_11011,N_11902);
nand U12669 (N_12669,N_11267,N_11009);
and U12670 (N_12670,N_11364,N_11646);
nand U12671 (N_12671,N_11582,N_11650);
and U12672 (N_12672,N_11150,N_11109);
or U12673 (N_12673,N_11066,N_11117);
nor U12674 (N_12674,N_11009,N_11495);
or U12675 (N_12675,N_11585,N_11743);
nand U12676 (N_12676,N_11053,N_11410);
or U12677 (N_12677,N_11273,N_11513);
nor U12678 (N_12678,N_11498,N_11411);
nor U12679 (N_12679,N_11402,N_11105);
xnor U12680 (N_12680,N_11720,N_11797);
or U12681 (N_12681,N_11421,N_11886);
nor U12682 (N_12682,N_11340,N_11847);
nand U12683 (N_12683,N_11192,N_11669);
nor U12684 (N_12684,N_11118,N_11903);
or U12685 (N_12685,N_11225,N_11154);
or U12686 (N_12686,N_11331,N_11939);
nor U12687 (N_12687,N_11967,N_11915);
nor U12688 (N_12688,N_11806,N_11639);
or U12689 (N_12689,N_11852,N_11870);
or U12690 (N_12690,N_11054,N_11515);
and U12691 (N_12691,N_11882,N_11385);
and U12692 (N_12692,N_11474,N_11418);
and U12693 (N_12693,N_11845,N_11410);
nor U12694 (N_12694,N_11776,N_11473);
nor U12695 (N_12695,N_11983,N_11574);
nand U12696 (N_12696,N_11519,N_11180);
nand U12697 (N_12697,N_11495,N_11205);
or U12698 (N_12698,N_11166,N_11463);
nor U12699 (N_12699,N_11550,N_11185);
and U12700 (N_12700,N_11654,N_11900);
nor U12701 (N_12701,N_11224,N_11533);
and U12702 (N_12702,N_11534,N_11420);
xor U12703 (N_12703,N_11003,N_11894);
nor U12704 (N_12704,N_11768,N_11428);
nor U12705 (N_12705,N_11733,N_11370);
or U12706 (N_12706,N_11295,N_11197);
nor U12707 (N_12707,N_11222,N_11500);
and U12708 (N_12708,N_11448,N_11363);
and U12709 (N_12709,N_11769,N_11473);
nor U12710 (N_12710,N_11104,N_11546);
and U12711 (N_12711,N_11721,N_11059);
nand U12712 (N_12712,N_11329,N_11622);
xnor U12713 (N_12713,N_11222,N_11942);
and U12714 (N_12714,N_11062,N_11362);
or U12715 (N_12715,N_11025,N_11716);
and U12716 (N_12716,N_11130,N_11621);
and U12717 (N_12717,N_11337,N_11087);
or U12718 (N_12718,N_11844,N_11340);
or U12719 (N_12719,N_11330,N_11966);
and U12720 (N_12720,N_11647,N_11965);
or U12721 (N_12721,N_11345,N_11035);
nand U12722 (N_12722,N_11831,N_11642);
nor U12723 (N_12723,N_11568,N_11958);
or U12724 (N_12724,N_11834,N_11031);
xor U12725 (N_12725,N_11610,N_11791);
nand U12726 (N_12726,N_11252,N_11516);
nand U12727 (N_12727,N_11988,N_11369);
nand U12728 (N_12728,N_11134,N_11696);
nand U12729 (N_12729,N_11155,N_11681);
or U12730 (N_12730,N_11529,N_11100);
nor U12731 (N_12731,N_11584,N_11539);
nor U12732 (N_12732,N_11270,N_11040);
and U12733 (N_12733,N_11133,N_11538);
and U12734 (N_12734,N_11273,N_11758);
or U12735 (N_12735,N_11110,N_11688);
or U12736 (N_12736,N_11467,N_11528);
nor U12737 (N_12737,N_11934,N_11178);
or U12738 (N_12738,N_11638,N_11100);
xnor U12739 (N_12739,N_11347,N_11216);
nor U12740 (N_12740,N_11225,N_11316);
nand U12741 (N_12741,N_11680,N_11450);
nor U12742 (N_12742,N_11091,N_11515);
xnor U12743 (N_12743,N_11161,N_11169);
or U12744 (N_12744,N_11764,N_11531);
and U12745 (N_12745,N_11848,N_11350);
nor U12746 (N_12746,N_11959,N_11132);
nand U12747 (N_12747,N_11606,N_11311);
or U12748 (N_12748,N_11603,N_11473);
and U12749 (N_12749,N_11754,N_11132);
nand U12750 (N_12750,N_11688,N_11773);
and U12751 (N_12751,N_11551,N_11467);
or U12752 (N_12752,N_11049,N_11808);
or U12753 (N_12753,N_11448,N_11346);
or U12754 (N_12754,N_11798,N_11587);
and U12755 (N_12755,N_11187,N_11964);
or U12756 (N_12756,N_11090,N_11687);
and U12757 (N_12757,N_11906,N_11103);
and U12758 (N_12758,N_11872,N_11996);
nor U12759 (N_12759,N_11402,N_11031);
xnor U12760 (N_12760,N_11365,N_11868);
or U12761 (N_12761,N_11962,N_11283);
nand U12762 (N_12762,N_11761,N_11085);
nor U12763 (N_12763,N_11008,N_11586);
nand U12764 (N_12764,N_11962,N_11483);
nor U12765 (N_12765,N_11091,N_11997);
nand U12766 (N_12766,N_11658,N_11935);
nor U12767 (N_12767,N_11403,N_11859);
or U12768 (N_12768,N_11692,N_11562);
or U12769 (N_12769,N_11315,N_11333);
nor U12770 (N_12770,N_11554,N_11562);
and U12771 (N_12771,N_11886,N_11485);
nor U12772 (N_12772,N_11096,N_11132);
xor U12773 (N_12773,N_11769,N_11461);
and U12774 (N_12774,N_11478,N_11625);
and U12775 (N_12775,N_11164,N_11765);
or U12776 (N_12776,N_11684,N_11941);
nor U12777 (N_12777,N_11449,N_11173);
or U12778 (N_12778,N_11154,N_11616);
nor U12779 (N_12779,N_11584,N_11153);
nor U12780 (N_12780,N_11663,N_11089);
nand U12781 (N_12781,N_11566,N_11167);
xnor U12782 (N_12782,N_11311,N_11769);
or U12783 (N_12783,N_11303,N_11218);
or U12784 (N_12784,N_11276,N_11415);
and U12785 (N_12785,N_11544,N_11054);
nand U12786 (N_12786,N_11313,N_11213);
or U12787 (N_12787,N_11137,N_11961);
nand U12788 (N_12788,N_11227,N_11217);
nor U12789 (N_12789,N_11496,N_11661);
nand U12790 (N_12790,N_11973,N_11847);
nand U12791 (N_12791,N_11703,N_11359);
nor U12792 (N_12792,N_11325,N_11868);
or U12793 (N_12793,N_11039,N_11984);
xor U12794 (N_12794,N_11966,N_11937);
nor U12795 (N_12795,N_11414,N_11262);
or U12796 (N_12796,N_11684,N_11525);
nor U12797 (N_12797,N_11052,N_11724);
and U12798 (N_12798,N_11719,N_11407);
and U12799 (N_12799,N_11270,N_11299);
and U12800 (N_12800,N_11212,N_11790);
or U12801 (N_12801,N_11873,N_11768);
nand U12802 (N_12802,N_11145,N_11171);
nor U12803 (N_12803,N_11589,N_11100);
and U12804 (N_12804,N_11397,N_11273);
or U12805 (N_12805,N_11119,N_11330);
xnor U12806 (N_12806,N_11077,N_11720);
or U12807 (N_12807,N_11555,N_11848);
nand U12808 (N_12808,N_11732,N_11746);
and U12809 (N_12809,N_11770,N_11742);
nor U12810 (N_12810,N_11449,N_11937);
nand U12811 (N_12811,N_11161,N_11311);
and U12812 (N_12812,N_11170,N_11531);
or U12813 (N_12813,N_11106,N_11428);
nor U12814 (N_12814,N_11362,N_11044);
or U12815 (N_12815,N_11799,N_11828);
and U12816 (N_12816,N_11992,N_11895);
nor U12817 (N_12817,N_11297,N_11520);
nand U12818 (N_12818,N_11137,N_11394);
or U12819 (N_12819,N_11919,N_11331);
xnor U12820 (N_12820,N_11662,N_11332);
or U12821 (N_12821,N_11509,N_11680);
or U12822 (N_12822,N_11215,N_11265);
nand U12823 (N_12823,N_11258,N_11023);
nand U12824 (N_12824,N_11904,N_11892);
and U12825 (N_12825,N_11288,N_11005);
and U12826 (N_12826,N_11486,N_11501);
xnor U12827 (N_12827,N_11455,N_11855);
nand U12828 (N_12828,N_11244,N_11490);
nand U12829 (N_12829,N_11198,N_11210);
nand U12830 (N_12830,N_11768,N_11077);
and U12831 (N_12831,N_11600,N_11725);
nand U12832 (N_12832,N_11841,N_11155);
nor U12833 (N_12833,N_11443,N_11300);
nor U12834 (N_12834,N_11294,N_11343);
and U12835 (N_12835,N_11266,N_11522);
and U12836 (N_12836,N_11477,N_11301);
and U12837 (N_12837,N_11720,N_11332);
nand U12838 (N_12838,N_11728,N_11499);
and U12839 (N_12839,N_11021,N_11254);
nor U12840 (N_12840,N_11854,N_11989);
or U12841 (N_12841,N_11986,N_11474);
nor U12842 (N_12842,N_11332,N_11344);
nand U12843 (N_12843,N_11667,N_11657);
or U12844 (N_12844,N_11759,N_11301);
xor U12845 (N_12845,N_11387,N_11695);
xnor U12846 (N_12846,N_11638,N_11970);
nand U12847 (N_12847,N_11121,N_11212);
and U12848 (N_12848,N_11500,N_11835);
or U12849 (N_12849,N_11734,N_11737);
and U12850 (N_12850,N_11297,N_11880);
nand U12851 (N_12851,N_11889,N_11233);
and U12852 (N_12852,N_11618,N_11914);
or U12853 (N_12853,N_11147,N_11799);
and U12854 (N_12854,N_11406,N_11597);
or U12855 (N_12855,N_11047,N_11458);
nand U12856 (N_12856,N_11902,N_11024);
and U12857 (N_12857,N_11800,N_11657);
nor U12858 (N_12858,N_11541,N_11069);
and U12859 (N_12859,N_11523,N_11349);
nor U12860 (N_12860,N_11943,N_11401);
and U12861 (N_12861,N_11275,N_11479);
or U12862 (N_12862,N_11513,N_11150);
or U12863 (N_12863,N_11384,N_11584);
or U12864 (N_12864,N_11843,N_11657);
nand U12865 (N_12865,N_11734,N_11246);
nand U12866 (N_12866,N_11081,N_11940);
nor U12867 (N_12867,N_11537,N_11818);
or U12868 (N_12868,N_11793,N_11362);
and U12869 (N_12869,N_11666,N_11832);
nand U12870 (N_12870,N_11133,N_11214);
or U12871 (N_12871,N_11272,N_11579);
nand U12872 (N_12872,N_11150,N_11895);
nand U12873 (N_12873,N_11919,N_11451);
or U12874 (N_12874,N_11400,N_11157);
and U12875 (N_12875,N_11592,N_11297);
nand U12876 (N_12876,N_11473,N_11167);
or U12877 (N_12877,N_11046,N_11049);
and U12878 (N_12878,N_11829,N_11585);
nor U12879 (N_12879,N_11907,N_11412);
or U12880 (N_12880,N_11506,N_11681);
or U12881 (N_12881,N_11237,N_11792);
and U12882 (N_12882,N_11422,N_11525);
or U12883 (N_12883,N_11408,N_11692);
nand U12884 (N_12884,N_11569,N_11597);
nand U12885 (N_12885,N_11115,N_11414);
and U12886 (N_12886,N_11996,N_11710);
nand U12887 (N_12887,N_11719,N_11336);
and U12888 (N_12888,N_11630,N_11021);
xor U12889 (N_12889,N_11436,N_11332);
nor U12890 (N_12890,N_11259,N_11570);
and U12891 (N_12891,N_11111,N_11927);
nor U12892 (N_12892,N_11177,N_11505);
nand U12893 (N_12893,N_11041,N_11956);
nand U12894 (N_12894,N_11757,N_11398);
nor U12895 (N_12895,N_11074,N_11803);
nor U12896 (N_12896,N_11292,N_11374);
and U12897 (N_12897,N_11566,N_11486);
and U12898 (N_12898,N_11508,N_11902);
nor U12899 (N_12899,N_11372,N_11358);
xor U12900 (N_12900,N_11404,N_11082);
nand U12901 (N_12901,N_11294,N_11719);
nand U12902 (N_12902,N_11002,N_11917);
nor U12903 (N_12903,N_11833,N_11078);
xor U12904 (N_12904,N_11259,N_11270);
and U12905 (N_12905,N_11097,N_11504);
nand U12906 (N_12906,N_11302,N_11431);
or U12907 (N_12907,N_11581,N_11594);
nand U12908 (N_12908,N_11580,N_11568);
nor U12909 (N_12909,N_11567,N_11547);
nand U12910 (N_12910,N_11706,N_11265);
and U12911 (N_12911,N_11600,N_11049);
and U12912 (N_12912,N_11028,N_11026);
or U12913 (N_12913,N_11896,N_11764);
nor U12914 (N_12914,N_11358,N_11160);
or U12915 (N_12915,N_11415,N_11028);
xnor U12916 (N_12916,N_11285,N_11938);
or U12917 (N_12917,N_11432,N_11662);
and U12918 (N_12918,N_11973,N_11540);
xnor U12919 (N_12919,N_11884,N_11399);
nor U12920 (N_12920,N_11780,N_11875);
or U12921 (N_12921,N_11990,N_11470);
and U12922 (N_12922,N_11210,N_11362);
xor U12923 (N_12923,N_11541,N_11114);
and U12924 (N_12924,N_11615,N_11318);
or U12925 (N_12925,N_11362,N_11435);
nor U12926 (N_12926,N_11617,N_11501);
xor U12927 (N_12927,N_11913,N_11322);
and U12928 (N_12928,N_11944,N_11007);
or U12929 (N_12929,N_11297,N_11047);
and U12930 (N_12930,N_11435,N_11529);
or U12931 (N_12931,N_11679,N_11953);
xnor U12932 (N_12932,N_11002,N_11108);
nand U12933 (N_12933,N_11904,N_11340);
and U12934 (N_12934,N_11014,N_11762);
xor U12935 (N_12935,N_11034,N_11851);
and U12936 (N_12936,N_11727,N_11364);
and U12937 (N_12937,N_11376,N_11519);
and U12938 (N_12938,N_11608,N_11513);
nor U12939 (N_12939,N_11495,N_11556);
and U12940 (N_12940,N_11773,N_11190);
and U12941 (N_12941,N_11879,N_11668);
nand U12942 (N_12942,N_11135,N_11598);
or U12943 (N_12943,N_11444,N_11965);
and U12944 (N_12944,N_11689,N_11526);
and U12945 (N_12945,N_11843,N_11485);
or U12946 (N_12946,N_11824,N_11304);
xor U12947 (N_12947,N_11251,N_11825);
nand U12948 (N_12948,N_11422,N_11113);
nand U12949 (N_12949,N_11081,N_11952);
nor U12950 (N_12950,N_11260,N_11151);
and U12951 (N_12951,N_11097,N_11926);
nand U12952 (N_12952,N_11157,N_11278);
nor U12953 (N_12953,N_11213,N_11206);
and U12954 (N_12954,N_11209,N_11686);
or U12955 (N_12955,N_11662,N_11537);
nand U12956 (N_12956,N_11623,N_11319);
and U12957 (N_12957,N_11035,N_11072);
nor U12958 (N_12958,N_11270,N_11743);
or U12959 (N_12959,N_11176,N_11316);
nor U12960 (N_12960,N_11989,N_11090);
nor U12961 (N_12961,N_11430,N_11274);
nand U12962 (N_12962,N_11678,N_11131);
nand U12963 (N_12963,N_11952,N_11303);
and U12964 (N_12964,N_11028,N_11231);
nor U12965 (N_12965,N_11746,N_11962);
nor U12966 (N_12966,N_11015,N_11471);
xnor U12967 (N_12967,N_11518,N_11663);
nand U12968 (N_12968,N_11679,N_11967);
nand U12969 (N_12969,N_11754,N_11347);
and U12970 (N_12970,N_11722,N_11730);
nor U12971 (N_12971,N_11635,N_11918);
nand U12972 (N_12972,N_11797,N_11106);
nand U12973 (N_12973,N_11656,N_11038);
nand U12974 (N_12974,N_11633,N_11968);
nor U12975 (N_12975,N_11495,N_11647);
nor U12976 (N_12976,N_11171,N_11160);
or U12977 (N_12977,N_11089,N_11825);
nor U12978 (N_12978,N_11652,N_11633);
and U12979 (N_12979,N_11547,N_11912);
nand U12980 (N_12980,N_11230,N_11022);
or U12981 (N_12981,N_11607,N_11756);
nand U12982 (N_12982,N_11960,N_11242);
nor U12983 (N_12983,N_11064,N_11675);
and U12984 (N_12984,N_11725,N_11139);
xor U12985 (N_12985,N_11244,N_11263);
nor U12986 (N_12986,N_11857,N_11124);
nand U12987 (N_12987,N_11827,N_11445);
xor U12988 (N_12988,N_11958,N_11734);
nor U12989 (N_12989,N_11738,N_11218);
nand U12990 (N_12990,N_11638,N_11138);
or U12991 (N_12991,N_11414,N_11055);
nor U12992 (N_12992,N_11837,N_11196);
nand U12993 (N_12993,N_11601,N_11590);
nand U12994 (N_12994,N_11602,N_11708);
and U12995 (N_12995,N_11838,N_11154);
nor U12996 (N_12996,N_11510,N_11275);
and U12997 (N_12997,N_11354,N_11681);
and U12998 (N_12998,N_11547,N_11262);
and U12999 (N_12999,N_11921,N_11655);
nand U13000 (N_13000,N_12380,N_12893);
nor U13001 (N_13001,N_12370,N_12153);
nor U13002 (N_13002,N_12693,N_12514);
nand U13003 (N_13003,N_12906,N_12409);
xnor U13004 (N_13004,N_12467,N_12272);
xor U13005 (N_13005,N_12349,N_12899);
and U13006 (N_13006,N_12322,N_12260);
nor U13007 (N_13007,N_12085,N_12532);
nand U13008 (N_13008,N_12989,N_12655);
nor U13009 (N_13009,N_12821,N_12478);
and U13010 (N_13010,N_12427,N_12143);
or U13011 (N_13011,N_12844,N_12545);
nand U13012 (N_13012,N_12887,N_12807);
or U13013 (N_13013,N_12238,N_12820);
and U13014 (N_13014,N_12160,N_12193);
and U13015 (N_13015,N_12399,N_12988);
nand U13016 (N_13016,N_12895,N_12750);
or U13017 (N_13017,N_12882,N_12840);
nor U13018 (N_13018,N_12069,N_12410);
nor U13019 (N_13019,N_12635,N_12862);
nand U13020 (N_13020,N_12429,N_12256);
nor U13021 (N_13021,N_12659,N_12582);
or U13022 (N_13022,N_12047,N_12498);
and U13023 (N_13023,N_12401,N_12691);
nor U13024 (N_13024,N_12888,N_12363);
nor U13025 (N_13025,N_12152,N_12639);
nor U13026 (N_13026,N_12034,N_12088);
or U13027 (N_13027,N_12967,N_12361);
and U13028 (N_13028,N_12879,N_12802);
nand U13029 (N_13029,N_12800,N_12938);
and U13030 (N_13030,N_12516,N_12930);
nand U13031 (N_13031,N_12289,N_12051);
nor U13032 (N_13032,N_12412,N_12651);
or U13033 (N_13033,N_12298,N_12027);
and U13034 (N_13034,N_12884,N_12985);
or U13035 (N_13035,N_12687,N_12058);
nand U13036 (N_13036,N_12759,N_12373);
or U13037 (N_13037,N_12019,N_12515);
nand U13038 (N_13038,N_12479,N_12053);
nand U13039 (N_13039,N_12773,N_12061);
or U13040 (N_13040,N_12346,N_12199);
and U13041 (N_13041,N_12350,N_12837);
or U13042 (N_13042,N_12677,N_12036);
nor U13043 (N_13043,N_12149,N_12777);
nand U13044 (N_13044,N_12682,N_12179);
and U13045 (N_13045,N_12225,N_12233);
or U13046 (N_13046,N_12081,N_12523);
nor U13047 (N_13047,N_12738,N_12797);
nor U13048 (N_13048,N_12236,N_12858);
nand U13049 (N_13049,N_12445,N_12644);
nand U13050 (N_13050,N_12245,N_12269);
or U13051 (N_13051,N_12737,N_12181);
and U13052 (N_13052,N_12836,N_12414);
nand U13053 (N_13053,N_12137,N_12084);
nor U13054 (N_13054,N_12045,N_12535);
nand U13055 (N_13055,N_12506,N_12568);
and U13056 (N_13056,N_12135,N_12130);
nand U13057 (N_13057,N_12709,N_12698);
nand U13058 (N_13058,N_12195,N_12933);
or U13059 (N_13059,N_12966,N_12267);
and U13060 (N_13060,N_12794,N_12360);
and U13061 (N_13061,N_12724,N_12287);
and U13062 (N_13062,N_12321,N_12940);
and U13063 (N_13063,N_12352,N_12652);
or U13064 (N_13064,N_12086,N_12851);
and U13065 (N_13065,N_12757,N_12695);
and U13066 (N_13066,N_12390,N_12681);
nor U13067 (N_13067,N_12751,N_12441);
nand U13068 (N_13068,N_12336,N_12089);
nand U13069 (N_13069,N_12871,N_12774);
nor U13070 (N_13070,N_12839,N_12743);
nand U13071 (N_13071,N_12834,N_12041);
or U13072 (N_13072,N_12620,N_12325);
and U13073 (N_13073,N_12144,N_12224);
nor U13074 (N_13074,N_12163,N_12612);
nand U13075 (N_13075,N_12883,N_12700);
and U13076 (N_13076,N_12301,N_12355);
nor U13077 (N_13077,N_12252,N_12830);
nor U13078 (N_13078,N_12952,N_12936);
and U13079 (N_13079,N_12408,N_12462);
nand U13080 (N_13080,N_12665,N_12753);
or U13081 (N_13081,N_12641,N_12011);
or U13082 (N_13082,N_12769,N_12673);
and U13083 (N_13083,N_12923,N_12662);
nand U13084 (N_13084,N_12071,N_12075);
nand U13085 (N_13085,N_12579,N_12021);
nor U13086 (N_13086,N_12881,N_12132);
nand U13087 (N_13087,N_12067,N_12495);
and U13088 (N_13088,N_12459,N_12196);
xor U13089 (N_13089,N_12022,N_12920);
nand U13090 (N_13090,N_12768,N_12124);
xnor U13091 (N_13091,N_12359,N_12904);
xor U13092 (N_13092,N_12250,N_12118);
nand U13093 (N_13093,N_12799,N_12500);
or U13094 (N_13094,N_12065,N_12537);
xnor U13095 (N_13095,N_12295,N_12310);
nand U13096 (N_13096,N_12551,N_12527);
nand U13097 (N_13097,N_12974,N_12491);
nor U13098 (N_13098,N_12793,N_12939);
or U13099 (N_13099,N_12365,N_12469);
nor U13100 (N_13100,N_12718,N_12372);
or U13101 (N_13101,N_12848,N_12158);
and U13102 (N_13102,N_12012,N_12711);
nor U13103 (N_13103,N_12969,N_12549);
nor U13104 (N_13104,N_12042,N_12726);
nor U13105 (N_13105,N_12804,N_12550);
and U13106 (N_13106,N_12131,N_12770);
or U13107 (N_13107,N_12020,N_12761);
or U13108 (N_13108,N_12645,N_12622);
and U13109 (N_13109,N_12186,N_12430);
and U13110 (N_13110,N_12251,N_12521);
or U13111 (N_13111,N_12120,N_12439);
nor U13112 (N_13112,N_12141,N_12099);
and U13113 (N_13113,N_12949,N_12362);
or U13114 (N_13114,N_12980,N_12388);
or U13115 (N_13115,N_12648,N_12182);
nand U13116 (N_13116,N_12745,N_12729);
nor U13117 (N_13117,N_12072,N_12063);
or U13118 (N_13118,N_12782,N_12519);
and U13119 (N_13119,N_12492,N_12323);
nand U13120 (N_13120,N_12091,N_12147);
nand U13121 (N_13121,N_12722,N_12766);
nor U13122 (N_13122,N_12563,N_12873);
nor U13123 (N_13123,N_12859,N_12314);
and U13124 (N_13124,N_12383,N_12932);
nand U13125 (N_13125,N_12822,N_12284);
or U13126 (N_13126,N_12771,N_12438);
or U13127 (N_13127,N_12092,N_12292);
nand U13128 (N_13128,N_12960,N_12159);
and U13129 (N_13129,N_12087,N_12801);
xor U13130 (N_13130,N_12157,N_12531);
nand U13131 (N_13131,N_12483,N_12207);
nand U13132 (N_13132,N_12277,N_12133);
nand U13133 (N_13133,N_12569,N_12249);
and U13134 (N_13134,N_12714,N_12843);
xnor U13135 (N_13135,N_12451,N_12596);
nand U13136 (N_13136,N_12235,N_12232);
nand U13137 (N_13137,N_12431,N_12209);
nor U13138 (N_13138,N_12869,N_12134);
nand U13139 (N_13139,N_12538,N_12338);
or U13140 (N_13140,N_12607,N_12449);
nor U13141 (N_13141,N_12922,N_12496);
and U13142 (N_13142,N_12198,N_12668);
nor U13143 (N_13143,N_12094,N_12337);
and U13144 (N_13144,N_12534,N_12995);
and U13145 (N_13145,N_12201,N_12572);
nor U13146 (N_13146,N_12202,N_12402);
or U13147 (N_13147,N_12795,N_12678);
nand U13148 (N_13148,N_12630,N_12744);
nor U13149 (N_13149,N_12046,N_12672);
nor U13150 (N_13150,N_12339,N_12145);
and U13151 (N_13151,N_12647,N_12205);
or U13152 (N_13152,N_12657,N_12817);
xor U13153 (N_13153,N_12707,N_12078);
and U13154 (N_13154,N_12642,N_12356);
or U13155 (N_13155,N_12405,N_12927);
and U13156 (N_13156,N_12216,N_12164);
nor U13157 (N_13157,N_12594,N_12841);
and U13158 (N_13158,N_12288,N_12981);
and U13159 (N_13159,N_12393,N_12090);
and U13160 (N_13160,N_12669,N_12253);
nor U13161 (N_13161,N_12796,N_12990);
nand U13162 (N_13162,N_12096,N_12508);
nand U13163 (N_13163,N_12611,N_12471);
nand U13164 (N_13164,N_12139,N_12870);
nor U13165 (N_13165,N_12931,N_12845);
nor U13166 (N_13166,N_12343,N_12230);
or U13167 (N_13167,N_12958,N_12993);
nor U13168 (N_13168,N_12320,N_12357);
nor U13169 (N_13169,N_12313,N_12876);
nand U13170 (N_13170,N_12852,N_12789);
nor U13171 (N_13171,N_12875,N_12849);
or U13172 (N_13172,N_12779,N_12917);
nand U13173 (N_13173,N_12161,N_12097);
nor U13174 (N_13174,N_12241,N_12690);
xnor U13175 (N_13175,N_12111,N_12348);
nor U13176 (N_13176,N_12294,N_12555);
nand U13177 (N_13177,N_12853,N_12998);
nand U13178 (N_13178,N_12727,N_12752);
nand U13179 (N_13179,N_12663,N_12608);
or U13180 (N_13180,N_12083,N_12542);
nor U13181 (N_13181,N_12615,N_12248);
nand U13182 (N_13182,N_12947,N_12983);
nand U13183 (N_13183,N_12525,N_12286);
and U13184 (N_13184,N_12300,N_12586);
and U13185 (N_13185,N_12942,N_12890);
and U13186 (N_13186,N_12315,N_12470);
nand U13187 (N_13187,N_12268,N_12577);
xor U13188 (N_13188,N_12511,N_12805);
and U13189 (N_13189,N_12055,N_12435);
nor U13190 (N_13190,N_12505,N_12835);
nand U13191 (N_13191,N_12452,N_12100);
nand U13192 (N_13192,N_12877,N_12842);
and U13193 (N_13193,N_12279,N_12244);
nand U13194 (N_13194,N_12378,N_12311);
nor U13195 (N_13195,N_12661,N_12103);
nor U13196 (N_13196,N_12627,N_12464);
nand U13197 (N_13197,N_12746,N_12602);
nand U13198 (N_13198,N_12318,N_12860);
nand U13199 (N_13199,N_12258,N_12623);
or U13200 (N_13200,N_12977,N_12706);
nand U13201 (N_13201,N_12214,N_12961);
and U13202 (N_13202,N_12271,N_12580);
and U13203 (N_13203,N_12710,N_12255);
or U13204 (N_13204,N_12048,N_12861);
nand U13205 (N_13205,N_12562,N_12674);
nor U13206 (N_13206,N_12331,N_12762);
nor U13207 (N_13207,N_12490,N_12351);
nor U13208 (N_13208,N_12598,N_12121);
nand U13209 (N_13209,N_12327,N_12929);
and U13210 (N_13210,N_12686,N_12038);
or U13211 (N_13211,N_12398,N_12283);
nand U13212 (N_13212,N_12114,N_12760);
nand U13213 (N_13213,N_12599,N_12493);
or U13214 (N_13214,N_12358,N_12581);
and U13215 (N_13215,N_12776,N_12062);
xor U13216 (N_13216,N_12951,N_12221);
xnor U13217 (N_13217,N_12175,N_12909);
or U13218 (N_13218,N_12812,N_12468);
xor U13219 (N_13219,N_12043,N_12210);
and U13220 (N_13220,N_12340,N_12824);
nand U13221 (N_13221,N_12200,N_12437);
and U13222 (N_13222,N_12347,N_12656);
xor U13223 (N_13223,N_12765,N_12015);
nor U13224 (N_13224,N_12878,N_12806);
or U13225 (N_13225,N_12274,N_12013);
nand U13226 (N_13226,N_12101,N_12509);
and U13227 (N_13227,N_12108,N_12787);
and U13228 (N_13228,N_12962,N_12780);
nor U13229 (N_13229,N_12685,N_12831);
nand U13230 (N_13230,N_12044,N_12671);
nor U13231 (N_13231,N_12965,N_12458);
nand U13232 (N_13232,N_12573,N_12915);
or U13233 (N_13233,N_12826,N_12595);
or U13234 (N_13234,N_12725,N_12326);
or U13235 (N_13235,N_12242,N_12057);
or U13236 (N_13236,N_12785,N_12334);
and U13237 (N_13237,N_12499,N_12539);
xor U13238 (N_13238,N_12997,N_12625);
nand U13239 (N_13239,N_12544,N_12166);
and U13240 (N_13240,N_12421,N_12455);
nand U13241 (N_13241,N_12619,N_12733);
or U13242 (N_13242,N_12703,N_12259);
nand U13243 (N_13243,N_12956,N_12174);
or U13244 (N_13244,N_12963,N_12764);
xnor U13245 (N_13245,N_12775,N_12285);
nand U13246 (N_13246,N_12624,N_12529);
nor U13247 (N_13247,N_12228,N_12129);
or U13248 (N_13248,N_12654,N_12017);
and U13249 (N_13249,N_12171,N_12172);
and U13250 (N_13250,N_12999,N_12628);
xnor U13251 (N_13251,N_12254,N_12823);
xnor U13252 (N_13252,N_12561,N_12080);
nor U13253 (N_13253,N_12902,N_12604);
nand U13254 (N_13254,N_12303,N_12184);
nand U13255 (N_13255,N_12699,N_12548);
nor U13256 (N_13256,N_12387,N_12112);
nand U13257 (N_13257,N_12741,N_12676);
or U13258 (N_13258,N_12975,N_12151);
nand U13259 (N_13259,N_12637,N_12928);
or U13260 (N_13260,N_12005,N_12991);
or U13261 (N_13261,N_12070,N_12600);
or U13262 (N_13262,N_12375,N_12461);
nand U13263 (N_13263,N_12472,N_12049);
and U13264 (N_13264,N_12423,N_12324);
or U13265 (N_13265,N_12863,N_12211);
nand U13266 (N_13266,N_12404,N_12865);
nand U13267 (N_13267,N_12425,N_12246);
nand U13268 (N_13268,N_12328,N_12978);
nand U13269 (N_13269,N_12004,N_12723);
or U13270 (N_13270,N_12546,N_12109);
nor U13271 (N_13271,N_12220,N_12033);
and U13272 (N_13272,N_12457,N_12169);
and U13273 (N_13273,N_12275,N_12098);
nand U13274 (N_13274,N_12125,N_12397);
xor U13275 (N_13275,N_12689,N_12215);
or U13276 (N_13276,N_12282,N_12456);
nor U13277 (N_13277,N_12305,N_12803);
xor U13278 (N_13278,N_12068,N_12023);
and U13279 (N_13279,N_12696,N_12424);
or U13280 (N_13280,N_12463,N_12266);
nand U13281 (N_13281,N_12748,N_12156);
nand U13282 (N_13282,N_12811,N_12583);
and U13283 (N_13283,N_12554,N_12778);
nor U13284 (N_13284,N_12261,N_12717);
nor U13285 (N_13285,N_12610,N_12454);
or U13286 (N_13286,N_12721,N_12374);
nand U13287 (N_13287,N_12605,N_12413);
nand U13288 (N_13288,N_12050,N_12994);
nand U13289 (N_13289,N_12477,N_12880);
or U13290 (N_13290,N_12576,N_12466);
nand U13291 (N_13291,N_12148,N_12631);
or U13292 (N_13292,N_12827,N_12411);
nand U13293 (N_13293,N_12908,N_12460);
nor U13294 (N_13294,N_12480,N_12578);
or U13295 (N_13295,N_12433,N_12574);
nand U13296 (N_13296,N_12896,N_12913);
nand U13297 (N_13297,N_12740,N_12032);
nor U13298 (N_13298,N_12392,N_12638);
or U13299 (N_13299,N_12575,N_12688);
nor U13300 (N_13300,N_12867,N_12154);
xor U13301 (N_13301,N_12319,N_12052);
and U13302 (N_13302,N_12567,N_12025);
and U13303 (N_13303,N_12924,N_12552);
and U13304 (N_13304,N_12907,N_12064);
xor U13305 (N_13305,N_12633,N_12217);
nor U13306 (N_13306,N_12828,N_12926);
nor U13307 (N_13307,N_12482,N_12713);
nor U13308 (N_13308,N_12382,N_12781);
and U13309 (N_13309,N_12912,N_12732);
nor U13310 (N_13310,N_12979,N_12223);
and U13311 (N_13311,N_12592,N_12609);
or U13312 (N_13312,N_12443,N_12520);
and U13313 (N_13313,N_12407,N_12712);
and U13314 (N_13314,N_12856,N_12872);
nand U13315 (N_13315,N_12307,N_12127);
nand U13316 (N_13316,N_12749,N_12833);
and U13317 (N_13317,N_12585,N_12658);
or U13318 (N_13318,N_12716,N_12814);
and U13319 (N_13319,N_12030,N_12296);
xnor U13320 (N_13320,N_12024,N_12968);
nor U13321 (N_13321,N_12697,N_12524);
xor U13322 (N_13322,N_12168,N_12889);
nor U13323 (N_13323,N_12420,N_12584);
and U13324 (N_13324,N_12728,N_12708);
and U13325 (N_13325,N_12874,N_12191);
nand U13326 (N_13326,N_12026,N_12178);
and U13327 (N_13327,N_12082,N_12559);
and U13328 (N_13328,N_12953,N_12791);
and U13329 (N_13329,N_12588,N_12465);
xnor U13330 (N_13330,N_12996,N_12416);
or U13331 (N_13331,N_12507,N_12731);
nand U13332 (N_13332,N_12395,N_12194);
nand U13333 (N_13333,N_12818,N_12116);
and U13334 (N_13334,N_12403,N_12864);
and U13335 (N_13335,N_12060,N_12517);
nand U13336 (N_13336,N_12257,N_12140);
xnor U13337 (N_13337,N_12891,N_12187);
or U13338 (N_13338,N_12798,N_12447);
nand U13339 (N_13339,N_12957,N_12591);
nor U13340 (N_13340,N_12142,N_12948);
and U13341 (N_13341,N_12901,N_12110);
nand U13342 (N_13342,N_12557,N_12680);
nand U13343 (N_13343,N_12342,N_12825);
and U13344 (N_13344,N_12964,N_12730);
nand U13345 (N_13345,N_12854,N_12453);
and U13346 (N_13346,N_12474,N_12332);
nor U13347 (N_13347,N_12014,N_12815);
nor U13348 (N_13348,N_12415,N_12855);
nor U13349 (N_13349,N_12646,N_12077);
and U13350 (N_13350,N_12095,N_12304);
nor U13351 (N_13351,N_12008,N_12903);
and U13352 (N_13352,N_12219,N_12291);
and U13353 (N_13353,N_12396,N_12119);
nor U13354 (N_13354,N_12945,N_12813);
xor U13355 (N_13355,N_12278,N_12054);
or U13356 (N_13356,N_12073,N_12434);
nor U13357 (N_13357,N_12944,N_12316);
xor U13358 (N_13358,N_12028,N_12720);
nor U13359 (N_13359,N_12756,N_12715);
or U13360 (N_13360,N_12487,N_12675);
or U13361 (N_13361,N_12003,N_12653);
or U13362 (N_13362,N_12501,N_12281);
xor U13363 (N_13363,N_12504,N_12218);
and U13364 (N_13364,N_12701,N_12203);
and U13365 (N_13365,N_12422,N_12180);
or U13366 (N_13366,N_12543,N_12792);
nand U13367 (N_13367,N_12170,N_12719);
xor U13368 (N_13368,N_12666,N_12526);
and U13369 (N_13369,N_12237,N_12808);
nor U13370 (N_13370,N_12897,N_12384);
nand U13371 (N_13371,N_12037,N_12767);
nor U13372 (N_13372,N_12105,N_12263);
or U13373 (N_13373,N_12226,N_12059);
or U13374 (N_13374,N_12231,N_12850);
and U13375 (N_13375,N_12039,N_12829);
nor U13376 (N_13376,N_12177,N_12809);
nand U13377 (N_13377,N_12943,N_12162);
nor U13378 (N_13378,N_12911,N_12113);
and U13379 (N_13379,N_12866,N_12273);
or U13380 (N_13380,N_12632,N_12547);
or U13381 (N_13381,N_12734,N_12485);
or U13382 (N_13382,N_12312,N_12742);
nor U13383 (N_13383,N_12763,N_12208);
and U13384 (N_13384,N_12971,N_12819);
nor U13385 (N_13385,N_12885,N_12970);
nor U13386 (N_13386,N_12418,N_12093);
nor U13387 (N_13387,N_12213,N_12364);
or U13388 (N_13388,N_12128,N_12367);
and U13389 (N_13389,N_12146,N_12556);
xor U13390 (N_13390,N_12810,N_12040);
nand U13391 (N_13391,N_12503,N_12494);
xor U13392 (N_13392,N_12914,N_12497);
xor U13393 (N_13393,N_12558,N_12341);
xnor U13394 (N_13394,N_12984,N_12959);
or U13395 (N_13395,N_12502,N_12353);
nand U13396 (N_13396,N_12345,N_12389);
nor U13397 (N_13397,N_12603,N_12354);
nor U13398 (N_13398,N_12270,N_12264);
nor U13399 (N_13399,N_12564,N_12150);
or U13400 (N_13400,N_12694,N_12954);
nor U13401 (N_13401,N_12918,N_12649);
or U13402 (N_13402,N_12533,N_12650);
xor U13403 (N_13403,N_12079,N_12570);
nand U13404 (N_13404,N_12847,N_12029);
nor U13405 (N_13405,N_12104,N_12475);
or U13406 (N_13406,N_12406,N_12016);
nand U13407 (N_13407,N_12747,N_12643);
xnor U13408 (N_13408,N_12905,N_12280);
nand U13409 (N_13409,N_12790,N_12394);
or U13410 (N_13410,N_12381,N_12919);
nand U13411 (N_13411,N_12868,N_12530);
and U13412 (N_13412,N_12426,N_12617);
nor U13413 (N_13413,N_12670,N_12243);
or U13414 (N_13414,N_12783,N_12484);
or U13415 (N_13415,N_12597,N_12206);
xnor U13416 (N_13416,N_12009,N_12772);
nand U13417 (N_13417,N_12925,N_12440);
and U13418 (N_13418,N_12473,N_12369);
or U13419 (N_13419,N_12512,N_12227);
or U13420 (N_13420,N_12138,N_12590);
nor U13421 (N_13421,N_12636,N_12736);
or U13422 (N_13422,N_12986,N_12031);
xor U13423 (N_13423,N_12618,N_12391);
or U13424 (N_13424,N_12987,N_12973);
nand U13425 (N_13425,N_12754,N_12432);
or U13426 (N_13426,N_12007,N_12634);
and U13427 (N_13427,N_12679,N_12385);
or U13428 (N_13428,N_12684,N_12265);
nor U13429 (N_13429,N_12982,N_12167);
and U13430 (N_13430,N_12076,N_12816);
or U13431 (N_13431,N_12522,N_12066);
nand U13432 (N_13432,N_12955,N_12419);
or U13433 (N_13433,N_12934,N_12115);
nor U13434 (N_13434,N_12553,N_12941);
xnor U13435 (N_13435,N_12513,N_12309);
or U13436 (N_13436,N_12329,N_12239);
xnor U13437 (N_13437,N_12386,N_12702);
or U13438 (N_13438,N_12155,N_12188);
and U13439 (N_13439,N_12784,N_12122);
and U13440 (N_13440,N_12262,N_12489);
or U13441 (N_13441,N_12333,N_12212);
nand U13442 (N_13442,N_12536,N_12123);
nand U13443 (N_13443,N_12571,N_12107);
nor U13444 (N_13444,N_12000,N_12488);
or U13445 (N_13445,N_12593,N_12330);
or U13446 (N_13446,N_12892,N_12613);
xor U13447 (N_13447,N_12616,N_12240);
nor U13448 (N_13448,N_12894,N_12587);
nor U13449 (N_13449,N_12614,N_12626);
and U13450 (N_13450,N_12481,N_12376);
or U13451 (N_13451,N_12935,N_12299);
nor U13452 (N_13452,N_12229,N_12377);
nand U13453 (N_13453,N_12126,N_12335);
nor U13454 (N_13454,N_12222,N_12117);
and U13455 (N_13455,N_12667,N_12560);
nand U13456 (N_13456,N_12518,N_12189);
nand U13457 (N_13457,N_12898,N_12510);
nor U13458 (N_13458,N_12629,N_12035);
xor U13459 (N_13459,N_12276,N_12946);
xor U13460 (N_13460,N_12442,N_12366);
nand U13461 (N_13461,N_12247,N_12417);
and U13462 (N_13462,N_12102,N_12010);
and U13463 (N_13463,N_12735,N_12541);
nand U13464 (N_13464,N_12832,N_12606);
or U13465 (N_13465,N_12185,N_12446);
nor U13466 (N_13466,N_12916,N_12290);
and U13467 (N_13467,N_12704,N_12106);
nor U13468 (N_13468,N_12293,N_12234);
or U13469 (N_13469,N_12739,N_12921);
nand U13470 (N_13470,N_12565,N_12660);
and U13471 (N_13471,N_12621,N_12183);
nand U13472 (N_13472,N_12297,N_12190);
nand U13473 (N_13473,N_12857,N_12976);
or U13474 (N_13474,N_12900,N_12683);
nor U13475 (N_13475,N_12692,N_12308);
and U13476 (N_13476,N_12018,N_12136);
nor U13477 (N_13477,N_12192,N_12197);
nand U13478 (N_13478,N_12448,N_12758);
and U13479 (N_13479,N_12306,N_12950);
and U13480 (N_13480,N_12788,N_12786);
xor U13481 (N_13481,N_12705,N_12371);
nand U13482 (N_13482,N_12486,N_12176);
and U13483 (N_13483,N_12379,N_12540);
or U13484 (N_13484,N_12992,N_12910);
xor U13485 (N_13485,N_12450,N_12566);
or U13486 (N_13486,N_12428,N_12640);
xnor U13487 (N_13487,N_12436,N_12074);
or U13488 (N_13488,N_12528,N_12001);
xnor U13489 (N_13489,N_12664,N_12317);
nor U13490 (N_13490,N_12601,N_12002);
nor U13491 (N_13491,N_12006,N_12755);
xor U13492 (N_13492,N_12838,N_12173);
or U13493 (N_13493,N_12937,N_12302);
and U13494 (N_13494,N_12165,N_12400);
and U13495 (N_13495,N_12846,N_12204);
nand U13496 (N_13496,N_12589,N_12972);
or U13497 (N_13497,N_12444,N_12368);
and U13498 (N_13498,N_12886,N_12476);
nand U13499 (N_13499,N_12344,N_12056);
nand U13500 (N_13500,N_12023,N_12153);
or U13501 (N_13501,N_12053,N_12214);
nand U13502 (N_13502,N_12187,N_12260);
xnor U13503 (N_13503,N_12996,N_12776);
and U13504 (N_13504,N_12046,N_12157);
nand U13505 (N_13505,N_12095,N_12853);
nand U13506 (N_13506,N_12558,N_12592);
nand U13507 (N_13507,N_12302,N_12050);
nand U13508 (N_13508,N_12463,N_12202);
and U13509 (N_13509,N_12678,N_12358);
nand U13510 (N_13510,N_12847,N_12962);
nand U13511 (N_13511,N_12298,N_12965);
nand U13512 (N_13512,N_12043,N_12932);
and U13513 (N_13513,N_12608,N_12722);
or U13514 (N_13514,N_12021,N_12565);
xnor U13515 (N_13515,N_12364,N_12356);
nand U13516 (N_13516,N_12440,N_12866);
and U13517 (N_13517,N_12417,N_12630);
nor U13518 (N_13518,N_12650,N_12017);
nand U13519 (N_13519,N_12872,N_12280);
nor U13520 (N_13520,N_12266,N_12308);
nand U13521 (N_13521,N_12223,N_12509);
or U13522 (N_13522,N_12280,N_12698);
nor U13523 (N_13523,N_12700,N_12478);
nor U13524 (N_13524,N_12969,N_12081);
or U13525 (N_13525,N_12260,N_12079);
nand U13526 (N_13526,N_12292,N_12470);
or U13527 (N_13527,N_12742,N_12031);
or U13528 (N_13528,N_12777,N_12525);
or U13529 (N_13529,N_12608,N_12619);
and U13530 (N_13530,N_12102,N_12550);
or U13531 (N_13531,N_12289,N_12054);
nor U13532 (N_13532,N_12253,N_12447);
nor U13533 (N_13533,N_12629,N_12404);
or U13534 (N_13534,N_12113,N_12094);
or U13535 (N_13535,N_12349,N_12487);
nor U13536 (N_13536,N_12844,N_12839);
nand U13537 (N_13537,N_12436,N_12866);
or U13538 (N_13538,N_12120,N_12725);
or U13539 (N_13539,N_12592,N_12372);
nor U13540 (N_13540,N_12579,N_12129);
nor U13541 (N_13541,N_12391,N_12686);
or U13542 (N_13542,N_12291,N_12241);
nand U13543 (N_13543,N_12877,N_12528);
or U13544 (N_13544,N_12563,N_12329);
or U13545 (N_13545,N_12121,N_12696);
and U13546 (N_13546,N_12233,N_12067);
and U13547 (N_13547,N_12981,N_12027);
nor U13548 (N_13548,N_12791,N_12812);
nand U13549 (N_13549,N_12824,N_12696);
nand U13550 (N_13550,N_12525,N_12249);
or U13551 (N_13551,N_12811,N_12130);
and U13552 (N_13552,N_12053,N_12778);
and U13553 (N_13553,N_12307,N_12045);
nand U13554 (N_13554,N_12737,N_12959);
and U13555 (N_13555,N_12786,N_12327);
nor U13556 (N_13556,N_12338,N_12503);
or U13557 (N_13557,N_12240,N_12894);
nor U13558 (N_13558,N_12079,N_12961);
nor U13559 (N_13559,N_12700,N_12300);
nor U13560 (N_13560,N_12190,N_12109);
nor U13561 (N_13561,N_12512,N_12991);
nor U13562 (N_13562,N_12018,N_12011);
nor U13563 (N_13563,N_12512,N_12901);
or U13564 (N_13564,N_12011,N_12465);
or U13565 (N_13565,N_12203,N_12143);
nand U13566 (N_13566,N_12879,N_12753);
nand U13567 (N_13567,N_12578,N_12446);
nand U13568 (N_13568,N_12617,N_12511);
nor U13569 (N_13569,N_12798,N_12863);
xnor U13570 (N_13570,N_12571,N_12656);
and U13571 (N_13571,N_12092,N_12483);
and U13572 (N_13572,N_12858,N_12738);
and U13573 (N_13573,N_12496,N_12175);
xor U13574 (N_13574,N_12012,N_12505);
and U13575 (N_13575,N_12415,N_12499);
and U13576 (N_13576,N_12817,N_12883);
nor U13577 (N_13577,N_12678,N_12339);
or U13578 (N_13578,N_12505,N_12572);
or U13579 (N_13579,N_12598,N_12569);
nor U13580 (N_13580,N_12727,N_12160);
nor U13581 (N_13581,N_12839,N_12064);
and U13582 (N_13582,N_12957,N_12349);
xor U13583 (N_13583,N_12149,N_12189);
nand U13584 (N_13584,N_12693,N_12782);
or U13585 (N_13585,N_12379,N_12279);
and U13586 (N_13586,N_12927,N_12237);
xor U13587 (N_13587,N_12047,N_12347);
nand U13588 (N_13588,N_12880,N_12853);
and U13589 (N_13589,N_12526,N_12472);
or U13590 (N_13590,N_12695,N_12239);
or U13591 (N_13591,N_12290,N_12758);
nand U13592 (N_13592,N_12489,N_12113);
and U13593 (N_13593,N_12487,N_12095);
nand U13594 (N_13594,N_12606,N_12224);
nand U13595 (N_13595,N_12179,N_12054);
xor U13596 (N_13596,N_12005,N_12326);
and U13597 (N_13597,N_12951,N_12427);
and U13598 (N_13598,N_12361,N_12952);
nor U13599 (N_13599,N_12300,N_12673);
nor U13600 (N_13600,N_12286,N_12052);
or U13601 (N_13601,N_12827,N_12700);
and U13602 (N_13602,N_12807,N_12330);
nand U13603 (N_13603,N_12682,N_12774);
nand U13604 (N_13604,N_12105,N_12102);
nand U13605 (N_13605,N_12943,N_12230);
nor U13606 (N_13606,N_12988,N_12039);
nor U13607 (N_13607,N_12540,N_12772);
and U13608 (N_13608,N_12995,N_12001);
and U13609 (N_13609,N_12840,N_12853);
and U13610 (N_13610,N_12967,N_12584);
xnor U13611 (N_13611,N_12513,N_12171);
and U13612 (N_13612,N_12968,N_12002);
and U13613 (N_13613,N_12318,N_12695);
and U13614 (N_13614,N_12876,N_12073);
or U13615 (N_13615,N_12736,N_12690);
or U13616 (N_13616,N_12222,N_12585);
nor U13617 (N_13617,N_12903,N_12359);
nor U13618 (N_13618,N_12827,N_12080);
nand U13619 (N_13619,N_12758,N_12249);
nand U13620 (N_13620,N_12392,N_12204);
and U13621 (N_13621,N_12092,N_12240);
and U13622 (N_13622,N_12002,N_12867);
nand U13623 (N_13623,N_12452,N_12769);
or U13624 (N_13624,N_12231,N_12422);
or U13625 (N_13625,N_12162,N_12095);
and U13626 (N_13626,N_12431,N_12851);
or U13627 (N_13627,N_12339,N_12664);
nand U13628 (N_13628,N_12899,N_12246);
or U13629 (N_13629,N_12973,N_12880);
nand U13630 (N_13630,N_12278,N_12875);
nand U13631 (N_13631,N_12874,N_12217);
and U13632 (N_13632,N_12235,N_12674);
nor U13633 (N_13633,N_12419,N_12178);
nor U13634 (N_13634,N_12612,N_12314);
nor U13635 (N_13635,N_12333,N_12930);
and U13636 (N_13636,N_12769,N_12009);
and U13637 (N_13637,N_12312,N_12875);
and U13638 (N_13638,N_12762,N_12619);
or U13639 (N_13639,N_12682,N_12770);
and U13640 (N_13640,N_12115,N_12656);
nor U13641 (N_13641,N_12386,N_12542);
nor U13642 (N_13642,N_12796,N_12106);
or U13643 (N_13643,N_12572,N_12879);
xor U13644 (N_13644,N_12869,N_12704);
nand U13645 (N_13645,N_12284,N_12571);
and U13646 (N_13646,N_12782,N_12623);
and U13647 (N_13647,N_12903,N_12194);
or U13648 (N_13648,N_12127,N_12242);
and U13649 (N_13649,N_12287,N_12948);
and U13650 (N_13650,N_12204,N_12327);
or U13651 (N_13651,N_12127,N_12258);
xor U13652 (N_13652,N_12430,N_12914);
and U13653 (N_13653,N_12249,N_12791);
or U13654 (N_13654,N_12021,N_12996);
nor U13655 (N_13655,N_12014,N_12901);
nor U13656 (N_13656,N_12714,N_12656);
nand U13657 (N_13657,N_12520,N_12118);
nor U13658 (N_13658,N_12776,N_12487);
nand U13659 (N_13659,N_12696,N_12689);
nand U13660 (N_13660,N_12275,N_12821);
xnor U13661 (N_13661,N_12795,N_12425);
and U13662 (N_13662,N_12894,N_12219);
nor U13663 (N_13663,N_12089,N_12161);
nor U13664 (N_13664,N_12788,N_12729);
nand U13665 (N_13665,N_12927,N_12565);
or U13666 (N_13666,N_12427,N_12481);
and U13667 (N_13667,N_12778,N_12434);
or U13668 (N_13668,N_12192,N_12375);
or U13669 (N_13669,N_12312,N_12722);
nor U13670 (N_13670,N_12798,N_12502);
and U13671 (N_13671,N_12143,N_12047);
or U13672 (N_13672,N_12903,N_12448);
nand U13673 (N_13673,N_12826,N_12381);
xor U13674 (N_13674,N_12444,N_12473);
nand U13675 (N_13675,N_12562,N_12679);
nand U13676 (N_13676,N_12078,N_12578);
or U13677 (N_13677,N_12969,N_12511);
nand U13678 (N_13678,N_12936,N_12916);
or U13679 (N_13679,N_12788,N_12395);
nand U13680 (N_13680,N_12090,N_12234);
and U13681 (N_13681,N_12648,N_12805);
or U13682 (N_13682,N_12525,N_12633);
or U13683 (N_13683,N_12938,N_12017);
nand U13684 (N_13684,N_12344,N_12025);
and U13685 (N_13685,N_12166,N_12267);
nor U13686 (N_13686,N_12856,N_12647);
or U13687 (N_13687,N_12795,N_12654);
and U13688 (N_13688,N_12481,N_12217);
nor U13689 (N_13689,N_12155,N_12579);
or U13690 (N_13690,N_12613,N_12279);
or U13691 (N_13691,N_12851,N_12592);
and U13692 (N_13692,N_12826,N_12648);
xnor U13693 (N_13693,N_12794,N_12002);
xor U13694 (N_13694,N_12775,N_12869);
and U13695 (N_13695,N_12693,N_12375);
or U13696 (N_13696,N_12540,N_12289);
or U13697 (N_13697,N_12306,N_12551);
nor U13698 (N_13698,N_12449,N_12989);
and U13699 (N_13699,N_12112,N_12984);
and U13700 (N_13700,N_12524,N_12559);
and U13701 (N_13701,N_12146,N_12023);
nor U13702 (N_13702,N_12210,N_12783);
nand U13703 (N_13703,N_12098,N_12862);
nand U13704 (N_13704,N_12797,N_12072);
xor U13705 (N_13705,N_12946,N_12138);
or U13706 (N_13706,N_12737,N_12537);
and U13707 (N_13707,N_12497,N_12749);
nand U13708 (N_13708,N_12878,N_12307);
nor U13709 (N_13709,N_12834,N_12343);
nand U13710 (N_13710,N_12484,N_12011);
and U13711 (N_13711,N_12800,N_12290);
xnor U13712 (N_13712,N_12244,N_12818);
and U13713 (N_13713,N_12851,N_12723);
or U13714 (N_13714,N_12449,N_12393);
and U13715 (N_13715,N_12286,N_12224);
and U13716 (N_13716,N_12948,N_12288);
nand U13717 (N_13717,N_12393,N_12737);
nor U13718 (N_13718,N_12509,N_12669);
nand U13719 (N_13719,N_12202,N_12459);
or U13720 (N_13720,N_12223,N_12872);
nor U13721 (N_13721,N_12809,N_12245);
xor U13722 (N_13722,N_12393,N_12707);
nand U13723 (N_13723,N_12203,N_12582);
nor U13724 (N_13724,N_12880,N_12734);
nor U13725 (N_13725,N_12486,N_12583);
or U13726 (N_13726,N_12213,N_12833);
or U13727 (N_13727,N_12748,N_12886);
nor U13728 (N_13728,N_12699,N_12011);
or U13729 (N_13729,N_12415,N_12733);
or U13730 (N_13730,N_12974,N_12715);
or U13731 (N_13731,N_12321,N_12522);
or U13732 (N_13732,N_12754,N_12745);
or U13733 (N_13733,N_12190,N_12293);
nand U13734 (N_13734,N_12400,N_12850);
nor U13735 (N_13735,N_12462,N_12697);
or U13736 (N_13736,N_12485,N_12935);
nand U13737 (N_13737,N_12287,N_12487);
xor U13738 (N_13738,N_12816,N_12571);
nor U13739 (N_13739,N_12234,N_12211);
nand U13740 (N_13740,N_12461,N_12464);
and U13741 (N_13741,N_12057,N_12104);
nand U13742 (N_13742,N_12071,N_12064);
nor U13743 (N_13743,N_12511,N_12169);
xor U13744 (N_13744,N_12146,N_12121);
nand U13745 (N_13745,N_12093,N_12519);
or U13746 (N_13746,N_12242,N_12028);
nand U13747 (N_13747,N_12268,N_12206);
nand U13748 (N_13748,N_12243,N_12689);
nand U13749 (N_13749,N_12816,N_12556);
nor U13750 (N_13750,N_12047,N_12997);
and U13751 (N_13751,N_12579,N_12701);
nand U13752 (N_13752,N_12759,N_12987);
nand U13753 (N_13753,N_12557,N_12814);
and U13754 (N_13754,N_12338,N_12086);
and U13755 (N_13755,N_12060,N_12881);
nor U13756 (N_13756,N_12849,N_12217);
or U13757 (N_13757,N_12397,N_12181);
or U13758 (N_13758,N_12921,N_12236);
nand U13759 (N_13759,N_12853,N_12394);
and U13760 (N_13760,N_12116,N_12642);
or U13761 (N_13761,N_12994,N_12865);
nor U13762 (N_13762,N_12224,N_12331);
nand U13763 (N_13763,N_12016,N_12849);
nor U13764 (N_13764,N_12903,N_12351);
nor U13765 (N_13765,N_12620,N_12919);
xnor U13766 (N_13766,N_12580,N_12358);
nor U13767 (N_13767,N_12499,N_12791);
nor U13768 (N_13768,N_12974,N_12580);
and U13769 (N_13769,N_12578,N_12888);
and U13770 (N_13770,N_12994,N_12532);
nor U13771 (N_13771,N_12610,N_12222);
nor U13772 (N_13772,N_12609,N_12398);
nor U13773 (N_13773,N_12949,N_12334);
xor U13774 (N_13774,N_12171,N_12577);
and U13775 (N_13775,N_12896,N_12751);
nor U13776 (N_13776,N_12401,N_12139);
or U13777 (N_13777,N_12581,N_12773);
nand U13778 (N_13778,N_12447,N_12530);
or U13779 (N_13779,N_12825,N_12324);
and U13780 (N_13780,N_12923,N_12357);
nor U13781 (N_13781,N_12429,N_12392);
nand U13782 (N_13782,N_12143,N_12137);
or U13783 (N_13783,N_12477,N_12837);
or U13784 (N_13784,N_12940,N_12514);
xnor U13785 (N_13785,N_12063,N_12631);
xor U13786 (N_13786,N_12974,N_12021);
or U13787 (N_13787,N_12029,N_12743);
xor U13788 (N_13788,N_12998,N_12383);
nor U13789 (N_13789,N_12232,N_12794);
nor U13790 (N_13790,N_12158,N_12250);
nor U13791 (N_13791,N_12643,N_12409);
xor U13792 (N_13792,N_12549,N_12274);
xnor U13793 (N_13793,N_12453,N_12930);
nand U13794 (N_13794,N_12058,N_12130);
or U13795 (N_13795,N_12651,N_12265);
xnor U13796 (N_13796,N_12577,N_12798);
nor U13797 (N_13797,N_12559,N_12411);
nand U13798 (N_13798,N_12592,N_12097);
nand U13799 (N_13799,N_12367,N_12805);
nand U13800 (N_13800,N_12029,N_12209);
xnor U13801 (N_13801,N_12233,N_12366);
and U13802 (N_13802,N_12790,N_12562);
nand U13803 (N_13803,N_12305,N_12490);
and U13804 (N_13804,N_12760,N_12983);
and U13805 (N_13805,N_12953,N_12673);
nor U13806 (N_13806,N_12078,N_12651);
nand U13807 (N_13807,N_12169,N_12707);
nor U13808 (N_13808,N_12976,N_12750);
and U13809 (N_13809,N_12304,N_12194);
or U13810 (N_13810,N_12899,N_12664);
or U13811 (N_13811,N_12713,N_12606);
nand U13812 (N_13812,N_12572,N_12100);
nand U13813 (N_13813,N_12594,N_12434);
or U13814 (N_13814,N_12058,N_12225);
or U13815 (N_13815,N_12471,N_12947);
or U13816 (N_13816,N_12066,N_12377);
nor U13817 (N_13817,N_12849,N_12526);
and U13818 (N_13818,N_12231,N_12879);
and U13819 (N_13819,N_12684,N_12755);
or U13820 (N_13820,N_12928,N_12271);
xnor U13821 (N_13821,N_12773,N_12746);
nor U13822 (N_13822,N_12563,N_12166);
and U13823 (N_13823,N_12817,N_12502);
xor U13824 (N_13824,N_12089,N_12309);
xor U13825 (N_13825,N_12430,N_12346);
or U13826 (N_13826,N_12384,N_12232);
and U13827 (N_13827,N_12859,N_12581);
nand U13828 (N_13828,N_12348,N_12848);
or U13829 (N_13829,N_12959,N_12207);
nand U13830 (N_13830,N_12932,N_12624);
and U13831 (N_13831,N_12594,N_12174);
nand U13832 (N_13832,N_12168,N_12394);
and U13833 (N_13833,N_12146,N_12000);
and U13834 (N_13834,N_12379,N_12741);
xnor U13835 (N_13835,N_12523,N_12705);
or U13836 (N_13836,N_12197,N_12713);
xnor U13837 (N_13837,N_12091,N_12988);
or U13838 (N_13838,N_12503,N_12403);
and U13839 (N_13839,N_12106,N_12175);
nand U13840 (N_13840,N_12688,N_12988);
nand U13841 (N_13841,N_12749,N_12745);
nor U13842 (N_13842,N_12354,N_12760);
or U13843 (N_13843,N_12349,N_12533);
or U13844 (N_13844,N_12912,N_12725);
xor U13845 (N_13845,N_12228,N_12022);
and U13846 (N_13846,N_12710,N_12136);
nor U13847 (N_13847,N_12080,N_12093);
nand U13848 (N_13848,N_12940,N_12889);
nor U13849 (N_13849,N_12839,N_12364);
nand U13850 (N_13850,N_12567,N_12983);
and U13851 (N_13851,N_12073,N_12123);
nand U13852 (N_13852,N_12755,N_12711);
and U13853 (N_13853,N_12739,N_12745);
nand U13854 (N_13854,N_12174,N_12069);
nor U13855 (N_13855,N_12160,N_12387);
nor U13856 (N_13856,N_12082,N_12976);
nor U13857 (N_13857,N_12480,N_12581);
or U13858 (N_13858,N_12183,N_12585);
nor U13859 (N_13859,N_12556,N_12545);
nand U13860 (N_13860,N_12047,N_12394);
or U13861 (N_13861,N_12980,N_12891);
nor U13862 (N_13862,N_12520,N_12155);
nor U13863 (N_13863,N_12329,N_12364);
and U13864 (N_13864,N_12716,N_12494);
xor U13865 (N_13865,N_12532,N_12318);
and U13866 (N_13866,N_12648,N_12300);
nand U13867 (N_13867,N_12261,N_12502);
and U13868 (N_13868,N_12797,N_12860);
nor U13869 (N_13869,N_12628,N_12224);
and U13870 (N_13870,N_12480,N_12279);
nor U13871 (N_13871,N_12935,N_12388);
xor U13872 (N_13872,N_12832,N_12919);
nand U13873 (N_13873,N_12668,N_12022);
nand U13874 (N_13874,N_12529,N_12411);
nor U13875 (N_13875,N_12153,N_12760);
or U13876 (N_13876,N_12967,N_12949);
xnor U13877 (N_13877,N_12338,N_12301);
nor U13878 (N_13878,N_12084,N_12935);
or U13879 (N_13879,N_12001,N_12025);
nor U13880 (N_13880,N_12957,N_12533);
or U13881 (N_13881,N_12322,N_12085);
nand U13882 (N_13882,N_12798,N_12864);
xor U13883 (N_13883,N_12111,N_12641);
nand U13884 (N_13884,N_12012,N_12588);
nand U13885 (N_13885,N_12333,N_12944);
nand U13886 (N_13886,N_12484,N_12444);
and U13887 (N_13887,N_12750,N_12690);
xor U13888 (N_13888,N_12583,N_12130);
and U13889 (N_13889,N_12220,N_12448);
nor U13890 (N_13890,N_12678,N_12418);
and U13891 (N_13891,N_12555,N_12468);
nor U13892 (N_13892,N_12332,N_12276);
or U13893 (N_13893,N_12854,N_12867);
and U13894 (N_13894,N_12392,N_12379);
nor U13895 (N_13895,N_12982,N_12451);
and U13896 (N_13896,N_12733,N_12549);
or U13897 (N_13897,N_12469,N_12244);
nor U13898 (N_13898,N_12940,N_12950);
nand U13899 (N_13899,N_12568,N_12022);
xor U13900 (N_13900,N_12509,N_12923);
and U13901 (N_13901,N_12531,N_12250);
or U13902 (N_13902,N_12599,N_12502);
xor U13903 (N_13903,N_12006,N_12183);
and U13904 (N_13904,N_12342,N_12412);
or U13905 (N_13905,N_12778,N_12873);
nand U13906 (N_13906,N_12842,N_12641);
nand U13907 (N_13907,N_12282,N_12320);
nand U13908 (N_13908,N_12688,N_12331);
nor U13909 (N_13909,N_12801,N_12341);
nor U13910 (N_13910,N_12092,N_12501);
nand U13911 (N_13911,N_12853,N_12448);
nor U13912 (N_13912,N_12877,N_12050);
and U13913 (N_13913,N_12308,N_12286);
nand U13914 (N_13914,N_12421,N_12526);
nor U13915 (N_13915,N_12811,N_12545);
and U13916 (N_13916,N_12388,N_12134);
or U13917 (N_13917,N_12623,N_12967);
xnor U13918 (N_13918,N_12987,N_12441);
nand U13919 (N_13919,N_12000,N_12370);
nand U13920 (N_13920,N_12128,N_12255);
or U13921 (N_13921,N_12464,N_12245);
nor U13922 (N_13922,N_12469,N_12537);
or U13923 (N_13923,N_12449,N_12527);
and U13924 (N_13924,N_12726,N_12853);
xor U13925 (N_13925,N_12744,N_12612);
or U13926 (N_13926,N_12601,N_12667);
nor U13927 (N_13927,N_12793,N_12054);
nor U13928 (N_13928,N_12109,N_12907);
or U13929 (N_13929,N_12612,N_12257);
nor U13930 (N_13930,N_12970,N_12597);
nor U13931 (N_13931,N_12193,N_12723);
nand U13932 (N_13932,N_12079,N_12534);
nor U13933 (N_13933,N_12098,N_12730);
nand U13934 (N_13934,N_12246,N_12800);
or U13935 (N_13935,N_12231,N_12712);
or U13936 (N_13936,N_12000,N_12722);
nor U13937 (N_13937,N_12269,N_12601);
or U13938 (N_13938,N_12807,N_12958);
nor U13939 (N_13939,N_12613,N_12103);
and U13940 (N_13940,N_12361,N_12258);
nand U13941 (N_13941,N_12748,N_12166);
nand U13942 (N_13942,N_12403,N_12558);
nand U13943 (N_13943,N_12162,N_12946);
or U13944 (N_13944,N_12213,N_12505);
and U13945 (N_13945,N_12258,N_12546);
or U13946 (N_13946,N_12926,N_12905);
or U13947 (N_13947,N_12445,N_12945);
nor U13948 (N_13948,N_12369,N_12658);
and U13949 (N_13949,N_12914,N_12354);
nand U13950 (N_13950,N_12268,N_12375);
or U13951 (N_13951,N_12966,N_12792);
or U13952 (N_13952,N_12806,N_12672);
xor U13953 (N_13953,N_12587,N_12691);
or U13954 (N_13954,N_12354,N_12763);
nor U13955 (N_13955,N_12771,N_12370);
and U13956 (N_13956,N_12947,N_12514);
xor U13957 (N_13957,N_12263,N_12163);
nor U13958 (N_13958,N_12281,N_12324);
nor U13959 (N_13959,N_12684,N_12162);
nand U13960 (N_13960,N_12904,N_12737);
nor U13961 (N_13961,N_12667,N_12959);
xor U13962 (N_13962,N_12578,N_12979);
nor U13963 (N_13963,N_12799,N_12052);
and U13964 (N_13964,N_12944,N_12871);
nand U13965 (N_13965,N_12637,N_12504);
nand U13966 (N_13966,N_12006,N_12074);
and U13967 (N_13967,N_12648,N_12524);
nor U13968 (N_13968,N_12308,N_12700);
nand U13969 (N_13969,N_12506,N_12524);
and U13970 (N_13970,N_12262,N_12931);
or U13971 (N_13971,N_12304,N_12810);
xnor U13972 (N_13972,N_12177,N_12778);
nor U13973 (N_13973,N_12493,N_12086);
and U13974 (N_13974,N_12644,N_12381);
or U13975 (N_13975,N_12289,N_12136);
and U13976 (N_13976,N_12410,N_12514);
or U13977 (N_13977,N_12656,N_12058);
nor U13978 (N_13978,N_12983,N_12978);
and U13979 (N_13979,N_12359,N_12657);
nand U13980 (N_13980,N_12000,N_12884);
or U13981 (N_13981,N_12270,N_12575);
or U13982 (N_13982,N_12535,N_12204);
nor U13983 (N_13983,N_12843,N_12166);
nor U13984 (N_13984,N_12153,N_12692);
or U13985 (N_13985,N_12506,N_12320);
and U13986 (N_13986,N_12404,N_12709);
nand U13987 (N_13987,N_12908,N_12288);
nand U13988 (N_13988,N_12802,N_12651);
nand U13989 (N_13989,N_12135,N_12588);
or U13990 (N_13990,N_12819,N_12630);
xor U13991 (N_13991,N_12464,N_12646);
nor U13992 (N_13992,N_12505,N_12035);
xnor U13993 (N_13993,N_12877,N_12183);
and U13994 (N_13994,N_12204,N_12988);
xnor U13995 (N_13995,N_12829,N_12203);
nor U13996 (N_13996,N_12419,N_12525);
or U13997 (N_13997,N_12872,N_12980);
and U13998 (N_13998,N_12171,N_12498);
nor U13999 (N_13999,N_12376,N_12746);
and U14000 (N_14000,N_13809,N_13907);
nand U14001 (N_14001,N_13670,N_13377);
nand U14002 (N_14002,N_13689,N_13880);
or U14003 (N_14003,N_13889,N_13634);
and U14004 (N_14004,N_13112,N_13373);
nor U14005 (N_14005,N_13939,N_13938);
nor U14006 (N_14006,N_13335,N_13448);
nand U14007 (N_14007,N_13769,N_13862);
nor U14008 (N_14008,N_13339,N_13606);
nand U14009 (N_14009,N_13585,N_13187);
or U14010 (N_14010,N_13516,N_13416);
xnor U14011 (N_14011,N_13561,N_13831);
or U14012 (N_14012,N_13249,N_13099);
and U14013 (N_14013,N_13386,N_13613);
or U14014 (N_14014,N_13124,N_13009);
and U14015 (N_14015,N_13289,N_13847);
and U14016 (N_14016,N_13250,N_13379);
nor U14017 (N_14017,N_13559,N_13288);
or U14018 (N_14018,N_13533,N_13669);
and U14019 (N_14019,N_13956,N_13801);
and U14020 (N_14020,N_13624,N_13403);
nor U14021 (N_14021,N_13142,N_13216);
nand U14022 (N_14022,N_13678,N_13025);
and U14023 (N_14023,N_13190,N_13159);
xnor U14024 (N_14024,N_13193,N_13055);
nor U14025 (N_14025,N_13942,N_13444);
nand U14026 (N_14026,N_13401,N_13426);
nor U14027 (N_14027,N_13034,N_13465);
or U14028 (N_14028,N_13572,N_13825);
or U14029 (N_14029,N_13716,N_13684);
or U14030 (N_14030,N_13368,N_13970);
or U14031 (N_14031,N_13863,N_13798);
and U14032 (N_14032,N_13109,N_13525);
and U14033 (N_14033,N_13311,N_13214);
or U14034 (N_14034,N_13361,N_13421);
nor U14035 (N_14035,N_13419,N_13677);
or U14036 (N_14036,N_13095,N_13537);
or U14037 (N_14037,N_13207,N_13692);
nor U14038 (N_14038,N_13732,N_13553);
nand U14039 (N_14039,N_13005,N_13481);
and U14040 (N_14040,N_13261,N_13902);
nand U14041 (N_14041,N_13567,N_13340);
or U14042 (N_14042,N_13500,N_13474);
or U14043 (N_14043,N_13449,N_13594);
nand U14044 (N_14044,N_13351,N_13700);
nor U14045 (N_14045,N_13575,N_13138);
nor U14046 (N_14046,N_13222,N_13768);
and U14047 (N_14047,N_13355,N_13713);
nor U14048 (N_14048,N_13735,N_13948);
or U14049 (N_14049,N_13484,N_13274);
and U14050 (N_14050,N_13196,N_13223);
or U14051 (N_14051,N_13758,N_13996);
or U14052 (N_14052,N_13369,N_13746);
nand U14053 (N_14053,N_13599,N_13165);
or U14054 (N_14054,N_13062,N_13727);
nand U14055 (N_14055,N_13084,N_13934);
xor U14056 (N_14056,N_13856,N_13330);
nor U14057 (N_14057,N_13304,N_13579);
nor U14058 (N_14058,N_13649,N_13944);
or U14059 (N_14059,N_13263,N_13707);
or U14060 (N_14060,N_13621,N_13359);
or U14061 (N_14061,N_13155,N_13991);
and U14062 (N_14062,N_13558,N_13935);
xnor U14063 (N_14063,N_13008,N_13059);
and U14064 (N_14064,N_13329,N_13682);
xnor U14065 (N_14065,N_13845,N_13246);
nor U14066 (N_14066,N_13676,N_13331);
and U14067 (N_14067,N_13745,N_13589);
and U14068 (N_14068,N_13919,N_13975);
or U14069 (N_14069,N_13770,N_13276);
nand U14070 (N_14070,N_13116,N_13305);
and U14071 (N_14071,N_13296,N_13799);
or U14072 (N_14072,N_13367,N_13595);
nor U14073 (N_14073,N_13945,N_13573);
and U14074 (N_14074,N_13076,N_13097);
and U14075 (N_14075,N_13171,N_13683);
nor U14076 (N_14076,N_13679,N_13393);
nand U14077 (N_14077,N_13480,N_13236);
and U14078 (N_14078,N_13588,N_13774);
or U14079 (N_14079,N_13545,N_13904);
nor U14080 (N_14080,N_13178,N_13168);
xor U14081 (N_14081,N_13779,N_13378);
and U14082 (N_14082,N_13805,N_13362);
nand U14083 (N_14083,N_13139,N_13674);
and U14084 (N_14084,N_13734,N_13217);
or U14085 (N_14085,N_13836,N_13583);
and U14086 (N_14086,N_13892,N_13953);
or U14087 (N_14087,N_13645,N_13255);
nor U14088 (N_14088,N_13875,N_13894);
and U14089 (N_14089,N_13166,N_13636);
nand U14090 (N_14090,N_13722,N_13611);
nor U14091 (N_14091,N_13463,N_13952);
nand U14092 (N_14092,N_13495,N_13219);
and U14093 (N_14093,N_13389,N_13253);
xor U14094 (N_14094,N_13134,N_13812);
nand U14095 (N_14095,N_13024,N_13663);
and U14096 (N_14096,N_13597,N_13036);
nand U14097 (N_14097,N_13307,N_13642);
and U14098 (N_14098,N_13900,N_13681);
or U14099 (N_14099,N_13915,N_13056);
nand U14100 (N_14100,N_13789,N_13264);
nor U14101 (N_14101,N_13917,N_13065);
and U14102 (N_14102,N_13306,N_13404);
and U14103 (N_14103,N_13167,N_13327);
and U14104 (N_14104,N_13666,N_13273);
and U14105 (N_14105,N_13882,N_13612);
or U14106 (N_14106,N_13365,N_13826);
nor U14107 (N_14107,N_13643,N_13494);
nor U14108 (N_14108,N_13651,N_13865);
and U14109 (N_14109,N_13529,N_13506);
xnor U14110 (N_14110,N_13020,N_13081);
and U14111 (N_14111,N_13800,N_13936);
or U14112 (N_14112,N_13511,N_13164);
and U14113 (N_14113,N_13225,N_13502);
nor U14114 (N_14114,N_13456,N_13728);
or U14115 (N_14115,N_13272,N_13245);
xnor U14116 (N_14116,N_13408,N_13292);
xor U14117 (N_14117,N_13980,N_13156);
and U14118 (N_14118,N_13177,N_13091);
and U14119 (N_14119,N_13406,N_13487);
nor U14120 (N_14120,N_13507,N_13132);
nand U14121 (N_14121,N_13834,N_13792);
nand U14122 (N_14122,N_13280,N_13411);
and U14123 (N_14123,N_13927,N_13957);
and U14124 (N_14124,N_13647,N_13937);
nand U14125 (N_14125,N_13392,N_13780);
nand U14126 (N_14126,N_13230,N_13822);
or U14127 (N_14127,N_13041,N_13173);
nand U14128 (N_14128,N_13486,N_13547);
or U14129 (N_14129,N_13371,N_13194);
nand U14130 (N_14130,N_13775,N_13299);
nand U14131 (N_14131,N_13120,N_13382);
and U14132 (N_14132,N_13424,N_13873);
nor U14133 (N_14133,N_13777,N_13069);
nor U14134 (N_14134,N_13538,N_13748);
or U14135 (N_14135,N_13323,N_13951);
nor U14136 (N_14136,N_13283,N_13357);
nand U14137 (N_14137,N_13137,N_13765);
nor U14138 (N_14138,N_13557,N_13428);
or U14139 (N_14139,N_13201,N_13491);
or U14140 (N_14140,N_13560,N_13662);
or U14141 (N_14141,N_13910,N_13600);
or U14142 (N_14142,N_13787,N_13628);
or U14143 (N_14143,N_13224,N_13657);
and U14144 (N_14144,N_13539,N_13268);
nor U14145 (N_14145,N_13893,N_13535);
nor U14146 (N_14146,N_13554,N_13923);
xor U14147 (N_14147,N_13072,N_13672);
nor U14148 (N_14148,N_13012,N_13832);
nor U14149 (N_14149,N_13520,N_13314);
or U14150 (N_14150,N_13218,N_13860);
and U14151 (N_14151,N_13650,N_13309);
or U14152 (N_14152,N_13644,N_13531);
or U14153 (N_14153,N_13696,N_13269);
nand U14154 (N_14154,N_13198,N_13442);
or U14155 (N_14155,N_13417,N_13852);
or U14156 (N_14156,N_13047,N_13969);
xnor U14157 (N_14157,N_13631,N_13067);
nand U14158 (N_14158,N_13958,N_13383);
nor U14159 (N_14159,N_13586,N_13267);
or U14160 (N_14160,N_13011,N_13083);
and U14161 (N_14161,N_13629,N_13429);
or U14162 (N_14162,N_13790,N_13452);
nor U14163 (N_14163,N_13234,N_13914);
and U14164 (N_14164,N_13850,N_13740);
and U14165 (N_14165,N_13710,N_13615);
xnor U14166 (N_14166,N_13046,N_13211);
nor U14167 (N_14167,N_13374,N_13764);
or U14168 (N_14168,N_13755,N_13861);
nand U14169 (N_14169,N_13431,N_13568);
or U14170 (N_14170,N_13625,N_13455);
or U14171 (N_14171,N_13782,N_13473);
nand U14172 (N_14172,N_13685,N_13133);
or U14173 (N_14173,N_13648,N_13400);
or U14174 (N_14174,N_13318,N_13415);
and U14175 (N_14175,N_13310,N_13375);
nor U14176 (N_14176,N_13381,N_13576);
or U14177 (N_14177,N_13844,N_13496);
nand U14178 (N_14178,N_13736,N_13867);
nor U14179 (N_14179,N_13313,N_13719);
and U14180 (N_14180,N_13571,N_13089);
nand U14181 (N_14181,N_13227,N_13503);
xor U14182 (N_14182,N_13675,N_13590);
nor U14183 (N_14183,N_13086,N_13646);
and U14184 (N_14184,N_13848,N_13891);
nand U14185 (N_14185,N_13752,N_13698);
or U14186 (N_14186,N_13427,N_13810);
or U14187 (N_14187,N_13665,N_13453);
and U14188 (N_14188,N_13301,N_13121);
nand U14189 (N_14189,N_13048,N_13353);
nand U14190 (N_14190,N_13058,N_13163);
nor U14191 (N_14191,N_13475,N_13932);
nand U14192 (N_14192,N_13906,N_13260);
or U14193 (N_14193,N_13610,N_13818);
nand U14194 (N_14194,N_13738,N_13001);
nand U14195 (N_14195,N_13410,N_13434);
nand U14196 (N_14196,N_13930,N_13045);
nor U14197 (N_14197,N_13857,N_13877);
nand U14198 (N_14198,N_13580,N_13528);
and U14199 (N_14199,N_13360,N_13023);
nor U14200 (N_14200,N_13987,N_13786);
and U14201 (N_14201,N_13108,N_13690);
nor U14202 (N_14202,N_13989,N_13941);
nand U14203 (N_14203,N_13796,N_13823);
or U14204 (N_14204,N_13243,N_13785);
nor U14205 (N_14205,N_13843,N_13140);
xor U14206 (N_14206,N_13115,N_13551);
nor U14207 (N_14207,N_13947,N_13215);
nand U14208 (N_14208,N_13791,N_13043);
and U14209 (N_14209,N_13897,N_13440);
or U14210 (N_14210,N_13596,N_13467);
xnor U14211 (N_14211,N_13051,N_13184);
and U14212 (N_14212,N_13524,N_13688);
nor U14213 (N_14213,N_13985,N_13354);
nand U14214 (N_14214,N_13117,N_13704);
or U14215 (N_14215,N_13721,N_13497);
nand U14216 (N_14216,N_13074,N_13298);
nand U14217 (N_14217,N_13813,N_13839);
xnor U14218 (N_14218,N_13820,N_13441);
xor U14219 (N_14219,N_13639,N_13518);
and U14220 (N_14220,N_13909,N_13622);
nand U14221 (N_14221,N_13443,N_13986);
nand U14222 (N_14222,N_13447,N_13652);
or U14223 (N_14223,N_13438,N_13271);
and U14224 (N_14224,N_13181,N_13835);
xor U14225 (N_14225,N_13244,N_13235);
nand U14226 (N_14226,N_13995,N_13238);
or U14227 (N_14227,N_13584,N_13922);
or U14228 (N_14228,N_13127,N_13686);
nor U14229 (N_14229,N_13854,N_13064);
nor U14230 (N_14230,N_13912,N_13326);
xnor U14231 (N_14231,N_13285,N_13028);
or U14232 (N_14232,N_13101,N_13756);
nand U14233 (N_14233,N_13931,N_13691);
and U14234 (N_14234,N_13437,N_13398);
and U14235 (N_14235,N_13007,N_13717);
and U14236 (N_14236,N_13469,N_13035);
and U14237 (N_14237,N_13290,N_13933);
xnor U14238 (N_14238,N_13080,N_13037);
nor U14239 (N_14239,N_13226,N_13213);
xor U14240 (N_14240,N_13982,N_13180);
nand U14241 (N_14241,N_13352,N_13436);
xor U14242 (N_14242,N_13057,N_13546);
nor U14243 (N_14243,N_13508,N_13103);
and U14244 (N_14244,N_13004,N_13630);
and U14245 (N_14245,N_13967,N_13366);
and U14246 (N_14246,N_13702,N_13370);
nor U14247 (N_14247,N_13905,N_13804);
and U14248 (N_14248,N_13961,N_13940);
and U14249 (N_14249,N_13040,N_13087);
nand U14250 (N_14250,N_13794,N_13760);
and U14251 (N_14251,N_13693,N_13846);
and U14252 (N_14252,N_13345,N_13018);
and U14253 (N_14253,N_13485,N_13966);
or U14254 (N_14254,N_13618,N_13153);
and U14255 (N_14255,N_13191,N_13974);
and U14256 (N_14256,N_13499,N_13432);
nor U14257 (N_14257,N_13021,N_13154);
nand U14258 (N_14258,N_13212,N_13459);
or U14259 (N_14259,N_13993,N_13100);
xnor U14260 (N_14260,N_13827,N_13013);
nor U14261 (N_14261,N_13252,N_13152);
nand U14262 (N_14262,N_13478,N_13536);
and U14263 (N_14263,N_13385,N_13281);
nor U14264 (N_14264,N_13162,N_13141);
nand U14265 (N_14265,N_13916,N_13924);
and U14266 (N_14266,N_13270,N_13476);
or U14267 (N_14267,N_13075,N_13256);
and U14268 (N_14268,N_13092,N_13349);
nand U14269 (N_14269,N_13188,N_13482);
nor U14270 (N_14270,N_13587,N_13189);
or U14271 (N_14271,N_13414,N_13853);
nand U14272 (N_14272,N_13753,N_13921);
nand U14273 (N_14273,N_13413,N_13635);
nand U14274 (N_14274,N_13763,N_13284);
or U14275 (N_14275,N_13896,N_13471);
xor U14276 (N_14276,N_13322,N_13556);
and U14277 (N_14277,N_13457,N_13706);
or U14278 (N_14278,N_13808,N_13607);
nand U14279 (N_14279,N_13718,N_13241);
nand U14280 (N_14280,N_13422,N_13347);
nor U14281 (N_14281,N_13185,N_13015);
nor U14282 (N_14282,N_13202,N_13807);
nand U14283 (N_14283,N_13602,N_13870);
nor U14284 (N_14284,N_13883,N_13821);
and U14285 (N_14285,N_13510,N_13811);
or U14286 (N_14286,N_13391,N_13170);
nor U14287 (N_14287,N_13950,N_13376);
nor U14288 (N_14288,N_13237,N_13477);
and U14289 (N_14289,N_13614,N_13145);
and U14290 (N_14290,N_13161,N_13498);
nand U14291 (N_14291,N_13550,N_13562);
nor U14292 (N_14292,N_13963,N_13275);
nor U14293 (N_14293,N_13955,N_13293);
xor U14294 (N_14294,N_13078,N_13439);
or U14295 (N_14295,N_13123,N_13715);
or U14296 (N_14296,N_13183,N_13016);
or U14297 (N_14297,N_13819,N_13501);
or U14298 (N_14298,N_13131,N_13460);
nand U14299 (N_14299,N_13454,N_13694);
and U14300 (N_14300,N_13527,N_13726);
or U14301 (N_14301,N_13402,N_13458);
or U14302 (N_14302,N_13129,N_13490);
xnor U14303 (N_14303,N_13027,N_13879);
nand U14304 (N_14304,N_13797,N_13130);
nand U14305 (N_14305,N_13751,N_13147);
xor U14306 (N_14306,N_13747,N_13061);
nor U14307 (N_14307,N_13543,N_13981);
xor U14308 (N_14308,N_13781,N_13592);
nand U14309 (N_14309,N_13344,N_13795);
and U14310 (N_14310,N_13569,N_13017);
and U14311 (N_14311,N_13977,N_13638);
nand U14312 (N_14312,N_13988,N_13591);
nor U14313 (N_14313,N_13363,N_13701);
or U14314 (N_14314,N_13332,N_13603);
nand U14315 (N_14315,N_13971,N_13829);
or U14316 (N_14316,N_13070,N_13898);
nand U14317 (N_14317,N_13493,N_13492);
or U14318 (N_14318,N_13451,N_13783);
or U14319 (N_14319,N_13540,N_13895);
and U14320 (N_14320,N_13549,N_13890);
nand U14321 (N_14321,N_13157,N_13817);
and U14322 (N_14322,N_13287,N_13384);
xnor U14323 (N_14323,N_13343,N_13090);
nand U14324 (N_14324,N_13888,N_13869);
or U14325 (N_14325,N_13654,N_13815);
nand U14326 (N_14326,N_13205,N_13548);
xnor U14327 (N_14327,N_13208,N_13578);
or U14328 (N_14328,N_13514,N_13342);
nand U14329 (N_14329,N_13144,N_13899);
and U14330 (N_14330,N_13802,N_13876);
xor U14331 (N_14331,N_13029,N_13723);
and U14332 (N_14332,N_13151,N_13731);
nor U14333 (N_14333,N_13446,N_13623);
or U14334 (N_14334,N_13570,N_13259);
nor U14335 (N_14335,N_13824,N_13000);
xnor U14336 (N_14336,N_13965,N_13350);
nand U14337 (N_14337,N_13228,N_13122);
and U14338 (N_14338,N_13049,N_13976);
or U14339 (N_14339,N_13978,N_13240);
nor U14340 (N_14340,N_13302,N_13082);
nand U14341 (N_14341,N_13433,N_13461);
and U14342 (N_14342,N_13866,N_13220);
and U14343 (N_14343,N_13757,N_13042);
and U14344 (N_14344,N_13929,N_13999);
or U14345 (N_14345,N_13641,N_13405);
nor U14346 (N_14346,N_13113,N_13574);
nand U14347 (N_14347,N_13088,N_13052);
nor U14348 (N_14348,N_13946,N_13338);
and U14349 (N_14349,N_13660,N_13601);
and U14350 (N_14350,N_13534,N_13172);
or U14351 (N_14351,N_13324,N_13544);
and U14352 (N_14352,N_13039,N_13632);
or U14353 (N_14353,N_13759,N_13872);
and U14354 (N_14354,N_13593,N_13388);
nor U14355 (N_14355,N_13730,N_13530);
and U14356 (N_14356,N_13068,N_13054);
and U14357 (N_14357,N_13192,N_13864);
nor U14358 (N_14358,N_13488,N_13356);
or U14359 (N_14359,N_13149,N_13766);
or U14360 (N_14360,N_13640,N_13093);
nor U14361 (N_14361,N_13773,N_13229);
nor U14362 (N_14362,N_13334,N_13725);
or U14363 (N_14363,N_13221,N_13003);
nor U14364 (N_14364,N_13328,N_13282);
or U14365 (N_14365,N_13291,N_13085);
nand U14366 (N_14366,N_13908,N_13239);
or U14367 (N_14367,N_13771,N_13364);
and U14368 (N_14368,N_13541,N_13175);
and U14369 (N_14369,N_13489,N_13526);
and U14370 (N_14370,N_13079,N_13680);
nor U14371 (N_14371,N_13949,N_13992);
xor U14372 (N_14372,N_13146,N_13118);
or U14373 (N_14373,N_13729,N_13317);
nor U14374 (N_14374,N_13136,N_13742);
or U14375 (N_14375,N_13918,N_13295);
nor U14376 (N_14376,N_13203,N_13582);
and U14377 (N_14377,N_13210,N_13430);
or U14378 (N_14378,N_13712,N_13960);
nor U14379 (N_14379,N_13814,N_13412);
nand U14380 (N_14380,N_13656,N_13668);
nor U14381 (N_14381,N_13911,N_13390);
or U14382 (N_14382,N_13744,N_13903);
and U14383 (N_14383,N_13828,N_13248);
nor U14384 (N_14384,N_13855,N_13697);
nor U14385 (N_14385,N_13671,N_13687);
nand U14386 (N_14386,N_13337,N_13784);
nand U14387 (N_14387,N_13445,N_13581);
nand U14388 (N_14388,N_13504,N_13659);
or U14389 (N_14389,N_13022,N_13286);
or U14390 (N_14390,N_13886,N_13830);
xnor U14391 (N_14391,N_13470,N_13619);
nand U14392 (N_14392,N_13566,N_13479);
and U14393 (N_14393,N_13653,N_13655);
or U14394 (N_14394,N_13358,N_13110);
or U14395 (N_14395,N_13407,N_13232);
or U14396 (N_14396,N_13251,N_13954);
and U14397 (N_14397,N_13160,N_13257);
or U14398 (N_14398,N_13014,N_13920);
nor U14399 (N_14399,N_13038,N_13994);
and U14400 (N_14400,N_13928,N_13703);
nand U14401 (N_14401,N_13754,N_13626);
xor U14402 (N_14402,N_13277,N_13209);
nor U14403 (N_14403,N_13107,N_13564);
or U14404 (N_14404,N_13032,N_13925);
nand U14405 (N_14405,N_13519,N_13464);
nor U14406 (N_14406,N_13833,N_13341);
xnor U14407 (N_14407,N_13066,N_13604);
xnor U14408 (N_14408,N_13266,N_13840);
or U14409 (N_14409,N_13767,N_13523);
xnor U14410 (N_14410,N_13724,N_13803);
or U14411 (N_14411,N_13838,N_13319);
or U14412 (N_14412,N_13750,N_13968);
nor U14413 (N_14413,N_13472,N_13204);
or U14414 (N_14414,N_13265,N_13806);
and U14415 (N_14415,N_13709,N_13399);
nand U14416 (N_14416,N_13174,N_13577);
nand U14417 (N_14417,N_13565,N_13901);
nor U14418 (N_14418,N_13387,N_13114);
nand U14419 (N_14419,N_13658,N_13073);
nand U14420 (N_14420,N_13699,N_13466);
and U14421 (N_14421,N_13943,N_13150);
and U14422 (N_14422,N_13044,N_13837);
or U14423 (N_14423,N_13515,N_13125);
or U14424 (N_14424,N_13315,N_13695);
and U14425 (N_14425,N_13336,N_13435);
and U14426 (N_14426,N_13321,N_13885);
nor U14427 (N_14427,N_13409,N_13262);
nor U14428 (N_14428,N_13031,N_13094);
or U14429 (N_14429,N_13111,N_13871);
and U14430 (N_14430,N_13851,N_13617);
nor U14431 (N_14431,N_13984,N_13608);
xnor U14432 (N_14432,N_13002,N_13868);
xor U14433 (N_14433,N_13661,N_13542);
nand U14434 (N_14434,N_13395,N_13998);
nor U14435 (N_14435,N_13605,N_13522);
and U14436 (N_14436,N_13096,N_13749);
and U14437 (N_14437,N_13010,N_13788);
or U14438 (N_14438,N_13997,N_13926);
nor U14439 (N_14439,N_13616,N_13521);
xnor U14440 (N_14440,N_13552,N_13761);
nor U14441 (N_14441,N_13849,N_13294);
or U14442 (N_14442,N_13633,N_13555);
or U14443 (N_14443,N_13913,N_13881);
nor U14444 (N_14444,N_13513,N_13962);
xor U14445 (N_14445,N_13316,N_13667);
xnor U14446 (N_14446,N_13148,N_13199);
and U14447 (N_14447,N_13026,N_13483);
nand U14448 (N_14448,N_13098,N_13418);
or U14449 (N_14449,N_13019,N_13972);
and U14450 (N_14450,N_13664,N_13609);
nand U14451 (N_14451,N_13673,N_13637);
nor U14452 (N_14452,N_13179,N_13517);
nand U14453 (N_14453,N_13380,N_13197);
xnor U14454 (N_14454,N_13119,N_13762);
xor U14455 (N_14455,N_13816,N_13104);
nor U14456 (N_14456,N_13303,N_13006);
nand U14457 (N_14457,N_13887,N_13060);
and U14458 (N_14458,N_13397,N_13102);
nor U14459 (N_14459,N_13512,N_13308);
nor U14460 (N_14460,N_13983,N_13973);
nand U14461 (N_14461,N_13776,N_13053);
or U14462 (N_14462,N_13105,N_13186);
and U14463 (N_14463,N_13563,N_13206);
nor U14464 (N_14464,N_13705,N_13325);
or U14465 (N_14465,N_13106,N_13396);
or U14466 (N_14466,N_13462,N_13964);
nand U14467 (N_14467,N_13297,N_13312);
and U14468 (N_14468,N_13050,N_13135);
and U14469 (N_14469,N_13420,N_13195);
xnor U14470 (N_14470,N_13346,N_13841);
or U14471 (N_14471,N_13884,N_13077);
nor U14472 (N_14472,N_13033,N_13200);
and U14473 (N_14473,N_13468,N_13030);
and U14474 (N_14474,N_13279,N_13242);
xnor U14475 (N_14475,N_13532,N_13143);
or U14476 (N_14476,N_13505,N_13450);
nand U14477 (N_14477,N_13627,N_13737);
or U14478 (N_14478,N_13509,N_13300);
and U14479 (N_14479,N_13254,N_13258);
nand U14480 (N_14480,N_13182,N_13071);
nand U14481 (N_14481,N_13741,N_13394);
nor U14482 (N_14482,N_13423,N_13169);
nand U14483 (N_14483,N_13720,N_13714);
nand U14484 (N_14484,N_13959,N_13425);
or U14485 (N_14485,N_13158,N_13842);
or U14486 (N_14486,N_13063,N_13320);
or U14487 (N_14487,N_13778,N_13247);
xor U14488 (N_14488,N_13878,N_13739);
nand U14489 (N_14489,N_13278,N_13372);
or U14490 (N_14490,N_13874,N_13859);
nor U14491 (N_14491,N_13333,N_13711);
xnor U14492 (N_14492,N_13176,N_13990);
nor U14493 (N_14493,N_13979,N_13858);
nand U14494 (N_14494,N_13743,N_13620);
nand U14495 (N_14495,N_13708,N_13793);
and U14496 (N_14496,N_13128,N_13772);
nor U14497 (N_14497,N_13233,N_13598);
and U14498 (N_14498,N_13348,N_13126);
and U14499 (N_14499,N_13733,N_13231);
or U14500 (N_14500,N_13095,N_13622);
or U14501 (N_14501,N_13753,N_13017);
and U14502 (N_14502,N_13110,N_13450);
or U14503 (N_14503,N_13016,N_13920);
and U14504 (N_14504,N_13022,N_13297);
nand U14505 (N_14505,N_13652,N_13395);
nand U14506 (N_14506,N_13107,N_13706);
or U14507 (N_14507,N_13374,N_13779);
xor U14508 (N_14508,N_13998,N_13769);
or U14509 (N_14509,N_13527,N_13878);
xnor U14510 (N_14510,N_13449,N_13986);
nor U14511 (N_14511,N_13213,N_13376);
and U14512 (N_14512,N_13443,N_13567);
or U14513 (N_14513,N_13317,N_13810);
nor U14514 (N_14514,N_13854,N_13918);
and U14515 (N_14515,N_13877,N_13830);
or U14516 (N_14516,N_13132,N_13494);
xnor U14517 (N_14517,N_13860,N_13782);
nand U14518 (N_14518,N_13742,N_13089);
or U14519 (N_14519,N_13007,N_13654);
nand U14520 (N_14520,N_13093,N_13548);
nand U14521 (N_14521,N_13100,N_13771);
or U14522 (N_14522,N_13407,N_13523);
nand U14523 (N_14523,N_13929,N_13294);
nor U14524 (N_14524,N_13510,N_13220);
and U14525 (N_14525,N_13024,N_13146);
and U14526 (N_14526,N_13861,N_13403);
or U14527 (N_14527,N_13491,N_13133);
or U14528 (N_14528,N_13028,N_13639);
or U14529 (N_14529,N_13358,N_13996);
nor U14530 (N_14530,N_13495,N_13287);
and U14531 (N_14531,N_13638,N_13254);
xor U14532 (N_14532,N_13958,N_13279);
nor U14533 (N_14533,N_13717,N_13028);
nand U14534 (N_14534,N_13695,N_13722);
and U14535 (N_14535,N_13548,N_13337);
nor U14536 (N_14536,N_13919,N_13619);
and U14537 (N_14537,N_13746,N_13641);
nand U14538 (N_14538,N_13893,N_13969);
and U14539 (N_14539,N_13259,N_13693);
nor U14540 (N_14540,N_13777,N_13034);
nand U14541 (N_14541,N_13021,N_13684);
nand U14542 (N_14542,N_13759,N_13342);
and U14543 (N_14543,N_13058,N_13100);
or U14544 (N_14544,N_13594,N_13171);
xor U14545 (N_14545,N_13048,N_13325);
and U14546 (N_14546,N_13785,N_13653);
and U14547 (N_14547,N_13102,N_13579);
or U14548 (N_14548,N_13221,N_13070);
and U14549 (N_14549,N_13360,N_13181);
or U14550 (N_14550,N_13900,N_13555);
or U14551 (N_14551,N_13791,N_13649);
or U14552 (N_14552,N_13024,N_13460);
nor U14553 (N_14553,N_13880,N_13441);
nand U14554 (N_14554,N_13765,N_13541);
nor U14555 (N_14555,N_13709,N_13746);
and U14556 (N_14556,N_13915,N_13597);
or U14557 (N_14557,N_13381,N_13813);
or U14558 (N_14558,N_13610,N_13462);
or U14559 (N_14559,N_13627,N_13390);
nand U14560 (N_14560,N_13987,N_13173);
nand U14561 (N_14561,N_13779,N_13859);
nand U14562 (N_14562,N_13789,N_13601);
nor U14563 (N_14563,N_13337,N_13021);
nand U14564 (N_14564,N_13161,N_13155);
nor U14565 (N_14565,N_13213,N_13589);
nand U14566 (N_14566,N_13153,N_13810);
and U14567 (N_14567,N_13268,N_13290);
or U14568 (N_14568,N_13185,N_13244);
nor U14569 (N_14569,N_13456,N_13921);
xor U14570 (N_14570,N_13312,N_13689);
or U14571 (N_14571,N_13349,N_13011);
or U14572 (N_14572,N_13065,N_13293);
nand U14573 (N_14573,N_13784,N_13296);
or U14574 (N_14574,N_13308,N_13692);
nor U14575 (N_14575,N_13342,N_13414);
nor U14576 (N_14576,N_13960,N_13560);
xor U14577 (N_14577,N_13773,N_13094);
or U14578 (N_14578,N_13016,N_13049);
nand U14579 (N_14579,N_13319,N_13218);
and U14580 (N_14580,N_13549,N_13105);
nand U14581 (N_14581,N_13358,N_13277);
nor U14582 (N_14582,N_13134,N_13998);
nor U14583 (N_14583,N_13739,N_13003);
and U14584 (N_14584,N_13279,N_13678);
and U14585 (N_14585,N_13025,N_13796);
and U14586 (N_14586,N_13915,N_13169);
xnor U14587 (N_14587,N_13871,N_13833);
and U14588 (N_14588,N_13242,N_13395);
and U14589 (N_14589,N_13986,N_13677);
nand U14590 (N_14590,N_13907,N_13364);
nand U14591 (N_14591,N_13410,N_13132);
nor U14592 (N_14592,N_13590,N_13827);
nor U14593 (N_14593,N_13375,N_13305);
nand U14594 (N_14594,N_13810,N_13177);
and U14595 (N_14595,N_13840,N_13036);
or U14596 (N_14596,N_13997,N_13486);
nand U14597 (N_14597,N_13243,N_13263);
nor U14598 (N_14598,N_13168,N_13434);
nand U14599 (N_14599,N_13252,N_13913);
nand U14600 (N_14600,N_13915,N_13032);
xnor U14601 (N_14601,N_13916,N_13500);
nand U14602 (N_14602,N_13155,N_13999);
or U14603 (N_14603,N_13389,N_13329);
nand U14604 (N_14604,N_13400,N_13307);
and U14605 (N_14605,N_13830,N_13696);
and U14606 (N_14606,N_13227,N_13363);
or U14607 (N_14607,N_13381,N_13638);
nor U14608 (N_14608,N_13886,N_13908);
or U14609 (N_14609,N_13270,N_13625);
nand U14610 (N_14610,N_13820,N_13910);
nand U14611 (N_14611,N_13618,N_13405);
nor U14612 (N_14612,N_13851,N_13296);
and U14613 (N_14613,N_13114,N_13883);
nand U14614 (N_14614,N_13483,N_13774);
and U14615 (N_14615,N_13970,N_13520);
nor U14616 (N_14616,N_13044,N_13473);
nand U14617 (N_14617,N_13908,N_13469);
nor U14618 (N_14618,N_13537,N_13784);
nor U14619 (N_14619,N_13439,N_13383);
nand U14620 (N_14620,N_13113,N_13070);
nor U14621 (N_14621,N_13794,N_13284);
or U14622 (N_14622,N_13956,N_13208);
xnor U14623 (N_14623,N_13966,N_13023);
and U14624 (N_14624,N_13847,N_13311);
nor U14625 (N_14625,N_13307,N_13335);
nor U14626 (N_14626,N_13567,N_13002);
and U14627 (N_14627,N_13791,N_13245);
nor U14628 (N_14628,N_13405,N_13503);
nand U14629 (N_14629,N_13471,N_13332);
and U14630 (N_14630,N_13357,N_13948);
or U14631 (N_14631,N_13731,N_13039);
nand U14632 (N_14632,N_13749,N_13775);
nand U14633 (N_14633,N_13205,N_13565);
nor U14634 (N_14634,N_13408,N_13067);
nand U14635 (N_14635,N_13014,N_13444);
and U14636 (N_14636,N_13308,N_13217);
and U14637 (N_14637,N_13689,N_13936);
or U14638 (N_14638,N_13639,N_13086);
or U14639 (N_14639,N_13872,N_13793);
or U14640 (N_14640,N_13182,N_13023);
and U14641 (N_14641,N_13306,N_13714);
or U14642 (N_14642,N_13347,N_13561);
and U14643 (N_14643,N_13235,N_13827);
nand U14644 (N_14644,N_13719,N_13738);
nand U14645 (N_14645,N_13329,N_13579);
nand U14646 (N_14646,N_13420,N_13066);
or U14647 (N_14647,N_13454,N_13965);
nor U14648 (N_14648,N_13500,N_13862);
or U14649 (N_14649,N_13090,N_13487);
nor U14650 (N_14650,N_13343,N_13977);
or U14651 (N_14651,N_13449,N_13959);
and U14652 (N_14652,N_13166,N_13711);
xnor U14653 (N_14653,N_13907,N_13827);
nand U14654 (N_14654,N_13314,N_13693);
xor U14655 (N_14655,N_13707,N_13712);
nor U14656 (N_14656,N_13604,N_13972);
nand U14657 (N_14657,N_13919,N_13652);
and U14658 (N_14658,N_13861,N_13683);
and U14659 (N_14659,N_13624,N_13096);
or U14660 (N_14660,N_13790,N_13812);
or U14661 (N_14661,N_13608,N_13083);
xor U14662 (N_14662,N_13153,N_13877);
nor U14663 (N_14663,N_13920,N_13624);
nor U14664 (N_14664,N_13843,N_13354);
nor U14665 (N_14665,N_13817,N_13343);
xnor U14666 (N_14666,N_13240,N_13825);
nand U14667 (N_14667,N_13180,N_13678);
and U14668 (N_14668,N_13809,N_13690);
and U14669 (N_14669,N_13540,N_13154);
nand U14670 (N_14670,N_13205,N_13074);
nor U14671 (N_14671,N_13256,N_13851);
and U14672 (N_14672,N_13636,N_13526);
or U14673 (N_14673,N_13812,N_13828);
and U14674 (N_14674,N_13946,N_13476);
nand U14675 (N_14675,N_13836,N_13638);
nor U14676 (N_14676,N_13962,N_13698);
or U14677 (N_14677,N_13727,N_13361);
and U14678 (N_14678,N_13944,N_13289);
or U14679 (N_14679,N_13424,N_13582);
nand U14680 (N_14680,N_13093,N_13260);
nor U14681 (N_14681,N_13458,N_13275);
nor U14682 (N_14682,N_13103,N_13327);
or U14683 (N_14683,N_13379,N_13493);
nor U14684 (N_14684,N_13130,N_13944);
or U14685 (N_14685,N_13120,N_13995);
nand U14686 (N_14686,N_13059,N_13307);
nor U14687 (N_14687,N_13033,N_13355);
or U14688 (N_14688,N_13687,N_13386);
and U14689 (N_14689,N_13275,N_13106);
xor U14690 (N_14690,N_13420,N_13159);
nand U14691 (N_14691,N_13655,N_13241);
nand U14692 (N_14692,N_13912,N_13701);
nor U14693 (N_14693,N_13498,N_13438);
nor U14694 (N_14694,N_13921,N_13106);
or U14695 (N_14695,N_13140,N_13313);
or U14696 (N_14696,N_13494,N_13249);
nor U14697 (N_14697,N_13537,N_13786);
xnor U14698 (N_14698,N_13079,N_13948);
nand U14699 (N_14699,N_13511,N_13915);
nand U14700 (N_14700,N_13532,N_13816);
nor U14701 (N_14701,N_13975,N_13457);
xnor U14702 (N_14702,N_13654,N_13241);
and U14703 (N_14703,N_13223,N_13662);
nor U14704 (N_14704,N_13457,N_13335);
and U14705 (N_14705,N_13494,N_13244);
nand U14706 (N_14706,N_13722,N_13861);
and U14707 (N_14707,N_13221,N_13562);
nor U14708 (N_14708,N_13129,N_13170);
nand U14709 (N_14709,N_13091,N_13740);
or U14710 (N_14710,N_13559,N_13177);
nand U14711 (N_14711,N_13093,N_13931);
or U14712 (N_14712,N_13758,N_13003);
and U14713 (N_14713,N_13576,N_13684);
and U14714 (N_14714,N_13286,N_13170);
nor U14715 (N_14715,N_13403,N_13119);
xor U14716 (N_14716,N_13789,N_13260);
and U14717 (N_14717,N_13310,N_13299);
xnor U14718 (N_14718,N_13308,N_13391);
nor U14719 (N_14719,N_13401,N_13446);
nor U14720 (N_14720,N_13575,N_13616);
nor U14721 (N_14721,N_13168,N_13396);
and U14722 (N_14722,N_13592,N_13568);
nor U14723 (N_14723,N_13134,N_13921);
nand U14724 (N_14724,N_13668,N_13269);
nand U14725 (N_14725,N_13817,N_13903);
nor U14726 (N_14726,N_13974,N_13057);
nor U14727 (N_14727,N_13896,N_13539);
nand U14728 (N_14728,N_13431,N_13987);
and U14729 (N_14729,N_13858,N_13778);
or U14730 (N_14730,N_13416,N_13212);
or U14731 (N_14731,N_13662,N_13887);
nand U14732 (N_14732,N_13077,N_13674);
xor U14733 (N_14733,N_13966,N_13723);
xnor U14734 (N_14734,N_13586,N_13890);
and U14735 (N_14735,N_13249,N_13280);
nor U14736 (N_14736,N_13649,N_13785);
xnor U14737 (N_14737,N_13122,N_13681);
nand U14738 (N_14738,N_13172,N_13987);
nand U14739 (N_14739,N_13979,N_13972);
nand U14740 (N_14740,N_13607,N_13878);
or U14741 (N_14741,N_13606,N_13977);
xor U14742 (N_14742,N_13796,N_13652);
and U14743 (N_14743,N_13690,N_13718);
nor U14744 (N_14744,N_13960,N_13943);
and U14745 (N_14745,N_13885,N_13886);
nand U14746 (N_14746,N_13603,N_13785);
nand U14747 (N_14747,N_13844,N_13296);
and U14748 (N_14748,N_13800,N_13281);
or U14749 (N_14749,N_13114,N_13680);
or U14750 (N_14750,N_13026,N_13357);
xor U14751 (N_14751,N_13575,N_13869);
xor U14752 (N_14752,N_13906,N_13064);
and U14753 (N_14753,N_13983,N_13853);
or U14754 (N_14754,N_13273,N_13932);
nand U14755 (N_14755,N_13263,N_13166);
nor U14756 (N_14756,N_13871,N_13682);
and U14757 (N_14757,N_13540,N_13763);
nor U14758 (N_14758,N_13694,N_13821);
or U14759 (N_14759,N_13541,N_13062);
and U14760 (N_14760,N_13802,N_13359);
nor U14761 (N_14761,N_13490,N_13518);
and U14762 (N_14762,N_13358,N_13278);
or U14763 (N_14763,N_13597,N_13703);
or U14764 (N_14764,N_13982,N_13845);
or U14765 (N_14765,N_13302,N_13538);
xnor U14766 (N_14766,N_13410,N_13832);
nor U14767 (N_14767,N_13654,N_13511);
xnor U14768 (N_14768,N_13226,N_13933);
nand U14769 (N_14769,N_13538,N_13655);
xor U14770 (N_14770,N_13357,N_13125);
or U14771 (N_14771,N_13646,N_13233);
or U14772 (N_14772,N_13263,N_13257);
nor U14773 (N_14773,N_13750,N_13360);
and U14774 (N_14774,N_13368,N_13450);
or U14775 (N_14775,N_13836,N_13075);
nor U14776 (N_14776,N_13850,N_13732);
nand U14777 (N_14777,N_13105,N_13062);
or U14778 (N_14778,N_13246,N_13235);
and U14779 (N_14779,N_13336,N_13805);
nor U14780 (N_14780,N_13616,N_13240);
nand U14781 (N_14781,N_13749,N_13795);
and U14782 (N_14782,N_13062,N_13299);
and U14783 (N_14783,N_13447,N_13075);
or U14784 (N_14784,N_13378,N_13362);
nand U14785 (N_14785,N_13137,N_13973);
nand U14786 (N_14786,N_13722,N_13583);
xnor U14787 (N_14787,N_13617,N_13089);
or U14788 (N_14788,N_13203,N_13569);
or U14789 (N_14789,N_13134,N_13975);
or U14790 (N_14790,N_13457,N_13471);
and U14791 (N_14791,N_13782,N_13623);
and U14792 (N_14792,N_13843,N_13799);
or U14793 (N_14793,N_13469,N_13543);
nor U14794 (N_14794,N_13004,N_13717);
xor U14795 (N_14795,N_13111,N_13669);
or U14796 (N_14796,N_13145,N_13143);
nand U14797 (N_14797,N_13048,N_13072);
nand U14798 (N_14798,N_13906,N_13494);
or U14799 (N_14799,N_13762,N_13554);
nor U14800 (N_14800,N_13467,N_13584);
and U14801 (N_14801,N_13130,N_13662);
or U14802 (N_14802,N_13870,N_13111);
and U14803 (N_14803,N_13510,N_13972);
nor U14804 (N_14804,N_13088,N_13909);
nor U14805 (N_14805,N_13535,N_13082);
nor U14806 (N_14806,N_13153,N_13048);
or U14807 (N_14807,N_13439,N_13792);
or U14808 (N_14808,N_13706,N_13517);
xor U14809 (N_14809,N_13709,N_13942);
nor U14810 (N_14810,N_13137,N_13609);
nor U14811 (N_14811,N_13963,N_13113);
or U14812 (N_14812,N_13583,N_13522);
or U14813 (N_14813,N_13532,N_13724);
nand U14814 (N_14814,N_13461,N_13189);
nand U14815 (N_14815,N_13850,N_13155);
nor U14816 (N_14816,N_13311,N_13131);
nand U14817 (N_14817,N_13643,N_13958);
or U14818 (N_14818,N_13012,N_13077);
nand U14819 (N_14819,N_13204,N_13153);
nor U14820 (N_14820,N_13123,N_13563);
nor U14821 (N_14821,N_13687,N_13358);
and U14822 (N_14822,N_13340,N_13755);
nor U14823 (N_14823,N_13977,N_13530);
xnor U14824 (N_14824,N_13709,N_13886);
nand U14825 (N_14825,N_13871,N_13916);
and U14826 (N_14826,N_13442,N_13459);
nor U14827 (N_14827,N_13310,N_13714);
and U14828 (N_14828,N_13133,N_13608);
nand U14829 (N_14829,N_13025,N_13827);
or U14830 (N_14830,N_13150,N_13780);
and U14831 (N_14831,N_13917,N_13056);
or U14832 (N_14832,N_13787,N_13054);
nor U14833 (N_14833,N_13097,N_13883);
xor U14834 (N_14834,N_13479,N_13319);
or U14835 (N_14835,N_13871,N_13551);
nand U14836 (N_14836,N_13533,N_13778);
nand U14837 (N_14837,N_13803,N_13368);
and U14838 (N_14838,N_13175,N_13032);
nor U14839 (N_14839,N_13808,N_13157);
nor U14840 (N_14840,N_13583,N_13729);
and U14841 (N_14841,N_13229,N_13732);
and U14842 (N_14842,N_13025,N_13051);
and U14843 (N_14843,N_13259,N_13289);
nor U14844 (N_14844,N_13610,N_13112);
xor U14845 (N_14845,N_13389,N_13279);
nor U14846 (N_14846,N_13586,N_13507);
xnor U14847 (N_14847,N_13092,N_13999);
nor U14848 (N_14848,N_13192,N_13332);
nor U14849 (N_14849,N_13904,N_13668);
nand U14850 (N_14850,N_13932,N_13239);
or U14851 (N_14851,N_13808,N_13948);
nor U14852 (N_14852,N_13075,N_13403);
and U14853 (N_14853,N_13308,N_13239);
nand U14854 (N_14854,N_13459,N_13104);
or U14855 (N_14855,N_13773,N_13364);
nor U14856 (N_14856,N_13973,N_13014);
and U14857 (N_14857,N_13292,N_13265);
nor U14858 (N_14858,N_13191,N_13450);
nand U14859 (N_14859,N_13542,N_13716);
nand U14860 (N_14860,N_13702,N_13190);
nor U14861 (N_14861,N_13612,N_13409);
nand U14862 (N_14862,N_13028,N_13136);
nand U14863 (N_14863,N_13796,N_13511);
nand U14864 (N_14864,N_13516,N_13602);
and U14865 (N_14865,N_13736,N_13202);
nor U14866 (N_14866,N_13968,N_13811);
or U14867 (N_14867,N_13043,N_13137);
nand U14868 (N_14868,N_13901,N_13135);
nor U14869 (N_14869,N_13468,N_13315);
or U14870 (N_14870,N_13798,N_13919);
or U14871 (N_14871,N_13513,N_13582);
and U14872 (N_14872,N_13257,N_13663);
nand U14873 (N_14873,N_13391,N_13253);
nand U14874 (N_14874,N_13176,N_13302);
nand U14875 (N_14875,N_13831,N_13839);
or U14876 (N_14876,N_13256,N_13444);
or U14877 (N_14877,N_13828,N_13410);
and U14878 (N_14878,N_13185,N_13914);
nand U14879 (N_14879,N_13871,N_13679);
nor U14880 (N_14880,N_13058,N_13916);
or U14881 (N_14881,N_13561,N_13732);
nand U14882 (N_14882,N_13284,N_13872);
nand U14883 (N_14883,N_13079,N_13900);
nor U14884 (N_14884,N_13544,N_13883);
or U14885 (N_14885,N_13625,N_13104);
nand U14886 (N_14886,N_13093,N_13516);
or U14887 (N_14887,N_13400,N_13082);
xnor U14888 (N_14888,N_13546,N_13397);
nand U14889 (N_14889,N_13109,N_13950);
nor U14890 (N_14890,N_13808,N_13419);
nand U14891 (N_14891,N_13675,N_13164);
nand U14892 (N_14892,N_13835,N_13212);
xor U14893 (N_14893,N_13319,N_13357);
nand U14894 (N_14894,N_13390,N_13689);
or U14895 (N_14895,N_13909,N_13351);
or U14896 (N_14896,N_13772,N_13424);
nand U14897 (N_14897,N_13411,N_13900);
xnor U14898 (N_14898,N_13930,N_13667);
and U14899 (N_14899,N_13370,N_13794);
nor U14900 (N_14900,N_13626,N_13638);
xnor U14901 (N_14901,N_13294,N_13302);
nor U14902 (N_14902,N_13641,N_13837);
and U14903 (N_14903,N_13984,N_13300);
xor U14904 (N_14904,N_13008,N_13814);
and U14905 (N_14905,N_13853,N_13499);
nor U14906 (N_14906,N_13440,N_13745);
nand U14907 (N_14907,N_13769,N_13957);
nand U14908 (N_14908,N_13079,N_13015);
or U14909 (N_14909,N_13743,N_13591);
nand U14910 (N_14910,N_13256,N_13144);
or U14911 (N_14911,N_13312,N_13302);
and U14912 (N_14912,N_13615,N_13985);
and U14913 (N_14913,N_13083,N_13230);
nor U14914 (N_14914,N_13507,N_13985);
or U14915 (N_14915,N_13816,N_13334);
nor U14916 (N_14916,N_13121,N_13311);
or U14917 (N_14917,N_13997,N_13689);
and U14918 (N_14918,N_13335,N_13430);
and U14919 (N_14919,N_13141,N_13082);
or U14920 (N_14920,N_13607,N_13215);
xnor U14921 (N_14921,N_13988,N_13789);
and U14922 (N_14922,N_13851,N_13459);
nand U14923 (N_14923,N_13892,N_13244);
xnor U14924 (N_14924,N_13043,N_13069);
and U14925 (N_14925,N_13876,N_13277);
or U14926 (N_14926,N_13834,N_13312);
nand U14927 (N_14927,N_13326,N_13492);
nor U14928 (N_14928,N_13991,N_13305);
or U14929 (N_14929,N_13722,N_13985);
and U14930 (N_14930,N_13663,N_13701);
and U14931 (N_14931,N_13619,N_13544);
nand U14932 (N_14932,N_13907,N_13746);
and U14933 (N_14933,N_13674,N_13525);
and U14934 (N_14934,N_13699,N_13558);
xnor U14935 (N_14935,N_13641,N_13379);
or U14936 (N_14936,N_13300,N_13862);
and U14937 (N_14937,N_13117,N_13884);
or U14938 (N_14938,N_13707,N_13332);
nor U14939 (N_14939,N_13186,N_13157);
nand U14940 (N_14940,N_13504,N_13400);
nor U14941 (N_14941,N_13549,N_13278);
xor U14942 (N_14942,N_13312,N_13057);
or U14943 (N_14943,N_13767,N_13764);
and U14944 (N_14944,N_13644,N_13961);
or U14945 (N_14945,N_13854,N_13219);
or U14946 (N_14946,N_13555,N_13559);
nand U14947 (N_14947,N_13521,N_13635);
nor U14948 (N_14948,N_13268,N_13679);
nand U14949 (N_14949,N_13294,N_13626);
and U14950 (N_14950,N_13374,N_13106);
nor U14951 (N_14951,N_13246,N_13048);
and U14952 (N_14952,N_13788,N_13580);
and U14953 (N_14953,N_13098,N_13266);
and U14954 (N_14954,N_13526,N_13225);
and U14955 (N_14955,N_13024,N_13561);
and U14956 (N_14956,N_13409,N_13903);
xnor U14957 (N_14957,N_13105,N_13191);
or U14958 (N_14958,N_13096,N_13097);
and U14959 (N_14959,N_13339,N_13822);
or U14960 (N_14960,N_13177,N_13084);
nand U14961 (N_14961,N_13229,N_13372);
and U14962 (N_14962,N_13462,N_13070);
nor U14963 (N_14963,N_13242,N_13516);
and U14964 (N_14964,N_13973,N_13958);
nand U14965 (N_14965,N_13564,N_13400);
nor U14966 (N_14966,N_13005,N_13170);
nand U14967 (N_14967,N_13260,N_13375);
nor U14968 (N_14968,N_13960,N_13450);
nand U14969 (N_14969,N_13319,N_13766);
xnor U14970 (N_14970,N_13179,N_13640);
and U14971 (N_14971,N_13260,N_13696);
nand U14972 (N_14972,N_13775,N_13059);
and U14973 (N_14973,N_13448,N_13609);
xnor U14974 (N_14974,N_13337,N_13485);
and U14975 (N_14975,N_13639,N_13926);
and U14976 (N_14976,N_13528,N_13418);
and U14977 (N_14977,N_13693,N_13591);
nand U14978 (N_14978,N_13286,N_13402);
and U14979 (N_14979,N_13727,N_13477);
or U14980 (N_14980,N_13643,N_13660);
or U14981 (N_14981,N_13895,N_13577);
nand U14982 (N_14982,N_13981,N_13149);
nand U14983 (N_14983,N_13402,N_13411);
nor U14984 (N_14984,N_13006,N_13134);
nand U14985 (N_14985,N_13793,N_13477);
nor U14986 (N_14986,N_13987,N_13363);
and U14987 (N_14987,N_13169,N_13681);
nand U14988 (N_14988,N_13808,N_13528);
or U14989 (N_14989,N_13895,N_13946);
or U14990 (N_14990,N_13894,N_13191);
nor U14991 (N_14991,N_13957,N_13345);
and U14992 (N_14992,N_13730,N_13969);
nand U14993 (N_14993,N_13522,N_13660);
nor U14994 (N_14994,N_13216,N_13176);
nand U14995 (N_14995,N_13191,N_13112);
nand U14996 (N_14996,N_13681,N_13932);
xnor U14997 (N_14997,N_13169,N_13898);
nor U14998 (N_14998,N_13922,N_13666);
and U14999 (N_14999,N_13953,N_13769);
xor UO_0 (O_0,N_14168,N_14545);
xnor UO_1 (O_1,N_14529,N_14247);
and UO_2 (O_2,N_14226,N_14124);
nor UO_3 (O_3,N_14570,N_14763);
and UO_4 (O_4,N_14645,N_14276);
or UO_5 (O_5,N_14634,N_14860);
nand UO_6 (O_6,N_14986,N_14602);
nor UO_7 (O_7,N_14130,N_14591);
or UO_8 (O_8,N_14918,N_14017);
nand UO_9 (O_9,N_14141,N_14428);
xnor UO_10 (O_10,N_14958,N_14354);
nand UO_11 (O_11,N_14207,N_14535);
nand UO_12 (O_12,N_14861,N_14619);
nor UO_13 (O_13,N_14352,N_14189);
or UO_14 (O_14,N_14974,N_14639);
and UO_15 (O_15,N_14195,N_14914);
or UO_16 (O_16,N_14801,N_14555);
nor UO_17 (O_17,N_14956,N_14922);
and UO_18 (O_18,N_14364,N_14016);
and UO_19 (O_19,N_14900,N_14253);
nand UO_20 (O_20,N_14393,N_14777);
or UO_21 (O_21,N_14912,N_14264);
xnor UO_22 (O_22,N_14669,N_14131);
nor UO_23 (O_23,N_14877,N_14950);
nor UO_24 (O_24,N_14427,N_14811);
and UO_25 (O_25,N_14710,N_14698);
nand UO_26 (O_26,N_14548,N_14625);
or UO_27 (O_27,N_14653,N_14337);
nor UO_28 (O_28,N_14030,N_14353);
nand UO_29 (O_29,N_14332,N_14758);
xor UO_30 (O_30,N_14411,N_14789);
and UO_31 (O_31,N_14584,N_14951);
nand UO_32 (O_32,N_14783,N_14971);
nand UO_33 (O_33,N_14129,N_14671);
or UO_34 (O_34,N_14288,N_14851);
or UO_35 (O_35,N_14357,N_14507);
or UO_36 (O_36,N_14641,N_14581);
nor UO_37 (O_37,N_14450,N_14659);
and UO_38 (O_38,N_14724,N_14178);
nor UO_39 (O_39,N_14980,N_14234);
nor UO_40 (O_40,N_14933,N_14681);
and UO_41 (O_41,N_14749,N_14240);
nor UO_42 (O_42,N_14533,N_14492);
nor UO_43 (O_43,N_14668,N_14314);
nand UO_44 (O_44,N_14819,N_14485);
nor UO_45 (O_45,N_14560,N_14887);
and UO_46 (O_46,N_14556,N_14365);
and UO_47 (O_47,N_14143,N_14344);
or UO_48 (O_48,N_14839,N_14519);
or UO_49 (O_49,N_14814,N_14932);
nand UO_50 (O_50,N_14330,N_14678);
nor UO_51 (O_51,N_14133,N_14685);
nand UO_52 (O_52,N_14417,N_14916);
or UO_53 (O_53,N_14559,N_14282);
and UO_54 (O_54,N_14132,N_14757);
nand UO_55 (O_55,N_14805,N_14707);
nor UO_56 (O_56,N_14847,N_14728);
or UO_57 (O_57,N_14984,N_14386);
nor UO_58 (O_58,N_14660,N_14487);
and UO_59 (O_59,N_14745,N_14292);
nand UO_60 (O_60,N_14670,N_14077);
and UO_61 (O_61,N_14173,N_14713);
and UO_62 (O_62,N_14488,N_14187);
nand UO_63 (O_63,N_14520,N_14009);
nor UO_64 (O_64,N_14667,N_14339);
and UO_65 (O_65,N_14246,N_14804);
nor UO_66 (O_66,N_14055,N_14585);
and UO_67 (O_67,N_14829,N_14748);
or UO_68 (O_68,N_14780,N_14408);
and UO_69 (O_69,N_14291,N_14894);
or UO_70 (O_70,N_14144,N_14044);
or UO_71 (O_71,N_14033,N_14062);
nand UO_72 (O_72,N_14441,N_14303);
or UO_73 (O_73,N_14875,N_14005);
and UO_74 (O_74,N_14733,N_14161);
nor UO_75 (O_75,N_14395,N_14380);
or UO_76 (O_76,N_14997,N_14614);
nand UO_77 (O_77,N_14147,N_14924);
or UO_78 (O_78,N_14474,N_14273);
nor UO_79 (O_79,N_14673,N_14772);
xnor UO_80 (O_80,N_14409,N_14775);
nand UO_81 (O_81,N_14606,N_14630);
xnor UO_82 (O_82,N_14731,N_14072);
or UO_83 (O_83,N_14531,N_14215);
nor UO_84 (O_84,N_14172,N_14830);
xnor UO_85 (O_85,N_14915,N_14939);
or UO_86 (O_86,N_14640,N_14238);
or UO_87 (O_87,N_14167,N_14508);
nor UO_88 (O_88,N_14065,N_14137);
and UO_89 (O_89,N_14266,N_14469);
nand UO_90 (O_90,N_14631,N_14836);
xnor UO_91 (O_91,N_14690,N_14320);
or UO_92 (O_92,N_14732,N_14891);
and UO_93 (O_93,N_14032,N_14381);
and UO_94 (O_94,N_14113,N_14200);
and UO_95 (O_95,N_14414,N_14211);
and UO_96 (O_96,N_14813,N_14175);
or UO_97 (O_97,N_14318,N_14217);
and UO_98 (O_98,N_14686,N_14424);
and UO_99 (O_99,N_14903,N_14854);
or UO_100 (O_100,N_14633,N_14007);
nand UO_101 (O_101,N_14623,N_14184);
nor UO_102 (O_102,N_14791,N_14899);
xor UO_103 (O_103,N_14735,N_14837);
nor UO_104 (O_104,N_14890,N_14437);
nor UO_105 (O_105,N_14391,N_14704);
nor UO_106 (O_106,N_14637,N_14263);
and UO_107 (O_107,N_14081,N_14527);
or UO_108 (O_108,N_14886,N_14573);
nor UO_109 (O_109,N_14265,N_14934);
and UO_110 (O_110,N_14553,N_14790);
xor UO_111 (O_111,N_14458,N_14236);
and UO_112 (O_112,N_14957,N_14832);
xor UO_113 (O_113,N_14868,N_14080);
or UO_114 (O_114,N_14475,N_14093);
and UO_115 (O_115,N_14193,N_14087);
nor UO_116 (O_116,N_14691,N_14094);
nand UO_117 (O_117,N_14587,N_14097);
nand UO_118 (O_118,N_14838,N_14786);
nor UO_119 (O_119,N_14426,N_14084);
and UO_120 (O_120,N_14150,N_14151);
nor UO_121 (O_121,N_14245,N_14756);
nand UO_122 (O_122,N_14595,N_14235);
nor UO_123 (O_123,N_14003,N_14542);
nor UO_124 (O_124,N_14059,N_14621);
nand UO_125 (O_125,N_14781,N_14734);
nand UO_126 (O_126,N_14898,N_14251);
nor UO_127 (O_127,N_14578,N_14361);
nand UO_128 (O_128,N_14242,N_14255);
nand UO_129 (O_129,N_14586,N_14947);
or UO_130 (O_130,N_14104,N_14367);
xnor UO_131 (O_131,N_14466,N_14078);
nand UO_132 (O_132,N_14122,N_14943);
and UO_133 (O_133,N_14759,N_14917);
nand UO_134 (O_134,N_14479,N_14889);
or UO_135 (O_135,N_14374,N_14712);
nor UO_136 (O_136,N_14356,N_14326);
xnor UO_137 (O_137,N_14074,N_14418);
nand UO_138 (O_138,N_14788,N_14463);
nor UO_139 (O_139,N_14779,N_14461);
nand UO_140 (O_140,N_14138,N_14909);
nand UO_141 (O_141,N_14224,N_14216);
or UO_142 (O_142,N_14363,N_14403);
xor UO_143 (O_143,N_14261,N_14905);
and UO_144 (O_144,N_14577,N_14278);
xor UO_145 (O_145,N_14117,N_14054);
nor UO_146 (O_146,N_14528,N_14831);
and UO_147 (O_147,N_14599,N_14135);
xnor UO_148 (O_148,N_14402,N_14991);
and UO_149 (O_149,N_14858,N_14176);
nand UO_150 (O_150,N_14302,N_14720);
nand UO_151 (O_151,N_14664,N_14638);
nand UO_152 (O_152,N_14692,N_14809);
or UO_153 (O_153,N_14038,N_14551);
nand UO_154 (O_154,N_14794,N_14256);
and UO_155 (O_155,N_14512,N_14041);
or UO_156 (O_156,N_14383,N_14058);
and UO_157 (O_157,N_14020,N_14445);
or UO_158 (O_158,N_14796,N_14243);
and UO_159 (O_159,N_14162,N_14680);
or UO_160 (O_160,N_14257,N_14422);
nor UO_161 (O_161,N_14787,N_14483);
or UO_162 (O_162,N_14321,N_14636);
or UO_163 (O_163,N_14331,N_14310);
nor UO_164 (O_164,N_14852,N_14675);
and UO_165 (O_165,N_14747,N_14572);
nor UO_166 (O_166,N_14160,N_14995);
nor UO_167 (O_167,N_14514,N_14872);
and UO_168 (O_168,N_14270,N_14406);
and UO_169 (O_169,N_14632,N_14694);
or UO_170 (O_170,N_14827,N_14362);
nor UO_171 (O_171,N_14598,N_14844);
nor UO_172 (O_172,N_14299,N_14448);
and UO_173 (O_173,N_14945,N_14800);
and UO_174 (O_174,N_14388,N_14272);
and UO_175 (O_175,N_14120,N_14396);
or UO_176 (O_176,N_14254,N_14481);
or UO_177 (O_177,N_14857,N_14769);
nor UO_178 (O_178,N_14695,N_14994);
nor UO_179 (O_179,N_14377,N_14333);
or UO_180 (O_180,N_14973,N_14765);
or UO_181 (O_181,N_14152,N_14999);
and UO_182 (O_182,N_14768,N_14760);
xnor UO_183 (O_183,N_14296,N_14451);
or UO_184 (O_184,N_14742,N_14503);
nor UO_185 (O_185,N_14169,N_14594);
nor UO_186 (O_186,N_14824,N_14157);
and UO_187 (O_187,N_14287,N_14334);
or UO_188 (O_188,N_14676,N_14060);
and UO_189 (O_189,N_14738,N_14223);
and UO_190 (O_190,N_14620,N_14795);
xor UO_191 (O_191,N_14806,N_14295);
or UO_192 (O_192,N_14027,N_14218);
nand UO_193 (O_193,N_14725,N_14646);
nor UO_194 (O_194,N_14534,N_14644);
or UO_195 (O_195,N_14412,N_14908);
nor UO_196 (O_196,N_14473,N_14118);
or UO_197 (O_197,N_14051,N_14439);
nor UO_198 (O_198,N_14037,N_14496);
or UO_199 (O_199,N_14359,N_14823);
and UO_200 (O_200,N_14154,N_14944);
nor UO_201 (O_201,N_14721,N_14754);
or UO_202 (O_202,N_14378,N_14842);
or UO_203 (O_203,N_14177,N_14355);
nand UO_204 (O_204,N_14373,N_14139);
and UO_205 (O_205,N_14179,N_14232);
or UO_206 (O_206,N_14289,N_14726);
or UO_207 (O_207,N_14576,N_14202);
or UO_208 (O_208,N_14521,N_14456);
and UO_209 (O_209,N_14658,N_14816);
or UO_210 (O_210,N_14629,N_14979);
nand UO_211 (O_211,N_14880,N_14014);
nor UO_212 (O_212,N_14106,N_14284);
xor UO_213 (O_213,N_14182,N_14543);
xnor UO_214 (O_214,N_14350,N_14906);
xor UO_215 (O_215,N_14047,N_14329);
nand UO_216 (O_216,N_14866,N_14476);
and UO_217 (O_217,N_14817,N_14582);
nand UO_218 (O_218,N_14090,N_14369);
xnor UO_219 (O_219,N_14657,N_14693);
nand UO_220 (O_220,N_14622,N_14046);
xnor UO_221 (O_221,N_14125,N_14384);
nand UO_222 (O_222,N_14468,N_14848);
and UO_223 (O_223,N_14647,N_14541);
xnor UO_224 (O_224,N_14913,N_14011);
nor UO_225 (O_225,N_14761,N_14275);
nor UO_226 (O_226,N_14677,N_14401);
nand UO_227 (O_227,N_14394,N_14068);
xnor UO_228 (O_228,N_14864,N_14605);
and UO_229 (O_229,N_14233,N_14064);
and UO_230 (O_230,N_14981,N_14313);
xnor UO_231 (O_231,N_14642,N_14882);
and UO_232 (O_232,N_14100,N_14849);
nand UO_233 (O_233,N_14870,N_14983);
or UO_234 (O_234,N_14716,N_14687);
or UO_235 (O_235,N_14440,N_14510);
nand UO_236 (O_236,N_14244,N_14221);
and UO_237 (O_237,N_14290,N_14904);
nor UO_238 (O_238,N_14271,N_14379);
and UO_239 (O_239,N_14322,N_14833);
nand UO_240 (O_240,N_14815,N_14400);
and UO_241 (O_241,N_14937,N_14070);
nor UO_242 (O_242,N_14478,N_14938);
and UO_243 (O_243,N_14338,N_14764);
xnor UO_244 (O_244,N_14034,N_14785);
or UO_245 (O_245,N_14336,N_14102);
or UO_246 (O_246,N_14085,N_14967);
and UO_247 (O_247,N_14259,N_14111);
or UO_248 (O_248,N_14031,N_14910);
nor UO_249 (O_249,N_14569,N_14746);
nand UO_250 (O_250,N_14523,N_14134);
nor UO_251 (O_251,N_14323,N_14782);
nor UO_252 (O_252,N_14546,N_14715);
and UO_253 (O_253,N_14180,N_14762);
nor UO_254 (O_254,N_14316,N_14285);
and UO_255 (O_255,N_14115,N_14453);
nor UO_256 (O_256,N_14392,N_14855);
nor UO_257 (O_257,N_14506,N_14375);
nor UO_258 (O_258,N_14513,N_14304);
nand UO_259 (O_259,N_14490,N_14752);
and UO_260 (O_260,N_14048,N_14489);
and UO_261 (O_261,N_14750,N_14867);
xnor UO_262 (O_262,N_14718,N_14229);
nand UO_263 (O_263,N_14568,N_14434);
or UO_264 (O_264,N_14472,N_14108);
nand UO_265 (O_265,N_14883,N_14425);
or UO_266 (O_266,N_14500,N_14696);
nand UO_267 (O_267,N_14042,N_14818);
nor UO_268 (O_268,N_14828,N_14420);
and UO_269 (O_269,N_14279,N_14464);
xnor UO_270 (O_270,N_14194,N_14069);
nor UO_271 (O_271,N_14444,N_14351);
xnor UO_272 (O_272,N_14486,N_14459);
nor UO_273 (O_273,N_14926,N_14557);
nand UO_274 (O_274,N_14793,N_14089);
nand UO_275 (O_275,N_14530,N_14484);
nand UO_276 (O_276,N_14063,N_14258);
or UO_277 (O_277,N_14969,N_14006);
or UO_278 (O_278,N_14148,N_14843);
nand UO_279 (O_279,N_14502,N_14537);
nor UO_280 (O_280,N_14571,N_14992);
nor UO_281 (O_281,N_14975,N_14429);
and UO_282 (O_282,N_14421,N_14191);
nor UO_283 (O_283,N_14965,N_14840);
nand UO_284 (O_284,N_14990,N_14753);
and UO_285 (O_285,N_14156,N_14228);
nand UO_286 (O_286,N_14371,N_14146);
and UO_287 (O_287,N_14755,N_14550);
or UO_288 (O_288,N_14928,N_14812);
nand UO_289 (O_289,N_14423,N_14185);
and UO_290 (O_290,N_14405,N_14600);
or UO_291 (O_291,N_14153,N_14635);
or UO_292 (O_292,N_14589,N_14022);
or UO_293 (O_293,N_14911,N_14652);
and UO_294 (O_294,N_14563,N_14988);
nor UO_295 (O_295,N_14149,N_14730);
or UO_296 (O_296,N_14346,N_14210);
and UO_297 (O_297,N_14091,N_14225);
or UO_298 (O_298,N_14711,N_14802);
and UO_299 (O_299,N_14192,N_14501);
nor UO_300 (O_300,N_14109,N_14532);
nand UO_301 (O_301,N_14612,N_14035);
xnor UO_302 (O_302,N_14015,N_14722);
nand UO_303 (O_303,N_14613,N_14368);
nand UO_304 (O_304,N_14230,N_14624);
nor UO_305 (O_305,N_14499,N_14964);
and UO_306 (O_306,N_14136,N_14049);
and UO_307 (O_307,N_14166,N_14925);
nand UO_308 (O_308,N_14312,N_14145);
nor UO_309 (O_309,N_14198,N_14547);
and UO_310 (O_310,N_14099,N_14204);
and UO_311 (O_311,N_14454,N_14250);
or UO_312 (O_312,N_14603,N_14159);
nand UO_313 (O_313,N_14404,N_14666);
nor UO_314 (O_314,N_14107,N_14447);
nor UO_315 (O_315,N_14307,N_14430);
and UO_316 (O_316,N_14061,N_14205);
and UO_317 (O_317,N_14165,N_14057);
or UO_318 (O_318,N_14873,N_14626);
and UO_319 (O_319,N_14053,N_14714);
xnor UO_320 (O_320,N_14438,N_14522);
and UO_321 (O_321,N_14209,N_14701);
or UO_322 (O_322,N_14655,N_14723);
nand UO_323 (O_323,N_14052,N_14993);
or UO_324 (O_324,N_14729,N_14862);
and UO_325 (O_325,N_14865,N_14366);
nor UO_326 (O_326,N_14277,N_14498);
nor UO_327 (O_327,N_14949,N_14110);
nor UO_328 (O_328,N_14298,N_14222);
and UO_329 (O_329,N_14850,N_14515);
nand UO_330 (O_330,N_14608,N_14931);
nand UO_331 (O_331,N_14398,N_14241);
nor UO_332 (O_332,N_14416,N_14884);
nor UO_333 (O_333,N_14708,N_14126);
nor UO_334 (O_334,N_14385,N_14778);
xor UO_335 (O_335,N_14494,N_14524);
nand UO_336 (O_336,N_14895,N_14114);
and UO_337 (O_337,N_14203,N_14040);
nand UO_338 (O_338,N_14504,N_14206);
nand UO_339 (O_339,N_14219,N_14082);
and UO_340 (O_340,N_14662,N_14803);
or UO_341 (O_341,N_14897,N_14674);
nand UO_342 (O_342,N_14497,N_14163);
nor UO_343 (O_343,N_14432,N_14766);
or UO_344 (O_344,N_14306,N_14846);
or UO_345 (O_345,N_14083,N_14583);
nand UO_346 (O_346,N_14538,N_14705);
nand UO_347 (O_347,N_14663,N_14018);
and UO_348 (O_348,N_14703,N_14590);
and UO_349 (O_349,N_14342,N_14561);
nand UO_350 (O_350,N_14592,N_14656);
nand UO_351 (O_351,N_14121,N_14942);
nand UO_352 (O_352,N_14056,N_14907);
nor UO_353 (O_353,N_14460,N_14863);
nor UO_354 (O_354,N_14281,N_14328);
nor UO_355 (O_355,N_14387,N_14930);
or UO_356 (O_356,N_14227,N_14317);
nor UO_357 (O_357,N_14349,N_14740);
or UO_358 (O_358,N_14881,N_14360);
nor UO_359 (O_359,N_14024,N_14955);
or UO_360 (O_360,N_14260,N_14076);
and UO_361 (O_361,N_14617,N_14845);
xor UO_362 (O_362,N_14319,N_14340);
and UO_363 (O_363,N_14170,N_14155);
or UO_364 (O_364,N_14183,N_14452);
nand UO_365 (O_365,N_14433,N_14536);
and UO_366 (O_366,N_14719,N_14376);
nor UO_367 (O_367,N_14682,N_14039);
and UO_368 (O_368,N_14477,N_14700);
and UO_369 (O_369,N_14158,N_14294);
xnor UO_370 (O_370,N_14826,N_14023);
or UO_371 (O_371,N_14188,N_14935);
xnor UO_372 (O_372,N_14982,N_14086);
nor UO_373 (O_373,N_14609,N_14593);
or UO_374 (O_374,N_14208,N_14397);
or UO_375 (O_375,N_14597,N_14878);
xnor UO_376 (O_376,N_14142,N_14834);
or UO_377 (O_377,N_14088,N_14098);
or UO_378 (O_378,N_14019,N_14615);
nand UO_379 (O_379,N_14171,N_14902);
nand UO_380 (O_380,N_14921,N_14564);
nand UO_381 (O_381,N_14526,N_14252);
nor UO_382 (O_382,N_14071,N_14961);
nor UO_383 (O_383,N_14067,N_14509);
and UO_384 (O_384,N_14262,N_14987);
and UO_385 (O_385,N_14885,N_14249);
and UO_386 (O_386,N_14297,N_14618);
or UO_387 (O_387,N_14744,N_14004);
or UO_388 (O_388,N_14231,N_14341);
or UO_389 (O_389,N_14467,N_14105);
or UO_390 (O_390,N_14628,N_14575);
or UO_391 (O_391,N_14237,N_14996);
xnor UO_392 (O_392,N_14968,N_14066);
nand UO_393 (O_393,N_14807,N_14859);
nand UO_394 (O_394,N_14610,N_14799);
nand UO_395 (O_395,N_14470,N_14588);
and UO_396 (O_396,N_14960,N_14140);
nand UO_397 (O_397,N_14267,N_14737);
xor UO_398 (O_398,N_14976,N_14308);
xnor UO_399 (O_399,N_14689,N_14627);
nand UO_400 (O_400,N_14443,N_14050);
or UO_401 (O_401,N_14293,N_14309);
nor UO_402 (O_402,N_14199,N_14948);
nand UO_403 (O_403,N_14648,N_14953);
nor UO_404 (O_404,N_14869,N_14554);
nand UO_405 (O_405,N_14954,N_14482);
xor UO_406 (O_406,N_14776,N_14574);
nand UO_407 (O_407,N_14212,N_14325);
or UO_408 (O_408,N_14491,N_14562);
or UO_409 (O_409,N_14672,N_14717);
nand UO_410 (O_410,N_14239,N_14410);
nor UO_411 (O_411,N_14684,N_14311);
nor UO_412 (O_412,N_14305,N_14213);
and UO_413 (O_413,N_14511,N_14856);
and UO_414 (O_414,N_14679,N_14029);
nor UO_415 (O_415,N_14181,N_14001);
nor UO_416 (O_416,N_14516,N_14095);
or UO_417 (O_417,N_14616,N_14419);
nand UO_418 (O_418,N_14315,N_14335);
xor UO_419 (O_419,N_14214,N_14566);
nor UO_420 (O_420,N_14036,N_14343);
nor UO_421 (O_421,N_14596,N_14455);
nand UO_422 (O_422,N_14449,N_14822);
nand UO_423 (O_423,N_14301,N_14941);
or UO_424 (O_424,N_14190,N_14517);
nor UO_425 (O_425,N_14390,N_14480);
and UO_426 (O_426,N_14654,N_14079);
or UO_427 (O_427,N_14407,N_14446);
or UO_428 (O_428,N_14601,N_14286);
or UO_429 (O_429,N_14442,N_14382);
and UO_430 (O_430,N_14021,N_14579);
or UO_431 (O_431,N_14751,N_14248);
or UO_432 (O_432,N_14736,N_14505);
nor UO_433 (O_433,N_14825,N_14493);
nor UO_434 (O_434,N_14820,N_14853);
or UO_435 (O_435,N_14457,N_14415);
and UO_436 (O_436,N_14946,N_14972);
nand UO_437 (O_437,N_14116,N_14977);
xnor UO_438 (O_438,N_14989,N_14348);
xor UO_439 (O_439,N_14611,N_14345);
or UO_440 (O_440,N_14013,N_14539);
and UO_441 (O_441,N_14952,N_14518);
nor UO_442 (O_442,N_14739,N_14936);
or UO_443 (O_443,N_14665,N_14835);
and UO_444 (O_444,N_14300,N_14196);
nor UO_445 (O_445,N_14413,N_14043);
or UO_446 (O_446,N_14970,N_14073);
and UO_447 (O_447,N_14770,N_14651);
nand UO_448 (O_448,N_14808,N_14280);
nand UO_449 (O_449,N_14959,N_14119);
xnor UO_450 (O_450,N_14727,N_14798);
xnor UO_451 (O_451,N_14540,N_14565);
nand UO_452 (O_452,N_14580,N_14879);
nor UO_453 (O_453,N_14709,N_14370);
or UO_454 (O_454,N_14893,N_14901);
or UO_455 (O_455,N_14028,N_14940);
nor UO_456 (O_456,N_14892,N_14186);
nor UO_457 (O_457,N_14164,N_14792);
nor UO_458 (O_458,N_14607,N_14399);
or UO_459 (O_459,N_14929,N_14324);
nand UO_460 (O_460,N_14462,N_14174);
nand UO_461 (O_461,N_14874,N_14347);
and UO_462 (O_462,N_14963,N_14841);
or UO_463 (O_463,N_14784,N_14389);
and UO_464 (O_464,N_14888,N_14000);
nand UO_465 (O_465,N_14075,N_14767);
xor UO_466 (O_466,N_14197,N_14871);
nand UO_467 (O_467,N_14797,N_14743);
xor UO_468 (O_468,N_14092,N_14604);
nor UO_469 (O_469,N_14127,N_14096);
nand UO_470 (O_470,N_14465,N_14103);
or UO_471 (O_471,N_14558,N_14220);
nand UO_472 (O_472,N_14985,N_14372);
nand UO_473 (O_473,N_14327,N_14525);
nor UO_474 (O_474,N_14008,N_14128);
or UO_475 (O_475,N_14688,N_14773);
nand UO_476 (O_476,N_14702,N_14045);
and UO_477 (O_477,N_14661,N_14966);
and UO_478 (O_478,N_14549,N_14919);
nand UO_479 (O_479,N_14026,N_14706);
or UO_480 (O_480,N_14201,N_14923);
nor UO_481 (O_481,N_14274,N_14699);
nor UO_482 (O_482,N_14649,N_14431);
or UO_483 (O_483,N_14810,N_14269);
and UO_484 (O_484,N_14101,N_14012);
and UO_485 (O_485,N_14697,N_14495);
nor UO_486 (O_486,N_14567,N_14112);
nand UO_487 (O_487,N_14821,N_14650);
and UO_488 (O_488,N_14002,N_14552);
nand UO_489 (O_489,N_14774,N_14876);
nand UO_490 (O_490,N_14010,N_14544);
nor UO_491 (O_491,N_14436,N_14962);
nand UO_492 (O_492,N_14920,N_14927);
and UO_493 (O_493,N_14435,N_14643);
nor UO_494 (O_494,N_14683,N_14358);
or UO_495 (O_495,N_14268,N_14283);
nand UO_496 (O_496,N_14998,N_14771);
and UO_497 (O_497,N_14978,N_14025);
nand UO_498 (O_498,N_14123,N_14896);
nand UO_499 (O_499,N_14741,N_14471);
nand UO_500 (O_500,N_14342,N_14601);
and UO_501 (O_501,N_14772,N_14730);
nor UO_502 (O_502,N_14031,N_14129);
nor UO_503 (O_503,N_14000,N_14209);
xor UO_504 (O_504,N_14712,N_14737);
nand UO_505 (O_505,N_14593,N_14168);
or UO_506 (O_506,N_14003,N_14035);
nor UO_507 (O_507,N_14131,N_14393);
or UO_508 (O_508,N_14306,N_14188);
nand UO_509 (O_509,N_14459,N_14815);
xor UO_510 (O_510,N_14378,N_14257);
nand UO_511 (O_511,N_14995,N_14848);
nand UO_512 (O_512,N_14357,N_14790);
xor UO_513 (O_513,N_14767,N_14036);
and UO_514 (O_514,N_14869,N_14099);
and UO_515 (O_515,N_14723,N_14344);
and UO_516 (O_516,N_14454,N_14730);
nand UO_517 (O_517,N_14855,N_14784);
and UO_518 (O_518,N_14862,N_14563);
nand UO_519 (O_519,N_14430,N_14783);
and UO_520 (O_520,N_14444,N_14087);
or UO_521 (O_521,N_14240,N_14791);
xor UO_522 (O_522,N_14403,N_14450);
xor UO_523 (O_523,N_14613,N_14697);
or UO_524 (O_524,N_14981,N_14704);
nand UO_525 (O_525,N_14546,N_14119);
or UO_526 (O_526,N_14158,N_14624);
nor UO_527 (O_527,N_14872,N_14652);
or UO_528 (O_528,N_14474,N_14592);
or UO_529 (O_529,N_14550,N_14967);
or UO_530 (O_530,N_14290,N_14669);
nor UO_531 (O_531,N_14643,N_14029);
nand UO_532 (O_532,N_14026,N_14927);
or UO_533 (O_533,N_14659,N_14537);
and UO_534 (O_534,N_14102,N_14189);
nand UO_535 (O_535,N_14580,N_14669);
nor UO_536 (O_536,N_14148,N_14545);
and UO_537 (O_537,N_14807,N_14040);
or UO_538 (O_538,N_14335,N_14509);
nand UO_539 (O_539,N_14273,N_14521);
and UO_540 (O_540,N_14736,N_14157);
or UO_541 (O_541,N_14301,N_14850);
nor UO_542 (O_542,N_14751,N_14446);
or UO_543 (O_543,N_14980,N_14883);
and UO_544 (O_544,N_14933,N_14215);
and UO_545 (O_545,N_14021,N_14341);
or UO_546 (O_546,N_14487,N_14407);
or UO_547 (O_547,N_14661,N_14852);
or UO_548 (O_548,N_14244,N_14880);
or UO_549 (O_549,N_14967,N_14072);
or UO_550 (O_550,N_14625,N_14076);
or UO_551 (O_551,N_14797,N_14596);
or UO_552 (O_552,N_14932,N_14790);
and UO_553 (O_553,N_14391,N_14385);
and UO_554 (O_554,N_14370,N_14209);
nand UO_555 (O_555,N_14224,N_14005);
nor UO_556 (O_556,N_14904,N_14519);
and UO_557 (O_557,N_14851,N_14540);
nand UO_558 (O_558,N_14479,N_14846);
and UO_559 (O_559,N_14020,N_14967);
nor UO_560 (O_560,N_14996,N_14206);
and UO_561 (O_561,N_14754,N_14255);
or UO_562 (O_562,N_14946,N_14498);
nor UO_563 (O_563,N_14881,N_14174);
nand UO_564 (O_564,N_14287,N_14475);
and UO_565 (O_565,N_14983,N_14280);
and UO_566 (O_566,N_14176,N_14187);
nor UO_567 (O_567,N_14492,N_14871);
nand UO_568 (O_568,N_14772,N_14995);
nand UO_569 (O_569,N_14993,N_14912);
nand UO_570 (O_570,N_14187,N_14711);
and UO_571 (O_571,N_14522,N_14136);
nor UO_572 (O_572,N_14284,N_14611);
nand UO_573 (O_573,N_14133,N_14160);
xnor UO_574 (O_574,N_14044,N_14395);
nor UO_575 (O_575,N_14865,N_14981);
nor UO_576 (O_576,N_14761,N_14314);
nor UO_577 (O_577,N_14116,N_14786);
and UO_578 (O_578,N_14391,N_14988);
nand UO_579 (O_579,N_14906,N_14605);
nand UO_580 (O_580,N_14685,N_14395);
nand UO_581 (O_581,N_14899,N_14472);
nand UO_582 (O_582,N_14284,N_14390);
nor UO_583 (O_583,N_14614,N_14906);
and UO_584 (O_584,N_14269,N_14676);
nor UO_585 (O_585,N_14303,N_14898);
or UO_586 (O_586,N_14166,N_14738);
nand UO_587 (O_587,N_14146,N_14865);
and UO_588 (O_588,N_14925,N_14750);
and UO_589 (O_589,N_14738,N_14484);
nand UO_590 (O_590,N_14099,N_14828);
and UO_591 (O_591,N_14025,N_14220);
or UO_592 (O_592,N_14898,N_14006);
or UO_593 (O_593,N_14211,N_14714);
nor UO_594 (O_594,N_14594,N_14022);
nor UO_595 (O_595,N_14465,N_14484);
nor UO_596 (O_596,N_14739,N_14900);
or UO_597 (O_597,N_14212,N_14294);
nor UO_598 (O_598,N_14978,N_14438);
nand UO_599 (O_599,N_14188,N_14681);
or UO_600 (O_600,N_14782,N_14860);
nand UO_601 (O_601,N_14446,N_14007);
or UO_602 (O_602,N_14667,N_14862);
nand UO_603 (O_603,N_14131,N_14035);
and UO_604 (O_604,N_14484,N_14054);
nand UO_605 (O_605,N_14167,N_14216);
nand UO_606 (O_606,N_14293,N_14108);
or UO_607 (O_607,N_14989,N_14882);
xor UO_608 (O_608,N_14722,N_14423);
and UO_609 (O_609,N_14798,N_14556);
and UO_610 (O_610,N_14087,N_14387);
and UO_611 (O_611,N_14948,N_14965);
nor UO_612 (O_612,N_14761,N_14558);
and UO_613 (O_613,N_14136,N_14072);
xnor UO_614 (O_614,N_14128,N_14817);
xnor UO_615 (O_615,N_14085,N_14264);
or UO_616 (O_616,N_14935,N_14468);
or UO_617 (O_617,N_14288,N_14330);
nand UO_618 (O_618,N_14094,N_14767);
and UO_619 (O_619,N_14181,N_14918);
nor UO_620 (O_620,N_14815,N_14374);
nor UO_621 (O_621,N_14907,N_14645);
xor UO_622 (O_622,N_14626,N_14989);
or UO_623 (O_623,N_14302,N_14050);
and UO_624 (O_624,N_14770,N_14753);
nor UO_625 (O_625,N_14399,N_14382);
nand UO_626 (O_626,N_14010,N_14333);
nand UO_627 (O_627,N_14950,N_14900);
or UO_628 (O_628,N_14600,N_14651);
nand UO_629 (O_629,N_14615,N_14897);
and UO_630 (O_630,N_14753,N_14464);
nand UO_631 (O_631,N_14018,N_14747);
nor UO_632 (O_632,N_14816,N_14265);
xor UO_633 (O_633,N_14756,N_14752);
nor UO_634 (O_634,N_14741,N_14182);
xor UO_635 (O_635,N_14691,N_14529);
nor UO_636 (O_636,N_14199,N_14723);
xnor UO_637 (O_637,N_14036,N_14698);
xor UO_638 (O_638,N_14281,N_14716);
and UO_639 (O_639,N_14253,N_14872);
or UO_640 (O_640,N_14109,N_14187);
xor UO_641 (O_641,N_14641,N_14352);
xnor UO_642 (O_642,N_14452,N_14882);
nor UO_643 (O_643,N_14627,N_14649);
and UO_644 (O_644,N_14605,N_14759);
nand UO_645 (O_645,N_14528,N_14909);
nand UO_646 (O_646,N_14390,N_14319);
and UO_647 (O_647,N_14296,N_14125);
or UO_648 (O_648,N_14497,N_14648);
nand UO_649 (O_649,N_14965,N_14499);
nor UO_650 (O_650,N_14792,N_14486);
nand UO_651 (O_651,N_14318,N_14471);
nand UO_652 (O_652,N_14259,N_14803);
and UO_653 (O_653,N_14308,N_14834);
or UO_654 (O_654,N_14692,N_14277);
and UO_655 (O_655,N_14203,N_14490);
and UO_656 (O_656,N_14888,N_14460);
and UO_657 (O_657,N_14899,N_14029);
and UO_658 (O_658,N_14652,N_14510);
or UO_659 (O_659,N_14542,N_14495);
xor UO_660 (O_660,N_14604,N_14817);
nand UO_661 (O_661,N_14241,N_14931);
nor UO_662 (O_662,N_14961,N_14770);
or UO_663 (O_663,N_14743,N_14116);
nor UO_664 (O_664,N_14128,N_14656);
nand UO_665 (O_665,N_14942,N_14547);
nand UO_666 (O_666,N_14913,N_14488);
and UO_667 (O_667,N_14037,N_14246);
nor UO_668 (O_668,N_14079,N_14794);
nor UO_669 (O_669,N_14245,N_14917);
nand UO_670 (O_670,N_14539,N_14631);
or UO_671 (O_671,N_14458,N_14154);
nor UO_672 (O_672,N_14937,N_14981);
nand UO_673 (O_673,N_14420,N_14084);
nand UO_674 (O_674,N_14478,N_14673);
or UO_675 (O_675,N_14157,N_14714);
nor UO_676 (O_676,N_14044,N_14541);
or UO_677 (O_677,N_14468,N_14358);
nand UO_678 (O_678,N_14471,N_14837);
nand UO_679 (O_679,N_14826,N_14069);
and UO_680 (O_680,N_14003,N_14264);
nand UO_681 (O_681,N_14937,N_14306);
nor UO_682 (O_682,N_14126,N_14650);
xnor UO_683 (O_683,N_14317,N_14381);
and UO_684 (O_684,N_14713,N_14716);
or UO_685 (O_685,N_14401,N_14823);
nand UO_686 (O_686,N_14973,N_14169);
or UO_687 (O_687,N_14438,N_14780);
and UO_688 (O_688,N_14773,N_14463);
xnor UO_689 (O_689,N_14234,N_14746);
nand UO_690 (O_690,N_14336,N_14282);
and UO_691 (O_691,N_14781,N_14965);
or UO_692 (O_692,N_14240,N_14365);
nand UO_693 (O_693,N_14041,N_14105);
and UO_694 (O_694,N_14134,N_14124);
nor UO_695 (O_695,N_14291,N_14962);
nand UO_696 (O_696,N_14664,N_14209);
nor UO_697 (O_697,N_14406,N_14888);
and UO_698 (O_698,N_14299,N_14467);
nand UO_699 (O_699,N_14447,N_14467);
or UO_700 (O_700,N_14938,N_14041);
and UO_701 (O_701,N_14513,N_14985);
nor UO_702 (O_702,N_14821,N_14878);
xnor UO_703 (O_703,N_14838,N_14394);
or UO_704 (O_704,N_14953,N_14024);
or UO_705 (O_705,N_14445,N_14920);
and UO_706 (O_706,N_14433,N_14572);
nand UO_707 (O_707,N_14959,N_14982);
nand UO_708 (O_708,N_14073,N_14888);
or UO_709 (O_709,N_14620,N_14609);
nand UO_710 (O_710,N_14131,N_14354);
and UO_711 (O_711,N_14037,N_14240);
nor UO_712 (O_712,N_14059,N_14002);
and UO_713 (O_713,N_14225,N_14849);
nor UO_714 (O_714,N_14398,N_14954);
nor UO_715 (O_715,N_14588,N_14463);
nor UO_716 (O_716,N_14649,N_14112);
nand UO_717 (O_717,N_14418,N_14035);
nor UO_718 (O_718,N_14152,N_14363);
and UO_719 (O_719,N_14526,N_14678);
and UO_720 (O_720,N_14812,N_14967);
nor UO_721 (O_721,N_14284,N_14670);
nor UO_722 (O_722,N_14848,N_14173);
or UO_723 (O_723,N_14541,N_14899);
and UO_724 (O_724,N_14848,N_14884);
nor UO_725 (O_725,N_14398,N_14691);
nand UO_726 (O_726,N_14282,N_14806);
or UO_727 (O_727,N_14502,N_14993);
xor UO_728 (O_728,N_14931,N_14083);
nand UO_729 (O_729,N_14650,N_14686);
or UO_730 (O_730,N_14246,N_14300);
or UO_731 (O_731,N_14907,N_14255);
nor UO_732 (O_732,N_14434,N_14387);
and UO_733 (O_733,N_14287,N_14579);
or UO_734 (O_734,N_14794,N_14816);
or UO_735 (O_735,N_14475,N_14225);
or UO_736 (O_736,N_14888,N_14074);
or UO_737 (O_737,N_14766,N_14433);
xor UO_738 (O_738,N_14620,N_14069);
nand UO_739 (O_739,N_14366,N_14009);
nand UO_740 (O_740,N_14528,N_14873);
and UO_741 (O_741,N_14560,N_14636);
and UO_742 (O_742,N_14881,N_14030);
nand UO_743 (O_743,N_14808,N_14725);
nand UO_744 (O_744,N_14087,N_14943);
and UO_745 (O_745,N_14013,N_14375);
nand UO_746 (O_746,N_14851,N_14866);
nand UO_747 (O_747,N_14748,N_14011);
and UO_748 (O_748,N_14768,N_14829);
or UO_749 (O_749,N_14503,N_14463);
nor UO_750 (O_750,N_14813,N_14759);
and UO_751 (O_751,N_14486,N_14313);
xnor UO_752 (O_752,N_14070,N_14110);
or UO_753 (O_753,N_14209,N_14361);
or UO_754 (O_754,N_14717,N_14470);
or UO_755 (O_755,N_14713,N_14923);
and UO_756 (O_756,N_14469,N_14300);
or UO_757 (O_757,N_14293,N_14151);
and UO_758 (O_758,N_14786,N_14825);
or UO_759 (O_759,N_14909,N_14213);
and UO_760 (O_760,N_14759,N_14325);
xnor UO_761 (O_761,N_14769,N_14952);
nor UO_762 (O_762,N_14658,N_14700);
nand UO_763 (O_763,N_14708,N_14640);
nand UO_764 (O_764,N_14595,N_14800);
and UO_765 (O_765,N_14278,N_14024);
or UO_766 (O_766,N_14971,N_14622);
or UO_767 (O_767,N_14053,N_14405);
and UO_768 (O_768,N_14092,N_14383);
xnor UO_769 (O_769,N_14864,N_14635);
nand UO_770 (O_770,N_14527,N_14997);
or UO_771 (O_771,N_14758,N_14783);
nor UO_772 (O_772,N_14299,N_14688);
xor UO_773 (O_773,N_14666,N_14070);
and UO_774 (O_774,N_14779,N_14102);
nand UO_775 (O_775,N_14457,N_14011);
nand UO_776 (O_776,N_14960,N_14389);
nor UO_777 (O_777,N_14838,N_14843);
nand UO_778 (O_778,N_14325,N_14923);
and UO_779 (O_779,N_14396,N_14234);
and UO_780 (O_780,N_14016,N_14847);
and UO_781 (O_781,N_14306,N_14567);
or UO_782 (O_782,N_14754,N_14981);
and UO_783 (O_783,N_14074,N_14898);
nor UO_784 (O_784,N_14680,N_14721);
nor UO_785 (O_785,N_14957,N_14763);
and UO_786 (O_786,N_14172,N_14623);
nand UO_787 (O_787,N_14381,N_14377);
nand UO_788 (O_788,N_14571,N_14619);
or UO_789 (O_789,N_14438,N_14216);
nand UO_790 (O_790,N_14261,N_14994);
xor UO_791 (O_791,N_14283,N_14029);
xnor UO_792 (O_792,N_14143,N_14263);
nand UO_793 (O_793,N_14499,N_14807);
or UO_794 (O_794,N_14755,N_14800);
and UO_795 (O_795,N_14551,N_14887);
nor UO_796 (O_796,N_14464,N_14871);
nand UO_797 (O_797,N_14814,N_14880);
or UO_798 (O_798,N_14449,N_14969);
nand UO_799 (O_799,N_14395,N_14999);
and UO_800 (O_800,N_14383,N_14481);
nor UO_801 (O_801,N_14209,N_14995);
nand UO_802 (O_802,N_14393,N_14775);
and UO_803 (O_803,N_14266,N_14311);
nor UO_804 (O_804,N_14233,N_14361);
and UO_805 (O_805,N_14017,N_14857);
or UO_806 (O_806,N_14122,N_14324);
nand UO_807 (O_807,N_14644,N_14236);
and UO_808 (O_808,N_14030,N_14611);
nand UO_809 (O_809,N_14193,N_14399);
nor UO_810 (O_810,N_14308,N_14050);
and UO_811 (O_811,N_14014,N_14497);
and UO_812 (O_812,N_14227,N_14319);
nor UO_813 (O_813,N_14641,N_14840);
xor UO_814 (O_814,N_14740,N_14396);
and UO_815 (O_815,N_14971,N_14829);
or UO_816 (O_816,N_14713,N_14220);
nor UO_817 (O_817,N_14482,N_14122);
and UO_818 (O_818,N_14320,N_14998);
and UO_819 (O_819,N_14423,N_14601);
nand UO_820 (O_820,N_14301,N_14952);
or UO_821 (O_821,N_14583,N_14254);
nand UO_822 (O_822,N_14192,N_14051);
or UO_823 (O_823,N_14837,N_14604);
xnor UO_824 (O_824,N_14637,N_14445);
nand UO_825 (O_825,N_14853,N_14367);
nand UO_826 (O_826,N_14148,N_14897);
nor UO_827 (O_827,N_14264,N_14570);
or UO_828 (O_828,N_14017,N_14392);
xnor UO_829 (O_829,N_14466,N_14665);
and UO_830 (O_830,N_14798,N_14995);
or UO_831 (O_831,N_14948,N_14539);
nor UO_832 (O_832,N_14948,N_14546);
xor UO_833 (O_833,N_14115,N_14123);
and UO_834 (O_834,N_14545,N_14630);
or UO_835 (O_835,N_14586,N_14280);
xnor UO_836 (O_836,N_14547,N_14834);
nor UO_837 (O_837,N_14363,N_14255);
nor UO_838 (O_838,N_14082,N_14338);
xnor UO_839 (O_839,N_14189,N_14515);
nor UO_840 (O_840,N_14708,N_14401);
nor UO_841 (O_841,N_14832,N_14927);
or UO_842 (O_842,N_14485,N_14254);
nor UO_843 (O_843,N_14426,N_14392);
and UO_844 (O_844,N_14636,N_14007);
nor UO_845 (O_845,N_14973,N_14881);
nand UO_846 (O_846,N_14786,N_14824);
nand UO_847 (O_847,N_14534,N_14701);
xnor UO_848 (O_848,N_14749,N_14798);
and UO_849 (O_849,N_14936,N_14651);
and UO_850 (O_850,N_14268,N_14169);
or UO_851 (O_851,N_14226,N_14385);
or UO_852 (O_852,N_14061,N_14885);
xnor UO_853 (O_853,N_14554,N_14082);
or UO_854 (O_854,N_14053,N_14850);
and UO_855 (O_855,N_14066,N_14162);
and UO_856 (O_856,N_14197,N_14408);
nand UO_857 (O_857,N_14621,N_14732);
nand UO_858 (O_858,N_14750,N_14327);
or UO_859 (O_859,N_14704,N_14270);
xor UO_860 (O_860,N_14727,N_14773);
nand UO_861 (O_861,N_14099,N_14607);
and UO_862 (O_862,N_14332,N_14338);
nand UO_863 (O_863,N_14320,N_14434);
nand UO_864 (O_864,N_14553,N_14635);
nand UO_865 (O_865,N_14704,N_14920);
nor UO_866 (O_866,N_14173,N_14715);
xor UO_867 (O_867,N_14816,N_14684);
nor UO_868 (O_868,N_14769,N_14120);
nor UO_869 (O_869,N_14185,N_14833);
and UO_870 (O_870,N_14228,N_14056);
xnor UO_871 (O_871,N_14837,N_14715);
and UO_872 (O_872,N_14000,N_14245);
nand UO_873 (O_873,N_14518,N_14763);
and UO_874 (O_874,N_14544,N_14382);
and UO_875 (O_875,N_14875,N_14597);
or UO_876 (O_876,N_14552,N_14553);
and UO_877 (O_877,N_14215,N_14256);
and UO_878 (O_878,N_14165,N_14389);
nor UO_879 (O_879,N_14878,N_14705);
xor UO_880 (O_880,N_14164,N_14235);
and UO_881 (O_881,N_14449,N_14950);
and UO_882 (O_882,N_14782,N_14784);
and UO_883 (O_883,N_14649,N_14139);
or UO_884 (O_884,N_14628,N_14015);
or UO_885 (O_885,N_14223,N_14935);
xor UO_886 (O_886,N_14625,N_14332);
nand UO_887 (O_887,N_14166,N_14894);
nor UO_888 (O_888,N_14447,N_14181);
xnor UO_889 (O_889,N_14414,N_14127);
and UO_890 (O_890,N_14080,N_14951);
nand UO_891 (O_891,N_14223,N_14995);
nor UO_892 (O_892,N_14436,N_14563);
nand UO_893 (O_893,N_14513,N_14736);
nand UO_894 (O_894,N_14726,N_14921);
xor UO_895 (O_895,N_14975,N_14042);
and UO_896 (O_896,N_14573,N_14191);
nand UO_897 (O_897,N_14225,N_14447);
and UO_898 (O_898,N_14578,N_14262);
nor UO_899 (O_899,N_14804,N_14442);
xor UO_900 (O_900,N_14380,N_14929);
nand UO_901 (O_901,N_14001,N_14581);
nand UO_902 (O_902,N_14722,N_14833);
or UO_903 (O_903,N_14030,N_14776);
nand UO_904 (O_904,N_14878,N_14466);
nand UO_905 (O_905,N_14724,N_14112);
and UO_906 (O_906,N_14482,N_14618);
and UO_907 (O_907,N_14734,N_14010);
and UO_908 (O_908,N_14981,N_14799);
and UO_909 (O_909,N_14455,N_14298);
and UO_910 (O_910,N_14468,N_14477);
nand UO_911 (O_911,N_14429,N_14906);
and UO_912 (O_912,N_14039,N_14006);
or UO_913 (O_913,N_14814,N_14556);
or UO_914 (O_914,N_14968,N_14179);
and UO_915 (O_915,N_14019,N_14836);
xor UO_916 (O_916,N_14785,N_14120);
nand UO_917 (O_917,N_14711,N_14406);
nand UO_918 (O_918,N_14670,N_14105);
or UO_919 (O_919,N_14619,N_14588);
and UO_920 (O_920,N_14293,N_14503);
xnor UO_921 (O_921,N_14325,N_14589);
or UO_922 (O_922,N_14378,N_14785);
or UO_923 (O_923,N_14967,N_14399);
and UO_924 (O_924,N_14351,N_14449);
and UO_925 (O_925,N_14513,N_14446);
and UO_926 (O_926,N_14326,N_14684);
nor UO_927 (O_927,N_14510,N_14203);
nand UO_928 (O_928,N_14412,N_14133);
nand UO_929 (O_929,N_14292,N_14868);
nand UO_930 (O_930,N_14457,N_14849);
nor UO_931 (O_931,N_14690,N_14917);
or UO_932 (O_932,N_14678,N_14037);
xor UO_933 (O_933,N_14491,N_14237);
or UO_934 (O_934,N_14000,N_14297);
or UO_935 (O_935,N_14926,N_14793);
and UO_936 (O_936,N_14596,N_14393);
nand UO_937 (O_937,N_14731,N_14912);
and UO_938 (O_938,N_14143,N_14956);
or UO_939 (O_939,N_14211,N_14759);
nor UO_940 (O_940,N_14235,N_14715);
or UO_941 (O_941,N_14158,N_14104);
or UO_942 (O_942,N_14015,N_14143);
nor UO_943 (O_943,N_14490,N_14108);
nor UO_944 (O_944,N_14992,N_14578);
nor UO_945 (O_945,N_14126,N_14763);
nand UO_946 (O_946,N_14850,N_14636);
and UO_947 (O_947,N_14630,N_14572);
nor UO_948 (O_948,N_14578,N_14271);
nor UO_949 (O_949,N_14950,N_14841);
or UO_950 (O_950,N_14311,N_14924);
or UO_951 (O_951,N_14251,N_14333);
and UO_952 (O_952,N_14560,N_14462);
nand UO_953 (O_953,N_14744,N_14300);
nor UO_954 (O_954,N_14921,N_14845);
and UO_955 (O_955,N_14842,N_14032);
and UO_956 (O_956,N_14440,N_14198);
or UO_957 (O_957,N_14330,N_14077);
or UO_958 (O_958,N_14220,N_14928);
nand UO_959 (O_959,N_14867,N_14226);
nand UO_960 (O_960,N_14718,N_14832);
or UO_961 (O_961,N_14946,N_14854);
nand UO_962 (O_962,N_14207,N_14634);
and UO_963 (O_963,N_14666,N_14697);
nor UO_964 (O_964,N_14016,N_14046);
and UO_965 (O_965,N_14589,N_14557);
xor UO_966 (O_966,N_14682,N_14654);
or UO_967 (O_967,N_14446,N_14984);
or UO_968 (O_968,N_14039,N_14513);
xnor UO_969 (O_969,N_14628,N_14089);
or UO_970 (O_970,N_14730,N_14317);
nand UO_971 (O_971,N_14267,N_14103);
and UO_972 (O_972,N_14436,N_14537);
and UO_973 (O_973,N_14726,N_14291);
or UO_974 (O_974,N_14048,N_14259);
nor UO_975 (O_975,N_14675,N_14217);
and UO_976 (O_976,N_14644,N_14497);
nor UO_977 (O_977,N_14998,N_14650);
nand UO_978 (O_978,N_14571,N_14008);
nand UO_979 (O_979,N_14604,N_14071);
or UO_980 (O_980,N_14631,N_14464);
nand UO_981 (O_981,N_14580,N_14651);
and UO_982 (O_982,N_14884,N_14476);
nor UO_983 (O_983,N_14070,N_14744);
nand UO_984 (O_984,N_14717,N_14685);
nand UO_985 (O_985,N_14099,N_14583);
nand UO_986 (O_986,N_14787,N_14364);
or UO_987 (O_987,N_14232,N_14199);
nor UO_988 (O_988,N_14539,N_14649);
nor UO_989 (O_989,N_14747,N_14000);
or UO_990 (O_990,N_14031,N_14764);
and UO_991 (O_991,N_14007,N_14956);
xnor UO_992 (O_992,N_14633,N_14135);
or UO_993 (O_993,N_14607,N_14082);
nand UO_994 (O_994,N_14449,N_14763);
or UO_995 (O_995,N_14047,N_14972);
and UO_996 (O_996,N_14353,N_14888);
xor UO_997 (O_997,N_14738,N_14561);
nand UO_998 (O_998,N_14941,N_14383);
or UO_999 (O_999,N_14532,N_14296);
or UO_1000 (O_1000,N_14618,N_14528);
nand UO_1001 (O_1001,N_14084,N_14741);
and UO_1002 (O_1002,N_14012,N_14180);
nor UO_1003 (O_1003,N_14298,N_14631);
nand UO_1004 (O_1004,N_14737,N_14189);
nor UO_1005 (O_1005,N_14515,N_14981);
nand UO_1006 (O_1006,N_14506,N_14491);
or UO_1007 (O_1007,N_14443,N_14620);
nor UO_1008 (O_1008,N_14636,N_14783);
and UO_1009 (O_1009,N_14532,N_14649);
or UO_1010 (O_1010,N_14938,N_14219);
or UO_1011 (O_1011,N_14708,N_14632);
and UO_1012 (O_1012,N_14535,N_14417);
nand UO_1013 (O_1013,N_14215,N_14150);
and UO_1014 (O_1014,N_14814,N_14530);
nand UO_1015 (O_1015,N_14014,N_14965);
nor UO_1016 (O_1016,N_14234,N_14316);
and UO_1017 (O_1017,N_14489,N_14344);
nor UO_1018 (O_1018,N_14012,N_14578);
nor UO_1019 (O_1019,N_14929,N_14086);
nor UO_1020 (O_1020,N_14397,N_14562);
or UO_1021 (O_1021,N_14137,N_14857);
and UO_1022 (O_1022,N_14297,N_14885);
nor UO_1023 (O_1023,N_14066,N_14890);
nor UO_1024 (O_1024,N_14613,N_14597);
nor UO_1025 (O_1025,N_14464,N_14517);
nor UO_1026 (O_1026,N_14695,N_14429);
xor UO_1027 (O_1027,N_14788,N_14226);
or UO_1028 (O_1028,N_14919,N_14293);
nand UO_1029 (O_1029,N_14244,N_14250);
nand UO_1030 (O_1030,N_14025,N_14545);
nand UO_1031 (O_1031,N_14013,N_14426);
and UO_1032 (O_1032,N_14180,N_14797);
xnor UO_1033 (O_1033,N_14136,N_14859);
nor UO_1034 (O_1034,N_14852,N_14176);
nor UO_1035 (O_1035,N_14721,N_14698);
and UO_1036 (O_1036,N_14788,N_14742);
nand UO_1037 (O_1037,N_14261,N_14900);
or UO_1038 (O_1038,N_14355,N_14450);
or UO_1039 (O_1039,N_14310,N_14512);
and UO_1040 (O_1040,N_14713,N_14603);
nor UO_1041 (O_1041,N_14935,N_14948);
or UO_1042 (O_1042,N_14005,N_14710);
or UO_1043 (O_1043,N_14553,N_14739);
nand UO_1044 (O_1044,N_14649,N_14484);
and UO_1045 (O_1045,N_14070,N_14111);
xnor UO_1046 (O_1046,N_14425,N_14598);
nor UO_1047 (O_1047,N_14610,N_14592);
or UO_1048 (O_1048,N_14535,N_14981);
or UO_1049 (O_1049,N_14876,N_14070);
nand UO_1050 (O_1050,N_14506,N_14589);
nor UO_1051 (O_1051,N_14910,N_14052);
nand UO_1052 (O_1052,N_14961,N_14996);
and UO_1053 (O_1053,N_14357,N_14179);
or UO_1054 (O_1054,N_14869,N_14855);
nand UO_1055 (O_1055,N_14978,N_14263);
nor UO_1056 (O_1056,N_14103,N_14495);
nand UO_1057 (O_1057,N_14833,N_14402);
and UO_1058 (O_1058,N_14212,N_14329);
and UO_1059 (O_1059,N_14301,N_14017);
nand UO_1060 (O_1060,N_14424,N_14996);
xnor UO_1061 (O_1061,N_14185,N_14391);
and UO_1062 (O_1062,N_14948,N_14337);
nor UO_1063 (O_1063,N_14141,N_14296);
or UO_1064 (O_1064,N_14469,N_14588);
nor UO_1065 (O_1065,N_14094,N_14510);
or UO_1066 (O_1066,N_14127,N_14380);
nor UO_1067 (O_1067,N_14939,N_14967);
or UO_1068 (O_1068,N_14859,N_14103);
nand UO_1069 (O_1069,N_14829,N_14167);
xor UO_1070 (O_1070,N_14602,N_14106);
or UO_1071 (O_1071,N_14927,N_14907);
and UO_1072 (O_1072,N_14272,N_14262);
nor UO_1073 (O_1073,N_14997,N_14197);
nand UO_1074 (O_1074,N_14251,N_14949);
nor UO_1075 (O_1075,N_14425,N_14579);
nor UO_1076 (O_1076,N_14740,N_14244);
or UO_1077 (O_1077,N_14083,N_14657);
or UO_1078 (O_1078,N_14068,N_14500);
xnor UO_1079 (O_1079,N_14188,N_14938);
nand UO_1080 (O_1080,N_14129,N_14843);
nand UO_1081 (O_1081,N_14399,N_14376);
nand UO_1082 (O_1082,N_14239,N_14909);
nand UO_1083 (O_1083,N_14385,N_14043);
nor UO_1084 (O_1084,N_14908,N_14035);
and UO_1085 (O_1085,N_14364,N_14812);
xor UO_1086 (O_1086,N_14088,N_14219);
and UO_1087 (O_1087,N_14433,N_14265);
and UO_1088 (O_1088,N_14446,N_14176);
nor UO_1089 (O_1089,N_14602,N_14130);
and UO_1090 (O_1090,N_14198,N_14144);
nand UO_1091 (O_1091,N_14188,N_14843);
and UO_1092 (O_1092,N_14652,N_14051);
or UO_1093 (O_1093,N_14602,N_14190);
nand UO_1094 (O_1094,N_14496,N_14776);
and UO_1095 (O_1095,N_14822,N_14992);
nand UO_1096 (O_1096,N_14527,N_14170);
and UO_1097 (O_1097,N_14606,N_14359);
nor UO_1098 (O_1098,N_14589,N_14159);
nor UO_1099 (O_1099,N_14732,N_14675);
nand UO_1100 (O_1100,N_14617,N_14144);
nand UO_1101 (O_1101,N_14690,N_14026);
and UO_1102 (O_1102,N_14469,N_14903);
and UO_1103 (O_1103,N_14688,N_14385);
and UO_1104 (O_1104,N_14352,N_14503);
and UO_1105 (O_1105,N_14295,N_14537);
or UO_1106 (O_1106,N_14799,N_14663);
xor UO_1107 (O_1107,N_14314,N_14465);
or UO_1108 (O_1108,N_14559,N_14605);
xnor UO_1109 (O_1109,N_14739,N_14551);
nand UO_1110 (O_1110,N_14707,N_14611);
or UO_1111 (O_1111,N_14240,N_14389);
and UO_1112 (O_1112,N_14543,N_14097);
and UO_1113 (O_1113,N_14496,N_14114);
and UO_1114 (O_1114,N_14860,N_14715);
xnor UO_1115 (O_1115,N_14404,N_14481);
or UO_1116 (O_1116,N_14353,N_14630);
and UO_1117 (O_1117,N_14267,N_14219);
or UO_1118 (O_1118,N_14343,N_14457);
or UO_1119 (O_1119,N_14694,N_14584);
and UO_1120 (O_1120,N_14391,N_14499);
nor UO_1121 (O_1121,N_14564,N_14378);
nor UO_1122 (O_1122,N_14462,N_14852);
and UO_1123 (O_1123,N_14845,N_14860);
nor UO_1124 (O_1124,N_14753,N_14045);
or UO_1125 (O_1125,N_14713,N_14851);
nor UO_1126 (O_1126,N_14331,N_14658);
nand UO_1127 (O_1127,N_14105,N_14047);
nor UO_1128 (O_1128,N_14132,N_14948);
nor UO_1129 (O_1129,N_14550,N_14598);
nor UO_1130 (O_1130,N_14700,N_14936);
or UO_1131 (O_1131,N_14651,N_14947);
and UO_1132 (O_1132,N_14836,N_14292);
nor UO_1133 (O_1133,N_14560,N_14969);
nand UO_1134 (O_1134,N_14003,N_14783);
and UO_1135 (O_1135,N_14191,N_14985);
nand UO_1136 (O_1136,N_14718,N_14507);
and UO_1137 (O_1137,N_14425,N_14707);
or UO_1138 (O_1138,N_14608,N_14005);
xnor UO_1139 (O_1139,N_14592,N_14034);
nor UO_1140 (O_1140,N_14925,N_14857);
nor UO_1141 (O_1141,N_14797,N_14876);
or UO_1142 (O_1142,N_14037,N_14716);
nand UO_1143 (O_1143,N_14343,N_14291);
nand UO_1144 (O_1144,N_14454,N_14147);
nand UO_1145 (O_1145,N_14792,N_14462);
nand UO_1146 (O_1146,N_14679,N_14066);
and UO_1147 (O_1147,N_14129,N_14981);
nor UO_1148 (O_1148,N_14350,N_14023);
xnor UO_1149 (O_1149,N_14692,N_14311);
or UO_1150 (O_1150,N_14651,N_14000);
or UO_1151 (O_1151,N_14855,N_14199);
nor UO_1152 (O_1152,N_14812,N_14466);
nor UO_1153 (O_1153,N_14512,N_14274);
nor UO_1154 (O_1154,N_14984,N_14110);
and UO_1155 (O_1155,N_14908,N_14538);
nor UO_1156 (O_1156,N_14416,N_14941);
or UO_1157 (O_1157,N_14174,N_14763);
nand UO_1158 (O_1158,N_14510,N_14645);
or UO_1159 (O_1159,N_14650,N_14782);
or UO_1160 (O_1160,N_14757,N_14496);
or UO_1161 (O_1161,N_14780,N_14990);
and UO_1162 (O_1162,N_14400,N_14406);
or UO_1163 (O_1163,N_14395,N_14865);
nand UO_1164 (O_1164,N_14380,N_14338);
nor UO_1165 (O_1165,N_14025,N_14159);
xnor UO_1166 (O_1166,N_14773,N_14028);
or UO_1167 (O_1167,N_14126,N_14172);
nor UO_1168 (O_1168,N_14103,N_14665);
or UO_1169 (O_1169,N_14914,N_14265);
or UO_1170 (O_1170,N_14985,N_14824);
nand UO_1171 (O_1171,N_14873,N_14837);
nand UO_1172 (O_1172,N_14113,N_14629);
or UO_1173 (O_1173,N_14889,N_14966);
and UO_1174 (O_1174,N_14611,N_14408);
nor UO_1175 (O_1175,N_14922,N_14683);
nor UO_1176 (O_1176,N_14528,N_14481);
or UO_1177 (O_1177,N_14608,N_14576);
nand UO_1178 (O_1178,N_14000,N_14241);
nand UO_1179 (O_1179,N_14050,N_14492);
and UO_1180 (O_1180,N_14863,N_14650);
xor UO_1181 (O_1181,N_14585,N_14493);
nor UO_1182 (O_1182,N_14825,N_14512);
nand UO_1183 (O_1183,N_14550,N_14671);
nor UO_1184 (O_1184,N_14022,N_14743);
and UO_1185 (O_1185,N_14118,N_14824);
nor UO_1186 (O_1186,N_14757,N_14424);
nand UO_1187 (O_1187,N_14288,N_14867);
and UO_1188 (O_1188,N_14205,N_14350);
or UO_1189 (O_1189,N_14323,N_14367);
nand UO_1190 (O_1190,N_14126,N_14553);
nor UO_1191 (O_1191,N_14666,N_14128);
nor UO_1192 (O_1192,N_14600,N_14010);
and UO_1193 (O_1193,N_14311,N_14432);
nor UO_1194 (O_1194,N_14269,N_14722);
nor UO_1195 (O_1195,N_14596,N_14896);
nor UO_1196 (O_1196,N_14806,N_14026);
and UO_1197 (O_1197,N_14823,N_14300);
or UO_1198 (O_1198,N_14914,N_14049);
or UO_1199 (O_1199,N_14221,N_14023);
or UO_1200 (O_1200,N_14300,N_14757);
nand UO_1201 (O_1201,N_14236,N_14540);
nand UO_1202 (O_1202,N_14065,N_14109);
nor UO_1203 (O_1203,N_14610,N_14844);
nor UO_1204 (O_1204,N_14454,N_14103);
or UO_1205 (O_1205,N_14873,N_14233);
nand UO_1206 (O_1206,N_14742,N_14543);
nand UO_1207 (O_1207,N_14026,N_14428);
and UO_1208 (O_1208,N_14874,N_14988);
xnor UO_1209 (O_1209,N_14458,N_14971);
xor UO_1210 (O_1210,N_14229,N_14161);
xor UO_1211 (O_1211,N_14290,N_14293);
nor UO_1212 (O_1212,N_14032,N_14194);
or UO_1213 (O_1213,N_14448,N_14209);
and UO_1214 (O_1214,N_14280,N_14399);
xnor UO_1215 (O_1215,N_14214,N_14854);
or UO_1216 (O_1216,N_14780,N_14819);
and UO_1217 (O_1217,N_14843,N_14922);
nand UO_1218 (O_1218,N_14086,N_14287);
or UO_1219 (O_1219,N_14862,N_14265);
xnor UO_1220 (O_1220,N_14645,N_14650);
and UO_1221 (O_1221,N_14471,N_14467);
nand UO_1222 (O_1222,N_14478,N_14959);
nand UO_1223 (O_1223,N_14754,N_14429);
nor UO_1224 (O_1224,N_14653,N_14065);
nor UO_1225 (O_1225,N_14169,N_14178);
and UO_1226 (O_1226,N_14748,N_14344);
or UO_1227 (O_1227,N_14766,N_14675);
xor UO_1228 (O_1228,N_14808,N_14569);
nor UO_1229 (O_1229,N_14103,N_14216);
and UO_1230 (O_1230,N_14527,N_14671);
or UO_1231 (O_1231,N_14118,N_14783);
and UO_1232 (O_1232,N_14178,N_14416);
or UO_1233 (O_1233,N_14984,N_14425);
or UO_1234 (O_1234,N_14718,N_14888);
or UO_1235 (O_1235,N_14056,N_14786);
nor UO_1236 (O_1236,N_14938,N_14510);
and UO_1237 (O_1237,N_14522,N_14779);
or UO_1238 (O_1238,N_14194,N_14065);
xnor UO_1239 (O_1239,N_14672,N_14718);
xor UO_1240 (O_1240,N_14072,N_14557);
nand UO_1241 (O_1241,N_14686,N_14183);
nor UO_1242 (O_1242,N_14914,N_14350);
nand UO_1243 (O_1243,N_14604,N_14369);
and UO_1244 (O_1244,N_14167,N_14022);
nand UO_1245 (O_1245,N_14113,N_14067);
xnor UO_1246 (O_1246,N_14937,N_14568);
and UO_1247 (O_1247,N_14468,N_14455);
nand UO_1248 (O_1248,N_14112,N_14286);
or UO_1249 (O_1249,N_14289,N_14639);
and UO_1250 (O_1250,N_14836,N_14674);
nor UO_1251 (O_1251,N_14292,N_14871);
and UO_1252 (O_1252,N_14937,N_14234);
nand UO_1253 (O_1253,N_14014,N_14531);
nor UO_1254 (O_1254,N_14053,N_14420);
nor UO_1255 (O_1255,N_14164,N_14870);
xor UO_1256 (O_1256,N_14779,N_14980);
or UO_1257 (O_1257,N_14856,N_14641);
or UO_1258 (O_1258,N_14884,N_14146);
or UO_1259 (O_1259,N_14794,N_14775);
nor UO_1260 (O_1260,N_14227,N_14691);
nand UO_1261 (O_1261,N_14500,N_14250);
and UO_1262 (O_1262,N_14709,N_14488);
and UO_1263 (O_1263,N_14213,N_14144);
nand UO_1264 (O_1264,N_14128,N_14124);
nand UO_1265 (O_1265,N_14025,N_14776);
and UO_1266 (O_1266,N_14967,N_14733);
nand UO_1267 (O_1267,N_14670,N_14841);
xor UO_1268 (O_1268,N_14330,N_14935);
nor UO_1269 (O_1269,N_14753,N_14633);
nand UO_1270 (O_1270,N_14180,N_14978);
or UO_1271 (O_1271,N_14059,N_14990);
or UO_1272 (O_1272,N_14673,N_14738);
nand UO_1273 (O_1273,N_14516,N_14560);
nand UO_1274 (O_1274,N_14159,N_14683);
nand UO_1275 (O_1275,N_14436,N_14010);
and UO_1276 (O_1276,N_14814,N_14458);
nand UO_1277 (O_1277,N_14779,N_14786);
or UO_1278 (O_1278,N_14709,N_14459);
xor UO_1279 (O_1279,N_14240,N_14528);
or UO_1280 (O_1280,N_14360,N_14726);
nand UO_1281 (O_1281,N_14534,N_14375);
nand UO_1282 (O_1282,N_14729,N_14588);
and UO_1283 (O_1283,N_14112,N_14554);
or UO_1284 (O_1284,N_14961,N_14184);
or UO_1285 (O_1285,N_14113,N_14934);
or UO_1286 (O_1286,N_14956,N_14316);
nor UO_1287 (O_1287,N_14875,N_14646);
nand UO_1288 (O_1288,N_14333,N_14142);
and UO_1289 (O_1289,N_14296,N_14664);
and UO_1290 (O_1290,N_14407,N_14296);
nor UO_1291 (O_1291,N_14820,N_14625);
and UO_1292 (O_1292,N_14348,N_14870);
and UO_1293 (O_1293,N_14986,N_14686);
and UO_1294 (O_1294,N_14386,N_14977);
nor UO_1295 (O_1295,N_14138,N_14570);
xnor UO_1296 (O_1296,N_14978,N_14540);
or UO_1297 (O_1297,N_14685,N_14401);
or UO_1298 (O_1298,N_14863,N_14364);
or UO_1299 (O_1299,N_14542,N_14106);
nor UO_1300 (O_1300,N_14329,N_14046);
or UO_1301 (O_1301,N_14588,N_14377);
nor UO_1302 (O_1302,N_14533,N_14978);
and UO_1303 (O_1303,N_14252,N_14411);
nand UO_1304 (O_1304,N_14748,N_14016);
nand UO_1305 (O_1305,N_14527,N_14380);
and UO_1306 (O_1306,N_14919,N_14608);
nor UO_1307 (O_1307,N_14009,N_14923);
or UO_1308 (O_1308,N_14874,N_14568);
nor UO_1309 (O_1309,N_14205,N_14027);
and UO_1310 (O_1310,N_14954,N_14715);
xnor UO_1311 (O_1311,N_14760,N_14545);
nand UO_1312 (O_1312,N_14453,N_14432);
or UO_1313 (O_1313,N_14047,N_14554);
or UO_1314 (O_1314,N_14420,N_14782);
nand UO_1315 (O_1315,N_14306,N_14237);
nor UO_1316 (O_1316,N_14444,N_14094);
and UO_1317 (O_1317,N_14127,N_14714);
nor UO_1318 (O_1318,N_14358,N_14550);
nand UO_1319 (O_1319,N_14128,N_14294);
or UO_1320 (O_1320,N_14419,N_14683);
nand UO_1321 (O_1321,N_14907,N_14271);
and UO_1322 (O_1322,N_14533,N_14487);
or UO_1323 (O_1323,N_14547,N_14353);
or UO_1324 (O_1324,N_14637,N_14754);
xnor UO_1325 (O_1325,N_14887,N_14890);
nand UO_1326 (O_1326,N_14918,N_14132);
or UO_1327 (O_1327,N_14688,N_14926);
xnor UO_1328 (O_1328,N_14688,N_14256);
nand UO_1329 (O_1329,N_14911,N_14419);
nor UO_1330 (O_1330,N_14120,N_14155);
and UO_1331 (O_1331,N_14809,N_14059);
nor UO_1332 (O_1332,N_14240,N_14502);
nand UO_1333 (O_1333,N_14064,N_14446);
and UO_1334 (O_1334,N_14393,N_14174);
nor UO_1335 (O_1335,N_14102,N_14073);
and UO_1336 (O_1336,N_14908,N_14686);
nor UO_1337 (O_1337,N_14004,N_14430);
and UO_1338 (O_1338,N_14501,N_14000);
nor UO_1339 (O_1339,N_14115,N_14805);
or UO_1340 (O_1340,N_14321,N_14369);
nor UO_1341 (O_1341,N_14185,N_14974);
xor UO_1342 (O_1342,N_14443,N_14548);
and UO_1343 (O_1343,N_14439,N_14829);
nor UO_1344 (O_1344,N_14989,N_14576);
nor UO_1345 (O_1345,N_14242,N_14890);
xnor UO_1346 (O_1346,N_14868,N_14343);
xor UO_1347 (O_1347,N_14289,N_14085);
and UO_1348 (O_1348,N_14730,N_14820);
and UO_1349 (O_1349,N_14106,N_14191);
xnor UO_1350 (O_1350,N_14223,N_14120);
or UO_1351 (O_1351,N_14686,N_14800);
xnor UO_1352 (O_1352,N_14548,N_14313);
xnor UO_1353 (O_1353,N_14964,N_14949);
or UO_1354 (O_1354,N_14473,N_14440);
nand UO_1355 (O_1355,N_14600,N_14860);
nor UO_1356 (O_1356,N_14038,N_14197);
nand UO_1357 (O_1357,N_14136,N_14567);
and UO_1358 (O_1358,N_14844,N_14797);
nand UO_1359 (O_1359,N_14845,N_14922);
nand UO_1360 (O_1360,N_14278,N_14564);
and UO_1361 (O_1361,N_14852,N_14348);
nor UO_1362 (O_1362,N_14006,N_14858);
nor UO_1363 (O_1363,N_14819,N_14446);
xor UO_1364 (O_1364,N_14472,N_14558);
and UO_1365 (O_1365,N_14297,N_14881);
nor UO_1366 (O_1366,N_14883,N_14688);
or UO_1367 (O_1367,N_14166,N_14680);
nor UO_1368 (O_1368,N_14875,N_14624);
xor UO_1369 (O_1369,N_14721,N_14384);
and UO_1370 (O_1370,N_14767,N_14581);
or UO_1371 (O_1371,N_14142,N_14929);
nor UO_1372 (O_1372,N_14600,N_14997);
nand UO_1373 (O_1373,N_14288,N_14127);
nor UO_1374 (O_1374,N_14713,N_14690);
nor UO_1375 (O_1375,N_14687,N_14271);
nor UO_1376 (O_1376,N_14107,N_14524);
nand UO_1377 (O_1377,N_14463,N_14055);
xnor UO_1378 (O_1378,N_14653,N_14807);
or UO_1379 (O_1379,N_14663,N_14710);
and UO_1380 (O_1380,N_14832,N_14665);
nand UO_1381 (O_1381,N_14555,N_14156);
or UO_1382 (O_1382,N_14974,N_14476);
nor UO_1383 (O_1383,N_14638,N_14620);
nor UO_1384 (O_1384,N_14564,N_14056);
or UO_1385 (O_1385,N_14069,N_14551);
xnor UO_1386 (O_1386,N_14805,N_14517);
nand UO_1387 (O_1387,N_14853,N_14841);
or UO_1388 (O_1388,N_14475,N_14049);
nand UO_1389 (O_1389,N_14844,N_14724);
or UO_1390 (O_1390,N_14739,N_14329);
and UO_1391 (O_1391,N_14473,N_14798);
nor UO_1392 (O_1392,N_14047,N_14293);
and UO_1393 (O_1393,N_14407,N_14006);
xor UO_1394 (O_1394,N_14686,N_14338);
nand UO_1395 (O_1395,N_14061,N_14254);
nor UO_1396 (O_1396,N_14746,N_14627);
xor UO_1397 (O_1397,N_14645,N_14029);
nor UO_1398 (O_1398,N_14866,N_14736);
nor UO_1399 (O_1399,N_14243,N_14031);
nand UO_1400 (O_1400,N_14009,N_14673);
nand UO_1401 (O_1401,N_14165,N_14286);
nor UO_1402 (O_1402,N_14833,N_14027);
or UO_1403 (O_1403,N_14211,N_14460);
nor UO_1404 (O_1404,N_14187,N_14578);
or UO_1405 (O_1405,N_14780,N_14504);
nor UO_1406 (O_1406,N_14231,N_14735);
or UO_1407 (O_1407,N_14489,N_14866);
nand UO_1408 (O_1408,N_14863,N_14459);
or UO_1409 (O_1409,N_14593,N_14989);
and UO_1410 (O_1410,N_14258,N_14698);
nor UO_1411 (O_1411,N_14445,N_14168);
nor UO_1412 (O_1412,N_14324,N_14262);
and UO_1413 (O_1413,N_14633,N_14245);
and UO_1414 (O_1414,N_14145,N_14082);
and UO_1415 (O_1415,N_14890,N_14354);
xnor UO_1416 (O_1416,N_14444,N_14244);
nor UO_1417 (O_1417,N_14804,N_14177);
or UO_1418 (O_1418,N_14234,N_14695);
and UO_1419 (O_1419,N_14766,N_14774);
or UO_1420 (O_1420,N_14207,N_14632);
and UO_1421 (O_1421,N_14982,N_14016);
and UO_1422 (O_1422,N_14950,N_14009);
or UO_1423 (O_1423,N_14723,N_14977);
or UO_1424 (O_1424,N_14937,N_14802);
nand UO_1425 (O_1425,N_14582,N_14304);
and UO_1426 (O_1426,N_14545,N_14849);
or UO_1427 (O_1427,N_14800,N_14987);
or UO_1428 (O_1428,N_14859,N_14712);
nand UO_1429 (O_1429,N_14809,N_14386);
and UO_1430 (O_1430,N_14173,N_14088);
or UO_1431 (O_1431,N_14419,N_14726);
and UO_1432 (O_1432,N_14885,N_14386);
nand UO_1433 (O_1433,N_14670,N_14484);
or UO_1434 (O_1434,N_14431,N_14792);
xnor UO_1435 (O_1435,N_14322,N_14376);
and UO_1436 (O_1436,N_14641,N_14070);
or UO_1437 (O_1437,N_14203,N_14119);
and UO_1438 (O_1438,N_14238,N_14980);
nand UO_1439 (O_1439,N_14878,N_14225);
or UO_1440 (O_1440,N_14828,N_14647);
and UO_1441 (O_1441,N_14391,N_14014);
or UO_1442 (O_1442,N_14815,N_14605);
and UO_1443 (O_1443,N_14514,N_14595);
nand UO_1444 (O_1444,N_14038,N_14033);
nand UO_1445 (O_1445,N_14336,N_14179);
nand UO_1446 (O_1446,N_14594,N_14397);
xor UO_1447 (O_1447,N_14436,N_14422);
and UO_1448 (O_1448,N_14301,N_14722);
or UO_1449 (O_1449,N_14137,N_14241);
or UO_1450 (O_1450,N_14040,N_14079);
xor UO_1451 (O_1451,N_14672,N_14362);
nor UO_1452 (O_1452,N_14097,N_14900);
or UO_1453 (O_1453,N_14611,N_14287);
nand UO_1454 (O_1454,N_14094,N_14593);
or UO_1455 (O_1455,N_14851,N_14131);
or UO_1456 (O_1456,N_14950,N_14764);
nor UO_1457 (O_1457,N_14539,N_14449);
nor UO_1458 (O_1458,N_14544,N_14479);
or UO_1459 (O_1459,N_14760,N_14541);
nor UO_1460 (O_1460,N_14085,N_14044);
and UO_1461 (O_1461,N_14458,N_14464);
xor UO_1462 (O_1462,N_14146,N_14101);
nor UO_1463 (O_1463,N_14248,N_14939);
and UO_1464 (O_1464,N_14603,N_14104);
xnor UO_1465 (O_1465,N_14055,N_14189);
and UO_1466 (O_1466,N_14909,N_14833);
nand UO_1467 (O_1467,N_14782,N_14409);
nor UO_1468 (O_1468,N_14318,N_14044);
and UO_1469 (O_1469,N_14533,N_14180);
and UO_1470 (O_1470,N_14429,N_14175);
or UO_1471 (O_1471,N_14439,N_14075);
or UO_1472 (O_1472,N_14391,N_14926);
xor UO_1473 (O_1473,N_14699,N_14811);
nor UO_1474 (O_1474,N_14773,N_14319);
nor UO_1475 (O_1475,N_14277,N_14343);
nand UO_1476 (O_1476,N_14527,N_14190);
and UO_1477 (O_1477,N_14524,N_14639);
nand UO_1478 (O_1478,N_14813,N_14282);
or UO_1479 (O_1479,N_14406,N_14485);
xnor UO_1480 (O_1480,N_14927,N_14344);
or UO_1481 (O_1481,N_14585,N_14180);
nand UO_1482 (O_1482,N_14759,N_14794);
xnor UO_1483 (O_1483,N_14109,N_14014);
and UO_1484 (O_1484,N_14364,N_14404);
or UO_1485 (O_1485,N_14530,N_14402);
nand UO_1486 (O_1486,N_14787,N_14370);
and UO_1487 (O_1487,N_14531,N_14994);
nand UO_1488 (O_1488,N_14883,N_14553);
nand UO_1489 (O_1489,N_14857,N_14968);
or UO_1490 (O_1490,N_14409,N_14279);
nor UO_1491 (O_1491,N_14302,N_14793);
nand UO_1492 (O_1492,N_14795,N_14971);
nand UO_1493 (O_1493,N_14331,N_14259);
nor UO_1494 (O_1494,N_14646,N_14489);
nor UO_1495 (O_1495,N_14883,N_14314);
and UO_1496 (O_1496,N_14396,N_14872);
or UO_1497 (O_1497,N_14016,N_14093);
and UO_1498 (O_1498,N_14122,N_14355);
nand UO_1499 (O_1499,N_14959,N_14767);
or UO_1500 (O_1500,N_14741,N_14236);
and UO_1501 (O_1501,N_14102,N_14390);
and UO_1502 (O_1502,N_14346,N_14585);
and UO_1503 (O_1503,N_14886,N_14446);
or UO_1504 (O_1504,N_14597,N_14626);
and UO_1505 (O_1505,N_14810,N_14870);
or UO_1506 (O_1506,N_14600,N_14046);
nand UO_1507 (O_1507,N_14301,N_14417);
xor UO_1508 (O_1508,N_14617,N_14827);
or UO_1509 (O_1509,N_14960,N_14566);
nand UO_1510 (O_1510,N_14617,N_14175);
nor UO_1511 (O_1511,N_14021,N_14536);
xnor UO_1512 (O_1512,N_14780,N_14894);
nor UO_1513 (O_1513,N_14554,N_14236);
nor UO_1514 (O_1514,N_14459,N_14527);
nor UO_1515 (O_1515,N_14879,N_14974);
nor UO_1516 (O_1516,N_14976,N_14921);
nand UO_1517 (O_1517,N_14780,N_14084);
and UO_1518 (O_1518,N_14132,N_14182);
nand UO_1519 (O_1519,N_14817,N_14794);
nand UO_1520 (O_1520,N_14084,N_14340);
nor UO_1521 (O_1521,N_14827,N_14222);
nor UO_1522 (O_1522,N_14577,N_14321);
nor UO_1523 (O_1523,N_14708,N_14511);
xnor UO_1524 (O_1524,N_14343,N_14951);
nand UO_1525 (O_1525,N_14778,N_14984);
or UO_1526 (O_1526,N_14181,N_14416);
xnor UO_1527 (O_1527,N_14343,N_14105);
nand UO_1528 (O_1528,N_14969,N_14887);
nor UO_1529 (O_1529,N_14102,N_14178);
and UO_1530 (O_1530,N_14355,N_14820);
nand UO_1531 (O_1531,N_14999,N_14616);
or UO_1532 (O_1532,N_14267,N_14855);
nand UO_1533 (O_1533,N_14293,N_14173);
nand UO_1534 (O_1534,N_14443,N_14516);
nor UO_1535 (O_1535,N_14645,N_14361);
nor UO_1536 (O_1536,N_14964,N_14716);
nand UO_1537 (O_1537,N_14692,N_14121);
nand UO_1538 (O_1538,N_14807,N_14580);
or UO_1539 (O_1539,N_14553,N_14376);
xnor UO_1540 (O_1540,N_14707,N_14005);
nand UO_1541 (O_1541,N_14335,N_14225);
nand UO_1542 (O_1542,N_14023,N_14697);
or UO_1543 (O_1543,N_14161,N_14955);
and UO_1544 (O_1544,N_14771,N_14979);
nor UO_1545 (O_1545,N_14256,N_14697);
or UO_1546 (O_1546,N_14603,N_14148);
nor UO_1547 (O_1547,N_14205,N_14139);
nand UO_1548 (O_1548,N_14179,N_14907);
nor UO_1549 (O_1549,N_14369,N_14010);
nand UO_1550 (O_1550,N_14196,N_14860);
xor UO_1551 (O_1551,N_14275,N_14784);
and UO_1552 (O_1552,N_14934,N_14624);
and UO_1553 (O_1553,N_14237,N_14086);
and UO_1554 (O_1554,N_14685,N_14080);
and UO_1555 (O_1555,N_14389,N_14383);
and UO_1556 (O_1556,N_14084,N_14391);
nor UO_1557 (O_1557,N_14844,N_14388);
and UO_1558 (O_1558,N_14429,N_14675);
and UO_1559 (O_1559,N_14668,N_14442);
or UO_1560 (O_1560,N_14465,N_14144);
nor UO_1561 (O_1561,N_14201,N_14047);
or UO_1562 (O_1562,N_14057,N_14782);
xnor UO_1563 (O_1563,N_14265,N_14299);
nor UO_1564 (O_1564,N_14045,N_14783);
nor UO_1565 (O_1565,N_14379,N_14206);
or UO_1566 (O_1566,N_14304,N_14351);
nor UO_1567 (O_1567,N_14856,N_14061);
xnor UO_1568 (O_1568,N_14617,N_14917);
nor UO_1569 (O_1569,N_14787,N_14468);
nor UO_1570 (O_1570,N_14110,N_14288);
and UO_1571 (O_1571,N_14832,N_14924);
and UO_1572 (O_1572,N_14845,N_14043);
and UO_1573 (O_1573,N_14598,N_14634);
nand UO_1574 (O_1574,N_14516,N_14783);
or UO_1575 (O_1575,N_14364,N_14888);
nand UO_1576 (O_1576,N_14997,N_14712);
and UO_1577 (O_1577,N_14595,N_14495);
and UO_1578 (O_1578,N_14295,N_14224);
nand UO_1579 (O_1579,N_14124,N_14792);
nor UO_1580 (O_1580,N_14620,N_14055);
xor UO_1581 (O_1581,N_14145,N_14592);
or UO_1582 (O_1582,N_14134,N_14580);
or UO_1583 (O_1583,N_14730,N_14731);
nor UO_1584 (O_1584,N_14740,N_14248);
or UO_1585 (O_1585,N_14786,N_14563);
or UO_1586 (O_1586,N_14148,N_14027);
or UO_1587 (O_1587,N_14005,N_14273);
nand UO_1588 (O_1588,N_14215,N_14901);
and UO_1589 (O_1589,N_14573,N_14744);
nor UO_1590 (O_1590,N_14287,N_14214);
nand UO_1591 (O_1591,N_14850,N_14634);
nor UO_1592 (O_1592,N_14817,N_14075);
nand UO_1593 (O_1593,N_14215,N_14957);
nor UO_1594 (O_1594,N_14196,N_14786);
nand UO_1595 (O_1595,N_14823,N_14294);
nor UO_1596 (O_1596,N_14607,N_14679);
or UO_1597 (O_1597,N_14498,N_14724);
or UO_1598 (O_1598,N_14415,N_14303);
nand UO_1599 (O_1599,N_14463,N_14895);
and UO_1600 (O_1600,N_14841,N_14407);
and UO_1601 (O_1601,N_14295,N_14055);
nor UO_1602 (O_1602,N_14931,N_14181);
xor UO_1603 (O_1603,N_14333,N_14165);
and UO_1604 (O_1604,N_14219,N_14093);
nor UO_1605 (O_1605,N_14423,N_14021);
xnor UO_1606 (O_1606,N_14395,N_14271);
nor UO_1607 (O_1607,N_14983,N_14243);
nand UO_1608 (O_1608,N_14076,N_14602);
nand UO_1609 (O_1609,N_14646,N_14422);
or UO_1610 (O_1610,N_14740,N_14883);
nand UO_1611 (O_1611,N_14702,N_14046);
and UO_1612 (O_1612,N_14605,N_14996);
and UO_1613 (O_1613,N_14004,N_14136);
and UO_1614 (O_1614,N_14267,N_14778);
or UO_1615 (O_1615,N_14854,N_14297);
and UO_1616 (O_1616,N_14047,N_14726);
or UO_1617 (O_1617,N_14373,N_14937);
or UO_1618 (O_1618,N_14605,N_14664);
nand UO_1619 (O_1619,N_14372,N_14100);
nand UO_1620 (O_1620,N_14948,N_14802);
and UO_1621 (O_1621,N_14050,N_14324);
xnor UO_1622 (O_1622,N_14449,N_14345);
xnor UO_1623 (O_1623,N_14932,N_14682);
and UO_1624 (O_1624,N_14639,N_14598);
nand UO_1625 (O_1625,N_14969,N_14756);
nand UO_1626 (O_1626,N_14658,N_14894);
and UO_1627 (O_1627,N_14345,N_14019);
and UO_1628 (O_1628,N_14943,N_14831);
and UO_1629 (O_1629,N_14031,N_14267);
nor UO_1630 (O_1630,N_14100,N_14823);
or UO_1631 (O_1631,N_14764,N_14220);
nand UO_1632 (O_1632,N_14527,N_14144);
nand UO_1633 (O_1633,N_14467,N_14604);
xor UO_1634 (O_1634,N_14481,N_14421);
nand UO_1635 (O_1635,N_14907,N_14172);
nor UO_1636 (O_1636,N_14761,N_14196);
and UO_1637 (O_1637,N_14751,N_14442);
nor UO_1638 (O_1638,N_14254,N_14986);
and UO_1639 (O_1639,N_14606,N_14960);
or UO_1640 (O_1640,N_14876,N_14465);
nand UO_1641 (O_1641,N_14859,N_14097);
nand UO_1642 (O_1642,N_14211,N_14349);
nand UO_1643 (O_1643,N_14453,N_14326);
nand UO_1644 (O_1644,N_14134,N_14229);
and UO_1645 (O_1645,N_14000,N_14997);
xnor UO_1646 (O_1646,N_14919,N_14278);
and UO_1647 (O_1647,N_14267,N_14808);
nor UO_1648 (O_1648,N_14144,N_14653);
nand UO_1649 (O_1649,N_14686,N_14397);
nand UO_1650 (O_1650,N_14524,N_14205);
and UO_1651 (O_1651,N_14882,N_14102);
nor UO_1652 (O_1652,N_14358,N_14300);
xnor UO_1653 (O_1653,N_14495,N_14852);
or UO_1654 (O_1654,N_14502,N_14791);
nand UO_1655 (O_1655,N_14640,N_14621);
and UO_1656 (O_1656,N_14012,N_14269);
or UO_1657 (O_1657,N_14717,N_14874);
or UO_1658 (O_1658,N_14083,N_14559);
and UO_1659 (O_1659,N_14372,N_14151);
or UO_1660 (O_1660,N_14598,N_14733);
and UO_1661 (O_1661,N_14231,N_14342);
nor UO_1662 (O_1662,N_14092,N_14412);
nand UO_1663 (O_1663,N_14667,N_14767);
nor UO_1664 (O_1664,N_14944,N_14415);
nor UO_1665 (O_1665,N_14842,N_14831);
or UO_1666 (O_1666,N_14615,N_14070);
xnor UO_1667 (O_1667,N_14149,N_14664);
and UO_1668 (O_1668,N_14250,N_14417);
or UO_1669 (O_1669,N_14213,N_14849);
nand UO_1670 (O_1670,N_14663,N_14008);
or UO_1671 (O_1671,N_14569,N_14749);
nand UO_1672 (O_1672,N_14169,N_14478);
and UO_1673 (O_1673,N_14819,N_14345);
and UO_1674 (O_1674,N_14353,N_14528);
or UO_1675 (O_1675,N_14985,N_14063);
and UO_1676 (O_1676,N_14685,N_14472);
xnor UO_1677 (O_1677,N_14845,N_14590);
and UO_1678 (O_1678,N_14345,N_14710);
nand UO_1679 (O_1679,N_14085,N_14035);
or UO_1680 (O_1680,N_14243,N_14276);
or UO_1681 (O_1681,N_14539,N_14203);
or UO_1682 (O_1682,N_14012,N_14844);
nor UO_1683 (O_1683,N_14490,N_14936);
nand UO_1684 (O_1684,N_14310,N_14200);
nor UO_1685 (O_1685,N_14442,N_14607);
nand UO_1686 (O_1686,N_14395,N_14338);
nand UO_1687 (O_1687,N_14189,N_14980);
or UO_1688 (O_1688,N_14753,N_14439);
or UO_1689 (O_1689,N_14059,N_14918);
and UO_1690 (O_1690,N_14917,N_14654);
and UO_1691 (O_1691,N_14133,N_14621);
or UO_1692 (O_1692,N_14472,N_14210);
and UO_1693 (O_1693,N_14448,N_14116);
or UO_1694 (O_1694,N_14938,N_14123);
and UO_1695 (O_1695,N_14794,N_14075);
xor UO_1696 (O_1696,N_14838,N_14278);
nand UO_1697 (O_1697,N_14873,N_14399);
nand UO_1698 (O_1698,N_14435,N_14738);
xor UO_1699 (O_1699,N_14304,N_14720);
nand UO_1700 (O_1700,N_14265,N_14685);
or UO_1701 (O_1701,N_14135,N_14621);
nor UO_1702 (O_1702,N_14562,N_14886);
nor UO_1703 (O_1703,N_14928,N_14508);
and UO_1704 (O_1704,N_14850,N_14269);
nand UO_1705 (O_1705,N_14448,N_14428);
and UO_1706 (O_1706,N_14559,N_14381);
xor UO_1707 (O_1707,N_14155,N_14096);
nand UO_1708 (O_1708,N_14262,N_14773);
nor UO_1709 (O_1709,N_14534,N_14368);
xor UO_1710 (O_1710,N_14187,N_14841);
xnor UO_1711 (O_1711,N_14119,N_14761);
nand UO_1712 (O_1712,N_14594,N_14031);
and UO_1713 (O_1713,N_14055,N_14085);
xor UO_1714 (O_1714,N_14207,N_14325);
nand UO_1715 (O_1715,N_14027,N_14171);
and UO_1716 (O_1716,N_14907,N_14888);
nand UO_1717 (O_1717,N_14842,N_14144);
nand UO_1718 (O_1718,N_14988,N_14735);
nor UO_1719 (O_1719,N_14049,N_14817);
nor UO_1720 (O_1720,N_14379,N_14502);
or UO_1721 (O_1721,N_14779,N_14258);
nor UO_1722 (O_1722,N_14419,N_14106);
nand UO_1723 (O_1723,N_14330,N_14372);
and UO_1724 (O_1724,N_14132,N_14597);
nor UO_1725 (O_1725,N_14894,N_14809);
nand UO_1726 (O_1726,N_14794,N_14664);
nor UO_1727 (O_1727,N_14461,N_14682);
and UO_1728 (O_1728,N_14715,N_14911);
or UO_1729 (O_1729,N_14779,N_14358);
nand UO_1730 (O_1730,N_14627,N_14319);
nor UO_1731 (O_1731,N_14728,N_14060);
nand UO_1732 (O_1732,N_14221,N_14388);
nand UO_1733 (O_1733,N_14617,N_14963);
or UO_1734 (O_1734,N_14024,N_14844);
or UO_1735 (O_1735,N_14995,N_14989);
and UO_1736 (O_1736,N_14340,N_14207);
or UO_1737 (O_1737,N_14124,N_14836);
or UO_1738 (O_1738,N_14441,N_14014);
nor UO_1739 (O_1739,N_14409,N_14624);
and UO_1740 (O_1740,N_14162,N_14993);
nor UO_1741 (O_1741,N_14556,N_14503);
nor UO_1742 (O_1742,N_14281,N_14869);
nor UO_1743 (O_1743,N_14198,N_14874);
nor UO_1744 (O_1744,N_14687,N_14872);
nor UO_1745 (O_1745,N_14269,N_14378);
nand UO_1746 (O_1746,N_14469,N_14099);
or UO_1747 (O_1747,N_14923,N_14766);
or UO_1748 (O_1748,N_14329,N_14887);
and UO_1749 (O_1749,N_14788,N_14188);
nand UO_1750 (O_1750,N_14412,N_14086);
nand UO_1751 (O_1751,N_14049,N_14345);
or UO_1752 (O_1752,N_14448,N_14947);
nand UO_1753 (O_1753,N_14733,N_14263);
nand UO_1754 (O_1754,N_14614,N_14211);
nand UO_1755 (O_1755,N_14298,N_14785);
and UO_1756 (O_1756,N_14929,N_14785);
or UO_1757 (O_1757,N_14259,N_14126);
nand UO_1758 (O_1758,N_14768,N_14517);
nor UO_1759 (O_1759,N_14987,N_14156);
nor UO_1760 (O_1760,N_14144,N_14608);
nor UO_1761 (O_1761,N_14179,N_14792);
and UO_1762 (O_1762,N_14697,N_14012);
nor UO_1763 (O_1763,N_14213,N_14285);
nand UO_1764 (O_1764,N_14297,N_14183);
nor UO_1765 (O_1765,N_14566,N_14985);
or UO_1766 (O_1766,N_14188,N_14680);
xnor UO_1767 (O_1767,N_14207,N_14800);
and UO_1768 (O_1768,N_14752,N_14098);
nor UO_1769 (O_1769,N_14946,N_14182);
nor UO_1770 (O_1770,N_14034,N_14703);
nor UO_1771 (O_1771,N_14184,N_14936);
nand UO_1772 (O_1772,N_14780,N_14969);
nand UO_1773 (O_1773,N_14351,N_14959);
or UO_1774 (O_1774,N_14616,N_14452);
nand UO_1775 (O_1775,N_14963,N_14007);
and UO_1776 (O_1776,N_14790,N_14924);
and UO_1777 (O_1777,N_14561,N_14075);
nor UO_1778 (O_1778,N_14305,N_14518);
and UO_1779 (O_1779,N_14921,N_14171);
or UO_1780 (O_1780,N_14474,N_14250);
or UO_1781 (O_1781,N_14904,N_14252);
or UO_1782 (O_1782,N_14437,N_14966);
nand UO_1783 (O_1783,N_14608,N_14571);
nand UO_1784 (O_1784,N_14636,N_14416);
nor UO_1785 (O_1785,N_14022,N_14058);
and UO_1786 (O_1786,N_14020,N_14642);
nand UO_1787 (O_1787,N_14636,N_14988);
and UO_1788 (O_1788,N_14762,N_14382);
or UO_1789 (O_1789,N_14697,N_14562);
and UO_1790 (O_1790,N_14375,N_14390);
xor UO_1791 (O_1791,N_14132,N_14520);
xnor UO_1792 (O_1792,N_14663,N_14445);
nand UO_1793 (O_1793,N_14581,N_14381);
and UO_1794 (O_1794,N_14140,N_14945);
xor UO_1795 (O_1795,N_14982,N_14315);
nor UO_1796 (O_1796,N_14813,N_14046);
or UO_1797 (O_1797,N_14825,N_14908);
nand UO_1798 (O_1798,N_14926,N_14555);
and UO_1799 (O_1799,N_14824,N_14449);
or UO_1800 (O_1800,N_14939,N_14562);
or UO_1801 (O_1801,N_14905,N_14123);
nor UO_1802 (O_1802,N_14303,N_14668);
nand UO_1803 (O_1803,N_14587,N_14030);
and UO_1804 (O_1804,N_14280,N_14160);
nor UO_1805 (O_1805,N_14757,N_14994);
nor UO_1806 (O_1806,N_14686,N_14238);
or UO_1807 (O_1807,N_14445,N_14862);
nor UO_1808 (O_1808,N_14812,N_14235);
nand UO_1809 (O_1809,N_14563,N_14759);
and UO_1810 (O_1810,N_14631,N_14262);
nand UO_1811 (O_1811,N_14345,N_14395);
or UO_1812 (O_1812,N_14938,N_14173);
and UO_1813 (O_1813,N_14908,N_14005);
or UO_1814 (O_1814,N_14558,N_14845);
nor UO_1815 (O_1815,N_14660,N_14545);
and UO_1816 (O_1816,N_14220,N_14115);
xnor UO_1817 (O_1817,N_14692,N_14819);
or UO_1818 (O_1818,N_14053,N_14707);
nor UO_1819 (O_1819,N_14858,N_14600);
and UO_1820 (O_1820,N_14663,N_14390);
nor UO_1821 (O_1821,N_14742,N_14926);
xor UO_1822 (O_1822,N_14959,N_14026);
xnor UO_1823 (O_1823,N_14801,N_14026);
and UO_1824 (O_1824,N_14370,N_14793);
xnor UO_1825 (O_1825,N_14564,N_14211);
nor UO_1826 (O_1826,N_14723,N_14743);
xor UO_1827 (O_1827,N_14662,N_14761);
or UO_1828 (O_1828,N_14894,N_14057);
and UO_1829 (O_1829,N_14373,N_14389);
and UO_1830 (O_1830,N_14389,N_14633);
or UO_1831 (O_1831,N_14149,N_14096);
or UO_1832 (O_1832,N_14166,N_14828);
xnor UO_1833 (O_1833,N_14697,N_14098);
nor UO_1834 (O_1834,N_14110,N_14080);
and UO_1835 (O_1835,N_14819,N_14289);
and UO_1836 (O_1836,N_14596,N_14033);
nand UO_1837 (O_1837,N_14437,N_14275);
and UO_1838 (O_1838,N_14916,N_14920);
nor UO_1839 (O_1839,N_14830,N_14688);
nor UO_1840 (O_1840,N_14626,N_14908);
or UO_1841 (O_1841,N_14340,N_14165);
nor UO_1842 (O_1842,N_14042,N_14918);
nand UO_1843 (O_1843,N_14256,N_14300);
nand UO_1844 (O_1844,N_14416,N_14841);
nor UO_1845 (O_1845,N_14522,N_14471);
nor UO_1846 (O_1846,N_14609,N_14331);
and UO_1847 (O_1847,N_14480,N_14331);
xnor UO_1848 (O_1848,N_14587,N_14502);
or UO_1849 (O_1849,N_14456,N_14094);
nand UO_1850 (O_1850,N_14149,N_14365);
or UO_1851 (O_1851,N_14505,N_14840);
nor UO_1852 (O_1852,N_14455,N_14221);
nor UO_1853 (O_1853,N_14268,N_14126);
nor UO_1854 (O_1854,N_14610,N_14289);
nor UO_1855 (O_1855,N_14166,N_14374);
and UO_1856 (O_1856,N_14541,N_14801);
nand UO_1857 (O_1857,N_14229,N_14689);
or UO_1858 (O_1858,N_14583,N_14204);
nor UO_1859 (O_1859,N_14867,N_14738);
nor UO_1860 (O_1860,N_14428,N_14979);
and UO_1861 (O_1861,N_14583,N_14377);
xnor UO_1862 (O_1862,N_14947,N_14236);
or UO_1863 (O_1863,N_14735,N_14486);
or UO_1864 (O_1864,N_14896,N_14692);
nor UO_1865 (O_1865,N_14121,N_14807);
or UO_1866 (O_1866,N_14614,N_14807);
and UO_1867 (O_1867,N_14200,N_14754);
nand UO_1868 (O_1868,N_14365,N_14106);
and UO_1869 (O_1869,N_14282,N_14570);
nor UO_1870 (O_1870,N_14317,N_14275);
and UO_1871 (O_1871,N_14885,N_14067);
and UO_1872 (O_1872,N_14771,N_14240);
and UO_1873 (O_1873,N_14184,N_14322);
and UO_1874 (O_1874,N_14544,N_14326);
or UO_1875 (O_1875,N_14607,N_14830);
nand UO_1876 (O_1876,N_14962,N_14567);
or UO_1877 (O_1877,N_14195,N_14737);
and UO_1878 (O_1878,N_14398,N_14983);
or UO_1879 (O_1879,N_14953,N_14091);
and UO_1880 (O_1880,N_14315,N_14220);
xnor UO_1881 (O_1881,N_14668,N_14897);
and UO_1882 (O_1882,N_14932,N_14045);
nand UO_1883 (O_1883,N_14199,N_14167);
and UO_1884 (O_1884,N_14558,N_14398);
xnor UO_1885 (O_1885,N_14452,N_14913);
nand UO_1886 (O_1886,N_14784,N_14206);
nor UO_1887 (O_1887,N_14962,N_14598);
nand UO_1888 (O_1888,N_14991,N_14636);
xor UO_1889 (O_1889,N_14091,N_14232);
and UO_1890 (O_1890,N_14976,N_14119);
nor UO_1891 (O_1891,N_14150,N_14205);
xnor UO_1892 (O_1892,N_14431,N_14484);
nand UO_1893 (O_1893,N_14199,N_14069);
nor UO_1894 (O_1894,N_14160,N_14417);
and UO_1895 (O_1895,N_14345,N_14712);
nand UO_1896 (O_1896,N_14903,N_14482);
nor UO_1897 (O_1897,N_14627,N_14274);
nand UO_1898 (O_1898,N_14262,N_14230);
nor UO_1899 (O_1899,N_14337,N_14435);
xnor UO_1900 (O_1900,N_14871,N_14926);
and UO_1901 (O_1901,N_14578,N_14770);
or UO_1902 (O_1902,N_14556,N_14980);
or UO_1903 (O_1903,N_14355,N_14509);
xor UO_1904 (O_1904,N_14721,N_14466);
or UO_1905 (O_1905,N_14274,N_14061);
nand UO_1906 (O_1906,N_14728,N_14823);
or UO_1907 (O_1907,N_14201,N_14679);
or UO_1908 (O_1908,N_14228,N_14529);
nand UO_1909 (O_1909,N_14530,N_14832);
nand UO_1910 (O_1910,N_14855,N_14156);
nand UO_1911 (O_1911,N_14905,N_14586);
and UO_1912 (O_1912,N_14100,N_14699);
xor UO_1913 (O_1913,N_14368,N_14376);
or UO_1914 (O_1914,N_14025,N_14328);
nand UO_1915 (O_1915,N_14270,N_14617);
nand UO_1916 (O_1916,N_14006,N_14554);
nor UO_1917 (O_1917,N_14814,N_14539);
nor UO_1918 (O_1918,N_14284,N_14282);
nor UO_1919 (O_1919,N_14252,N_14369);
and UO_1920 (O_1920,N_14555,N_14324);
or UO_1921 (O_1921,N_14138,N_14086);
or UO_1922 (O_1922,N_14969,N_14515);
xnor UO_1923 (O_1923,N_14907,N_14316);
or UO_1924 (O_1924,N_14561,N_14999);
and UO_1925 (O_1925,N_14178,N_14315);
or UO_1926 (O_1926,N_14191,N_14167);
or UO_1927 (O_1927,N_14733,N_14786);
and UO_1928 (O_1928,N_14556,N_14305);
nand UO_1929 (O_1929,N_14049,N_14105);
nor UO_1930 (O_1930,N_14941,N_14940);
and UO_1931 (O_1931,N_14431,N_14938);
and UO_1932 (O_1932,N_14020,N_14246);
nand UO_1933 (O_1933,N_14696,N_14711);
or UO_1934 (O_1934,N_14453,N_14814);
nand UO_1935 (O_1935,N_14128,N_14781);
nor UO_1936 (O_1936,N_14184,N_14361);
and UO_1937 (O_1937,N_14769,N_14485);
xor UO_1938 (O_1938,N_14788,N_14211);
nor UO_1939 (O_1939,N_14428,N_14540);
xnor UO_1940 (O_1940,N_14511,N_14489);
xnor UO_1941 (O_1941,N_14093,N_14922);
nor UO_1942 (O_1942,N_14520,N_14409);
nand UO_1943 (O_1943,N_14833,N_14980);
nand UO_1944 (O_1944,N_14865,N_14547);
or UO_1945 (O_1945,N_14338,N_14947);
xor UO_1946 (O_1946,N_14679,N_14005);
nand UO_1947 (O_1947,N_14439,N_14100);
nand UO_1948 (O_1948,N_14073,N_14833);
nor UO_1949 (O_1949,N_14348,N_14088);
nand UO_1950 (O_1950,N_14073,N_14793);
or UO_1951 (O_1951,N_14889,N_14954);
xor UO_1952 (O_1952,N_14969,N_14399);
or UO_1953 (O_1953,N_14321,N_14921);
and UO_1954 (O_1954,N_14495,N_14356);
nor UO_1955 (O_1955,N_14057,N_14582);
nor UO_1956 (O_1956,N_14628,N_14336);
nor UO_1957 (O_1957,N_14418,N_14535);
xor UO_1958 (O_1958,N_14397,N_14196);
or UO_1959 (O_1959,N_14946,N_14617);
and UO_1960 (O_1960,N_14030,N_14232);
nor UO_1961 (O_1961,N_14443,N_14642);
nand UO_1962 (O_1962,N_14354,N_14054);
and UO_1963 (O_1963,N_14508,N_14713);
nand UO_1964 (O_1964,N_14267,N_14210);
nor UO_1965 (O_1965,N_14426,N_14627);
and UO_1966 (O_1966,N_14787,N_14652);
and UO_1967 (O_1967,N_14295,N_14692);
xor UO_1968 (O_1968,N_14453,N_14663);
and UO_1969 (O_1969,N_14457,N_14779);
or UO_1970 (O_1970,N_14709,N_14002);
and UO_1971 (O_1971,N_14887,N_14877);
and UO_1972 (O_1972,N_14075,N_14375);
nor UO_1973 (O_1973,N_14936,N_14336);
and UO_1974 (O_1974,N_14366,N_14405);
or UO_1975 (O_1975,N_14423,N_14849);
xnor UO_1976 (O_1976,N_14451,N_14230);
nor UO_1977 (O_1977,N_14715,N_14979);
and UO_1978 (O_1978,N_14933,N_14883);
xor UO_1979 (O_1979,N_14177,N_14390);
nor UO_1980 (O_1980,N_14162,N_14172);
and UO_1981 (O_1981,N_14388,N_14532);
or UO_1982 (O_1982,N_14335,N_14559);
nand UO_1983 (O_1983,N_14399,N_14919);
nor UO_1984 (O_1984,N_14985,N_14681);
nor UO_1985 (O_1985,N_14229,N_14539);
or UO_1986 (O_1986,N_14367,N_14710);
or UO_1987 (O_1987,N_14841,N_14240);
nand UO_1988 (O_1988,N_14308,N_14630);
nand UO_1989 (O_1989,N_14973,N_14403);
nor UO_1990 (O_1990,N_14878,N_14863);
nand UO_1991 (O_1991,N_14558,N_14834);
and UO_1992 (O_1992,N_14614,N_14353);
nand UO_1993 (O_1993,N_14359,N_14897);
and UO_1994 (O_1994,N_14859,N_14568);
nand UO_1995 (O_1995,N_14096,N_14169);
nand UO_1996 (O_1996,N_14276,N_14691);
and UO_1997 (O_1997,N_14990,N_14646);
nand UO_1998 (O_1998,N_14561,N_14778);
or UO_1999 (O_1999,N_14153,N_14291);
endmodule