module basic_2500_25000_3000_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_2108,In_295);
xnor U1 (N_1,In_1945,In_428);
and U2 (N_2,In_4,In_1442);
or U3 (N_3,In_1234,In_583);
and U4 (N_4,In_685,In_780);
and U5 (N_5,In_970,In_1158);
nor U6 (N_6,In_1178,In_807);
xor U7 (N_7,In_2481,In_547);
nand U8 (N_8,In_610,In_1530);
nor U9 (N_9,In_515,In_2176);
and U10 (N_10,In_2412,In_200);
xor U11 (N_11,In_1220,In_108);
nor U12 (N_12,In_765,In_803);
and U13 (N_13,In_837,In_2456);
nand U14 (N_14,In_2064,In_1705);
xnor U15 (N_15,In_170,In_60);
nand U16 (N_16,In_865,In_142);
xor U17 (N_17,In_1842,In_1672);
xnor U18 (N_18,In_1685,In_2076);
or U19 (N_19,In_898,In_1908);
nand U20 (N_20,In_644,In_1302);
nor U21 (N_21,In_2220,In_221);
or U22 (N_22,In_975,In_3);
nand U23 (N_23,In_946,In_1494);
xor U24 (N_24,In_116,In_914);
or U25 (N_25,In_825,In_399);
nand U26 (N_26,In_1077,In_431);
nor U27 (N_27,In_1728,In_408);
nor U28 (N_28,In_1098,In_2249);
and U29 (N_29,In_944,In_796);
xnor U30 (N_30,In_378,In_2016);
xor U31 (N_31,In_1104,In_709);
or U32 (N_32,In_1512,In_1833);
nor U33 (N_33,In_1412,In_467);
xor U34 (N_34,In_852,In_2235);
nor U35 (N_35,In_2202,In_1271);
and U36 (N_36,In_527,In_1827);
and U37 (N_37,In_380,In_5);
nand U38 (N_38,In_2476,In_1191);
or U39 (N_39,In_1469,In_1625);
xnor U40 (N_40,In_1974,In_647);
and U41 (N_41,In_419,In_1056);
nand U42 (N_42,In_1181,In_146);
nand U43 (N_43,In_1041,In_614);
nand U44 (N_44,In_1004,In_371);
and U45 (N_45,In_1830,In_294);
and U46 (N_46,In_630,In_1207);
and U47 (N_47,In_654,In_1358);
or U48 (N_48,In_443,In_293);
and U49 (N_49,In_902,In_1978);
xnor U50 (N_50,In_2029,In_45);
nor U51 (N_51,In_954,In_1863);
nand U52 (N_52,In_2082,In_2281);
xnor U53 (N_53,In_2437,In_262);
nand U54 (N_54,In_1367,In_2393);
nand U55 (N_55,In_1722,In_469);
or U56 (N_56,In_2363,In_1179);
nor U57 (N_57,In_1228,In_2037);
and U58 (N_58,In_696,In_2439);
nor U59 (N_59,In_1920,In_1541);
and U60 (N_60,In_1421,In_171);
xor U61 (N_61,In_1548,In_779);
nand U62 (N_62,In_2424,In_957);
nor U63 (N_63,In_1912,In_2332);
nand U64 (N_64,In_772,In_396);
nand U65 (N_65,In_115,In_1951);
nand U66 (N_66,In_2465,In_1617);
and U67 (N_67,In_2318,In_543);
and U68 (N_68,In_912,In_1235);
nor U69 (N_69,In_1509,In_1006);
xor U70 (N_70,In_690,In_1484);
nor U71 (N_71,In_1382,In_1594);
nor U72 (N_72,In_1648,In_474);
and U73 (N_73,In_2356,In_776);
nand U74 (N_74,In_2100,In_480);
nor U75 (N_75,In_149,In_287);
or U76 (N_76,In_1458,In_1330);
nor U77 (N_77,In_175,In_1420);
nand U78 (N_78,In_205,In_1200);
or U79 (N_79,In_2373,In_129);
or U80 (N_80,In_1433,In_1918);
and U81 (N_81,In_1331,In_2197);
xor U82 (N_82,In_593,In_1873);
or U83 (N_83,In_44,In_1516);
xor U84 (N_84,In_305,In_2366);
and U85 (N_85,In_26,In_2451);
or U86 (N_86,In_1835,In_1649);
or U87 (N_87,In_896,In_7);
xnor U88 (N_88,In_1667,In_2312);
or U89 (N_89,In_227,In_2168);
xor U90 (N_90,In_1927,In_49);
nand U91 (N_91,In_2189,In_1535);
nand U92 (N_92,In_665,In_587);
or U93 (N_93,In_2063,In_1904);
or U94 (N_94,In_877,In_1301);
and U95 (N_95,In_465,In_1069);
xor U96 (N_96,In_1139,In_2129);
xor U97 (N_97,In_851,In_854);
xor U98 (N_98,In_1946,In_1965);
and U99 (N_99,In_281,In_2389);
nor U100 (N_100,In_76,In_471);
nor U101 (N_101,In_525,In_2116);
nand U102 (N_102,In_1710,In_2205);
and U103 (N_103,In_695,In_1928);
or U104 (N_104,In_284,In_1989);
xor U105 (N_105,In_1320,In_1487);
nor U106 (N_106,In_198,In_2104);
xnor U107 (N_107,In_2313,In_2039);
and U108 (N_108,In_787,In_359);
xnor U109 (N_109,In_158,In_345);
nand U110 (N_110,In_2369,In_922);
xor U111 (N_111,In_123,In_2409);
nor U112 (N_112,In_2232,In_1346);
nand U113 (N_113,In_212,In_415);
xnor U114 (N_114,In_1733,In_2198);
nor U115 (N_115,In_135,In_1399);
xnor U116 (N_116,In_2098,In_669);
or U117 (N_117,In_1604,In_1773);
xor U118 (N_118,In_1226,In_1144);
nor U119 (N_119,In_2478,In_566);
or U120 (N_120,In_1278,In_1100);
and U121 (N_121,In_1520,In_2419);
and U122 (N_122,In_707,In_2335);
and U123 (N_123,In_866,In_1919);
xor U124 (N_124,In_22,In_1527);
nor U125 (N_125,In_1824,In_417);
or U126 (N_126,In_1299,In_252);
and U127 (N_127,In_2338,In_475);
xor U128 (N_128,In_2275,In_1394);
or U129 (N_129,In_895,In_762);
or U130 (N_130,In_2190,In_1641);
nor U131 (N_131,In_1291,In_2117);
nor U132 (N_132,In_2449,In_2483);
nand U133 (N_133,In_804,In_521);
xnor U134 (N_134,In_260,In_1470);
or U135 (N_135,In_1380,In_2009);
and U136 (N_136,In_801,In_1603);
or U137 (N_137,In_853,In_1001);
and U138 (N_138,In_1342,In_2336);
or U139 (N_139,In_245,In_1038);
nor U140 (N_140,In_2239,In_2223);
xor U141 (N_141,In_1184,In_65);
nand U142 (N_142,In_847,In_1467);
or U143 (N_143,In_760,In_829);
and U144 (N_144,In_435,In_1032);
xnor U145 (N_145,In_2413,In_2096);
nor U146 (N_146,In_2459,In_2150);
nand U147 (N_147,In_487,In_328);
and U148 (N_148,In_1955,In_1730);
or U149 (N_149,In_2055,In_160);
nand U150 (N_150,In_588,In_1998);
xor U151 (N_151,In_1498,In_1085);
xor U152 (N_152,In_2301,In_98);
and U153 (N_153,In_1752,In_1504);
and U154 (N_154,In_2420,In_908);
and U155 (N_155,In_483,In_1122);
and U156 (N_156,In_1531,In_2148);
xor U157 (N_157,In_11,In_447);
nand U158 (N_158,In_1258,In_256);
nand U159 (N_159,In_210,In_2159);
nand U160 (N_160,In_1057,In_826);
or U161 (N_161,In_697,In_1473);
nor U162 (N_162,In_2273,In_2217);
nand U163 (N_163,In_927,In_1429);
nor U164 (N_164,In_1087,In_2472);
or U165 (N_165,In_1961,In_2475);
and U166 (N_166,In_1883,In_699);
and U167 (N_167,In_1761,In_657);
and U168 (N_168,In_1969,In_661);
or U169 (N_169,In_140,In_463);
and U170 (N_170,In_2090,In_1642);
xnor U171 (N_171,In_503,In_1763);
xor U172 (N_172,In_2042,In_455);
nand U173 (N_173,In_1990,In_157);
and U174 (N_174,In_77,In_1236);
nor U175 (N_175,In_1223,In_1203);
and U176 (N_176,In_2374,In_53);
nor U177 (N_177,In_2361,In_74);
nor U178 (N_178,In_1187,In_1999);
xor U179 (N_179,In_2262,In_1225);
nand U180 (N_180,In_304,In_2357);
nand U181 (N_181,In_64,In_1408);
nand U182 (N_182,In_2378,In_1160);
and U183 (N_183,In_1556,In_2382);
or U184 (N_184,In_1062,In_290);
and U185 (N_185,In_353,In_504);
nor U186 (N_186,In_1340,In_978);
nand U187 (N_187,In_1680,In_127);
or U188 (N_188,In_1798,In_1443);
and U189 (N_189,In_1885,In_692);
and U190 (N_190,In_917,In_1149);
xor U191 (N_191,In_1022,In_2006);
nor U192 (N_192,In_2349,In_2028);
nand U193 (N_193,In_1310,In_1852);
xor U194 (N_194,In_2395,In_189);
or U195 (N_195,In_546,In_143);
nand U196 (N_196,In_2422,In_237);
nand U197 (N_197,In_1933,In_1159);
and U198 (N_198,In_731,In_524);
nand U199 (N_199,In_1309,In_1546);
xnor U200 (N_200,In_403,In_235);
or U201 (N_201,In_2041,In_892);
and U202 (N_202,In_381,In_1640);
nand U203 (N_203,In_2071,In_213);
and U204 (N_204,In_1699,In_1661);
and U205 (N_205,In_2225,In_1284);
nand U206 (N_206,In_2048,In_1524);
xnor U207 (N_207,In_1703,In_2464);
or U208 (N_208,In_1192,In_509);
or U209 (N_209,In_2206,In_2125);
xor U210 (N_210,In_169,In_1567);
nand U211 (N_211,In_664,In_1084);
or U212 (N_212,In_1717,In_1956);
xor U213 (N_213,In_956,In_174);
nand U214 (N_214,In_1911,In_1652);
xor U215 (N_215,In_1706,In_1485);
nand U216 (N_216,In_1026,In_2490);
nor U217 (N_217,In_1079,In_202);
nor U218 (N_218,In_1736,In_2498);
and U219 (N_219,In_2046,In_651);
and U220 (N_220,In_105,In_686);
or U221 (N_221,In_869,In_1479);
xor U222 (N_222,In_1583,In_1448);
nor U223 (N_223,In_1683,In_1256);
nor U224 (N_224,In_1314,In_6);
nor U225 (N_225,In_1459,In_1799);
and U226 (N_226,In_832,In_1180);
xnor U227 (N_227,In_1324,In_1749);
nor U228 (N_228,In_1046,In_1003);
and U229 (N_229,In_58,In_2107);
xnor U230 (N_230,In_163,In_1629);
nand U231 (N_231,In_1950,In_1000);
or U232 (N_232,In_1844,In_1150);
or U233 (N_233,In_2011,In_633);
nor U234 (N_234,In_735,In_1905);
nand U235 (N_235,In_632,In_747);
and U236 (N_236,In_2103,In_59);
nor U237 (N_237,In_891,In_2201);
nand U238 (N_238,In_1177,In_671);
xor U239 (N_239,In_313,In_1211);
xor U240 (N_240,In_715,In_1468);
nand U241 (N_241,In_2179,In_1080);
and U242 (N_242,In_2400,In_1886);
or U243 (N_243,In_589,In_2178);
nor U244 (N_244,In_1311,In_1014);
xor U245 (N_245,In_1671,In_18);
xor U246 (N_246,In_1409,In_1522);
and U247 (N_247,In_2147,In_1186);
and U248 (N_248,In_1106,In_529);
nand U249 (N_249,In_1901,In_2371);
nor U250 (N_250,In_2185,In_337);
or U251 (N_251,In_1845,In_1916);
and U252 (N_252,In_377,In_2362);
or U253 (N_253,In_1690,In_2341);
nor U254 (N_254,In_1765,In_1850);
nor U255 (N_255,In_1917,In_1797);
and U256 (N_256,In_862,In_1692);
xnor U257 (N_257,In_1633,In_1616);
and U258 (N_258,In_1049,In_1726);
xor U259 (N_259,In_1746,In_2200);
nor U260 (N_260,In_1925,In_1086);
or U261 (N_261,In_2061,In_910);
nor U262 (N_262,In_2416,In_823);
xor U263 (N_263,In_2181,In_2334);
nor U264 (N_264,In_1313,In_254);
and U265 (N_265,In_783,In_2146);
nand U266 (N_266,In_191,In_288);
and U267 (N_267,In_2385,In_830);
nor U268 (N_268,In_950,In_512);
or U269 (N_269,In_439,In_2345);
nand U270 (N_270,In_424,In_1294);
or U271 (N_271,In_1823,In_656);
xor U272 (N_272,In_476,In_725);
xnor U273 (N_273,In_2145,In_2322);
nor U274 (N_274,In_1668,In_613);
and U275 (N_275,In_239,In_1374);
xor U276 (N_276,In_1591,In_2126);
nand U277 (N_277,In_1618,In_2492);
nor U278 (N_278,In_2019,In_1357);
nor U279 (N_279,In_742,In_2152);
nor U280 (N_280,In_1689,In_1146);
nand U281 (N_281,In_2018,In_2443);
or U282 (N_282,In_1489,In_1027);
and U283 (N_283,In_980,In_343);
xnor U284 (N_284,In_2056,In_279);
and U285 (N_285,In_429,In_2445);
xor U286 (N_286,In_1768,In_995);
xor U287 (N_287,In_813,In_1913);
and U288 (N_288,In_1859,In_1549);
nand U289 (N_289,In_1876,In_2162);
nor U290 (N_290,In_2268,In_615);
xnor U291 (N_291,In_1624,In_993);
nor U292 (N_292,In_183,In_984);
nand U293 (N_293,In_1052,In_1204);
nor U294 (N_294,In_727,In_704);
or U295 (N_295,In_1949,In_56);
and U296 (N_296,In_440,In_1719);
or U297 (N_297,In_1126,In_50);
nor U298 (N_298,In_2236,In_38);
nand U299 (N_299,In_1663,In_2105);
or U300 (N_300,In_1188,In_25);
xnor U301 (N_301,In_426,In_582);
and U302 (N_302,In_2058,In_1893);
or U303 (N_303,In_1317,In_2226);
nor U304 (N_304,In_700,In_2234);
and U305 (N_305,In_1152,In_1569);
and U306 (N_306,In_296,In_1995);
or U307 (N_307,In_2031,In_2370);
or U308 (N_308,In_1804,In_687);
or U309 (N_309,In_2122,In_868);
or U310 (N_310,In_448,In_2032);
nor U311 (N_311,In_1450,In_596);
and U312 (N_312,In_1163,In_1816);
nor U313 (N_313,In_1643,In_2277);
or U314 (N_314,In_1721,In_2325);
and U315 (N_315,In_1560,In_2184);
or U316 (N_316,In_13,In_969);
or U317 (N_317,In_2073,In_1);
nor U318 (N_318,In_1197,In_433);
nand U319 (N_319,In_2388,In_1350);
nand U320 (N_320,In_2279,In_99);
or U321 (N_321,In_121,In_2091);
or U322 (N_322,In_757,In_620);
or U323 (N_323,In_208,In_1981);
nor U324 (N_324,In_277,In_802);
or U325 (N_325,In_2462,In_1557);
and U326 (N_326,In_1767,In_89);
xnor U327 (N_327,In_2045,In_2130);
nor U328 (N_328,In_929,In_2414);
or U329 (N_329,In_1147,In_2066);
and U330 (N_330,In_1500,In_1243);
xor U331 (N_331,In_712,In_93);
xnor U332 (N_332,In_23,In_2311);
or U333 (N_333,In_1345,In_1456);
xnor U334 (N_334,In_1865,In_1738);
nor U335 (N_335,In_1304,In_268);
or U336 (N_336,In_387,In_2120);
or U337 (N_337,In_986,In_1670);
nor U338 (N_338,In_621,In_39);
nor U339 (N_339,In_1053,In_358);
and U340 (N_340,In_31,In_1170);
and U341 (N_341,In_1064,In_2381);
and U342 (N_342,In_1347,In_658);
nor U343 (N_343,In_798,In_2187);
and U344 (N_344,In_2013,In_85);
and U345 (N_345,In_2119,In_368);
nor U346 (N_346,In_113,In_2208);
nand U347 (N_347,In_2421,In_849);
or U348 (N_348,In_1471,In_563);
xor U349 (N_349,In_1411,In_1343);
xor U350 (N_350,In_1877,In_2278);
nor U351 (N_351,In_2106,In_1262);
nand U352 (N_352,In_1169,In_1395);
nand U353 (N_353,In_324,In_1472);
nor U354 (N_354,In_518,In_2078);
or U355 (N_355,In_446,In_2323);
and U356 (N_356,In_159,In_2427);
and U357 (N_357,In_2435,In_261);
or U358 (N_358,In_231,In_739);
or U359 (N_359,In_926,In_2215);
xor U360 (N_360,In_681,In_1483);
xnor U361 (N_361,In_1327,In_1040);
nor U362 (N_362,In_1289,In_2316);
xnor U363 (N_363,In_1227,In_545);
nor U364 (N_364,In_1452,In_166);
nand U365 (N_365,In_920,In_679);
nor U366 (N_366,In_609,In_1402);
xnor U367 (N_367,In_1586,In_1682);
nand U368 (N_368,In_2229,In_1803);
or U369 (N_369,In_1050,In_114);
and U370 (N_370,In_1679,In_1171);
nand U371 (N_371,In_81,In_1849);
xnor U372 (N_372,In_1283,In_1932);
and U373 (N_373,In_398,In_2497);
nor U374 (N_374,In_1577,In_1611);
xnor U375 (N_375,In_1502,In_556);
nor U376 (N_376,In_393,In_740);
xor U377 (N_377,In_182,In_1862);
or U378 (N_378,In_1547,In_1240);
and U379 (N_379,In_1786,In_1599);
xnor U380 (N_380,In_2228,In_473);
and U381 (N_381,In_599,In_2191);
nor U382 (N_382,In_1102,In_834);
nor U383 (N_383,In_1977,In_1476);
nor U384 (N_384,In_250,In_1348);
and U385 (N_385,In_2401,In_1581);
nor U386 (N_386,In_1646,In_1691);
xnor U387 (N_387,In_126,In_1488);
or U388 (N_388,In_133,In_622);
nand U389 (N_389,In_557,In_2326);
xor U390 (N_390,In_989,In_2469);
and U391 (N_391,In_2077,In_360);
and U392 (N_392,In_331,In_1011);
or U393 (N_393,In_1954,In_2167);
xor U394 (N_394,In_2070,In_1012);
nand U395 (N_395,In_96,In_312);
and U396 (N_396,In_531,In_522);
or U397 (N_397,In_2180,In_1597);
and U398 (N_398,In_1229,In_1116);
and U399 (N_399,In_382,In_238);
or U400 (N_400,In_228,In_966);
nor U401 (N_401,In_1248,In_502);
nor U402 (N_402,In_1678,In_676);
xor U403 (N_403,In_1941,In_222);
nor U404 (N_404,In_2259,In_413);
and U405 (N_405,In_310,In_323);
and U406 (N_406,In_62,In_1462);
xor U407 (N_407,In_2118,In_2230);
and U408 (N_408,In_80,In_1495);
xnor U409 (N_409,In_1819,In_1215);
xor U410 (N_410,In_2330,In_1501);
nand U411 (N_411,In_1906,In_913);
xor U412 (N_412,In_1434,In_1492);
xor U413 (N_413,In_1461,In_2059);
nor U414 (N_414,In_844,In_840);
xnor U415 (N_415,In_741,In_156);
nor U416 (N_416,In_909,In_842);
nand U417 (N_417,In_960,In_2491);
xnor U418 (N_418,In_462,In_1743);
nand U419 (N_419,In_2034,In_790);
nor U420 (N_420,In_2315,In_2247);
xnor U421 (N_421,In_1426,In_2350);
or U422 (N_422,In_1005,In_2319);
and U423 (N_423,In_190,In_384);
nand U424 (N_424,In_1953,In_1938);
xor U425 (N_425,In_1851,In_893);
nand U426 (N_426,In_164,In_1265);
xor U427 (N_427,In_1994,In_220);
nand U428 (N_428,In_333,In_2170);
xor U429 (N_429,In_2132,In_619);
nor U430 (N_430,In_544,In_778);
or U431 (N_431,In_449,In_247);
nand U432 (N_432,In_1435,In_500);
nor U433 (N_433,In_2367,In_362);
or U434 (N_434,In_2254,In_2068);
nor U435 (N_435,In_2177,In_1963);
or U436 (N_436,In_63,In_918);
xor U437 (N_437,In_265,In_1114);
nor U438 (N_438,In_1282,In_214);
nand U439 (N_439,In_1323,In_95);
xnor U440 (N_440,In_1054,In_520);
nor U441 (N_441,In_488,In_2347);
or U442 (N_442,In_1529,In_1131);
or U443 (N_443,In_1300,In_263);
nand U444 (N_444,In_653,In_2460);
xnor U445 (N_445,In_1538,In_885);
nand U446 (N_446,In_1151,In_2231);
nor U447 (N_447,In_477,In_1909);
nor U448 (N_448,In_977,In_1045);
and U449 (N_449,In_1758,In_339);
and U450 (N_450,In_1112,In_625);
nand U451 (N_451,In_1727,In_873);
nand U452 (N_452,In_1021,In_2099);
or U453 (N_453,In_703,In_623);
or U454 (N_454,In_150,In_2305);
nor U455 (N_455,In_2255,In_2284);
nor U456 (N_456,In_1337,In_781);
and U457 (N_457,In_363,In_627);
or U458 (N_458,In_2065,In_109);
xor U459 (N_459,In_1811,In_1944);
or U460 (N_460,In_1148,In_1189);
nand U461 (N_461,In_1238,In_643);
nor U462 (N_462,In_1587,In_2408);
or U463 (N_463,In_1800,In_2165);
nand U464 (N_464,In_1864,In_1414);
nor U465 (N_465,In_1066,In_508);
nand U466 (N_466,In_2218,In_1219);
and U467 (N_467,In_1601,In_1821);
xor U468 (N_468,In_955,In_1540);
nand U469 (N_469,In_2199,In_894);
or U470 (N_470,In_1894,In_1725);
or U471 (N_471,In_364,In_2440);
and U472 (N_472,In_1401,In_2292);
and U473 (N_473,In_901,In_1390);
and U474 (N_474,In_2372,In_843);
xor U475 (N_475,In_1630,In_370);
nor U476 (N_476,In_600,In_594);
xor U477 (N_477,In_1936,In_2141);
nand U478 (N_478,In_2377,In_2487);
or U479 (N_479,In_1335,In_732);
or U480 (N_480,In_1428,In_1874);
nor U481 (N_481,In_2471,In_2423);
nor U482 (N_482,In_1183,In_234);
nor U483 (N_483,In_1687,In_201);
or U484 (N_484,In_822,In_994);
xor U485 (N_485,In_1083,In_870);
nor U486 (N_486,In_973,In_819);
and U487 (N_487,In_1868,In_29);
xor U488 (N_488,In_267,In_236);
nand U489 (N_489,In_1326,In_729);
nor U490 (N_490,In_2390,In_2457);
or U491 (N_491,In_1206,In_2030);
nand U492 (N_492,In_1355,In_1552);
or U493 (N_493,In_327,In_2174);
or U494 (N_494,In_875,In_280);
xnor U495 (N_495,In_481,In_1771);
nand U496 (N_496,In_1718,In_253);
nor U497 (N_497,In_1028,In_558);
xnor U498 (N_498,In_1364,In_1043);
and U499 (N_499,In_888,In_2441);
nand U500 (N_500,In_2317,In_1782);
nor U501 (N_501,N_430,N_38);
and U502 (N_502,In_1855,In_356);
and U503 (N_503,In_232,In_376);
or U504 (N_504,N_349,In_180);
nand U505 (N_505,N_132,In_12);
and U506 (N_506,In_925,N_64);
nor U507 (N_507,In_2410,In_492);
nand U508 (N_508,In_666,In_2488);
or U509 (N_509,In_111,In_2436);
or U510 (N_510,In_2482,In_292);
and U511 (N_511,In_32,In_1880);
and U512 (N_512,In_1713,In_2036);
or U513 (N_513,In_1195,In_1055);
or U514 (N_514,In_464,In_325);
xor U515 (N_515,In_1332,In_2138);
or U516 (N_516,In_2425,In_2328);
xnor U517 (N_517,N_150,In_1034);
and U518 (N_518,In_2113,N_499);
nand U519 (N_519,In_1871,N_42);
nor U520 (N_520,In_650,In_1973);
xor U521 (N_521,In_395,N_37);
xnor U522 (N_522,In_1554,In_43);
nand U523 (N_523,In_595,In_2387);
nor U524 (N_524,In_736,In_422);
or U525 (N_525,In_1542,In_1677);
nor U526 (N_526,N_121,In_2020);
and U527 (N_527,In_2265,In_1292);
or U528 (N_528,In_2392,In_2084);
nor U529 (N_529,In_660,N_229);
xnor U530 (N_530,In_1250,In_72);
or U531 (N_531,In_1360,In_517);
nor U532 (N_532,In_981,In_2222);
or U533 (N_533,In_1349,N_290);
xor U534 (N_534,N_367,In_514);
nand U535 (N_535,N_66,In_86);
and U536 (N_536,N_376,In_1937);
or U537 (N_537,In_900,In_1942);
and U538 (N_538,N_346,In_1628);
and U539 (N_539,N_2,In_996);
nor U540 (N_540,N_396,N_300);
nand U541 (N_541,In_2384,In_1482);
xor U542 (N_542,In_2297,N_352);
xor U543 (N_543,In_2430,In_1334);
and U544 (N_544,In_693,N_303);
nand U545 (N_545,In_1993,N_149);
or U546 (N_546,In_106,In_1297);
nor U547 (N_547,In_352,In_2308);
nor U548 (N_548,In_911,In_1121);
nor U549 (N_549,In_1082,N_464);
or U550 (N_550,In_1627,N_250);
and U551 (N_551,In_315,In_1070);
or U552 (N_552,N_240,In_1344);
nor U553 (N_553,N_14,In_1029);
and U554 (N_554,N_392,In_711);
nor U555 (N_555,In_1232,In_2344);
xor U556 (N_556,In_1729,In_2196);
nand U557 (N_557,N_408,In_1605);
nand U558 (N_558,In_2479,In_300);
nand U559 (N_559,N_412,In_1766);
xor U560 (N_560,In_2022,In_2288);
xor U561 (N_561,In_173,In_329);
and U562 (N_562,In_1035,In_857);
nor U563 (N_563,In_2486,In_678);
xor U564 (N_564,N_432,In_1276);
nor U565 (N_565,N_404,N_36);
xnor U566 (N_566,In_2299,In_1373);
or U567 (N_567,In_2203,In_2133);
nor U568 (N_568,In_2343,In_1902);
nand U569 (N_569,N_124,N_11);
nand U570 (N_570,In_1796,In_2067);
nor U571 (N_571,In_698,In_1202);
or U572 (N_572,In_73,In_733);
and U573 (N_573,In_1198,In_1665);
and U574 (N_574,In_1510,In_1580);
nand U575 (N_575,In_1315,In_921);
xor U576 (N_576,In_1205,N_466);
xnor U577 (N_577,In_774,In_1793);
or U578 (N_578,N_163,In_494);
nand U579 (N_579,In_2248,In_1059);
nor U580 (N_580,In_308,In_2428);
nor U581 (N_581,In_874,In_1002);
and U582 (N_582,In_1818,N_217);
nand U583 (N_583,In_1762,In_340);
nor U584 (N_584,In_344,In_988);
and U585 (N_585,In_2327,In_2450);
xor U586 (N_586,N_147,In_1631);
xnor U587 (N_587,In_1734,N_288);
and U588 (N_588,In_1105,In_391);
xnor U589 (N_589,In_2000,In_1715);
or U590 (N_590,In_1785,In_1269);
or U591 (N_591,In_705,In_2153);
xnor U592 (N_592,In_412,In_668);
and U593 (N_593,In_203,In_562);
or U594 (N_594,N_273,N_277);
nor U595 (N_595,In_354,In_427);
nand U596 (N_596,In_987,N_207);
xnor U597 (N_597,In_905,In_2015);
xnor U598 (N_598,In_1825,In_217);
xor U599 (N_599,In_320,In_601);
or U600 (N_600,In_1295,In_225);
nor U601 (N_601,In_1707,N_206);
nor U602 (N_602,In_1988,In_629);
nor U603 (N_603,In_876,In_1562);
nor U604 (N_604,In_1201,In_1389);
nand U605 (N_605,In_1274,In_1199);
or U606 (N_606,N_71,N_84);
nor U607 (N_607,In_1720,N_443);
xnor U608 (N_608,In_964,In_1268);
nor U609 (N_609,In_916,N_281);
and U610 (N_610,In_2368,In_1422);
or U611 (N_611,In_75,In_2014);
or U612 (N_612,In_1111,In_2227);
or U613 (N_613,In_2245,N_323);
xnor U614 (N_614,In_88,In_1848);
and U615 (N_615,In_2142,In_2287);
xor U616 (N_616,N_63,In_789);
or U617 (N_617,N_427,In_1709);
nor U618 (N_618,In_507,In_357);
xnor U619 (N_619,In_949,In_1024);
or U620 (N_620,In_1675,In_1417);
and U621 (N_621,N_265,In_341);
nand U622 (N_622,N_454,In_2195);
nand U623 (N_623,In_1579,In_16);
nor U624 (N_624,In_2035,In_2359);
nand U625 (N_625,In_937,In_734);
or U626 (N_626,In_338,In_1506);
nand U627 (N_627,In_2467,In_677);
or U628 (N_628,N_377,In_1593);
and U629 (N_629,In_197,N_347);
nand U630 (N_630,N_119,N_48);
and U631 (N_631,In_1384,N_449);
nor U632 (N_632,In_1213,N_284);
xnor U633 (N_633,N_162,In_450);
nor U634 (N_634,In_1133,N_228);
nor U635 (N_635,In_1656,N_4);
nand U636 (N_636,In_1834,In_1051);
xor U637 (N_637,N_212,In_1097);
nand U638 (N_638,In_1783,In_1645);
xnor U639 (N_639,In_172,N_258);
and U640 (N_640,N_424,In_634);
and U641 (N_641,In_84,In_516);
or U642 (N_642,In_472,In_569);
xnor U643 (N_643,In_1020,In_2240);
nor U644 (N_644,In_348,In_680);
and U645 (N_645,In_1257,N_494);
and U646 (N_646,In_2353,In_2480);
or U647 (N_647,N_157,N_190);
nand U648 (N_648,In_147,In_2060);
nand U649 (N_649,In_999,In_1044);
nor U650 (N_650,N_21,N_421);
or U651 (N_651,N_272,In_2038);
nor U652 (N_652,In_2139,In_638);
or U653 (N_653,N_282,In_1806);
xor U654 (N_654,In_1638,In_1288);
xor U655 (N_655,N_123,In_141);
xnor U656 (N_656,In_537,In_94);
xnor U657 (N_657,In_2194,In_773);
and U658 (N_658,N_101,In_1947);
nand U659 (N_659,In_1514,In_886);
xnor U660 (N_660,N_165,In_1067);
or U661 (N_661,In_2360,In_1175);
nand U662 (N_662,N_231,N_302);
nor U663 (N_663,In_1030,N_364);
and U664 (N_664,N_24,In_1636);
nor U665 (N_665,In_952,N_468);
or U666 (N_666,N_374,In_1737);
nor U667 (N_667,N_293,In_1157);
nor U668 (N_668,In_1481,In_753);
nor U669 (N_669,N_387,N_398);
nand U670 (N_670,In_846,In_2172);
and U671 (N_671,In_1790,In_2112);
xor U672 (N_672,In_1437,In_2340);
nand U673 (N_673,In_967,In_549);
nand U674 (N_674,In_365,N_481);
xnor U675 (N_675,In_1634,In_1971);
and U676 (N_676,In_1425,In_758);
nor U677 (N_677,In_2442,N_200);
or U678 (N_678,In_2092,N_27);
or U679 (N_679,N_373,In_1867);
nand U680 (N_680,In_1696,In_744);
or U681 (N_681,N_275,In_1789);
xnor U682 (N_682,In_1209,N_345);
or U683 (N_683,N_260,In_1772);
or U684 (N_684,In_1351,N_113);
and U685 (N_685,In_584,N_471);
nor U686 (N_686,In_97,N_16);
and U687 (N_687,N_498,In_1430);
or U688 (N_688,In_2094,In_1585);
xor U689 (N_689,In_185,In_2256);
nand U690 (N_690,N_313,In_1418);
or U691 (N_691,N_356,N_423);
xnor U692 (N_692,In_720,In_1780);
nor U693 (N_693,In_456,N_314);
or U694 (N_694,N_386,In_764);
nor U695 (N_695,In_1129,N_67);
or U696 (N_696,In_1217,In_1466);
xor U697 (N_697,N_270,In_592);
or U698 (N_698,In_880,In_240);
and U699 (N_699,N_224,In_1493);
xnor U700 (N_700,In_1025,In_1312);
xor U701 (N_701,In_1644,In_1153);
or U702 (N_702,In_66,N_378);
nand U703 (N_703,In_1457,N_419);
or U704 (N_704,N_246,In_1352);
or U705 (N_705,In_1463,In_606);
xor U706 (N_706,In_270,N_239);
and U707 (N_707,In_2025,In_940);
nor U708 (N_708,In_906,In_1415);
nor U709 (N_709,N_203,In_2110);
and U710 (N_710,In_799,In_1132);
and U711 (N_711,In_2285,N_400);
nor U712 (N_712,In_1814,In_972);
nand U713 (N_713,In_2383,N_75);
and U714 (N_714,In_1582,In_743);
xor U715 (N_715,N_6,In_1651);
or U716 (N_716,In_1935,In_55);
and U717 (N_717,N_204,In_1120);
nor U718 (N_718,In_723,In_810);
xor U719 (N_719,In_2164,In_1794);
nor U720 (N_720,N_46,In_390);
or U721 (N_721,N_74,In_1009);
nand U722 (N_722,In_2431,In_410);
nand U723 (N_723,In_1805,In_2243);
and U724 (N_724,N_480,N_18);
nand U725 (N_725,In_2274,N_294);
and U726 (N_726,In_1559,In_649);
and U727 (N_727,N_331,N_316);
nand U728 (N_728,In_934,In_809);
nand U729 (N_729,In_691,In_2216);
or U730 (N_730,In_1613,N_197);
or U731 (N_731,In_120,N_333);
nor U732 (N_732,In_1831,In_1503);
and U733 (N_733,In_899,In_1185);
nor U734 (N_734,N_256,In_125);
xnor U735 (N_735,In_2135,In_1403);
and U736 (N_736,N_429,In_1801);
or U737 (N_737,In_285,In_1218);
nand U738 (N_738,N_127,N_366);
nor U739 (N_739,In_1659,In_1673);
or U740 (N_740,In_2396,In_1764);
and U741 (N_741,In_401,In_2171);
nand U742 (N_742,In_598,N_334);
nor U743 (N_743,In_2251,N_436);
nor U744 (N_744,In_1832,In_2175);
nor U745 (N_745,In_1870,In_881);
and U746 (N_746,N_226,In_1103);
xnor U747 (N_747,In_501,In_2499);
nor U748 (N_748,In_2237,In_1396);
nand U749 (N_749,In_2188,In_548);
or U750 (N_750,In_188,N_178);
nor U751 (N_751,N_188,In_1891);
or U752 (N_752,In_1325,In_959);
and U753 (N_753,N_418,In_1976);
and U754 (N_754,In_1230,In_258);
nor U755 (N_755,In_1698,In_2415);
and U756 (N_756,In_1252,N_153);
or U757 (N_757,In_1637,In_2026);
and U758 (N_758,N_122,In_2365);
or U759 (N_759,In_46,N_193);
nand U760 (N_760,In_2418,In_1626);
nand U761 (N_761,In_1809,In_1109);
and U762 (N_762,In_48,N_33);
and U763 (N_763,In_1254,In_769);
and U764 (N_764,N_393,In_1957);
or U765 (N_765,N_286,N_311);
nor U766 (N_766,In_1381,N_96);
nand U767 (N_767,In_561,In_580);
and U768 (N_768,In_1259,In_1376);
xor U769 (N_769,N_493,N_342);
and U770 (N_770,N_26,In_1078);
nor U771 (N_771,In_784,In_1247);
nor U772 (N_772,In_1695,In_1210);
nor U773 (N_773,In_1486,In_2017);
nand U774 (N_774,N_492,In_1118);
and U775 (N_775,N_299,In_564);
nand U776 (N_776,In_2010,In_571);
nor U777 (N_777,In_2270,In_420);
nor U778 (N_778,In_871,In_1899);
nor U779 (N_779,In_418,N_138);
xor U780 (N_780,N_191,In_430);
xor U781 (N_781,In_2339,In_863);
or U782 (N_782,In_118,In_400);
nand U783 (N_783,In_2040,In_1371);
and U784 (N_784,In_1924,N_13);
nand U785 (N_785,In_642,In_1164);
or U786 (N_786,N_221,In_1436);
and U787 (N_787,In_28,In_1194);
nor U788 (N_788,In_2295,In_1943);
nor U789 (N_789,In_1071,In_510);
nand U790 (N_790,In_2298,In_1694);
or U791 (N_791,In_1890,In_289);
and U792 (N_792,In_800,N_431);
xor U793 (N_793,In_2257,In_2002);
or U794 (N_794,In_2386,In_997);
or U795 (N_795,In_194,In_983);
nor U796 (N_796,In_306,In_1856);
xor U797 (N_797,In_374,In_574);
and U798 (N_798,In_538,N_319);
nor U799 (N_799,In_1190,In_1750);
or U800 (N_800,In_461,N_372);
nand U801 (N_801,In_36,In_982);
nor U802 (N_802,N_135,In_2405);
nand U803 (N_803,In_2302,In_662);
and U804 (N_804,In_1033,N_202);
xnor U805 (N_805,In_1101,In_1658);
and U806 (N_806,In_168,In_2069);
nor U807 (N_807,N_199,In_795);
xnor U808 (N_808,In_1321,N_308);
or U809 (N_809,N_496,In_737);
xnor U810 (N_810,N_434,N_335);
or U811 (N_811,In_1964,N_56);
xor U812 (N_812,In_617,In_1817);
xnor U813 (N_813,N_171,N_358);
nor U814 (N_814,In_152,In_2250);
nor U815 (N_815,In_2057,N_459);
nand U816 (N_816,N_369,In_1166);
nor U817 (N_817,In_104,In_565);
or U818 (N_818,In_1654,N_109);
xnor U819 (N_819,N_394,N_60);
nor U820 (N_820,In_1550,In_416);
or U821 (N_821,In_421,In_355);
xor U822 (N_822,In_155,In_533);
nor U823 (N_823,In_570,In_831);
or U824 (N_824,In_248,In_1701);
nand U825 (N_825,In_1915,In_388);
or U826 (N_826,In_385,N_179);
xnor U827 (N_827,In_342,N_415);
and U828 (N_828,In_266,N_365);
or U829 (N_829,In_1124,In_1369);
and U830 (N_830,N_309,In_534);
or U831 (N_831,In_1296,In_1760);
xnor U832 (N_832,In_47,N_88);
and U833 (N_833,N_482,In_451);
nand U834 (N_834,In_1096,In_763);
nand U835 (N_835,In_2209,In_15);
or U836 (N_836,In_1404,In_848);
or U837 (N_837,In_1776,In_1480);
and U838 (N_838,In_785,In_1511);
and U839 (N_839,In_162,In_1031);
and U840 (N_840,N_474,In_317);
nor U841 (N_841,In_2286,In_675);
nor U842 (N_842,In_40,In_1145);
or U843 (N_843,In_2444,In_771);
and U844 (N_844,In_1791,N_106);
or U845 (N_845,In_602,In_560);
xor U846 (N_846,In_2242,In_1273);
nor U847 (N_847,In_2411,In_833);
and U848 (N_848,In_491,N_100);
nand U849 (N_849,In_457,In_264);
or U850 (N_850,In_759,N_159);
or U851 (N_851,In_674,In_1316);
nand U852 (N_852,In_2252,In_2221);
nand U853 (N_853,In_2429,In_714);
and U854 (N_854,In_2062,In_1019);
xor U855 (N_855,N_475,In_1251);
and U856 (N_856,In_943,In_1253);
nor U857 (N_857,In_1839,N_389);
xnor U858 (N_858,In_1881,N_130);
nor U859 (N_859,In_728,N_220);
xor U860 (N_860,In_1431,In_1119);
xnor U861 (N_861,In_68,N_79);
or U862 (N_862,In_1565,In_2127);
nand U863 (N_863,In_1441,In_122);
and U864 (N_864,In_1224,In_1008);
and U865 (N_865,N_420,In_667);
and U866 (N_866,In_1878,In_1449);
and U867 (N_867,In_301,N_255);
and U868 (N_868,In_211,In_1275);
xor U869 (N_869,In_1445,N_336);
and U870 (N_870,In_2086,In_176);
xor U871 (N_871,N_457,N_218);
and U872 (N_872,N_166,N_55);
or U873 (N_873,In_1246,In_192);
or U874 (N_874,In_1307,In_452);
nor U875 (N_875,In_1775,In_523);
nand U876 (N_876,In_2044,N_329);
and U877 (N_877,In_1543,N_289);
nand U878 (N_878,In_856,In_193);
nor U879 (N_879,N_73,In_1154);
nand U880 (N_880,In_1362,In_286);
xnor U881 (N_881,N_370,In_486);
nor U882 (N_882,In_373,In_444);
nand U883 (N_883,N_360,N_237);
nor U884 (N_884,N_355,In_1237);
and U885 (N_885,N_411,In_1934);
xnor U886 (N_886,In_1042,N_136);
nor U887 (N_887,In_1134,In_466);
or U888 (N_888,In_2211,In_470);
nand U889 (N_889,In_827,In_441);
or U890 (N_890,In_1807,In_1702);
or U891 (N_891,N_350,In_69);
nand U892 (N_892,In_724,In_423);
nor U893 (N_893,In_1372,N_144);
xor U894 (N_894,N_187,In_1387);
xnor U895 (N_895,In_2154,In_495);
or U896 (N_896,N_92,In_948);
xor U897 (N_897,In_297,In_1093);
or U898 (N_898,In_17,In_1176);
nand U899 (N_899,In_1829,In_1013);
or U900 (N_900,In_867,In_639);
xor U901 (N_901,N_458,In_1711);
and U902 (N_902,In_1576,In_748);
nand U903 (N_903,In_1967,In_710);
nand U904 (N_904,In_92,In_786);
xor U905 (N_905,N_315,N_340);
nand U906 (N_906,In_1474,N_437);
or U907 (N_907,In_1465,In_1322);
or U908 (N_908,In_1091,In_752);
and U909 (N_909,In_536,In_719);
and U910 (N_910,In_1666,In_2417);
nand U911 (N_911,In_1681,N_463);
nand U912 (N_912,In_414,In_2291);
nor U913 (N_913,In_1532,In_2331);
nor U914 (N_914,In_42,In_992);
nor U915 (N_915,In_1975,In_1889);
nor U916 (N_916,In_2233,In_219);
or U917 (N_917,In_70,N_263);
nand U918 (N_918,In_1704,In_1095);
and U919 (N_919,In_1897,In_51);
or U920 (N_920,In_930,In_878);
xnor U921 (N_921,N_253,In_616);
xnor U922 (N_922,N_269,In_2136);
nand U923 (N_923,In_2212,In_497);
and U924 (N_924,In_1968,In_2158);
nand U925 (N_925,In_2204,In_1910);
or U926 (N_926,In_2053,In_1647);
nand U927 (N_927,In_2276,N_152);
and U928 (N_928,N_205,N_426);
and U929 (N_929,In_1076,N_126);
xnor U930 (N_930,In_688,In_1923);
nand U931 (N_931,N_167,In_1406);
nand U932 (N_932,In_755,N_452);
nor U933 (N_933,In_2402,N_461);
nand U934 (N_934,In_1810,In_1016);
or U935 (N_935,In_2182,In_57);
or U936 (N_936,In_335,In_1279);
and U937 (N_937,In_1308,In_1359);
or U938 (N_938,In_302,In_2093);
or U939 (N_939,N_368,In_2470);
nor U940 (N_940,In_392,N_19);
xnor U941 (N_941,In_1287,N_22);
xnor U942 (N_942,In_181,N_158);
nor U943 (N_943,N_484,In_2054);
or U944 (N_944,In_1110,In_1519);
or U945 (N_945,N_467,N_72);
xnor U946 (N_946,In_1860,N_417);
and U947 (N_947,In_2324,In_434);
nand U948 (N_948,In_572,In_226);
xor U949 (N_949,In_1478,In_1117);
nor U950 (N_950,In_586,In_1997);
nor U951 (N_951,In_394,In_1222);
xor U952 (N_952,In_1375,In_459);
xor U953 (N_953,In_1379,In_1914);
nand U954 (N_954,In_1270,In_1982);
nor U955 (N_955,In_2001,In_824);
nor U956 (N_956,In_1578,In_1828);
or U957 (N_957,In_186,In_389);
or U958 (N_958,In_482,In_1958);
xor U959 (N_959,In_367,In_1242);
nand U960 (N_960,In_1341,N_142);
xor U961 (N_961,In_579,N_95);
or U962 (N_962,In_555,In_953);
and U963 (N_963,In_788,N_343);
and U964 (N_964,In_1898,N_438);
nand U965 (N_965,In_1820,In_1753);
nor U966 (N_966,In_1162,In_1061);
or U967 (N_967,N_103,N_268);
and U968 (N_968,In_139,In_540);
nor U969 (N_969,In_1137,N_453);
and U970 (N_970,In_672,In_131);
xor U971 (N_971,N_439,In_117);
or U972 (N_972,In_806,In_1972);
and U973 (N_973,In_1018,In_887);
and U974 (N_974,N_180,In_1697);
and U975 (N_975,In_144,In_2137);
or U976 (N_976,In_947,In_2253);
or U977 (N_977,In_1523,In_1127);
and U978 (N_978,N_194,In_1221);
nand U979 (N_979,In_2114,In_607);
or U980 (N_980,In_2426,N_91);
or U981 (N_981,In_938,In_2358);
xnor U982 (N_982,N_155,N_85);
xnor U983 (N_983,N_40,In_2333);
xor U984 (N_984,In_708,N_58);
and U985 (N_985,N_98,In_2246);
nor U986 (N_986,In_1385,In_1802);
and U987 (N_987,In_1328,N_225);
xor U988 (N_988,In_1065,In_539);
nand U989 (N_989,In_1650,In_1888);
nand U990 (N_990,In_604,In_904);
nor U991 (N_991,In_971,In_1074);
xor U992 (N_992,In_751,In_165);
or U993 (N_993,In_1700,In_468);
nor U994 (N_994,In_2021,In_541);
nor U995 (N_995,N_216,N_43);
nor U996 (N_996,N_89,N_76);
xnor U997 (N_997,In_154,In_2463);
and U998 (N_998,In_568,In_931);
xor U999 (N_999,In_933,N_223);
or U1000 (N_1000,N_670,N_249);
or U1001 (N_1001,N_755,N_445);
nor U1002 (N_1002,In_1378,In_1795);
or U1003 (N_1003,In_1688,N_732);
nor U1004 (N_1004,In_990,N_83);
and U1005 (N_1005,In_1533,In_79);
nand U1006 (N_1006,N_446,N_865);
or U1007 (N_1007,In_1970,In_979);
xnor U1008 (N_1008,In_1777,N_371);
or U1009 (N_1009,N_690,In_243);
nand U1010 (N_1010,In_2214,In_2023);
or U1011 (N_1011,In_850,N_108);
or U1012 (N_1012,In_618,N_818);
nand U1013 (N_1013,N_678,N_762);
nand U1014 (N_1014,N_754,N_17);
nor U1015 (N_1015,In_273,N_134);
or U1016 (N_1016,In_637,In_883);
xnor U1017 (N_1017,In_34,In_1039);
xor U1018 (N_1018,In_839,N_561);
nor U1019 (N_1019,In_2432,In_2394);
nor U1020 (N_1020,In_1285,N_861);
nor U1021 (N_1021,N_325,N_705);
or U1022 (N_1022,In_1156,In_490);
or U1023 (N_1023,In_1770,In_1172);
or U1024 (N_1024,In_1477,N_7);
xnor U1025 (N_1025,N_515,In_2097);
nor U1026 (N_1026,In_1290,In_1089);
nand U1027 (N_1027,N_222,In_1930);
or U1028 (N_1028,In_9,N_631);
or U1029 (N_1029,N_362,In_496);
or U1030 (N_1030,N_534,N_950);
xnor U1031 (N_1031,In_2004,In_1193);
nand U1032 (N_1032,In_2033,In_1419);
or U1033 (N_1033,In_2391,N_578);
nand U1034 (N_1034,N_327,In_10);
and U1035 (N_1035,N_501,N_612);
nor U1036 (N_1036,N_626,In_1036);
nand U1037 (N_1037,N_778,In_730);
nor U1038 (N_1038,N_788,N_835);
and U1039 (N_1039,In_1455,In_103);
or U1040 (N_1040,In_1060,In_2484);
xnor U1041 (N_1041,N_886,N_568);
xor U1042 (N_1042,N_99,In_726);
xor U1043 (N_1043,N_455,In_1841);
nor U1044 (N_1044,N_864,N_956);
xnor U1045 (N_1045,In_1491,N_603);
nand U1046 (N_1046,N_198,N_552);
nor U1047 (N_1047,In_2329,N_539);
or U1048 (N_1048,In_1716,N_947);
nor U1049 (N_1049,N_326,N_332);
or U1050 (N_1050,In_1245,In_506);
nor U1051 (N_1051,In_1398,N_757);
or U1052 (N_1052,N_767,N_86);
xnor U1053 (N_1053,N_857,N_405);
or U1054 (N_1054,In_350,N_709);
xor U1055 (N_1055,N_576,N_610);
or U1056 (N_1056,In_1610,In_184);
or U1057 (N_1057,In_136,In_1196);
nand U1058 (N_1058,N_456,N_133);
nand U1059 (N_1059,In_1413,In_215);
xor U1060 (N_1060,N_242,In_326);
xnor U1061 (N_1061,In_1361,N_264);
nand U1062 (N_1062,N_845,N_891);
xor U1063 (N_1063,N_906,N_805);
and U1064 (N_1064,N_676,In_1368);
nor U1065 (N_1065,N_605,In_8);
nand U1066 (N_1066,N_954,N_295);
or U1067 (N_1067,In_551,N_177);
nor U1068 (N_1068,In_1212,In_2155);
nand U1069 (N_1069,In_2043,N_556);
nand U1070 (N_1070,N_796,N_549);
nor U1071 (N_1071,In_673,N_962);
nor U1072 (N_1072,In_1424,N_617);
nand U1073 (N_1073,In_2307,N_661);
nand U1074 (N_1074,In_2321,N_514);
nor U1075 (N_1075,In_2397,N_233);
xor U1076 (N_1076,In_2087,In_2406);
and U1077 (N_1077,N_710,In_1598);
or U1078 (N_1078,In_861,N_248);
and U1079 (N_1079,In_1853,N_599);
xor U1080 (N_1080,N_518,In_1526);
or U1081 (N_1081,In_845,N_719);
and U1082 (N_1082,N_406,In_1551);
xor U1083 (N_1083,N_384,In_1573);
and U1084 (N_1084,N_298,In_347);
and U1085 (N_1085,In_2380,In_1072);
or U1086 (N_1086,In_838,N_554);
and U1087 (N_1087,In_2348,In_145);
or U1088 (N_1088,N_809,N_381);
and U1089 (N_1089,In_859,N_792);
xor U1090 (N_1090,In_1143,N_143);
nand U1091 (N_1091,N_82,N_760);
and U1092 (N_1092,In_1607,N_651);
xor U1093 (N_1093,In_138,In_372);
nor U1094 (N_1094,In_351,N_638);
xor U1095 (N_1095,In_976,In_409);
nand U1096 (N_1096,N_978,In_605);
nor U1097 (N_1097,In_218,N_245);
nand U1098 (N_1098,N_833,In_553);
or U1099 (N_1099,In_1099,N_585);
xnor U1100 (N_1100,N_118,N_211);
nor U1101 (N_1101,N_450,N_695);
nor U1102 (N_1102,In_689,N_877);
and U1103 (N_1103,In_1553,N_746);
or U1104 (N_1104,In_130,In_2012);
or U1105 (N_1105,N_15,N_232);
nor U1106 (N_1106,In_1048,In_1985);
nand U1107 (N_1107,In_722,N_61);
or U1108 (N_1108,In_1353,In_1714);
xor U1109 (N_1109,In_624,In_1778);
and U1110 (N_1110,In_1286,In_207);
nand U1111 (N_1111,N_976,In_1826);
xor U1112 (N_1112,N_201,In_2375);
xor U1113 (N_1113,N_44,N_45);
nor U1114 (N_1114,N_380,N_699);
and U1115 (N_1115,In_1555,In_1453);
xnor U1116 (N_1116,In_1588,N_530);
nor U1117 (N_1117,In_1854,N_572);
xnor U1118 (N_1118,N_824,In_923);
nor U1119 (N_1119,In_505,In_1216);
nor U1120 (N_1120,In_2115,In_2485);
nand U1121 (N_1121,In_438,N_409);
nand U1122 (N_1122,N_600,N_989);
xnor U1123 (N_1123,N_953,N_799);
or U1124 (N_1124,In_2272,In_1952);
xor U1125 (N_1125,In_2244,In_319);
and U1126 (N_1126,In_2143,In_1521);
nor U1127 (N_1127,In_112,In_1676);
xor U1128 (N_1128,N_966,N_562);
or U1129 (N_1129,N_519,In_535);
nor U1130 (N_1130,In_2399,In_1537);
nand U1131 (N_1131,N_442,N_748);
nand U1132 (N_1132,N_227,N_555);
nor U1133 (N_1133,N_606,In_1241);
xor U1134 (N_1134,N_707,N_852);
or U1135 (N_1135,N_219,In_2224);
nor U1136 (N_1136,N_543,N_497);
or U1137 (N_1137,N_960,In_107);
or U1138 (N_1138,In_2260,In_961);
xnor U1139 (N_1139,In_761,In_1336);
xnor U1140 (N_1140,N_291,In_291);
nand U1141 (N_1141,In_1980,In_101);
nor U1142 (N_1142,N_731,In_663);
and U1143 (N_1143,N_479,N_914);
xor U1144 (N_1144,N_62,N_483);
xnor U1145 (N_1145,In_1660,In_1319);
and U1146 (N_1146,N_648,N_995);
and U1147 (N_1147,N_783,N_306);
nand U1148 (N_1148,N_643,In_2448);
nand U1149 (N_1149,N_321,In_1277);
nand U1150 (N_1150,N_957,In_577);
and U1151 (N_1151,N_850,In_1363);
nor U1152 (N_1152,In_246,In_336);
and U1153 (N_1153,In_1393,N_832);
and U1154 (N_1154,N_587,In_2140);
nor U1155 (N_1155,In_1451,In_2101);
or U1156 (N_1156,In_1929,In_1123);
nand U1157 (N_1157,N_759,In_1356);
xor U1158 (N_1158,N_522,N_972);
nor U1159 (N_1159,N_428,In_1808);
nor U1160 (N_1160,In_2337,N_949);
and U1161 (N_1161,In_1879,N_535);
and U1162 (N_1162,In_1566,In_2309);
xor U1163 (N_1163,N_513,N_701);
and U1164 (N_1164,In_1872,In_1427);
or U1165 (N_1165,In_1574,N_997);
nand U1166 (N_1166,In_128,N_730);
xor U1167 (N_1167,In_2452,In_1847);
xnor U1168 (N_1168,In_67,In_1255);
nor U1169 (N_1169,In_1564,In_2314);
nor U1170 (N_1170,In_1575,In_187);
nor U1171 (N_1171,In_1858,In_756);
nand U1172 (N_1172,N_283,In_167);
or U1173 (N_1173,In_775,In_1544);
nand U1174 (N_1174,In_2407,In_2193);
and U1175 (N_1175,N_688,N_734);
xnor U1176 (N_1176,N_107,In_1815);
and U1177 (N_1177,In_1386,N_564);
or U1178 (N_1178,N_681,In_1708);
xnor U1179 (N_1179,In_445,N_271);
nand U1180 (N_1180,N_184,In_2074);
nand U1181 (N_1181,In_1742,N_868);
nand U1182 (N_1182,In_1838,N_684);
nor U1183 (N_1183,N_69,N_862);
nor U1184 (N_1184,In_2124,N_904);
and U1185 (N_1185,N_673,N_821);
nor U1186 (N_1186,In_897,In_1657);
nand U1187 (N_1187,In_1108,N_234);
nor U1188 (N_1188,In_640,In_1570);
or U1189 (N_1189,In_608,N_140);
nand U1190 (N_1190,N_717,In_2473);
nor U1191 (N_1191,In_1921,In_71);
nand U1192 (N_1192,In_1094,In_1590);
nor U1193 (N_1193,In_2128,N_943);
or U1194 (N_1194,N_570,N_892);
and U1195 (N_1195,In_499,N_769);
nor U1196 (N_1196,N_680,In_1907);
xnor U1197 (N_1197,N_341,N_932);
nand U1198 (N_1198,In_706,In_805);
nand U1199 (N_1199,N_540,N_51);
nor U1200 (N_1200,N_980,N_448);
nor U1201 (N_1201,N_975,N_758);
nand U1202 (N_1202,N_842,In_782);
xor U1203 (N_1203,N_878,In_1755);
nor U1204 (N_1204,In_882,N_847);
nand U1205 (N_1205,In_1505,In_489);
xnor U1206 (N_1206,N_738,In_334);
or U1207 (N_1207,In_1589,In_1735);
nor U1208 (N_1208,N_819,N_322);
nor U1209 (N_1209,N_351,N_831);
and U1210 (N_1210,In_242,In_1788);
and U1211 (N_1211,N_683,In_383);
nand U1212 (N_1212,N_628,In_2280);
nand U1213 (N_1213,In_2192,N_729);
nor U1214 (N_1214,N_981,In_1940);
nor U1215 (N_1215,N_279,N_992);
and U1216 (N_1216,N_607,In_1774);
xor U1217 (N_1217,N_623,In_2003);
xnor U1218 (N_1218,N_383,N_413);
nand U1219 (N_1219,N_874,N_888);
nand U1220 (N_1220,N_689,N_971);
nand U1221 (N_1221,In_1088,N_723);
and U1222 (N_1222,N_982,N_385);
xor U1223 (N_1223,N_935,In_1572);
nand U1224 (N_1224,In_1759,In_836);
and U1225 (N_1225,In_2294,In_683);
or U1226 (N_1226,N_667,N_893);
and U1227 (N_1227,N_565,N_524);
xnor U1228 (N_1228,N_987,In_1446);
nand U1229 (N_1229,In_1740,In_2398);
and U1230 (N_1230,In_1892,N_141);
and U1231 (N_1231,N_65,N_804);
or U1232 (N_1232,In_178,In_1208);
nand U1233 (N_1233,In_2123,N_490);
nand U1234 (N_1234,N_318,N_918);
nand U1235 (N_1235,N_708,N_10);
nand U1236 (N_1236,N_189,In_1047);
xor U1237 (N_1237,N_642,In_945);
or U1238 (N_1238,N_724,N_715);
nand U1239 (N_1239,N_485,N_656);
nand U1240 (N_1240,N_998,In_199);
nand U1241 (N_1241,N_553,N_973);
xor U1242 (N_1242,In_1595,N_802);
nor U1243 (N_1243,N_296,In_379);
xor U1244 (N_1244,In_432,In_2005);
and U1245 (N_1245,N_173,In_1686);
nor U1246 (N_1246,N_57,In_750);
nand U1247 (N_1247,N_595,In_1438);
nand U1248 (N_1248,N_915,N_660);
or U1249 (N_1249,In_532,N_907);
nand U1250 (N_1250,In_928,In_1397);
or U1251 (N_1251,In_132,N_722);
or U1252 (N_1252,N_968,N_580);
nor U1253 (N_1253,In_204,N_324);
nor U1254 (N_1254,In_209,N_958);
nand U1255 (N_1255,N_860,In_889);
and U1256 (N_1256,N_486,N_985);
nor U1257 (N_1257,N_646,In_2095);
nor U1258 (N_1258,In_626,In_890);
and U1259 (N_1259,In_817,N_23);
nand U1260 (N_1260,N_922,N_172);
xor U1261 (N_1261,In_1233,In_575);
or U1262 (N_1262,In_1318,N_274);
nand U1263 (N_1263,N_698,In_276);
nor U1264 (N_1264,In_307,In_2157);
or U1265 (N_1265,In_2296,In_2007);
or U1266 (N_1266,N_615,In_1639);
and U1267 (N_1267,N_790,N_756);
nand U1268 (N_1268,In_1405,N_669);
or U1269 (N_1269,In_2434,In_612);
and U1270 (N_1270,N_505,In_1620);
xnor U1271 (N_1271,N_337,In_1068);
nor U1272 (N_1272,In_858,N_54);
xnor U1273 (N_1273,N_192,In_1987);
or U1274 (N_1274,In_397,In_1264);
or U1275 (N_1275,In_2151,N_569);
nand U1276 (N_1276,N_797,N_435);
and U1277 (N_1277,N_712,N_97);
nor U1278 (N_1278,N_267,In_119);
xor U1279 (N_1279,N_838,N_251);
and U1280 (N_1280,N_622,In_1926);
xnor U1281 (N_1281,N_739,In_1623);
and U1282 (N_1282,N_728,N_440);
nor U1283 (N_1283,In_314,N_208);
xor U1284 (N_1284,In_2080,In_2310);
xnor U1285 (N_1285,In_2008,In_2149);
xor U1286 (N_1286,In_2495,N_34);
or U1287 (N_1287,In_821,N_93);
nand U1288 (N_1288,N_601,In_578);
and U1289 (N_1289,N_720,In_1161);
or U1290 (N_1290,N_90,N_774);
and U1291 (N_1291,N_596,N_996);
nand U1292 (N_1292,In_257,In_196);
nand U1293 (N_1293,In_860,In_1787);
nor U1294 (N_1294,In_1130,In_229);
or U1295 (N_1295,In_2282,N_476);
xor U1296 (N_1296,In_793,In_811);
nand U1297 (N_1297,In_321,N_117);
nand U1298 (N_1298,In_274,N_616);
xnor U1299 (N_1299,N_633,N_800);
nand U1300 (N_1300,In_407,N_955);
nor U1301 (N_1301,In_808,N_911);
and U1302 (N_1302,N_557,N_28);
or U1303 (N_1303,N_29,N_115);
nand U1304 (N_1304,In_1515,In_2183);
and U1305 (N_1305,N_830,N_532);
and U1306 (N_1306,In_1354,In_2266);
xor U1307 (N_1307,In_316,In_1609);
xor U1308 (N_1308,In_1939,In_153);
or U1309 (N_1309,In_100,N_551);
or U1310 (N_1310,N_897,In_659);
nand U1311 (N_1311,In_1884,In_2446);
and U1312 (N_1312,N_872,N_338);
and U1313 (N_1313,N_307,N_414);
or U1314 (N_1314,In_1015,In_2261);
nand U1315 (N_1315,N_948,In_1377);
nand U1316 (N_1316,N_841,N_923);
xnor U1317 (N_1317,In_14,N_292);
and U1318 (N_1318,N_647,N_913);
nand U1319 (N_1319,In_1263,N_743);
nor U1320 (N_1320,In_1744,In_309);
nand U1321 (N_1321,N_741,N_694);
xnor U1322 (N_1322,N_546,In_1454);
nor U1323 (N_1323,N_969,N_105);
and U1324 (N_1324,In_919,In_2144);
nor U1325 (N_1325,In_2024,In_648);
nand U1326 (N_1326,N_94,N_196);
nor U1327 (N_1327,N_590,N_939);
nor U1328 (N_1328,N_77,N_851);
nand U1329 (N_1329,In_1731,In_87);
and U1330 (N_1330,In_1584,In_1558);
nor U1331 (N_1331,N_991,N_702);
nand U1332 (N_1332,In_1167,N_733);
and U1333 (N_1333,N_685,N_469);
nand U1334 (N_1334,N_776,In_1895);
and U1335 (N_1335,N_547,N_844);
and U1336 (N_1336,In_1664,N_397);
and U1337 (N_1337,In_1983,N_938);
nor U1338 (N_1338,N_706,N_447);
or U1339 (N_1339,N_745,N_550);
or U1340 (N_1340,N_873,In_641);
nand U1341 (N_1341,N_825,N_793);
or U1342 (N_1342,In_1023,N_473);
nor U1343 (N_1343,N_640,N_591);
nand U1344 (N_1344,In_2493,N_3);
nand U1345 (N_1345,In_567,In_991);
and U1346 (N_1346,N_937,In_716);
and U1347 (N_1347,N_236,N_828);
or U1348 (N_1348,In_1693,N_999);
or U1349 (N_1349,In_519,N_990);
nand U1350 (N_1350,In_1614,N_653);
nor U1351 (N_1351,N_312,N_49);
nand U1352 (N_1352,In_597,N_182);
nand U1353 (N_1353,In_1092,N_185);
nand U1354 (N_1354,N_161,In_812);
or U1355 (N_1355,N_988,In_1075);
xnor U1356 (N_1356,N_794,N_391);
or U1357 (N_1357,In_1781,In_1517);
nand U1358 (N_1358,N_361,In_1769);
and U1359 (N_1359,N_657,In_1303);
or U1360 (N_1360,N_478,In_1513);
and U1361 (N_1361,In_402,N_771);
and U1362 (N_1362,In_820,N_276);
and U1363 (N_1363,N_379,N_696);
xor U1364 (N_1364,N_183,N_639);
or U1365 (N_1365,N_959,In_2351);
nand U1366 (N_1366,In_1392,In_1128);
xor U1367 (N_1367,In_958,In_1545);
xor U1368 (N_1368,N_686,In_590);
nand U1369 (N_1369,In_224,In_1410);
nor U1370 (N_1370,In_816,N_619);
nor U1371 (N_1371,N_856,In_749);
nand U1372 (N_1372,N_545,In_1366);
or U1373 (N_1373,In_1400,In_2454);
nand U1374 (N_1374,In_1606,N_986);
and U1375 (N_1375,N_930,In_939);
and U1376 (N_1376,In_1900,In_1846);
nor U1377 (N_1377,In_576,In_1081);
and U1378 (N_1378,In_1338,In_1857);
nor U1379 (N_1379,N_837,N_931);
and U1380 (N_1380,In_968,N_876);
and U1381 (N_1381,N_713,In_1922);
nand U1382 (N_1382,In_1090,In_35);
xor U1383 (N_1383,In_2433,N_399);
nand U1384 (N_1384,N_772,In_528);
xnor U1385 (N_1385,In_1010,In_2156);
nor U1386 (N_1386,N_855,In_37);
or U1387 (N_1387,N_301,In_137);
or U1388 (N_1388,N_944,In_1444);
and U1389 (N_1389,In_2173,N_462);
nand U1390 (N_1390,N_905,In_1756);
or U1391 (N_1391,N_261,In_2072);
nor U1392 (N_1392,N_840,N_588);
xnor U1393 (N_1393,N_806,N_593);
nand U1394 (N_1394,N_353,In_655);
nor U1395 (N_1395,N_579,In_2271);
and U1396 (N_1396,N_47,N_674);
nand U1397 (N_1397,N_320,N_487);
and U1398 (N_1398,In_453,N_247);
nand U1399 (N_1399,N_567,In_2085);
and U1400 (N_1400,N_297,N_508);
xnor U1401 (N_1401,In_241,N_544);
nand U1402 (N_1402,In_2355,N_787);
and U1403 (N_1403,N_951,In_1391);
nand U1404 (N_1404,N_330,N_359);
nor U1405 (N_1405,In_1138,In_1464);
or U1406 (N_1406,In_91,In_682);
nor U1407 (N_1407,N_721,In_206);
or U1408 (N_1408,N_727,N_909);
nand U1409 (N_1409,N_898,N_945);
or U1410 (N_1410,In_2303,N_675);
nand U1411 (N_1411,N_889,N_736);
xor U1412 (N_1412,In_2121,In_259);
and U1413 (N_1413,N_903,N_773);
nor U1414 (N_1414,In_652,In_1007);
nor U1415 (N_1415,In_754,N_620);
nor U1416 (N_1416,N_714,N_649);
and U1417 (N_1417,In_962,In_278);
xor U1418 (N_1418,N_170,N_536);
xor U1419 (N_1419,In_1843,In_386);
nor U1420 (N_1420,N_598,In_1959);
or U1421 (N_1421,In_1779,In_1896);
or U1422 (N_1422,N_940,In_815);
nand U1423 (N_1423,In_2496,In_124);
nand U1424 (N_1424,N_589,In_2027);
nand U1425 (N_1425,In_1272,In_526);
nor U1426 (N_1426,In_454,N_781);
and U1427 (N_1427,In_1407,N_816);
or U1428 (N_1428,N_735,In_552);
nand U1429 (N_1429,N_102,In_27);
nand U1430 (N_1430,N_503,N_994);
nor U1431 (N_1431,N_416,In_2458);
and U1432 (N_1432,N_652,N_716);
xor U1433 (N_1433,N_894,N_339);
or U1434 (N_1434,In_701,In_1168);
nand U1435 (N_1435,In_2293,In_2352);
nand U1436 (N_1436,N_401,N_866);
nand U1437 (N_1437,N_285,In_405);
nand U1438 (N_1438,N_81,In_1662);
nand U1439 (N_1439,In_1723,In_770);
and U1440 (N_1440,N_146,In_1960);
nor U1441 (N_1441,In_330,In_1655);
and U1442 (N_1442,N_859,N_933);
xnor U1443 (N_1443,In_1986,N_650);
and U1444 (N_1444,N_843,N_506);
and U1445 (N_1445,N_472,In_791);
and U1446 (N_1446,In_1267,N_899);
xor U1447 (N_1447,N_820,N_520);
xor U1448 (N_1448,In_646,N_541);
nor U1449 (N_1449,N_70,N_789);
xnor U1450 (N_1450,N_703,N_533);
or U1451 (N_1451,In_1518,N_125);
nand U1452 (N_1452,In_283,N_895);
xor U1453 (N_1453,In_1293,In_794);
nor U1454 (N_1454,N_896,In_1903);
and U1455 (N_1455,N_692,N_668);
nand U1456 (N_1456,N_636,In_1507);
xnor U1457 (N_1457,In_1748,N_243);
or U1458 (N_1458,In_1534,In_1966);
or U1459 (N_1459,In_61,N_31);
or U1460 (N_1460,N_654,In_303);
nand U1461 (N_1461,N_410,In_2075);
nand U1462 (N_1462,In_161,N_846);
or U1463 (N_1463,In_1383,N_558);
and U1464 (N_1464,N_983,N_8);
and U1465 (N_1465,N_849,In_195);
and U1466 (N_1466,N_700,In_2283);
or U1467 (N_1467,N_687,N_444);
xor U1468 (N_1468,In_718,N_934);
and U1469 (N_1469,In_511,N_900);
xor U1470 (N_1470,In_2267,In_33);
and U1471 (N_1471,N_168,In_1107);
xnor U1472 (N_1472,N_967,N_869);
nor U1473 (N_1473,N_502,N_697);
or U1474 (N_1474,In_965,In_1724);
nor U1475 (N_1475,N_363,In_2466);
and U1476 (N_1476,In_1596,In_2364);
nor U1477 (N_1477,In_251,N_691);
xor U1478 (N_1478,N_495,N_910);
xor U1479 (N_1479,In_349,N_827);
and U1480 (N_1480,N_110,N_753);
or U1481 (N_1481,N_765,N_304);
nor U1482 (N_1482,In_1669,In_2160);
and U1483 (N_1483,N_890,In_738);
nand U1484 (N_1484,N_621,N_181);
nor U1485 (N_1485,N_763,N_592);
and U1486 (N_1486,N_214,In_1214);
nor U1487 (N_1487,N_637,N_659);
nor U1488 (N_1488,In_299,N_186);
xnor U1489 (N_1489,In_585,In_1499);
nor U1490 (N_1490,N_504,In_1416);
xor U1491 (N_1491,In_2161,In_864);
nor U1492 (N_1492,In_1822,N_764);
nand U1493 (N_1493,In_102,N_521);
xor U1494 (N_1494,In_19,N_238);
or U1495 (N_1495,In_932,N_791);
nor U1496 (N_1496,In_2477,In_1712);
xnor U1497 (N_1497,N_12,N_516);
xnor U1498 (N_1498,N_925,N_305);
xor U1499 (N_1499,N_655,N_965);
and U1500 (N_1500,N_1260,In_41);
and U1501 (N_1501,In_1125,N_884);
nand U1502 (N_1502,N_1323,N_834);
or U1503 (N_1503,N_1482,N_1443);
or U1504 (N_1504,In_2047,N_1052);
or U1505 (N_1505,N_1269,N_53);
or U1506 (N_1506,N_777,N_1177);
xnor U1507 (N_1507,N_1301,N_1470);
nand U1508 (N_1508,N_1079,N_1174);
nand U1509 (N_1509,N_1330,N_1355);
and U1510 (N_1510,N_1200,In_1173);
nor U1511 (N_1511,In_52,N_677);
and U1512 (N_1512,In_1136,N_1005);
or U1513 (N_1513,N_1387,N_1137);
or U1514 (N_1514,N_1149,N_823);
nor U1515 (N_1515,In_375,In_2376);
and U1516 (N_1516,In_2186,N_1311);
and U1517 (N_1517,In_406,N_581);
or U1518 (N_1518,N_525,N_807);
nor U1519 (N_1519,N_1155,N_460);
nand U1520 (N_1520,N_1440,N_512);
nor U1521 (N_1521,In_216,N_1435);
nand U1522 (N_1522,N_1036,N_597);
or U1523 (N_1523,N_1153,In_1261);
nor U1524 (N_1524,N_1172,N_1432);
nand U1525 (N_1525,N_120,N_974);
or U1526 (N_1526,N_87,N_858);
xnor U1527 (N_1527,N_1389,N_527);
xnor U1528 (N_1528,In_1632,In_1635);
nor U1529 (N_1529,N_357,N_465);
nand U1530 (N_1530,N_1442,N_1407);
and U1531 (N_1531,In_2304,N_815);
xor U1532 (N_1532,N_577,N_129);
and U1533 (N_1533,N_682,N_1170);
nor U1534 (N_1534,N_1481,N_1233);
or U1535 (N_1535,N_1126,N_936);
and U1536 (N_1536,In_2494,In_1836);
or U1537 (N_1537,N_537,N_230);
and U1538 (N_1538,N_1077,N_531);
nand U1539 (N_1539,N_1277,In_2238);
nand U1540 (N_1540,N_1019,N_1000);
xnor U1541 (N_1541,In_275,N_1264);
or U1542 (N_1542,N_1123,N_1050);
nand U1543 (N_1543,In_768,N_1043);
or U1544 (N_1544,N_52,In_1561);
or U1545 (N_1545,In_2052,N_1478);
nand U1546 (N_1546,N_1082,N_35);
nor U1547 (N_1547,N_1109,N_407);
and U1548 (N_1548,N_1038,N_1376);
xnor U1549 (N_1549,N_1015,In_361);
xor U1550 (N_1550,N_1310,In_2489);
nand U1551 (N_1551,N_1493,In_2354);
or U1552 (N_1552,In_404,N_390);
xor U1553 (N_1553,In_2379,N_1122);
nor U1554 (N_1554,N_1114,N_1142);
and U1555 (N_1555,N_1430,N_441);
and U1556 (N_1556,N_25,N_1445);
xor U1557 (N_1557,In_1615,In_1266);
nand U1558 (N_1558,In_20,In_573);
and U1559 (N_1559,N_1255,N_1437);
xnor U1560 (N_1560,N_433,N_630);
and U1561 (N_1561,In_702,In_884);
xnor U1562 (N_1562,N_1162,N_1);
or U1563 (N_1563,N_801,N_1148);
and U1564 (N_1564,In_2213,N_266);
xnor U1565 (N_1565,In_721,In_1370);
nor U1566 (N_1566,N_30,In_855);
nand U1567 (N_1567,In_2269,In_818);
xor U1568 (N_1568,N_1163,In_272);
and U1569 (N_1569,In_21,N_1419);
or U1570 (N_1570,N_1468,N_1349);
and U1571 (N_1571,N_1438,N_1318);
nor U1572 (N_1572,N_644,In_636);
nand U1573 (N_1573,N_870,N_826);
nand U1574 (N_1574,In_0,N_1007);
nor U1575 (N_1575,In_670,N_1199);
nand U1576 (N_1576,N_1307,In_2089);
nand U1577 (N_1577,N_244,N_1409);
nor U1578 (N_1578,N_1104,N_1495);
xnor U1579 (N_1579,N_1476,In_1979);
and U1580 (N_1580,N_1124,In_1165);
or U1581 (N_1581,N_1106,N_1395);
xnor U1582 (N_1582,N_116,In_1460);
xnor U1583 (N_1583,N_1127,N_917);
xnor U1584 (N_1584,In_1741,N_1382);
or U1585 (N_1585,N_928,N_1188);
or U1586 (N_1586,N_1203,N_1096);
or U1587 (N_1587,N_1384,In_2131);
nor U1588 (N_1588,N_1088,N_1178);
nor U1589 (N_1589,N_1029,N_1378);
nand U1590 (N_1590,N_1207,N_1267);
xor U1591 (N_1591,N_1282,N_1185);
and U1592 (N_1592,N_1131,N_766);
nand U1593 (N_1593,In_828,N_779);
and U1594 (N_1594,N_1371,In_177);
xor U1595 (N_1595,N_871,In_2049);
or U1596 (N_1596,N_1021,N_1105);
and U1597 (N_1597,In_2300,In_1249);
and U1598 (N_1598,In_2134,In_935);
nand U1599 (N_1599,In_282,N_151);
and U1600 (N_1600,N_586,N_1164);
nand U1601 (N_1601,In_1298,In_151);
and U1602 (N_1602,In_1563,In_1244);
nor U1603 (N_1603,N_1014,N_1464);
and U1604 (N_1604,N_1173,N_1219);
or U1605 (N_1605,In_559,In_1962);
xor U1606 (N_1606,N_1003,N_1253);
xnor U1607 (N_1607,N_1192,N_1097);
xor U1608 (N_1608,N_1487,N_1074);
nor U1609 (N_1609,In_694,In_1239);
xor U1610 (N_1610,N_786,N_1313);
nor U1611 (N_1611,In_713,N_635);
nand U1612 (N_1612,N_902,N_566);
and U1613 (N_1613,N_1364,N_1008);
and U1614 (N_1614,N_1471,In_425);
nor U1615 (N_1615,N_1449,N_1402);
and U1616 (N_1616,N_112,N_1211);
nand U1617 (N_1617,N_725,N_1386);
nor U1618 (N_1618,N_1280,N_1147);
nand U1619 (N_1619,N_1010,N_1224);
nor U1620 (N_1620,N_1337,N_1473);
nand U1621 (N_1621,In_1861,N_139);
nand U1622 (N_1622,In_2111,N_1319);
nand U1623 (N_1623,In_942,N_1499);
and U1624 (N_1624,N_1216,N_1227);
nor U1625 (N_1625,N_1416,N_1099);
or U1626 (N_1626,N_1314,In_1497);
nor U1627 (N_1627,In_2241,N_1228);
nor U1628 (N_1628,N_1210,N_1257);
or U1629 (N_1629,In_554,In_2210);
nor U1630 (N_1630,N_1071,In_1602);
nor U1631 (N_1631,N_1394,N_970);
xnor U1632 (N_1632,N_1370,In_814);
nor U1633 (N_1633,N_1143,N_344);
or U1634 (N_1634,N_213,In_233);
nand U1635 (N_1635,In_915,N_1362);
or U1636 (N_1636,N_1201,N_1139);
nand U1637 (N_1637,N_614,N_1235);
nand U1638 (N_1638,N_1133,N_1463);
and U1639 (N_1639,N_1278,N_348);
nor U1640 (N_1640,In_311,N_1299);
xor U1641 (N_1641,In_611,N_1102);
and U1642 (N_1642,N_812,N_1193);
nor U1643 (N_1643,In_1508,N_704);
nor U1644 (N_1644,In_1592,N_1061);
nor U1645 (N_1645,N_403,N_164);
and U1646 (N_1646,N_317,N_1369);
xor U1647 (N_1647,N_1455,N_0);
xnor U1648 (N_1648,N_148,N_1294);
and U1649 (N_1649,In_2081,N_761);
nor U1650 (N_1650,In_1991,N_665);
and U1651 (N_1651,N_1275,N_604);
nor U1652 (N_1652,N_1348,N_1251);
and U1653 (N_1653,In_1339,In_2088);
nor U1654 (N_1654,In_1739,In_1329);
or U1655 (N_1655,N_287,N_1453);
nor U1656 (N_1656,N_1424,N_1128);
and U1657 (N_1657,N_1169,N_538);
or U1658 (N_1658,N_1171,N_919);
nor U1659 (N_1659,N_1191,N_1067);
or U1660 (N_1660,N_529,N_1297);
and U1661 (N_1661,N_50,N_1334);
nor U1662 (N_1662,N_1009,N_1321);
xnor U1663 (N_1663,N_1373,N_1232);
nand U1664 (N_1664,N_881,N_658);
xnor U1665 (N_1665,N_1347,N_1031);
nor U1666 (N_1666,N_582,In_2079);
nor U1667 (N_1667,N_1475,In_1875);
nand U1668 (N_1668,N_1156,N_1136);
nand U1669 (N_1669,N_671,N_1087);
or U1670 (N_1670,N_542,In_2109);
and U1671 (N_1671,In_1231,N_1144);
xnor U1672 (N_1672,N_354,N_1064);
xor U1673 (N_1673,In_1115,N_1439);
nand U1674 (N_1674,In_269,N_500);
xnor U1675 (N_1675,N_1306,N_1249);
nor U1676 (N_1676,In_1423,N_1022);
and U1677 (N_1677,N_111,N_1418);
xnor U1678 (N_1678,N_488,N_1065);
xor U1679 (N_1679,In_797,N_879);
and U1680 (N_1680,N_740,In_591);
and U1681 (N_1681,In_134,N_618);
and U1682 (N_1682,In_2264,N_1085);
or U1683 (N_1683,N_1119,N_875);
nand U1684 (N_1684,N_1316,N_1187);
nand U1685 (N_1685,In_148,N_1161);
nand U1686 (N_1686,In_271,N_1035);
and U1687 (N_1687,N_1190,In_1528);
xor U1688 (N_1688,N_1168,N_1302);
nand U1689 (N_1689,N_1483,N_1115);
xor U1690 (N_1690,N_1154,N_780);
nor U1691 (N_1691,N_1381,In_498);
and U1692 (N_1692,N_310,N_509);
nand U1693 (N_1693,N_1477,In_835);
nand U1694 (N_1694,N_775,N_813);
nand U1695 (N_1695,N_1125,N_1324);
nand U1696 (N_1696,N_768,N_920);
and U1697 (N_1697,N_517,In_2083);
xor U1698 (N_1698,N_375,N_1240);
nand U1699 (N_1699,N_1412,In_631);
xnor U1700 (N_1700,N_726,N_1237);
nor U1701 (N_1701,In_530,N_1141);
xnor U1702 (N_1702,N_853,N_1157);
nor U1703 (N_1703,N_784,N_1268);
nor U1704 (N_1704,N_1265,N_1095);
xnor U1705 (N_1705,N_1338,N_1048);
nor U1706 (N_1706,N_1377,N_836);
xnor U1707 (N_1707,N_1456,N_882);
nand U1708 (N_1708,N_829,In_1866);
xor U1709 (N_1709,N_209,N_1180);
and U1710 (N_1710,N_1182,N_672);
nor U1711 (N_1711,N_1421,N_1243);
or U1712 (N_1712,In_2207,N_1289);
nand U1713 (N_1713,N_663,N_1335);
xor U1714 (N_1714,N_1375,In_318);
nand U1715 (N_1715,In_2447,N_1341);
or U1716 (N_1716,N_750,In_2453);
xnor U1717 (N_1717,N_609,N_693);
nand U1718 (N_1718,N_1030,In_230);
or U1719 (N_1719,In_1732,N_1111);
xor U1720 (N_1720,N_1049,N_548);
and U1721 (N_1721,N_382,N_1283);
or U1722 (N_1722,In_2289,In_1140);
nand U1723 (N_1723,N_451,In_1037);
xnor U1724 (N_1724,N_629,N_1189);
nand U1725 (N_1725,N_1120,In_479);
xor U1726 (N_1726,N_1217,N_1056);
or U1727 (N_1727,N_1293,N_1223);
nor U1728 (N_1728,N_1057,N_1467);
nor U1729 (N_1729,In_581,N_1285);
nand U1730 (N_1730,N_1261,N_1046);
nor U1731 (N_1731,In_1784,N_215);
nor U1732 (N_1732,N_1436,N_1206);
xnor U1733 (N_1733,N_1315,In_255);
nand U1734 (N_1734,N_885,N_395);
nand U1735 (N_1735,N_1051,In_603);
nand U1736 (N_1736,N_1460,N_156);
nor U1737 (N_1737,N_1300,In_1113);
or U1738 (N_1738,In_951,N_1028);
xnor U1739 (N_1739,N_1037,N_1291);
and U1740 (N_1740,N_1469,N_1452);
nand U1741 (N_1741,N_131,N_839);
nand U1742 (N_1742,N_1359,In_460);
nor U1743 (N_1743,N_946,N_1336);
nand U1744 (N_1744,N_1413,N_1252);
xor U1745 (N_1745,N_1428,N_1184);
nor U1746 (N_1746,In_90,In_493);
xor U1747 (N_1747,N_1247,In_1608);
nor U1748 (N_1748,N_883,N_511);
and U1749 (N_1749,In_1887,In_244);
and U1750 (N_1750,N_1086,N_744);
or U1751 (N_1751,N_489,N_916);
or U1752 (N_1752,In_369,N_5);
xor U1753 (N_1753,N_1461,N_1399);
nand U1754 (N_1754,N_747,N_1308);
xor U1755 (N_1755,In_766,In_1141);
and U1756 (N_1756,N_1360,N_563);
or U1757 (N_1757,In_1142,N_632);
or U1758 (N_1758,N_921,N_1462);
or U1759 (N_1759,In_1984,N_280);
nand U1760 (N_1760,N_1198,N_1118);
or U1761 (N_1761,In_2290,N_1352);
xnor U1762 (N_1762,In_1388,N_718);
or U1763 (N_1763,N_1140,N_1179);
nand U1764 (N_1764,N_1103,In_879);
nor U1765 (N_1765,In_628,N_1298);
and U1766 (N_1766,N_1447,N_627);
and U1767 (N_1767,In_1612,N_1411);
nand U1768 (N_1768,N_941,N_1112);
and U1769 (N_1769,N_1368,N_470);
or U1770 (N_1770,N_1374,N_863);
xnor U1771 (N_1771,N_560,N_1006);
or U1772 (N_1772,N_1072,N_1151);
xnor U1773 (N_1773,N_1250,N_1342);
and U1774 (N_1774,N_1379,N_1351);
nand U1775 (N_1775,N_1328,N_1215);
nand U1776 (N_1776,N_1242,N_1183);
nand U1777 (N_1777,In_1432,N_634);
or U1778 (N_1778,N_1152,N_1290);
xnor U1779 (N_1779,In_1496,N_1309);
nor U1780 (N_1780,In_2438,N_1066);
or U1781 (N_1781,N_1466,N_1357);
and U1782 (N_1782,In_717,N_1134);
or U1783 (N_1783,N_1167,N_1304);
and U1784 (N_1784,N_1098,N_584);
nand U1785 (N_1785,In_2461,N_402);
nand U1786 (N_1786,N_1132,In_110);
and U1787 (N_1787,In_1622,N_1108);
and U1788 (N_1788,N_422,N_594);
xnor U1789 (N_1789,In_1571,N_1488);
or U1790 (N_1790,In_1539,N_1405);
nor U1791 (N_1791,N_174,N_1117);
and U1792 (N_1792,N_1209,N_1013);
nor U1793 (N_1793,In_2,N_1404);
nand U1794 (N_1794,In_1058,N_1146);
and U1795 (N_1795,In_1063,N_1055);
and U1796 (N_1796,N_1248,In_484);
and U1797 (N_1797,N_1459,N_908);
nor U1798 (N_1798,N_78,In_1813);
and U1799 (N_1799,N_59,N_1365);
xor U1800 (N_1800,N_1479,N_1480);
xor U1801 (N_1801,N_1281,N_257);
nor U1802 (N_1802,N_1230,In_366);
and U1803 (N_1803,In_2342,N_1286);
xor U1804 (N_1804,N_1084,N_1083);
nor U1805 (N_1805,N_1353,In_332);
and U1806 (N_1806,In_924,In_78);
nand U1807 (N_1807,N_1166,In_1992);
nand U1808 (N_1808,N_1231,In_767);
and U1809 (N_1809,N_742,In_411);
xor U1810 (N_1810,N_1401,In_1812);
or U1811 (N_1811,In_903,In_30);
xnor U1812 (N_1812,N_1040,N_1059);
and U1813 (N_1813,N_770,N_608);
or U1814 (N_1814,In_513,N_1288);
xnor U1815 (N_1815,N_1380,N_1214);
and U1816 (N_1816,N_1327,In_437);
nor U1817 (N_1817,N_262,N_1069);
and U1818 (N_1818,N_848,N_624);
or U1819 (N_1819,N_1121,N_1110);
nor U1820 (N_1820,N_1089,In_2102);
nand U1821 (N_1821,In_458,In_1490);
nor U1822 (N_1822,N_1236,N_1238);
and U1823 (N_1823,N_573,N_1062);
and U1824 (N_1824,N_1091,N_1017);
and U1825 (N_1825,N_785,N_1457);
nor U1826 (N_1826,N_1033,N_1354);
xor U1827 (N_1827,In_1475,N_1465);
nor U1828 (N_1828,N_964,N_1047);
xnor U1829 (N_1829,N_176,N_810);
and U1830 (N_1830,N_803,N_641);
or U1831 (N_1831,N_1486,In_223);
or U1832 (N_1832,In_2468,N_1498);
nor U1833 (N_1833,In_872,In_1619);
xor U1834 (N_1834,In_442,N_979);
xnor U1835 (N_1835,N_1295,N_1361);
and U1836 (N_1836,N_880,N_1444);
nand U1837 (N_1837,N_175,N_1410);
or U1838 (N_1838,N_1212,N_137);
xnor U1839 (N_1839,N_1372,N_1241);
and U1840 (N_1840,In_1996,In_1536);
xnor U1841 (N_1841,N_507,N_80);
xor U1842 (N_1842,N_1490,N_1181);
and U1843 (N_1843,In_1600,N_1060);
and U1844 (N_1844,N_1417,In_1182);
nand U1845 (N_1845,N_1345,N_571);
nor U1846 (N_1846,N_1329,In_1792);
nor U1847 (N_1847,N_1333,In_745);
xnor U1848 (N_1848,N_1326,N_1239);
and U1849 (N_1849,In_1757,N_1363);
nand U1850 (N_1850,In_1568,N_195);
and U1851 (N_1851,N_425,N_1305);
nand U1852 (N_1852,N_1397,N_752);
and U1853 (N_1853,In_1440,N_1346);
xor U1854 (N_1854,N_1340,N_1350);
xor U1855 (N_1855,N_1150,N_1011);
and U1856 (N_1856,In_1174,N_751);
nor U1857 (N_1857,In_907,N_1358);
or U1858 (N_1858,In_1747,N_154);
nor U1859 (N_1859,N_1303,N_1018);
nand U1860 (N_1860,N_666,In_2169);
and U1861 (N_1861,N_1393,N_510);
nand U1862 (N_1862,N_1234,N_1070);
xnor U1863 (N_1863,N_1023,In_54);
and U1864 (N_1864,N_1012,N_1408);
nand U1865 (N_1865,In_684,N_1080);
or U1866 (N_1866,N_1398,In_1155);
nand U1867 (N_1867,N_1165,N_1415);
xnor U1868 (N_1868,N_1220,N_1202);
xnor U1869 (N_1869,N_160,In_1837);
nand U1870 (N_1870,N_1196,N_1276);
nor U1871 (N_1871,N_737,N_1054);
nor U1872 (N_1872,In_2219,N_1312);
and U1873 (N_1873,In_1931,N_41);
and U1874 (N_1874,N_1063,N_1039);
and U1875 (N_1875,N_1279,N_1317);
or U1876 (N_1876,N_1383,N_993);
nor U1877 (N_1877,In_2051,N_1058);
and U1878 (N_1878,In_322,In_1280);
nand U1879 (N_1879,In_346,N_798);
and U1880 (N_1880,N_1497,In_2050);
nor U1881 (N_1881,N_1366,N_1076);
nor U1882 (N_1882,In_83,N_1472);
nor U1883 (N_1883,N_1422,N_662);
nand U1884 (N_1884,N_1458,N_1053);
or U1885 (N_1885,N_1429,N_526);
nor U1886 (N_1886,In_746,N_388);
or U1887 (N_1887,N_1263,N_477);
or U1888 (N_1888,N_1426,N_952);
nor U1889 (N_1889,N_1130,N_1222);
nor U1890 (N_1890,N_32,N_1175);
or U1891 (N_1891,In_542,N_811);
nand U1892 (N_1892,N_942,In_2320);
xor U1893 (N_1893,In_1674,N_1474);
nor U1894 (N_1894,N_711,N_1414);
and U1895 (N_1895,N_1068,N_1266);
nand U1896 (N_1896,N_1396,N_1256);
and U1897 (N_1897,In_635,N_1274);
xnor U1898 (N_1898,N_1259,N_20);
nor U1899 (N_1899,In_82,In_1365);
nor U1900 (N_1900,N_679,In_1869);
and U1901 (N_1901,N_114,N_1073);
or U1902 (N_1902,N_491,In_550);
xnor U1903 (N_1903,In_941,N_1425);
xnor U1904 (N_1904,N_782,In_1017);
and U1905 (N_1905,In_1260,N_1101);
nor U1906 (N_1906,N_254,N_1245);
or U1907 (N_1907,N_1041,N_39);
nand U1908 (N_1908,N_1129,N_1258);
nand U1909 (N_1909,N_1208,N_1025);
or U1910 (N_1910,N_602,N_328);
nor U1911 (N_1911,N_1001,N_1221);
nor U1912 (N_1912,In_1135,N_1244);
xnor U1913 (N_1913,In_24,In_1306);
nor U1914 (N_1914,N_1094,N_1107);
nor U1915 (N_1915,N_1491,In_998);
or U1916 (N_1916,N_1400,N_822);
nor U1917 (N_1917,N_528,N_145);
nand U1918 (N_1918,N_1044,N_1420);
nand U1919 (N_1919,In_2258,N_523);
and U1920 (N_1920,N_1045,In_179);
and U1921 (N_1921,N_1160,N_1385);
nand U1922 (N_1922,In_1745,N_1213);
nor U1923 (N_1923,N_1138,In_1754);
or U1924 (N_1924,N_1296,N_817);
nor U1925 (N_1925,N_575,N_1496);
xor U1926 (N_1926,In_1621,N_1434);
and U1927 (N_1927,N_645,In_792);
nand U1928 (N_1928,N_1135,In_436);
xnor U1929 (N_1929,In_1447,N_1406);
or U1930 (N_1930,N_1431,N_1331);
and U1931 (N_1931,N_1032,In_485);
or U1932 (N_1932,In_936,In_2163);
nand U1933 (N_1933,In_2404,N_1100);
xor U1934 (N_1934,N_574,N_1034);
and U1935 (N_1935,N_1262,N_1284);
nor U1936 (N_1936,N_1494,N_961);
nor U1937 (N_1937,N_1090,In_478);
nand U1938 (N_1938,N_1081,N_749);
nor U1939 (N_1939,N_241,In_1751);
or U1940 (N_1940,N_795,In_1653);
and U1941 (N_1941,N_128,N_1344);
nand U1942 (N_1942,N_1320,In_2346);
xor U1943 (N_1943,N_1403,In_1333);
xnor U1944 (N_1944,N_1343,N_613);
nand U1945 (N_1945,N_1392,N_1195);
xnor U1946 (N_1946,N_1205,N_1226);
or U1947 (N_1947,N_1042,N_1454);
and U1948 (N_1948,N_977,N_104);
and U1949 (N_1949,In_2403,In_2306);
nand U1950 (N_1950,In_1073,In_974);
xor U1951 (N_1951,In_841,N_169);
nand U1952 (N_1952,N_1485,N_1332);
xor U1953 (N_1953,In_1439,N_1391);
xnor U1954 (N_1954,N_625,In_985);
xor U1955 (N_1955,N_1002,In_1840);
xor U1956 (N_1956,N_887,N_1441);
nor U1957 (N_1957,N_1292,N_1254);
and U1958 (N_1958,N_926,N_559);
and U1959 (N_1959,N_1446,N_1027);
xor U1960 (N_1960,N_912,N_901);
or U1961 (N_1961,N_1075,N_1489);
and U1962 (N_1962,N_252,N_1218);
xor U1963 (N_1963,N_1390,In_2166);
and U1964 (N_1964,N_1186,In_1882);
xnor U1965 (N_1965,N_927,N_924);
or U1966 (N_1966,N_808,In_1305);
nor U1967 (N_1967,N_1020,N_1356);
nor U1968 (N_1968,N_1145,N_1427);
nand U1969 (N_1969,N_664,N_929);
or U1970 (N_1970,N_854,N_1004);
or U1971 (N_1971,N_984,N_68);
and U1972 (N_1972,In_298,In_2455);
and U1973 (N_1973,In_1684,N_1273);
or U1974 (N_1974,N_1451,N_1158);
xor U1975 (N_1975,N_1113,N_1024);
nand U1976 (N_1976,N_1325,N_1287);
nor U1977 (N_1977,N_1423,N_1197);
or U1978 (N_1978,N_1194,N_235);
xor U1979 (N_1979,N_611,N_1272);
xor U1980 (N_1980,In_645,N_1270);
and U1981 (N_1981,In_1525,In_249);
xnor U1982 (N_1982,N_1016,N_1116);
or U1983 (N_1983,N_1339,N_814);
and U1984 (N_1984,N_278,N_1367);
nand U1985 (N_1985,N_1433,N_867);
or U1986 (N_1986,N_1159,N_210);
or U1987 (N_1987,N_1450,In_2263);
or U1988 (N_1988,N_1092,N_1322);
nor U1989 (N_1989,In_777,In_2474);
nor U1990 (N_1990,N_1225,N_1026);
xor U1991 (N_1991,N_1078,N_259);
and U1992 (N_1992,In_1281,N_583);
nand U1993 (N_1993,N_1246,N_963);
nor U1994 (N_1994,N_1204,N_9);
nor U1995 (N_1995,N_1093,N_1492);
and U1996 (N_1996,N_1484,N_1176);
nand U1997 (N_1997,N_1388,N_1229);
nand U1998 (N_1998,In_963,N_1271);
or U1999 (N_1999,In_1948,N_1448);
nand U2000 (N_2000,N_1657,N_1725);
and U2001 (N_2001,N_1849,N_1708);
or U2002 (N_2002,N_1642,N_1518);
and U2003 (N_2003,N_1886,N_1775);
nand U2004 (N_2004,N_1617,N_1624);
xor U2005 (N_2005,N_1771,N_1830);
and U2006 (N_2006,N_1804,N_1580);
and U2007 (N_2007,N_1542,N_1773);
or U2008 (N_2008,N_1680,N_1789);
nand U2009 (N_2009,N_1838,N_1857);
and U2010 (N_2010,N_1908,N_1807);
nor U2011 (N_2011,N_1893,N_1998);
nor U2012 (N_2012,N_1803,N_1595);
or U2013 (N_2013,N_1841,N_1974);
and U2014 (N_2014,N_1983,N_1628);
nor U2015 (N_2015,N_1932,N_1823);
or U2016 (N_2016,N_1770,N_1952);
and U2017 (N_2017,N_1612,N_1977);
nor U2018 (N_2018,N_1697,N_1829);
nor U2019 (N_2019,N_1756,N_1751);
xor U2020 (N_2020,N_1967,N_1722);
xor U2021 (N_2021,N_1997,N_1860);
and U2022 (N_2022,N_1545,N_1840);
or U2023 (N_2023,N_1676,N_1909);
nor U2024 (N_2024,N_1723,N_1558);
xor U2025 (N_2025,N_1635,N_1970);
or U2026 (N_2026,N_1714,N_1815);
xnor U2027 (N_2027,N_1702,N_1929);
xor U2028 (N_2028,N_1587,N_1761);
nand U2029 (N_2029,N_1647,N_1832);
nor U2030 (N_2030,N_1745,N_1623);
or U2031 (N_2031,N_1957,N_1851);
nor U2032 (N_2032,N_1837,N_1910);
or U2033 (N_2033,N_1781,N_1821);
nor U2034 (N_2034,N_1561,N_1596);
xnor U2035 (N_2035,N_1964,N_1514);
xnor U2036 (N_2036,N_1577,N_1520);
xnor U2037 (N_2037,N_1777,N_1716);
nand U2038 (N_2038,N_1986,N_1724);
or U2039 (N_2039,N_1704,N_1573);
nor U2040 (N_2040,N_1755,N_1950);
and U2041 (N_2041,N_1850,N_1913);
xnor U2042 (N_2042,N_1728,N_1656);
nand U2043 (N_2043,N_1567,N_1504);
nor U2044 (N_2044,N_1948,N_1634);
and U2045 (N_2045,N_1574,N_1827);
nand U2046 (N_2046,N_1616,N_1906);
nor U2047 (N_2047,N_1794,N_1800);
nand U2048 (N_2048,N_1625,N_1707);
or U2049 (N_2049,N_1575,N_1584);
xnor U2050 (N_2050,N_1674,N_1890);
nor U2051 (N_2051,N_1801,N_1779);
xnor U2052 (N_2052,N_1926,N_1626);
nand U2053 (N_2053,N_1615,N_1870);
xor U2054 (N_2054,N_1865,N_1774);
xor U2055 (N_2055,N_1813,N_1836);
nor U2056 (N_2056,N_1638,N_1738);
nor U2057 (N_2057,N_1592,N_1569);
or U2058 (N_2058,N_1548,N_1802);
or U2059 (N_2059,N_1784,N_1931);
xnor U2060 (N_2060,N_1519,N_1793);
nor U2061 (N_2061,N_1792,N_1904);
or U2062 (N_2062,N_1619,N_1663);
and U2063 (N_2063,N_1609,N_1975);
nor U2064 (N_2064,N_1798,N_1532);
nand U2065 (N_2065,N_1854,N_1922);
nand U2066 (N_2066,N_1503,N_1696);
xor U2067 (N_2067,N_1705,N_1679);
or U2068 (N_2068,N_1658,N_1896);
nand U2069 (N_2069,N_1842,N_1633);
xor U2070 (N_2070,N_1848,N_1563);
nand U2071 (N_2071,N_1956,N_1509);
nand U2072 (N_2072,N_1750,N_1666);
and U2073 (N_2073,N_1991,N_1690);
nor U2074 (N_2074,N_1866,N_1919);
nand U2075 (N_2075,N_1530,N_1820);
nand U2076 (N_2076,N_1748,N_1954);
nor U2077 (N_2077,N_1976,N_1987);
nand U2078 (N_2078,N_1889,N_1698);
nand U2079 (N_2079,N_1984,N_1576);
nand U2080 (N_2080,N_1783,N_1734);
xor U2081 (N_2081,N_1701,N_1729);
or U2082 (N_2082,N_1949,N_1564);
and U2083 (N_2083,N_1808,N_1868);
or U2084 (N_2084,N_1601,N_1999);
nand U2085 (N_2085,N_1877,N_1901);
xnor U2086 (N_2086,N_1883,N_1659);
or U2087 (N_2087,N_1557,N_1796);
or U2088 (N_2088,N_1879,N_1521);
nor U2089 (N_2089,N_1858,N_1819);
xor U2090 (N_2090,N_1882,N_1640);
xnor U2091 (N_2091,N_1535,N_1852);
nor U2092 (N_2092,N_1531,N_1699);
nand U2093 (N_2093,N_1550,N_1989);
nand U2094 (N_2094,N_1718,N_1822);
and U2095 (N_2095,N_1539,N_1799);
or U2096 (N_2096,N_1892,N_1715);
nand U2097 (N_2097,N_1874,N_1591);
nor U2098 (N_2098,N_1953,N_1873);
nand U2099 (N_2099,N_1670,N_1544);
nor U2100 (N_2100,N_1758,N_1627);
xnor U2101 (N_2101,N_1712,N_1689);
or U2102 (N_2102,N_1675,N_1809);
nor U2103 (N_2103,N_1523,N_1711);
and U2104 (N_2104,N_1747,N_1673);
or U2105 (N_2105,N_1568,N_1920);
and U2106 (N_2106,N_1856,N_1762);
or U2107 (N_2107,N_1862,N_1934);
nand U2108 (N_2108,N_1655,N_1528);
nor U2109 (N_2109,N_1846,N_1586);
nand U2110 (N_2110,N_1565,N_1894);
nor U2111 (N_2111,N_1912,N_1691);
or U2112 (N_2112,N_1958,N_1853);
and U2113 (N_2113,N_1502,N_1996);
nor U2114 (N_2114,N_1706,N_1915);
or U2115 (N_2115,N_1583,N_1646);
nand U2116 (N_2116,N_1988,N_1553);
or U2117 (N_2117,N_1622,N_1500);
xnor U2118 (N_2118,N_1772,N_1598);
and U2119 (N_2119,N_1769,N_1517);
and U2120 (N_2120,N_1533,N_1631);
nor U2121 (N_2121,N_1613,N_1888);
xnor U2122 (N_2122,N_1639,N_1516);
xnor U2123 (N_2123,N_1787,N_1993);
and U2124 (N_2124,N_1597,N_1744);
xor U2125 (N_2125,N_1562,N_1749);
xor U2126 (N_2126,N_1884,N_1962);
nand U2127 (N_2127,N_1982,N_1643);
or U2128 (N_2128,N_1936,N_1717);
nand U2129 (N_2129,N_1570,N_1703);
or U2130 (N_2130,N_1981,N_1505);
and U2131 (N_2131,N_1942,N_1736);
xor U2132 (N_2132,N_1719,N_1861);
and U2133 (N_2133,N_1961,N_1925);
or U2134 (N_2134,N_1682,N_1540);
and U2135 (N_2135,N_1688,N_1695);
nand U2136 (N_2136,N_1585,N_1881);
nor U2137 (N_2137,N_1891,N_1733);
and U2138 (N_2138,N_1660,N_1606);
nand U2139 (N_2139,N_1864,N_1692);
or U2140 (N_2140,N_1581,N_1551);
nand U2141 (N_2141,N_1914,N_1526);
xnor U2142 (N_2142,N_1946,N_1590);
or U2143 (N_2143,N_1522,N_1875);
nand U2144 (N_2144,N_1721,N_1795);
xor U2145 (N_2145,N_1940,N_1572);
nor U2146 (N_2146,N_1720,N_1555);
or U2147 (N_2147,N_1979,N_1778);
and U2148 (N_2148,N_1806,N_1652);
nor U2149 (N_2149,N_1525,N_1900);
or U2150 (N_2150,N_1947,N_1895);
xor U2151 (N_2151,N_1939,N_1911);
nor U2152 (N_2152,N_1898,N_1651);
nand U2153 (N_2153,N_1742,N_1945);
nor U2154 (N_2154,N_1527,N_1757);
and U2155 (N_2155,N_1935,N_1899);
xnor U2156 (N_2156,N_1785,N_1589);
or U2157 (N_2157,N_1620,N_1880);
nor U2158 (N_2158,N_1629,N_1863);
xnor U2159 (N_2159,N_1855,N_1671);
and U2160 (N_2160,N_1737,N_1661);
xnor U2161 (N_2161,N_1578,N_1944);
or U2162 (N_2162,N_1985,N_1594);
nand U2163 (N_2163,N_1746,N_1872);
nand U2164 (N_2164,N_1788,N_1759);
or U2165 (N_2165,N_1951,N_1905);
xor U2166 (N_2166,N_1978,N_1876);
nor U2167 (N_2167,N_1782,N_1554);
nand U2168 (N_2168,N_1669,N_1990);
xnor U2169 (N_2169,N_1513,N_1818);
or U2170 (N_2170,N_1645,N_1752);
xnor U2171 (N_2171,N_1928,N_1681);
nor U2172 (N_2172,N_1930,N_1790);
xnor U2173 (N_2173,N_1650,N_1963);
xnor U2174 (N_2174,N_1959,N_1684);
and U2175 (N_2175,N_1686,N_1938);
xor U2176 (N_2176,N_1867,N_1869);
xor U2177 (N_2177,N_1965,N_1839);
and U2178 (N_2178,N_1602,N_1667);
nand U2179 (N_2179,N_1743,N_1537);
nor U2180 (N_2180,N_1834,N_1971);
and U2181 (N_2181,N_1507,N_1560);
nor U2182 (N_2182,N_1741,N_1644);
and U2183 (N_2183,N_1677,N_1672);
xor U2184 (N_2184,N_1921,N_1897);
xnor U2185 (N_2185,N_1731,N_1511);
nor U2186 (N_2186,N_1828,N_1538);
nand U2187 (N_2187,N_1600,N_1685);
or U2188 (N_2188,N_1943,N_1835);
xnor U2189 (N_2189,N_1763,N_1764);
xnor U2190 (N_2190,N_1824,N_1871);
nor U2191 (N_2191,N_1559,N_1501);
xnor U2192 (N_2192,N_1833,N_1515);
xnor U2193 (N_2193,N_1767,N_1710);
nor U2194 (N_2194,N_1766,N_1923);
nand U2195 (N_2195,N_1927,N_1776);
xor U2196 (N_2196,N_1730,N_1780);
and U2197 (N_2197,N_1887,N_1924);
xnor U2198 (N_2198,N_1916,N_1753);
and U2199 (N_2199,N_1811,N_1621);
and U2200 (N_2200,N_1665,N_1649);
xnor U2201 (N_2201,N_1786,N_1844);
or U2202 (N_2202,N_1847,N_1524);
or U2203 (N_2203,N_1588,N_1885);
xnor U2204 (N_2204,N_1817,N_1641);
nand U2205 (N_2205,N_1536,N_1740);
xor U2206 (N_2206,N_1648,N_1726);
xor U2207 (N_2207,N_1825,N_1727);
nor U2208 (N_2208,N_1812,N_1664);
or U2209 (N_2209,N_1814,N_1994);
xnor U2210 (N_2210,N_1797,N_1843);
and U2211 (N_2211,N_1845,N_1632);
nor U2212 (N_2212,N_1739,N_1582);
xor U2213 (N_2213,N_1546,N_1610);
nor U2214 (N_2214,N_1995,N_1552);
or U2215 (N_2215,N_1603,N_1566);
nand U2216 (N_2216,N_1732,N_1668);
nand U2217 (N_2217,N_1653,N_1637);
xnor U2218 (N_2218,N_1918,N_1549);
or U2219 (N_2219,N_1754,N_1907);
and U2220 (N_2220,N_1608,N_1508);
or U2221 (N_2221,N_1678,N_1654);
nand U2222 (N_2222,N_1917,N_1709);
xnor U2223 (N_2223,N_1810,N_1972);
xor U2224 (N_2224,N_1968,N_1611);
nand U2225 (N_2225,N_1826,N_1980);
nor U2226 (N_2226,N_1937,N_1683);
nor U2227 (N_2227,N_1614,N_1902);
nand U2228 (N_2228,N_1604,N_1941);
nand U2229 (N_2229,N_1662,N_1966);
nor U2230 (N_2230,N_1541,N_1607);
nand U2231 (N_2231,N_1512,N_1687);
xor U2232 (N_2232,N_1510,N_1630);
xnor U2233 (N_2233,N_1992,N_1636);
nor U2234 (N_2234,N_1955,N_1933);
and U2235 (N_2235,N_1831,N_1735);
and U2236 (N_2236,N_1791,N_1713);
nor U2237 (N_2237,N_1605,N_1816);
or U2238 (N_2238,N_1859,N_1760);
nand U2239 (N_2239,N_1805,N_1599);
nor U2240 (N_2240,N_1765,N_1571);
nor U2241 (N_2241,N_1973,N_1543);
or U2242 (N_2242,N_1618,N_1878);
nor U2243 (N_2243,N_1693,N_1556);
and U2244 (N_2244,N_1768,N_1700);
or U2245 (N_2245,N_1903,N_1969);
nand U2246 (N_2246,N_1694,N_1960);
and U2247 (N_2247,N_1547,N_1593);
or U2248 (N_2248,N_1534,N_1506);
or U2249 (N_2249,N_1529,N_1579);
nor U2250 (N_2250,N_1712,N_1898);
and U2251 (N_2251,N_1824,N_1555);
nand U2252 (N_2252,N_1541,N_1724);
and U2253 (N_2253,N_1768,N_1522);
nor U2254 (N_2254,N_1726,N_1710);
or U2255 (N_2255,N_1590,N_1746);
nor U2256 (N_2256,N_1881,N_1942);
or U2257 (N_2257,N_1540,N_1788);
and U2258 (N_2258,N_1708,N_1988);
xnor U2259 (N_2259,N_1509,N_1819);
xnor U2260 (N_2260,N_1862,N_1894);
xor U2261 (N_2261,N_1820,N_1753);
xnor U2262 (N_2262,N_1819,N_1560);
xnor U2263 (N_2263,N_1994,N_1686);
nor U2264 (N_2264,N_1865,N_1952);
nor U2265 (N_2265,N_1641,N_1999);
nand U2266 (N_2266,N_1612,N_1803);
nor U2267 (N_2267,N_1643,N_1564);
and U2268 (N_2268,N_1695,N_1592);
nand U2269 (N_2269,N_1562,N_1993);
nor U2270 (N_2270,N_1731,N_1762);
xnor U2271 (N_2271,N_1779,N_1873);
and U2272 (N_2272,N_1823,N_1614);
nand U2273 (N_2273,N_1864,N_1881);
xor U2274 (N_2274,N_1617,N_1651);
xor U2275 (N_2275,N_1846,N_1908);
and U2276 (N_2276,N_1555,N_1915);
nand U2277 (N_2277,N_1796,N_1688);
and U2278 (N_2278,N_1542,N_1774);
nand U2279 (N_2279,N_1531,N_1757);
xor U2280 (N_2280,N_1645,N_1678);
nand U2281 (N_2281,N_1544,N_1827);
and U2282 (N_2282,N_1633,N_1517);
xor U2283 (N_2283,N_1762,N_1626);
nand U2284 (N_2284,N_1751,N_1514);
and U2285 (N_2285,N_1779,N_1805);
nand U2286 (N_2286,N_1810,N_1548);
nand U2287 (N_2287,N_1516,N_1514);
xnor U2288 (N_2288,N_1500,N_1813);
nor U2289 (N_2289,N_1597,N_1829);
xor U2290 (N_2290,N_1705,N_1672);
nor U2291 (N_2291,N_1723,N_1600);
nor U2292 (N_2292,N_1810,N_1989);
nand U2293 (N_2293,N_1765,N_1981);
or U2294 (N_2294,N_1536,N_1785);
nor U2295 (N_2295,N_1909,N_1860);
or U2296 (N_2296,N_1607,N_1650);
nand U2297 (N_2297,N_1744,N_1731);
and U2298 (N_2298,N_1716,N_1667);
or U2299 (N_2299,N_1517,N_1618);
nand U2300 (N_2300,N_1917,N_1904);
nand U2301 (N_2301,N_1917,N_1521);
nor U2302 (N_2302,N_1598,N_1569);
and U2303 (N_2303,N_1747,N_1664);
or U2304 (N_2304,N_1804,N_1764);
xor U2305 (N_2305,N_1574,N_1813);
xor U2306 (N_2306,N_1749,N_1910);
and U2307 (N_2307,N_1785,N_1755);
nor U2308 (N_2308,N_1704,N_1567);
nand U2309 (N_2309,N_1831,N_1895);
nor U2310 (N_2310,N_1913,N_1952);
nor U2311 (N_2311,N_1735,N_1817);
nor U2312 (N_2312,N_1726,N_1777);
nor U2313 (N_2313,N_1722,N_1993);
and U2314 (N_2314,N_1956,N_1676);
xor U2315 (N_2315,N_1648,N_1871);
or U2316 (N_2316,N_1799,N_1579);
xor U2317 (N_2317,N_1720,N_1523);
nand U2318 (N_2318,N_1883,N_1979);
or U2319 (N_2319,N_1770,N_1850);
nor U2320 (N_2320,N_1704,N_1622);
xor U2321 (N_2321,N_1634,N_1827);
or U2322 (N_2322,N_1676,N_1777);
or U2323 (N_2323,N_1852,N_1993);
or U2324 (N_2324,N_1719,N_1808);
nand U2325 (N_2325,N_1733,N_1516);
xor U2326 (N_2326,N_1753,N_1957);
nor U2327 (N_2327,N_1727,N_1657);
or U2328 (N_2328,N_1630,N_1662);
and U2329 (N_2329,N_1705,N_1624);
xor U2330 (N_2330,N_1611,N_1842);
or U2331 (N_2331,N_1983,N_1878);
nor U2332 (N_2332,N_1602,N_1579);
or U2333 (N_2333,N_1572,N_1962);
nand U2334 (N_2334,N_1725,N_1888);
xnor U2335 (N_2335,N_1969,N_1782);
or U2336 (N_2336,N_1587,N_1776);
nor U2337 (N_2337,N_1657,N_1894);
nor U2338 (N_2338,N_1524,N_1501);
xnor U2339 (N_2339,N_1952,N_1670);
nor U2340 (N_2340,N_1515,N_1705);
or U2341 (N_2341,N_1637,N_1607);
nand U2342 (N_2342,N_1631,N_1980);
or U2343 (N_2343,N_1623,N_1596);
xor U2344 (N_2344,N_1988,N_1501);
and U2345 (N_2345,N_1693,N_1573);
and U2346 (N_2346,N_1618,N_1637);
nand U2347 (N_2347,N_1994,N_1685);
or U2348 (N_2348,N_1633,N_1630);
nand U2349 (N_2349,N_1699,N_1799);
nand U2350 (N_2350,N_1879,N_1596);
or U2351 (N_2351,N_1805,N_1864);
or U2352 (N_2352,N_1607,N_1635);
nand U2353 (N_2353,N_1568,N_1865);
xnor U2354 (N_2354,N_1698,N_1901);
and U2355 (N_2355,N_1692,N_1695);
or U2356 (N_2356,N_1590,N_1685);
nand U2357 (N_2357,N_1880,N_1662);
xor U2358 (N_2358,N_1835,N_1692);
nor U2359 (N_2359,N_1809,N_1899);
or U2360 (N_2360,N_1527,N_1917);
nand U2361 (N_2361,N_1535,N_1761);
xor U2362 (N_2362,N_1692,N_1654);
xor U2363 (N_2363,N_1881,N_1934);
and U2364 (N_2364,N_1520,N_1762);
xnor U2365 (N_2365,N_1913,N_1542);
nor U2366 (N_2366,N_1531,N_1979);
xor U2367 (N_2367,N_1508,N_1683);
and U2368 (N_2368,N_1746,N_1812);
xor U2369 (N_2369,N_1787,N_1837);
nor U2370 (N_2370,N_1784,N_1744);
xor U2371 (N_2371,N_1535,N_1554);
nand U2372 (N_2372,N_1988,N_1717);
and U2373 (N_2373,N_1743,N_1882);
nor U2374 (N_2374,N_1552,N_1919);
or U2375 (N_2375,N_1770,N_1686);
or U2376 (N_2376,N_1995,N_1795);
or U2377 (N_2377,N_1721,N_1903);
and U2378 (N_2378,N_1949,N_1527);
xnor U2379 (N_2379,N_1866,N_1678);
or U2380 (N_2380,N_1913,N_1837);
nor U2381 (N_2381,N_1819,N_1730);
xnor U2382 (N_2382,N_1832,N_1632);
xnor U2383 (N_2383,N_1711,N_1823);
nor U2384 (N_2384,N_1793,N_1596);
and U2385 (N_2385,N_1913,N_1513);
nor U2386 (N_2386,N_1907,N_1518);
and U2387 (N_2387,N_1770,N_1902);
nor U2388 (N_2388,N_1841,N_1781);
and U2389 (N_2389,N_1985,N_1539);
nand U2390 (N_2390,N_1599,N_1938);
nor U2391 (N_2391,N_1919,N_1557);
nor U2392 (N_2392,N_1837,N_1792);
or U2393 (N_2393,N_1812,N_1501);
or U2394 (N_2394,N_1755,N_1770);
nor U2395 (N_2395,N_1590,N_1692);
nand U2396 (N_2396,N_1571,N_1619);
and U2397 (N_2397,N_1676,N_1563);
xor U2398 (N_2398,N_1906,N_1843);
nand U2399 (N_2399,N_1703,N_1606);
and U2400 (N_2400,N_1518,N_1533);
xor U2401 (N_2401,N_1625,N_1649);
xor U2402 (N_2402,N_1856,N_1563);
nor U2403 (N_2403,N_1905,N_1638);
nand U2404 (N_2404,N_1946,N_1944);
nor U2405 (N_2405,N_1953,N_1570);
nand U2406 (N_2406,N_1894,N_1948);
or U2407 (N_2407,N_1875,N_1960);
and U2408 (N_2408,N_1762,N_1938);
nand U2409 (N_2409,N_1900,N_1773);
nand U2410 (N_2410,N_1592,N_1637);
xor U2411 (N_2411,N_1556,N_1632);
nand U2412 (N_2412,N_1719,N_1918);
and U2413 (N_2413,N_1573,N_1526);
or U2414 (N_2414,N_1704,N_1869);
nand U2415 (N_2415,N_1865,N_1586);
nor U2416 (N_2416,N_1616,N_1796);
nor U2417 (N_2417,N_1784,N_1634);
nand U2418 (N_2418,N_1999,N_1794);
nor U2419 (N_2419,N_1878,N_1680);
nand U2420 (N_2420,N_1990,N_1795);
or U2421 (N_2421,N_1993,N_1678);
xor U2422 (N_2422,N_1916,N_1640);
nor U2423 (N_2423,N_1554,N_1839);
xor U2424 (N_2424,N_1558,N_1861);
xnor U2425 (N_2425,N_1736,N_1518);
nand U2426 (N_2426,N_1851,N_1930);
and U2427 (N_2427,N_1526,N_1768);
nor U2428 (N_2428,N_1501,N_1526);
xor U2429 (N_2429,N_1568,N_1759);
and U2430 (N_2430,N_1902,N_1906);
or U2431 (N_2431,N_1518,N_1589);
nor U2432 (N_2432,N_1898,N_1920);
and U2433 (N_2433,N_1972,N_1733);
or U2434 (N_2434,N_1981,N_1599);
or U2435 (N_2435,N_1656,N_1561);
nand U2436 (N_2436,N_1693,N_1976);
xnor U2437 (N_2437,N_1851,N_1769);
and U2438 (N_2438,N_1764,N_1705);
xor U2439 (N_2439,N_1911,N_1913);
nand U2440 (N_2440,N_1714,N_1575);
nand U2441 (N_2441,N_1862,N_1982);
or U2442 (N_2442,N_1993,N_1614);
nor U2443 (N_2443,N_1561,N_1515);
nand U2444 (N_2444,N_1908,N_1792);
or U2445 (N_2445,N_1741,N_1653);
and U2446 (N_2446,N_1802,N_1540);
nand U2447 (N_2447,N_1800,N_1577);
nor U2448 (N_2448,N_1701,N_1984);
nand U2449 (N_2449,N_1806,N_1993);
or U2450 (N_2450,N_1600,N_1541);
and U2451 (N_2451,N_1600,N_1845);
nor U2452 (N_2452,N_1648,N_1579);
nand U2453 (N_2453,N_1732,N_1859);
nor U2454 (N_2454,N_1524,N_1809);
xnor U2455 (N_2455,N_1676,N_1688);
nand U2456 (N_2456,N_1641,N_1542);
nor U2457 (N_2457,N_1796,N_1772);
and U2458 (N_2458,N_1956,N_1677);
nor U2459 (N_2459,N_1909,N_1555);
or U2460 (N_2460,N_1546,N_1551);
xor U2461 (N_2461,N_1503,N_1510);
nand U2462 (N_2462,N_1845,N_1995);
or U2463 (N_2463,N_1606,N_1537);
and U2464 (N_2464,N_1665,N_1593);
nand U2465 (N_2465,N_1920,N_1556);
xnor U2466 (N_2466,N_1815,N_1840);
or U2467 (N_2467,N_1741,N_1951);
nor U2468 (N_2468,N_1542,N_1974);
xnor U2469 (N_2469,N_1689,N_1551);
or U2470 (N_2470,N_1689,N_1703);
and U2471 (N_2471,N_1904,N_1901);
nand U2472 (N_2472,N_1692,N_1702);
or U2473 (N_2473,N_1958,N_1760);
nand U2474 (N_2474,N_1667,N_1660);
nand U2475 (N_2475,N_1870,N_1969);
or U2476 (N_2476,N_1963,N_1562);
and U2477 (N_2477,N_1615,N_1926);
nor U2478 (N_2478,N_1998,N_1626);
nand U2479 (N_2479,N_1613,N_1505);
nor U2480 (N_2480,N_1942,N_1869);
xnor U2481 (N_2481,N_1800,N_1842);
xor U2482 (N_2482,N_1780,N_1721);
nand U2483 (N_2483,N_1884,N_1823);
xor U2484 (N_2484,N_1568,N_1990);
nor U2485 (N_2485,N_1576,N_1629);
nor U2486 (N_2486,N_1773,N_1945);
and U2487 (N_2487,N_1895,N_1817);
xor U2488 (N_2488,N_1950,N_1506);
nand U2489 (N_2489,N_1675,N_1980);
nand U2490 (N_2490,N_1760,N_1960);
nand U2491 (N_2491,N_1670,N_1876);
xnor U2492 (N_2492,N_1591,N_1807);
nor U2493 (N_2493,N_1736,N_1878);
nor U2494 (N_2494,N_1524,N_1563);
and U2495 (N_2495,N_1582,N_1829);
and U2496 (N_2496,N_1504,N_1945);
nand U2497 (N_2497,N_1942,N_1788);
nand U2498 (N_2498,N_1848,N_1541);
and U2499 (N_2499,N_1727,N_1685);
or U2500 (N_2500,N_2193,N_2147);
and U2501 (N_2501,N_2338,N_2075);
and U2502 (N_2502,N_2080,N_2146);
nand U2503 (N_2503,N_2163,N_2391);
nand U2504 (N_2504,N_2003,N_2475);
and U2505 (N_2505,N_2089,N_2038);
xnor U2506 (N_2506,N_2417,N_2226);
nor U2507 (N_2507,N_2235,N_2133);
xnor U2508 (N_2508,N_2271,N_2024);
nand U2509 (N_2509,N_2433,N_2451);
xor U2510 (N_2510,N_2355,N_2119);
nand U2511 (N_2511,N_2060,N_2251);
nor U2512 (N_2512,N_2044,N_2374);
nand U2513 (N_2513,N_2078,N_2107);
nor U2514 (N_2514,N_2328,N_2412);
xor U2515 (N_2515,N_2331,N_2394);
nand U2516 (N_2516,N_2437,N_2238);
nand U2517 (N_2517,N_2208,N_2365);
or U2518 (N_2518,N_2117,N_2164);
or U2519 (N_2519,N_2349,N_2291);
nand U2520 (N_2520,N_2076,N_2282);
nand U2521 (N_2521,N_2316,N_2178);
xnor U2522 (N_2522,N_2279,N_2330);
or U2523 (N_2523,N_2401,N_2306);
and U2524 (N_2524,N_2430,N_2145);
xor U2525 (N_2525,N_2113,N_2327);
nor U2526 (N_2526,N_2422,N_2440);
nor U2527 (N_2527,N_2166,N_2028);
nor U2528 (N_2528,N_2065,N_2399);
nand U2529 (N_2529,N_2213,N_2177);
and U2530 (N_2530,N_2441,N_2491);
nand U2531 (N_2531,N_2037,N_2383);
and U2532 (N_2532,N_2258,N_2116);
and U2533 (N_2533,N_2369,N_2049);
nand U2534 (N_2534,N_2175,N_2159);
and U2535 (N_2535,N_2153,N_2325);
and U2536 (N_2536,N_2479,N_2463);
or U2537 (N_2537,N_2449,N_2368);
and U2538 (N_2538,N_2157,N_2406);
nor U2539 (N_2539,N_2442,N_2287);
xnor U2540 (N_2540,N_2446,N_2319);
xor U2541 (N_2541,N_2496,N_2305);
nand U2542 (N_2542,N_2309,N_2444);
or U2543 (N_2543,N_2231,N_2040);
or U2544 (N_2544,N_2455,N_2335);
nor U2545 (N_2545,N_2301,N_2035);
nor U2546 (N_2546,N_2141,N_2372);
nor U2547 (N_2547,N_2280,N_2160);
and U2548 (N_2548,N_2459,N_2105);
and U2549 (N_2549,N_2033,N_2450);
and U2550 (N_2550,N_2064,N_2452);
and U2551 (N_2551,N_2434,N_2248);
nand U2552 (N_2552,N_2244,N_2285);
and U2553 (N_2553,N_2484,N_2268);
or U2554 (N_2554,N_2172,N_2012);
or U2555 (N_2555,N_2314,N_2182);
nand U2556 (N_2556,N_2091,N_2296);
nand U2557 (N_2557,N_2099,N_2181);
nand U2558 (N_2558,N_2067,N_2302);
or U2559 (N_2559,N_2400,N_2135);
or U2560 (N_2560,N_2404,N_2418);
xor U2561 (N_2561,N_2468,N_2015);
nand U2562 (N_2562,N_2056,N_2267);
and U2563 (N_2563,N_2345,N_2266);
or U2564 (N_2564,N_2256,N_2168);
nor U2565 (N_2565,N_2408,N_2167);
and U2566 (N_2566,N_2447,N_2224);
and U2567 (N_2567,N_2197,N_2432);
or U2568 (N_2568,N_2337,N_2252);
xor U2569 (N_2569,N_2209,N_2128);
xor U2570 (N_2570,N_2095,N_2051);
or U2571 (N_2571,N_2201,N_2162);
and U2572 (N_2572,N_2289,N_2478);
and U2573 (N_2573,N_2409,N_2216);
and U2574 (N_2574,N_2386,N_2294);
or U2575 (N_2575,N_2069,N_2087);
nand U2576 (N_2576,N_2101,N_2017);
or U2577 (N_2577,N_2005,N_2428);
and U2578 (N_2578,N_2344,N_2411);
xnor U2579 (N_2579,N_2126,N_2247);
xor U2580 (N_2580,N_2315,N_2169);
xnor U2581 (N_2581,N_2072,N_2390);
nor U2582 (N_2582,N_2388,N_2299);
or U2583 (N_2583,N_2096,N_2023);
xor U2584 (N_2584,N_2058,N_2048);
xor U2585 (N_2585,N_2321,N_2237);
or U2586 (N_2586,N_2403,N_2332);
and U2587 (N_2587,N_2260,N_2363);
or U2588 (N_2588,N_2382,N_2132);
xnor U2589 (N_2589,N_2274,N_2032);
nor U2590 (N_2590,N_2492,N_2151);
nor U2591 (N_2591,N_2234,N_2293);
and U2592 (N_2592,N_2298,N_2174);
and U2593 (N_2593,N_2109,N_2010);
and U2594 (N_2594,N_2240,N_2376);
and U2595 (N_2595,N_2469,N_2002);
xor U2596 (N_2596,N_2407,N_2343);
nand U2597 (N_2597,N_2150,N_2124);
xnor U2598 (N_2598,N_2071,N_2473);
and U2599 (N_2599,N_2053,N_2477);
xnor U2600 (N_2600,N_2094,N_2199);
and U2601 (N_2601,N_2220,N_2125);
or U2602 (N_2602,N_2066,N_2192);
or U2603 (N_2603,N_2140,N_2253);
nor U2604 (N_2604,N_2063,N_2190);
nor U2605 (N_2605,N_2474,N_2004);
and U2606 (N_2606,N_2270,N_2171);
and U2607 (N_2607,N_2022,N_2384);
nor U2608 (N_2608,N_2106,N_2269);
nor U2609 (N_2609,N_2081,N_2367);
xor U2610 (N_2610,N_2018,N_2079);
or U2611 (N_2611,N_2110,N_2215);
or U2612 (N_2612,N_2453,N_2273);
and U2613 (N_2613,N_2308,N_2183);
nand U2614 (N_2614,N_2290,N_2414);
nand U2615 (N_2615,N_2431,N_2427);
or U2616 (N_2616,N_2462,N_2458);
nor U2617 (N_2617,N_2137,N_2499);
nor U2618 (N_2618,N_2131,N_2230);
or U2619 (N_2619,N_2186,N_2217);
nand U2620 (N_2620,N_2052,N_2118);
xor U2621 (N_2621,N_2385,N_2340);
nor U2622 (N_2622,N_2250,N_2445);
xor U2623 (N_2623,N_2472,N_2487);
or U2624 (N_2624,N_2239,N_2439);
nand U2625 (N_2625,N_2136,N_2229);
nor U2626 (N_2626,N_2185,N_2416);
nand U2627 (N_2627,N_2364,N_2413);
or U2628 (N_2628,N_2352,N_2195);
nand U2629 (N_2629,N_2254,N_2262);
xor U2630 (N_2630,N_2465,N_2225);
and U2631 (N_2631,N_2377,N_2456);
nor U2632 (N_2632,N_2104,N_2351);
nor U2633 (N_2633,N_2149,N_2467);
or U2634 (N_2634,N_2156,N_2127);
nand U2635 (N_2635,N_2210,N_2361);
or U2636 (N_2636,N_2233,N_2317);
nand U2637 (N_2637,N_2341,N_2189);
or U2638 (N_2638,N_2265,N_2144);
and U2639 (N_2639,N_2421,N_2281);
nor U2640 (N_2640,N_2191,N_2042);
nor U2641 (N_2641,N_2366,N_2333);
and U2642 (N_2642,N_2152,N_2312);
nor U2643 (N_2643,N_2054,N_2389);
or U2644 (N_2644,N_2026,N_2470);
or U2645 (N_2645,N_2373,N_2143);
or U2646 (N_2646,N_2495,N_2221);
nand U2647 (N_2647,N_2086,N_2165);
nor U2648 (N_2648,N_2203,N_2129);
nor U2649 (N_2649,N_2227,N_2405);
xnor U2650 (N_2650,N_2120,N_2448);
xor U2651 (N_2651,N_2288,N_2395);
or U2652 (N_2652,N_2139,N_2357);
or U2653 (N_2653,N_2311,N_2329);
and U2654 (N_2654,N_2030,N_2180);
or U2655 (N_2655,N_2381,N_2050);
and U2656 (N_2656,N_2438,N_2284);
nor U2657 (N_2657,N_2036,N_2222);
and U2658 (N_2658,N_2255,N_2276);
nand U2659 (N_2659,N_2092,N_2425);
and U2660 (N_2660,N_2241,N_2059);
nand U2661 (N_2661,N_2008,N_2375);
and U2662 (N_2662,N_2300,N_2490);
nand U2663 (N_2663,N_2236,N_2443);
or U2664 (N_2664,N_2188,N_2007);
nand U2665 (N_2665,N_2457,N_2326);
and U2666 (N_2666,N_2039,N_2387);
or U2667 (N_2667,N_2034,N_2098);
and U2668 (N_2668,N_2077,N_2393);
nand U2669 (N_2669,N_2336,N_2114);
or U2670 (N_2670,N_2275,N_2093);
xnor U2671 (N_2671,N_2423,N_2379);
or U2672 (N_2672,N_2354,N_2173);
xor U2673 (N_2673,N_2295,N_2378);
xor U2674 (N_2674,N_2424,N_2031);
nand U2675 (N_2675,N_2426,N_2027);
nor U2676 (N_2676,N_2283,N_2212);
and U2677 (N_2677,N_2214,N_2481);
or U2678 (N_2678,N_2057,N_2420);
and U2679 (N_2679,N_2380,N_2161);
and U2680 (N_2680,N_2346,N_2097);
nor U2681 (N_2681,N_2303,N_2219);
nand U2682 (N_2682,N_2277,N_2055);
xnor U2683 (N_2683,N_2198,N_2324);
and U2684 (N_2684,N_2045,N_2006);
nand U2685 (N_2685,N_2461,N_2370);
nand U2686 (N_2686,N_2242,N_2435);
nand U2687 (N_2687,N_2176,N_2476);
xor U2688 (N_2688,N_2011,N_2187);
nand U2689 (N_2689,N_2029,N_2232);
nand U2690 (N_2690,N_2115,N_2158);
xor U2691 (N_2691,N_2206,N_2202);
and U2692 (N_2692,N_2436,N_2360);
nor U2693 (N_2693,N_2154,N_2488);
nor U2694 (N_2694,N_2342,N_2392);
xnor U2695 (N_2695,N_2471,N_2323);
xor U2696 (N_2696,N_2334,N_2429);
nand U2697 (N_2697,N_2419,N_2320);
and U2698 (N_2698,N_2085,N_2243);
xor U2699 (N_2699,N_2350,N_2371);
xnor U2700 (N_2700,N_2070,N_2396);
nor U2701 (N_2701,N_2398,N_2259);
nand U2702 (N_2702,N_2196,N_2402);
xor U2703 (N_2703,N_2073,N_2041);
nand U2704 (N_2704,N_2486,N_2123);
nand U2705 (N_2705,N_2090,N_2194);
nand U2706 (N_2706,N_2348,N_2061);
nor U2707 (N_2707,N_2264,N_2020);
or U2708 (N_2708,N_2088,N_2043);
nor U2709 (N_2709,N_2102,N_2211);
xor U2710 (N_2710,N_2019,N_2485);
xnor U2711 (N_2711,N_2494,N_2155);
nor U2712 (N_2712,N_2480,N_2359);
or U2713 (N_2713,N_2497,N_2410);
xnor U2714 (N_2714,N_2246,N_2228);
xnor U2715 (N_2715,N_2310,N_2257);
and U2716 (N_2716,N_2205,N_2130);
or U2717 (N_2717,N_2014,N_2103);
or U2718 (N_2718,N_2074,N_2307);
nand U2719 (N_2719,N_2218,N_2313);
xor U2720 (N_2720,N_2272,N_2112);
or U2721 (N_2721,N_2356,N_2084);
nand U2722 (N_2722,N_2466,N_2184);
and U2723 (N_2723,N_2122,N_2142);
xor U2724 (N_2724,N_2000,N_2362);
or U2725 (N_2725,N_2062,N_2397);
nor U2726 (N_2726,N_2498,N_2318);
and U2727 (N_2727,N_2068,N_2249);
nor U2728 (N_2728,N_2100,N_2223);
and U2729 (N_2729,N_2415,N_2482);
xnor U2730 (N_2730,N_2489,N_2046);
nor U2731 (N_2731,N_2358,N_2286);
nand U2732 (N_2732,N_2001,N_2460);
xor U2733 (N_2733,N_2111,N_2322);
nand U2734 (N_2734,N_2047,N_2134);
nor U2735 (N_2735,N_2025,N_2464);
xor U2736 (N_2736,N_2016,N_2454);
nand U2737 (N_2737,N_2148,N_2138);
nor U2738 (N_2738,N_2021,N_2082);
and U2739 (N_2739,N_2493,N_2292);
xor U2740 (N_2740,N_2339,N_2009);
or U2741 (N_2741,N_2179,N_2483);
nor U2742 (N_2742,N_2170,N_2304);
or U2743 (N_2743,N_2121,N_2083);
nor U2744 (N_2744,N_2347,N_2278);
and U2745 (N_2745,N_2200,N_2297);
or U2746 (N_2746,N_2263,N_2013);
and U2747 (N_2747,N_2245,N_2207);
nand U2748 (N_2748,N_2353,N_2261);
xnor U2749 (N_2749,N_2204,N_2108);
nand U2750 (N_2750,N_2284,N_2459);
xor U2751 (N_2751,N_2160,N_2194);
nor U2752 (N_2752,N_2105,N_2059);
or U2753 (N_2753,N_2460,N_2080);
nor U2754 (N_2754,N_2216,N_2038);
and U2755 (N_2755,N_2438,N_2104);
xnor U2756 (N_2756,N_2419,N_2295);
or U2757 (N_2757,N_2265,N_2287);
xor U2758 (N_2758,N_2070,N_2287);
nand U2759 (N_2759,N_2199,N_2323);
and U2760 (N_2760,N_2115,N_2059);
nand U2761 (N_2761,N_2332,N_2232);
nor U2762 (N_2762,N_2256,N_2336);
nand U2763 (N_2763,N_2325,N_2011);
or U2764 (N_2764,N_2416,N_2114);
and U2765 (N_2765,N_2363,N_2353);
nor U2766 (N_2766,N_2239,N_2005);
and U2767 (N_2767,N_2016,N_2161);
nand U2768 (N_2768,N_2484,N_2408);
or U2769 (N_2769,N_2274,N_2174);
and U2770 (N_2770,N_2082,N_2054);
and U2771 (N_2771,N_2388,N_2305);
or U2772 (N_2772,N_2350,N_2323);
nand U2773 (N_2773,N_2092,N_2241);
nor U2774 (N_2774,N_2087,N_2056);
nor U2775 (N_2775,N_2117,N_2183);
or U2776 (N_2776,N_2449,N_2270);
or U2777 (N_2777,N_2218,N_2454);
xnor U2778 (N_2778,N_2481,N_2194);
and U2779 (N_2779,N_2213,N_2493);
nor U2780 (N_2780,N_2224,N_2129);
and U2781 (N_2781,N_2294,N_2447);
nor U2782 (N_2782,N_2439,N_2417);
and U2783 (N_2783,N_2415,N_2131);
nand U2784 (N_2784,N_2368,N_2429);
nor U2785 (N_2785,N_2146,N_2101);
xor U2786 (N_2786,N_2133,N_2456);
and U2787 (N_2787,N_2221,N_2326);
and U2788 (N_2788,N_2168,N_2381);
and U2789 (N_2789,N_2216,N_2032);
or U2790 (N_2790,N_2131,N_2099);
nor U2791 (N_2791,N_2046,N_2091);
xnor U2792 (N_2792,N_2486,N_2194);
xor U2793 (N_2793,N_2007,N_2216);
and U2794 (N_2794,N_2253,N_2259);
xnor U2795 (N_2795,N_2014,N_2052);
xnor U2796 (N_2796,N_2187,N_2299);
xor U2797 (N_2797,N_2469,N_2158);
xnor U2798 (N_2798,N_2286,N_2213);
xnor U2799 (N_2799,N_2095,N_2338);
and U2800 (N_2800,N_2058,N_2042);
nor U2801 (N_2801,N_2130,N_2227);
xor U2802 (N_2802,N_2480,N_2244);
nor U2803 (N_2803,N_2349,N_2214);
and U2804 (N_2804,N_2118,N_2462);
and U2805 (N_2805,N_2222,N_2236);
nor U2806 (N_2806,N_2410,N_2452);
xnor U2807 (N_2807,N_2196,N_2052);
nor U2808 (N_2808,N_2479,N_2122);
and U2809 (N_2809,N_2048,N_2316);
or U2810 (N_2810,N_2173,N_2373);
xor U2811 (N_2811,N_2359,N_2033);
or U2812 (N_2812,N_2014,N_2371);
or U2813 (N_2813,N_2147,N_2288);
or U2814 (N_2814,N_2217,N_2057);
nor U2815 (N_2815,N_2270,N_2306);
or U2816 (N_2816,N_2246,N_2053);
or U2817 (N_2817,N_2419,N_2480);
nand U2818 (N_2818,N_2490,N_2332);
nand U2819 (N_2819,N_2497,N_2279);
xor U2820 (N_2820,N_2117,N_2111);
and U2821 (N_2821,N_2444,N_2453);
or U2822 (N_2822,N_2246,N_2304);
nand U2823 (N_2823,N_2271,N_2407);
xor U2824 (N_2824,N_2228,N_2368);
or U2825 (N_2825,N_2126,N_2429);
and U2826 (N_2826,N_2194,N_2231);
or U2827 (N_2827,N_2095,N_2433);
and U2828 (N_2828,N_2383,N_2350);
and U2829 (N_2829,N_2455,N_2215);
or U2830 (N_2830,N_2265,N_2269);
xor U2831 (N_2831,N_2442,N_2170);
and U2832 (N_2832,N_2062,N_2326);
nor U2833 (N_2833,N_2356,N_2383);
or U2834 (N_2834,N_2406,N_2334);
and U2835 (N_2835,N_2304,N_2124);
xnor U2836 (N_2836,N_2214,N_2220);
and U2837 (N_2837,N_2255,N_2291);
or U2838 (N_2838,N_2043,N_2473);
nor U2839 (N_2839,N_2175,N_2408);
xnor U2840 (N_2840,N_2158,N_2330);
xnor U2841 (N_2841,N_2488,N_2460);
or U2842 (N_2842,N_2260,N_2321);
nand U2843 (N_2843,N_2274,N_2178);
nor U2844 (N_2844,N_2270,N_2123);
xnor U2845 (N_2845,N_2148,N_2111);
or U2846 (N_2846,N_2492,N_2052);
xnor U2847 (N_2847,N_2212,N_2289);
nor U2848 (N_2848,N_2056,N_2471);
xnor U2849 (N_2849,N_2479,N_2274);
nand U2850 (N_2850,N_2045,N_2019);
or U2851 (N_2851,N_2268,N_2192);
xor U2852 (N_2852,N_2151,N_2001);
nand U2853 (N_2853,N_2296,N_2343);
nand U2854 (N_2854,N_2177,N_2498);
nand U2855 (N_2855,N_2126,N_2402);
and U2856 (N_2856,N_2132,N_2241);
and U2857 (N_2857,N_2457,N_2233);
nand U2858 (N_2858,N_2029,N_2138);
nor U2859 (N_2859,N_2302,N_2339);
or U2860 (N_2860,N_2163,N_2051);
nand U2861 (N_2861,N_2248,N_2477);
or U2862 (N_2862,N_2417,N_2173);
or U2863 (N_2863,N_2277,N_2256);
nand U2864 (N_2864,N_2262,N_2275);
xor U2865 (N_2865,N_2006,N_2034);
and U2866 (N_2866,N_2153,N_2392);
nand U2867 (N_2867,N_2094,N_2219);
nor U2868 (N_2868,N_2065,N_2108);
xor U2869 (N_2869,N_2013,N_2068);
nor U2870 (N_2870,N_2497,N_2176);
xnor U2871 (N_2871,N_2346,N_2251);
nor U2872 (N_2872,N_2047,N_2116);
and U2873 (N_2873,N_2012,N_2372);
or U2874 (N_2874,N_2076,N_2148);
or U2875 (N_2875,N_2363,N_2379);
xnor U2876 (N_2876,N_2415,N_2232);
xor U2877 (N_2877,N_2418,N_2364);
nand U2878 (N_2878,N_2298,N_2321);
nand U2879 (N_2879,N_2060,N_2225);
or U2880 (N_2880,N_2388,N_2479);
and U2881 (N_2881,N_2065,N_2097);
and U2882 (N_2882,N_2424,N_2258);
nor U2883 (N_2883,N_2364,N_2080);
or U2884 (N_2884,N_2198,N_2441);
and U2885 (N_2885,N_2438,N_2332);
and U2886 (N_2886,N_2049,N_2429);
and U2887 (N_2887,N_2213,N_2175);
xnor U2888 (N_2888,N_2354,N_2135);
nand U2889 (N_2889,N_2333,N_2132);
xor U2890 (N_2890,N_2366,N_2410);
and U2891 (N_2891,N_2397,N_2470);
and U2892 (N_2892,N_2284,N_2306);
and U2893 (N_2893,N_2460,N_2326);
xor U2894 (N_2894,N_2136,N_2232);
and U2895 (N_2895,N_2266,N_2088);
and U2896 (N_2896,N_2016,N_2068);
or U2897 (N_2897,N_2248,N_2390);
nand U2898 (N_2898,N_2062,N_2080);
and U2899 (N_2899,N_2372,N_2364);
or U2900 (N_2900,N_2327,N_2030);
xor U2901 (N_2901,N_2127,N_2483);
xor U2902 (N_2902,N_2112,N_2399);
nand U2903 (N_2903,N_2054,N_2319);
and U2904 (N_2904,N_2145,N_2173);
xor U2905 (N_2905,N_2470,N_2124);
or U2906 (N_2906,N_2060,N_2434);
nor U2907 (N_2907,N_2383,N_2180);
and U2908 (N_2908,N_2162,N_2251);
nor U2909 (N_2909,N_2425,N_2285);
or U2910 (N_2910,N_2392,N_2309);
nor U2911 (N_2911,N_2182,N_2237);
and U2912 (N_2912,N_2356,N_2487);
nor U2913 (N_2913,N_2369,N_2367);
and U2914 (N_2914,N_2404,N_2258);
nand U2915 (N_2915,N_2420,N_2390);
xor U2916 (N_2916,N_2081,N_2049);
or U2917 (N_2917,N_2223,N_2013);
xor U2918 (N_2918,N_2151,N_2211);
nor U2919 (N_2919,N_2325,N_2397);
nand U2920 (N_2920,N_2015,N_2315);
nor U2921 (N_2921,N_2213,N_2418);
or U2922 (N_2922,N_2276,N_2259);
nor U2923 (N_2923,N_2381,N_2373);
or U2924 (N_2924,N_2149,N_2239);
xnor U2925 (N_2925,N_2064,N_2077);
xnor U2926 (N_2926,N_2303,N_2455);
and U2927 (N_2927,N_2491,N_2201);
nor U2928 (N_2928,N_2132,N_2419);
nor U2929 (N_2929,N_2439,N_2075);
or U2930 (N_2930,N_2105,N_2289);
or U2931 (N_2931,N_2332,N_2122);
and U2932 (N_2932,N_2382,N_2091);
xor U2933 (N_2933,N_2359,N_2344);
and U2934 (N_2934,N_2208,N_2085);
nor U2935 (N_2935,N_2363,N_2029);
nand U2936 (N_2936,N_2038,N_2116);
and U2937 (N_2937,N_2130,N_2268);
nor U2938 (N_2938,N_2354,N_2225);
and U2939 (N_2939,N_2446,N_2415);
nor U2940 (N_2940,N_2216,N_2128);
and U2941 (N_2941,N_2024,N_2170);
and U2942 (N_2942,N_2027,N_2450);
nand U2943 (N_2943,N_2102,N_2144);
or U2944 (N_2944,N_2107,N_2421);
nor U2945 (N_2945,N_2134,N_2280);
nor U2946 (N_2946,N_2155,N_2241);
nand U2947 (N_2947,N_2133,N_2372);
and U2948 (N_2948,N_2308,N_2315);
or U2949 (N_2949,N_2386,N_2315);
xnor U2950 (N_2950,N_2233,N_2161);
or U2951 (N_2951,N_2112,N_2039);
nor U2952 (N_2952,N_2349,N_2227);
and U2953 (N_2953,N_2314,N_2437);
nand U2954 (N_2954,N_2475,N_2351);
nand U2955 (N_2955,N_2384,N_2216);
nor U2956 (N_2956,N_2342,N_2295);
nand U2957 (N_2957,N_2095,N_2019);
nand U2958 (N_2958,N_2088,N_2305);
or U2959 (N_2959,N_2175,N_2226);
and U2960 (N_2960,N_2341,N_2365);
and U2961 (N_2961,N_2415,N_2343);
nand U2962 (N_2962,N_2471,N_2151);
nor U2963 (N_2963,N_2440,N_2095);
or U2964 (N_2964,N_2405,N_2269);
nor U2965 (N_2965,N_2237,N_2332);
xor U2966 (N_2966,N_2390,N_2160);
nor U2967 (N_2967,N_2037,N_2312);
or U2968 (N_2968,N_2296,N_2036);
xnor U2969 (N_2969,N_2453,N_2270);
nor U2970 (N_2970,N_2212,N_2430);
or U2971 (N_2971,N_2227,N_2364);
nor U2972 (N_2972,N_2310,N_2392);
nor U2973 (N_2973,N_2215,N_2387);
nor U2974 (N_2974,N_2312,N_2014);
or U2975 (N_2975,N_2038,N_2486);
xor U2976 (N_2976,N_2088,N_2359);
nor U2977 (N_2977,N_2299,N_2122);
nor U2978 (N_2978,N_2023,N_2341);
nand U2979 (N_2979,N_2074,N_2013);
nor U2980 (N_2980,N_2192,N_2333);
or U2981 (N_2981,N_2160,N_2312);
nand U2982 (N_2982,N_2229,N_2114);
nor U2983 (N_2983,N_2363,N_2403);
nor U2984 (N_2984,N_2125,N_2214);
or U2985 (N_2985,N_2261,N_2490);
xor U2986 (N_2986,N_2170,N_2082);
nand U2987 (N_2987,N_2431,N_2325);
nor U2988 (N_2988,N_2051,N_2307);
xor U2989 (N_2989,N_2296,N_2346);
or U2990 (N_2990,N_2162,N_2222);
nand U2991 (N_2991,N_2047,N_2093);
and U2992 (N_2992,N_2096,N_2043);
and U2993 (N_2993,N_2169,N_2256);
or U2994 (N_2994,N_2250,N_2044);
nand U2995 (N_2995,N_2180,N_2495);
nand U2996 (N_2996,N_2103,N_2210);
nand U2997 (N_2997,N_2315,N_2178);
nand U2998 (N_2998,N_2437,N_2177);
xor U2999 (N_2999,N_2136,N_2446);
and U3000 (N_3000,N_2685,N_2866);
nor U3001 (N_3001,N_2793,N_2500);
and U3002 (N_3002,N_2507,N_2799);
nor U3003 (N_3003,N_2669,N_2970);
xor U3004 (N_3004,N_2791,N_2630);
xnor U3005 (N_3005,N_2573,N_2895);
or U3006 (N_3006,N_2883,N_2703);
xor U3007 (N_3007,N_2702,N_2504);
or U3008 (N_3008,N_2602,N_2898);
nand U3009 (N_3009,N_2706,N_2789);
or U3010 (N_3010,N_2779,N_2939);
and U3011 (N_3011,N_2731,N_2931);
and U3012 (N_3012,N_2603,N_2869);
xnor U3013 (N_3013,N_2567,N_2528);
xor U3014 (N_3014,N_2981,N_2548);
nand U3015 (N_3015,N_2966,N_2655);
xor U3016 (N_3016,N_2677,N_2776);
and U3017 (N_3017,N_2783,N_2599);
and U3018 (N_3018,N_2620,N_2916);
and U3019 (N_3019,N_2950,N_2597);
xnor U3020 (N_3020,N_2834,N_2541);
and U3021 (N_3021,N_2634,N_2800);
and U3022 (N_3022,N_2814,N_2594);
nor U3023 (N_3023,N_2907,N_2721);
or U3024 (N_3024,N_2593,N_2554);
nand U3025 (N_3025,N_2980,N_2524);
or U3026 (N_3026,N_2804,N_2932);
xor U3027 (N_3027,N_2662,N_2707);
nor U3028 (N_3028,N_2592,N_2945);
and U3029 (N_3029,N_2969,N_2775);
xor U3030 (N_3030,N_2736,N_2838);
nor U3031 (N_3031,N_2515,N_2823);
nand U3032 (N_3032,N_2739,N_2583);
and U3033 (N_3033,N_2718,N_2608);
nand U3034 (N_3034,N_2660,N_2965);
and U3035 (N_3035,N_2624,N_2732);
and U3036 (N_3036,N_2742,N_2816);
and U3037 (N_3037,N_2896,N_2714);
nand U3038 (N_3038,N_2615,N_2882);
or U3039 (N_3039,N_2790,N_2581);
nand U3040 (N_3040,N_2847,N_2688);
nor U3041 (N_3041,N_2754,N_2934);
nor U3042 (N_3042,N_2664,N_2935);
or U3043 (N_3043,N_2854,N_2505);
and U3044 (N_3044,N_2535,N_2533);
and U3045 (N_3045,N_2610,N_2788);
nor U3046 (N_3046,N_2880,N_2698);
or U3047 (N_3047,N_2958,N_2606);
xnor U3048 (N_3048,N_2991,N_2760);
and U3049 (N_3049,N_2792,N_2753);
or U3050 (N_3050,N_2873,N_2650);
xor U3051 (N_3051,N_2727,N_2673);
xor U3052 (N_3052,N_2512,N_2946);
or U3053 (N_3053,N_2879,N_2519);
nand U3054 (N_3054,N_2918,N_2808);
nor U3055 (N_3055,N_2740,N_2700);
nand U3056 (N_3056,N_2928,N_2711);
nand U3057 (N_3057,N_2552,N_2770);
and U3058 (N_3058,N_2737,N_2676);
nor U3059 (N_3059,N_2961,N_2848);
nor U3060 (N_3060,N_2794,N_2513);
nand U3061 (N_3061,N_2805,N_2510);
xor U3062 (N_3062,N_2871,N_2623);
nand U3063 (N_3063,N_2622,N_2645);
nor U3064 (N_3064,N_2837,N_2972);
or U3065 (N_3065,N_2810,N_2647);
or U3066 (N_3066,N_2734,N_2690);
and U3067 (N_3067,N_2643,N_2547);
nor U3068 (N_3068,N_2941,N_2876);
and U3069 (N_3069,N_2526,N_2521);
or U3070 (N_3070,N_2828,N_2614);
xor U3071 (N_3071,N_2658,N_2682);
nand U3072 (N_3072,N_2644,N_2699);
and U3073 (N_3073,N_2832,N_2944);
xor U3074 (N_3074,N_2953,N_2830);
nand U3075 (N_3075,N_2988,N_2891);
nand U3076 (N_3076,N_2766,N_2723);
and U3077 (N_3077,N_2708,N_2910);
or U3078 (N_3078,N_2557,N_2514);
xor U3079 (N_3079,N_2843,N_2661);
nor U3080 (N_3080,N_2815,N_2929);
xnor U3081 (N_3081,N_2963,N_2726);
nand U3082 (N_3082,N_2822,N_2582);
nor U3083 (N_3083,N_2782,N_2983);
xor U3084 (N_3084,N_2888,N_2671);
nand U3085 (N_3085,N_2956,N_2984);
nand U3086 (N_3086,N_2856,N_2572);
and U3087 (N_3087,N_2884,N_2577);
or U3088 (N_3088,N_2564,N_2553);
xnor U3089 (N_3089,N_2659,N_2917);
nand U3090 (N_3090,N_2860,N_2600);
or U3091 (N_3091,N_2738,N_2691);
nand U3092 (N_3092,N_2839,N_2976);
xnor U3093 (N_3093,N_2584,N_2508);
or U3094 (N_3094,N_2914,N_2818);
or U3095 (N_3095,N_2536,N_2806);
and U3096 (N_3096,N_2601,N_2679);
and U3097 (N_3097,N_2563,N_2777);
xor U3098 (N_3098,N_2820,N_2803);
xor U3099 (N_3099,N_2619,N_2696);
or U3100 (N_3100,N_2947,N_2587);
nor U3101 (N_3101,N_2865,N_2892);
and U3102 (N_3102,N_2973,N_2885);
and U3103 (N_3103,N_2750,N_2666);
nand U3104 (N_3104,N_2921,N_2545);
or U3105 (N_3105,N_2641,N_2616);
nand U3106 (N_3106,N_2844,N_2765);
nand U3107 (N_3107,N_2943,N_2652);
xor U3108 (N_3108,N_2518,N_2653);
nor U3109 (N_3109,N_2825,N_2640);
and U3110 (N_3110,N_2618,N_2925);
nor U3111 (N_3111,N_2933,N_2751);
nand U3112 (N_3112,N_2670,N_2719);
nor U3113 (N_3113,N_2511,N_2809);
or U3114 (N_3114,N_2938,N_2665);
and U3115 (N_3115,N_2772,N_2850);
nor U3116 (N_3116,N_2561,N_2555);
and U3117 (N_3117,N_2683,N_2530);
nor U3118 (N_3118,N_2802,N_2786);
or U3119 (N_3119,N_2836,N_2798);
xnor U3120 (N_3120,N_2975,N_2648);
and U3121 (N_3121,N_2784,N_2900);
and U3122 (N_3122,N_2773,N_2657);
nor U3123 (N_3123,N_2940,N_2764);
xor U3124 (N_3124,N_2638,N_2951);
or U3125 (N_3125,N_2542,N_2912);
or U3126 (N_3126,N_2558,N_2748);
and U3127 (N_3127,N_2845,N_2565);
xnor U3128 (N_3128,N_2566,N_2857);
nand U3129 (N_3129,N_2853,N_2957);
nand U3130 (N_3130,N_2801,N_2893);
nor U3131 (N_3131,N_2831,N_2813);
nor U3132 (N_3132,N_2855,N_2632);
xor U3133 (N_3133,N_2543,N_2859);
nor U3134 (N_3134,N_2967,N_2654);
xnor U3135 (N_3135,N_2626,N_2590);
and U3136 (N_3136,N_2827,N_2894);
or U3137 (N_3137,N_2756,N_2501);
and U3138 (N_3138,N_2897,N_2908);
nor U3139 (N_3139,N_2550,N_2846);
or U3140 (N_3140,N_2874,N_2715);
nand U3141 (N_3141,N_2529,N_2864);
and U3142 (N_3142,N_2964,N_2675);
xnor U3143 (N_3143,N_2716,N_2639);
or U3144 (N_3144,N_2663,N_2523);
and U3145 (N_3145,N_2559,N_2995);
or U3146 (N_3146,N_2960,N_2588);
or U3147 (N_3147,N_2977,N_2628);
and U3148 (N_3148,N_2686,N_2911);
and U3149 (N_3149,N_2769,N_2781);
or U3150 (N_3150,N_2642,N_2717);
nor U3151 (N_3151,N_2927,N_2605);
nand U3152 (N_3152,N_2684,N_2858);
nor U3153 (N_3153,N_2817,N_2704);
nor U3154 (N_3154,N_2695,N_2520);
nand U3155 (N_3155,N_2625,N_2901);
xor U3156 (N_3156,N_2534,N_2771);
and U3157 (N_3157,N_2758,N_2978);
and U3158 (N_3158,N_2621,N_2595);
or U3159 (N_3159,N_2612,N_2668);
or U3160 (N_3160,N_2959,N_2861);
or U3161 (N_3161,N_2752,N_2955);
nor U3162 (N_3162,N_2755,N_2949);
nand U3163 (N_3163,N_2607,N_2948);
or U3164 (N_3164,N_2899,N_2926);
xnor U3165 (N_3165,N_2701,N_2531);
nor U3166 (N_3166,N_2906,N_2749);
and U3167 (N_3167,N_2937,N_2913);
and U3168 (N_3168,N_2870,N_2591);
xnor U3169 (N_3169,N_2611,N_2835);
xor U3170 (N_3170,N_2778,N_2637);
nand U3171 (N_3171,N_2598,N_2841);
nor U3172 (N_3172,N_2730,N_2886);
nand U3173 (N_3173,N_2936,N_2728);
nor U3174 (N_3174,N_2763,N_2852);
nand U3175 (N_3175,N_2924,N_2902);
nand U3176 (N_3176,N_2881,N_2979);
xor U3177 (N_3177,N_2585,N_2575);
and U3178 (N_3178,N_2517,N_2712);
nand U3179 (N_3179,N_2586,N_2785);
or U3180 (N_3180,N_2889,N_2672);
nor U3181 (N_3181,N_2849,N_2743);
nor U3182 (N_3182,N_2952,N_2851);
nand U3183 (N_3183,N_2747,N_2705);
or U3184 (N_3184,N_2887,N_2689);
or U3185 (N_3185,N_2819,N_2503);
and U3186 (N_3186,N_2506,N_2992);
and U3187 (N_3187,N_2560,N_2971);
nand U3188 (N_3188,N_2627,N_2741);
nand U3189 (N_3189,N_2746,N_2811);
xnor U3190 (N_3190,N_2930,N_2720);
nor U3191 (N_3191,N_2633,N_2631);
nand U3192 (N_3192,N_2905,N_2525);
and U3193 (N_3193,N_2875,N_2544);
or U3194 (N_3194,N_2968,N_2868);
xor U3195 (N_3195,N_2768,N_2826);
or U3196 (N_3196,N_2985,N_2556);
xor U3197 (N_3197,N_2589,N_2878);
and U3198 (N_3198,N_2527,N_2986);
nor U3199 (N_3199,N_2571,N_2812);
and U3200 (N_3200,N_2993,N_2574);
or U3201 (N_3201,N_2797,N_2942);
or U3202 (N_3202,N_2516,N_2569);
nor U3203 (N_3203,N_2745,N_2609);
or U3204 (N_3204,N_2999,N_2694);
or U3205 (N_3205,N_2646,N_2909);
xor U3206 (N_3206,N_2962,N_2502);
nand U3207 (N_3207,N_2725,N_2997);
nor U3208 (N_3208,N_2681,N_2903);
or U3209 (N_3209,N_2733,N_2551);
or U3210 (N_3210,N_2570,N_2509);
nor U3211 (N_3211,N_2920,N_2998);
xor U3212 (N_3212,N_2915,N_2767);
nor U3213 (N_3213,N_2890,N_2987);
nand U3214 (N_3214,N_2678,N_2613);
and U3215 (N_3215,N_2989,N_2693);
nand U3216 (N_3216,N_2635,N_2774);
xnor U3217 (N_3217,N_2568,N_2821);
nand U3218 (N_3218,N_2636,N_2576);
xor U3219 (N_3219,N_2762,N_2872);
nor U3220 (N_3220,N_2722,N_2829);
and U3221 (N_3221,N_2994,N_2629);
nand U3222 (N_3222,N_2796,N_2759);
xnor U3223 (N_3223,N_2562,N_2862);
nor U3224 (N_3224,N_2824,N_2990);
xnor U3225 (N_3225,N_2579,N_2724);
nand U3226 (N_3226,N_2596,N_2709);
or U3227 (N_3227,N_2537,N_2974);
and U3228 (N_3228,N_2649,N_2538);
and U3229 (N_3229,N_2807,N_2667);
nor U3230 (N_3230,N_2546,N_2744);
xor U3231 (N_3231,N_2580,N_2840);
nand U3232 (N_3232,N_2713,N_2617);
or U3233 (N_3233,N_2729,N_2522);
xnor U3234 (N_3234,N_2757,N_2863);
nand U3235 (N_3235,N_2680,N_2687);
nor U3236 (N_3236,N_2833,N_2651);
and U3237 (N_3237,N_2982,N_2922);
xnor U3238 (N_3238,N_2919,N_2532);
xnor U3239 (N_3239,N_2842,N_2604);
nor U3240 (N_3240,N_2877,N_2710);
nand U3241 (N_3241,N_2549,N_2656);
and U3242 (N_3242,N_2867,N_2923);
nand U3243 (N_3243,N_2692,N_2735);
or U3244 (N_3244,N_2996,N_2787);
and U3245 (N_3245,N_2795,N_2697);
and U3246 (N_3246,N_2674,N_2540);
xnor U3247 (N_3247,N_2761,N_2954);
nand U3248 (N_3248,N_2578,N_2780);
nor U3249 (N_3249,N_2904,N_2539);
or U3250 (N_3250,N_2840,N_2715);
nor U3251 (N_3251,N_2792,N_2919);
nor U3252 (N_3252,N_2505,N_2708);
nor U3253 (N_3253,N_2889,N_2984);
nor U3254 (N_3254,N_2842,N_2916);
nor U3255 (N_3255,N_2542,N_2721);
or U3256 (N_3256,N_2978,N_2815);
xor U3257 (N_3257,N_2889,N_2568);
and U3258 (N_3258,N_2863,N_2614);
nand U3259 (N_3259,N_2993,N_2892);
nand U3260 (N_3260,N_2907,N_2799);
xnor U3261 (N_3261,N_2501,N_2854);
xnor U3262 (N_3262,N_2904,N_2959);
nor U3263 (N_3263,N_2819,N_2665);
or U3264 (N_3264,N_2668,N_2542);
nor U3265 (N_3265,N_2596,N_2863);
nand U3266 (N_3266,N_2906,N_2857);
or U3267 (N_3267,N_2861,N_2815);
xnor U3268 (N_3268,N_2829,N_2826);
nand U3269 (N_3269,N_2554,N_2619);
nor U3270 (N_3270,N_2820,N_2968);
or U3271 (N_3271,N_2692,N_2657);
or U3272 (N_3272,N_2917,N_2989);
nor U3273 (N_3273,N_2946,N_2587);
xor U3274 (N_3274,N_2864,N_2743);
or U3275 (N_3275,N_2661,N_2576);
or U3276 (N_3276,N_2562,N_2763);
nor U3277 (N_3277,N_2561,N_2545);
nand U3278 (N_3278,N_2506,N_2608);
xor U3279 (N_3279,N_2501,N_2601);
and U3280 (N_3280,N_2912,N_2803);
xor U3281 (N_3281,N_2649,N_2562);
or U3282 (N_3282,N_2986,N_2662);
or U3283 (N_3283,N_2892,N_2516);
nand U3284 (N_3284,N_2833,N_2766);
xor U3285 (N_3285,N_2959,N_2754);
or U3286 (N_3286,N_2727,N_2746);
xnor U3287 (N_3287,N_2565,N_2607);
xnor U3288 (N_3288,N_2573,N_2501);
nor U3289 (N_3289,N_2888,N_2625);
xor U3290 (N_3290,N_2850,N_2594);
nand U3291 (N_3291,N_2658,N_2524);
xor U3292 (N_3292,N_2786,N_2835);
nor U3293 (N_3293,N_2756,N_2550);
nor U3294 (N_3294,N_2835,N_2666);
or U3295 (N_3295,N_2675,N_2633);
xnor U3296 (N_3296,N_2778,N_2563);
nor U3297 (N_3297,N_2815,N_2955);
and U3298 (N_3298,N_2583,N_2865);
nor U3299 (N_3299,N_2755,N_2883);
and U3300 (N_3300,N_2894,N_2815);
or U3301 (N_3301,N_2534,N_2596);
and U3302 (N_3302,N_2907,N_2560);
nor U3303 (N_3303,N_2832,N_2825);
nor U3304 (N_3304,N_2692,N_2874);
or U3305 (N_3305,N_2955,N_2639);
xor U3306 (N_3306,N_2900,N_2723);
nand U3307 (N_3307,N_2989,N_2986);
and U3308 (N_3308,N_2559,N_2793);
nor U3309 (N_3309,N_2715,N_2720);
nor U3310 (N_3310,N_2933,N_2865);
xnor U3311 (N_3311,N_2785,N_2786);
or U3312 (N_3312,N_2753,N_2937);
nand U3313 (N_3313,N_2697,N_2555);
or U3314 (N_3314,N_2542,N_2659);
and U3315 (N_3315,N_2682,N_2970);
or U3316 (N_3316,N_2559,N_2908);
or U3317 (N_3317,N_2962,N_2969);
or U3318 (N_3318,N_2792,N_2694);
nand U3319 (N_3319,N_2855,N_2971);
nor U3320 (N_3320,N_2946,N_2863);
and U3321 (N_3321,N_2850,N_2928);
nor U3322 (N_3322,N_2867,N_2524);
and U3323 (N_3323,N_2974,N_2916);
xnor U3324 (N_3324,N_2783,N_2835);
and U3325 (N_3325,N_2792,N_2787);
or U3326 (N_3326,N_2877,N_2730);
nand U3327 (N_3327,N_2882,N_2942);
nor U3328 (N_3328,N_2810,N_2754);
nor U3329 (N_3329,N_2632,N_2670);
nor U3330 (N_3330,N_2678,N_2627);
or U3331 (N_3331,N_2582,N_2787);
xnor U3332 (N_3332,N_2711,N_2713);
nor U3333 (N_3333,N_2778,N_2727);
xnor U3334 (N_3334,N_2738,N_2957);
or U3335 (N_3335,N_2908,N_2869);
nand U3336 (N_3336,N_2818,N_2879);
xnor U3337 (N_3337,N_2569,N_2723);
nor U3338 (N_3338,N_2967,N_2624);
nand U3339 (N_3339,N_2880,N_2787);
or U3340 (N_3340,N_2815,N_2617);
nor U3341 (N_3341,N_2962,N_2669);
nor U3342 (N_3342,N_2959,N_2797);
or U3343 (N_3343,N_2544,N_2695);
xnor U3344 (N_3344,N_2640,N_2541);
and U3345 (N_3345,N_2846,N_2952);
xnor U3346 (N_3346,N_2518,N_2992);
and U3347 (N_3347,N_2865,N_2698);
nor U3348 (N_3348,N_2789,N_2840);
or U3349 (N_3349,N_2845,N_2668);
xnor U3350 (N_3350,N_2561,N_2650);
and U3351 (N_3351,N_2782,N_2660);
and U3352 (N_3352,N_2514,N_2828);
nand U3353 (N_3353,N_2763,N_2560);
nand U3354 (N_3354,N_2654,N_2685);
nand U3355 (N_3355,N_2868,N_2611);
nor U3356 (N_3356,N_2865,N_2956);
nand U3357 (N_3357,N_2902,N_2611);
nand U3358 (N_3358,N_2909,N_2687);
or U3359 (N_3359,N_2680,N_2679);
xnor U3360 (N_3360,N_2936,N_2572);
xnor U3361 (N_3361,N_2550,N_2904);
xnor U3362 (N_3362,N_2901,N_2692);
xor U3363 (N_3363,N_2747,N_2749);
or U3364 (N_3364,N_2563,N_2889);
xnor U3365 (N_3365,N_2606,N_2568);
nand U3366 (N_3366,N_2996,N_2953);
nor U3367 (N_3367,N_2674,N_2697);
nor U3368 (N_3368,N_2782,N_2852);
nor U3369 (N_3369,N_2696,N_2853);
and U3370 (N_3370,N_2956,N_2864);
nand U3371 (N_3371,N_2825,N_2698);
or U3372 (N_3372,N_2846,N_2728);
nand U3373 (N_3373,N_2804,N_2598);
and U3374 (N_3374,N_2500,N_2668);
xnor U3375 (N_3375,N_2755,N_2668);
and U3376 (N_3376,N_2738,N_2922);
nand U3377 (N_3377,N_2993,N_2762);
or U3378 (N_3378,N_2990,N_2656);
and U3379 (N_3379,N_2996,N_2693);
or U3380 (N_3380,N_2744,N_2585);
and U3381 (N_3381,N_2516,N_2824);
or U3382 (N_3382,N_2560,N_2993);
nor U3383 (N_3383,N_2523,N_2681);
nand U3384 (N_3384,N_2943,N_2633);
and U3385 (N_3385,N_2946,N_2623);
and U3386 (N_3386,N_2662,N_2603);
nor U3387 (N_3387,N_2897,N_2525);
or U3388 (N_3388,N_2566,N_2651);
nand U3389 (N_3389,N_2650,N_2937);
or U3390 (N_3390,N_2720,N_2986);
xnor U3391 (N_3391,N_2659,N_2805);
and U3392 (N_3392,N_2521,N_2703);
or U3393 (N_3393,N_2804,N_2845);
and U3394 (N_3394,N_2887,N_2876);
nor U3395 (N_3395,N_2581,N_2817);
xor U3396 (N_3396,N_2590,N_2535);
and U3397 (N_3397,N_2698,N_2745);
nand U3398 (N_3398,N_2902,N_2775);
xor U3399 (N_3399,N_2584,N_2622);
nand U3400 (N_3400,N_2947,N_2762);
nand U3401 (N_3401,N_2847,N_2862);
nor U3402 (N_3402,N_2619,N_2604);
nand U3403 (N_3403,N_2977,N_2996);
nor U3404 (N_3404,N_2564,N_2773);
xor U3405 (N_3405,N_2585,N_2941);
and U3406 (N_3406,N_2731,N_2980);
and U3407 (N_3407,N_2829,N_2801);
nand U3408 (N_3408,N_2867,N_2804);
nand U3409 (N_3409,N_2661,N_2865);
nor U3410 (N_3410,N_2943,N_2989);
nand U3411 (N_3411,N_2937,N_2856);
or U3412 (N_3412,N_2982,N_2630);
and U3413 (N_3413,N_2842,N_2926);
and U3414 (N_3414,N_2979,N_2540);
or U3415 (N_3415,N_2786,N_2569);
and U3416 (N_3416,N_2672,N_2609);
or U3417 (N_3417,N_2517,N_2948);
or U3418 (N_3418,N_2710,N_2978);
or U3419 (N_3419,N_2765,N_2661);
and U3420 (N_3420,N_2842,N_2616);
and U3421 (N_3421,N_2615,N_2521);
and U3422 (N_3422,N_2523,N_2720);
nor U3423 (N_3423,N_2645,N_2985);
or U3424 (N_3424,N_2895,N_2516);
or U3425 (N_3425,N_2775,N_2989);
or U3426 (N_3426,N_2896,N_2706);
and U3427 (N_3427,N_2704,N_2842);
or U3428 (N_3428,N_2729,N_2639);
or U3429 (N_3429,N_2975,N_2621);
nor U3430 (N_3430,N_2913,N_2681);
nand U3431 (N_3431,N_2547,N_2798);
nand U3432 (N_3432,N_2976,N_2851);
xnor U3433 (N_3433,N_2943,N_2862);
or U3434 (N_3434,N_2619,N_2543);
nor U3435 (N_3435,N_2759,N_2898);
nand U3436 (N_3436,N_2613,N_2846);
nor U3437 (N_3437,N_2763,N_2546);
and U3438 (N_3438,N_2632,N_2643);
nand U3439 (N_3439,N_2909,N_2892);
nand U3440 (N_3440,N_2804,N_2590);
or U3441 (N_3441,N_2573,N_2528);
nor U3442 (N_3442,N_2947,N_2633);
nand U3443 (N_3443,N_2550,N_2690);
xor U3444 (N_3444,N_2525,N_2770);
nand U3445 (N_3445,N_2678,N_2982);
nand U3446 (N_3446,N_2989,N_2928);
nand U3447 (N_3447,N_2712,N_2989);
nand U3448 (N_3448,N_2669,N_2577);
nand U3449 (N_3449,N_2784,N_2750);
nand U3450 (N_3450,N_2724,N_2816);
nand U3451 (N_3451,N_2586,N_2862);
and U3452 (N_3452,N_2813,N_2522);
nor U3453 (N_3453,N_2671,N_2777);
nor U3454 (N_3454,N_2749,N_2981);
nor U3455 (N_3455,N_2627,N_2942);
nor U3456 (N_3456,N_2711,N_2532);
xnor U3457 (N_3457,N_2921,N_2608);
nor U3458 (N_3458,N_2601,N_2847);
xor U3459 (N_3459,N_2776,N_2570);
and U3460 (N_3460,N_2645,N_2683);
xor U3461 (N_3461,N_2642,N_2720);
nor U3462 (N_3462,N_2953,N_2539);
or U3463 (N_3463,N_2850,N_2837);
xnor U3464 (N_3464,N_2909,N_2630);
xnor U3465 (N_3465,N_2722,N_2595);
xor U3466 (N_3466,N_2796,N_2951);
xor U3467 (N_3467,N_2524,N_2506);
xor U3468 (N_3468,N_2906,N_2723);
or U3469 (N_3469,N_2869,N_2634);
nor U3470 (N_3470,N_2694,N_2610);
nand U3471 (N_3471,N_2989,N_2792);
nand U3472 (N_3472,N_2535,N_2739);
nor U3473 (N_3473,N_2994,N_2834);
xnor U3474 (N_3474,N_2829,N_2695);
or U3475 (N_3475,N_2759,N_2573);
or U3476 (N_3476,N_2992,N_2578);
xnor U3477 (N_3477,N_2793,N_2660);
xnor U3478 (N_3478,N_2650,N_2668);
nor U3479 (N_3479,N_2594,N_2994);
or U3480 (N_3480,N_2718,N_2529);
nand U3481 (N_3481,N_2644,N_2875);
xnor U3482 (N_3482,N_2633,N_2823);
xnor U3483 (N_3483,N_2614,N_2637);
nand U3484 (N_3484,N_2588,N_2675);
or U3485 (N_3485,N_2519,N_2711);
nand U3486 (N_3486,N_2939,N_2694);
nand U3487 (N_3487,N_2665,N_2575);
nor U3488 (N_3488,N_2744,N_2568);
or U3489 (N_3489,N_2672,N_2698);
and U3490 (N_3490,N_2580,N_2809);
and U3491 (N_3491,N_2727,N_2618);
and U3492 (N_3492,N_2943,N_2895);
xnor U3493 (N_3493,N_2813,N_2925);
nor U3494 (N_3494,N_2910,N_2552);
and U3495 (N_3495,N_2681,N_2961);
and U3496 (N_3496,N_2815,N_2641);
and U3497 (N_3497,N_2895,N_2528);
or U3498 (N_3498,N_2753,N_2854);
xnor U3499 (N_3499,N_2656,N_2534);
xor U3500 (N_3500,N_3058,N_3092);
and U3501 (N_3501,N_3018,N_3355);
and U3502 (N_3502,N_3363,N_3081);
nor U3503 (N_3503,N_3195,N_3272);
or U3504 (N_3504,N_3332,N_3020);
nor U3505 (N_3505,N_3388,N_3215);
or U3506 (N_3506,N_3105,N_3167);
nand U3507 (N_3507,N_3139,N_3153);
xor U3508 (N_3508,N_3032,N_3224);
xnor U3509 (N_3509,N_3364,N_3226);
or U3510 (N_3510,N_3422,N_3119);
or U3511 (N_3511,N_3108,N_3383);
xor U3512 (N_3512,N_3181,N_3262);
and U3513 (N_3513,N_3396,N_3314);
nand U3514 (N_3514,N_3008,N_3243);
xnor U3515 (N_3515,N_3354,N_3234);
and U3516 (N_3516,N_3285,N_3039);
xnor U3517 (N_3517,N_3009,N_3391);
and U3518 (N_3518,N_3397,N_3325);
and U3519 (N_3519,N_3407,N_3085);
and U3520 (N_3520,N_3466,N_3434);
and U3521 (N_3521,N_3436,N_3442);
and U3522 (N_3522,N_3437,N_3278);
nor U3523 (N_3523,N_3468,N_3074);
xnor U3524 (N_3524,N_3155,N_3250);
and U3525 (N_3525,N_3275,N_3118);
or U3526 (N_3526,N_3412,N_3140);
nand U3527 (N_3527,N_3003,N_3327);
nand U3528 (N_3528,N_3190,N_3471);
or U3529 (N_3529,N_3143,N_3337);
and U3530 (N_3530,N_3241,N_3300);
nor U3531 (N_3531,N_3304,N_3473);
or U3532 (N_3532,N_3417,N_3485);
nor U3533 (N_3533,N_3191,N_3295);
or U3534 (N_3534,N_3086,N_3141);
nor U3535 (N_3535,N_3299,N_3414);
or U3536 (N_3536,N_3494,N_3024);
nand U3537 (N_3537,N_3330,N_3015);
or U3538 (N_3538,N_3258,N_3308);
nand U3539 (N_3539,N_3274,N_3227);
and U3540 (N_3540,N_3264,N_3446);
nor U3541 (N_3541,N_3331,N_3377);
or U3542 (N_3542,N_3328,N_3373);
nand U3543 (N_3543,N_3060,N_3429);
and U3544 (N_3544,N_3135,N_3161);
nor U3545 (N_3545,N_3448,N_3265);
nor U3546 (N_3546,N_3075,N_3114);
or U3547 (N_3547,N_3115,N_3045);
nor U3548 (N_3548,N_3061,N_3362);
xor U3549 (N_3549,N_3482,N_3251);
xor U3550 (N_3550,N_3145,N_3342);
and U3551 (N_3551,N_3177,N_3217);
nor U3552 (N_3552,N_3212,N_3253);
nand U3553 (N_3553,N_3340,N_3451);
or U3554 (N_3554,N_3420,N_3378);
and U3555 (N_3555,N_3293,N_3172);
or U3556 (N_3556,N_3033,N_3384);
and U3557 (N_3557,N_3360,N_3110);
nor U3558 (N_3558,N_3409,N_3333);
nor U3559 (N_3559,N_3049,N_3102);
nor U3560 (N_3560,N_3284,N_3270);
nor U3561 (N_3561,N_3151,N_3395);
nor U3562 (N_3562,N_3126,N_3123);
nand U3563 (N_3563,N_3089,N_3438);
and U3564 (N_3564,N_3146,N_3310);
nor U3565 (N_3565,N_3210,N_3221);
xor U3566 (N_3566,N_3326,N_3324);
nor U3567 (N_3567,N_3184,N_3113);
and U3568 (N_3568,N_3339,N_3180);
and U3569 (N_3569,N_3367,N_3256);
nand U3570 (N_3570,N_3399,N_3164);
xnor U3571 (N_3571,N_3338,N_3286);
nor U3572 (N_3572,N_3387,N_3385);
and U3573 (N_3573,N_3239,N_3276);
and U3574 (N_3574,N_3321,N_3219);
nor U3575 (N_3575,N_3044,N_3431);
nand U3576 (N_3576,N_3109,N_3347);
nand U3577 (N_3577,N_3163,N_3398);
or U3578 (N_3578,N_3148,N_3366);
xnor U3579 (N_3579,N_3159,N_3288);
nand U3580 (N_3580,N_3218,N_3400);
and U3581 (N_3581,N_3281,N_3273);
and U3582 (N_3582,N_3068,N_3296);
nor U3583 (N_3583,N_3090,N_3361);
nor U3584 (N_3584,N_3402,N_3376);
nand U3585 (N_3585,N_3025,N_3200);
nand U3586 (N_3586,N_3306,N_3059);
nor U3587 (N_3587,N_3271,N_3392);
or U3588 (N_3588,N_3419,N_3460);
nor U3589 (N_3589,N_3433,N_3100);
xor U3590 (N_3590,N_3229,N_3470);
xnor U3591 (N_3591,N_3223,N_3449);
nor U3592 (N_3592,N_3290,N_3173);
or U3593 (N_3593,N_3474,N_3487);
nand U3594 (N_3594,N_3078,N_3477);
xor U3595 (N_3595,N_3323,N_3403);
nand U3596 (N_3596,N_3370,N_3443);
or U3597 (N_3597,N_3000,N_3201);
or U3598 (N_3598,N_3231,N_3406);
or U3599 (N_3599,N_3206,N_3149);
or U3600 (N_3600,N_3182,N_3205);
or U3601 (N_3601,N_3103,N_3080);
and U3602 (N_3602,N_3185,N_3382);
and U3603 (N_3603,N_3386,N_3237);
nor U3604 (N_3604,N_3111,N_3415);
or U3605 (N_3605,N_3405,N_3309);
nor U3606 (N_3606,N_3193,N_3246);
and U3607 (N_3607,N_3097,N_3475);
nand U3608 (N_3608,N_3079,N_3315);
nor U3609 (N_3609,N_3244,N_3313);
xnor U3610 (N_3610,N_3496,N_3104);
or U3611 (N_3611,N_3101,N_3374);
xnor U3612 (N_3612,N_3359,N_3152);
or U3613 (N_3613,N_3302,N_3428);
nand U3614 (N_3614,N_3390,N_3194);
nor U3615 (N_3615,N_3432,N_3445);
xor U3616 (N_3616,N_3322,N_3425);
and U3617 (N_3617,N_3413,N_3121);
and U3618 (N_3618,N_3444,N_3063);
xor U3619 (N_3619,N_3187,N_3014);
nand U3620 (N_3620,N_3174,N_3418);
nor U3621 (N_3621,N_3001,N_3156);
nor U3622 (N_3622,N_3381,N_3052);
and U3623 (N_3623,N_3497,N_3458);
xor U3624 (N_3624,N_3055,N_3481);
and U3625 (N_3625,N_3165,N_3358);
and U3626 (N_3626,N_3027,N_3457);
nor U3627 (N_3627,N_3401,N_3357);
and U3628 (N_3628,N_3245,N_3125);
nor U3629 (N_3629,N_3236,N_3248);
or U3630 (N_3630,N_3053,N_3178);
and U3631 (N_3631,N_3346,N_3454);
nor U3632 (N_3632,N_3169,N_3352);
and U3633 (N_3633,N_3465,N_3077);
nor U3634 (N_3634,N_3380,N_3269);
or U3635 (N_3635,N_3051,N_3120);
nor U3636 (N_3636,N_3137,N_3450);
xor U3637 (N_3637,N_3435,N_3179);
or U3638 (N_3638,N_3127,N_3176);
nor U3639 (N_3639,N_3283,N_3461);
nand U3640 (N_3640,N_3479,N_3233);
nor U3641 (N_3641,N_3301,N_3073);
xnor U3642 (N_3642,N_3260,N_3307);
xnor U3643 (N_3643,N_3011,N_3082);
or U3644 (N_3644,N_3211,N_3144);
and U3645 (N_3645,N_3188,N_3131);
or U3646 (N_3646,N_3375,N_3368);
nand U3647 (N_3647,N_3472,N_3069);
nand U3648 (N_3648,N_3006,N_3026);
nand U3649 (N_3649,N_3087,N_3186);
xnor U3650 (N_3650,N_3096,N_3279);
and U3651 (N_3651,N_3335,N_3136);
and U3652 (N_3652,N_3094,N_3037);
or U3653 (N_3653,N_3343,N_3491);
or U3654 (N_3654,N_3192,N_3305);
or U3655 (N_3655,N_3235,N_3430);
or U3656 (N_3656,N_3336,N_3005);
or U3657 (N_3657,N_3099,N_3289);
xnor U3658 (N_3658,N_3088,N_3266);
nand U3659 (N_3659,N_3469,N_3122);
xnor U3660 (N_3660,N_3257,N_3222);
nand U3661 (N_3661,N_3066,N_3345);
nand U3662 (N_3662,N_3204,N_3083);
nor U3663 (N_3663,N_3416,N_3132);
or U3664 (N_3664,N_3440,N_3456);
nand U3665 (N_3665,N_3452,N_3054);
and U3666 (N_3666,N_3394,N_3389);
or U3667 (N_3667,N_3207,N_3404);
nand U3668 (N_3668,N_3411,N_3356);
nand U3669 (N_3669,N_3214,N_3147);
nor U3670 (N_3670,N_3040,N_3316);
xnor U3671 (N_3671,N_3424,N_3130);
or U3672 (N_3672,N_3490,N_3280);
nor U3673 (N_3673,N_3017,N_3162);
and U3674 (N_3674,N_3166,N_3303);
and U3675 (N_3675,N_3463,N_3171);
and U3676 (N_3676,N_3483,N_3216);
and U3677 (N_3677,N_3042,N_3455);
nand U3678 (N_3678,N_3209,N_3203);
and U3679 (N_3679,N_3028,N_3220);
nor U3680 (N_3680,N_3029,N_3124);
xor U3681 (N_3681,N_3261,N_3294);
xnor U3682 (N_3682,N_3098,N_3369);
or U3683 (N_3683,N_3268,N_3493);
xor U3684 (N_3684,N_3050,N_3007);
nand U3685 (N_3685,N_3016,N_3072);
nand U3686 (N_3686,N_3255,N_3318);
nand U3687 (N_3687,N_3202,N_3478);
and U3688 (N_3688,N_3439,N_3071);
nor U3689 (N_3689,N_3311,N_3351);
and U3690 (N_3690,N_3070,N_3480);
and U3691 (N_3691,N_3117,N_3057);
nand U3692 (N_3692,N_3441,N_3213);
xor U3693 (N_3693,N_3030,N_3199);
or U3694 (N_3694,N_3393,N_3189);
nand U3695 (N_3695,N_3160,N_3486);
nand U3696 (N_3696,N_3043,N_3022);
or U3697 (N_3697,N_3196,N_3154);
and U3698 (N_3698,N_3031,N_3208);
xor U3699 (N_3699,N_3348,N_3067);
nor U3700 (N_3700,N_3365,N_3046);
and U3701 (N_3701,N_3168,N_3112);
nand U3702 (N_3702,N_3426,N_3464);
xor U3703 (N_3703,N_3263,N_3242);
or U3704 (N_3704,N_3021,N_3349);
xor U3705 (N_3705,N_3353,N_3423);
nand U3706 (N_3706,N_3427,N_3372);
or U3707 (N_3707,N_3129,N_3116);
or U3708 (N_3708,N_3467,N_3408);
xor U3709 (N_3709,N_3459,N_3107);
and U3710 (N_3710,N_3056,N_3198);
or U3711 (N_3711,N_3095,N_3462);
nand U3712 (N_3712,N_3488,N_3133);
nor U3713 (N_3713,N_3228,N_3492);
and U3714 (N_3714,N_3065,N_3238);
nand U3715 (N_3715,N_3498,N_3254);
nor U3716 (N_3716,N_3225,N_3453);
and U3717 (N_3717,N_3476,N_3175);
xor U3718 (N_3718,N_3170,N_3240);
nor U3719 (N_3719,N_3350,N_3230);
nand U3720 (N_3720,N_3319,N_3041);
nor U3721 (N_3721,N_3267,N_3499);
and U3722 (N_3722,N_3048,N_3091);
xor U3723 (N_3723,N_3138,N_3287);
or U3724 (N_3724,N_3004,N_3034);
nand U3725 (N_3725,N_3371,N_3232);
and U3726 (N_3726,N_3247,N_3019);
or U3727 (N_3727,N_3142,N_3023);
nand U3728 (N_3728,N_3329,N_3197);
or U3729 (N_3729,N_3047,N_3334);
xor U3730 (N_3730,N_3344,N_3012);
nor U3731 (N_3731,N_3489,N_3084);
or U3732 (N_3732,N_3277,N_3035);
xor U3733 (N_3733,N_3134,N_3128);
and U3734 (N_3734,N_3291,N_3317);
xor U3735 (N_3735,N_3106,N_3076);
and U3736 (N_3736,N_3410,N_3038);
xnor U3737 (N_3737,N_3158,N_3282);
or U3738 (N_3738,N_3379,N_3447);
and U3739 (N_3739,N_3421,N_3298);
nor U3740 (N_3740,N_3002,N_3062);
xnor U3741 (N_3741,N_3150,N_3157);
nand U3742 (N_3742,N_3093,N_3320);
and U3743 (N_3743,N_3013,N_3297);
or U3744 (N_3744,N_3341,N_3259);
nor U3745 (N_3745,N_3312,N_3183);
xor U3746 (N_3746,N_3484,N_3252);
and U3747 (N_3747,N_3036,N_3010);
and U3748 (N_3748,N_3064,N_3495);
or U3749 (N_3749,N_3249,N_3292);
or U3750 (N_3750,N_3199,N_3356);
and U3751 (N_3751,N_3430,N_3014);
nor U3752 (N_3752,N_3348,N_3147);
xnor U3753 (N_3753,N_3115,N_3030);
or U3754 (N_3754,N_3059,N_3141);
nor U3755 (N_3755,N_3368,N_3175);
nand U3756 (N_3756,N_3110,N_3405);
xor U3757 (N_3757,N_3336,N_3360);
xor U3758 (N_3758,N_3059,N_3010);
and U3759 (N_3759,N_3472,N_3021);
nor U3760 (N_3760,N_3492,N_3280);
and U3761 (N_3761,N_3191,N_3333);
and U3762 (N_3762,N_3080,N_3135);
or U3763 (N_3763,N_3155,N_3061);
and U3764 (N_3764,N_3495,N_3033);
nor U3765 (N_3765,N_3418,N_3052);
nand U3766 (N_3766,N_3076,N_3158);
xnor U3767 (N_3767,N_3380,N_3181);
xnor U3768 (N_3768,N_3192,N_3145);
or U3769 (N_3769,N_3484,N_3113);
nor U3770 (N_3770,N_3121,N_3103);
and U3771 (N_3771,N_3126,N_3066);
and U3772 (N_3772,N_3229,N_3303);
or U3773 (N_3773,N_3117,N_3340);
nor U3774 (N_3774,N_3106,N_3209);
or U3775 (N_3775,N_3044,N_3276);
nor U3776 (N_3776,N_3454,N_3233);
and U3777 (N_3777,N_3470,N_3222);
or U3778 (N_3778,N_3297,N_3238);
and U3779 (N_3779,N_3032,N_3039);
or U3780 (N_3780,N_3480,N_3458);
xnor U3781 (N_3781,N_3407,N_3193);
nor U3782 (N_3782,N_3014,N_3204);
nand U3783 (N_3783,N_3022,N_3329);
nor U3784 (N_3784,N_3143,N_3321);
and U3785 (N_3785,N_3167,N_3282);
or U3786 (N_3786,N_3477,N_3451);
nor U3787 (N_3787,N_3008,N_3194);
nand U3788 (N_3788,N_3275,N_3018);
or U3789 (N_3789,N_3262,N_3326);
nor U3790 (N_3790,N_3291,N_3238);
or U3791 (N_3791,N_3356,N_3227);
nand U3792 (N_3792,N_3184,N_3004);
and U3793 (N_3793,N_3054,N_3182);
nor U3794 (N_3794,N_3222,N_3085);
nand U3795 (N_3795,N_3017,N_3170);
and U3796 (N_3796,N_3421,N_3294);
or U3797 (N_3797,N_3066,N_3164);
and U3798 (N_3798,N_3374,N_3104);
nor U3799 (N_3799,N_3336,N_3016);
nor U3800 (N_3800,N_3355,N_3436);
xnor U3801 (N_3801,N_3147,N_3116);
nor U3802 (N_3802,N_3179,N_3307);
or U3803 (N_3803,N_3128,N_3299);
nor U3804 (N_3804,N_3446,N_3404);
xnor U3805 (N_3805,N_3169,N_3155);
xor U3806 (N_3806,N_3163,N_3216);
xor U3807 (N_3807,N_3085,N_3134);
nand U3808 (N_3808,N_3432,N_3122);
nand U3809 (N_3809,N_3036,N_3336);
and U3810 (N_3810,N_3167,N_3178);
nor U3811 (N_3811,N_3220,N_3260);
xnor U3812 (N_3812,N_3290,N_3183);
nand U3813 (N_3813,N_3077,N_3426);
nand U3814 (N_3814,N_3044,N_3469);
or U3815 (N_3815,N_3190,N_3133);
or U3816 (N_3816,N_3143,N_3469);
or U3817 (N_3817,N_3278,N_3383);
nand U3818 (N_3818,N_3082,N_3295);
or U3819 (N_3819,N_3363,N_3259);
nor U3820 (N_3820,N_3404,N_3415);
nor U3821 (N_3821,N_3055,N_3185);
nand U3822 (N_3822,N_3378,N_3016);
or U3823 (N_3823,N_3211,N_3467);
and U3824 (N_3824,N_3019,N_3340);
and U3825 (N_3825,N_3410,N_3349);
xnor U3826 (N_3826,N_3026,N_3021);
xnor U3827 (N_3827,N_3263,N_3265);
nor U3828 (N_3828,N_3283,N_3451);
and U3829 (N_3829,N_3059,N_3233);
and U3830 (N_3830,N_3315,N_3437);
or U3831 (N_3831,N_3304,N_3074);
nor U3832 (N_3832,N_3232,N_3029);
or U3833 (N_3833,N_3322,N_3250);
nor U3834 (N_3834,N_3196,N_3135);
xor U3835 (N_3835,N_3233,N_3298);
or U3836 (N_3836,N_3365,N_3476);
xnor U3837 (N_3837,N_3078,N_3373);
nand U3838 (N_3838,N_3089,N_3094);
nand U3839 (N_3839,N_3054,N_3309);
and U3840 (N_3840,N_3213,N_3099);
nor U3841 (N_3841,N_3408,N_3207);
xor U3842 (N_3842,N_3029,N_3003);
nand U3843 (N_3843,N_3068,N_3471);
or U3844 (N_3844,N_3484,N_3444);
and U3845 (N_3845,N_3070,N_3437);
and U3846 (N_3846,N_3376,N_3129);
or U3847 (N_3847,N_3209,N_3232);
or U3848 (N_3848,N_3114,N_3045);
nor U3849 (N_3849,N_3455,N_3482);
nor U3850 (N_3850,N_3196,N_3046);
or U3851 (N_3851,N_3103,N_3345);
xnor U3852 (N_3852,N_3386,N_3209);
nor U3853 (N_3853,N_3297,N_3023);
or U3854 (N_3854,N_3183,N_3042);
or U3855 (N_3855,N_3162,N_3395);
nand U3856 (N_3856,N_3402,N_3355);
nand U3857 (N_3857,N_3431,N_3024);
xor U3858 (N_3858,N_3002,N_3475);
or U3859 (N_3859,N_3166,N_3219);
or U3860 (N_3860,N_3298,N_3230);
nand U3861 (N_3861,N_3472,N_3019);
xor U3862 (N_3862,N_3165,N_3272);
nand U3863 (N_3863,N_3450,N_3082);
nand U3864 (N_3864,N_3422,N_3239);
or U3865 (N_3865,N_3246,N_3269);
nand U3866 (N_3866,N_3042,N_3154);
or U3867 (N_3867,N_3411,N_3466);
or U3868 (N_3868,N_3078,N_3086);
or U3869 (N_3869,N_3413,N_3497);
xnor U3870 (N_3870,N_3352,N_3275);
or U3871 (N_3871,N_3204,N_3218);
and U3872 (N_3872,N_3020,N_3389);
nand U3873 (N_3873,N_3223,N_3393);
and U3874 (N_3874,N_3092,N_3493);
nand U3875 (N_3875,N_3215,N_3015);
or U3876 (N_3876,N_3174,N_3333);
nand U3877 (N_3877,N_3222,N_3427);
xor U3878 (N_3878,N_3447,N_3304);
nand U3879 (N_3879,N_3006,N_3278);
xor U3880 (N_3880,N_3441,N_3283);
nand U3881 (N_3881,N_3257,N_3390);
or U3882 (N_3882,N_3308,N_3171);
or U3883 (N_3883,N_3122,N_3294);
nor U3884 (N_3884,N_3002,N_3370);
or U3885 (N_3885,N_3285,N_3257);
nor U3886 (N_3886,N_3129,N_3397);
and U3887 (N_3887,N_3278,N_3082);
or U3888 (N_3888,N_3451,N_3472);
nor U3889 (N_3889,N_3217,N_3254);
nand U3890 (N_3890,N_3083,N_3377);
and U3891 (N_3891,N_3034,N_3341);
and U3892 (N_3892,N_3002,N_3399);
xor U3893 (N_3893,N_3411,N_3445);
xnor U3894 (N_3894,N_3080,N_3159);
xnor U3895 (N_3895,N_3234,N_3161);
and U3896 (N_3896,N_3484,N_3133);
and U3897 (N_3897,N_3215,N_3120);
and U3898 (N_3898,N_3323,N_3452);
xor U3899 (N_3899,N_3070,N_3193);
xor U3900 (N_3900,N_3269,N_3058);
or U3901 (N_3901,N_3480,N_3128);
nor U3902 (N_3902,N_3345,N_3123);
xor U3903 (N_3903,N_3449,N_3235);
and U3904 (N_3904,N_3481,N_3495);
and U3905 (N_3905,N_3140,N_3316);
and U3906 (N_3906,N_3318,N_3116);
and U3907 (N_3907,N_3254,N_3209);
or U3908 (N_3908,N_3386,N_3202);
nand U3909 (N_3909,N_3480,N_3362);
nor U3910 (N_3910,N_3159,N_3116);
nand U3911 (N_3911,N_3360,N_3409);
nand U3912 (N_3912,N_3160,N_3438);
and U3913 (N_3913,N_3126,N_3414);
xor U3914 (N_3914,N_3382,N_3294);
and U3915 (N_3915,N_3228,N_3412);
nand U3916 (N_3916,N_3063,N_3484);
or U3917 (N_3917,N_3124,N_3112);
nor U3918 (N_3918,N_3067,N_3269);
or U3919 (N_3919,N_3225,N_3113);
nand U3920 (N_3920,N_3277,N_3168);
or U3921 (N_3921,N_3302,N_3165);
and U3922 (N_3922,N_3202,N_3378);
nand U3923 (N_3923,N_3172,N_3180);
xor U3924 (N_3924,N_3116,N_3165);
and U3925 (N_3925,N_3359,N_3160);
or U3926 (N_3926,N_3047,N_3099);
and U3927 (N_3927,N_3350,N_3366);
nand U3928 (N_3928,N_3444,N_3318);
xor U3929 (N_3929,N_3161,N_3444);
or U3930 (N_3930,N_3181,N_3264);
nand U3931 (N_3931,N_3158,N_3404);
and U3932 (N_3932,N_3301,N_3104);
and U3933 (N_3933,N_3119,N_3455);
and U3934 (N_3934,N_3298,N_3002);
and U3935 (N_3935,N_3343,N_3320);
or U3936 (N_3936,N_3219,N_3307);
and U3937 (N_3937,N_3290,N_3140);
or U3938 (N_3938,N_3232,N_3215);
and U3939 (N_3939,N_3091,N_3130);
nand U3940 (N_3940,N_3334,N_3078);
and U3941 (N_3941,N_3057,N_3139);
nor U3942 (N_3942,N_3415,N_3064);
xnor U3943 (N_3943,N_3085,N_3212);
nand U3944 (N_3944,N_3319,N_3433);
or U3945 (N_3945,N_3134,N_3064);
nor U3946 (N_3946,N_3178,N_3307);
or U3947 (N_3947,N_3435,N_3261);
nand U3948 (N_3948,N_3349,N_3314);
nor U3949 (N_3949,N_3132,N_3014);
xor U3950 (N_3950,N_3406,N_3133);
nand U3951 (N_3951,N_3284,N_3436);
and U3952 (N_3952,N_3241,N_3020);
nor U3953 (N_3953,N_3119,N_3290);
xnor U3954 (N_3954,N_3045,N_3145);
xnor U3955 (N_3955,N_3307,N_3209);
or U3956 (N_3956,N_3105,N_3355);
nand U3957 (N_3957,N_3100,N_3262);
nand U3958 (N_3958,N_3360,N_3291);
nor U3959 (N_3959,N_3320,N_3351);
and U3960 (N_3960,N_3069,N_3471);
and U3961 (N_3961,N_3159,N_3462);
and U3962 (N_3962,N_3323,N_3146);
or U3963 (N_3963,N_3010,N_3255);
and U3964 (N_3964,N_3198,N_3261);
nor U3965 (N_3965,N_3026,N_3304);
xor U3966 (N_3966,N_3187,N_3233);
xor U3967 (N_3967,N_3103,N_3171);
xnor U3968 (N_3968,N_3423,N_3480);
and U3969 (N_3969,N_3134,N_3306);
xnor U3970 (N_3970,N_3093,N_3169);
and U3971 (N_3971,N_3339,N_3027);
nor U3972 (N_3972,N_3016,N_3045);
nor U3973 (N_3973,N_3237,N_3376);
nor U3974 (N_3974,N_3394,N_3050);
nand U3975 (N_3975,N_3037,N_3168);
xnor U3976 (N_3976,N_3283,N_3050);
xnor U3977 (N_3977,N_3026,N_3028);
xor U3978 (N_3978,N_3185,N_3110);
and U3979 (N_3979,N_3116,N_3197);
or U3980 (N_3980,N_3379,N_3005);
or U3981 (N_3981,N_3328,N_3486);
nor U3982 (N_3982,N_3310,N_3043);
nor U3983 (N_3983,N_3491,N_3428);
xnor U3984 (N_3984,N_3313,N_3484);
or U3985 (N_3985,N_3470,N_3210);
nand U3986 (N_3986,N_3247,N_3484);
nand U3987 (N_3987,N_3290,N_3478);
or U3988 (N_3988,N_3406,N_3156);
and U3989 (N_3989,N_3209,N_3125);
and U3990 (N_3990,N_3030,N_3155);
nor U3991 (N_3991,N_3496,N_3351);
nor U3992 (N_3992,N_3142,N_3127);
xnor U3993 (N_3993,N_3212,N_3485);
nor U3994 (N_3994,N_3185,N_3170);
nor U3995 (N_3995,N_3456,N_3330);
nand U3996 (N_3996,N_3092,N_3397);
and U3997 (N_3997,N_3216,N_3123);
or U3998 (N_3998,N_3403,N_3240);
nand U3999 (N_3999,N_3250,N_3438);
or U4000 (N_4000,N_3951,N_3520);
and U4001 (N_4001,N_3871,N_3767);
or U4002 (N_4002,N_3642,N_3672);
nor U4003 (N_4003,N_3911,N_3541);
nor U4004 (N_4004,N_3762,N_3724);
and U4005 (N_4005,N_3573,N_3514);
or U4006 (N_4006,N_3879,N_3568);
or U4007 (N_4007,N_3868,N_3974);
nand U4008 (N_4008,N_3622,N_3554);
or U4009 (N_4009,N_3846,N_3935);
and U4010 (N_4010,N_3667,N_3722);
xor U4011 (N_4011,N_3854,N_3768);
or U4012 (N_4012,N_3753,N_3612);
xnor U4013 (N_4013,N_3836,N_3534);
nand U4014 (N_4014,N_3602,N_3660);
nand U4015 (N_4015,N_3536,N_3609);
or U4016 (N_4016,N_3979,N_3988);
nand U4017 (N_4017,N_3574,N_3699);
nand U4018 (N_4018,N_3645,N_3616);
nand U4019 (N_4019,N_3530,N_3511);
nand U4020 (N_4020,N_3505,N_3682);
xnor U4021 (N_4021,N_3857,N_3590);
xnor U4022 (N_4022,N_3973,N_3926);
or U4023 (N_4023,N_3500,N_3748);
and U4024 (N_4024,N_3819,N_3631);
nor U4025 (N_4025,N_3607,N_3987);
xnor U4026 (N_4026,N_3847,N_3833);
nor U4027 (N_4027,N_3501,N_3962);
xor U4028 (N_4028,N_3910,N_3659);
and U4029 (N_4029,N_3653,N_3579);
nand U4030 (N_4030,N_3878,N_3998);
nand U4031 (N_4031,N_3595,N_3900);
nor U4032 (N_4032,N_3688,N_3882);
or U4033 (N_4033,N_3877,N_3634);
or U4034 (N_4034,N_3733,N_3725);
nand U4035 (N_4035,N_3632,N_3508);
nor U4036 (N_4036,N_3807,N_3796);
nor U4037 (N_4037,N_3611,N_3542);
or U4038 (N_4038,N_3557,N_3975);
nor U4039 (N_4039,N_3740,N_3739);
or U4040 (N_4040,N_3537,N_3841);
nor U4041 (N_4041,N_3775,N_3670);
nand U4042 (N_4042,N_3799,N_3647);
nor U4043 (N_4043,N_3738,N_3745);
nor U4044 (N_4044,N_3756,N_3897);
xnor U4045 (N_4045,N_3872,N_3695);
xnor U4046 (N_4046,N_3548,N_3842);
nor U4047 (N_4047,N_3896,N_3582);
and U4048 (N_4048,N_3583,N_3652);
and U4049 (N_4049,N_3571,N_3736);
nor U4050 (N_4050,N_3933,N_3845);
nor U4051 (N_4051,N_3665,N_3808);
and U4052 (N_4052,N_3726,N_3706);
nor U4053 (N_4053,N_3860,N_3608);
and U4054 (N_4054,N_3886,N_3522);
or U4055 (N_4055,N_3676,N_3664);
xnor U4056 (N_4056,N_3742,N_3884);
or U4057 (N_4057,N_3965,N_3918);
or U4058 (N_4058,N_3627,N_3957);
and U4059 (N_4059,N_3707,N_3787);
nand U4060 (N_4060,N_3635,N_3892);
nand U4061 (N_4061,N_3912,N_3732);
nor U4062 (N_4062,N_3749,N_3856);
nand U4063 (N_4063,N_3598,N_3779);
xnor U4064 (N_4064,N_3949,N_3853);
and U4065 (N_4065,N_3790,N_3914);
nor U4066 (N_4066,N_3778,N_3967);
or U4067 (N_4067,N_3629,N_3773);
nor U4068 (N_4068,N_3902,N_3690);
or U4069 (N_4069,N_3633,N_3939);
nor U4070 (N_4070,N_3813,N_3662);
nor U4071 (N_4071,N_3937,N_3521);
xor U4072 (N_4072,N_3874,N_3989);
and U4073 (N_4073,N_3889,N_3519);
nor U4074 (N_4074,N_3771,N_3596);
and U4075 (N_4075,N_3980,N_3531);
xnor U4076 (N_4076,N_3524,N_3785);
and U4077 (N_4077,N_3552,N_3862);
xor U4078 (N_4078,N_3948,N_3620);
nor U4079 (N_4079,N_3700,N_3977);
and U4080 (N_4080,N_3539,N_3936);
or U4081 (N_4081,N_3512,N_3619);
nor U4082 (N_4082,N_3945,N_3705);
and U4083 (N_4083,N_3716,N_3708);
nand U4084 (N_4084,N_3529,N_3567);
nand U4085 (N_4085,N_3625,N_3502);
or U4086 (N_4086,N_3562,N_3769);
xor U4087 (N_4087,N_3824,N_3817);
xnor U4088 (N_4088,N_3990,N_3992);
nand U4089 (N_4089,N_3650,N_3592);
nor U4090 (N_4090,N_3802,N_3535);
or U4091 (N_4091,N_3932,N_3995);
xnor U4092 (N_4092,N_3666,N_3919);
nand U4093 (N_4093,N_3747,N_3798);
nor U4094 (N_4094,N_3735,N_3513);
and U4095 (N_4095,N_3526,N_3834);
or U4096 (N_4096,N_3680,N_3674);
and U4097 (N_4097,N_3822,N_3823);
nand U4098 (N_4098,N_3533,N_3963);
and U4099 (N_4099,N_3538,N_3528);
nand U4100 (N_4100,N_3844,N_3786);
nor U4101 (N_4101,N_3576,N_3744);
and U4102 (N_4102,N_3811,N_3876);
nor U4103 (N_4103,N_3614,N_3848);
or U4104 (N_4104,N_3924,N_3907);
nor U4105 (N_4105,N_3656,N_3651);
xor U4106 (N_4106,N_3774,N_3546);
nor U4107 (N_4107,N_3859,N_3503);
or U4108 (N_4108,N_3594,N_3560);
nor U4109 (N_4109,N_3961,N_3928);
nor U4110 (N_4110,N_3584,N_3960);
xnor U4111 (N_4111,N_3555,N_3639);
and U4112 (N_4112,N_3899,N_3814);
nor U4113 (N_4113,N_3850,N_3578);
or U4114 (N_4114,N_3941,N_3603);
or U4115 (N_4115,N_3718,N_3757);
or U4116 (N_4116,N_3999,N_3991);
and U4117 (N_4117,N_3646,N_3921);
and U4118 (N_4118,N_3809,N_3580);
or U4119 (N_4119,N_3515,N_3587);
nand U4120 (N_4120,N_3835,N_3766);
and U4121 (N_4121,N_3678,N_3687);
nor U4122 (N_4122,N_3806,N_3628);
or U4123 (N_4123,N_3715,N_3610);
or U4124 (N_4124,N_3597,N_3981);
and U4125 (N_4125,N_3543,N_3916);
or U4126 (N_4126,N_3908,N_3764);
nor U4127 (N_4127,N_3689,N_3818);
or U4128 (N_4128,N_3801,N_3940);
nor U4129 (N_4129,N_3586,N_3870);
nand U4130 (N_4130,N_3968,N_3922);
nand U4131 (N_4131,N_3805,N_3750);
nor U4132 (N_4132,N_3923,N_3517);
nor U4133 (N_4133,N_3885,N_3605);
and U4134 (N_4134,N_3506,N_3626);
xor U4135 (N_4135,N_3955,N_3730);
xor U4136 (N_4136,N_3971,N_3559);
or U4137 (N_4137,N_3997,N_3780);
nand U4138 (N_4138,N_3901,N_3741);
and U4139 (N_4139,N_3697,N_3723);
nor U4140 (N_4140,N_3832,N_3701);
or U4141 (N_4141,N_3952,N_3864);
nor U4142 (N_4142,N_3729,N_3821);
and U4143 (N_4143,N_3930,N_3869);
nor U4144 (N_4144,N_3863,N_3934);
xor U4145 (N_4145,N_3585,N_3804);
and U4146 (N_4146,N_3712,N_3770);
and U4147 (N_4147,N_3601,N_3589);
or U4148 (N_4148,N_3691,N_3649);
nor U4149 (N_4149,N_3615,N_3840);
and U4150 (N_4150,N_3710,N_3743);
nand U4151 (N_4151,N_3684,N_3721);
nand U4152 (N_4152,N_3637,N_3925);
nor U4153 (N_4153,N_3719,N_3976);
nand U4154 (N_4154,N_3958,N_3713);
nor U4155 (N_4155,N_3772,N_3570);
xnor U4156 (N_4156,N_3669,N_3903);
or U4157 (N_4157,N_3793,N_3668);
and U4158 (N_4158,N_3891,N_3827);
nand U4159 (N_4159,N_3890,N_3964);
nor U4160 (N_4160,N_3826,N_3830);
nor U4161 (N_4161,N_3504,N_3881);
and U4162 (N_4162,N_3569,N_3581);
xor U4163 (N_4163,N_3895,N_3759);
nand U4164 (N_4164,N_3692,N_3643);
nand U4165 (N_4165,N_3946,N_3913);
nor U4166 (N_4166,N_3624,N_3509);
nand U4167 (N_4167,N_3898,N_3993);
or U4168 (N_4168,N_3800,N_3956);
and U4169 (N_4169,N_3905,N_3852);
or U4170 (N_4170,N_3711,N_3788);
nor U4171 (N_4171,N_3544,N_3588);
or U4172 (N_4172,N_3858,N_3686);
xor U4173 (N_4173,N_3763,N_3904);
xor U4174 (N_4174,N_3888,N_3969);
or U4175 (N_4175,N_3752,N_3755);
nand U4176 (N_4176,N_3549,N_3641);
and U4177 (N_4177,N_3754,N_3783);
xor U4178 (N_4178,N_3865,N_3915);
xor U4179 (N_4179,N_3781,N_3657);
nand U4180 (N_4180,N_3654,N_3673);
xnor U4181 (N_4181,N_3617,N_3606);
nor U4182 (N_4182,N_3867,N_3621);
or U4183 (N_4183,N_3599,N_3855);
and U4184 (N_4184,N_3825,N_3618);
and U4185 (N_4185,N_3683,N_3640);
or U4186 (N_4186,N_3986,N_3816);
and U4187 (N_4187,N_3746,N_3677);
xor U4188 (N_4188,N_3734,N_3685);
nand U4189 (N_4189,N_3681,N_3709);
nand U4190 (N_4190,N_3839,N_3970);
nor U4191 (N_4191,N_3828,N_3810);
nor U4192 (N_4192,N_3547,N_3572);
xor U4193 (N_4193,N_3812,N_3727);
nor U4194 (N_4194,N_3703,N_3658);
and U4195 (N_4195,N_3765,N_3532);
xor U4196 (N_4196,N_3873,N_3943);
and U4197 (N_4197,N_3613,N_3556);
and U4198 (N_4198,N_3604,N_3558);
nand U4199 (N_4199,N_3887,N_3954);
and U4200 (N_4200,N_3523,N_3815);
nand U4201 (N_4201,N_3953,N_3663);
xnor U4202 (N_4202,N_3829,N_3545);
nand U4203 (N_4203,N_3671,N_3917);
nand U4204 (N_4204,N_3507,N_3527);
nor U4205 (N_4205,N_3655,N_3861);
nand U4206 (N_4206,N_3564,N_3577);
or U4207 (N_4207,N_3920,N_3894);
xnor U4208 (N_4208,N_3893,N_3983);
nand U4209 (N_4209,N_3931,N_3797);
or U4210 (N_4210,N_3978,N_3820);
or U4211 (N_4211,N_3794,N_3883);
xnor U4212 (N_4212,N_3837,N_3696);
nor U4213 (N_4213,N_3760,N_3942);
nand U4214 (N_4214,N_3525,N_3906);
xor U4215 (N_4215,N_3575,N_3803);
nor U4216 (N_4216,N_3792,N_3630);
and U4217 (N_4217,N_3866,N_3994);
nor U4218 (N_4218,N_3551,N_3784);
or U4219 (N_4219,N_3758,N_3563);
and U4220 (N_4220,N_3591,N_3984);
nand U4221 (N_4221,N_3623,N_3518);
and U4222 (N_4222,N_3791,N_3927);
and U4223 (N_4223,N_3661,N_3789);
xor U4224 (N_4224,N_3944,N_3720);
or U4225 (N_4225,N_3875,N_3929);
xor U4226 (N_4226,N_3838,N_3761);
xor U4227 (N_4227,N_3731,N_3714);
nor U4228 (N_4228,N_3694,N_3516);
nand U4229 (N_4229,N_3648,N_3831);
or U4230 (N_4230,N_3737,N_3553);
or U4231 (N_4231,N_3795,N_3849);
or U4232 (N_4232,N_3947,N_3704);
or U4233 (N_4233,N_3693,N_3959);
nor U4234 (N_4234,N_3982,N_3566);
and U4235 (N_4235,N_3510,N_3717);
or U4236 (N_4236,N_3550,N_3675);
xor U4237 (N_4237,N_3777,N_3966);
and U4238 (N_4238,N_3728,N_3950);
nand U4239 (N_4239,N_3938,N_3600);
nor U4240 (N_4240,N_3638,N_3679);
xnor U4241 (N_4241,N_3644,N_3540);
and U4242 (N_4242,N_3909,N_3776);
nand U4243 (N_4243,N_3880,N_3593);
and U4244 (N_4244,N_3751,N_3636);
or U4245 (N_4245,N_3851,N_3972);
xnor U4246 (N_4246,N_3565,N_3782);
and U4247 (N_4247,N_3698,N_3996);
xor U4248 (N_4248,N_3843,N_3985);
xor U4249 (N_4249,N_3702,N_3561);
and U4250 (N_4250,N_3835,N_3708);
or U4251 (N_4251,N_3899,N_3514);
and U4252 (N_4252,N_3768,N_3727);
and U4253 (N_4253,N_3525,N_3929);
or U4254 (N_4254,N_3755,N_3792);
xnor U4255 (N_4255,N_3757,N_3551);
nor U4256 (N_4256,N_3764,N_3939);
xnor U4257 (N_4257,N_3610,N_3651);
or U4258 (N_4258,N_3540,N_3632);
nor U4259 (N_4259,N_3841,N_3838);
or U4260 (N_4260,N_3914,N_3785);
or U4261 (N_4261,N_3820,N_3676);
or U4262 (N_4262,N_3951,N_3675);
nor U4263 (N_4263,N_3530,N_3872);
nand U4264 (N_4264,N_3522,N_3708);
or U4265 (N_4265,N_3790,N_3771);
nand U4266 (N_4266,N_3862,N_3669);
nor U4267 (N_4267,N_3875,N_3554);
nor U4268 (N_4268,N_3821,N_3917);
and U4269 (N_4269,N_3713,N_3861);
or U4270 (N_4270,N_3859,N_3898);
nand U4271 (N_4271,N_3741,N_3888);
and U4272 (N_4272,N_3507,N_3587);
xor U4273 (N_4273,N_3795,N_3559);
nand U4274 (N_4274,N_3957,N_3851);
xor U4275 (N_4275,N_3970,N_3928);
nor U4276 (N_4276,N_3564,N_3644);
and U4277 (N_4277,N_3769,N_3956);
nand U4278 (N_4278,N_3784,N_3686);
and U4279 (N_4279,N_3620,N_3747);
xor U4280 (N_4280,N_3590,N_3597);
nor U4281 (N_4281,N_3653,N_3813);
xor U4282 (N_4282,N_3778,N_3965);
and U4283 (N_4283,N_3914,N_3585);
nand U4284 (N_4284,N_3531,N_3751);
xnor U4285 (N_4285,N_3537,N_3653);
nor U4286 (N_4286,N_3513,N_3614);
nand U4287 (N_4287,N_3798,N_3767);
nand U4288 (N_4288,N_3905,N_3938);
xor U4289 (N_4289,N_3947,N_3892);
nor U4290 (N_4290,N_3821,N_3940);
or U4291 (N_4291,N_3947,N_3758);
or U4292 (N_4292,N_3588,N_3706);
or U4293 (N_4293,N_3856,N_3929);
nand U4294 (N_4294,N_3907,N_3726);
nor U4295 (N_4295,N_3726,N_3895);
xnor U4296 (N_4296,N_3942,N_3812);
nor U4297 (N_4297,N_3868,N_3972);
xor U4298 (N_4298,N_3768,N_3719);
nand U4299 (N_4299,N_3533,N_3954);
nor U4300 (N_4300,N_3703,N_3579);
nor U4301 (N_4301,N_3988,N_3719);
xnor U4302 (N_4302,N_3592,N_3849);
and U4303 (N_4303,N_3566,N_3651);
and U4304 (N_4304,N_3638,N_3855);
nand U4305 (N_4305,N_3799,N_3721);
or U4306 (N_4306,N_3667,N_3904);
and U4307 (N_4307,N_3555,N_3813);
or U4308 (N_4308,N_3569,N_3997);
or U4309 (N_4309,N_3565,N_3577);
nand U4310 (N_4310,N_3852,N_3788);
and U4311 (N_4311,N_3807,N_3542);
or U4312 (N_4312,N_3585,N_3730);
xor U4313 (N_4313,N_3953,N_3617);
and U4314 (N_4314,N_3845,N_3617);
nor U4315 (N_4315,N_3823,N_3921);
nand U4316 (N_4316,N_3946,N_3606);
nor U4317 (N_4317,N_3551,N_3528);
and U4318 (N_4318,N_3537,N_3535);
or U4319 (N_4319,N_3770,N_3656);
nor U4320 (N_4320,N_3835,N_3930);
or U4321 (N_4321,N_3909,N_3880);
and U4322 (N_4322,N_3713,N_3869);
nand U4323 (N_4323,N_3867,N_3620);
nand U4324 (N_4324,N_3673,N_3623);
nand U4325 (N_4325,N_3901,N_3691);
xor U4326 (N_4326,N_3828,N_3926);
and U4327 (N_4327,N_3553,N_3551);
or U4328 (N_4328,N_3816,N_3718);
nand U4329 (N_4329,N_3542,N_3580);
or U4330 (N_4330,N_3659,N_3768);
and U4331 (N_4331,N_3750,N_3870);
and U4332 (N_4332,N_3567,N_3748);
and U4333 (N_4333,N_3763,N_3970);
or U4334 (N_4334,N_3801,N_3948);
and U4335 (N_4335,N_3841,N_3552);
xnor U4336 (N_4336,N_3788,N_3699);
nor U4337 (N_4337,N_3697,N_3908);
nand U4338 (N_4338,N_3767,N_3586);
nand U4339 (N_4339,N_3846,N_3961);
or U4340 (N_4340,N_3907,N_3902);
nand U4341 (N_4341,N_3602,N_3905);
and U4342 (N_4342,N_3855,N_3629);
nand U4343 (N_4343,N_3707,N_3538);
or U4344 (N_4344,N_3582,N_3805);
or U4345 (N_4345,N_3840,N_3565);
or U4346 (N_4346,N_3841,N_3568);
nor U4347 (N_4347,N_3997,N_3595);
or U4348 (N_4348,N_3759,N_3829);
and U4349 (N_4349,N_3693,N_3748);
or U4350 (N_4350,N_3762,N_3680);
nand U4351 (N_4351,N_3962,N_3710);
xnor U4352 (N_4352,N_3554,N_3671);
nor U4353 (N_4353,N_3753,N_3852);
nor U4354 (N_4354,N_3502,N_3710);
xor U4355 (N_4355,N_3842,N_3641);
or U4356 (N_4356,N_3966,N_3788);
and U4357 (N_4357,N_3594,N_3660);
or U4358 (N_4358,N_3949,N_3938);
and U4359 (N_4359,N_3537,N_3917);
xor U4360 (N_4360,N_3800,N_3960);
xor U4361 (N_4361,N_3784,N_3796);
nor U4362 (N_4362,N_3892,N_3624);
and U4363 (N_4363,N_3583,N_3642);
or U4364 (N_4364,N_3633,N_3831);
and U4365 (N_4365,N_3731,N_3789);
xnor U4366 (N_4366,N_3981,N_3994);
nand U4367 (N_4367,N_3712,N_3697);
nor U4368 (N_4368,N_3868,N_3895);
nand U4369 (N_4369,N_3510,N_3550);
xnor U4370 (N_4370,N_3765,N_3865);
nand U4371 (N_4371,N_3648,N_3526);
nand U4372 (N_4372,N_3582,N_3909);
nor U4373 (N_4373,N_3665,N_3751);
or U4374 (N_4374,N_3674,N_3938);
xnor U4375 (N_4375,N_3863,N_3747);
xor U4376 (N_4376,N_3904,N_3601);
or U4377 (N_4377,N_3859,N_3825);
nor U4378 (N_4378,N_3905,N_3870);
xor U4379 (N_4379,N_3778,N_3824);
and U4380 (N_4380,N_3802,N_3828);
and U4381 (N_4381,N_3779,N_3927);
nor U4382 (N_4382,N_3738,N_3653);
xnor U4383 (N_4383,N_3989,N_3942);
nand U4384 (N_4384,N_3604,N_3776);
or U4385 (N_4385,N_3556,N_3843);
or U4386 (N_4386,N_3829,N_3897);
nor U4387 (N_4387,N_3922,N_3628);
or U4388 (N_4388,N_3744,N_3960);
or U4389 (N_4389,N_3991,N_3867);
nand U4390 (N_4390,N_3602,N_3730);
xor U4391 (N_4391,N_3552,N_3810);
nand U4392 (N_4392,N_3556,N_3915);
and U4393 (N_4393,N_3654,N_3852);
and U4394 (N_4394,N_3849,N_3995);
nor U4395 (N_4395,N_3936,N_3646);
nand U4396 (N_4396,N_3652,N_3707);
xor U4397 (N_4397,N_3794,N_3530);
or U4398 (N_4398,N_3616,N_3665);
or U4399 (N_4399,N_3538,N_3725);
and U4400 (N_4400,N_3862,N_3728);
xnor U4401 (N_4401,N_3642,N_3658);
and U4402 (N_4402,N_3656,N_3871);
or U4403 (N_4403,N_3656,N_3531);
or U4404 (N_4404,N_3805,N_3759);
or U4405 (N_4405,N_3662,N_3694);
nand U4406 (N_4406,N_3725,N_3970);
nor U4407 (N_4407,N_3674,N_3739);
nor U4408 (N_4408,N_3819,N_3786);
nand U4409 (N_4409,N_3745,N_3551);
nand U4410 (N_4410,N_3729,N_3944);
nor U4411 (N_4411,N_3843,N_3869);
nand U4412 (N_4412,N_3532,N_3625);
nor U4413 (N_4413,N_3694,N_3915);
and U4414 (N_4414,N_3854,N_3875);
or U4415 (N_4415,N_3625,N_3770);
xnor U4416 (N_4416,N_3810,N_3532);
nor U4417 (N_4417,N_3809,N_3572);
nand U4418 (N_4418,N_3846,N_3605);
nor U4419 (N_4419,N_3691,N_3628);
xnor U4420 (N_4420,N_3688,N_3843);
xor U4421 (N_4421,N_3656,N_3650);
or U4422 (N_4422,N_3674,N_3791);
or U4423 (N_4423,N_3631,N_3732);
xor U4424 (N_4424,N_3665,N_3689);
nand U4425 (N_4425,N_3757,N_3581);
xor U4426 (N_4426,N_3557,N_3635);
and U4427 (N_4427,N_3544,N_3784);
nor U4428 (N_4428,N_3746,N_3828);
nand U4429 (N_4429,N_3543,N_3512);
or U4430 (N_4430,N_3549,N_3741);
nand U4431 (N_4431,N_3561,N_3781);
xnor U4432 (N_4432,N_3879,N_3694);
xor U4433 (N_4433,N_3711,N_3964);
and U4434 (N_4434,N_3536,N_3938);
nand U4435 (N_4435,N_3997,N_3547);
xor U4436 (N_4436,N_3646,N_3836);
nor U4437 (N_4437,N_3870,N_3690);
nor U4438 (N_4438,N_3817,N_3877);
and U4439 (N_4439,N_3933,N_3675);
nand U4440 (N_4440,N_3629,N_3858);
and U4441 (N_4441,N_3573,N_3570);
xor U4442 (N_4442,N_3677,N_3543);
xnor U4443 (N_4443,N_3868,N_3961);
nand U4444 (N_4444,N_3945,N_3952);
xnor U4445 (N_4445,N_3842,N_3592);
nor U4446 (N_4446,N_3578,N_3508);
and U4447 (N_4447,N_3932,N_3726);
and U4448 (N_4448,N_3989,N_3802);
and U4449 (N_4449,N_3554,N_3861);
and U4450 (N_4450,N_3645,N_3864);
or U4451 (N_4451,N_3810,N_3974);
nand U4452 (N_4452,N_3561,N_3600);
or U4453 (N_4453,N_3852,N_3631);
and U4454 (N_4454,N_3552,N_3595);
xor U4455 (N_4455,N_3684,N_3870);
and U4456 (N_4456,N_3722,N_3839);
nor U4457 (N_4457,N_3647,N_3802);
nand U4458 (N_4458,N_3879,N_3857);
or U4459 (N_4459,N_3593,N_3673);
xor U4460 (N_4460,N_3651,N_3565);
or U4461 (N_4461,N_3595,N_3691);
or U4462 (N_4462,N_3557,N_3683);
nor U4463 (N_4463,N_3842,N_3653);
nor U4464 (N_4464,N_3863,N_3630);
xor U4465 (N_4465,N_3590,N_3515);
xor U4466 (N_4466,N_3562,N_3583);
xnor U4467 (N_4467,N_3997,N_3802);
nor U4468 (N_4468,N_3840,N_3718);
or U4469 (N_4469,N_3915,N_3943);
or U4470 (N_4470,N_3508,N_3791);
nor U4471 (N_4471,N_3840,N_3734);
xor U4472 (N_4472,N_3880,N_3722);
nor U4473 (N_4473,N_3949,N_3769);
xnor U4474 (N_4474,N_3517,N_3653);
nand U4475 (N_4475,N_3963,N_3517);
nor U4476 (N_4476,N_3948,N_3602);
nand U4477 (N_4477,N_3511,N_3817);
xor U4478 (N_4478,N_3703,N_3953);
xor U4479 (N_4479,N_3661,N_3527);
and U4480 (N_4480,N_3732,N_3522);
and U4481 (N_4481,N_3707,N_3874);
nor U4482 (N_4482,N_3769,N_3790);
xor U4483 (N_4483,N_3681,N_3554);
xor U4484 (N_4484,N_3760,N_3862);
nor U4485 (N_4485,N_3978,N_3869);
or U4486 (N_4486,N_3514,N_3887);
nor U4487 (N_4487,N_3712,N_3830);
or U4488 (N_4488,N_3682,N_3897);
or U4489 (N_4489,N_3644,N_3648);
xor U4490 (N_4490,N_3901,N_3558);
xor U4491 (N_4491,N_3667,N_3653);
and U4492 (N_4492,N_3911,N_3670);
nand U4493 (N_4493,N_3804,N_3767);
nor U4494 (N_4494,N_3937,N_3783);
nand U4495 (N_4495,N_3622,N_3661);
nor U4496 (N_4496,N_3983,N_3863);
nand U4497 (N_4497,N_3659,N_3653);
or U4498 (N_4498,N_3911,N_3623);
or U4499 (N_4499,N_3777,N_3533);
and U4500 (N_4500,N_4196,N_4276);
and U4501 (N_4501,N_4390,N_4401);
nand U4502 (N_4502,N_4074,N_4095);
nand U4503 (N_4503,N_4473,N_4223);
nand U4504 (N_4504,N_4475,N_4203);
nor U4505 (N_4505,N_4462,N_4251);
nor U4506 (N_4506,N_4310,N_4319);
nor U4507 (N_4507,N_4094,N_4149);
or U4508 (N_4508,N_4138,N_4249);
xnor U4509 (N_4509,N_4481,N_4033);
nor U4510 (N_4510,N_4262,N_4266);
xnor U4511 (N_4511,N_4093,N_4122);
or U4512 (N_4512,N_4349,N_4120);
nand U4513 (N_4513,N_4205,N_4381);
nor U4514 (N_4514,N_4028,N_4082);
nand U4515 (N_4515,N_4044,N_4143);
and U4516 (N_4516,N_4380,N_4375);
and U4517 (N_4517,N_4161,N_4274);
nor U4518 (N_4518,N_4468,N_4283);
nor U4519 (N_4519,N_4499,N_4063);
and U4520 (N_4520,N_4053,N_4377);
nand U4521 (N_4521,N_4440,N_4422);
nor U4522 (N_4522,N_4035,N_4119);
xor U4523 (N_4523,N_4087,N_4491);
xnor U4524 (N_4524,N_4216,N_4024);
nor U4525 (N_4525,N_4474,N_4465);
nor U4526 (N_4526,N_4423,N_4011);
or U4527 (N_4527,N_4148,N_4088);
nor U4528 (N_4528,N_4313,N_4346);
nand U4529 (N_4529,N_4434,N_4043);
and U4530 (N_4530,N_4201,N_4306);
nand U4531 (N_4531,N_4212,N_4384);
and U4532 (N_4532,N_4322,N_4186);
or U4533 (N_4533,N_4117,N_4493);
and U4534 (N_4534,N_4029,N_4092);
nor U4535 (N_4535,N_4037,N_4027);
and U4536 (N_4536,N_4382,N_4219);
nand U4537 (N_4537,N_4160,N_4421);
and U4538 (N_4538,N_4100,N_4016);
or U4539 (N_4539,N_4064,N_4168);
nand U4540 (N_4540,N_4188,N_4000);
xor U4541 (N_4541,N_4228,N_4356);
nor U4542 (N_4542,N_4080,N_4438);
xnor U4543 (N_4543,N_4008,N_4348);
xor U4544 (N_4544,N_4159,N_4393);
or U4545 (N_4545,N_4208,N_4420);
and U4546 (N_4546,N_4373,N_4385);
or U4547 (N_4547,N_4333,N_4255);
or U4548 (N_4548,N_4351,N_4139);
xor U4549 (N_4549,N_4050,N_4362);
or U4550 (N_4550,N_4153,N_4197);
nor U4551 (N_4551,N_4206,N_4394);
or U4552 (N_4552,N_4290,N_4467);
nand U4553 (N_4553,N_4146,N_4166);
nor U4554 (N_4554,N_4032,N_4400);
or U4555 (N_4555,N_4102,N_4075);
nor U4556 (N_4556,N_4311,N_4357);
nor U4557 (N_4557,N_4424,N_4309);
xnor U4558 (N_4558,N_4198,N_4314);
nand U4559 (N_4559,N_4226,N_4361);
and U4560 (N_4560,N_4018,N_4089);
xor U4561 (N_4561,N_4469,N_4360);
nand U4562 (N_4562,N_4013,N_4183);
and U4563 (N_4563,N_4471,N_4222);
nor U4564 (N_4564,N_4456,N_4218);
nor U4565 (N_4565,N_4452,N_4334);
and U4566 (N_4566,N_4070,N_4023);
and U4567 (N_4567,N_4046,N_4060);
nor U4568 (N_4568,N_4134,N_4487);
nor U4569 (N_4569,N_4337,N_4038);
nand U4570 (N_4570,N_4057,N_4441);
nor U4571 (N_4571,N_4479,N_4386);
xor U4572 (N_4572,N_4358,N_4405);
nor U4573 (N_4573,N_4325,N_4258);
nand U4574 (N_4574,N_4498,N_4454);
xnor U4575 (N_4575,N_4254,N_4131);
nand U4576 (N_4576,N_4289,N_4485);
and U4577 (N_4577,N_4442,N_4107);
xnor U4578 (N_4578,N_4365,N_4245);
or U4579 (N_4579,N_4066,N_4132);
nand U4580 (N_4580,N_4190,N_4340);
xnor U4581 (N_4581,N_4253,N_4073);
and U4582 (N_4582,N_4490,N_4045);
or U4583 (N_4583,N_4252,N_4430);
nand U4584 (N_4584,N_4301,N_4416);
nor U4585 (N_4585,N_4352,N_4432);
nand U4586 (N_4586,N_4118,N_4484);
or U4587 (N_4587,N_4446,N_4085);
nor U4588 (N_4588,N_4112,N_4178);
xor U4589 (N_4589,N_4268,N_4215);
xnor U4590 (N_4590,N_4303,N_4002);
xor U4591 (N_4591,N_4181,N_4185);
and U4592 (N_4592,N_4154,N_4124);
and U4593 (N_4593,N_4081,N_4447);
and U4594 (N_4594,N_4317,N_4101);
xor U4595 (N_4595,N_4437,N_4388);
xnor U4596 (N_4596,N_4329,N_4391);
xor U4597 (N_4597,N_4478,N_4034);
or U4598 (N_4598,N_4343,N_4236);
and U4599 (N_4599,N_4022,N_4477);
nand U4600 (N_4600,N_4169,N_4463);
nand U4601 (N_4601,N_4195,N_4129);
or U4602 (N_4602,N_4439,N_4091);
nand U4603 (N_4603,N_4244,N_4246);
nand U4604 (N_4604,N_4009,N_4071);
xnor U4605 (N_4605,N_4040,N_4224);
and U4606 (N_4606,N_4305,N_4242);
or U4607 (N_4607,N_4058,N_4459);
or U4608 (N_4608,N_4488,N_4453);
xnor U4609 (N_4609,N_4199,N_4157);
or U4610 (N_4610,N_4059,N_4299);
nor U4611 (N_4611,N_4072,N_4426);
or U4612 (N_4612,N_4025,N_4297);
nor U4613 (N_4613,N_4372,N_4248);
or U4614 (N_4614,N_4472,N_4363);
or U4615 (N_4615,N_4189,N_4285);
nor U4616 (N_4616,N_4338,N_4328);
or U4617 (N_4617,N_4217,N_4123);
or U4618 (N_4618,N_4204,N_4069);
and U4619 (N_4619,N_4211,N_4282);
and U4620 (N_4620,N_4121,N_4062);
xor U4621 (N_4621,N_4494,N_4470);
or U4622 (N_4622,N_4003,N_4261);
nor U4623 (N_4623,N_4109,N_4387);
or U4624 (N_4624,N_4135,N_4292);
nand U4625 (N_4625,N_4144,N_4172);
and U4626 (N_4626,N_4193,N_4331);
and U4627 (N_4627,N_4140,N_4460);
nand U4628 (N_4628,N_4404,N_4096);
xor U4629 (N_4629,N_4200,N_4409);
and U4630 (N_4630,N_4184,N_4298);
nor U4631 (N_4631,N_4152,N_4145);
nand U4632 (N_4632,N_4210,N_4445);
xor U4633 (N_4633,N_4304,N_4496);
xnor U4634 (N_4634,N_4374,N_4202);
or U4635 (N_4635,N_4231,N_4302);
xnor U4636 (N_4636,N_4378,N_4015);
and U4637 (N_4637,N_4483,N_4407);
and U4638 (N_4638,N_4017,N_4489);
nand U4639 (N_4639,N_4455,N_4326);
and U4640 (N_4640,N_4175,N_4449);
or U4641 (N_4641,N_4402,N_4240);
or U4642 (N_4642,N_4376,N_4256);
nand U4643 (N_4643,N_4312,N_4339);
xnor U4644 (N_4644,N_4243,N_4280);
or U4645 (N_4645,N_4171,N_4392);
nand U4646 (N_4646,N_4300,N_4250);
or U4647 (N_4647,N_4207,N_4234);
nand U4648 (N_4648,N_4359,N_4174);
or U4649 (N_4649,N_4213,N_4464);
nor U4650 (N_4650,N_4412,N_4347);
or U4651 (N_4651,N_4461,N_4030);
nand U4652 (N_4652,N_4395,N_4238);
nand U4653 (N_4653,N_4130,N_4307);
nor U4654 (N_4654,N_4270,N_4187);
or U4655 (N_4655,N_4427,N_4042);
nor U4656 (N_4656,N_4371,N_4061);
xor U4657 (N_4657,N_4086,N_4497);
or U4658 (N_4658,N_4429,N_4342);
nor U4659 (N_4659,N_4230,N_4180);
and U4660 (N_4660,N_4012,N_4495);
xor U4661 (N_4661,N_4265,N_4067);
and U4662 (N_4662,N_4316,N_4019);
and U4663 (N_4663,N_4006,N_4237);
or U4664 (N_4664,N_4191,N_4476);
nand U4665 (N_4665,N_4021,N_4323);
or U4666 (N_4666,N_4235,N_4332);
nand U4667 (N_4667,N_4128,N_4369);
xnor U4668 (N_4668,N_4182,N_4039);
xnor U4669 (N_4669,N_4098,N_4155);
or U4670 (N_4670,N_4115,N_4167);
and U4671 (N_4671,N_4173,N_4133);
nor U4672 (N_4672,N_4403,N_4417);
and U4673 (N_4673,N_4247,N_4041);
nand U4674 (N_4674,N_4368,N_4137);
nand U4675 (N_4675,N_4435,N_4010);
nor U4676 (N_4676,N_4327,N_4036);
nand U4677 (N_4677,N_4433,N_4111);
or U4678 (N_4678,N_4320,N_4431);
or U4679 (N_4679,N_4458,N_4296);
and U4680 (N_4680,N_4354,N_4177);
and U4681 (N_4681,N_4284,N_4466);
xnor U4682 (N_4682,N_4103,N_4396);
and U4683 (N_4683,N_4104,N_4277);
or U4684 (N_4684,N_4125,N_4335);
xor U4685 (N_4685,N_4083,N_4379);
nor U4686 (N_4686,N_4436,N_4220);
and U4687 (N_4687,N_4054,N_4065);
nand U4688 (N_4688,N_4451,N_4271);
and U4689 (N_4689,N_4269,N_4076);
nor U4690 (N_4690,N_4286,N_4162);
or U4691 (N_4691,N_4194,N_4055);
or U4692 (N_4692,N_4482,N_4221);
xor U4693 (N_4693,N_4272,N_4367);
and U4694 (N_4694,N_4275,N_4084);
and U4695 (N_4695,N_4179,N_4324);
xor U4696 (N_4696,N_4389,N_4411);
or U4697 (N_4697,N_4287,N_4068);
and U4698 (N_4698,N_4142,N_4136);
or U4699 (N_4699,N_4214,N_4090);
xnor U4700 (N_4700,N_4364,N_4443);
or U4701 (N_4701,N_4229,N_4056);
xnor U4702 (N_4702,N_4233,N_4397);
nand U4703 (N_4703,N_4049,N_4077);
nor U4704 (N_4704,N_4418,N_4031);
nor U4705 (N_4705,N_4330,N_4165);
nand U4706 (N_4706,N_4047,N_4383);
or U4707 (N_4707,N_4415,N_4048);
nand U4708 (N_4708,N_4273,N_4370);
and U4709 (N_4709,N_4164,N_4163);
nor U4710 (N_4710,N_4005,N_4486);
xnor U4711 (N_4711,N_4225,N_4414);
and U4712 (N_4712,N_4116,N_4051);
nand U4713 (N_4713,N_4239,N_4156);
nand U4714 (N_4714,N_4492,N_4291);
xnor U4715 (N_4715,N_4126,N_4026);
nor U4716 (N_4716,N_4295,N_4267);
nand U4717 (N_4717,N_4114,N_4288);
nor U4718 (N_4718,N_4241,N_4308);
xor U4719 (N_4719,N_4448,N_4350);
nor U4720 (N_4720,N_4020,N_4158);
xor U4721 (N_4721,N_4004,N_4419);
nand U4722 (N_4722,N_4232,N_4353);
or U4723 (N_4723,N_4176,N_4294);
and U4724 (N_4724,N_4151,N_4408);
xor U4725 (N_4725,N_4257,N_4341);
nor U4726 (N_4726,N_4259,N_4318);
and U4727 (N_4727,N_4260,N_4227);
nor U4728 (N_4728,N_4263,N_4293);
and U4729 (N_4729,N_4078,N_4110);
xnor U4730 (N_4730,N_4079,N_4209);
or U4731 (N_4731,N_4113,N_4105);
nor U4732 (N_4732,N_4127,N_4450);
xor U4733 (N_4733,N_4147,N_4366);
and U4734 (N_4734,N_4192,N_4355);
xnor U4735 (N_4735,N_4344,N_4170);
and U4736 (N_4736,N_4141,N_4444);
and U4737 (N_4737,N_4106,N_4279);
nor U4738 (N_4738,N_4345,N_4398);
or U4739 (N_4739,N_4099,N_4321);
nand U4740 (N_4740,N_4007,N_4150);
nor U4741 (N_4741,N_4457,N_4336);
nand U4742 (N_4742,N_4281,N_4052);
nand U4743 (N_4743,N_4425,N_4410);
and U4744 (N_4744,N_4278,N_4097);
and U4745 (N_4745,N_4428,N_4406);
xor U4746 (N_4746,N_4399,N_4001);
or U4747 (N_4747,N_4264,N_4014);
or U4748 (N_4748,N_4413,N_4108);
xor U4749 (N_4749,N_4315,N_4480);
and U4750 (N_4750,N_4245,N_4167);
nand U4751 (N_4751,N_4325,N_4464);
nor U4752 (N_4752,N_4058,N_4308);
nand U4753 (N_4753,N_4234,N_4298);
and U4754 (N_4754,N_4460,N_4031);
nand U4755 (N_4755,N_4392,N_4356);
or U4756 (N_4756,N_4327,N_4330);
xor U4757 (N_4757,N_4024,N_4392);
nand U4758 (N_4758,N_4019,N_4449);
and U4759 (N_4759,N_4468,N_4325);
nor U4760 (N_4760,N_4025,N_4068);
nor U4761 (N_4761,N_4290,N_4128);
nor U4762 (N_4762,N_4044,N_4218);
xnor U4763 (N_4763,N_4475,N_4109);
nor U4764 (N_4764,N_4126,N_4428);
or U4765 (N_4765,N_4263,N_4215);
xnor U4766 (N_4766,N_4057,N_4341);
nor U4767 (N_4767,N_4065,N_4288);
and U4768 (N_4768,N_4039,N_4280);
or U4769 (N_4769,N_4150,N_4234);
xnor U4770 (N_4770,N_4116,N_4415);
and U4771 (N_4771,N_4373,N_4266);
or U4772 (N_4772,N_4036,N_4226);
and U4773 (N_4773,N_4344,N_4039);
xor U4774 (N_4774,N_4200,N_4477);
xnor U4775 (N_4775,N_4046,N_4220);
or U4776 (N_4776,N_4055,N_4448);
and U4777 (N_4777,N_4281,N_4440);
nand U4778 (N_4778,N_4090,N_4296);
nor U4779 (N_4779,N_4307,N_4439);
xnor U4780 (N_4780,N_4339,N_4256);
and U4781 (N_4781,N_4174,N_4055);
nor U4782 (N_4782,N_4380,N_4398);
nor U4783 (N_4783,N_4480,N_4332);
nor U4784 (N_4784,N_4388,N_4361);
and U4785 (N_4785,N_4183,N_4471);
nor U4786 (N_4786,N_4350,N_4290);
nor U4787 (N_4787,N_4405,N_4239);
and U4788 (N_4788,N_4295,N_4274);
nand U4789 (N_4789,N_4298,N_4247);
nand U4790 (N_4790,N_4119,N_4109);
nand U4791 (N_4791,N_4154,N_4287);
and U4792 (N_4792,N_4263,N_4094);
and U4793 (N_4793,N_4376,N_4492);
or U4794 (N_4794,N_4149,N_4165);
and U4795 (N_4795,N_4252,N_4446);
nand U4796 (N_4796,N_4040,N_4228);
and U4797 (N_4797,N_4038,N_4234);
xnor U4798 (N_4798,N_4105,N_4324);
or U4799 (N_4799,N_4415,N_4177);
nand U4800 (N_4800,N_4079,N_4463);
or U4801 (N_4801,N_4086,N_4363);
and U4802 (N_4802,N_4173,N_4490);
xnor U4803 (N_4803,N_4491,N_4012);
nand U4804 (N_4804,N_4239,N_4191);
nand U4805 (N_4805,N_4450,N_4067);
nor U4806 (N_4806,N_4299,N_4190);
xnor U4807 (N_4807,N_4390,N_4057);
and U4808 (N_4808,N_4342,N_4192);
nor U4809 (N_4809,N_4043,N_4131);
nand U4810 (N_4810,N_4465,N_4264);
or U4811 (N_4811,N_4040,N_4001);
and U4812 (N_4812,N_4153,N_4100);
nand U4813 (N_4813,N_4133,N_4467);
or U4814 (N_4814,N_4069,N_4479);
or U4815 (N_4815,N_4380,N_4254);
and U4816 (N_4816,N_4121,N_4437);
and U4817 (N_4817,N_4099,N_4312);
nor U4818 (N_4818,N_4137,N_4217);
nor U4819 (N_4819,N_4167,N_4021);
nor U4820 (N_4820,N_4444,N_4304);
or U4821 (N_4821,N_4219,N_4062);
nand U4822 (N_4822,N_4344,N_4340);
nand U4823 (N_4823,N_4334,N_4150);
xor U4824 (N_4824,N_4493,N_4096);
xnor U4825 (N_4825,N_4295,N_4272);
nor U4826 (N_4826,N_4360,N_4102);
xor U4827 (N_4827,N_4379,N_4290);
xor U4828 (N_4828,N_4052,N_4481);
nand U4829 (N_4829,N_4197,N_4316);
and U4830 (N_4830,N_4169,N_4443);
nor U4831 (N_4831,N_4278,N_4221);
nand U4832 (N_4832,N_4365,N_4067);
nor U4833 (N_4833,N_4206,N_4048);
nand U4834 (N_4834,N_4365,N_4447);
and U4835 (N_4835,N_4296,N_4391);
and U4836 (N_4836,N_4361,N_4287);
or U4837 (N_4837,N_4285,N_4081);
nor U4838 (N_4838,N_4201,N_4203);
and U4839 (N_4839,N_4373,N_4228);
and U4840 (N_4840,N_4415,N_4386);
or U4841 (N_4841,N_4360,N_4426);
xor U4842 (N_4842,N_4304,N_4473);
and U4843 (N_4843,N_4073,N_4254);
nor U4844 (N_4844,N_4205,N_4068);
or U4845 (N_4845,N_4060,N_4030);
and U4846 (N_4846,N_4308,N_4152);
xnor U4847 (N_4847,N_4149,N_4415);
and U4848 (N_4848,N_4338,N_4296);
nand U4849 (N_4849,N_4217,N_4262);
xnor U4850 (N_4850,N_4423,N_4279);
xnor U4851 (N_4851,N_4218,N_4119);
or U4852 (N_4852,N_4275,N_4348);
or U4853 (N_4853,N_4284,N_4118);
xor U4854 (N_4854,N_4480,N_4108);
xor U4855 (N_4855,N_4458,N_4230);
xor U4856 (N_4856,N_4057,N_4250);
or U4857 (N_4857,N_4079,N_4297);
nor U4858 (N_4858,N_4310,N_4344);
and U4859 (N_4859,N_4002,N_4054);
nand U4860 (N_4860,N_4045,N_4496);
nand U4861 (N_4861,N_4463,N_4477);
xnor U4862 (N_4862,N_4371,N_4408);
xor U4863 (N_4863,N_4262,N_4344);
xor U4864 (N_4864,N_4377,N_4229);
nor U4865 (N_4865,N_4462,N_4028);
and U4866 (N_4866,N_4287,N_4122);
nand U4867 (N_4867,N_4264,N_4163);
or U4868 (N_4868,N_4106,N_4405);
or U4869 (N_4869,N_4117,N_4107);
nand U4870 (N_4870,N_4498,N_4190);
xnor U4871 (N_4871,N_4272,N_4437);
nand U4872 (N_4872,N_4006,N_4202);
nand U4873 (N_4873,N_4340,N_4132);
nor U4874 (N_4874,N_4414,N_4481);
xnor U4875 (N_4875,N_4238,N_4303);
xnor U4876 (N_4876,N_4078,N_4492);
xor U4877 (N_4877,N_4251,N_4012);
nand U4878 (N_4878,N_4220,N_4179);
or U4879 (N_4879,N_4210,N_4151);
or U4880 (N_4880,N_4218,N_4426);
nor U4881 (N_4881,N_4147,N_4263);
nor U4882 (N_4882,N_4189,N_4427);
xor U4883 (N_4883,N_4230,N_4210);
and U4884 (N_4884,N_4441,N_4311);
or U4885 (N_4885,N_4338,N_4051);
nand U4886 (N_4886,N_4052,N_4261);
nor U4887 (N_4887,N_4188,N_4233);
nor U4888 (N_4888,N_4248,N_4173);
xor U4889 (N_4889,N_4199,N_4172);
xor U4890 (N_4890,N_4335,N_4472);
or U4891 (N_4891,N_4023,N_4343);
and U4892 (N_4892,N_4352,N_4149);
or U4893 (N_4893,N_4063,N_4253);
nand U4894 (N_4894,N_4010,N_4491);
nand U4895 (N_4895,N_4031,N_4278);
or U4896 (N_4896,N_4015,N_4414);
nand U4897 (N_4897,N_4006,N_4236);
or U4898 (N_4898,N_4254,N_4427);
nand U4899 (N_4899,N_4464,N_4252);
and U4900 (N_4900,N_4004,N_4250);
nand U4901 (N_4901,N_4413,N_4372);
nor U4902 (N_4902,N_4203,N_4294);
nand U4903 (N_4903,N_4018,N_4161);
and U4904 (N_4904,N_4059,N_4069);
nand U4905 (N_4905,N_4301,N_4442);
nor U4906 (N_4906,N_4312,N_4394);
nand U4907 (N_4907,N_4147,N_4303);
or U4908 (N_4908,N_4061,N_4208);
nor U4909 (N_4909,N_4349,N_4203);
nor U4910 (N_4910,N_4442,N_4081);
and U4911 (N_4911,N_4479,N_4446);
and U4912 (N_4912,N_4218,N_4329);
xor U4913 (N_4913,N_4425,N_4218);
xor U4914 (N_4914,N_4147,N_4112);
and U4915 (N_4915,N_4376,N_4386);
xnor U4916 (N_4916,N_4312,N_4477);
and U4917 (N_4917,N_4393,N_4023);
and U4918 (N_4918,N_4087,N_4345);
nand U4919 (N_4919,N_4354,N_4135);
nand U4920 (N_4920,N_4230,N_4396);
or U4921 (N_4921,N_4429,N_4001);
xor U4922 (N_4922,N_4125,N_4347);
nand U4923 (N_4923,N_4419,N_4343);
nand U4924 (N_4924,N_4140,N_4381);
nor U4925 (N_4925,N_4369,N_4486);
and U4926 (N_4926,N_4274,N_4172);
and U4927 (N_4927,N_4205,N_4428);
nor U4928 (N_4928,N_4473,N_4000);
nand U4929 (N_4929,N_4289,N_4329);
or U4930 (N_4930,N_4141,N_4095);
and U4931 (N_4931,N_4051,N_4440);
or U4932 (N_4932,N_4132,N_4446);
xor U4933 (N_4933,N_4216,N_4269);
and U4934 (N_4934,N_4273,N_4461);
and U4935 (N_4935,N_4199,N_4113);
nor U4936 (N_4936,N_4256,N_4187);
nor U4937 (N_4937,N_4192,N_4013);
and U4938 (N_4938,N_4322,N_4256);
nand U4939 (N_4939,N_4157,N_4409);
xnor U4940 (N_4940,N_4274,N_4048);
or U4941 (N_4941,N_4385,N_4439);
and U4942 (N_4942,N_4217,N_4364);
or U4943 (N_4943,N_4072,N_4452);
nor U4944 (N_4944,N_4482,N_4458);
and U4945 (N_4945,N_4420,N_4045);
or U4946 (N_4946,N_4197,N_4062);
xnor U4947 (N_4947,N_4474,N_4054);
or U4948 (N_4948,N_4496,N_4057);
or U4949 (N_4949,N_4156,N_4191);
or U4950 (N_4950,N_4328,N_4392);
xnor U4951 (N_4951,N_4252,N_4206);
xnor U4952 (N_4952,N_4322,N_4105);
and U4953 (N_4953,N_4384,N_4273);
or U4954 (N_4954,N_4326,N_4348);
nor U4955 (N_4955,N_4359,N_4376);
or U4956 (N_4956,N_4208,N_4198);
and U4957 (N_4957,N_4020,N_4494);
nand U4958 (N_4958,N_4282,N_4308);
and U4959 (N_4959,N_4341,N_4260);
xnor U4960 (N_4960,N_4035,N_4037);
and U4961 (N_4961,N_4120,N_4373);
nor U4962 (N_4962,N_4412,N_4109);
or U4963 (N_4963,N_4367,N_4190);
nand U4964 (N_4964,N_4194,N_4481);
nor U4965 (N_4965,N_4126,N_4019);
or U4966 (N_4966,N_4363,N_4423);
or U4967 (N_4967,N_4288,N_4319);
nand U4968 (N_4968,N_4165,N_4181);
xnor U4969 (N_4969,N_4048,N_4384);
xnor U4970 (N_4970,N_4494,N_4314);
nand U4971 (N_4971,N_4190,N_4001);
nand U4972 (N_4972,N_4110,N_4226);
or U4973 (N_4973,N_4426,N_4176);
and U4974 (N_4974,N_4295,N_4293);
and U4975 (N_4975,N_4239,N_4103);
nor U4976 (N_4976,N_4452,N_4301);
xnor U4977 (N_4977,N_4049,N_4214);
or U4978 (N_4978,N_4200,N_4128);
or U4979 (N_4979,N_4139,N_4460);
xnor U4980 (N_4980,N_4195,N_4337);
and U4981 (N_4981,N_4159,N_4491);
and U4982 (N_4982,N_4306,N_4216);
nand U4983 (N_4983,N_4264,N_4316);
nand U4984 (N_4984,N_4257,N_4295);
nand U4985 (N_4985,N_4051,N_4111);
or U4986 (N_4986,N_4089,N_4289);
and U4987 (N_4987,N_4050,N_4017);
xor U4988 (N_4988,N_4315,N_4202);
nand U4989 (N_4989,N_4181,N_4393);
nand U4990 (N_4990,N_4151,N_4260);
nand U4991 (N_4991,N_4127,N_4184);
or U4992 (N_4992,N_4054,N_4440);
and U4993 (N_4993,N_4233,N_4406);
or U4994 (N_4994,N_4294,N_4328);
or U4995 (N_4995,N_4357,N_4070);
xnor U4996 (N_4996,N_4364,N_4129);
or U4997 (N_4997,N_4273,N_4355);
or U4998 (N_4998,N_4140,N_4319);
or U4999 (N_4999,N_4139,N_4035);
nand U5000 (N_5000,N_4833,N_4558);
nor U5001 (N_5001,N_4592,N_4873);
nand U5002 (N_5002,N_4756,N_4682);
or U5003 (N_5003,N_4965,N_4759);
or U5004 (N_5004,N_4565,N_4834);
xnor U5005 (N_5005,N_4802,N_4821);
or U5006 (N_5006,N_4786,N_4654);
xnor U5007 (N_5007,N_4712,N_4905);
xnor U5008 (N_5008,N_4723,N_4947);
nand U5009 (N_5009,N_4711,N_4553);
nand U5010 (N_5010,N_4622,N_4569);
nor U5011 (N_5011,N_4754,N_4710);
and U5012 (N_5012,N_4840,N_4535);
and U5013 (N_5013,N_4640,N_4696);
and U5014 (N_5014,N_4828,N_4740);
nor U5015 (N_5015,N_4531,N_4987);
nor U5016 (N_5016,N_4566,N_4601);
or U5017 (N_5017,N_4637,N_4581);
nand U5018 (N_5018,N_4559,N_4706);
or U5019 (N_5019,N_4629,N_4670);
xnor U5020 (N_5020,N_4609,N_4934);
or U5021 (N_5021,N_4877,N_4746);
and U5022 (N_5022,N_4839,N_4530);
or U5023 (N_5023,N_4634,N_4509);
or U5024 (N_5024,N_4832,N_4971);
xor U5025 (N_5025,N_4969,N_4763);
nand U5026 (N_5026,N_4510,N_4924);
and U5027 (N_5027,N_4577,N_4517);
and U5028 (N_5028,N_4861,N_4527);
nand U5029 (N_5029,N_4796,N_4625);
nor U5030 (N_5030,N_4812,N_4819);
or U5031 (N_5031,N_4643,N_4894);
or U5032 (N_5032,N_4513,N_4518);
or U5033 (N_5033,N_4881,N_4829);
nand U5034 (N_5034,N_4809,N_4998);
nand U5035 (N_5035,N_4695,N_4820);
or U5036 (N_5036,N_4739,N_4899);
nand U5037 (N_5037,N_4795,N_4727);
or U5038 (N_5038,N_4742,N_4792);
nor U5039 (N_5039,N_4946,N_4794);
nor U5040 (N_5040,N_4658,N_4758);
and U5041 (N_5041,N_4891,N_4850);
and U5042 (N_5042,N_4648,N_4836);
xor U5043 (N_5043,N_4661,N_4719);
nand U5044 (N_5044,N_4816,N_4540);
nor U5045 (N_5045,N_4608,N_4551);
or U5046 (N_5046,N_4798,N_4731);
or U5047 (N_5047,N_4961,N_4726);
xor U5048 (N_5048,N_4503,N_4656);
xor U5049 (N_5049,N_4584,N_4514);
nand U5050 (N_5050,N_4979,N_4589);
xnor U5051 (N_5051,N_4564,N_4898);
xor U5052 (N_5052,N_4882,N_4767);
nor U5053 (N_5053,N_4659,N_4966);
nand U5054 (N_5054,N_4732,N_4957);
and U5055 (N_5055,N_4849,N_4766);
xor U5056 (N_5056,N_4871,N_4649);
and U5057 (N_5057,N_4920,N_4826);
nor U5058 (N_5058,N_4642,N_4962);
xnor U5059 (N_5059,N_4932,N_4691);
xnor U5060 (N_5060,N_4978,N_4500);
and U5061 (N_5061,N_4782,N_4800);
or U5062 (N_5062,N_4702,N_4557);
nand U5063 (N_5063,N_4853,N_4940);
nor U5064 (N_5064,N_4542,N_4990);
or U5065 (N_5065,N_4699,N_4674);
or U5066 (N_5066,N_4543,N_4997);
and U5067 (N_5067,N_4597,N_4607);
nor U5068 (N_5068,N_4799,N_4679);
nand U5069 (N_5069,N_4952,N_4512);
and U5070 (N_5070,N_4573,N_4628);
nor U5071 (N_5071,N_4841,N_4830);
xor U5072 (N_5072,N_4626,N_4996);
nor U5073 (N_5073,N_4912,N_4842);
and U5074 (N_5074,N_4753,N_4835);
and U5075 (N_5075,N_4669,N_4817);
nand U5076 (N_5076,N_4874,N_4526);
xnor U5077 (N_5077,N_4694,N_4621);
and U5078 (N_5078,N_4580,N_4908);
and U5079 (N_5079,N_4730,N_4568);
nor U5080 (N_5080,N_4775,N_4744);
xor U5081 (N_5081,N_4970,N_4595);
or U5082 (N_5082,N_4761,N_4505);
nor U5083 (N_5083,N_4982,N_4715);
or U5084 (N_5084,N_4603,N_4806);
nor U5085 (N_5085,N_4883,N_4537);
nor U5086 (N_5086,N_4552,N_4975);
or U5087 (N_5087,N_4964,N_4837);
nor U5088 (N_5088,N_4716,N_4684);
xor U5089 (N_5089,N_4630,N_4714);
nand U5090 (N_5090,N_4522,N_4504);
or U5091 (N_5091,N_4973,N_4534);
and U5092 (N_5092,N_4538,N_4765);
and U5093 (N_5093,N_4937,N_4536);
nand U5094 (N_5094,N_4751,N_4879);
nor U5095 (N_5095,N_4797,N_4993);
and U5096 (N_5096,N_4728,N_4989);
nor U5097 (N_5097,N_4617,N_4638);
nand U5098 (N_5098,N_4651,N_4635);
xor U5099 (N_5099,N_4749,N_4612);
nor U5100 (N_5100,N_4664,N_4515);
nor U5101 (N_5101,N_4539,N_4680);
nand U5102 (N_5102,N_4914,N_4668);
nand U5103 (N_5103,N_4523,N_4843);
nand U5104 (N_5104,N_4945,N_4532);
xor U5105 (N_5105,N_4783,N_4951);
nor U5106 (N_5106,N_4662,N_4867);
xor U5107 (N_5107,N_4547,N_4824);
nand U5108 (N_5108,N_4949,N_4771);
or U5109 (N_5109,N_4655,N_4582);
xor U5110 (N_5110,N_4926,N_4687);
and U5111 (N_5111,N_4610,N_4616);
nor U5112 (N_5112,N_4752,N_4698);
and U5113 (N_5113,N_4546,N_4585);
and U5114 (N_5114,N_4933,N_4735);
nand U5115 (N_5115,N_4521,N_4560);
nand U5116 (N_5116,N_4992,N_4645);
nor U5117 (N_5117,N_4893,N_4845);
nand U5118 (N_5118,N_4789,N_4942);
or U5119 (N_5119,N_4922,N_4941);
xor U5120 (N_5120,N_4929,N_4895);
and U5121 (N_5121,N_4676,N_4620);
and U5122 (N_5122,N_4683,N_4697);
xor U5123 (N_5123,N_4921,N_4672);
xor U5124 (N_5124,N_4639,N_4653);
xnor U5125 (N_5125,N_4738,N_4903);
nor U5126 (N_5126,N_4575,N_4562);
xnor U5127 (N_5127,N_4686,N_4884);
nand U5128 (N_5128,N_4692,N_4856);
nand U5129 (N_5129,N_4600,N_4598);
xnor U5130 (N_5130,N_4950,N_4844);
xnor U5131 (N_5131,N_4769,N_4704);
nor U5132 (N_5132,N_4803,N_4948);
or U5133 (N_5133,N_4613,N_4804);
or U5134 (N_5134,N_4611,N_4596);
and U5135 (N_5135,N_4707,N_4848);
nor U5136 (N_5136,N_4958,N_4980);
or U5137 (N_5137,N_4915,N_4541);
nand U5138 (N_5138,N_4713,N_4918);
and U5139 (N_5139,N_4868,N_4745);
and U5140 (N_5140,N_4548,N_4801);
xnor U5141 (N_5141,N_4519,N_4827);
and U5142 (N_5142,N_4590,N_4737);
xnor U5143 (N_5143,N_4693,N_4785);
and U5144 (N_5144,N_4857,N_4507);
nor U5145 (N_5145,N_4793,N_4623);
xnor U5146 (N_5146,N_4708,N_4703);
nor U5147 (N_5147,N_4994,N_4591);
or U5148 (N_5148,N_4846,N_4570);
or U5149 (N_5149,N_4773,N_4864);
nor U5150 (N_5150,N_4561,N_4677);
or U5151 (N_5151,N_4917,N_4520);
or U5152 (N_5152,N_4901,N_4675);
and U5153 (N_5153,N_4619,N_4866);
and U5154 (N_5154,N_4902,N_4574);
nor U5155 (N_5155,N_4847,N_4885);
xnor U5156 (N_5156,N_4762,N_4855);
nand U5157 (N_5157,N_4776,N_4784);
nand U5158 (N_5158,N_4974,N_4927);
nand U5159 (N_5159,N_4823,N_4939);
nand U5160 (N_5160,N_4681,N_4913);
nand U5161 (N_5161,N_4916,N_4545);
nor U5162 (N_5162,N_4631,N_4814);
and U5163 (N_5163,N_4572,N_4831);
xor U5164 (N_5164,N_4606,N_4909);
nand U5165 (N_5165,N_4750,N_4741);
nand U5166 (N_5166,N_4859,N_4647);
nand U5167 (N_5167,N_4760,N_4602);
or U5168 (N_5168,N_4646,N_4944);
nor U5169 (N_5169,N_4890,N_4660);
or U5170 (N_5170,N_4747,N_4632);
xor U5171 (N_5171,N_4936,N_4636);
nand U5172 (N_5172,N_4910,N_4860);
and U5173 (N_5173,N_4550,N_4778);
nor U5174 (N_5174,N_4624,N_4709);
nand U5175 (N_5175,N_4985,N_4734);
xor U5176 (N_5176,N_4671,N_4981);
or U5177 (N_5177,N_4615,N_4721);
xnor U5178 (N_5178,N_4906,N_4960);
and U5179 (N_5179,N_4907,N_4586);
and U5180 (N_5180,N_4991,N_4854);
nor U5181 (N_5181,N_4822,N_4983);
and U5182 (N_5182,N_4583,N_4599);
nand U5183 (N_5183,N_4928,N_4665);
nand U5184 (N_5184,N_4666,N_4529);
and U5185 (N_5185,N_4544,N_4876);
or U5186 (N_5186,N_4862,N_4614);
and U5187 (N_5187,N_4777,N_4579);
and U5188 (N_5188,N_4787,N_4689);
xnor U5189 (N_5189,N_4650,N_4768);
or U5190 (N_5190,N_4511,N_4722);
or U5191 (N_5191,N_4549,N_4688);
xor U5192 (N_5192,N_4720,N_4725);
xnor U5193 (N_5193,N_4919,N_4815);
xor U5194 (N_5194,N_4995,N_4959);
nand U5195 (N_5195,N_4525,N_4892);
nor U5196 (N_5196,N_4588,N_4641);
nand U5197 (N_5197,N_4851,N_4972);
xnor U5198 (N_5198,N_4900,N_4911);
xnor U5199 (N_5199,N_4880,N_4984);
xnor U5200 (N_5200,N_4717,N_4808);
and U5201 (N_5201,N_4633,N_4930);
and U5202 (N_5202,N_4988,N_4805);
and U5203 (N_5203,N_4506,N_4685);
nor U5204 (N_5204,N_4652,N_4774);
and U5205 (N_5205,N_4764,N_4724);
nor U5206 (N_5206,N_4556,N_4571);
and U5207 (N_5207,N_4889,N_4878);
xor U5208 (N_5208,N_4770,N_4938);
nor U5209 (N_5209,N_4818,N_4502);
or U5210 (N_5210,N_4999,N_4858);
xor U5211 (N_5211,N_4963,N_4508);
nor U5212 (N_5212,N_4678,N_4955);
xnor U5213 (N_5213,N_4516,N_4886);
nand U5214 (N_5214,N_4594,N_4705);
nand U5215 (N_5215,N_4733,N_4852);
xor U5216 (N_5216,N_4605,N_4729);
nor U5217 (N_5217,N_4618,N_4810);
nor U5218 (N_5218,N_4870,N_4743);
and U5219 (N_5219,N_4567,N_4604);
or U5220 (N_5220,N_4931,N_4807);
or U5221 (N_5221,N_4813,N_4825);
nor U5222 (N_5222,N_4555,N_4790);
nand U5223 (N_5223,N_4953,N_4968);
or U5224 (N_5224,N_4501,N_4736);
nor U5225 (N_5225,N_4863,N_4967);
or U5226 (N_5226,N_4627,N_4875);
and U5227 (N_5227,N_4838,N_4667);
nand U5228 (N_5228,N_4673,N_4977);
nand U5229 (N_5229,N_4888,N_4897);
xor U5230 (N_5230,N_4663,N_4976);
nor U5231 (N_5231,N_4811,N_4700);
or U5232 (N_5232,N_4657,N_4718);
nor U5233 (N_5233,N_4956,N_4925);
and U5234 (N_5234,N_4780,N_4748);
xor U5235 (N_5235,N_4587,N_4869);
xnor U5236 (N_5236,N_4954,N_4524);
nand U5237 (N_5237,N_4923,N_4593);
and U5238 (N_5238,N_4644,N_4872);
or U5239 (N_5239,N_4701,N_4865);
nand U5240 (N_5240,N_4554,N_4779);
xor U5241 (N_5241,N_4690,N_4887);
nor U5242 (N_5242,N_4781,N_4772);
nand U5243 (N_5243,N_4943,N_4578);
nor U5244 (N_5244,N_4757,N_4986);
xnor U5245 (N_5245,N_4896,N_4791);
xor U5246 (N_5246,N_4563,N_4935);
nor U5247 (N_5247,N_4528,N_4755);
nor U5248 (N_5248,N_4788,N_4904);
or U5249 (N_5249,N_4576,N_4533);
nand U5250 (N_5250,N_4935,N_4839);
xor U5251 (N_5251,N_4712,N_4619);
nor U5252 (N_5252,N_4865,N_4671);
nor U5253 (N_5253,N_4552,N_4751);
or U5254 (N_5254,N_4909,N_4695);
and U5255 (N_5255,N_4534,N_4568);
nand U5256 (N_5256,N_4699,N_4988);
nand U5257 (N_5257,N_4907,N_4793);
and U5258 (N_5258,N_4976,N_4773);
xor U5259 (N_5259,N_4935,N_4803);
nor U5260 (N_5260,N_4652,N_4516);
nand U5261 (N_5261,N_4755,N_4968);
nand U5262 (N_5262,N_4955,N_4847);
xnor U5263 (N_5263,N_4803,N_4807);
nand U5264 (N_5264,N_4674,N_4867);
or U5265 (N_5265,N_4943,N_4884);
nand U5266 (N_5266,N_4592,N_4665);
xnor U5267 (N_5267,N_4865,N_4623);
and U5268 (N_5268,N_4846,N_4569);
xnor U5269 (N_5269,N_4889,N_4528);
and U5270 (N_5270,N_4825,N_4809);
and U5271 (N_5271,N_4519,N_4887);
or U5272 (N_5272,N_4572,N_4855);
nor U5273 (N_5273,N_4898,N_4608);
xor U5274 (N_5274,N_4835,N_4720);
nand U5275 (N_5275,N_4570,N_4901);
xnor U5276 (N_5276,N_4688,N_4856);
nand U5277 (N_5277,N_4773,N_4690);
xnor U5278 (N_5278,N_4771,N_4845);
xor U5279 (N_5279,N_4744,N_4612);
nor U5280 (N_5280,N_4918,N_4818);
nor U5281 (N_5281,N_4978,N_4879);
nand U5282 (N_5282,N_4800,N_4734);
nand U5283 (N_5283,N_4550,N_4791);
nand U5284 (N_5284,N_4644,N_4624);
nor U5285 (N_5285,N_4936,N_4854);
and U5286 (N_5286,N_4788,N_4839);
nor U5287 (N_5287,N_4826,N_4528);
xnor U5288 (N_5288,N_4946,N_4908);
or U5289 (N_5289,N_4884,N_4832);
and U5290 (N_5290,N_4804,N_4955);
nand U5291 (N_5291,N_4999,N_4668);
and U5292 (N_5292,N_4988,N_4912);
nand U5293 (N_5293,N_4923,N_4767);
nor U5294 (N_5294,N_4559,N_4582);
and U5295 (N_5295,N_4894,N_4541);
xor U5296 (N_5296,N_4699,N_4740);
or U5297 (N_5297,N_4796,N_4799);
or U5298 (N_5298,N_4753,N_4762);
xor U5299 (N_5299,N_4786,N_4956);
nand U5300 (N_5300,N_4541,N_4619);
nor U5301 (N_5301,N_4989,N_4761);
nand U5302 (N_5302,N_4660,N_4621);
nand U5303 (N_5303,N_4785,N_4863);
xor U5304 (N_5304,N_4705,N_4579);
or U5305 (N_5305,N_4517,N_4523);
nor U5306 (N_5306,N_4653,N_4866);
xor U5307 (N_5307,N_4873,N_4726);
or U5308 (N_5308,N_4894,N_4805);
nand U5309 (N_5309,N_4916,N_4558);
or U5310 (N_5310,N_4990,N_4763);
nor U5311 (N_5311,N_4792,N_4506);
and U5312 (N_5312,N_4668,N_4683);
xor U5313 (N_5313,N_4795,N_4602);
nor U5314 (N_5314,N_4776,N_4736);
nor U5315 (N_5315,N_4657,N_4593);
nand U5316 (N_5316,N_4912,N_4679);
and U5317 (N_5317,N_4865,N_4891);
or U5318 (N_5318,N_4902,N_4712);
or U5319 (N_5319,N_4876,N_4866);
nor U5320 (N_5320,N_4791,N_4564);
nand U5321 (N_5321,N_4963,N_4977);
or U5322 (N_5322,N_4747,N_4964);
xor U5323 (N_5323,N_4685,N_4532);
xor U5324 (N_5324,N_4912,N_4853);
xnor U5325 (N_5325,N_4692,N_4610);
nand U5326 (N_5326,N_4513,N_4582);
and U5327 (N_5327,N_4582,N_4660);
nand U5328 (N_5328,N_4790,N_4928);
xnor U5329 (N_5329,N_4573,N_4585);
or U5330 (N_5330,N_4935,N_4663);
or U5331 (N_5331,N_4752,N_4778);
and U5332 (N_5332,N_4612,N_4616);
and U5333 (N_5333,N_4585,N_4741);
or U5334 (N_5334,N_4822,N_4716);
or U5335 (N_5335,N_4545,N_4650);
nand U5336 (N_5336,N_4592,N_4986);
nor U5337 (N_5337,N_4517,N_4622);
nor U5338 (N_5338,N_4581,N_4690);
and U5339 (N_5339,N_4985,N_4732);
or U5340 (N_5340,N_4660,N_4697);
nand U5341 (N_5341,N_4997,N_4652);
nand U5342 (N_5342,N_4564,N_4571);
xor U5343 (N_5343,N_4541,N_4941);
and U5344 (N_5344,N_4838,N_4708);
xnor U5345 (N_5345,N_4977,N_4924);
and U5346 (N_5346,N_4934,N_4966);
xnor U5347 (N_5347,N_4754,N_4937);
nand U5348 (N_5348,N_4739,N_4762);
or U5349 (N_5349,N_4829,N_4766);
nand U5350 (N_5350,N_4730,N_4824);
nor U5351 (N_5351,N_4539,N_4669);
nand U5352 (N_5352,N_4999,N_4609);
xnor U5353 (N_5353,N_4751,N_4559);
xor U5354 (N_5354,N_4969,N_4649);
nand U5355 (N_5355,N_4940,N_4954);
nand U5356 (N_5356,N_4506,N_4666);
and U5357 (N_5357,N_4649,N_4831);
and U5358 (N_5358,N_4833,N_4703);
nor U5359 (N_5359,N_4641,N_4508);
nand U5360 (N_5360,N_4903,N_4841);
xnor U5361 (N_5361,N_4985,N_4547);
xnor U5362 (N_5362,N_4640,N_4758);
and U5363 (N_5363,N_4964,N_4821);
nand U5364 (N_5364,N_4793,N_4926);
and U5365 (N_5365,N_4727,N_4758);
nor U5366 (N_5366,N_4553,N_4799);
nand U5367 (N_5367,N_4806,N_4593);
nor U5368 (N_5368,N_4821,N_4908);
and U5369 (N_5369,N_4700,N_4547);
or U5370 (N_5370,N_4774,N_4817);
xor U5371 (N_5371,N_4725,N_4912);
xnor U5372 (N_5372,N_4547,N_4641);
or U5373 (N_5373,N_4550,N_4600);
nand U5374 (N_5374,N_4816,N_4649);
nor U5375 (N_5375,N_4953,N_4518);
xor U5376 (N_5376,N_4789,N_4962);
or U5377 (N_5377,N_4836,N_4860);
nand U5378 (N_5378,N_4959,N_4993);
and U5379 (N_5379,N_4573,N_4779);
nand U5380 (N_5380,N_4512,N_4671);
nor U5381 (N_5381,N_4551,N_4822);
nor U5382 (N_5382,N_4985,N_4798);
nand U5383 (N_5383,N_4663,N_4635);
nor U5384 (N_5384,N_4724,N_4851);
xnor U5385 (N_5385,N_4531,N_4962);
or U5386 (N_5386,N_4593,N_4938);
and U5387 (N_5387,N_4954,N_4851);
and U5388 (N_5388,N_4997,N_4772);
or U5389 (N_5389,N_4503,N_4513);
and U5390 (N_5390,N_4978,N_4764);
and U5391 (N_5391,N_4544,N_4972);
xor U5392 (N_5392,N_4762,N_4680);
and U5393 (N_5393,N_4789,N_4912);
or U5394 (N_5394,N_4857,N_4820);
nor U5395 (N_5395,N_4793,N_4695);
and U5396 (N_5396,N_4913,N_4615);
and U5397 (N_5397,N_4755,N_4704);
and U5398 (N_5398,N_4647,N_4640);
nor U5399 (N_5399,N_4574,N_4741);
and U5400 (N_5400,N_4662,N_4817);
xor U5401 (N_5401,N_4528,N_4604);
and U5402 (N_5402,N_4987,N_4522);
nor U5403 (N_5403,N_4712,N_4633);
nand U5404 (N_5404,N_4780,N_4747);
nor U5405 (N_5405,N_4762,N_4851);
nor U5406 (N_5406,N_4737,N_4867);
xnor U5407 (N_5407,N_4667,N_4846);
nor U5408 (N_5408,N_4768,N_4951);
xor U5409 (N_5409,N_4967,N_4935);
nor U5410 (N_5410,N_4598,N_4964);
nor U5411 (N_5411,N_4682,N_4932);
nand U5412 (N_5412,N_4798,N_4923);
or U5413 (N_5413,N_4618,N_4667);
and U5414 (N_5414,N_4646,N_4720);
nor U5415 (N_5415,N_4972,N_4651);
or U5416 (N_5416,N_4628,N_4500);
or U5417 (N_5417,N_4897,N_4853);
nor U5418 (N_5418,N_4664,N_4764);
and U5419 (N_5419,N_4975,N_4825);
nor U5420 (N_5420,N_4731,N_4802);
nand U5421 (N_5421,N_4934,N_4606);
and U5422 (N_5422,N_4789,N_4535);
xnor U5423 (N_5423,N_4547,N_4947);
nand U5424 (N_5424,N_4594,N_4709);
and U5425 (N_5425,N_4725,N_4599);
nor U5426 (N_5426,N_4731,N_4734);
xnor U5427 (N_5427,N_4623,N_4701);
nand U5428 (N_5428,N_4542,N_4809);
nand U5429 (N_5429,N_4678,N_4989);
xnor U5430 (N_5430,N_4511,N_4833);
nand U5431 (N_5431,N_4785,N_4659);
or U5432 (N_5432,N_4589,N_4641);
xnor U5433 (N_5433,N_4958,N_4585);
and U5434 (N_5434,N_4833,N_4961);
and U5435 (N_5435,N_4768,N_4816);
nor U5436 (N_5436,N_4618,N_4555);
xnor U5437 (N_5437,N_4691,N_4593);
nor U5438 (N_5438,N_4601,N_4791);
nor U5439 (N_5439,N_4687,N_4577);
and U5440 (N_5440,N_4609,N_4671);
xor U5441 (N_5441,N_4840,N_4835);
xor U5442 (N_5442,N_4694,N_4859);
nand U5443 (N_5443,N_4773,N_4972);
nor U5444 (N_5444,N_4751,N_4697);
xnor U5445 (N_5445,N_4515,N_4554);
nor U5446 (N_5446,N_4892,N_4540);
xnor U5447 (N_5447,N_4750,N_4814);
nand U5448 (N_5448,N_4516,N_4918);
nor U5449 (N_5449,N_4580,N_4590);
and U5450 (N_5450,N_4781,N_4522);
nor U5451 (N_5451,N_4794,N_4971);
nor U5452 (N_5452,N_4662,N_4758);
or U5453 (N_5453,N_4838,N_4643);
nor U5454 (N_5454,N_4668,N_4852);
xnor U5455 (N_5455,N_4824,N_4524);
xor U5456 (N_5456,N_4732,N_4866);
and U5457 (N_5457,N_4792,N_4682);
xor U5458 (N_5458,N_4875,N_4578);
or U5459 (N_5459,N_4638,N_4922);
xor U5460 (N_5460,N_4656,N_4897);
nor U5461 (N_5461,N_4667,N_4890);
xnor U5462 (N_5462,N_4968,N_4881);
and U5463 (N_5463,N_4508,N_4550);
nor U5464 (N_5464,N_4784,N_4610);
and U5465 (N_5465,N_4940,N_4666);
nand U5466 (N_5466,N_4844,N_4727);
nand U5467 (N_5467,N_4810,N_4667);
xor U5468 (N_5468,N_4525,N_4613);
and U5469 (N_5469,N_4565,N_4665);
or U5470 (N_5470,N_4776,N_4577);
nor U5471 (N_5471,N_4650,N_4660);
xnor U5472 (N_5472,N_4844,N_4593);
or U5473 (N_5473,N_4653,N_4641);
or U5474 (N_5474,N_4615,N_4825);
or U5475 (N_5475,N_4836,N_4615);
and U5476 (N_5476,N_4750,N_4677);
nor U5477 (N_5477,N_4652,N_4625);
xnor U5478 (N_5478,N_4565,N_4881);
nand U5479 (N_5479,N_4876,N_4529);
or U5480 (N_5480,N_4596,N_4646);
xor U5481 (N_5481,N_4802,N_4633);
and U5482 (N_5482,N_4750,N_4984);
or U5483 (N_5483,N_4887,N_4763);
nor U5484 (N_5484,N_4865,N_4593);
xnor U5485 (N_5485,N_4563,N_4789);
and U5486 (N_5486,N_4721,N_4929);
nand U5487 (N_5487,N_4860,N_4759);
and U5488 (N_5488,N_4892,N_4859);
or U5489 (N_5489,N_4606,N_4710);
or U5490 (N_5490,N_4901,N_4983);
or U5491 (N_5491,N_4835,N_4709);
and U5492 (N_5492,N_4828,N_4979);
and U5493 (N_5493,N_4748,N_4553);
xor U5494 (N_5494,N_4823,N_4627);
xor U5495 (N_5495,N_4886,N_4996);
xor U5496 (N_5496,N_4512,N_4975);
nand U5497 (N_5497,N_4875,N_4611);
nand U5498 (N_5498,N_4826,N_4730);
xor U5499 (N_5499,N_4936,N_4745);
nand U5500 (N_5500,N_5075,N_5237);
xor U5501 (N_5501,N_5066,N_5063);
xor U5502 (N_5502,N_5422,N_5133);
and U5503 (N_5503,N_5445,N_5331);
nor U5504 (N_5504,N_5395,N_5114);
nand U5505 (N_5505,N_5052,N_5396);
nor U5506 (N_5506,N_5421,N_5007);
xnor U5507 (N_5507,N_5130,N_5105);
or U5508 (N_5508,N_5429,N_5324);
xor U5509 (N_5509,N_5458,N_5224);
nand U5510 (N_5510,N_5243,N_5062);
nor U5511 (N_5511,N_5298,N_5081);
xnor U5512 (N_5512,N_5313,N_5356);
nand U5513 (N_5513,N_5078,N_5368);
nand U5514 (N_5514,N_5202,N_5467);
nor U5515 (N_5515,N_5154,N_5360);
or U5516 (N_5516,N_5046,N_5328);
or U5517 (N_5517,N_5333,N_5115);
or U5518 (N_5518,N_5284,N_5199);
and U5519 (N_5519,N_5000,N_5307);
nand U5520 (N_5520,N_5264,N_5393);
nand U5521 (N_5521,N_5170,N_5030);
or U5522 (N_5522,N_5197,N_5167);
nor U5523 (N_5523,N_5181,N_5265);
and U5524 (N_5524,N_5498,N_5097);
nand U5525 (N_5525,N_5025,N_5180);
nor U5526 (N_5526,N_5451,N_5306);
or U5527 (N_5527,N_5153,N_5029);
nor U5528 (N_5528,N_5339,N_5345);
and U5529 (N_5529,N_5372,N_5272);
or U5530 (N_5530,N_5300,N_5019);
and U5531 (N_5531,N_5236,N_5386);
nor U5532 (N_5532,N_5118,N_5367);
nand U5533 (N_5533,N_5485,N_5083);
xnor U5534 (N_5534,N_5214,N_5488);
nor U5535 (N_5535,N_5082,N_5493);
nand U5536 (N_5536,N_5369,N_5036);
xnor U5537 (N_5537,N_5431,N_5258);
and U5538 (N_5538,N_5125,N_5392);
nor U5539 (N_5539,N_5033,N_5428);
xor U5540 (N_5540,N_5413,N_5240);
xor U5541 (N_5541,N_5175,N_5303);
or U5542 (N_5542,N_5247,N_5337);
and U5543 (N_5543,N_5069,N_5201);
nor U5544 (N_5544,N_5065,N_5059);
or U5545 (N_5545,N_5011,N_5366);
nor U5546 (N_5546,N_5228,N_5352);
and U5547 (N_5547,N_5299,N_5136);
or U5548 (N_5548,N_5489,N_5461);
nor U5549 (N_5549,N_5497,N_5188);
and U5550 (N_5550,N_5219,N_5128);
and U5551 (N_5551,N_5206,N_5443);
nand U5552 (N_5552,N_5129,N_5285);
and U5553 (N_5553,N_5255,N_5267);
and U5554 (N_5554,N_5293,N_5268);
xor U5555 (N_5555,N_5326,N_5191);
nor U5556 (N_5556,N_5449,N_5408);
nand U5557 (N_5557,N_5354,N_5172);
and U5558 (N_5558,N_5143,N_5329);
nor U5559 (N_5559,N_5338,N_5430);
and U5560 (N_5560,N_5198,N_5117);
nor U5561 (N_5561,N_5295,N_5283);
and U5562 (N_5562,N_5390,N_5043);
nor U5563 (N_5563,N_5297,N_5023);
nor U5564 (N_5564,N_5041,N_5151);
nand U5565 (N_5565,N_5371,N_5270);
nor U5566 (N_5566,N_5391,N_5370);
and U5567 (N_5567,N_5279,N_5452);
and U5568 (N_5568,N_5402,N_5146);
xor U5569 (N_5569,N_5472,N_5200);
or U5570 (N_5570,N_5157,N_5420);
xor U5571 (N_5571,N_5212,N_5321);
and U5572 (N_5572,N_5335,N_5446);
xor U5573 (N_5573,N_5464,N_5499);
and U5574 (N_5574,N_5055,N_5310);
nor U5575 (N_5575,N_5194,N_5102);
or U5576 (N_5576,N_5348,N_5089);
nor U5577 (N_5577,N_5323,N_5232);
xnor U5578 (N_5578,N_5308,N_5113);
nor U5579 (N_5579,N_5330,N_5252);
or U5580 (N_5580,N_5207,N_5465);
nor U5581 (N_5581,N_5211,N_5296);
and U5582 (N_5582,N_5166,N_5058);
nor U5583 (N_5583,N_5222,N_5463);
nor U5584 (N_5584,N_5165,N_5406);
xnor U5585 (N_5585,N_5317,N_5042);
xor U5586 (N_5586,N_5477,N_5060);
nor U5587 (N_5587,N_5253,N_5226);
nor U5588 (N_5588,N_5459,N_5439);
nand U5589 (N_5589,N_5470,N_5084);
nand U5590 (N_5590,N_5450,N_5480);
xnor U5591 (N_5591,N_5022,N_5399);
and U5592 (N_5592,N_5203,N_5251);
nor U5593 (N_5593,N_5003,N_5478);
xnor U5594 (N_5594,N_5286,N_5238);
nor U5595 (N_5595,N_5009,N_5087);
and U5596 (N_5596,N_5466,N_5394);
xnor U5597 (N_5597,N_5432,N_5365);
or U5598 (N_5598,N_5134,N_5234);
xor U5599 (N_5599,N_5205,N_5173);
and U5600 (N_5600,N_5216,N_5273);
and U5601 (N_5601,N_5351,N_5483);
nand U5602 (N_5602,N_5319,N_5347);
or U5603 (N_5603,N_5401,N_5441);
xor U5604 (N_5604,N_5196,N_5373);
nand U5605 (N_5605,N_5103,N_5486);
and U5606 (N_5606,N_5256,N_5142);
xor U5607 (N_5607,N_5095,N_5168);
and U5608 (N_5608,N_5220,N_5344);
xor U5609 (N_5609,N_5111,N_5434);
or U5610 (N_5610,N_5229,N_5456);
nor U5611 (N_5611,N_5260,N_5290);
or U5612 (N_5612,N_5107,N_5379);
or U5613 (N_5613,N_5389,N_5479);
nand U5614 (N_5614,N_5495,N_5148);
or U5615 (N_5615,N_5015,N_5051);
nor U5616 (N_5616,N_5274,N_5026);
nand U5617 (N_5617,N_5437,N_5161);
or U5618 (N_5618,N_5494,N_5315);
nor U5619 (N_5619,N_5482,N_5375);
nand U5620 (N_5620,N_5487,N_5387);
or U5621 (N_5621,N_5176,N_5045);
or U5622 (N_5622,N_5223,N_5418);
or U5623 (N_5623,N_5187,N_5353);
nor U5624 (N_5624,N_5108,N_5008);
or U5625 (N_5625,N_5358,N_5204);
and U5626 (N_5626,N_5340,N_5316);
or U5627 (N_5627,N_5039,N_5179);
or U5628 (N_5628,N_5235,N_5416);
or U5629 (N_5629,N_5250,N_5332);
nor U5630 (N_5630,N_5318,N_5481);
and U5631 (N_5631,N_5417,N_5447);
nor U5632 (N_5632,N_5455,N_5044);
nor U5633 (N_5633,N_5271,N_5020);
or U5634 (N_5634,N_5309,N_5262);
nand U5635 (N_5635,N_5414,N_5169);
nor U5636 (N_5636,N_5491,N_5032);
xnor U5637 (N_5637,N_5248,N_5233);
xnor U5638 (N_5638,N_5110,N_5382);
nor U5639 (N_5639,N_5287,N_5050);
nor U5640 (N_5640,N_5218,N_5397);
or U5641 (N_5641,N_5355,N_5171);
nor U5642 (N_5642,N_5453,N_5124);
or U5643 (N_5643,N_5024,N_5440);
and U5644 (N_5644,N_5017,N_5341);
xor U5645 (N_5645,N_5412,N_5158);
or U5646 (N_5646,N_5056,N_5411);
nor U5647 (N_5647,N_5139,N_5469);
xor U5648 (N_5648,N_5037,N_5263);
or U5649 (N_5649,N_5266,N_5031);
and U5650 (N_5650,N_5048,N_5121);
xnor U5651 (N_5651,N_5028,N_5049);
xnor U5652 (N_5652,N_5438,N_5156);
nand U5653 (N_5653,N_5403,N_5246);
nand U5654 (N_5654,N_5278,N_5289);
and U5655 (N_5655,N_5213,N_5141);
xnor U5656 (N_5656,N_5182,N_5064);
nand U5657 (N_5657,N_5407,N_5164);
nor U5658 (N_5658,N_5070,N_5178);
nand U5659 (N_5659,N_5126,N_5071);
xor U5660 (N_5660,N_5342,N_5068);
and U5661 (N_5661,N_5090,N_5086);
or U5662 (N_5662,N_5160,N_5364);
or U5663 (N_5663,N_5006,N_5301);
xnor U5664 (N_5664,N_5275,N_5004);
and U5665 (N_5665,N_5484,N_5378);
nand U5666 (N_5666,N_5473,N_5314);
nand U5667 (N_5667,N_5190,N_5144);
or U5668 (N_5668,N_5005,N_5093);
xnor U5669 (N_5669,N_5014,N_5245);
xnor U5670 (N_5670,N_5409,N_5426);
nor U5671 (N_5671,N_5067,N_5415);
nand U5672 (N_5672,N_5127,N_5302);
or U5673 (N_5673,N_5027,N_5288);
or U5674 (N_5674,N_5383,N_5435);
and U5675 (N_5675,N_5122,N_5346);
xor U5676 (N_5676,N_5468,N_5098);
nor U5677 (N_5677,N_5092,N_5425);
or U5678 (N_5678,N_5076,N_5312);
or U5679 (N_5679,N_5311,N_5096);
or U5680 (N_5680,N_5462,N_5012);
xnor U5681 (N_5681,N_5040,N_5334);
and U5682 (N_5682,N_5325,N_5433);
nor U5683 (N_5683,N_5239,N_5244);
nor U5684 (N_5684,N_5150,N_5013);
nand U5685 (N_5685,N_5101,N_5010);
xnor U5686 (N_5686,N_5476,N_5147);
xor U5687 (N_5687,N_5361,N_5080);
nor U5688 (N_5688,N_5132,N_5116);
nor U5689 (N_5689,N_5381,N_5460);
or U5690 (N_5690,N_5419,N_5094);
nor U5691 (N_5691,N_5259,N_5357);
nand U5692 (N_5692,N_5292,N_5077);
xnor U5693 (N_5693,N_5119,N_5054);
nor U5694 (N_5694,N_5047,N_5380);
nor U5695 (N_5695,N_5405,N_5057);
and U5696 (N_5696,N_5189,N_5079);
or U5697 (N_5697,N_5257,N_5474);
or U5698 (N_5698,N_5195,N_5304);
and U5699 (N_5699,N_5336,N_5496);
nor U5700 (N_5700,N_5423,N_5074);
nand U5701 (N_5701,N_5002,N_5034);
or U5702 (N_5702,N_5149,N_5225);
and U5703 (N_5703,N_5221,N_5400);
nor U5704 (N_5704,N_5398,N_5230);
and U5705 (N_5705,N_5277,N_5209);
nand U5706 (N_5706,N_5282,N_5436);
xor U5707 (N_5707,N_5099,N_5091);
and U5708 (N_5708,N_5261,N_5376);
nor U5709 (N_5709,N_5457,N_5193);
or U5710 (N_5710,N_5320,N_5385);
nand U5711 (N_5711,N_5152,N_5448);
xor U5712 (N_5712,N_5018,N_5359);
nor U5713 (N_5713,N_5163,N_5276);
xnor U5714 (N_5714,N_5281,N_5185);
xnor U5715 (N_5715,N_5215,N_5294);
nand U5716 (N_5716,N_5242,N_5135);
xor U5717 (N_5717,N_5374,N_5343);
nor U5718 (N_5718,N_5492,N_5035);
nand U5719 (N_5719,N_5384,N_5322);
nand U5720 (N_5720,N_5377,N_5410);
and U5721 (N_5721,N_5475,N_5349);
xnor U5722 (N_5722,N_5177,N_5227);
nand U5723 (N_5723,N_5490,N_5280);
and U5724 (N_5724,N_5155,N_5363);
xor U5725 (N_5725,N_5073,N_5454);
or U5726 (N_5726,N_5210,N_5291);
nand U5727 (N_5727,N_5123,N_5145);
nor U5728 (N_5728,N_5104,N_5085);
nor U5729 (N_5729,N_5388,N_5109);
and U5730 (N_5730,N_5159,N_5038);
nand U5731 (N_5731,N_5138,N_5427);
nand U5732 (N_5732,N_5131,N_5140);
and U5733 (N_5733,N_5184,N_5305);
and U5734 (N_5734,N_5269,N_5362);
nor U5735 (N_5735,N_5061,N_5137);
or U5736 (N_5736,N_5088,N_5162);
and U5737 (N_5737,N_5106,N_5016);
and U5738 (N_5738,N_5021,N_5192);
and U5739 (N_5739,N_5471,N_5072);
and U5740 (N_5740,N_5404,N_5217);
and U5741 (N_5741,N_5100,N_5444);
or U5742 (N_5742,N_5186,N_5241);
nand U5743 (N_5743,N_5183,N_5249);
nor U5744 (N_5744,N_5001,N_5053);
nand U5745 (N_5745,N_5424,N_5231);
nand U5746 (N_5746,N_5174,N_5208);
nor U5747 (N_5747,N_5120,N_5350);
or U5748 (N_5748,N_5254,N_5112);
xnor U5749 (N_5749,N_5442,N_5327);
nand U5750 (N_5750,N_5038,N_5313);
and U5751 (N_5751,N_5084,N_5305);
and U5752 (N_5752,N_5291,N_5234);
xor U5753 (N_5753,N_5174,N_5135);
nor U5754 (N_5754,N_5035,N_5422);
nand U5755 (N_5755,N_5337,N_5411);
and U5756 (N_5756,N_5307,N_5448);
xnor U5757 (N_5757,N_5246,N_5252);
nor U5758 (N_5758,N_5260,N_5173);
or U5759 (N_5759,N_5417,N_5354);
and U5760 (N_5760,N_5305,N_5197);
and U5761 (N_5761,N_5431,N_5463);
or U5762 (N_5762,N_5103,N_5470);
and U5763 (N_5763,N_5057,N_5145);
and U5764 (N_5764,N_5455,N_5388);
and U5765 (N_5765,N_5275,N_5092);
xnor U5766 (N_5766,N_5054,N_5222);
xor U5767 (N_5767,N_5258,N_5142);
nor U5768 (N_5768,N_5036,N_5410);
and U5769 (N_5769,N_5052,N_5303);
nand U5770 (N_5770,N_5211,N_5339);
nor U5771 (N_5771,N_5332,N_5312);
and U5772 (N_5772,N_5109,N_5403);
nor U5773 (N_5773,N_5185,N_5166);
xor U5774 (N_5774,N_5451,N_5014);
or U5775 (N_5775,N_5200,N_5278);
and U5776 (N_5776,N_5399,N_5370);
nor U5777 (N_5777,N_5271,N_5410);
nand U5778 (N_5778,N_5044,N_5103);
or U5779 (N_5779,N_5146,N_5410);
and U5780 (N_5780,N_5395,N_5264);
or U5781 (N_5781,N_5060,N_5062);
or U5782 (N_5782,N_5350,N_5498);
nand U5783 (N_5783,N_5190,N_5121);
xnor U5784 (N_5784,N_5379,N_5348);
xor U5785 (N_5785,N_5490,N_5297);
nand U5786 (N_5786,N_5047,N_5167);
or U5787 (N_5787,N_5371,N_5152);
xnor U5788 (N_5788,N_5423,N_5111);
xor U5789 (N_5789,N_5342,N_5345);
and U5790 (N_5790,N_5204,N_5393);
xnor U5791 (N_5791,N_5159,N_5041);
xor U5792 (N_5792,N_5077,N_5432);
nor U5793 (N_5793,N_5240,N_5095);
nand U5794 (N_5794,N_5167,N_5400);
nand U5795 (N_5795,N_5197,N_5162);
or U5796 (N_5796,N_5498,N_5151);
or U5797 (N_5797,N_5351,N_5291);
nand U5798 (N_5798,N_5465,N_5034);
nand U5799 (N_5799,N_5342,N_5406);
and U5800 (N_5800,N_5422,N_5265);
and U5801 (N_5801,N_5396,N_5014);
nor U5802 (N_5802,N_5049,N_5474);
or U5803 (N_5803,N_5116,N_5490);
nor U5804 (N_5804,N_5375,N_5238);
nand U5805 (N_5805,N_5409,N_5334);
or U5806 (N_5806,N_5128,N_5020);
and U5807 (N_5807,N_5223,N_5173);
and U5808 (N_5808,N_5176,N_5098);
xnor U5809 (N_5809,N_5024,N_5035);
or U5810 (N_5810,N_5277,N_5307);
or U5811 (N_5811,N_5296,N_5439);
nor U5812 (N_5812,N_5051,N_5085);
or U5813 (N_5813,N_5462,N_5273);
and U5814 (N_5814,N_5402,N_5473);
or U5815 (N_5815,N_5007,N_5433);
xnor U5816 (N_5816,N_5095,N_5071);
xor U5817 (N_5817,N_5078,N_5198);
nor U5818 (N_5818,N_5042,N_5264);
or U5819 (N_5819,N_5199,N_5467);
or U5820 (N_5820,N_5037,N_5372);
or U5821 (N_5821,N_5368,N_5492);
nand U5822 (N_5822,N_5181,N_5325);
and U5823 (N_5823,N_5477,N_5242);
nor U5824 (N_5824,N_5080,N_5491);
nor U5825 (N_5825,N_5154,N_5343);
or U5826 (N_5826,N_5013,N_5042);
nor U5827 (N_5827,N_5362,N_5439);
xor U5828 (N_5828,N_5248,N_5114);
and U5829 (N_5829,N_5240,N_5146);
nand U5830 (N_5830,N_5236,N_5378);
xor U5831 (N_5831,N_5444,N_5291);
nand U5832 (N_5832,N_5305,N_5494);
nand U5833 (N_5833,N_5480,N_5320);
nand U5834 (N_5834,N_5200,N_5209);
xnor U5835 (N_5835,N_5256,N_5010);
xor U5836 (N_5836,N_5333,N_5069);
and U5837 (N_5837,N_5274,N_5477);
nand U5838 (N_5838,N_5334,N_5248);
nor U5839 (N_5839,N_5110,N_5146);
xnor U5840 (N_5840,N_5314,N_5219);
and U5841 (N_5841,N_5001,N_5334);
and U5842 (N_5842,N_5011,N_5235);
or U5843 (N_5843,N_5450,N_5393);
or U5844 (N_5844,N_5493,N_5372);
nor U5845 (N_5845,N_5374,N_5277);
nand U5846 (N_5846,N_5432,N_5478);
xnor U5847 (N_5847,N_5260,N_5131);
and U5848 (N_5848,N_5181,N_5187);
and U5849 (N_5849,N_5147,N_5282);
and U5850 (N_5850,N_5355,N_5375);
nand U5851 (N_5851,N_5070,N_5044);
and U5852 (N_5852,N_5341,N_5091);
nor U5853 (N_5853,N_5430,N_5094);
and U5854 (N_5854,N_5153,N_5384);
nor U5855 (N_5855,N_5115,N_5341);
or U5856 (N_5856,N_5380,N_5130);
nor U5857 (N_5857,N_5235,N_5499);
nor U5858 (N_5858,N_5029,N_5421);
or U5859 (N_5859,N_5280,N_5028);
or U5860 (N_5860,N_5079,N_5434);
or U5861 (N_5861,N_5057,N_5288);
nand U5862 (N_5862,N_5002,N_5335);
or U5863 (N_5863,N_5021,N_5245);
and U5864 (N_5864,N_5282,N_5221);
nand U5865 (N_5865,N_5418,N_5380);
or U5866 (N_5866,N_5402,N_5321);
or U5867 (N_5867,N_5206,N_5087);
and U5868 (N_5868,N_5253,N_5147);
nand U5869 (N_5869,N_5412,N_5061);
nand U5870 (N_5870,N_5332,N_5163);
nor U5871 (N_5871,N_5275,N_5273);
nor U5872 (N_5872,N_5459,N_5213);
xnor U5873 (N_5873,N_5054,N_5479);
nand U5874 (N_5874,N_5175,N_5183);
nor U5875 (N_5875,N_5150,N_5125);
xnor U5876 (N_5876,N_5153,N_5074);
nand U5877 (N_5877,N_5408,N_5027);
nand U5878 (N_5878,N_5177,N_5357);
and U5879 (N_5879,N_5381,N_5171);
xor U5880 (N_5880,N_5463,N_5477);
nor U5881 (N_5881,N_5473,N_5394);
or U5882 (N_5882,N_5429,N_5161);
nor U5883 (N_5883,N_5397,N_5149);
and U5884 (N_5884,N_5261,N_5128);
nand U5885 (N_5885,N_5207,N_5013);
nor U5886 (N_5886,N_5092,N_5189);
xor U5887 (N_5887,N_5139,N_5205);
or U5888 (N_5888,N_5046,N_5425);
nor U5889 (N_5889,N_5073,N_5175);
and U5890 (N_5890,N_5166,N_5443);
and U5891 (N_5891,N_5297,N_5217);
or U5892 (N_5892,N_5425,N_5274);
nand U5893 (N_5893,N_5277,N_5345);
xor U5894 (N_5894,N_5370,N_5129);
or U5895 (N_5895,N_5435,N_5434);
or U5896 (N_5896,N_5483,N_5038);
nand U5897 (N_5897,N_5276,N_5231);
nor U5898 (N_5898,N_5461,N_5246);
nor U5899 (N_5899,N_5230,N_5049);
and U5900 (N_5900,N_5228,N_5464);
or U5901 (N_5901,N_5205,N_5369);
xor U5902 (N_5902,N_5446,N_5490);
xnor U5903 (N_5903,N_5431,N_5437);
or U5904 (N_5904,N_5404,N_5020);
nor U5905 (N_5905,N_5129,N_5393);
nor U5906 (N_5906,N_5200,N_5364);
nor U5907 (N_5907,N_5340,N_5004);
xor U5908 (N_5908,N_5479,N_5268);
or U5909 (N_5909,N_5083,N_5410);
or U5910 (N_5910,N_5128,N_5114);
nand U5911 (N_5911,N_5255,N_5170);
or U5912 (N_5912,N_5293,N_5174);
nor U5913 (N_5913,N_5372,N_5313);
or U5914 (N_5914,N_5238,N_5121);
and U5915 (N_5915,N_5471,N_5192);
or U5916 (N_5916,N_5154,N_5132);
and U5917 (N_5917,N_5284,N_5305);
nand U5918 (N_5918,N_5056,N_5042);
xnor U5919 (N_5919,N_5333,N_5491);
xor U5920 (N_5920,N_5292,N_5097);
nand U5921 (N_5921,N_5083,N_5274);
nand U5922 (N_5922,N_5401,N_5008);
and U5923 (N_5923,N_5033,N_5228);
xnor U5924 (N_5924,N_5428,N_5191);
or U5925 (N_5925,N_5164,N_5061);
nor U5926 (N_5926,N_5169,N_5446);
nor U5927 (N_5927,N_5240,N_5465);
or U5928 (N_5928,N_5074,N_5293);
xor U5929 (N_5929,N_5342,N_5266);
and U5930 (N_5930,N_5445,N_5457);
and U5931 (N_5931,N_5420,N_5343);
and U5932 (N_5932,N_5400,N_5117);
nand U5933 (N_5933,N_5388,N_5376);
xnor U5934 (N_5934,N_5474,N_5112);
nor U5935 (N_5935,N_5371,N_5037);
xor U5936 (N_5936,N_5231,N_5445);
and U5937 (N_5937,N_5373,N_5125);
or U5938 (N_5938,N_5394,N_5299);
nand U5939 (N_5939,N_5312,N_5217);
nor U5940 (N_5940,N_5149,N_5444);
xor U5941 (N_5941,N_5268,N_5353);
nor U5942 (N_5942,N_5066,N_5394);
xnor U5943 (N_5943,N_5468,N_5135);
nor U5944 (N_5944,N_5287,N_5171);
nor U5945 (N_5945,N_5258,N_5226);
and U5946 (N_5946,N_5204,N_5377);
or U5947 (N_5947,N_5435,N_5166);
xor U5948 (N_5948,N_5442,N_5392);
xnor U5949 (N_5949,N_5362,N_5245);
xnor U5950 (N_5950,N_5377,N_5183);
xnor U5951 (N_5951,N_5113,N_5083);
nand U5952 (N_5952,N_5445,N_5198);
xnor U5953 (N_5953,N_5188,N_5098);
and U5954 (N_5954,N_5011,N_5313);
and U5955 (N_5955,N_5468,N_5474);
nor U5956 (N_5956,N_5451,N_5066);
and U5957 (N_5957,N_5036,N_5122);
or U5958 (N_5958,N_5265,N_5362);
or U5959 (N_5959,N_5113,N_5419);
xor U5960 (N_5960,N_5277,N_5290);
and U5961 (N_5961,N_5317,N_5099);
nand U5962 (N_5962,N_5157,N_5140);
or U5963 (N_5963,N_5165,N_5361);
nor U5964 (N_5964,N_5033,N_5278);
nor U5965 (N_5965,N_5149,N_5416);
xor U5966 (N_5966,N_5099,N_5415);
nor U5967 (N_5967,N_5340,N_5027);
xor U5968 (N_5968,N_5087,N_5470);
xor U5969 (N_5969,N_5129,N_5153);
nand U5970 (N_5970,N_5347,N_5024);
nand U5971 (N_5971,N_5077,N_5222);
nand U5972 (N_5972,N_5170,N_5105);
or U5973 (N_5973,N_5474,N_5311);
nand U5974 (N_5974,N_5211,N_5458);
nor U5975 (N_5975,N_5396,N_5128);
xor U5976 (N_5976,N_5079,N_5486);
and U5977 (N_5977,N_5475,N_5104);
or U5978 (N_5978,N_5055,N_5043);
xor U5979 (N_5979,N_5289,N_5343);
nand U5980 (N_5980,N_5184,N_5251);
xnor U5981 (N_5981,N_5197,N_5378);
nor U5982 (N_5982,N_5381,N_5396);
nand U5983 (N_5983,N_5174,N_5070);
or U5984 (N_5984,N_5363,N_5067);
or U5985 (N_5985,N_5093,N_5088);
or U5986 (N_5986,N_5245,N_5119);
xor U5987 (N_5987,N_5051,N_5183);
or U5988 (N_5988,N_5405,N_5306);
or U5989 (N_5989,N_5461,N_5317);
xor U5990 (N_5990,N_5036,N_5434);
or U5991 (N_5991,N_5151,N_5209);
and U5992 (N_5992,N_5004,N_5226);
or U5993 (N_5993,N_5258,N_5037);
xor U5994 (N_5994,N_5312,N_5003);
xnor U5995 (N_5995,N_5295,N_5278);
or U5996 (N_5996,N_5364,N_5084);
nor U5997 (N_5997,N_5297,N_5255);
or U5998 (N_5998,N_5081,N_5283);
nand U5999 (N_5999,N_5259,N_5063);
nand U6000 (N_6000,N_5569,N_5692);
nand U6001 (N_6001,N_5863,N_5638);
or U6002 (N_6002,N_5646,N_5576);
nor U6003 (N_6003,N_5525,N_5659);
and U6004 (N_6004,N_5568,N_5688);
or U6005 (N_6005,N_5864,N_5862);
nor U6006 (N_6006,N_5691,N_5809);
or U6007 (N_6007,N_5869,N_5747);
nand U6008 (N_6008,N_5765,N_5612);
nor U6009 (N_6009,N_5939,N_5535);
xnor U6010 (N_6010,N_5908,N_5741);
and U6011 (N_6011,N_5843,N_5935);
xor U6012 (N_6012,N_5918,N_5983);
xnor U6013 (N_6013,N_5859,N_5871);
xnor U6014 (N_6014,N_5721,N_5855);
xor U6015 (N_6015,N_5740,N_5616);
or U6016 (N_6016,N_5718,N_5946);
and U6017 (N_6017,N_5517,N_5522);
nor U6018 (N_6018,N_5686,N_5753);
or U6019 (N_6019,N_5713,N_5913);
xor U6020 (N_6020,N_5929,N_5565);
nor U6021 (N_6021,N_5647,N_5622);
or U6022 (N_6022,N_5743,N_5878);
nand U6023 (N_6023,N_5549,N_5722);
nand U6024 (N_6024,N_5528,N_5603);
nand U6025 (N_6025,N_5799,N_5866);
and U6026 (N_6026,N_5538,N_5769);
xor U6027 (N_6027,N_5557,N_5815);
and U6028 (N_6028,N_5635,N_5544);
or U6029 (N_6029,N_5999,N_5950);
or U6030 (N_6030,N_5602,N_5787);
nor U6031 (N_6031,N_5583,N_5841);
nor U6032 (N_6032,N_5888,N_5853);
or U6033 (N_6033,N_5847,N_5628);
xnor U6034 (N_6034,N_5987,N_5667);
nor U6035 (N_6035,N_5512,N_5954);
or U6036 (N_6036,N_5814,N_5566);
or U6037 (N_6037,N_5624,N_5955);
or U6038 (N_6038,N_5690,N_5744);
nor U6039 (N_6039,N_5840,N_5861);
and U6040 (N_6040,N_5529,N_5959);
and U6041 (N_6041,N_5904,N_5676);
nor U6042 (N_6042,N_5597,N_5778);
xor U6043 (N_6043,N_5651,N_5532);
xor U6044 (N_6044,N_5926,N_5848);
and U6045 (N_6045,N_5825,N_5501);
or U6046 (N_6046,N_5687,N_5613);
and U6047 (N_6047,N_5996,N_5754);
and U6048 (N_6048,N_5828,N_5974);
xor U6049 (N_6049,N_5988,N_5604);
or U6050 (N_6050,N_5877,N_5795);
and U6051 (N_6051,N_5821,N_5960);
nand U6052 (N_6052,N_5555,N_5502);
nor U6053 (N_6053,N_5984,N_5961);
and U6054 (N_6054,N_5867,N_5817);
xnor U6055 (N_6055,N_5886,N_5981);
or U6056 (N_6056,N_5641,N_5749);
and U6057 (N_6057,N_5806,N_5515);
nand U6058 (N_6058,N_5683,N_5581);
nand U6059 (N_6059,N_5763,N_5800);
nor U6060 (N_6060,N_5533,N_5601);
xor U6061 (N_6061,N_5591,N_5665);
and U6062 (N_6062,N_5547,N_5680);
nor U6063 (N_6063,N_5865,N_5678);
xor U6064 (N_6064,N_5643,N_5720);
or U6065 (N_6065,N_5776,N_5978);
or U6066 (N_6066,N_5664,N_5571);
or U6067 (N_6067,N_5923,N_5589);
or U6068 (N_6068,N_5975,N_5600);
and U6069 (N_6069,N_5541,N_5654);
xor U6070 (N_6070,N_5816,N_5531);
or U6071 (N_6071,N_5693,N_5971);
nor U6072 (N_6072,N_5938,N_5810);
and U6073 (N_6073,N_5898,N_5627);
nor U6074 (N_6074,N_5893,N_5605);
xor U6075 (N_6075,N_5916,N_5737);
nand U6076 (N_6076,N_5782,N_5656);
nor U6077 (N_6077,N_5586,N_5907);
or U6078 (N_6078,N_5868,N_5801);
or U6079 (N_6079,N_5719,N_5796);
nor U6080 (N_6080,N_5663,N_5573);
or U6081 (N_6081,N_5970,N_5653);
nand U6082 (N_6082,N_5882,N_5550);
or U6083 (N_6083,N_5579,N_5774);
and U6084 (N_6084,N_5542,N_5798);
and U6085 (N_6085,N_5995,N_5924);
or U6086 (N_6086,N_5900,N_5513);
nand U6087 (N_6087,N_5792,N_5596);
nand U6088 (N_6088,N_5773,N_5615);
or U6089 (N_6089,N_5844,N_5606);
and U6090 (N_6090,N_5756,N_5958);
or U6091 (N_6091,N_5732,N_5964);
nor U6092 (N_6092,N_5738,N_5558);
or U6093 (N_6093,N_5682,N_5887);
and U6094 (N_6094,N_5771,N_5534);
nand U6095 (N_6095,N_5514,N_5652);
and U6096 (N_6096,N_5742,N_5967);
and U6097 (N_6097,N_5715,N_5839);
xor U6098 (N_6098,N_5963,N_5642);
nand U6099 (N_6099,N_5824,N_5711);
and U6100 (N_6100,N_5927,N_5716);
nand U6101 (N_6101,N_5835,N_5519);
and U6102 (N_6102,N_5858,N_5873);
and U6103 (N_6103,N_5625,N_5649);
and U6104 (N_6104,N_5694,N_5758);
or U6105 (N_6105,N_5503,N_5508);
or U6106 (N_6106,N_5553,N_5751);
nand U6107 (N_6107,N_5791,N_5752);
nor U6108 (N_6108,N_5574,N_5832);
or U6109 (N_6109,N_5662,N_5933);
nand U6110 (N_6110,N_5731,N_5854);
xnor U6111 (N_6111,N_5903,N_5819);
and U6112 (N_6112,N_5607,N_5644);
nor U6113 (N_6113,N_5631,N_5993);
xor U6114 (N_6114,N_5895,N_5559);
or U6115 (N_6115,N_5634,N_5770);
and U6116 (N_6116,N_5872,N_5726);
and U6117 (N_6117,N_5714,N_5925);
nor U6118 (N_6118,N_5768,N_5932);
or U6119 (N_6119,N_5831,N_5965);
nand U6120 (N_6120,N_5704,N_5997);
nor U6121 (N_6121,N_5811,N_5702);
xnor U6122 (N_6122,N_5881,N_5640);
nand U6123 (N_6123,N_5560,N_5775);
nand U6124 (N_6124,N_5703,N_5906);
and U6125 (N_6125,N_5896,N_5725);
or U6126 (N_6126,N_5911,N_5618);
or U6127 (N_6127,N_5973,N_5750);
nand U6128 (N_6128,N_5707,N_5812);
nand U6129 (N_6129,N_5941,N_5966);
xnor U6130 (N_6130,N_5500,N_5745);
xnor U6131 (N_6131,N_5705,N_5919);
xor U6132 (N_6132,N_5505,N_5636);
nand U6133 (N_6133,N_5685,N_5951);
nand U6134 (N_6134,N_5793,N_5789);
nand U6135 (N_6135,N_5681,N_5985);
or U6136 (N_6136,N_5518,N_5823);
xor U6137 (N_6137,N_5708,N_5728);
and U6138 (N_6138,N_5998,N_5945);
nand U6139 (N_6139,N_5609,N_5546);
nand U6140 (N_6140,N_5953,N_5802);
and U6141 (N_6141,N_5524,N_5930);
or U6142 (N_6142,N_5599,N_5709);
nand U6143 (N_6143,N_5510,N_5590);
or U6144 (N_6144,N_5739,N_5784);
and U6145 (N_6145,N_5736,N_5915);
nor U6146 (N_6146,N_5991,N_5899);
nor U6147 (N_6147,N_5766,N_5539);
and U6148 (N_6148,N_5598,N_5761);
nor U6149 (N_6149,N_5675,N_5632);
nor U6150 (N_6150,N_5710,N_5757);
nor U6151 (N_6151,N_5548,N_5699);
or U6152 (N_6152,N_5584,N_5949);
nand U6153 (N_6153,N_5897,N_5875);
nor U6154 (N_6154,N_5734,N_5698);
xor U6155 (N_6155,N_5788,N_5626);
and U6156 (N_6156,N_5509,N_5593);
nor U6157 (N_6157,N_5696,N_5931);
and U6158 (N_6158,N_5504,N_5850);
and U6159 (N_6159,N_5672,N_5836);
nand U6160 (N_6160,N_5712,N_5660);
xor U6161 (N_6161,N_5820,N_5697);
and U6162 (N_6162,N_5575,N_5578);
and U6163 (N_6163,N_5564,N_5942);
or U6164 (N_6164,N_5822,N_5717);
nor U6165 (N_6165,N_5562,N_5608);
nor U6166 (N_6166,N_5706,N_5890);
and U6167 (N_6167,N_5689,N_5972);
nor U6168 (N_6168,N_5779,N_5992);
or U6169 (N_6169,N_5909,N_5670);
nand U6170 (N_6170,N_5679,N_5764);
nand U6171 (N_6171,N_5520,N_5804);
or U6172 (N_6172,N_5570,N_5914);
xor U6173 (N_6173,N_5797,N_5934);
nor U6174 (N_6174,N_5552,N_5860);
nand U6175 (N_6175,N_5645,N_5902);
nand U6176 (N_6176,N_5561,N_5577);
xor U6177 (N_6177,N_5813,N_5956);
xor U6178 (N_6178,N_5912,N_5982);
nand U6179 (N_6179,N_5610,N_5786);
nand U6180 (N_6180,N_5759,N_5648);
and U6181 (N_6181,N_5735,N_5968);
and U6182 (N_6182,N_5623,N_5582);
nand U6183 (N_6183,N_5587,N_5733);
and U6184 (N_6184,N_5668,N_5594);
or U6185 (N_6185,N_5620,N_5891);
nor U6186 (N_6186,N_5760,N_5976);
and U6187 (N_6187,N_5677,N_5633);
nand U6188 (N_6188,N_5723,N_5655);
and U6189 (N_6189,N_5940,N_5980);
nand U6190 (N_6190,N_5540,N_5666);
xor U6191 (N_6191,N_5943,N_5536);
and U6192 (N_6192,N_5794,N_5521);
xor U6193 (N_6193,N_5511,N_5572);
and U6194 (N_6194,N_5669,N_5880);
nand U6195 (N_6195,N_5962,N_5554);
nor U6196 (N_6196,N_5994,N_5684);
nor U6197 (N_6197,N_5830,N_5834);
nor U6198 (N_6198,N_5805,N_5990);
nand U6199 (N_6199,N_5772,N_5857);
xnor U6200 (N_6200,N_5630,N_5506);
and U6201 (N_6201,N_5889,N_5567);
or U6202 (N_6202,N_5874,N_5545);
nand U6203 (N_6203,N_5730,N_5701);
or U6204 (N_6204,N_5852,N_5658);
nand U6205 (N_6205,N_5846,N_5674);
nand U6206 (N_6206,N_5790,N_5762);
xor U6207 (N_6207,N_5910,N_5838);
nand U6208 (N_6208,N_5781,N_5833);
xor U6209 (N_6209,N_5944,N_5920);
xnor U6210 (N_6210,N_5894,N_5516);
or U6211 (N_6211,N_5695,N_5808);
xor U6212 (N_6212,N_5783,N_5884);
nand U6213 (N_6213,N_5885,N_5977);
nor U6214 (N_6214,N_5948,N_5621);
and U6215 (N_6215,N_5849,N_5947);
xor U6216 (N_6216,N_5588,N_5986);
xor U6217 (N_6217,N_5729,N_5507);
and U6218 (N_6218,N_5989,N_5551);
or U6219 (N_6219,N_5556,N_5657);
nor U6220 (N_6220,N_5936,N_5727);
and U6221 (N_6221,N_5957,N_5905);
and U6222 (N_6222,N_5879,N_5922);
nand U6223 (N_6223,N_5870,N_5724);
or U6224 (N_6224,N_5748,N_5917);
nor U6225 (N_6225,N_5611,N_5818);
nand U6226 (N_6226,N_5614,N_5671);
and U6227 (N_6227,N_5807,N_5921);
or U6228 (N_6228,N_5937,N_5523);
and U6229 (N_6229,N_5979,N_5803);
nor U6230 (N_6230,N_5526,N_5543);
xnor U6231 (N_6231,N_5537,N_5700);
xnor U6232 (N_6232,N_5785,N_5767);
nand U6233 (N_6233,N_5755,N_5876);
xnor U6234 (N_6234,N_5619,N_5585);
xor U6235 (N_6235,N_5592,N_5637);
xnor U6236 (N_6236,N_5856,N_5650);
and U6237 (N_6237,N_5826,N_5780);
xor U6238 (N_6238,N_5527,N_5842);
nand U6239 (N_6239,N_5901,N_5928);
or U6240 (N_6240,N_5580,N_5639);
xnor U6241 (N_6241,N_5629,N_5952);
nand U6242 (N_6242,N_5563,N_5892);
nor U6243 (N_6243,N_5673,N_5617);
or U6244 (N_6244,N_5530,N_5969);
xnor U6245 (N_6245,N_5827,N_5837);
and U6246 (N_6246,N_5746,N_5595);
or U6247 (N_6247,N_5883,N_5851);
and U6248 (N_6248,N_5661,N_5845);
and U6249 (N_6249,N_5829,N_5777);
nor U6250 (N_6250,N_5543,N_5896);
or U6251 (N_6251,N_5837,N_5746);
nand U6252 (N_6252,N_5911,N_5889);
or U6253 (N_6253,N_5934,N_5662);
xor U6254 (N_6254,N_5633,N_5685);
and U6255 (N_6255,N_5742,N_5582);
xnor U6256 (N_6256,N_5835,N_5917);
and U6257 (N_6257,N_5614,N_5962);
xnor U6258 (N_6258,N_5559,N_5983);
nand U6259 (N_6259,N_5702,N_5911);
or U6260 (N_6260,N_5719,N_5683);
and U6261 (N_6261,N_5607,N_5979);
and U6262 (N_6262,N_5851,N_5669);
xnor U6263 (N_6263,N_5737,N_5935);
and U6264 (N_6264,N_5884,N_5841);
and U6265 (N_6265,N_5836,N_5837);
or U6266 (N_6266,N_5752,N_5629);
xor U6267 (N_6267,N_5990,N_5710);
and U6268 (N_6268,N_5723,N_5553);
or U6269 (N_6269,N_5998,N_5523);
or U6270 (N_6270,N_5982,N_5704);
or U6271 (N_6271,N_5593,N_5763);
and U6272 (N_6272,N_5934,N_5801);
and U6273 (N_6273,N_5882,N_5767);
xnor U6274 (N_6274,N_5793,N_5812);
xnor U6275 (N_6275,N_5983,N_5544);
nor U6276 (N_6276,N_5858,N_5997);
nor U6277 (N_6277,N_5734,N_5948);
or U6278 (N_6278,N_5981,N_5656);
xnor U6279 (N_6279,N_5592,N_5717);
nand U6280 (N_6280,N_5547,N_5589);
or U6281 (N_6281,N_5912,N_5538);
and U6282 (N_6282,N_5798,N_5909);
or U6283 (N_6283,N_5870,N_5897);
nand U6284 (N_6284,N_5922,N_5522);
nand U6285 (N_6285,N_5533,N_5989);
or U6286 (N_6286,N_5603,N_5936);
xor U6287 (N_6287,N_5653,N_5731);
or U6288 (N_6288,N_5928,N_5770);
and U6289 (N_6289,N_5949,N_5536);
or U6290 (N_6290,N_5660,N_5530);
nand U6291 (N_6291,N_5689,N_5592);
nor U6292 (N_6292,N_5550,N_5781);
nor U6293 (N_6293,N_5848,N_5633);
xnor U6294 (N_6294,N_5885,N_5857);
and U6295 (N_6295,N_5629,N_5700);
xnor U6296 (N_6296,N_5550,N_5828);
or U6297 (N_6297,N_5850,N_5680);
nand U6298 (N_6298,N_5505,N_5940);
nand U6299 (N_6299,N_5626,N_5852);
nand U6300 (N_6300,N_5869,N_5640);
and U6301 (N_6301,N_5975,N_5680);
nand U6302 (N_6302,N_5614,N_5523);
and U6303 (N_6303,N_5971,N_5950);
and U6304 (N_6304,N_5651,N_5690);
nor U6305 (N_6305,N_5902,N_5826);
xor U6306 (N_6306,N_5805,N_5578);
or U6307 (N_6307,N_5812,N_5671);
xor U6308 (N_6308,N_5663,N_5562);
nor U6309 (N_6309,N_5655,N_5922);
xnor U6310 (N_6310,N_5919,N_5848);
or U6311 (N_6311,N_5575,N_5723);
nand U6312 (N_6312,N_5937,N_5832);
or U6313 (N_6313,N_5700,N_5916);
xnor U6314 (N_6314,N_5539,N_5950);
or U6315 (N_6315,N_5817,N_5837);
or U6316 (N_6316,N_5821,N_5988);
nor U6317 (N_6317,N_5918,N_5554);
nor U6318 (N_6318,N_5738,N_5759);
nand U6319 (N_6319,N_5562,N_5665);
or U6320 (N_6320,N_5873,N_5928);
xor U6321 (N_6321,N_5826,N_5810);
and U6322 (N_6322,N_5516,N_5773);
nor U6323 (N_6323,N_5509,N_5977);
nor U6324 (N_6324,N_5839,N_5819);
nor U6325 (N_6325,N_5998,N_5774);
nor U6326 (N_6326,N_5990,N_5585);
nor U6327 (N_6327,N_5911,N_5560);
nor U6328 (N_6328,N_5936,N_5620);
xnor U6329 (N_6329,N_5729,N_5542);
nand U6330 (N_6330,N_5656,N_5523);
or U6331 (N_6331,N_5698,N_5761);
xnor U6332 (N_6332,N_5525,N_5724);
xnor U6333 (N_6333,N_5652,N_5913);
and U6334 (N_6334,N_5779,N_5799);
xnor U6335 (N_6335,N_5545,N_5901);
nand U6336 (N_6336,N_5661,N_5689);
and U6337 (N_6337,N_5653,N_5785);
or U6338 (N_6338,N_5701,N_5667);
nand U6339 (N_6339,N_5593,N_5691);
xnor U6340 (N_6340,N_5702,N_5830);
xnor U6341 (N_6341,N_5513,N_5555);
xnor U6342 (N_6342,N_5947,N_5627);
xnor U6343 (N_6343,N_5949,N_5843);
nand U6344 (N_6344,N_5856,N_5799);
nand U6345 (N_6345,N_5849,N_5807);
or U6346 (N_6346,N_5928,N_5869);
xnor U6347 (N_6347,N_5583,N_5858);
and U6348 (N_6348,N_5827,N_5613);
and U6349 (N_6349,N_5703,N_5688);
nor U6350 (N_6350,N_5651,N_5806);
nand U6351 (N_6351,N_5587,N_5671);
or U6352 (N_6352,N_5548,N_5607);
xnor U6353 (N_6353,N_5696,N_5528);
xor U6354 (N_6354,N_5815,N_5790);
nand U6355 (N_6355,N_5639,N_5759);
nor U6356 (N_6356,N_5916,N_5993);
nand U6357 (N_6357,N_5852,N_5926);
or U6358 (N_6358,N_5847,N_5920);
and U6359 (N_6359,N_5572,N_5910);
or U6360 (N_6360,N_5658,N_5941);
nor U6361 (N_6361,N_5720,N_5611);
nand U6362 (N_6362,N_5907,N_5605);
nand U6363 (N_6363,N_5865,N_5805);
nor U6364 (N_6364,N_5621,N_5610);
xnor U6365 (N_6365,N_5563,N_5594);
xor U6366 (N_6366,N_5815,N_5867);
nand U6367 (N_6367,N_5741,N_5858);
nand U6368 (N_6368,N_5994,N_5597);
or U6369 (N_6369,N_5797,N_5837);
nor U6370 (N_6370,N_5864,N_5613);
or U6371 (N_6371,N_5732,N_5887);
and U6372 (N_6372,N_5600,N_5963);
nor U6373 (N_6373,N_5864,N_5536);
nand U6374 (N_6374,N_5571,N_5799);
xor U6375 (N_6375,N_5570,N_5685);
nand U6376 (N_6376,N_5799,N_5803);
xor U6377 (N_6377,N_5656,N_5963);
xnor U6378 (N_6378,N_5976,N_5888);
nor U6379 (N_6379,N_5541,N_5656);
xor U6380 (N_6380,N_5891,N_5875);
nand U6381 (N_6381,N_5704,N_5556);
nor U6382 (N_6382,N_5577,N_5951);
and U6383 (N_6383,N_5901,N_5875);
xor U6384 (N_6384,N_5779,N_5511);
xor U6385 (N_6385,N_5580,N_5519);
nand U6386 (N_6386,N_5814,N_5750);
or U6387 (N_6387,N_5817,N_5514);
xor U6388 (N_6388,N_5760,N_5779);
xnor U6389 (N_6389,N_5665,N_5655);
nor U6390 (N_6390,N_5705,N_5791);
or U6391 (N_6391,N_5558,N_5683);
nor U6392 (N_6392,N_5666,N_5839);
and U6393 (N_6393,N_5856,N_5790);
and U6394 (N_6394,N_5713,N_5824);
xor U6395 (N_6395,N_5811,N_5738);
nand U6396 (N_6396,N_5886,N_5757);
xnor U6397 (N_6397,N_5617,N_5514);
or U6398 (N_6398,N_5894,N_5662);
nor U6399 (N_6399,N_5535,N_5836);
and U6400 (N_6400,N_5709,N_5632);
and U6401 (N_6401,N_5926,N_5711);
and U6402 (N_6402,N_5503,N_5964);
nor U6403 (N_6403,N_5632,N_5714);
nor U6404 (N_6404,N_5545,N_5529);
nor U6405 (N_6405,N_5792,N_5721);
or U6406 (N_6406,N_5633,N_5793);
and U6407 (N_6407,N_5995,N_5623);
nand U6408 (N_6408,N_5775,N_5861);
nand U6409 (N_6409,N_5718,N_5573);
xor U6410 (N_6410,N_5513,N_5752);
xor U6411 (N_6411,N_5931,N_5906);
nand U6412 (N_6412,N_5962,N_5930);
xnor U6413 (N_6413,N_5896,N_5666);
or U6414 (N_6414,N_5781,N_5656);
xor U6415 (N_6415,N_5764,N_5752);
nand U6416 (N_6416,N_5763,N_5891);
or U6417 (N_6417,N_5696,N_5864);
or U6418 (N_6418,N_5844,N_5997);
nor U6419 (N_6419,N_5724,N_5521);
or U6420 (N_6420,N_5891,N_5633);
xor U6421 (N_6421,N_5734,N_5576);
xnor U6422 (N_6422,N_5865,N_5997);
nor U6423 (N_6423,N_5671,N_5674);
and U6424 (N_6424,N_5821,N_5803);
nor U6425 (N_6425,N_5728,N_5961);
nand U6426 (N_6426,N_5755,N_5682);
and U6427 (N_6427,N_5655,N_5516);
nand U6428 (N_6428,N_5873,N_5779);
or U6429 (N_6429,N_5833,N_5802);
nor U6430 (N_6430,N_5830,N_5959);
nand U6431 (N_6431,N_5741,N_5712);
nand U6432 (N_6432,N_5848,N_5539);
nand U6433 (N_6433,N_5805,N_5822);
nand U6434 (N_6434,N_5948,N_5884);
and U6435 (N_6435,N_5655,N_5830);
or U6436 (N_6436,N_5510,N_5721);
xnor U6437 (N_6437,N_5801,N_5927);
or U6438 (N_6438,N_5701,N_5590);
nand U6439 (N_6439,N_5762,N_5714);
and U6440 (N_6440,N_5526,N_5765);
nand U6441 (N_6441,N_5747,N_5955);
and U6442 (N_6442,N_5576,N_5948);
nor U6443 (N_6443,N_5556,N_5744);
xnor U6444 (N_6444,N_5844,N_5558);
nand U6445 (N_6445,N_5809,N_5880);
and U6446 (N_6446,N_5762,N_5786);
xnor U6447 (N_6447,N_5515,N_5900);
nand U6448 (N_6448,N_5691,N_5701);
nand U6449 (N_6449,N_5957,N_5920);
or U6450 (N_6450,N_5880,N_5958);
or U6451 (N_6451,N_5818,N_5553);
or U6452 (N_6452,N_5874,N_5594);
nand U6453 (N_6453,N_5787,N_5843);
xnor U6454 (N_6454,N_5838,N_5979);
nor U6455 (N_6455,N_5804,N_5990);
nor U6456 (N_6456,N_5905,N_5647);
nor U6457 (N_6457,N_5983,N_5851);
xor U6458 (N_6458,N_5500,N_5742);
xor U6459 (N_6459,N_5832,N_5841);
or U6460 (N_6460,N_5753,N_5919);
xnor U6461 (N_6461,N_5905,N_5574);
and U6462 (N_6462,N_5916,N_5712);
and U6463 (N_6463,N_5985,N_5543);
nand U6464 (N_6464,N_5978,N_5723);
or U6465 (N_6465,N_5521,N_5908);
or U6466 (N_6466,N_5732,N_5702);
or U6467 (N_6467,N_5950,N_5568);
xnor U6468 (N_6468,N_5830,N_5873);
xnor U6469 (N_6469,N_5561,N_5652);
or U6470 (N_6470,N_5516,N_5734);
nor U6471 (N_6471,N_5917,N_5957);
xnor U6472 (N_6472,N_5559,N_5614);
and U6473 (N_6473,N_5921,N_5926);
xnor U6474 (N_6474,N_5592,N_5771);
nand U6475 (N_6475,N_5881,N_5996);
nor U6476 (N_6476,N_5732,N_5855);
nand U6477 (N_6477,N_5968,N_5694);
or U6478 (N_6478,N_5721,N_5693);
xor U6479 (N_6479,N_5720,N_5621);
and U6480 (N_6480,N_5560,N_5987);
nand U6481 (N_6481,N_5506,N_5655);
or U6482 (N_6482,N_5902,N_5792);
nand U6483 (N_6483,N_5748,N_5713);
nand U6484 (N_6484,N_5644,N_5709);
or U6485 (N_6485,N_5621,N_5846);
nand U6486 (N_6486,N_5512,N_5951);
nor U6487 (N_6487,N_5595,N_5986);
nand U6488 (N_6488,N_5703,N_5572);
xor U6489 (N_6489,N_5703,N_5960);
or U6490 (N_6490,N_5619,N_5568);
or U6491 (N_6491,N_5879,N_5963);
and U6492 (N_6492,N_5755,N_5977);
nand U6493 (N_6493,N_5970,N_5512);
nand U6494 (N_6494,N_5729,N_5514);
nor U6495 (N_6495,N_5762,N_5727);
xor U6496 (N_6496,N_5755,N_5686);
xor U6497 (N_6497,N_5991,N_5815);
xor U6498 (N_6498,N_5619,N_5869);
nor U6499 (N_6499,N_5578,N_5945);
nand U6500 (N_6500,N_6065,N_6187);
xor U6501 (N_6501,N_6202,N_6472);
and U6502 (N_6502,N_6006,N_6115);
and U6503 (N_6503,N_6314,N_6124);
nor U6504 (N_6504,N_6342,N_6145);
xor U6505 (N_6505,N_6455,N_6397);
xor U6506 (N_6506,N_6110,N_6064);
or U6507 (N_6507,N_6400,N_6450);
nor U6508 (N_6508,N_6201,N_6204);
nor U6509 (N_6509,N_6088,N_6381);
nand U6510 (N_6510,N_6066,N_6112);
nand U6511 (N_6511,N_6285,N_6206);
xor U6512 (N_6512,N_6434,N_6490);
or U6513 (N_6513,N_6337,N_6485);
or U6514 (N_6514,N_6410,N_6248);
nor U6515 (N_6515,N_6407,N_6362);
xnor U6516 (N_6516,N_6002,N_6144);
nor U6517 (N_6517,N_6041,N_6383);
nand U6518 (N_6518,N_6252,N_6325);
xor U6519 (N_6519,N_6322,N_6469);
nand U6520 (N_6520,N_6113,N_6474);
or U6521 (N_6521,N_6104,N_6331);
nand U6522 (N_6522,N_6213,N_6257);
or U6523 (N_6523,N_6108,N_6329);
xnor U6524 (N_6524,N_6412,N_6173);
and U6525 (N_6525,N_6441,N_6417);
nor U6526 (N_6526,N_6424,N_6009);
or U6527 (N_6527,N_6270,N_6323);
and U6528 (N_6528,N_6050,N_6121);
nor U6529 (N_6529,N_6493,N_6142);
nand U6530 (N_6530,N_6303,N_6376);
nor U6531 (N_6531,N_6157,N_6276);
xnor U6532 (N_6532,N_6404,N_6373);
nand U6533 (N_6533,N_6127,N_6289);
and U6534 (N_6534,N_6359,N_6226);
and U6535 (N_6535,N_6413,N_6191);
nor U6536 (N_6536,N_6245,N_6258);
and U6537 (N_6537,N_6052,N_6176);
and U6538 (N_6538,N_6347,N_6100);
nor U6539 (N_6539,N_6487,N_6463);
nand U6540 (N_6540,N_6229,N_6475);
nor U6541 (N_6541,N_6156,N_6097);
or U6542 (N_6542,N_6221,N_6132);
nand U6543 (N_6543,N_6465,N_6283);
nand U6544 (N_6544,N_6265,N_6272);
xnor U6545 (N_6545,N_6266,N_6171);
nand U6546 (N_6546,N_6334,N_6443);
and U6547 (N_6547,N_6357,N_6260);
and U6548 (N_6548,N_6042,N_6014);
or U6549 (N_6549,N_6330,N_6162);
nor U6550 (N_6550,N_6118,N_6195);
and U6551 (N_6551,N_6131,N_6205);
or U6552 (N_6552,N_6192,N_6479);
nand U6553 (N_6553,N_6136,N_6354);
and U6554 (N_6554,N_6125,N_6387);
nand U6555 (N_6555,N_6103,N_6483);
nor U6556 (N_6556,N_6382,N_6054);
nand U6557 (N_6557,N_6175,N_6083);
or U6558 (N_6558,N_6003,N_6246);
nor U6559 (N_6559,N_6222,N_6232);
and U6560 (N_6560,N_6236,N_6071);
or U6561 (N_6561,N_6188,N_6420);
xor U6562 (N_6562,N_6026,N_6369);
nand U6563 (N_6563,N_6025,N_6250);
and U6564 (N_6564,N_6489,N_6361);
and U6565 (N_6565,N_6370,N_6279);
or U6566 (N_6566,N_6317,N_6137);
and U6567 (N_6567,N_6119,N_6299);
nor U6568 (N_6568,N_6368,N_6253);
nor U6569 (N_6569,N_6148,N_6307);
nand U6570 (N_6570,N_6291,N_6169);
nor U6571 (N_6571,N_6254,N_6320);
xor U6572 (N_6572,N_6379,N_6012);
nor U6573 (N_6573,N_6461,N_6480);
xor U6574 (N_6574,N_6139,N_6034);
xor U6575 (N_6575,N_6101,N_6219);
and U6576 (N_6576,N_6020,N_6439);
and U6577 (N_6577,N_6231,N_6084);
xnor U6578 (N_6578,N_6149,N_6055);
nand U6579 (N_6579,N_6058,N_6073);
nor U6580 (N_6580,N_6238,N_6053);
and U6581 (N_6581,N_6095,N_6022);
and U6582 (N_6582,N_6341,N_6416);
nand U6583 (N_6583,N_6288,N_6099);
or U6584 (N_6584,N_6405,N_6301);
or U6585 (N_6585,N_6399,N_6004);
and U6586 (N_6586,N_6349,N_6212);
nand U6587 (N_6587,N_6167,N_6306);
and U6588 (N_6588,N_6074,N_6182);
xor U6589 (N_6589,N_6057,N_6464);
or U6590 (N_6590,N_6403,N_6384);
nor U6591 (N_6591,N_6059,N_6114);
xnor U6592 (N_6592,N_6215,N_6036);
and U6593 (N_6593,N_6146,N_6249);
xnor U6594 (N_6594,N_6478,N_6079);
nand U6595 (N_6595,N_6346,N_6076);
nor U6596 (N_6596,N_6315,N_6126);
xor U6597 (N_6597,N_6452,N_6363);
nand U6598 (N_6598,N_6378,N_6459);
and U6599 (N_6599,N_6286,N_6326);
or U6600 (N_6600,N_6080,N_6495);
xor U6601 (N_6601,N_6062,N_6085);
and U6602 (N_6602,N_6388,N_6391);
nor U6603 (N_6603,N_6094,N_6335);
xnor U6604 (N_6604,N_6220,N_6154);
xnor U6605 (N_6605,N_6482,N_6268);
xnor U6606 (N_6606,N_6198,N_6300);
nand U6607 (N_6607,N_6061,N_6210);
nand U6608 (N_6608,N_6197,N_6375);
or U6609 (N_6609,N_6040,N_6422);
xnor U6610 (N_6610,N_6230,N_6029);
xor U6611 (N_6611,N_6409,N_6189);
or U6612 (N_6612,N_6395,N_6484);
nor U6613 (N_6613,N_6389,N_6033);
xor U6614 (N_6614,N_6351,N_6273);
or U6615 (N_6615,N_6164,N_6348);
or U6616 (N_6616,N_6393,N_6292);
nand U6617 (N_6617,N_6355,N_6454);
xnor U6618 (N_6618,N_6045,N_6037);
or U6619 (N_6619,N_6128,N_6043);
nand U6620 (N_6620,N_6366,N_6332);
nand U6621 (N_6621,N_6287,N_6435);
xor U6622 (N_6622,N_6486,N_6406);
xnor U6623 (N_6623,N_6150,N_6122);
nor U6624 (N_6624,N_6244,N_6436);
or U6625 (N_6625,N_6430,N_6470);
xor U6626 (N_6626,N_6089,N_6000);
nor U6627 (N_6627,N_6177,N_6019);
or U6628 (N_6628,N_6023,N_6477);
xor U6629 (N_6629,N_6001,N_6186);
and U6630 (N_6630,N_6365,N_6234);
and U6631 (N_6631,N_6318,N_6081);
and U6632 (N_6632,N_6179,N_6310);
nor U6633 (N_6633,N_6093,N_6488);
xnor U6634 (N_6634,N_6111,N_6432);
nor U6635 (N_6635,N_6135,N_6467);
nor U6636 (N_6636,N_6466,N_6374);
xor U6637 (N_6637,N_6453,N_6421);
nor U6638 (N_6638,N_6415,N_6345);
or U6639 (N_6639,N_6224,N_6172);
and U6640 (N_6640,N_6183,N_6414);
and U6641 (N_6641,N_6377,N_6242);
and U6642 (N_6642,N_6274,N_6446);
nand U6643 (N_6643,N_6438,N_6158);
or U6644 (N_6644,N_6035,N_6163);
or U6645 (N_6645,N_6178,N_6056);
nor U6646 (N_6646,N_6471,N_6473);
or U6647 (N_6647,N_6476,N_6356);
nand U6648 (N_6648,N_6321,N_6098);
or U6649 (N_6649,N_6067,N_6380);
and U6650 (N_6650,N_6336,N_6308);
xnor U6651 (N_6651,N_6251,N_6030);
or U6652 (N_6652,N_6394,N_6401);
nor U6653 (N_6653,N_6063,N_6133);
or U6654 (N_6654,N_6116,N_6046);
xor U6655 (N_6655,N_6199,N_6151);
or U6656 (N_6656,N_6225,N_6105);
and U6657 (N_6657,N_6134,N_6358);
and U6658 (N_6658,N_6256,N_6130);
nand U6659 (N_6659,N_6264,N_6051);
nand U6660 (N_6660,N_6075,N_6106);
nand U6661 (N_6661,N_6423,N_6143);
and U6662 (N_6662,N_6174,N_6155);
nand U6663 (N_6663,N_6316,N_6181);
nand U6664 (N_6664,N_6385,N_6360);
xnor U6665 (N_6665,N_6492,N_6497);
nand U6666 (N_6666,N_6458,N_6072);
xor U6667 (N_6667,N_6352,N_6223);
nand U6668 (N_6668,N_6152,N_6196);
or U6669 (N_6669,N_6218,N_6281);
nand U6670 (N_6670,N_6457,N_6109);
or U6671 (N_6671,N_6091,N_6038);
nand U6672 (N_6672,N_6451,N_6239);
and U6673 (N_6673,N_6305,N_6275);
xor U6674 (N_6674,N_6203,N_6429);
and U6675 (N_6675,N_6010,N_6468);
and U6676 (N_6676,N_6092,N_6017);
nor U6677 (N_6677,N_6324,N_6185);
nor U6678 (N_6678,N_6447,N_6170);
xnor U6679 (N_6679,N_6298,N_6462);
and U6680 (N_6680,N_6442,N_6312);
xnor U6681 (N_6681,N_6364,N_6096);
xor U6682 (N_6682,N_6005,N_6294);
or U6683 (N_6683,N_6241,N_6214);
nor U6684 (N_6684,N_6240,N_6481);
nor U6685 (N_6685,N_6184,N_6193);
nor U6686 (N_6686,N_6237,N_6090);
and U6687 (N_6687,N_6070,N_6044);
or U6688 (N_6688,N_6491,N_6433);
nor U6689 (N_6689,N_6086,N_6418);
and U6690 (N_6690,N_6069,N_6015);
and U6691 (N_6691,N_6117,N_6319);
nor U6692 (N_6692,N_6078,N_6428);
xor U6693 (N_6693,N_6333,N_6102);
nor U6694 (N_6694,N_6190,N_6153);
or U6695 (N_6695,N_6243,N_6129);
nand U6696 (N_6696,N_6261,N_6209);
and U6697 (N_6697,N_6278,N_6311);
and U6698 (N_6698,N_6018,N_6343);
and U6699 (N_6699,N_6233,N_6340);
nand U6700 (N_6700,N_6448,N_6262);
nor U6701 (N_6701,N_6168,N_6284);
nor U6702 (N_6702,N_6228,N_6082);
nor U6703 (N_6703,N_6039,N_6328);
nor U6704 (N_6704,N_6295,N_6293);
nand U6705 (N_6705,N_6445,N_6159);
nor U6706 (N_6706,N_6302,N_6499);
or U6707 (N_6707,N_6207,N_6049);
nor U6708 (N_6708,N_6280,N_6024);
xnor U6709 (N_6709,N_6032,N_6267);
or U6710 (N_6710,N_6277,N_6269);
nand U6711 (N_6711,N_6216,N_6255);
and U6712 (N_6712,N_6077,N_6282);
xnor U6713 (N_6713,N_6160,N_6297);
xor U6714 (N_6714,N_6408,N_6498);
nand U6715 (N_6715,N_6371,N_6211);
or U6716 (N_6716,N_6263,N_6016);
and U6717 (N_6717,N_6344,N_6427);
nor U6718 (N_6718,N_6031,N_6217);
xor U6719 (N_6719,N_6367,N_6437);
or U6720 (N_6720,N_6194,N_6313);
nor U6721 (N_6721,N_6008,N_6247);
and U6722 (N_6722,N_6147,N_6426);
and U6723 (N_6723,N_6296,N_6165);
nand U6724 (N_6724,N_6166,N_6123);
nand U6725 (N_6725,N_6290,N_6327);
xor U6726 (N_6726,N_6140,N_6411);
nand U6727 (N_6727,N_6259,N_6390);
nor U6728 (N_6728,N_6011,N_6460);
nand U6729 (N_6729,N_6386,N_6141);
and U6730 (N_6730,N_6007,N_6309);
and U6731 (N_6731,N_6496,N_6444);
nor U6732 (N_6732,N_6350,N_6494);
xnor U6733 (N_6733,N_6208,N_6087);
xnor U6734 (N_6734,N_6402,N_6027);
or U6735 (N_6735,N_6227,N_6068);
and U6736 (N_6736,N_6138,N_6372);
and U6737 (N_6737,N_6398,N_6271);
or U6738 (N_6738,N_6028,N_6419);
nand U6739 (N_6739,N_6339,N_6200);
and U6740 (N_6740,N_6180,N_6107);
and U6741 (N_6741,N_6060,N_6048);
nand U6742 (N_6742,N_6392,N_6021);
nor U6743 (N_6743,N_6449,N_6120);
nor U6744 (N_6744,N_6431,N_6161);
or U6745 (N_6745,N_6338,N_6235);
or U6746 (N_6746,N_6440,N_6456);
and U6747 (N_6747,N_6304,N_6353);
nand U6748 (N_6748,N_6425,N_6013);
nand U6749 (N_6749,N_6047,N_6396);
nor U6750 (N_6750,N_6200,N_6487);
xor U6751 (N_6751,N_6256,N_6212);
nand U6752 (N_6752,N_6119,N_6261);
xnor U6753 (N_6753,N_6445,N_6387);
nor U6754 (N_6754,N_6253,N_6098);
nand U6755 (N_6755,N_6272,N_6386);
and U6756 (N_6756,N_6194,N_6424);
or U6757 (N_6757,N_6360,N_6011);
nor U6758 (N_6758,N_6109,N_6448);
and U6759 (N_6759,N_6161,N_6342);
nand U6760 (N_6760,N_6430,N_6398);
or U6761 (N_6761,N_6231,N_6335);
or U6762 (N_6762,N_6218,N_6349);
xnor U6763 (N_6763,N_6185,N_6385);
nand U6764 (N_6764,N_6323,N_6476);
nand U6765 (N_6765,N_6242,N_6275);
and U6766 (N_6766,N_6134,N_6477);
or U6767 (N_6767,N_6021,N_6037);
nand U6768 (N_6768,N_6306,N_6082);
and U6769 (N_6769,N_6414,N_6287);
xnor U6770 (N_6770,N_6443,N_6144);
xor U6771 (N_6771,N_6000,N_6065);
and U6772 (N_6772,N_6417,N_6493);
nand U6773 (N_6773,N_6250,N_6203);
and U6774 (N_6774,N_6463,N_6358);
or U6775 (N_6775,N_6408,N_6093);
or U6776 (N_6776,N_6195,N_6175);
or U6777 (N_6777,N_6476,N_6148);
nor U6778 (N_6778,N_6449,N_6448);
nand U6779 (N_6779,N_6117,N_6285);
and U6780 (N_6780,N_6177,N_6261);
xor U6781 (N_6781,N_6392,N_6390);
nand U6782 (N_6782,N_6485,N_6054);
or U6783 (N_6783,N_6404,N_6268);
nor U6784 (N_6784,N_6387,N_6262);
xor U6785 (N_6785,N_6458,N_6446);
and U6786 (N_6786,N_6190,N_6237);
or U6787 (N_6787,N_6408,N_6073);
nor U6788 (N_6788,N_6451,N_6180);
and U6789 (N_6789,N_6146,N_6244);
xnor U6790 (N_6790,N_6207,N_6237);
xnor U6791 (N_6791,N_6140,N_6478);
and U6792 (N_6792,N_6222,N_6328);
nor U6793 (N_6793,N_6436,N_6125);
or U6794 (N_6794,N_6118,N_6270);
and U6795 (N_6795,N_6338,N_6005);
nor U6796 (N_6796,N_6273,N_6228);
nand U6797 (N_6797,N_6187,N_6339);
nor U6798 (N_6798,N_6348,N_6014);
and U6799 (N_6799,N_6156,N_6410);
or U6800 (N_6800,N_6153,N_6125);
or U6801 (N_6801,N_6213,N_6134);
nand U6802 (N_6802,N_6040,N_6085);
and U6803 (N_6803,N_6025,N_6365);
xnor U6804 (N_6804,N_6357,N_6128);
and U6805 (N_6805,N_6091,N_6370);
nand U6806 (N_6806,N_6415,N_6011);
and U6807 (N_6807,N_6060,N_6347);
nand U6808 (N_6808,N_6344,N_6381);
or U6809 (N_6809,N_6490,N_6358);
or U6810 (N_6810,N_6452,N_6275);
nor U6811 (N_6811,N_6279,N_6293);
and U6812 (N_6812,N_6490,N_6079);
nor U6813 (N_6813,N_6489,N_6088);
and U6814 (N_6814,N_6306,N_6039);
or U6815 (N_6815,N_6128,N_6445);
xor U6816 (N_6816,N_6332,N_6379);
and U6817 (N_6817,N_6170,N_6472);
nand U6818 (N_6818,N_6160,N_6134);
or U6819 (N_6819,N_6036,N_6356);
nand U6820 (N_6820,N_6057,N_6141);
or U6821 (N_6821,N_6383,N_6316);
xnor U6822 (N_6822,N_6417,N_6414);
or U6823 (N_6823,N_6345,N_6286);
nand U6824 (N_6824,N_6081,N_6160);
and U6825 (N_6825,N_6232,N_6277);
or U6826 (N_6826,N_6139,N_6293);
and U6827 (N_6827,N_6124,N_6417);
nor U6828 (N_6828,N_6064,N_6034);
xor U6829 (N_6829,N_6001,N_6343);
nand U6830 (N_6830,N_6427,N_6361);
and U6831 (N_6831,N_6298,N_6438);
and U6832 (N_6832,N_6254,N_6313);
nor U6833 (N_6833,N_6146,N_6168);
and U6834 (N_6834,N_6397,N_6247);
and U6835 (N_6835,N_6133,N_6306);
or U6836 (N_6836,N_6258,N_6181);
or U6837 (N_6837,N_6280,N_6058);
xnor U6838 (N_6838,N_6207,N_6227);
nand U6839 (N_6839,N_6150,N_6099);
or U6840 (N_6840,N_6466,N_6023);
nand U6841 (N_6841,N_6326,N_6259);
xnor U6842 (N_6842,N_6255,N_6156);
xor U6843 (N_6843,N_6213,N_6039);
nor U6844 (N_6844,N_6154,N_6455);
or U6845 (N_6845,N_6287,N_6103);
xor U6846 (N_6846,N_6319,N_6480);
nor U6847 (N_6847,N_6243,N_6362);
nor U6848 (N_6848,N_6051,N_6411);
nor U6849 (N_6849,N_6358,N_6056);
xnor U6850 (N_6850,N_6460,N_6144);
xnor U6851 (N_6851,N_6052,N_6391);
xnor U6852 (N_6852,N_6008,N_6198);
or U6853 (N_6853,N_6101,N_6036);
nand U6854 (N_6854,N_6252,N_6269);
nand U6855 (N_6855,N_6060,N_6097);
nand U6856 (N_6856,N_6097,N_6030);
and U6857 (N_6857,N_6026,N_6109);
or U6858 (N_6858,N_6255,N_6115);
or U6859 (N_6859,N_6218,N_6391);
xnor U6860 (N_6860,N_6222,N_6304);
or U6861 (N_6861,N_6049,N_6204);
nor U6862 (N_6862,N_6002,N_6062);
xnor U6863 (N_6863,N_6270,N_6495);
nand U6864 (N_6864,N_6116,N_6103);
or U6865 (N_6865,N_6360,N_6103);
or U6866 (N_6866,N_6231,N_6175);
nand U6867 (N_6867,N_6447,N_6289);
and U6868 (N_6868,N_6138,N_6307);
and U6869 (N_6869,N_6261,N_6017);
and U6870 (N_6870,N_6071,N_6162);
and U6871 (N_6871,N_6432,N_6364);
or U6872 (N_6872,N_6157,N_6124);
and U6873 (N_6873,N_6377,N_6245);
or U6874 (N_6874,N_6346,N_6290);
nand U6875 (N_6875,N_6115,N_6025);
and U6876 (N_6876,N_6077,N_6429);
nor U6877 (N_6877,N_6268,N_6058);
or U6878 (N_6878,N_6279,N_6479);
and U6879 (N_6879,N_6201,N_6060);
xor U6880 (N_6880,N_6025,N_6428);
nand U6881 (N_6881,N_6282,N_6248);
nor U6882 (N_6882,N_6314,N_6267);
xor U6883 (N_6883,N_6036,N_6343);
xor U6884 (N_6884,N_6202,N_6216);
and U6885 (N_6885,N_6036,N_6405);
nand U6886 (N_6886,N_6496,N_6400);
nor U6887 (N_6887,N_6016,N_6027);
nand U6888 (N_6888,N_6418,N_6286);
or U6889 (N_6889,N_6166,N_6103);
or U6890 (N_6890,N_6134,N_6034);
nand U6891 (N_6891,N_6005,N_6445);
nor U6892 (N_6892,N_6243,N_6434);
nor U6893 (N_6893,N_6073,N_6218);
nand U6894 (N_6894,N_6484,N_6411);
nor U6895 (N_6895,N_6455,N_6096);
nor U6896 (N_6896,N_6494,N_6423);
and U6897 (N_6897,N_6335,N_6397);
or U6898 (N_6898,N_6394,N_6235);
xnor U6899 (N_6899,N_6029,N_6224);
xnor U6900 (N_6900,N_6144,N_6140);
nand U6901 (N_6901,N_6412,N_6002);
nand U6902 (N_6902,N_6115,N_6366);
nor U6903 (N_6903,N_6015,N_6153);
xnor U6904 (N_6904,N_6080,N_6276);
or U6905 (N_6905,N_6189,N_6051);
or U6906 (N_6906,N_6234,N_6436);
or U6907 (N_6907,N_6112,N_6054);
xor U6908 (N_6908,N_6065,N_6334);
and U6909 (N_6909,N_6359,N_6267);
xor U6910 (N_6910,N_6240,N_6077);
xnor U6911 (N_6911,N_6434,N_6482);
nand U6912 (N_6912,N_6010,N_6003);
nand U6913 (N_6913,N_6082,N_6226);
or U6914 (N_6914,N_6006,N_6047);
and U6915 (N_6915,N_6309,N_6459);
nand U6916 (N_6916,N_6067,N_6428);
xnor U6917 (N_6917,N_6017,N_6476);
or U6918 (N_6918,N_6020,N_6193);
or U6919 (N_6919,N_6276,N_6491);
and U6920 (N_6920,N_6200,N_6173);
nor U6921 (N_6921,N_6426,N_6099);
nand U6922 (N_6922,N_6466,N_6220);
and U6923 (N_6923,N_6057,N_6143);
xor U6924 (N_6924,N_6209,N_6306);
or U6925 (N_6925,N_6185,N_6110);
and U6926 (N_6926,N_6084,N_6228);
and U6927 (N_6927,N_6057,N_6197);
xnor U6928 (N_6928,N_6093,N_6012);
or U6929 (N_6929,N_6208,N_6181);
nand U6930 (N_6930,N_6234,N_6273);
and U6931 (N_6931,N_6415,N_6486);
nand U6932 (N_6932,N_6297,N_6465);
and U6933 (N_6933,N_6392,N_6291);
and U6934 (N_6934,N_6074,N_6115);
and U6935 (N_6935,N_6203,N_6495);
and U6936 (N_6936,N_6487,N_6329);
nand U6937 (N_6937,N_6107,N_6339);
or U6938 (N_6938,N_6106,N_6042);
or U6939 (N_6939,N_6317,N_6245);
xnor U6940 (N_6940,N_6239,N_6010);
nand U6941 (N_6941,N_6328,N_6336);
or U6942 (N_6942,N_6480,N_6129);
nand U6943 (N_6943,N_6242,N_6364);
or U6944 (N_6944,N_6033,N_6290);
or U6945 (N_6945,N_6242,N_6241);
and U6946 (N_6946,N_6038,N_6451);
nand U6947 (N_6947,N_6371,N_6376);
nand U6948 (N_6948,N_6468,N_6228);
nor U6949 (N_6949,N_6129,N_6063);
and U6950 (N_6950,N_6132,N_6251);
nor U6951 (N_6951,N_6165,N_6026);
and U6952 (N_6952,N_6155,N_6352);
xor U6953 (N_6953,N_6069,N_6048);
xnor U6954 (N_6954,N_6128,N_6428);
and U6955 (N_6955,N_6321,N_6271);
xor U6956 (N_6956,N_6341,N_6393);
or U6957 (N_6957,N_6292,N_6108);
nor U6958 (N_6958,N_6364,N_6054);
xnor U6959 (N_6959,N_6280,N_6347);
and U6960 (N_6960,N_6037,N_6040);
or U6961 (N_6961,N_6482,N_6488);
nor U6962 (N_6962,N_6329,N_6335);
or U6963 (N_6963,N_6478,N_6337);
nor U6964 (N_6964,N_6194,N_6008);
or U6965 (N_6965,N_6230,N_6016);
xor U6966 (N_6966,N_6474,N_6200);
and U6967 (N_6967,N_6485,N_6142);
xor U6968 (N_6968,N_6390,N_6062);
nand U6969 (N_6969,N_6256,N_6016);
and U6970 (N_6970,N_6471,N_6046);
xor U6971 (N_6971,N_6040,N_6390);
xor U6972 (N_6972,N_6244,N_6240);
or U6973 (N_6973,N_6197,N_6182);
and U6974 (N_6974,N_6108,N_6303);
xor U6975 (N_6975,N_6100,N_6209);
nand U6976 (N_6976,N_6463,N_6416);
nand U6977 (N_6977,N_6137,N_6453);
nor U6978 (N_6978,N_6326,N_6428);
or U6979 (N_6979,N_6420,N_6204);
nor U6980 (N_6980,N_6490,N_6415);
nand U6981 (N_6981,N_6038,N_6342);
nor U6982 (N_6982,N_6049,N_6407);
or U6983 (N_6983,N_6485,N_6043);
xor U6984 (N_6984,N_6112,N_6169);
and U6985 (N_6985,N_6038,N_6200);
or U6986 (N_6986,N_6317,N_6026);
xnor U6987 (N_6987,N_6106,N_6438);
or U6988 (N_6988,N_6062,N_6141);
and U6989 (N_6989,N_6478,N_6137);
and U6990 (N_6990,N_6076,N_6439);
xor U6991 (N_6991,N_6115,N_6197);
or U6992 (N_6992,N_6417,N_6269);
xor U6993 (N_6993,N_6251,N_6040);
or U6994 (N_6994,N_6137,N_6152);
and U6995 (N_6995,N_6255,N_6024);
and U6996 (N_6996,N_6207,N_6292);
xor U6997 (N_6997,N_6087,N_6139);
and U6998 (N_6998,N_6226,N_6320);
or U6999 (N_6999,N_6487,N_6131);
or U7000 (N_7000,N_6751,N_6847);
and U7001 (N_7001,N_6698,N_6854);
or U7002 (N_7002,N_6578,N_6850);
xnor U7003 (N_7003,N_6870,N_6755);
nand U7004 (N_7004,N_6685,N_6846);
nand U7005 (N_7005,N_6745,N_6945);
and U7006 (N_7006,N_6862,N_6828);
xor U7007 (N_7007,N_6707,N_6598);
or U7008 (N_7008,N_6793,N_6797);
nor U7009 (N_7009,N_6577,N_6894);
nand U7010 (N_7010,N_6597,N_6939);
and U7011 (N_7011,N_6938,N_6557);
nor U7012 (N_7012,N_6771,N_6530);
and U7013 (N_7013,N_6822,N_6809);
nand U7014 (N_7014,N_6558,N_6935);
and U7015 (N_7015,N_6692,N_6853);
or U7016 (N_7016,N_6629,N_6591);
and U7017 (N_7017,N_6515,N_6933);
xor U7018 (N_7018,N_6959,N_6571);
and U7019 (N_7019,N_6925,N_6602);
nor U7020 (N_7020,N_6815,N_6690);
xnor U7021 (N_7021,N_6756,N_6529);
xor U7022 (N_7022,N_6647,N_6914);
and U7023 (N_7023,N_6615,N_6583);
xor U7024 (N_7024,N_6735,N_6812);
nand U7025 (N_7025,N_6818,N_6523);
xnor U7026 (N_7026,N_6506,N_6930);
nand U7027 (N_7027,N_6689,N_6540);
xor U7028 (N_7028,N_6678,N_6898);
xor U7029 (N_7029,N_6741,N_6669);
nor U7030 (N_7030,N_6842,N_6527);
nor U7031 (N_7031,N_6572,N_6519);
nand U7032 (N_7032,N_6663,N_6642);
nor U7033 (N_7033,N_6638,N_6708);
xnor U7034 (N_7034,N_6702,N_6559);
xnor U7035 (N_7035,N_6710,N_6623);
nor U7036 (N_7036,N_6758,N_6625);
xor U7037 (N_7037,N_6510,N_6538);
nor U7038 (N_7038,N_6810,N_6727);
nor U7039 (N_7039,N_6721,N_6742);
nand U7040 (N_7040,N_6730,N_6582);
xor U7041 (N_7041,N_6997,N_6715);
or U7042 (N_7042,N_6592,N_6525);
nand U7043 (N_7043,N_6973,N_6608);
and U7044 (N_7044,N_6983,N_6979);
or U7045 (N_7045,N_6986,N_6521);
and U7046 (N_7046,N_6993,N_6995);
nand U7047 (N_7047,N_6603,N_6605);
nand U7048 (N_7048,N_6996,N_6990);
and U7049 (N_7049,N_6904,N_6693);
nor U7050 (N_7050,N_6680,N_6874);
or U7051 (N_7051,N_6790,N_6794);
nand U7052 (N_7052,N_6942,N_6588);
or U7053 (N_7053,N_6891,N_6932);
nand U7054 (N_7054,N_6585,N_6550);
nand U7055 (N_7055,N_6596,N_6770);
nor U7056 (N_7056,N_6507,N_6781);
xor U7057 (N_7057,N_6576,N_6561);
nor U7058 (N_7058,N_6569,N_6662);
nand U7059 (N_7059,N_6875,N_6985);
nand U7060 (N_7060,N_6813,N_6711);
or U7061 (N_7061,N_6590,N_6659);
xor U7062 (N_7062,N_6726,N_6970);
nand U7063 (N_7063,N_6841,N_6881);
and U7064 (N_7064,N_6746,N_6518);
nand U7065 (N_7065,N_6859,N_6673);
and U7066 (N_7066,N_6505,N_6921);
nand U7067 (N_7067,N_6792,N_6587);
and U7068 (N_7068,N_6636,N_6593);
nor U7069 (N_7069,N_6905,N_6574);
and U7070 (N_7070,N_6533,N_6757);
xnor U7071 (N_7071,N_6691,N_6668);
nor U7072 (N_7072,N_6974,N_6762);
or U7073 (N_7073,N_6754,N_6796);
xor U7074 (N_7074,N_6806,N_6998);
or U7075 (N_7075,N_6761,N_6618);
xnor U7076 (N_7076,N_6679,N_6500);
and U7077 (N_7077,N_6705,N_6944);
nor U7078 (N_7078,N_6830,N_6736);
and U7079 (N_7079,N_6729,N_6855);
or U7080 (N_7080,N_6982,N_6612);
and U7081 (N_7081,N_6575,N_6787);
or U7082 (N_7082,N_6720,N_6706);
or U7083 (N_7083,N_6972,N_6656);
and U7084 (N_7084,N_6934,N_6980);
nand U7085 (N_7085,N_6873,N_6728);
xor U7086 (N_7086,N_6660,N_6774);
nor U7087 (N_7087,N_6955,N_6917);
and U7088 (N_7088,N_6637,N_6633);
nand U7089 (N_7089,N_6991,N_6851);
and U7090 (N_7090,N_6641,N_6544);
nand U7091 (N_7091,N_6655,N_6632);
or U7092 (N_7092,N_6867,N_6611);
and U7093 (N_7093,N_6789,N_6562);
and U7094 (N_7094,N_6504,N_6564);
or U7095 (N_7095,N_6665,N_6791);
nand U7096 (N_7096,N_6600,N_6560);
or U7097 (N_7097,N_6718,N_6953);
nand U7098 (N_7098,N_6620,N_6878);
and U7099 (N_7099,N_6613,N_6601);
nand U7100 (N_7100,N_6737,N_6956);
nand U7101 (N_7101,N_6951,N_6884);
nor U7102 (N_7102,N_6833,N_6831);
xnor U7103 (N_7103,N_6666,N_6918);
xnor U7104 (N_7104,N_6556,N_6783);
nor U7105 (N_7105,N_6604,N_6906);
nand U7106 (N_7106,N_6614,N_6820);
nor U7107 (N_7107,N_6536,N_6686);
xor U7108 (N_7108,N_6768,N_6976);
and U7109 (N_7109,N_6922,N_6753);
xor U7110 (N_7110,N_6988,N_6606);
xnor U7111 (N_7111,N_6740,N_6816);
or U7112 (N_7112,N_6883,N_6717);
xnor U7113 (N_7113,N_6843,N_6769);
and U7114 (N_7114,N_6779,N_6539);
and U7115 (N_7115,N_6724,N_6826);
nor U7116 (N_7116,N_6520,N_6936);
xor U7117 (N_7117,N_6941,N_6908);
nand U7118 (N_7118,N_6900,N_6772);
and U7119 (N_7119,N_6897,N_6876);
and U7120 (N_7120,N_6916,N_6651);
xnor U7121 (N_7121,N_6967,N_6927);
nor U7122 (N_7122,N_6631,N_6554);
nor U7123 (N_7123,N_6889,N_6759);
nor U7124 (N_7124,N_6987,N_6915);
nor U7125 (N_7125,N_6803,N_6895);
nor U7126 (N_7126,N_6716,N_6675);
or U7127 (N_7127,N_6589,N_6682);
xor U7128 (N_7128,N_6640,N_6750);
xnor U7129 (N_7129,N_6872,N_6627);
nand U7130 (N_7130,N_6885,N_6628);
nor U7131 (N_7131,N_6785,N_6966);
or U7132 (N_7132,N_6526,N_6565);
or U7133 (N_7133,N_6650,N_6825);
xnor U7134 (N_7134,N_6802,N_6634);
nand U7135 (N_7135,N_6765,N_6910);
and U7136 (N_7136,N_6777,N_6667);
xnor U7137 (N_7137,N_6811,N_6681);
nor U7138 (N_7138,N_6528,N_6880);
or U7139 (N_7139,N_6835,N_6952);
and U7140 (N_7140,N_6502,N_6743);
or U7141 (N_7141,N_6767,N_6548);
nand U7142 (N_7142,N_6696,N_6677);
or U7143 (N_7143,N_6929,N_6858);
nor U7144 (N_7144,N_6749,N_6547);
nor U7145 (N_7145,N_6849,N_6857);
nand U7146 (N_7146,N_6819,N_6863);
nor U7147 (N_7147,N_6653,N_6688);
or U7148 (N_7148,N_6645,N_6541);
or U7149 (N_7149,N_6845,N_6896);
xor U7150 (N_7150,N_6760,N_6887);
or U7151 (N_7151,N_6960,N_6657);
xnor U7152 (N_7152,N_6817,N_6839);
nand U7153 (N_7153,N_6840,N_6524);
nor U7154 (N_7154,N_6852,N_6599);
xor U7155 (N_7155,N_6763,N_6643);
nor U7156 (N_7156,N_6782,N_6940);
nor U7157 (N_7157,N_6994,N_6937);
xnor U7158 (N_7158,N_6902,N_6630);
xnor U7159 (N_7159,N_6664,N_6734);
nor U7160 (N_7160,N_6992,N_6617);
and U7161 (N_7161,N_6635,N_6676);
or U7162 (N_7162,N_6732,N_6877);
nand U7163 (N_7163,N_6568,N_6570);
and U7164 (N_7164,N_6701,N_6522);
nand U7165 (N_7165,N_6699,N_6646);
and U7166 (N_7166,N_6860,N_6962);
and U7167 (N_7167,N_6800,N_6981);
or U7168 (N_7168,N_6958,N_6517);
and U7169 (N_7169,N_6713,N_6697);
nand U7170 (N_7170,N_6748,N_6512);
nand U7171 (N_7171,N_6700,N_6695);
nor U7172 (N_7172,N_6581,N_6744);
nor U7173 (N_7173,N_6503,N_6683);
xnor U7174 (N_7174,N_6553,N_6514);
or U7175 (N_7175,N_6924,N_6652);
and U7176 (N_7176,N_6856,N_6829);
xnor U7177 (N_7177,N_6546,N_6892);
nor U7178 (N_7178,N_6607,N_6804);
or U7179 (N_7179,N_6709,N_6871);
and U7180 (N_7180,N_6784,N_6824);
xnor U7181 (N_7181,N_6739,N_6764);
nor U7182 (N_7182,N_6639,N_6622);
nor U7183 (N_7183,N_6722,N_6882);
or U7184 (N_7184,N_6926,N_6658);
and U7185 (N_7185,N_6621,N_6963);
or U7186 (N_7186,N_6965,N_6977);
or U7187 (N_7187,N_6670,N_6532);
or U7188 (N_7188,N_6805,N_6837);
nor U7189 (N_7189,N_6580,N_6516);
nand U7190 (N_7190,N_6555,N_6566);
xor U7191 (N_7191,N_6542,N_6868);
or U7192 (N_7192,N_6671,N_6567);
and U7193 (N_7193,N_6731,N_6594);
and U7194 (N_7194,N_6714,N_6513);
nor U7195 (N_7195,N_6788,N_6869);
or U7196 (N_7196,N_6919,N_6807);
nand U7197 (N_7197,N_6909,N_6511);
or U7198 (N_7198,N_6752,N_6674);
or U7199 (N_7199,N_6694,N_6975);
nand U7200 (N_7200,N_6899,N_6879);
nand U7201 (N_7201,N_6661,N_6961);
and U7202 (N_7202,N_6584,N_6644);
or U7203 (N_7203,N_6537,N_6703);
xnor U7204 (N_7204,N_6733,N_6948);
or U7205 (N_7205,N_6838,N_6920);
or U7206 (N_7206,N_6776,N_6535);
and U7207 (N_7207,N_6866,N_6549);
and U7208 (N_7208,N_6964,N_6672);
nor U7209 (N_7209,N_6801,N_6903);
or U7210 (N_7210,N_6949,N_6684);
xnor U7211 (N_7211,N_6907,N_6719);
nor U7212 (N_7212,N_6999,N_6778);
nor U7213 (N_7213,N_6954,N_6799);
nor U7214 (N_7214,N_6836,N_6648);
and U7215 (N_7215,N_6775,N_6821);
and U7216 (N_7216,N_6971,N_6579);
nand U7217 (N_7217,N_6814,N_6834);
nand U7218 (N_7218,N_6827,N_6534);
and U7219 (N_7219,N_6950,N_6508);
xnor U7220 (N_7220,N_6531,N_6619);
nor U7221 (N_7221,N_6928,N_6780);
and U7222 (N_7222,N_6723,N_6865);
nand U7223 (N_7223,N_6808,N_6563);
or U7224 (N_7224,N_6931,N_6911);
or U7225 (N_7225,N_6704,N_6861);
and U7226 (N_7226,N_6786,N_6823);
nor U7227 (N_7227,N_6616,N_6893);
nor U7228 (N_7228,N_6890,N_6864);
xor U7229 (N_7229,N_6984,N_6844);
or U7230 (N_7230,N_6946,N_6586);
xnor U7231 (N_7231,N_6654,N_6649);
nand U7232 (N_7232,N_6725,N_6798);
nor U7233 (N_7233,N_6947,N_6573);
nor U7234 (N_7234,N_6501,N_6545);
nor U7235 (N_7235,N_6886,N_6912);
xnor U7236 (N_7236,N_6978,N_6595);
xnor U7237 (N_7237,N_6712,N_6989);
xor U7238 (N_7238,N_6773,N_6968);
nor U7239 (N_7239,N_6738,N_6913);
xnor U7240 (N_7240,N_6795,N_6923);
nand U7241 (N_7241,N_6969,N_6832);
xnor U7242 (N_7242,N_6610,N_6509);
xnor U7243 (N_7243,N_6543,N_6551);
and U7244 (N_7244,N_6888,N_6943);
nor U7245 (N_7245,N_6848,N_6626);
xor U7246 (N_7246,N_6747,N_6552);
or U7247 (N_7247,N_6624,N_6687);
or U7248 (N_7248,N_6766,N_6957);
nand U7249 (N_7249,N_6901,N_6609);
and U7250 (N_7250,N_6985,N_6663);
nand U7251 (N_7251,N_6833,N_6881);
and U7252 (N_7252,N_6997,N_6944);
nand U7253 (N_7253,N_6710,N_6939);
or U7254 (N_7254,N_6687,N_6931);
or U7255 (N_7255,N_6617,N_6991);
nor U7256 (N_7256,N_6510,N_6967);
nor U7257 (N_7257,N_6826,N_6636);
or U7258 (N_7258,N_6952,N_6908);
xnor U7259 (N_7259,N_6703,N_6980);
or U7260 (N_7260,N_6983,N_6687);
or U7261 (N_7261,N_6906,N_6891);
nand U7262 (N_7262,N_6880,N_6640);
or U7263 (N_7263,N_6500,N_6690);
xor U7264 (N_7264,N_6533,N_6603);
or U7265 (N_7265,N_6652,N_6804);
or U7266 (N_7266,N_6745,N_6772);
or U7267 (N_7267,N_6538,N_6686);
and U7268 (N_7268,N_6905,N_6612);
and U7269 (N_7269,N_6567,N_6991);
and U7270 (N_7270,N_6712,N_6641);
xor U7271 (N_7271,N_6996,N_6797);
and U7272 (N_7272,N_6921,N_6755);
nand U7273 (N_7273,N_6841,N_6537);
xor U7274 (N_7274,N_6979,N_6691);
nor U7275 (N_7275,N_6516,N_6755);
or U7276 (N_7276,N_6693,N_6960);
xor U7277 (N_7277,N_6736,N_6995);
or U7278 (N_7278,N_6742,N_6971);
xor U7279 (N_7279,N_6894,N_6536);
nor U7280 (N_7280,N_6753,N_6521);
xor U7281 (N_7281,N_6572,N_6700);
and U7282 (N_7282,N_6938,N_6522);
xnor U7283 (N_7283,N_6720,N_6632);
nand U7284 (N_7284,N_6824,N_6906);
or U7285 (N_7285,N_6721,N_6705);
nor U7286 (N_7286,N_6530,N_6662);
and U7287 (N_7287,N_6673,N_6791);
xor U7288 (N_7288,N_6819,N_6515);
or U7289 (N_7289,N_6884,N_6537);
or U7290 (N_7290,N_6594,N_6873);
and U7291 (N_7291,N_6626,N_6939);
nand U7292 (N_7292,N_6511,N_6572);
xnor U7293 (N_7293,N_6906,N_6630);
and U7294 (N_7294,N_6868,N_6806);
or U7295 (N_7295,N_6573,N_6808);
nand U7296 (N_7296,N_6822,N_6500);
and U7297 (N_7297,N_6613,N_6741);
or U7298 (N_7298,N_6604,N_6883);
nand U7299 (N_7299,N_6660,N_6934);
nor U7300 (N_7300,N_6627,N_6798);
or U7301 (N_7301,N_6812,N_6695);
nand U7302 (N_7302,N_6670,N_6601);
or U7303 (N_7303,N_6949,N_6739);
nand U7304 (N_7304,N_6770,N_6962);
nor U7305 (N_7305,N_6915,N_6871);
nand U7306 (N_7306,N_6691,N_6542);
and U7307 (N_7307,N_6641,N_6748);
nor U7308 (N_7308,N_6603,N_6945);
nand U7309 (N_7309,N_6579,N_6787);
xor U7310 (N_7310,N_6924,N_6843);
or U7311 (N_7311,N_6975,N_6946);
or U7312 (N_7312,N_6611,N_6968);
nand U7313 (N_7313,N_6888,N_6845);
or U7314 (N_7314,N_6507,N_6874);
or U7315 (N_7315,N_6530,N_6743);
or U7316 (N_7316,N_6663,N_6762);
xor U7317 (N_7317,N_6573,N_6754);
xnor U7318 (N_7318,N_6729,N_6585);
nand U7319 (N_7319,N_6875,N_6759);
xnor U7320 (N_7320,N_6916,N_6934);
nor U7321 (N_7321,N_6849,N_6650);
and U7322 (N_7322,N_6941,N_6979);
nor U7323 (N_7323,N_6548,N_6926);
and U7324 (N_7324,N_6884,N_6671);
or U7325 (N_7325,N_6621,N_6824);
or U7326 (N_7326,N_6684,N_6978);
xor U7327 (N_7327,N_6961,N_6778);
or U7328 (N_7328,N_6993,N_6964);
or U7329 (N_7329,N_6942,N_6989);
nand U7330 (N_7330,N_6711,N_6789);
nand U7331 (N_7331,N_6894,N_6669);
nor U7332 (N_7332,N_6859,N_6952);
xnor U7333 (N_7333,N_6823,N_6654);
nor U7334 (N_7334,N_6564,N_6975);
and U7335 (N_7335,N_6897,N_6518);
or U7336 (N_7336,N_6625,N_6781);
xnor U7337 (N_7337,N_6681,N_6992);
xor U7338 (N_7338,N_6909,N_6649);
nand U7339 (N_7339,N_6701,N_6752);
nor U7340 (N_7340,N_6553,N_6962);
nand U7341 (N_7341,N_6903,N_6524);
or U7342 (N_7342,N_6922,N_6766);
nor U7343 (N_7343,N_6876,N_6809);
nand U7344 (N_7344,N_6813,N_6883);
nor U7345 (N_7345,N_6579,N_6793);
or U7346 (N_7346,N_6512,N_6978);
xnor U7347 (N_7347,N_6927,N_6586);
nand U7348 (N_7348,N_6736,N_6819);
and U7349 (N_7349,N_6524,N_6863);
or U7350 (N_7350,N_6577,N_6816);
and U7351 (N_7351,N_6846,N_6935);
nor U7352 (N_7352,N_6603,N_6699);
nor U7353 (N_7353,N_6552,N_6649);
nand U7354 (N_7354,N_6811,N_6892);
or U7355 (N_7355,N_6946,N_6839);
and U7356 (N_7356,N_6628,N_6590);
nor U7357 (N_7357,N_6677,N_6770);
or U7358 (N_7358,N_6922,N_6942);
or U7359 (N_7359,N_6922,N_6813);
nand U7360 (N_7360,N_6699,N_6628);
xnor U7361 (N_7361,N_6855,N_6645);
xor U7362 (N_7362,N_6962,N_6541);
and U7363 (N_7363,N_6946,N_6533);
or U7364 (N_7364,N_6787,N_6844);
nand U7365 (N_7365,N_6581,N_6707);
nand U7366 (N_7366,N_6655,N_6959);
and U7367 (N_7367,N_6690,N_6770);
xnor U7368 (N_7368,N_6634,N_6535);
xor U7369 (N_7369,N_6514,N_6965);
nand U7370 (N_7370,N_6949,N_6983);
and U7371 (N_7371,N_6768,N_6729);
and U7372 (N_7372,N_6925,N_6803);
nor U7373 (N_7373,N_6544,N_6513);
xor U7374 (N_7374,N_6673,N_6542);
nor U7375 (N_7375,N_6816,N_6612);
nand U7376 (N_7376,N_6617,N_6996);
xor U7377 (N_7377,N_6975,N_6644);
or U7378 (N_7378,N_6745,N_6564);
or U7379 (N_7379,N_6576,N_6719);
or U7380 (N_7380,N_6568,N_6804);
xnor U7381 (N_7381,N_6714,N_6933);
and U7382 (N_7382,N_6653,N_6593);
or U7383 (N_7383,N_6922,N_6684);
nand U7384 (N_7384,N_6531,N_6814);
nor U7385 (N_7385,N_6605,N_6734);
nor U7386 (N_7386,N_6722,N_6777);
nand U7387 (N_7387,N_6641,N_6596);
xnor U7388 (N_7388,N_6845,N_6753);
xnor U7389 (N_7389,N_6825,N_6972);
xnor U7390 (N_7390,N_6755,N_6761);
xor U7391 (N_7391,N_6768,N_6631);
nand U7392 (N_7392,N_6712,N_6852);
nor U7393 (N_7393,N_6947,N_6671);
or U7394 (N_7394,N_6897,N_6982);
nor U7395 (N_7395,N_6959,N_6738);
and U7396 (N_7396,N_6951,N_6575);
and U7397 (N_7397,N_6611,N_6647);
and U7398 (N_7398,N_6830,N_6928);
or U7399 (N_7399,N_6510,N_6524);
xor U7400 (N_7400,N_6750,N_6895);
or U7401 (N_7401,N_6504,N_6889);
and U7402 (N_7402,N_6983,N_6718);
nor U7403 (N_7403,N_6523,N_6569);
and U7404 (N_7404,N_6724,N_6656);
and U7405 (N_7405,N_6993,N_6792);
and U7406 (N_7406,N_6912,N_6795);
and U7407 (N_7407,N_6559,N_6866);
xnor U7408 (N_7408,N_6697,N_6605);
and U7409 (N_7409,N_6723,N_6555);
nand U7410 (N_7410,N_6745,N_6736);
xnor U7411 (N_7411,N_6773,N_6794);
xnor U7412 (N_7412,N_6920,N_6728);
nand U7413 (N_7413,N_6782,N_6609);
or U7414 (N_7414,N_6758,N_6959);
xnor U7415 (N_7415,N_6681,N_6819);
xnor U7416 (N_7416,N_6547,N_6579);
nor U7417 (N_7417,N_6505,N_6762);
nand U7418 (N_7418,N_6598,N_6626);
nand U7419 (N_7419,N_6561,N_6902);
and U7420 (N_7420,N_6948,N_6600);
nand U7421 (N_7421,N_6836,N_6589);
or U7422 (N_7422,N_6606,N_6738);
and U7423 (N_7423,N_6554,N_6984);
or U7424 (N_7424,N_6898,N_6673);
xor U7425 (N_7425,N_6969,N_6959);
or U7426 (N_7426,N_6852,N_6586);
or U7427 (N_7427,N_6955,N_6606);
and U7428 (N_7428,N_6678,N_6870);
and U7429 (N_7429,N_6647,N_6559);
xnor U7430 (N_7430,N_6533,N_6580);
nor U7431 (N_7431,N_6522,N_6798);
and U7432 (N_7432,N_6928,N_6854);
nand U7433 (N_7433,N_6996,N_6751);
and U7434 (N_7434,N_6737,N_6851);
nand U7435 (N_7435,N_6656,N_6837);
and U7436 (N_7436,N_6770,N_6881);
and U7437 (N_7437,N_6808,N_6977);
and U7438 (N_7438,N_6621,N_6883);
nand U7439 (N_7439,N_6712,N_6602);
xnor U7440 (N_7440,N_6518,N_6516);
nand U7441 (N_7441,N_6892,N_6815);
nand U7442 (N_7442,N_6618,N_6689);
and U7443 (N_7443,N_6808,N_6740);
nor U7444 (N_7444,N_6832,N_6813);
nor U7445 (N_7445,N_6795,N_6823);
and U7446 (N_7446,N_6613,N_6542);
nand U7447 (N_7447,N_6513,N_6592);
and U7448 (N_7448,N_6502,N_6857);
xnor U7449 (N_7449,N_6962,N_6731);
xor U7450 (N_7450,N_6834,N_6572);
nand U7451 (N_7451,N_6922,N_6948);
nor U7452 (N_7452,N_6560,N_6524);
xnor U7453 (N_7453,N_6883,N_6513);
or U7454 (N_7454,N_6865,N_6750);
xnor U7455 (N_7455,N_6747,N_6968);
or U7456 (N_7456,N_6996,N_6827);
or U7457 (N_7457,N_6936,N_6534);
or U7458 (N_7458,N_6683,N_6944);
nor U7459 (N_7459,N_6795,N_6683);
and U7460 (N_7460,N_6593,N_6833);
nand U7461 (N_7461,N_6613,N_6854);
or U7462 (N_7462,N_6938,N_6568);
xnor U7463 (N_7463,N_6926,N_6651);
or U7464 (N_7464,N_6822,N_6543);
or U7465 (N_7465,N_6586,N_6530);
nand U7466 (N_7466,N_6584,N_6948);
nor U7467 (N_7467,N_6543,N_6980);
and U7468 (N_7468,N_6654,N_6886);
nand U7469 (N_7469,N_6749,N_6760);
xnor U7470 (N_7470,N_6556,N_6822);
or U7471 (N_7471,N_6901,N_6679);
or U7472 (N_7472,N_6570,N_6665);
nor U7473 (N_7473,N_6718,N_6923);
nor U7474 (N_7474,N_6729,N_6870);
or U7475 (N_7475,N_6691,N_6999);
nor U7476 (N_7476,N_6531,N_6629);
or U7477 (N_7477,N_6927,N_6638);
nor U7478 (N_7478,N_6817,N_6707);
and U7479 (N_7479,N_6720,N_6826);
xor U7480 (N_7480,N_6662,N_6813);
and U7481 (N_7481,N_6650,N_6583);
nor U7482 (N_7482,N_6727,N_6973);
and U7483 (N_7483,N_6615,N_6856);
xor U7484 (N_7484,N_6701,N_6904);
nand U7485 (N_7485,N_6919,N_6956);
or U7486 (N_7486,N_6821,N_6883);
or U7487 (N_7487,N_6623,N_6860);
or U7488 (N_7488,N_6942,N_6728);
nor U7489 (N_7489,N_6505,N_6672);
or U7490 (N_7490,N_6634,N_6615);
nor U7491 (N_7491,N_6631,N_6725);
and U7492 (N_7492,N_6917,N_6768);
and U7493 (N_7493,N_6615,N_6793);
and U7494 (N_7494,N_6672,N_6628);
and U7495 (N_7495,N_6674,N_6892);
or U7496 (N_7496,N_6719,N_6725);
nand U7497 (N_7497,N_6762,N_6572);
or U7498 (N_7498,N_6554,N_6916);
nor U7499 (N_7499,N_6628,N_6605);
and U7500 (N_7500,N_7062,N_7268);
nor U7501 (N_7501,N_7419,N_7327);
nor U7502 (N_7502,N_7270,N_7398);
nand U7503 (N_7503,N_7138,N_7330);
or U7504 (N_7504,N_7305,N_7130);
or U7505 (N_7505,N_7284,N_7261);
or U7506 (N_7506,N_7162,N_7407);
nand U7507 (N_7507,N_7424,N_7223);
nand U7508 (N_7508,N_7390,N_7037);
xor U7509 (N_7509,N_7412,N_7059);
nor U7510 (N_7510,N_7166,N_7324);
or U7511 (N_7511,N_7131,N_7251);
xor U7512 (N_7512,N_7238,N_7426);
nor U7513 (N_7513,N_7181,N_7161);
nor U7514 (N_7514,N_7151,N_7114);
or U7515 (N_7515,N_7370,N_7143);
xnor U7516 (N_7516,N_7376,N_7217);
xor U7517 (N_7517,N_7319,N_7322);
nand U7518 (N_7518,N_7420,N_7447);
and U7519 (N_7519,N_7311,N_7208);
nand U7520 (N_7520,N_7448,N_7417);
and U7521 (N_7521,N_7460,N_7459);
and U7522 (N_7522,N_7084,N_7304);
or U7523 (N_7523,N_7487,N_7226);
xnor U7524 (N_7524,N_7446,N_7197);
or U7525 (N_7525,N_7016,N_7331);
or U7526 (N_7526,N_7203,N_7329);
nor U7527 (N_7527,N_7190,N_7338);
xor U7528 (N_7528,N_7485,N_7436);
or U7529 (N_7529,N_7336,N_7025);
nand U7530 (N_7530,N_7088,N_7442);
nor U7531 (N_7531,N_7320,N_7204);
or U7532 (N_7532,N_7389,N_7321);
or U7533 (N_7533,N_7076,N_7458);
nand U7534 (N_7534,N_7317,N_7428);
nor U7535 (N_7535,N_7402,N_7074);
nor U7536 (N_7536,N_7364,N_7072);
and U7537 (N_7537,N_7044,N_7054);
nand U7538 (N_7538,N_7355,N_7174);
nand U7539 (N_7539,N_7163,N_7094);
or U7540 (N_7540,N_7422,N_7388);
and U7541 (N_7541,N_7228,N_7403);
and U7542 (N_7542,N_7303,N_7385);
xor U7543 (N_7543,N_7150,N_7133);
nand U7544 (N_7544,N_7154,N_7050);
nor U7545 (N_7545,N_7078,N_7418);
and U7546 (N_7546,N_7058,N_7280);
or U7547 (N_7547,N_7325,N_7276);
nand U7548 (N_7548,N_7348,N_7469);
and U7549 (N_7549,N_7002,N_7010);
or U7550 (N_7550,N_7244,N_7356);
or U7551 (N_7551,N_7134,N_7269);
and U7552 (N_7552,N_7405,N_7452);
nand U7553 (N_7553,N_7290,N_7494);
xor U7554 (N_7554,N_7187,N_7308);
nor U7555 (N_7555,N_7107,N_7421);
or U7556 (N_7556,N_7252,N_7039);
and U7557 (N_7557,N_7431,N_7211);
or U7558 (N_7558,N_7333,N_7450);
and U7559 (N_7559,N_7394,N_7091);
or U7560 (N_7560,N_7430,N_7082);
or U7561 (N_7561,N_7079,N_7256);
xnor U7562 (N_7562,N_7409,N_7281);
nor U7563 (N_7563,N_7068,N_7127);
or U7564 (N_7564,N_7188,N_7158);
nor U7565 (N_7565,N_7298,N_7299);
nor U7566 (N_7566,N_7227,N_7310);
nor U7567 (N_7567,N_7083,N_7024);
xnor U7568 (N_7568,N_7247,N_7465);
xnor U7569 (N_7569,N_7140,N_7396);
and U7570 (N_7570,N_7195,N_7155);
nor U7571 (N_7571,N_7198,N_7001);
nand U7572 (N_7572,N_7199,N_7027);
nor U7573 (N_7573,N_7093,N_7326);
or U7574 (N_7574,N_7175,N_7361);
nand U7575 (N_7575,N_7480,N_7033);
xnor U7576 (N_7576,N_7391,N_7395);
and U7577 (N_7577,N_7171,N_7357);
nand U7578 (N_7578,N_7236,N_7495);
xor U7579 (N_7579,N_7372,N_7386);
or U7580 (N_7580,N_7359,N_7497);
xnor U7581 (N_7581,N_7449,N_7382);
and U7582 (N_7582,N_7440,N_7400);
or U7583 (N_7583,N_7439,N_7486);
and U7584 (N_7584,N_7354,N_7482);
and U7585 (N_7585,N_7471,N_7029);
or U7586 (N_7586,N_7491,N_7429);
or U7587 (N_7587,N_7119,N_7052);
or U7588 (N_7588,N_7490,N_7425);
or U7589 (N_7589,N_7224,N_7081);
or U7590 (N_7590,N_7410,N_7337);
nor U7591 (N_7591,N_7206,N_7036);
nor U7592 (N_7592,N_7470,N_7484);
nor U7593 (N_7593,N_7231,N_7103);
xnor U7594 (N_7594,N_7344,N_7248);
nor U7595 (N_7595,N_7352,N_7101);
xnor U7596 (N_7596,N_7069,N_7275);
or U7597 (N_7597,N_7136,N_7132);
nand U7598 (N_7598,N_7080,N_7179);
and U7599 (N_7599,N_7443,N_7472);
or U7600 (N_7600,N_7277,N_7205);
and U7601 (N_7601,N_7215,N_7477);
nor U7602 (N_7602,N_7295,N_7263);
xor U7603 (N_7603,N_7349,N_7200);
xnor U7604 (N_7604,N_7373,N_7479);
nor U7605 (N_7605,N_7099,N_7129);
or U7606 (N_7606,N_7413,N_7454);
or U7607 (N_7607,N_7250,N_7111);
or U7608 (N_7608,N_7225,N_7157);
nor U7609 (N_7609,N_7196,N_7384);
xor U7610 (N_7610,N_7245,N_7498);
nand U7611 (N_7611,N_7427,N_7021);
nor U7612 (N_7612,N_7255,N_7375);
and U7613 (N_7613,N_7009,N_7499);
or U7614 (N_7614,N_7264,N_7230);
nor U7615 (N_7615,N_7467,N_7489);
nand U7616 (N_7616,N_7014,N_7049);
and U7617 (N_7617,N_7401,N_7180);
xor U7618 (N_7618,N_7393,N_7260);
nand U7619 (N_7619,N_7381,N_7067);
xor U7620 (N_7620,N_7003,N_7377);
xor U7621 (N_7621,N_7464,N_7258);
xor U7622 (N_7622,N_7035,N_7241);
xor U7623 (N_7623,N_7306,N_7463);
or U7624 (N_7624,N_7026,N_7153);
nand U7625 (N_7625,N_7368,N_7095);
nand U7626 (N_7626,N_7071,N_7374);
xnor U7627 (N_7627,N_7432,N_7408);
or U7628 (N_7628,N_7307,N_7481);
nand U7629 (N_7629,N_7271,N_7122);
or U7630 (N_7630,N_7218,N_7367);
nand U7631 (N_7631,N_7488,N_7334);
nand U7632 (N_7632,N_7239,N_7047);
nand U7633 (N_7633,N_7221,N_7137);
and U7634 (N_7634,N_7005,N_7340);
xnor U7635 (N_7635,N_7173,N_7492);
and U7636 (N_7636,N_7202,N_7476);
or U7637 (N_7637,N_7462,N_7312);
xnor U7638 (N_7638,N_7193,N_7148);
xnor U7639 (N_7639,N_7272,N_7189);
or U7640 (N_7640,N_7214,N_7046);
or U7641 (N_7641,N_7040,N_7229);
xor U7642 (N_7642,N_7353,N_7493);
xnor U7643 (N_7643,N_7108,N_7316);
nor U7644 (N_7644,N_7273,N_7350);
xor U7645 (N_7645,N_7145,N_7249);
xor U7646 (N_7646,N_7456,N_7118);
xnor U7647 (N_7647,N_7423,N_7192);
xnor U7648 (N_7648,N_7028,N_7110);
nor U7649 (N_7649,N_7351,N_7013);
or U7650 (N_7650,N_7346,N_7406);
or U7651 (N_7651,N_7152,N_7387);
nand U7652 (N_7652,N_7115,N_7219);
nand U7653 (N_7653,N_7017,N_7339);
xor U7654 (N_7654,N_7043,N_7383);
or U7655 (N_7655,N_7222,N_7070);
or U7656 (N_7656,N_7116,N_7100);
xor U7657 (N_7657,N_7233,N_7345);
nor U7658 (N_7658,N_7300,N_7369);
or U7659 (N_7659,N_7042,N_7288);
and U7660 (N_7660,N_7360,N_7160);
xnor U7661 (N_7661,N_7109,N_7254);
xnor U7662 (N_7662,N_7146,N_7444);
or U7663 (N_7663,N_7022,N_7023);
xnor U7664 (N_7664,N_7285,N_7283);
nor U7665 (N_7665,N_7414,N_7121);
nor U7666 (N_7666,N_7191,N_7365);
nor U7667 (N_7667,N_7301,N_7262);
nand U7668 (N_7668,N_7057,N_7434);
nor U7669 (N_7669,N_7404,N_7282);
xor U7670 (N_7670,N_7451,N_7274);
and U7671 (N_7671,N_7096,N_7073);
nand U7672 (N_7672,N_7182,N_7184);
nor U7673 (N_7673,N_7041,N_7060);
xor U7674 (N_7674,N_7293,N_7253);
xnor U7675 (N_7675,N_7183,N_7149);
or U7676 (N_7676,N_7085,N_7455);
nand U7677 (N_7677,N_7030,N_7265);
and U7678 (N_7678,N_7415,N_7397);
nand U7679 (N_7679,N_7125,N_7380);
xnor U7680 (N_7680,N_7259,N_7411);
and U7681 (N_7681,N_7104,N_7102);
xor U7682 (N_7682,N_7437,N_7232);
xor U7683 (N_7683,N_7475,N_7315);
and U7684 (N_7684,N_7185,N_7332);
xnor U7685 (N_7685,N_7159,N_7178);
or U7686 (N_7686,N_7341,N_7213);
nor U7687 (N_7687,N_7065,N_7453);
and U7688 (N_7688,N_7018,N_7468);
xnor U7689 (N_7689,N_7092,N_7063);
xnor U7690 (N_7690,N_7242,N_7064);
nand U7691 (N_7691,N_7212,N_7055);
and U7692 (N_7692,N_7045,N_7004);
xor U7693 (N_7693,N_7313,N_7194);
and U7694 (N_7694,N_7363,N_7291);
nand U7695 (N_7695,N_7172,N_7209);
nor U7696 (N_7696,N_7012,N_7144);
and U7697 (N_7697,N_7240,N_7379);
or U7698 (N_7698,N_7289,N_7266);
and U7699 (N_7699,N_7032,N_7234);
or U7700 (N_7700,N_7164,N_7117);
nor U7701 (N_7701,N_7441,N_7020);
and U7702 (N_7702,N_7135,N_7483);
nand U7703 (N_7703,N_7019,N_7314);
nand U7704 (N_7704,N_7170,N_7106);
xor U7705 (N_7705,N_7257,N_7343);
or U7706 (N_7706,N_7015,N_7433);
or U7707 (N_7707,N_7077,N_7473);
nor U7708 (N_7708,N_7445,N_7392);
and U7709 (N_7709,N_7147,N_7287);
nand U7710 (N_7710,N_7156,N_7278);
nor U7711 (N_7711,N_7169,N_7098);
or U7712 (N_7712,N_7123,N_7097);
nand U7713 (N_7713,N_7165,N_7366);
or U7714 (N_7714,N_7362,N_7478);
xor U7715 (N_7715,N_7466,N_7168);
and U7716 (N_7716,N_7008,N_7011);
xnor U7717 (N_7717,N_7006,N_7038);
nor U7718 (N_7718,N_7237,N_7302);
xnor U7719 (N_7719,N_7113,N_7051);
or U7720 (N_7720,N_7496,N_7139);
and U7721 (N_7721,N_7089,N_7112);
or U7722 (N_7722,N_7086,N_7090);
or U7723 (N_7723,N_7358,N_7297);
and U7724 (N_7724,N_7034,N_7318);
nor U7725 (N_7725,N_7292,N_7056);
nand U7726 (N_7726,N_7461,N_7416);
or U7727 (N_7727,N_7371,N_7120);
or U7728 (N_7728,N_7347,N_7066);
nor U7729 (N_7729,N_7141,N_7128);
xor U7730 (N_7730,N_7210,N_7186);
and U7731 (N_7731,N_7061,N_7267);
xor U7732 (N_7732,N_7105,N_7294);
nand U7733 (N_7733,N_7309,N_7235);
nand U7734 (N_7734,N_7126,N_7279);
and U7735 (N_7735,N_7007,N_7207);
nor U7736 (N_7736,N_7438,N_7167);
and U7737 (N_7737,N_7177,N_7031);
nor U7738 (N_7738,N_7323,N_7474);
nand U7739 (N_7739,N_7243,N_7328);
nand U7740 (N_7740,N_7457,N_7435);
or U7741 (N_7741,N_7000,N_7075);
nand U7742 (N_7742,N_7087,N_7335);
nand U7743 (N_7743,N_7378,N_7053);
xnor U7744 (N_7744,N_7286,N_7176);
nand U7745 (N_7745,N_7124,N_7246);
and U7746 (N_7746,N_7399,N_7296);
nor U7747 (N_7747,N_7342,N_7220);
nand U7748 (N_7748,N_7142,N_7216);
nor U7749 (N_7749,N_7201,N_7048);
xor U7750 (N_7750,N_7364,N_7441);
and U7751 (N_7751,N_7479,N_7233);
nor U7752 (N_7752,N_7310,N_7105);
nor U7753 (N_7753,N_7335,N_7325);
and U7754 (N_7754,N_7316,N_7053);
or U7755 (N_7755,N_7220,N_7308);
and U7756 (N_7756,N_7193,N_7299);
xor U7757 (N_7757,N_7026,N_7307);
xor U7758 (N_7758,N_7001,N_7251);
nor U7759 (N_7759,N_7402,N_7053);
nand U7760 (N_7760,N_7054,N_7459);
or U7761 (N_7761,N_7138,N_7085);
or U7762 (N_7762,N_7391,N_7013);
xnor U7763 (N_7763,N_7093,N_7142);
xor U7764 (N_7764,N_7305,N_7293);
xor U7765 (N_7765,N_7209,N_7458);
nor U7766 (N_7766,N_7198,N_7299);
or U7767 (N_7767,N_7277,N_7004);
xnor U7768 (N_7768,N_7203,N_7463);
nand U7769 (N_7769,N_7022,N_7046);
xor U7770 (N_7770,N_7461,N_7045);
nor U7771 (N_7771,N_7396,N_7442);
or U7772 (N_7772,N_7166,N_7279);
nor U7773 (N_7773,N_7176,N_7141);
and U7774 (N_7774,N_7376,N_7466);
xnor U7775 (N_7775,N_7039,N_7185);
nor U7776 (N_7776,N_7047,N_7111);
or U7777 (N_7777,N_7406,N_7132);
or U7778 (N_7778,N_7406,N_7207);
xor U7779 (N_7779,N_7086,N_7295);
nor U7780 (N_7780,N_7349,N_7256);
nand U7781 (N_7781,N_7358,N_7493);
and U7782 (N_7782,N_7187,N_7311);
or U7783 (N_7783,N_7469,N_7386);
or U7784 (N_7784,N_7066,N_7467);
nor U7785 (N_7785,N_7248,N_7295);
and U7786 (N_7786,N_7193,N_7293);
nand U7787 (N_7787,N_7193,N_7354);
or U7788 (N_7788,N_7317,N_7178);
nor U7789 (N_7789,N_7486,N_7070);
or U7790 (N_7790,N_7347,N_7174);
xnor U7791 (N_7791,N_7204,N_7132);
nand U7792 (N_7792,N_7403,N_7020);
xor U7793 (N_7793,N_7209,N_7309);
nor U7794 (N_7794,N_7028,N_7355);
nand U7795 (N_7795,N_7109,N_7013);
xor U7796 (N_7796,N_7026,N_7167);
nand U7797 (N_7797,N_7139,N_7467);
and U7798 (N_7798,N_7424,N_7237);
and U7799 (N_7799,N_7175,N_7484);
xnor U7800 (N_7800,N_7403,N_7241);
nand U7801 (N_7801,N_7433,N_7103);
and U7802 (N_7802,N_7259,N_7261);
nor U7803 (N_7803,N_7002,N_7037);
xor U7804 (N_7804,N_7285,N_7499);
or U7805 (N_7805,N_7210,N_7071);
and U7806 (N_7806,N_7449,N_7026);
and U7807 (N_7807,N_7191,N_7348);
xnor U7808 (N_7808,N_7040,N_7450);
and U7809 (N_7809,N_7150,N_7483);
nor U7810 (N_7810,N_7410,N_7200);
and U7811 (N_7811,N_7142,N_7184);
nor U7812 (N_7812,N_7410,N_7352);
nand U7813 (N_7813,N_7245,N_7008);
nand U7814 (N_7814,N_7280,N_7154);
nor U7815 (N_7815,N_7479,N_7133);
or U7816 (N_7816,N_7446,N_7416);
nand U7817 (N_7817,N_7272,N_7438);
xor U7818 (N_7818,N_7388,N_7338);
nor U7819 (N_7819,N_7274,N_7330);
and U7820 (N_7820,N_7129,N_7387);
and U7821 (N_7821,N_7321,N_7377);
xor U7822 (N_7822,N_7179,N_7128);
nand U7823 (N_7823,N_7276,N_7250);
nand U7824 (N_7824,N_7203,N_7187);
and U7825 (N_7825,N_7018,N_7090);
xor U7826 (N_7826,N_7017,N_7110);
nor U7827 (N_7827,N_7286,N_7499);
and U7828 (N_7828,N_7015,N_7310);
nand U7829 (N_7829,N_7194,N_7425);
and U7830 (N_7830,N_7128,N_7011);
nand U7831 (N_7831,N_7083,N_7417);
nor U7832 (N_7832,N_7274,N_7069);
xor U7833 (N_7833,N_7145,N_7223);
and U7834 (N_7834,N_7498,N_7370);
xnor U7835 (N_7835,N_7328,N_7015);
xor U7836 (N_7836,N_7270,N_7359);
or U7837 (N_7837,N_7448,N_7278);
xnor U7838 (N_7838,N_7290,N_7450);
xnor U7839 (N_7839,N_7203,N_7003);
nand U7840 (N_7840,N_7175,N_7112);
nand U7841 (N_7841,N_7470,N_7373);
xor U7842 (N_7842,N_7249,N_7262);
nand U7843 (N_7843,N_7252,N_7075);
and U7844 (N_7844,N_7280,N_7372);
and U7845 (N_7845,N_7364,N_7134);
or U7846 (N_7846,N_7312,N_7191);
nand U7847 (N_7847,N_7055,N_7138);
and U7848 (N_7848,N_7261,N_7426);
and U7849 (N_7849,N_7239,N_7018);
or U7850 (N_7850,N_7245,N_7356);
xor U7851 (N_7851,N_7161,N_7294);
and U7852 (N_7852,N_7429,N_7438);
and U7853 (N_7853,N_7141,N_7368);
and U7854 (N_7854,N_7286,N_7366);
xnor U7855 (N_7855,N_7002,N_7213);
nor U7856 (N_7856,N_7094,N_7157);
and U7857 (N_7857,N_7244,N_7256);
and U7858 (N_7858,N_7488,N_7087);
nor U7859 (N_7859,N_7292,N_7034);
and U7860 (N_7860,N_7216,N_7004);
and U7861 (N_7861,N_7147,N_7386);
and U7862 (N_7862,N_7455,N_7462);
xor U7863 (N_7863,N_7190,N_7323);
xor U7864 (N_7864,N_7340,N_7157);
or U7865 (N_7865,N_7324,N_7355);
and U7866 (N_7866,N_7051,N_7447);
nor U7867 (N_7867,N_7091,N_7069);
and U7868 (N_7868,N_7291,N_7184);
nor U7869 (N_7869,N_7084,N_7485);
and U7870 (N_7870,N_7134,N_7236);
nor U7871 (N_7871,N_7302,N_7029);
nor U7872 (N_7872,N_7451,N_7067);
or U7873 (N_7873,N_7015,N_7008);
or U7874 (N_7874,N_7237,N_7028);
xnor U7875 (N_7875,N_7104,N_7179);
xor U7876 (N_7876,N_7263,N_7390);
or U7877 (N_7877,N_7359,N_7268);
or U7878 (N_7878,N_7343,N_7306);
and U7879 (N_7879,N_7428,N_7382);
nand U7880 (N_7880,N_7201,N_7347);
nand U7881 (N_7881,N_7431,N_7461);
and U7882 (N_7882,N_7071,N_7305);
or U7883 (N_7883,N_7160,N_7433);
and U7884 (N_7884,N_7352,N_7349);
nor U7885 (N_7885,N_7485,N_7040);
xor U7886 (N_7886,N_7394,N_7300);
and U7887 (N_7887,N_7269,N_7308);
and U7888 (N_7888,N_7176,N_7104);
nand U7889 (N_7889,N_7427,N_7269);
xor U7890 (N_7890,N_7095,N_7350);
xor U7891 (N_7891,N_7272,N_7079);
nand U7892 (N_7892,N_7265,N_7365);
xnor U7893 (N_7893,N_7288,N_7153);
nor U7894 (N_7894,N_7442,N_7195);
nand U7895 (N_7895,N_7404,N_7129);
or U7896 (N_7896,N_7025,N_7015);
nand U7897 (N_7897,N_7130,N_7072);
nor U7898 (N_7898,N_7236,N_7315);
nand U7899 (N_7899,N_7036,N_7100);
nor U7900 (N_7900,N_7244,N_7400);
or U7901 (N_7901,N_7258,N_7280);
and U7902 (N_7902,N_7396,N_7035);
nor U7903 (N_7903,N_7281,N_7406);
and U7904 (N_7904,N_7360,N_7455);
nand U7905 (N_7905,N_7474,N_7290);
nand U7906 (N_7906,N_7235,N_7411);
nor U7907 (N_7907,N_7232,N_7467);
nand U7908 (N_7908,N_7047,N_7052);
or U7909 (N_7909,N_7343,N_7483);
nand U7910 (N_7910,N_7339,N_7096);
xnor U7911 (N_7911,N_7418,N_7138);
nand U7912 (N_7912,N_7439,N_7276);
xor U7913 (N_7913,N_7428,N_7348);
xnor U7914 (N_7914,N_7243,N_7245);
xnor U7915 (N_7915,N_7000,N_7093);
nand U7916 (N_7916,N_7301,N_7192);
and U7917 (N_7917,N_7144,N_7180);
or U7918 (N_7918,N_7163,N_7178);
nor U7919 (N_7919,N_7245,N_7329);
nor U7920 (N_7920,N_7268,N_7199);
or U7921 (N_7921,N_7388,N_7170);
nand U7922 (N_7922,N_7368,N_7250);
and U7923 (N_7923,N_7165,N_7013);
and U7924 (N_7924,N_7268,N_7060);
xor U7925 (N_7925,N_7469,N_7358);
nand U7926 (N_7926,N_7255,N_7448);
xor U7927 (N_7927,N_7096,N_7199);
nand U7928 (N_7928,N_7441,N_7393);
or U7929 (N_7929,N_7109,N_7483);
or U7930 (N_7930,N_7145,N_7422);
nor U7931 (N_7931,N_7463,N_7168);
xor U7932 (N_7932,N_7249,N_7097);
nand U7933 (N_7933,N_7414,N_7191);
nand U7934 (N_7934,N_7378,N_7466);
or U7935 (N_7935,N_7108,N_7276);
and U7936 (N_7936,N_7055,N_7366);
and U7937 (N_7937,N_7070,N_7016);
nor U7938 (N_7938,N_7363,N_7472);
xor U7939 (N_7939,N_7210,N_7043);
and U7940 (N_7940,N_7003,N_7246);
or U7941 (N_7941,N_7234,N_7497);
nor U7942 (N_7942,N_7496,N_7113);
nor U7943 (N_7943,N_7063,N_7145);
xnor U7944 (N_7944,N_7238,N_7089);
nor U7945 (N_7945,N_7186,N_7343);
nand U7946 (N_7946,N_7174,N_7176);
xnor U7947 (N_7947,N_7223,N_7479);
nor U7948 (N_7948,N_7351,N_7192);
or U7949 (N_7949,N_7109,N_7294);
and U7950 (N_7950,N_7055,N_7259);
or U7951 (N_7951,N_7248,N_7491);
nor U7952 (N_7952,N_7372,N_7325);
nor U7953 (N_7953,N_7190,N_7493);
or U7954 (N_7954,N_7120,N_7318);
nand U7955 (N_7955,N_7378,N_7380);
and U7956 (N_7956,N_7222,N_7284);
nand U7957 (N_7957,N_7232,N_7203);
nand U7958 (N_7958,N_7053,N_7056);
nor U7959 (N_7959,N_7361,N_7125);
xnor U7960 (N_7960,N_7152,N_7364);
nor U7961 (N_7961,N_7037,N_7261);
and U7962 (N_7962,N_7270,N_7361);
or U7963 (N_7963,N_7104,N_7395);
and U7964 (N_7964,N_7440,N_7465);
or U7965 (N_7965,N_7294,N_7464);
nand U7966 (N_7966,N_7181,N_7152);
nor U7967 (N_7967,N_7378,N_7476);
nor U7968 (N_7968,N_7275,N_7381);
xor U7969 (N_7969,N_7015,N_7039);
xnor U7970 (N_7970,N_7223,N_7155);
or U7971 (N_7971,N_7005,N_7214);
nand U7972 (N_7972,N_7243,N_7236);
and U7973 (N_7973,N_7064,N_7215);
and U7974 (N_7974,N_7124,N_7035);
xnor U7975 (N_7975,N_7325,N_7316);
or U7976 (N_7976,N_7447,N_7432);
xor U7977 (N_7977,N_7049,N_7001);
nand U7978 (N_7978,N_7205,N_7157);
or U7979 (N_7979,N_7230,N_7237);
and U7980 (N_7980,N_7422,N_7444);
nor U7981 (N_7981,N_7455,N_7159);
and U7982 (N_7982,N_7140,N_7008);
nand U7983 (N_7983,N_7255,N_7385);
nor U7984 (N_7984,N_7263,N_7042);
or U7985 (N_7985,N_7417,N_7447);
nor U7986 (N_7986,N_7008,N_7262);
or U7987 (N_7987,N_7136,N_7467);
or U7988 (N_7988,N_7277,N_7439);
nor U7989 (N_7989,N_7392,N_7277);
nor U7990 (N_7990,N_7481,N_7190);
nor U7991 (N_7991,N_7144,N_7354);
xor U7992 (N_7992,N_7037,N_7204);
xnor U7993 (N_7993,N_7436,N_7451);
nand U7994 (N_7994,N_7400,N_7092);
and U7995 (N_7995,N_7116,N_7160);
and U7996 (N_7996,N_7285,N_7074);
nand U7997 (N_7997,N_7206,N_7004);
or U7998 (N_7998,N_7478,N_7100);
or U7999 (N_7999,N_7162,N_7096);
nand U8000 (N_8000,N_7914,N_7830);
nor U8001 (N_8001,N_7802,N_7674);
or U8002 (N_8002,N_7908,N_7934);
and U8003 (N_8003,N_7625,N_7671);
nor U8004 (N_8004,N_7616,N_7745);
xnor U8005 (N_8005,N_7893,N_7649);
nor U8006 (N_8006,N_7971,N_7856);
or U8007 (N_8007,N_7621,N_7896);
nor U8008 (N_8008,N_7955,N_7540);
xnor U8009 (N_8009,N_7619,N_7897);
nand U8010 (N_8010,N_7578,N_7819);
xor U8011 (N_8011,N_7562,N_7710);
and U8012 (N_8012,N_7620,N_7698);
nor U8013 (N_8013,N_7851,N_7536);
xnor U8014 (N_8014,N_7724,N_7505);
and U8015 (N_8015,N_7930,N_7550);
and U8016 (N_8016,N_7529,N_7503);
xor U8017 (N_8017,N_7785,N_7885);
or U8018 (N_8018,N_7855,N_7778);
xor U8019 (N_8019,N_7939,N_7718);
and U8020 (N_8020,N_7521,N_7976);
or U8021 (N_8021,N_7796,N_7563);
or U8022 (N_8022,N_7973,N_7808);
xnor U8023 (N_8023,N_7868,N_7803);
xnor U8024 (N_8024,N_7655,N_7932);
or U8025 (N_8025,N_7834,N_7782);
nor U8026 (N_8026,N_7570,N_7623);
nand U8027 (N_8027,N_7644,N_7588);
or U8028 (N_8028,N_7879,N_7717);
xor U8029 (N_8029,N_7573,N_7515);
or U8030 (N_8030,N_7615,N_7725);
or U8031 (N_8031,N_7987,N_7682);
xnor U8032 (N_8032,N_7813,N_7557);
and U8033 (N_8033,N_7635,N_7843);
xor U8034 (N_8034,N_7773,N_7846);
xnor U8035 (N_8035,N_7920,N_7837);
or U8036 (N_8036,N_7787,N_7989);
and U8037 (N_8037,N_7596,N_7753);
and U8038 (N_8038,N_7607,N_7978);
or U8039 (N_8039,N_7730,N_7881);
and U8040 (N_8040,N_7913,N_7757);
nor U8041 (N_8041,N_7888,N_7963);
nor U8042 (N_8042,N_7775,N_7765);
or U8043 (N_8043,N_7795,N_7760);
and U8044 (N_8044,N_7558,N_7501);
nor U8045 (N_8045,N_7952,N_7605);
xnor U8046 (N_8046,N_7680,N_7736);
nand U8047 (N_8047,N_7774,N_7887);
xor U8048 (N_8048,N_7611,N_7579);
xor U8049 (N_8049,N_7610,N_7903);
and U8050 (N_8050,N_7632,N_7829);
nor U8051 (N_8051,N_7666,N_7513);
nand U8052 (N_8052,N_7875,N_7945);
or U8053 (N_8053,N_7759,N_7617);
or U8054 (N_8054,N_7580,N_7953);
xnor U8055 (N_8055,N_7998,N_7788);
nand U8056 (N_8056,N_7962,N_7764);
nand U8057 (N_8057,N_7543,N_7949);
and U8058 (N_8058,N_7918,N_7958);
nand U8059 (N_8059,N_7713,N_7756);
or U8060 (N_8060,N_7721,N_7938);
or U8061 (N_8061,N_7701,N_7749);
xnor U8062 (N_8062,N_7544,N_7656);
nand U8063 (N_8063,N_7648,N_7694);
nand U8064 (N_8064,N_7676,N_7806);
nor U8065 (N_8065,N_7733,N_7612);
nor U8066 (N_8066,N_7595,N_7613);
nand U8067 (N_8067,N_7792,N_7811);
nand U8068 (N_8068,N_7568,N_7519);
xnor U8069 (N_8069,N_7793,N_7684);
and U8070 (N_8070,N_7997,N_7709);
xnor U8071 (N_8071,N_7891,N_7643);
nand U8072 (N_8072,N_7520,N_7950);
nand U8073 (N_8073,N_7751,N_7933);
xnor U8074 (N_8074,N_7640,N_7618);
nand U8075 (N_8075,N_7712,N_7797);
xnor U8076 (N_8076,N_7816,N_7946);
nor U8077 (N_8077,N_7772,N_7586);
xor U8078 (N_8078,N_7831,N_7700);
xnor U8079 (N_8079,N_7815,N_7780);
and U8080 (N_8080,N_7679,N_7912);
or U8081 (N_8081,N_7894,N_7907);
xor U8082 (N_8082,N_7556,N_7683);
nor U8083 (N_8083,N_7650,N_7661);
nor U8084 (N_8084,N_7669,N_7744);
nor U8085 (N_8085,N_7516,N_7690);
or U8086 (N_8086,N_7850,N_7585);
xor U8087 (N_8087,N_7645,N_7711);
or U8088 (N_8088,N_7905,N_7541);
xor U8089 (N_8089,N_7719,N_7532);
nor U8090 (N_8090,N_7731,N_7738);
nor U8091 (N_8091,N_7758,N_7705);
or U8092 (N_8092,N_7628,N_7985);
nor U8093 (N_8093,N_7860,N_7728);
or U8094 (N_8094,N_7518,N_7972);
xnor U8095 (N_8095,N_7553,N_7627);
or U8096 (N_8096,N_7993,N_7964);
or U8097 (N_8097,N_7981,N_7691);
xnor U8098 (N_8098,N_7892,N_7979);
xor U8099 (N_8099,N_7569,N_7692);
and U8100 (N_8100,N_7583,N_7707);
and U8101 (N_8101,N_7658,N_7906);
and U8102 (N_8102,N_7768,N_7857);
or U8103 (N_8103,N_7869,N_7871);
xnor U8104 (N_8104,N_7880,N_7741);
or U8105 (N_8105,N_7921,N_7576);
and U8106 (N_8106,N_7821,N_7672);
xor U8107 (N_8107,N_7873,N_7827);
nand U8108 (N_8108,N_7965,N_7783);
nor U8109 (N_8109,N_7755,N_7902);
or U8110 (N_8110,N_7589,N_7561);
and U8111 (N_8111,N_7864,N_7752);
or U8112 (N_8112,N_7748,N_7609);
and U8113 (N_8113,N_7631,N_7695);
nand U8114 (N_8114,N_7983,N_7577);
xor U8115 (N_8115,N_7899,N_7500);
or U8116 (N_8116,N_7948,N_7943);
nor U8117 (N_8117,N_7599,N_7708);
or U8118 (N_8118,N_7844,N_7988);
and U8119 (N_8119,N_7940,N_7863);
and U8120 (N_8120,N_7776,N_7872);
nor U8121 (N_8121,N_7750,N_7735);
and U8122 (N_8122,N_7944,N_7828);
and U8123 (N_8123,N_7936,N_7626);
nand U8124 (N_8124,N_7678,N_7699);
or U8125 (N_8125,N_7931,N_7598);
nor U8126 (N_8126,N_7928,N_7657);
or U8127 (N_8127,N_7592,N_7524);
and U8128 (N_8128,N_7954,N_7651);
xor U8129 (N_8129,N_7746,N_7591);
and U8130 (N_8130,N_7762,N_7587);
xnor U8131 (N_8131,N_7791,N_7847);
and U8132 (N_8132,N_7854,N_7539);
xnor U8133 (N_8133,N_7994,N_7689);
xor U8134 (N_8134,N_7805,N_7876);
xnor U8135 (N_8135,N_7923,N_7777);
or U8136 (N_8136,N_7686,N_7729);
and U8137 (N_8137,N_7883,N_7537);
nor U8138 (N_8138,N_7801,N_7977);
nor U8139 (N_8139,N_7859,N_7804);
and U8140 (N_8140,N_7722,N_7502);
and U8141 (N_8141,N_7526,N_7527);
nor U8142 (N_8142,N_7685,N_7966);
nand U8143 (N_8143,N_7866,N_7525);
nand U8144 (N_8144,N_7779,N_7662);
and U8145 (N_8145,N_7687,N_7771);
nand U8146 (N_8146,N_7726,N_7970);
or U8147 (N_8147,N_7975,N_7867);
or U8148 (N_8148,N_7984,N_7799);
nor U8149 (N_8149,N_7849,N_7734);
and U8150 (N_8150,N_7999,N_7737);
or U8151 (N_8151,N_7603,N_7600);
or U8152 (N_8152,N_7665,N_7660);
nor U8153 (N_8153,N_7647,N_7574);
and U8154 (N_8154,N_7900,N_7911);
xnor U8155 (N_8155,N_7812,N_7715);
nand U8156 (N_8156,N_7927,N_7681);
nor U8157 (N_8157,N_7861,N_7582);
and U8158 (N_8158,N_7739,N_7531);
or U8159 (N_8159,N_7693,N_7677);
nand U8160 (N_8160,N_7642,N_7670);
or U8161 (N_8161,N_7514,N_7663);
nand U8162 (N_8162,N_7538,N_7798);
nand U8163 (N_8163,N_7697,N_7742);
nor U8164 (N_8164,N_7982,N_7546);
xnor U8165 (N_8165,N_7786,N_7552);
nand U8166 (N_8166,N_7852,N_7545);
or U8167 (N_8167,N_7767,N_7720);
nand U8168 (N_8168,N_7836,N_7942);
nand U8169 (N_8169,N_7884,N_7549);
or U8170 (N_8170,N_7548,N_7703);
and U8171 (N_8171,N_7925,N_7528);
and U8172 (N_8172,N_7941,N_7575);
nand U8173 (N_8173,N_7947,N_7602);
nor U8174 (N_8174,N_7924,N_7507);
and U8175 (N_8175,N_7901,N_7889);
or U8176 (N_8176,N_7886,N_7995);
nor U8177 (N_8177,N_7727,N_7959);
xor U8178 (N_8178,N_7781,N_7633);
nor U8179 (N_8179,N_7668,N_7820);
xor U8180 (N_8180,N_7790,N_7858);
or U8181 (N_8181,N_7910,N_7996);
and U8182 (N_8182,N_7814,N_7853);
and U8183 (N_8183,N_7968,N_7555);
and U8184 (N_8184,N_7838,N_7817);
and U8185 (N_8185,N_7564,N_7675);
and U8186 (N_8186,N_7874,N_7696);
nor U8187 (N_8187,N_7723,N_7634);
or U8188 (N_8188,N_7862,N_7732);
nor U8189 (N_8189,N_7878,N_7594);
or U8190 (N_8190,N_7980,N_7990);
or U8191 (N_8191,N_7926,N_7547);
and U8192 (N_8192,N_7530,N_7706);
or U8193 (N_8193,N_7770,N_7825);
and U8194 (N_8194,N_7898,N_7824);
or U8195 (N_8195,N_7716,N_7840);
or U8196 (N_8196,N_7614,N_7915);
and U8197 (N_8197,N_7559,N_7673);
or U8198 (N_8198,N_7638,N_7935);
or U8199 (N_8199,N_7848,N_7877);
xnor U8200 (N_8200,N_7807,N_7512);
nor U8201 (N_8201,N_7654,N_7653);
and U8202 (N_8202,N_7581,N_7509);
nor U8203 (N_8203,N_7630,N_7809);
nand U8204 (N_8204,N_7646,N_7641);
nor U8205 (N_8205,N_7754,N_7818);
xnor U8206 (N_8206,N_7560,N_7624);
nand U8207 (N_8207,N_7637,N_7761);
nand U8208 (N_8208,N_7833,N_7702);
xor U8209 (N_8209,N_7533,N_7704);
or U8210 (N_8210,N_7504,N_7510);
or U8211 (N_8211,N_7909,N_7937);
nand U8212 (N_8212,N_7551,N_7572);
nor U8213 (N_8213,N_7511,N_7922);
xnor U8214 (N_8214,N_7542,N_7593);
nor U8215 (N_8215,N_7919,N_7810);
xor U8216 (N_8216,N_7784,N_7590);
xnor U8217 (N_8217,N_7839,N_7688);
xor U8218 (N_8218,N_7534,N_7535);
or U8219 (N_8219,N_7800,N_7608);
xor U8220 (N_8220,N_7992,N_7565);
xnor U8221 (N_8221,N_7584,N_7636);
xor U8222 (N_8222,N_7622,N_7917);
nand U8223 (N_8223,N_7961,N_7740);
or U8224 (N_8224,N_7794,N_7841);
and U8225 (N_8225,N_7714,N_7974);
or U8226 (N_8226,N_7606,N_7951);
nor U8227 (N_8227,N_7826,N_7566);
xor U8228 (N_8228,N_7763,N_7967);
and U8229 (N_8229,N_7916,N_7554);
xor U8230 (N_8230,N_7597,N_7747);
and U8231 (N_8231,N_7822,N_7956);
nand U8232 (N_8232,N_7639,N_7604);
xnor U8233 (N_8233,N_7517,N_7960);
or U8234 (N_8234,N_7506,N_7659);
nor U8235 (N_8235,N_7743,N_7845);
or U8236 (N_8236,N_7991,N_7567);
nor U8237 (N_8237,N_7865,N_7769);
nand U8238 (N_8238,N_7823,N_7832);
or U8239 (N_8239,N_7890,N_7842);
xnor U8240 (N_8240,N_7957,N_7522);
and U8241 (N_8241,N_7667,N_7895);
nor U8242 (N_8242,N_7789,N_7508);
or U8243 (N_8243,N_7986,N_7766);
nor U8244 (N_8244,N_7904,N_7652);
nand U8245 (N_8245,N_7601,N_7870);
or U8246 (N_8246,N_7969,N_7629);
and U8247 (N_8247,N_7835,N_7929);
xor U8248 (N_8248,N_7523,N_7882);
or U8249 (N_8249,N_7571,N_7664);
nand U8250 (N_8250,N_7814,N_7686);
and U8251 (N_8251,N_7529,N_7763);
and U8252 (N_8252,N_7938,N_7587);
or U8253 (N_8253,N_7840,N_7924);
or U8254 (N_8254,N_7840,N_7662);
and U8255 (N_8255,N_7630,N_7761);
nand U8256 (N_8256,N_7587,N_7627);
nand U8257 (N_8257,N_7732,N_7604);
or U8258 (N_8258,N_7909,N_7880);
or U8259 (N_8259,N_7662,N_7846);
nor U8260 (N_8260,N_7971,N_7934);
and U8261 (N_8261,N_7674,N_7950);
nand U8262 (N_8262,N_7656,N_7576);
nor U8263 (N_8263,N_7909,N_7908);
and U8264 (N_8264,N_7503,N_7755);
xor U8265 (N_8265,N_7577,N_7507);
nor U8266 (N_8266,N_7935,N_7621);
nand U8267 (N_8267,N_7564,N_7698);
or U8268 (N_8268,N_7599,N_7630);
nand U8269 (N_8269,N_7954,N_7699);
nor U8270 (N_8270,N_7580,N_7994);
nor U8271 (N_8271,N_7964,N_7693);
xnor U8272 (N_8272,N_7542,N_7902);
nor U8273 (N_8273,N_7618,N_7712);
or U8274 (N_8274,N_7914,N_7787);
or U8275 (N_8275,N_7729,N_7768);
xnor U8276 (N_8276,N_7966,N_7682);
xnor U8277 (N_8277,N_7501,N_7944);
nor U8278 (N_8278,N_7966,N_7736);
or U8279 (N_8279,N_7973,N_7587);
nor U8280 (N_8280,N_7579,N_7909);
xnor U8281 (N_8281,N_7754,N_7796);
xnor U8282 (N_8282,N_7571,N_7985);
nand U8283 (N_8283,N_7891,N_7912);
or U8284 (N_8284,N_7920,N_7913);
nand U8285 (N_8285,N_7911,N_7992);
and U8286 (N_8286,N_7665,N_7752);
nand U8287 (N_8287,N_7997,N_7769);
xnor U8288 (N_8288,N_7594,N_7932);
nand U8289 (N_8289,N_7864,N_7773);
nand U8290 (N_8290,N_7761,N_7756);
xor U8291 (N_8291,N_7647,N_7690);
or U8292 (N_8292,N_7724,N_7712);
and U8293 (N_8293,N_7515,N_7776);
or U8294 (N_8294,N_7593,N_7764);
and U8295 (N_8295,N_7958,N_7941);
xnor U8296 (N_8296,N_7559,N_7606);
xor U8297 (N_8297,N_7920,N_7609);
and U8298 (N_8298,N_7896,N_7859);
nand U8299 (N_8299,N_7624,N_7639);
nand U8300 (N_8300,N_7888,N_7713);
and U8301 (N_8301,N_7697,N_7773);
xnor U8302 (N_8302,N_7832,N_7879);
nor U8303 (N_8303,N_7732,N_7952);
and U8304 (N_8304,N_7693,N_7812);
or U8305 (N_8305,N_7824,N_7716);
nand U8306 (N_8306,N_7592,N_7681);
and U8307 (N_8307,N_7996,N_7936);
xnor U8308 (N_8308,N_7798,N_7860);
xor U8309 (N_8309,N_7656,N_7511);
nor U8310 (N_8310,N_7835,N_7804);
and U8311 (N_8311,N_7951,N_7987);
nor U8312 (N_8312,N_7692,N_7758);
or U8313 (N_8313,N_7577,N_7687);
and U8314 (N_8314,N_7796,N_7851);
nor U8315 (N_8315,N_7968,N_7619);
xor U8316 (N_8316,N_7768,N_7932);
nor U8317 (N_8317,N_7874,N_7697);
xnor U8318 (N_8318,N_7892,N_7779);
and U8319 (N_8319,N_7862,N_7699);
and U8320 (N_8320,N_7894,N_7620);
or U8321 (N_8321,N_7607,N_7525);
nor U8322 (N_8322,N_7794,N_7970);
or U8323 (N_8323,N_7768,N_7710);
or U8324 (N_8324,N_7791,N_7723);
or U8325 (N_8325,N_7732,N_7613);
nor U8326 (N_8326,N_7576,N_7777);
or U8327 (N_8327,N_7678,N_7631);
nand U8328 (N_8328,N_7912,N_7567);
xor U8329 (N_8329,N_7660,N_7995);
nand U8330 (N_8330,N_7588,N_7917);
or U8331 (N_8331,N_7948,N_7860);
or U8332 (N_8332,N_7544,N_7519);
and U8333 (N_8333,N_7695,N_7909);
or U8334 (N_8334,N_7894,N_7767);
xnor U8335 (N_8335,N_7563,N_7681);
nor U8336 (N_8336,N_7581,N_7609);
or U8337 (N_8337,N_7912,N_7586);
nor U8338 (N_8338,N_7684,N_7598);
or U8339 (N_8339,N_7987,N_7694);
or U8340 (N_8340,N_7895,N_7808);
nand U8341 (N_8341,N_7853,N_7698);
or U8342 (N_8342,N_7622,N_7641);
and U8343 (N_8343,N_7850,N_7797);
xnor U8344 (N_8344,N_7830,N_7704);
and U8345 (N_8345,N_7568,N_7536);
or U8346 (N_8346,N_7612,N_7884);
nand U8347 (N_8347,N_7936,N_7950);
xor U8348 (N_8348,N_7628,N_7856);
and U8349 (N_8349,N_7865,N_7943);
xnor U8350 (N_8350,N_7953,N_7634);
nor U8351 (N_8351,N_7507,N_7785);
and U8352 (N_8352,N_7623,N_7651);
xnor U8353 (N_8353,N_7805,N_7553);
and U8354 (N_8354,N_7677,N_7512);
nand U8355 (N_8355,N_7551,N_7665);
or U8356 (N_8356,N_7926,N_7764);
xor U8357 (N_8357,N_7812,N_7843);
nand U8358 (N_8358,N_7596,N_7799);
nor U8359 (N_8359,N_7697,N_7598);
nor U8360 (N_8360,N_7843,N_7511);
or U8361 (N_8361,N_7940,N_7724);
nand U8362 (N_8362,N_7666,N_7675);
nor U8363 (N_8363,N_7678,N_7915);
nor U8364 (N_8364,N_7614,N_7697);
and U8365 (N_8365,N_7968,N_7655);
nor U8366 (N_8366,N_7568,N_7777);
and U8367 (N_8367,N_7747,N_7653);
and U8368 (N_8368,N_7678,N_7668);
or U8369 (N_8369,N_7735,N_7985);
nor U8370 (N_8370,N_7822,N_7874);
nor U8371 (N_8371,N_7759,N_7512);
nand U8372 (N_8372,N_7669,N_7767);
and U8373 (N_8373,N_7775,N_7975);
nand U8374 (N_8374,N_7673,N_7943);
nand U8375 (N_8375,N_7944,N_7741);
nand U8376 (N_8376,N_7967,N_7900);
and U8377 (N_8377,N_7922,N_7934);
nor U8378 (N_8378,N_7933,N_7837);
or U8379 (N_8379,N_7877,N_7819);
xor U8380 (N_8380,N_7680,N_7632);
or U8381 (N_8381,N_7844,N_7977);
xnor U8382 (N_8382,N_7514,N_7968);
xor U8383 (N_8383,N_7671,N_7787);
xor U8384 (N_8384,N_7620,N_7592);
nor U8385 (N_8385,N_7616,N_7503);
nor U8386 (N_8386,N_7862,N_7521);
xor U8387 (N_8387,N_7838,N_7843);
nor U8388 (N_8388,N_7984,N_7975);
nand U8389 (N_8389,N_7741,N_7839);
xor U8390 (N_8390,N_7810,N_7845);
nor U8391 (N_8391,N_7716,N_7523);
nand U8392 (N_8392,N_7767,N_7933);
or U8393 (N_8393,N_7609,N_7799);
nand U8394 (N_8394,N_7569,N_7655);
and U8395 (N_8395,N_7889,N_7846);
and U8396 (N_8396,N_7939,N_7533);
nand U8397 (N_8397,N_7784,N_7938);
and U8398 (N_8398,N_7575,N_7613);
nor U8399 (N_8399,N_7501,N_7565);
or U8400 (N_8400,N_7661,N_7533);
nand U8401 (N_8401,N_7938,N_7921);
xnor U8402 (N_8402,N_7743,N_7882);
nand U8403 (N_8403,N_7616,N_7731);
and U8404 (N_8404,N_7534,N_7791);
nor U8405 (N_8405,N_7915,N_7600);
or U8406 (N_8406,N_7942,N_7771);
and U8407 (N_8407,N_7571,N_7540);
nor U8408 (N_8408,N_7891,N_7738);
or U8409 (N_8409,N_7830,N_7538);
xnor U8410 (N_8410,N_7790,N_7982);
or U8411 (N_8411,N_7724,N_7934);
nor U8412 (N_8412,N_7647,N_7585);
nand U8413 (N_8413,N_7540,N_7882);
xor U8414 (N_8414,N_7803,N_7931);
and U8415 (N_8415,N_7998,N_7534);
nand U8416 (N_8416,N_7627,N_7893);
xnor U8417 (N_8417,N_7771,N_7916);
or U8418 (N_8418,N_7644,N_7802);
nand U8419 (N_8419,N_7704,N_7658);
xor U8420 (N_8420,N_7558,N_7790);
nand U8421 (N_8421,N_7515,N_7632);
or U8422 (N_8422,N_7713,N_7726);
nor U8423 (N_8423,N_7705,N_7505);
and U8424 (N_8424,N_7985,N_7576);
nand U8425 (N_8425,N_7532,N_7774);
xnor U8426 (N_8426,N_7869,N_7537);
xnor U8427 (N_8427,N_7873,N_7869);
xor U8428 (N_8428,N_7995,N_7849);
and U8429 (N_8429,N_7796,N_7591);
xor U8430 (N_8430,N_7570,N_7672);
nand U8431 (N_8431,N_7960,N_7687);
xnor U8432 (N_8432,N_7566,N_7578);
and U8433 (N_8433,N_7991,N_7700);
and U8434 (N_8434,N_7939,N_7509);
and U8435 (N_8435,N_7744,N_7544);
nor U8436 (N_8436,N_7556,N_7893);
or U8437 (N_8437,N_7924,N_7930);
or U8438 (N_8438,N_7604,N_7758);
xnor U8439 (N_8439,N_7589,N_7983);
or U8440 (N_8440,N_7623,N_7911);
xnor U8441 (N_8441,N_7827,N_7737);
or U8442 (N_8442,N_7965,N_7876);
nand U8443 (N_8443,N_7611,N_7928);
and U8444 (N_8444,N_7923,N_7708);
nand U8445 (N_8445,N_7817,N_7834);
and U8446 (N_8446,N_7596,N_7632);
or U8447 (N_8447,N_7885,N_7636);
nand U8448 (N_8448,N_7563,N_7829);
nor U8449 (N_8449,N_7955,N_7854);
or U8450 (N_8450,N_7626,N_7564);
and U8451 (N_8451,N_7860,N_7554);
nor U8452 (N_8452,N_7534,N_7682);
xnor U8453 (N_8453,N_7788,N_7681);
xor U8454 (N_8454,N_7738,N_7769);
xor U8455 (N_8455,N_7655,N_7557);
nor U8456 (N_8456,N_7908,N_7878);
or U8457 (N_8457,N_7984,N_7546);
nand U8458 (N_8458,N_7738,N_7566);
nor U8459 (N_8459,N_7665,N_7722);
nand U8460 (N_8460,N_7703,N_7524);
or U8461 (N_8461,N_7650,N_7909);
and U8462 (N_8462,N_7731,N_7798);
xnor U8463 (N_8463,N_7988,N_7652);
xor U8464 (N_8464,N_7600,N_7508);
xor U8465 (N_8465,N_7974,N_7598);
nand U8466 (N_8466,N_7770,N_7513);
nand U8467 (N_8467,N_7657,N_7634);
xnor U8468 (N_8468,N_7505,N_7926);
and U8469 (N_8469,N_7883,N_7764);
or U8470 (N_8470,N_7993,N_7856);
and U8471 (N_8471,N_7714,N_7642);
nand U8472 (N_8472,N_7752,N_7608);
xor U8473 (N_8473,N_7570,N_7987);
xnor U8474 (N_8474,N_7622,N_7590);
or U8475 (N_8475,N_7840,N_7655);
nand U8476 (N_8476,N_7560,N_7879);
nor U8477 (N_8477,N_7853,N_7701);
or U8478 (N_8478,N_7652,N_7895);
nand U8479 (N_8479,N_7506,N_7884);
nand U8480 (N_8480,N_7519,N_7784);
and U8481 (N_8481,N_7965,N_7647);
nand U8482 (N_8482,N_7641,N_7778);
and U8483 (N_8483,N_7995,N_7639);
or U8484 (N_8484,N_7889,N_7979);
nand U8485 (N_8485,N_7532,N_7792);
xor U8486 (N_8486,N_7514,N_7528);
xnor U8487 (N_8487,N_7983,N_7622);
xor U8488 (N_8488,N_7873,N_7663);
and U8489 (N_8489,N_7917,N_7815);
nand U8490 (N_8490,N_7947,N_7642);
nand U8491 (N_8491,N_7745,N_7778);
and U8492 (N_8492,N_7750,N_7643);
and U8493 (N_8493,N_7662,N_7701);
nand U8494 (N_8494,N_7974,N_7697);
and U8495 (N_8495,N_7670,N_7632);
and U8496 (N_8496,N_7993,N_7806);
or U8497 (N_8497,N_7537,N_7733);
xnor U8498 (N_8498,N_7841,N_7672);
nand U8499 (N_8499,N_7987,N_7603);
or U8500 (N_8500,N_8382,N_8282);
nand U8501 (N_8501,N_8375,N_8286);
nand U8502 (N_8502,N_8099,N_8184);
nor U8503 (N_8503,N_8125,N_8157);
xnor U8504 (N_8504,N_8136,N_8002);
and U8505 (N_8505,N_8141,N_8485);
and U8506 (N_8506,N_8143,N_8399);
xor U8507 (N_8507,N_8460,N_8070);
and U8508 (N_8508,N_8358,N_8253);
nand U8509 (N_8509,N_8083,N_8271);
nor U8510 (N_8510,N_8440,N_8360);
and U8511 (N_8511,N_8024,N_8031);
nand U8512 (N_8512,N_8321,N_8110);
xor U8513 (N_8513,N_8473,N_8349);
nand U8514 (N_8514,N_8380,N_8322);
and U8515 (N_8515,N_8305,N_8295);
xor U8516 (N_8516,N_8425,N_8023);
nand U8517 (N_8517,N_8198,N_8032);
and U8518 (N_8518,N_8405,N_8145);
xnor U8519 (N_8519,N_8042,N_8272);
and U8520 (N_8520,N_8071,N_8302);
nor U8521 (N_8521,N_8325,N_8021);
xor U8522 (N_8522,N_8045,N_8087);
xnor U8523 (N_8523,N_8011,N_8117);
nand U8524 (N_8524,N_8338,N_8390);
xnor U8525 (N_8525,N_8014,N_8298);
and U8526 (N_8526,N_8151,N_8140);
xnor U8527 (N_8527,N_8212,N_8126);
nand U8528 (N_8528,N_8100,N_8447);
xor U8529 (N_8529,N_8268,N_8118);
or U8530 (N_8530,N_8420,N_8205);
nor U8531 (N_8531,N_8097,N_8211);
and U8532 (N_8532,N_8171,N_8057);
nand U8533 (N_8533,N_8478,N_8464);
or U8534 (N_8534,N_8038,N_8389);
or U8535 (N_8535,N_8467,N_8299);
and U8536 (N_8536,N_8189,N_8104);
and U8537 (N_8537,N_8444,N_8487);
nor U8538 (N_8538,N_8372,N_8159);
or U8539 (N_8539,N_8086,N_8498);
nand U8540 (N_8540,N_8028,N_8085);
xor U8541 (N_8541,N_8470,N_8328);
nor U8542 (N_8542,N_8000,N_8162);
nor U8543 (N_8543,N_8240,N_8155);
nor U8544 (N_8544,N_8278,N_8101);
and U8545 (N_8545,N_8292,N_8297);
xnor U8546 (N_8546,N_8401,N_8237);
nor U8547 (N_8547,N_8267,N_8483);
nor U8548 (N_8548,N_8041,N_8061);
nand U8549 (N_8549,N_8427,N_8105);
nand U8550 (N_8550,N_8130,N_8144);
xnor U8551 (N_8551,N_8453,N_8304);
or U8552 (N_8552,N_8471,N_8040);
xnor U8553 (N_8553,N_8074,N_8192);
nand U8554 (N_8554,N_8256,N_8030);
nor U8555 (N_8555,N_8003,N_8181);
and U8556 (N_8556,N_8497,N_8044);
xnor U8557 (N_8557,N_8309,N_8323);
or U8558 (N_8558,N_8046,N_8356);
and U8559 (N_8559,N_8452,N_8276);
xor U8560 (N_8560,N_8300,N_8343);
xnor U8561 (N_8561,N_8377,N_8182);
nand U8562 (N_8562,N_8076,N_8357);
or U8563 (N_8563,N_8482,N_8008);
and U8564 (N_8564,N_8465,N_8430);
and U8565 (N_8565,N_8163,N_8310);
xor U8566 (N_8566,N_8232,N_8345);
xor U8567 (N_8567,N_8426,N_8431);
or U8568 (N_8568,N_8314,N_8194);
nor U8569 (N_8569,N_8180,N_8006);
or U8570 (N_8570,N_8007,N_8206);
xnor U8571 (N_8571,N_8224,N_8026);
nor U8572 (N_8572,N_8201,N_8213);
nor U8573 (N_8573,N_8396,N_8436);
or U8574 (N_8574,N_8102,N_8387);
nor U8575 (N_8575,N_8226,N_8468);
nor U8576 (N_8576,N_8274,N_8318);
xor U8577 (N_8577,N_8039,N_8152);
nor U8578 (N_8578,N_8234,N_8403);
and U8579 (N_8579,N_8113,N_8033);
nor U8580 (N_8580,N_8219,N_8016);
xnor U8581 (N_8581,N_8209,N_8166);
or U8582 (N_8582,N_8019,N_8022);
xor U8583 (N_8583,N_8441,N_8429);
and U8584 (N_8584,N_8288,N_8348);
or U8585 (N_8585,N_8103,N_8280);
xor U8586 (N_8586,N_8443,N_8066);
nand U8587 (N_8587,N_8036,N_8269);
nor U8588 (N_8588,N_8190,N_8183);
nand U8589 (N_8589,N_8415,N_8456);
and U8590 (N_8590,N_8106,N_8439);
or U8591 (N_8591,N_8058,N_8174);
or U8592 (N_8592,N_8170,N_8012);
nand U8593 (N_8593,N_8463,N_8290);
or U8594 (N_8594,N_8250,N_8121);
or U8595 (N_8595,N_8404,N_8340);
or U8596 (N_8596,N_8249,N_8373);
and U8597 (N_8597,N_8147,N_8433);
nand U8598 (N_8598,N_8247,N_8413);
or U8599 (N_8599,N_8341,N_8359);
nand U8600 (N_8600,N_8394,N_8095);
xor U8601 (N_8601,N_8499,N_8411);
and U8602 (N_8602,N_8417,N_8385);
nor U8603 (N_8603,N_8203,N_8284);
or U8604 (N_8604,N_8197,N_8167);
nor U8605 (N_8605,N_8236,N_8037);
and U8606 (N_8606,N_8111,N_8052);
or U8607 (N_8607,N_8214,N_8260);
xor U8608 (N_8608,N_8296,N_8324);
and U8609 (N_8609,N_8369,N_8200);
or U8610 (N_8610,N_8418,N_8149);
nand U8611 (N_8611,N_8294,N_8313);
and U8612 (N_8612,N_8277,N_8017);
or U8613 (N_8613,N_8388,N_8090);
nor U8614 (N_8614,N_8367,N_8450);
xnor U8615 (N_8615,N_8075,N_8263);
nand U8616 (N_8616,N_8069,N_8080);
nand U8617 (N_8617,N_8225,N_8361);
nand U8618 (N_8618,N_8254,N_8491);
or U8619 (N_8619,N_8333,N_8091);
xor U8620 (N_8620,N_8207,N_8217);
and U8621 (N_8621,N_8476,N_8398);
xnor U8622 (N_8622,N_8025,N_8013);
and U8623 (N_8623,N_8336,N_8408);
and U8624 (N_8624,N_8005,N_8400);
or U8625 (N_8625,N_8352,N_8128);
nor U8626 (N_8626,N_8480,N_8275);
and U8627 (N_8627,N_8466,N_8034);
and U8628 (N_8628,N_8407,N_8156);
and U8629 (N_8629,N_8176,N_8489);
nand U8630 (N_8630,N_8457,N_8451);
and U8631 (N_8631,N_8368,N_8204);
and U8632 (N_8632,N_8273,N_8244);
nand U8633 (N_8633,N_8409,N_8172);
nand U8634 (N_8634,N_8437,N_8255);
and U8635 (N_8635,N_8216,N_8096);
xnor U8636 (N_8636,N_8406,N_8289);
nand U8637 (N_8637,N_8353,N_8379);
and U8638 (N_8638,N_8065,N_8494);
xnor U8639 (N_8639,N_8238,N_8371);
or U8640 (N_8640,N_8123,N_8208);
or U8641 (N_8641,N_8261,N_8291);
or U8642 (N_8642,N_8376,N_8119);
or U8643 (N_8643,N_8161,N_8412);
nor U8644 (N_8644,N_8374,N_8495);
nand U8645 (N_8645,N_8266,N_8312);
nand U8646 (N_8646,N_8461,N_8073);
or U8647 (N_8647,N_8384,N_8428);
and U8648 (N_8648,N_8316,N_8484);
xnor U8649 (N_8649,N_8093,N_8233);
nand U8650 (N_8650,N_8241,N_8293);
xor U8651 (N_8651,N_8397,N_8332);
xnor U8652 (N_8652,N_8009,N_8317);
xor U8653 (N_8653,N_8010,N_8004);
or U8654 (N_8654,N_8218,N_8112);
and U8655 (N_8655,N_8252,N_8001);
and U8656 (N_8656,N_8049,N_8445);
xnor U8657 (N_8657,N_8364,N_8424);
nand U8658 (N_8658,N_8175,N_8235);
nor U8659 (N_8659,N_8472,N_8048);
nand U8660 (N_8660,N_8285,N_8474);
nand U8661 (N_8661,N_8133,N_8239);
or U8662 (N_8662,N_8169,N_8094);
and U8663 (N_8663,N_8421,N_8281);
xnor U8664 (N_8664,N_8265,N_8077);
nand U8665 (N_8665,N_8381,N_8362);
nand U8666 (N_8666,N_8446,N_8221);
or U8667 (N_8667,N_8138,N_8060);
or U8668 (N_8668,N_8423,N_8186);
or U8669 (N_8669,N_8477,N_8088);
xor U8670 (N_8670,N_8243,N_8259);
xor U8671 (N_8671,N_8185,N_8168);
or U8672 (N_8672,N_8137,N_8462);
xor U8673 (N_8673,N_8109,N_8496);
xnor U8674 (N_8674,N_8363,N_8393);
and U8675 (N_8675,N_8245,N_8391);
or U8676 (N_8676,N_8246,N_8370);
xnor U8677 (N_8677,N_8050,N_8248);
nor U8678 (N_8678,N_8195,N_8416);
xor U8679 (N_8679,N_8178,N_8301);
or U8680 (N_8680,N_8355,N_8479);
xor U8681 (N_8681,N_8223,N_8230);
xnor U8682 (N_8682,N_8351,N_8366);
xnor U8683 (N_8683,N_8442,N_8222);
nand U8684 (N_8684,N_8064,N_8078);
xor U8685 (N_8685,N_8438,N_8308);
xnor U8686 (N_8686,N_8054,N_8220);
nor U8687 (N_8687,N_8434,N_8432);
nor U8688 (N_8688,N_8165,N_8350);
nand U8689 (N_8689,N_8191,N_8386);
nand U8690 (N_8690,N_8469,N_8383);
or U8691 (N_8691,N_8062,N_8056);
or U8692 (N_8692,N_8402,N_8067);
or U8693 (N_8693,N_8326,N_8481);
or U8694 (N_8694,N_8320,N_8081);
nor U8695 (N_8695,N_8029,N_8047);
xnor U8696 (N_8696,N_8459,N_8334);
nand U8697 (N_8697,N_8122,N_8392);
nand U8698 (N_8698,N_8173,N_8262);
or U8699 (N_8699,N_8327,N_8134);
nor U8700 (N_8700,N_8303,N_8492);
xor U8701 (N_8701,N_8229,N_8187);
nor U8702 (N_8702,N_8072,N_8132);
and U8703 (N_8703,N_8455,N_8177);
or U8704 (N_8704,N_8055,N_8135);
nand U8705 (N_8705,N_8129,N_8231);
nor U8706 (N_8706,N_8053,N_8330);
and U8707 (N_8707,N_8127,N_8116);
xor U8708 (N_8708,N_8458,N_8311);
nand U8709 (N_8709,N_8108,N_8329);
and U8710 (N_8710,N_8346,N_8270);
or U8711 (N_8711,N_8092,N_8114);
and U8712 (N_8712,N_8419,N_8154);
xnor U8713 (N_8713,N_8242,N_8339);
or U8714 (N_8714,N_8018,N_8258);
nor U8715 (N_8715,N_8414,N_8035);
and U8716 (N_8716,N_8027,N_8068);
xor U8717 (N_8717,N_8486,N_8410);
xnor U8718 (N_8718,N_8279,N_8059);
xor U8719 (N_8719,N_8210,N_8079);
nor U8720 (N_8720,N_8063,N_8365);
and U8721 (N_8721,N_8347,N_8488);
xnor U8722 (N_8722,N_8158,N_8084);
nand U8723 (N_8723,N_8082,N_8315);
nand U8724 (N_8724,N_8139,N_8454);
and U8725 (N_8725,N_8344,N_8493);
xnor U8726 (N_8726,N_8257,N_8227);
nor U8727 (N_8727,N_8264,N_8089);
nor U8728 (N_8728,N_8150,N_8307);
nor U8729 (N_8729,N_8107,N_8342);
or U8730 (N_8730,N_8422,N_8043);
xnor U8731 (N_8731,N_8475,N_8337);
and U8732 (N_8732,N_8306,N_8164);
nand U8733 (N_8733,N_8193,N_8287);
xnor U8734 (N_8734,N_8124,N_8435);
xnor U8735 (N_8735,N_8354,N_8020);
nand U8736 (N_8736,N_8115,N_8283);
xor U8737 (N_8737,N_8160,N_8251);
or U8738 (N_8738,N_8015,N_8131);
nor U8739 (N_8739,N_8199,N_8142);
xnor U8740 (N_8740,N_8490,N_8395);
xor U8741 (N_8741,N_8153,N_8196);
nand U8742 (N_8742,N_8148,N_8228);
nand U8743 (N_8743,N_8319,N_8098);
nand U8744 (N_8744,N_8448,N_8215);
or U8745 (N_8745,N_8202,N_8120);
and U8746 (N_8746,N_8331,N_8146);
xnor U8747 (N_8747,N_8179,N_8449);
and U8748 (N_8748,N_8051,N_8188);
or U8749 (N_8749,N_8335,N_8378);
nor U8750 (N_8750,N_8381,N_8146);
or U8751 (N_8751,N_8397,N_8032);
xnor U8752 (N_8752,N_8012,N_8297);
nor U8753 (N_8753,N_8371,N_8432);
or U8754 (N_8754,N_8477,N_8307);
xor U8755 (N_8755,N_8156,N_8215);
and U8756 (N_8756,N_8236,N_8304);
nor U8757 (N_8757,N_8380,N_8210);
and U8758 (N_8758,N_8393,N_8361);
or U8759 (N_8759,N_8216,N_8393);
nand U8760 (N_8760,N_8437,N_8186);
xnor U8761 (N_8761,N_8010,N_8446);
or U8762 (N_8762,N_8227,N_8275);
and U8763 (N_8763,N_8318,N_8439);
nor U8764 (N_8764,N_8389,N_8058);
nand U8765 (N_8765,N_8352,N_8403);
and U8766 (N_8766,N_8248,N_8214);
xor U8767 (N_8767,N_8125,N_8272);
nand U8768 (N_8768,N_8377,N_8453);
xor U8769 (N_8769,N_8215,N_8007);
or U8770 (N_8770,N_8168,N_8123);
or U8771 (N_8771,N_8389,N_8379);
nand U8772 (N_8772,N_8407,N_8448);
or U8773 (N_8773,N_8377,N_8083);
xor U8774 (N_8774,N_8123,N_8158);
nand U8775 (N_8775,N_8347,N_8154);
and U8776 (N_8776,N_8432,N_8478);
or U8777 (N_8777,N_8336,N_8299);
nor U8778 (N_8778,N_8094,N_8073);
or U8779 (N_8779,N_8351,N_8390);
nor U8780 (N_8780,N_8251,N_8413);
or U8781 (N_8781,N_8017,N_8142);
and U8782 (N_8782,N_8301,N_8480);
nand U8783 (N_8783,N_8375,N_8331);
nor U8784 (N_8784,N_8139,N_8293);
nor U8785 (N_8785,N_8016,N_8048);
and U8786 (N_8786,N_8372,N_8193);
or U8787 (N_8787,N_8204,N_8499);
nand U8788 (N_8788,N_8337,N_8133);
or U8789 (N_8789,N_8410,N_8117);
nand U8790 (N_8790,N_8384,N_8053);
nand U8791 (N_8791,N_8140,N_8428);
or U8792 (N_8792,N_8053,N_8014);
nor U8793 (N_8793,N_8394,N_8184);
or U8794 (N_8794,N_8166,N_8411);
nand U8795 (N_8795,N_8250,N_8107);
and U8796 (N_8796,N_8082,N_8104);
nor U8797 (N_8797,N_8435,N_8479);
nand U8798 (N_8798,N_8206,N_8190);
or U8799 (N_8799,N_8081,N_8191);
and U8800 (N_8800,N_8445,N_8193);
nor U8801 (N_8801,N_8447,N_8136);
xor U8802 (N_8802,N_8153,N_8223);
nor U8803 (N_8803,N_8157,N_8248);
xnor U8804 (N_8804,N_8366,N_8111);
or U8805 (N_8805,N_8271,N_8454);
and U8806 (N_8806,N_8281,N_8182);
and U8807 (N_8807,N_8255,N_8181);
or U8808 (N_8808,N_8181,N_8122);
xor U8809 (N_8809,N_8310,N_8222);
nor U8810 (N_8810,N_8227,N_8104);
nand U8811 (N_8811,N_8222,N_8388);
xor U8812 (N_8812,N_8457,N_8339);
xnor U8813 (N_8813,N_8433,N_8195);
nand U8814 (N_8814,N_8209,N_8113);
nor U8815 (N_8815,N_8466,N_8369);
xor U8816 (N_8816,N_8181,N_8071);
nand U8817 (N_8817,N_8234,N_8269);
and U8818 (N_8818,N_8337,N_8168);
nand U8819 (N_8819,N_8266,N_8268);
nand U8820 (N_8820,N_8056,N_8277);
nand U8821 (N_8821,N_8156,N_8391);
xor U8822 (N_8822,N_8074,N_8079);
nor U8823 (N_8823,N_8169,N_8379);
or U8824 (N_8824,N_8060,N_8366);
or U8825 (N_8825,N_8091,N_8214);
nand U8826 (N_8826,N_8285,N_8198);
and U8827 (N_8827,N_8459,N_8471);
or U8828 (N_8828,N_8181,N_8262);
nor U8829 (N_8829,N_8087,N_8300);
nand U8830 (N_8830,N_8379,N_8165);
and U8831 (N_8831,N_8451,N_8153);
nand U8832 (N_8832,N_8468,N_8391);
and U8833 (N_8833,N_8300,N_8178);
or U8834 (N_8834,N_8295,N_8105);
xor U8835 (N_8835,N_8374,N_8010);
nand U8836 (N_8836,N_8423,N_8309);
nand U8837 (N_8837,N_8069,N_8094);
and U8838 (N_8838,N_8160,N_8244);
or U8839 (N_8839,N_8379,N_8174);
nor U8840 (N_8840,N_8129,N_8152);
nor U8841 (N_8841,N_8338,N_8414);
xor U8842 (N_8842,N_8123,N_8349);
xnor U8843 (N_8843,N_8474,N_8188);
and U8844 (N_8844,N_8054,N_8364);
or U8845 (N_8845,N_8396,N_8427);
and U8846 (N_8846,N_8258,N_8021);
or U8847 (N_8847,N_8419,N_8110);
or U8848 (N_8848,N_8247,N_8320);
nor U8849 (N_8849,N_8096,N_8168);
or U8850 (N_8850,N_8347,N_8165);
nor U8851 (N_8851,N_8089,N_8063);
nor U8852 (N_8852,N_8108,N_8080);
and U8853 (N_8853,N_8269,N_8407);
nand U8854 (N_8854,N_8165,N_8393);
and U8855 (N_8855,N_8000,N_8072);
or U8856 (N_8856,N_8186,N_8008);
nand U8857 (N_8857,N_8150,N_8481);
nor U8858 (N_8858,N_8430,N_8124);
and U8859 (N_8859,N_8484,N_8442);
xor U8860 (N_8860,N_8378,N_8018);
xnor U8861 (N_8861,N_8381,N_8238);
nor U8862 (N_8862,N_8311,N_8400);
nor U8863 (N_8863,N_8004,N_8001);
nand U8864 (N_8864,N_8287,N_8420);
nand U8865 (N_8865,N_8214,N_8083);
xnor U8866 (N_8866,N_8193,N_8237);
or U8867 (N_8867,N_8048,N_8341);
nor U8868 (N_8868,N_8190,N_8334);
nor U8869 (N_8869,N_8340,N_8457);
xnor U8870 (N_8870,N_8174,N_8139);
or U8871 (N_8871,N_8468,N_8187);
or U8872 (N_8872,N_8365,N_8441);
and U8873 (N_8873,N_8040,N_8074);
nand U8874 (N_8874,N_8146,N_8440);
nand U8875 (N_8875,N_8321,N_8243);
xor U8876 (N_8876,N_8398,N_8262);
nor U8877 (N_8877,N_8132,N_8338);
or U8878 (N_8878,N_8494,N_8248);
xnor U8879 (N_8879,N_8218,N_8140);
nand U8880 (N_8880,N_8297,N_8221);
nor U8881 (N_8881,N_8348,N_8433);
or U8882 (N_8882,N_8326,N_8281);
or U8883 (N_8883,N_8094,N_8228);
nor U8884 (N_8884,N_8372,N_8291);
and U8885 (N_8885,N_8181,N_8032);
xor U8886 (N_8886,N_8388,N_8315);
or U8887 (N_8887,N_8379,N_8283);
xor U8888 (N_8888,N_8080,N_8028);
and U8889 (N_8889,N_8329,N_8320);
nor U8890 (N_8890,N_8330,N_8280);
nor U8891 (N_8891,N_8194,N_8279);
and U8892 (N_8892,N_8026,N_8284);
and U8893 (N_8893,N_8250,N_8326);
and U8894 (N_8894,N_8233,N_8450);
nor U8895 (N_8895,N_8036,N_8225);
xnor U8896 (N_8896,N_8212,N_8032);
xor U8897 (N_8897,N_8060,N_8377);
xor U8898 (N_8898,N_8412,N_8376);
nand U8899 (N_8899,N_8314,N_8479);
and U8900 (N_8900,N_8316,N_8256);
xor U8901 (N_8901,N_8026,N_8395);
xnor U8902 (N_8902,N_8255,N_8374);
nor U8903 (N_8903,N_8205,N_8299);
nand U8904 (N_8904,N_8021,N_8102);
or U8905 (N_8905,N_8015,N_8386);
xnor U8906 (N_8906,N_8260,N_8468);
xnor U8907 (N_8907,N_8030,N_8001);
nor U8908 (N_8908,N_8246,N_8182);
or U8909 (N_8909,N_8350,N_8349);
xnor U8910 (N_8910,N_8158,N_8473);
and U8911 (N_8911,N_8327,N_8222);
nor U8912 (N_8912,N_8388,N_8193);
xnor U8913 (N_8913,N_8311,N_8091);
xor U8914 (N_8914,N_8380,N_8454);
and U8915 (N_8915,N_8090,N_8025);
or U8916 (N_8916,N_8114,N_8421);
or U8917 (N_8917,N_8194,N_8078);
xnor U8918 (N_8918,N_8307,N_8373);
or U8919 (N_8919,N_8316,N_8173);
nor U8920 (N_8920,N_8448,N_8031);
nand U8921 (N_8921,N_8257,N_8341);
xor U8922 (N_8922,N_8410,N_8289);
and U8923 (N_8923,N_8325,N_8367);
and U8924 (N_8924,N_8039,N_8437);
nor U8925 (N_8925,N_8402,N_8423);
or U8926 (N_8926,N_8059,N_8062);
and U8927 (N_8927,N_8435,N_8351);
nand U8928 (N_8928,N_8497,N_8081);
or U8929 (N_8929,N_8473,N_8408);
and U8930 (N_8930,N_8099,N_8072);
nor U8931 (N_8931,N_8258,N_8244);
xnor U8932 (N_8932,N_8260,N_8199);
nand U8933 (N_8933,N_8057,N_8118);
nand U8934 (N_8934,N_8338,N_8095);
and U8935 (N_8935,N_8355,N_8319);
xor U8936 (N_8936,N_8072,N_8195);
and U8937 (N_8937,N_8414,N_8296);
or U8938 (N_8938,N_8185,N_8118);
or U8939 (N_8939,N_8488,N_8136);
nor U8940 (N_8940,N_8117,N_8475);
and U8941 (N_8941,N_8379,N_8072);
nor U8942 (N_8942,N_8005,N_8418);
nand U8943 (N_8943,N_8182,N_8395);
and U8944 (N_8944,N_8405,N_8261);
xor U8945 (N_8945,N_8347,N_8467);
nor U8946 (N_8946,N_8172,N_8299);
nand U8947 (N_8947,N_8170,N_8326);
nor U8948 (N_8948,N_8051,N_8278);
nor U8949 (N_8949,N_8139,N_8155);
nor U8950 (N_8950,N_8280,N_8425);
xnor U8951 (N_8951,N_8248,N_8189);
or U8952 (N_8952,N_8079,N_8082);
nor U8953 (N_8953,N_8428,N_8243);
xor U8954 (N_8954,N_8272,N_8011);
xor U8955 (N_8955,N_8301,N_8496);
nand U8956 (N_8956,N_8255,N_8211);
or U8957 (N_8957,N_8017,N_8297);
or U8958 (N_8958,N_8052,N_8320);
xnor U8959 (N_8959,N_8137,N_8141);
or U8960 (N_8960,N_8212,N_8284);
nor U8961 (N_8961,N_8260,N_8144);
and U8962 (N_8962,N_8444,N_8299);
or U8963 (N_8963,N_8308,N_8018);
and U8964 (N_8964,N_8480,N_8484);
nand U8965 (N_8965,N_8067,N_8391);
and U8966 (N_8966,N_8082,N_8437);
or U8967 (N_8967,N_8429,N_8030);
xnor U8968 (N_8968,N_8048,N_8357);
nand U8969 (N_8969,N_8424,N_8138);
nand U8970 (N_8970,N_8311,N_8385);
and U8971 (N_8971,N_8067,N_8253);
or U8972 (N_8972,N_8094,N_8145);
or U8973 (N_8973,N_8253,N_8290);
and U8974 (N_8974,N_8392,N_8150);
and U8975 (N_8975,N_8360,N_8366);
or U8976 (N_8976,N_8462,N_8154);
nor U8977 (N_8977,N_8167,N_8069);
nor U8978 (N_8978,N_8282,N_8146);
nor U8979 (N_8979,N_8298,N_8190);
xor U8980 (N_8980,N_8380,N_8109);
nor U8981 (N_8981,N_8175,N_8249);
nand U8982 (N_8982,N_8353,N_8454);
and U8983 (N_8983,N_8466,N_8029);
nor U8984 (N_8984,N_8134,N_8054);
nand U8985 (N_8985,N_8190,N_8014);
nor U8986 (N_8986,N_8186,N_8381);
or U8987 (N_8987,N_8445,N_8355);
nor U8988 (N_8988,N_8152,N_8119);
and U8989 (N_8989,N_8170,N_8122);
or U8990 (N_8990,N_8045,N_8439);
xnor U8991 (N_8991,N_8189,N_8383);
nand U8992 (N_8992,N_8041,N_8420);
and U8993 (N_8993,N_8054,N_8126);
xnor U8994 (N_8994,N_8111,N_8426);
or U8995 (N_8995,N_8376,N_8332);
and U8996 (N_8996,N_8102,N_8279);
nor U8997 (N_8997,N_8386,N_8260);
nor U8998 (N_8998,N_8336,N_8389);
xnor U8999 (N_8999,N_8383,N_8101);
nand U9000 (N_9000,N_8977,N_8716);
xnor U9001 (N_9001,N_8990,N_8546);
and U9002 (N_9002,N_8866,N_8572);
nand U9003 (N_9003,N_8800,N_8631);
nor U9004 (N_9004,N_8641,N_8931);
nand U9005 (N_9005,N_8764,N_8694);
xor U9006 (N_9006,N_8957,N_8865);
nor U9007 (N_9007,N_8830,N_8843);
nor U9008 (N_9008,N_8605,N_8891);
nand U9009 (N_9009,N_8821,N_8513);
xnor U9010 (N_9010,N_8775,N_8794);
xor U9011 (N_9011,N_8636,N_8619);
nand U9012 (N_9012,N_8786,N_8994);
nand U9013 (N_9013,N_8682,N_8556);
and U9014 (N_9014,N_8599,N_8791);
xor U9015 (N_9015,N_8778,N_8582);
or U9016 (N_9016,N_8686,N_8881);
nand U9017 (N_9017,N_8813,N_8644);
and U9018 (N_9018,N_8525,N_8779);
or U9019 (N_9019,N_8902,N_8624);
or U9020 (N_9020,N_8804,N_8630);
and U9021 (N_9021,N_8917,N_8934);
nand U9022 (N_9022,N_8561,N_8592);
xor U9023 (N_9023,N_8590,N_8846);
nand U9024 (N_9024,N_8862,N_8797);
nand U9025 (N_9025,N_8936,N_8999);
nor U9026 (N_9026,N_8538,N_8566);
nor U9027 (N_9027,N_8688,N_8770);
nor U9028 (N_9028,N_8623,N_8968);
or U9029 (N_9029,N_8913,N_8806);
or U9030 (N_9030,N_8628,N_8746);
and U9031 (N_9031,N_8693,N_8714);
nor U9032 (N_9032,N_8790,N_8594);
or U9033 (N_9033,N_8616,N_8926);
nor U9034 (N_9034,N_8659,N_8591);
nand U9035 (N_9035,N_8820,N_8986);
xnor U9036 (N_9036,N_8515,N_8838);
nor U9037 (N_9037,N_8912,N_8650);
nand U9038 (N_9038,N_8910,N_8577);
and U9039 (N_9039,N_8709,N_8647);
xnor U9040 (N_9040,N_8962,N_8530);
xnor U9041 (N_9041,N_8700,N_8763);
nor U9042 (N_9042,N_8985,N_8979);
or U9043 (N_9043,N_8924,N_8526);
or U9044 (N_9044,N_8640,N_8637);
xnor U9045 (N_9045,N_8516,N_8823);
xnor U9046 (N_9046,N_8504,N_8517);
nand U9047 (N_9047,N_8966,N_8803);
nand U9048 (N_9048,N_8726,N_8661);
and U9049 (N_9049,N_8998,N_8537);
xnor U9050 (N_9050,N_8654,N_8678);
and U9051 (N_9051,N_8787,N_8885);
and U9052 (N_9052,N_8964,N_8534);
or U9053 (N_9053,N_8508,N_8533);
and U9054 (N_9054,N_8564,N_8904);
xor U9055 (N_9055,N_8584,N_8992);
or U9056 (N_9056,N_8818,N_8849);
nor U9057 (N_9057,N_8603,N_8935);
and U9058 (N_9058,N_8684,N_8614);
nand U9059 (N_9059,N_8903,N_8805);
nor U9060 (N_9060,N_8872,N_8907);
or U9061 (N_9061,N_8959,N_8706);
nor U9062 (N_9062,N_8638,N_8698);
nor U9063 (N_9063,N_8595,N_8674);
xnor U9064 (N_9064,N_8544,N_8611);
nor U9065 (N_9065,N_8850,N_8841);
nor U9066 (N_9066,N_8555,N_8737);
and U9067 (N_9067,N_8652,N_8947);
or U9068 (N_9068,N_8699,N_8571);
or U9069 (N_9069,N_8932,N_8635);
or U9070 (N_9070,N_8601,N_8540);
nand U9071 (N_9071,N_8500,N_8919);
xnor U9072 (N_9072,N_8609,N_8593);
nand U9073 (N_9073,N_8923,N_8869);
nor U9074 (N_9074,N_8939,N_8824);
and U9075 (N_9075,N_8730,N_8503);
nor U9076 (N_9076,N_8626,N_8789);
nand U9077 (N_9077,N_8724,N_8646);
nand U9078 (N_9078,N_8672,N_8927);
nor U9079 (N_9079,N_8819,N_8657);
xor U9080 (N_9080,N_8745,N_8765);
xor U9081 (N_9081,N_8660,N_8612);
or U9082 (N_9082,N_8827,N_8760);
nand U9083 (N_9083,N_8993,N_8620);
nand U9084 (N_9084,N_8618,N_8875);
nor U9085 (N_9085,N_8666,N_8505);
and U9086 (N_9086,N_8523,N_8673);
nor U9087 (N_9087,N_8622,N_8855);
or U9088 (N_9088,N_8701,N_8961);
xor U9089 (N_9089,N_8648,N_8889);
xor U9090 (N_9090,N_8669,N_8906);
xor U9091 (N_9091,N_8656,N_8575);
nor U9092 (N_9092,N_8711,N_8835);
nor U9093 (N_9093,N_8653,N_8965);
nand U9094 (N_9094,N_8995,N_8877);
nand U9095 (N_9095,N_8574,N_8970);
nor U9096 (N_9096,N_8776,N_8983);
and U9097 (N_9097,N_8840,N_8617);
nor U9098 (N_9098,N_8920,N_8610);
xor U9099 (N_9099,N_8743,N_8596);
nor U9100 (N_9100,N_8867,N_8649);
or U9101 (N_9101,N_8502,N_8670);
and U9102 (N_9102,N_8958,N_8911);
and U9103 (N_9103,N_8704,N_8768);
nor U9104 (N_9104,N_8522,N_8832);
xnor U9105 (N_9105,N_8645,N_8944);
nor U9106 (N_9106,N_8836,N_8625);
nor U9107 (N_9107,N_8946,N_8784);
nor U9108 (N_9108,N_8676,N_8587);
or U9109 (N_9109,N_8722,N_8792);
or U9110 (N_9110,N_8973,N_8971);
and U9111 (N_9111,N_8607,N_8691);
xnor U9112 (N_9112,N_8736,N_8573);
nor U9113 (N_9113,N_8559,N_8597);
xnor U9114 (N_9114,N_8908,N_8578);
or U9115 (N_9115,N_8527,N_8529);
xnor U9116 (N_9116,N_8568,N_8520);
nor U9117 (N_9117,N_8532,N_8632);
nand U9118 (N_9118,N_8719,N_8557);
and U9119 (N_9119,N_8579,N_8738);
nand U9120 (N_9120,N_8960,N_8996);
nor U9121 (N_9121,N_8811,N_8747);
nand U9122 (N_9122,N_8543,N_8802);
and U9123 (N_9123,N_8752,N_8788);
xnor U9124 (N_9124,N_8535,N_8554);
nor U9125 (N_9125,N_8853,N_8602);
or U9126 (N_9126,N_8697,N_8703);
xnor U9127 (N_9127,N_8783,N_8812);
or U9128 (N_9128,N_8953,N_8583);
and U9129 (N_9129,N_8860,N_8880);
or U9130 (N_9130,N_8856,N_8518);
or U9131 (N_9131,N_8731,N_8615);
nand U9132 (N_9132,N_8884,N_8808);
xnor U9133 (N_9133,N_8796,N_8633);
or U9134 (N_9134,N_8943,N_8553);
nor U9135 (N_9135,N_8874,N_8748);
or U9136 (N_9136,N_8861,N_8954);
or U9137 (N_9137,N_8774,N_8948);
or U9138 (N_9138,N_8729,N_8545);
nor U9139 (N_9139,N_8909,N_8687);
xor U9140 (N_9140,N_8769,N_8664);
or U9141 (N_9141,N_8873,N_8740);
or U9142 (N_9142,N_8667,N_8829);
nor U9143 (N_9143,N_8930,N_8871);
and U9144 (N_9144,N_8689,N_8725);
or U9145 (N_9145,N_8870,N_8897);
xor U9146 (N_9146,N_8721,N_8772);
and U9147 (N_9147,N_8974,N_8825);
and U9148 (N_9148,N_8956,N_8929);
or U9149 (N_9149,N_8844,N_8549);
and U9150 (N_9150,N_8982,N_8708);
and U9151 (N_9151,N_8727,N_8780);
nor U9152 (N_9152,N_8901,N_8690);
nand U9153 (N_9153,N_8705,N_8834);
xnor U9154 (N_9154,N_8898,N_8679);
xor U9155 (N_9155,N_8933,N_8883);
or U9156 (N_9156,N_8570,N_8833);
or U9157 (N_9157,N_8950,N_8894);
nor U9158 (N_9158,N_8828,N_8581);
xor U9159 (N_9159,N_8782,N_8976);
nand U9160 (N_9160,N_8900,N_8887);
nor U9161 (N_9161,N_8680,N_8837);
nor U9162 (N_9162,N_8852,N_8755);
or U9163 (N_9163,N_8550,N_8519);
nand U9164 (N_9164,N_8878,N_8742);
xor U9165 (N_9165,N_8928,N_8773);
nor U9166 (N_9166,N_8562,N_8621);
or U9167 (N_9167,N_8524,N_8785);
nand U9168 (N_9168,N_8741,N_8600);
nand U9169 (N_9169,N_8864,N_8655);
and U9170 (N_9170,N_8634,N_8586);
and U9171 (N_9171,N_8857,N_8969);
or U9172 (N_9172,N_8799,N_8539);
nand U9173 (N_9173,N_8509,N_8845);
nor U9174 (N_9174,N_8980,N_8658);
and U9175 (N_9175,N_8952,N_8882);
and U9176 (N_9176,N_8938,N_8914);
nand U9177 (N_9177,N_8510,N_8576);
nor U9178 (N_9178,N_8826,N_8642);
nand U9179 (N_9179,N_8816,N_8754);
or U9180 (N_9180,N_8613,N_8810);
or U9181 (N_9181,N_8798,N_8542);
or U9182 (N_9182,N_8771,N_8942);
or U9183 (N_9183,N_8876,N_8848);
nand U9184 (N_9184,N_8847,N_8759);
or U9185 (N_9185,N_8681,N_8915);
nand U9186 (N_9186,N_8567,N_8558);
and U9187 (N_9187,N_8949,N_8922);
xnor U9188 (N_9188,N_8629,N_8551);
nand U9189 (N_9189,N_8733,N_8695);
and U9190 (N_9190,N_8528,N_8665);
and U9191 (N_9191,N_8989,N_8851);
nand U9192 (N_9192,N_8814,N_8945);
and U9193 (N_9193,N_8717,N_8758);
and U9194 (N_9194,N_8639,N_8916);
or U9195 (N_9195,N_8514,N_8580);
or U9196 (N_9196,N_8941,N_8892);
and U9197 (N_9197,N_8692,N_8735);
and U9198 (N_9198,N_8675,N_8507);
or U9199 (N_9199,N_8997,N_8750);
nor U9200 (N_9200,N_8720,N_8940);
nor U9201 (N_9201,N_8663,N_8547);
nor U9202 (N_9202,N_8668,N_8831);
nor U9203 (N_9203,N_8854,N_8627);
or U9204 (N_9204,N_8987,N_8988);
and U9205 (N_9205,N_8728,N_8552);
and U9206 (N_9206,N_8858,N_8951);
nand U9207 (N_9207,N_8606,N_8937);
nand U9208 (N_9208,N_8744,N_8879);
nand U9209 (N_9209,N_8588,N_8967);
nor U9210 (N_9210,N_8569,N_8817);
and U9211 (N_9211,N_8585,N_8757);
nand U9212 (N_9212,N_8712,N_8793);
and U9213 (N_9213,N_8512,N_8541);
or U9214 (N_9214,N_8896,N_8715);
nor U9215 (N_9215,N_8671,N_8696);
and U9216 (N_9216,N_8685,N_8886);
and U9217 (N_9217,N_8975,N_8815);
xnor U9218 (N_9218,N_8506,N_8565);
nor U9219 (N_9219,N_8766,N_8749);
nand U9220 (N_9220,N_8608,N_8707);
or U9221 (N_9221,N_8839,N_8761);
and U9222 (N_9222,N_8888,N_8723);
xnor U9223 (N_9223,N_8710,N_8801);
nand U9224 (N_9224,N_8795,N_8863);
xor U9225 (N_9225,N_8809,N_8662);
xor U9226 (N_9226,N_8756,N_8893);
xor U9227 (N_9227,N_8899,N_8842);
nand U9228 (N_9228,N_8548,N_8921);
or U9229 (N_9229,N_8683,N_8718);
nor U9230 (N_9230,N_8734,N_8781);
or U9231 (N_9231,N_8560,N_8732);
nor U9232 (N_9232,N_8739,N_8991);
nor U9233 (N_9233,N_8777,N_8981);
xnor U9234 (N_9234,N_8753,N_8589);
xor U9235 (N_9235,N_8511,N_8651);
and U9236 (N_9236,N_8501,N_8702);
or U9237 (N_9237,N_8767,N_8890);
or U9238 (N_9238,N_8751,N_8918);
xnor U9239 (N_9239,N_8677,N_8807);
and U9240 (N_9240,N_8859,N_8531);
nand U9241 (N_9241,N_8598,N_8604);
or U9242 (N_9242,N_8822,N_8905);
nor U9243 (N_9243,N_8536,N_8521);
nor U9244 (N_9244,N_8955,N_8972);
nand U9245 (N_9245,N_8643,N_8563);
and U9246 (N_9246,N_8963,N_8895);
nand U9247 (N_9247,N_8868,N_8925);
nand U9248 (N_9248,N_8713,N_8978);
xor U9249 (N_9249,N_8984,N_8762);
and U9250 (N_9250,N_8756,N_8878);
xnor U9251 (N_9251,N_8741,N_8618);
nor U9252 (N_9252,N_8791,N_8800);
nand U9253 (N_9253,N_8932,N_8726);
nand U9254 (N_9254,N_8755,N_8987);
or U9255 (N_9255,N_8556,N_8710);
and U9256 (N_9256,N_8875,N_8929);
or U9257 (N_9257,N_8570,N_8537);
and U9258 (N_9258,N_8608,N_8747);
nor U9259 (N_9259,N_8655,N_8687);
and U9260 (N_9260,N_8862,N_8938);
xnor U9261 (N_9261,N_8794,N_8822);
xor U9262 (N_9262,N_8985,N_8784);
and U9263 (N_9263,N_8871,N_8503);
nand U9264 (N_9264,N_8741,N_8913);
and U9265 (N_9265,N_8580,N_8530);
nor U9266 (N_9266,N_8913,N_8949);
nor U9267 (N_9267,N_8816,N_8556);
nor U9268 (N_9268,N_8980,N_8953);
nor U9269 (N_9269,N_8987,N_8968);
xor U9270 (N_9270,N_8907,N_8910);
and U9271 (N_9271,N_8553,N_8766);
nor U9272 (N_9272,N_8676,N_8842);
nor U9273 (N_9273,N_8852,N_8699);
nand U9274 (N_9274,N_8800,N_8900);
xor U9275 (N_9275,N_8530,N_8694);
and U9276 (N_9276,N_8794,N_8636);
nor U9277 (N_9277,N_8581,N_8817);
nand U9278 (N_9278,N_8672,N_8771);
nand U9279 (N_9279,N_8778,N_8812);
or U9280 (N_9280,N_8873,N_8616);
xnor U9281 (N_9281,N_8822,N_8552);
and U9282 (N_9282,N_8516,N_8826);
and U9283 (N_9283,N_8679,N_8846);
or U9284 (N_9284,N_8769,N_8576);
nand U9285 (N_9285,N_8723,N_8971);
or U9286 (N_9286,N_8504,N_8593);
and U9287 (N_9287,N_8583,N_8609);
or U9288 (N_9288,N_8621,N_8654);
xor U9289 (N_9289,N_8624,N_8773);
and U9290 (N_9290,N_8599,N_8516);
xnor U9291 (N_9291,N_8789,N_8679);
xnor U9292 (N_9292,N_8534,N_8966);
xnor U9293 (N_9293,N_8775,N_8622);
xor U9294 (N_9294,N_8645,N_8683);
xnor U9295 (N_9295,N_8989,N_8670);
xnor U9296 (N_9296,N_8691,N_8975);
or U9297 (N_9297,N_8890,N_8880);
nand U9298 (N_9298,N_8787,N_8827);
xor U9299 (N_9299,N_8589,N_8796);
and U9300 (N_9300,N_8611,N_8680);
nor U9301 (N_9301,N_8504,N_8549);
and U9302 (N_9302,N_8819,N_8794);
xor U9303 (N_9303,N_8759,N_8502);
and U9304 (N_9304,N_8640,N_8620);
nor U9305 (N_9305,N_8977,N_8954);
nor U9306 (N_9306,N_8572,N_8649);
nor U9307 (N_9307,N_8768,N_8815);
and U9308 (N_9308,N_8501,N_8885);
nand U9309 (N_9309,N_8653,N_8529);
and U9310 (N_9310,N_8979,N_8824);
nor U9311 (N_9311,N_8939,N_8876);
nor U9312 (N_9312,N_8603,N_8657);
nand U9313 (N_9313,N_8535,N_8502);
and U9314 (N_9314,N_8996,N_8855);
nor U9315 (N_9315,N_8607,N_8707);
and U9316 (N_9316,N_8762,N_8536);
nor U9317 (N_9317,N_8902,N_8940);
and U9318 (N_9318,N_8520,N_8786);
or U9319 (N_9319,N_8589,N_8516);
nand U9320 (N_9320,N_8962,N_8544);
nor U9321 (N_9321,N_8818,N_8915);
nor U9322 (N_9322,N_8628,N_8952);
or U9323 (N_9323,N_8762,N_8848);
and U9324 (N_9324,N_8544,N_8532);
and U9325 (N_9325,N_8727,N_8806);
or U9326 (N_9326,N_8815,N_8901);
nand U9327 (N_9327,N_8824,N_8928);
and U9328 (N_9328,N_8737,N_8671);
nand U9329 (N_9329,N_8817,N_8570);
nand U9330 (N_9330,N_8582,N_8525);
or U9331 (N_9331,N_8614,N_8903);
and U9332 (N_9332,N_8567,N_8694);
or U9333 (N_9333,N_8859,N_8535);
xor U9334 (N_9334,N_8509,N_8542);
nand U9335 (N_9335,N_8855,N_8892);
or U9336 (N_9336,N_8819,N_8648);
xor U9337 (N_9337,N_8765,N_8852);
xnor U9338 (N_9338,N_8634,N_8504);
or U9339 (N_9339,N_8825,N_8603);
or U9340 (N_9340,N_8769,N_8965);
nor U9341 (N_9341,N_8583,N_8929);
or U9342 (N_9342,N_8500,N_8834);
or U9343 (N_9343,N_8513,N_8827);
nor U9344 (N_9344,N_8606,N_8984);
nand U9345 (N_9345,N_8545,N_8506);
nand U9346 (N_9346,N_8896,N_8546);
and U9347 (N_9347,N_8992,N_8740);
xnor U9348 (N_9348,N_8696,N_8807);
xor U9349 (N_9349,N_8734,N_8889);
nand U9350 (N_9350,N_8733,N_8893);
xnor U9351 (N_9351,N_8854,N_8606);
xor U9352 (N_9352,N_8652,N_8500);
and U9353 (N_9353,N_8620,N_8578);
and U9354 (N_9354,N_8563,N_8738);
and U9355 (N_9355,N_8571,N_8982);
nand U9356 (N_9356,N_8646,N_8617);
or U9357 (N_9357,N_8531,N_8731);
xnor U9358 (N_9358,N_8971,N_8754);
xor U9359 (N_9359,N_8897,N_8911);
nand U9360 (N_9360,N_8846,N_8818);
or U9361 (N_9361,N_8544,N_8727);
and U9362 (N_9362,N_8621,N_8511);
and U9363 (N_9363,N_8706,N_8807);
xor U9364 (N_9364,N_8576,N_8663);
and U9365 (N_9365,N_8834,N_8594);
and U9366 (N_9366,N_8654,N_8993);
nand U9367 (N_9367,N_8650,N_8677);
nand U9368 (N_9368,N_8896,N_8921);
nand U9369 (N_9369,N_8999,N_8651);
or U9370 (N_9370,N_8797,N_8688);
nand U9371 (N_9371,N_8987,N_8585);
or U9372 (N_9372,N_8698,N_8724);
or U9373 (N_9373,N_8779,N_8553);
xor U9374 (N_9374,N_8596,N_8679);
xnor U9375 (N_9375,N_8761,N_8880);
and U9376 (N_9376,N_8911,N_8693);
and U9377 (N_9377,N_8997,N_8773);
nor U9378 (N_9378,N_8978,N_8779);
nor U9379 (N_9379,N_8962,N_8839);
or U9380 (N_9380,N_8923,N_8608);
and U9381 (N_9381,N_8979,N_8842);
or U9382 (N_9382,N_8590,N_8620);
or U9383 (N_9383,N_8726,N_8962);
or U9384 (N_9384,N_8566,N_8608);
and U9385 (N_9385,N_8671,N_8677);
and U9386 (N_9386,N_8994,N_8581);
and U9387 (N_9387,N_8818,N_8838);
nand U9388 (N_9388,N_8628,N_8524);
or U9389 (N_9389,N_8965,N_8689);
and U9390 (N_9390,N_8573,N_8975);
nand U9391 (N_9391,N_8995,N_8875);
and U9392 (N_9392,N_8936,N_8704);
xnor U9393 (N_9393,N_8751,N_8831);
and U9394 (N_9394,N_8597,N_8784);
xnor U9395 (N_9395,N_8893,N_8962);
or U9396 (N_9396,N_8793,N_8640);
and U9397 (N_9397,N_8644,N_8589);
and U9398 (N_9398,N_8799,N_8703);
or U9399 (N_9399,N_8894,N_8997);
or U9400 (N_9400,N_8654,N_8960);
and U9401 (N_9401,N_8599,N_8663);
nor U9402 (N_9402,N_8528,N_8505);
or U9403 (N_9403,N_8738,N_8862);
or U9404 (N_9404,N_8553,N_8995);
xor U9405 (N_9405,N_8543,N_8508);
nor U9406 (N_9406,N_8874,N_8782);
nor U9407 (N_9407,N_8794,N_8877);
and U9408 (N_9408,N_8575,N_8948);
and U9409 (N_9409,N_8969,N_8860);
or U9410 (N_9410,N_8714,N_8689);
and U9411 (N_9411,N_8915,N_8619);
xor U9412 (N_9412,N_8616,N_8737);
nor U9413 (N_9413,N_8708,N_8706);
and U9414 (N_9414,N_8872,N_8826);
or U9415 (N_9415,N_8600,N_8897);
nor U9416 (N_9416,N_8987,N_8933);
nor U9417 (N_9417,N_8545,N_8716);
xnor U9418 (N_9418,N_8505,N_8936);
xor U9419 (N_9419,N_8757,N_8894);
or U9420 (N_9420,N_8888,N_8502);
nand U9421 (N_9421,N_8901,N_8761);
xor U9422 (N_9422,N_8998,N_8753);
nor U9423 (N_9423,N_8577,N_8779);
and U9424 (N_9424,N_8759,N_8523);
xnor U9425 (N_9425,N_8838,N_8553);
nand U9426 (N_9426,N_8883,N_8527);
nor U9427 (N_9427,N_8602,N_8729);
nor U9428 (N_9428,N_8909,N_8608);
and U9429 (N_9429,N_8535,N_8523);
xor U9430 (N_9430,N_8694,N_8809);
and U9431 (N_9431,N_8510,N_8627);
nor U9432 (N_9432,N_8721,N_8870);
nand U9433 (N_9433,N_8808,N_8583);
or U9434 (N_9434,N_8557,N_8760);
nor U9435 (N_9435,N_8735,N_8970);
nand U9436 (N_9436,N_8514,N_8826);
or U9437 (N_9437,N_8810,N_8777);
or U9438 (N_9438,N_8942,N_8637);
nor U9439 (N_9439,N_8500,N_8936);
nand U9440 (N_9440,N_8856,N_8542);
nand U9441 (N_9441,N_8545,N_8649);
or U9442 (N_9442,N_8521,N_8792);
or U9443 (N_9443,N_8989,N_8788);
nand U9444 (N_9444,N_8925,N_8939);
nor U9445 (N_9445,N_8786,N_8617);
xor U9446 (N_9446,N_8591,N_8585);
and U9447 (N_9447,N_8609,N_8544);
nor U9448 (N_9448,N_8881,N_8982);
and U9449 (N_9449,N_8776,N_8960);
nor U9450 (N_9450,N_8961,N_8785);
xnor U9451 (N_9451,N_8913,N_8878);
nor U9452 (N_9452,N_8531,N_8943);
nand U9453 (N_9453,N_8680,N_8565);
nor U9454 (N_9454,N_8930,N_8545);
xor U9455 (N_9455,N_8756,N_8506);
nor U9456 (N_9456,N_8700,N_8723);
or U9457 (N_9457,N_8548,N_8506);
xnor U9458 (N_9458,N_8744,N_8956);
xnor U9459 (N_9459,N_8693,N_8757);
or U9460 (N_9460,N_8838,N_8923);
xor U9461 (N_9461,N_8801,N_8939);
nand U9462 (N_9462,N_8758,N_8970);
nand U9463 (N_9463,N_8986,N_8514);
and U9464 (N_9464,N_8557,N_8978);
nor U9465 (N_9465,N_8872,N_8614);
xnor U9466 (N_9466,N_8951,N_8940);
xor U9467 (N_9467,N_8659,N_8930);
and U9468 (N_9468,N_8573,N_8621);
and U9469 (N_9469,N_8632,N_8824);
xnor U9470 (N_9470,N_8975,N_8649);
xor U9471 (N_9471,N_8589,N_8743);
and U9472 (N_9472,N_8929,N_8777);
xor U9473 (N_9473,N_8568,N_8863);
nor U9474 (N_9474,N_8805,N_8625);
and U9475 (N_9475,N_8955,N_8918);
nand U9476 (N_9476,N_8774,N_8557);
and U9477 (N_9477,N_8535,N_8669);
and U9478 (N_9478,N_8875,N_8860);
nand U9479 (N_9479,N_8571,N_8776);
nand U9480 (N_9480,N_8549,N_8769);
or U9481 (N_9481,N_8744,N_8814);
nor U9482 (N_9482,N_8837,N_8640);
xor U9483 (N_9483,N_8640,N_8838);
and U9484 (N_9484,N_8940,N_8726);
and U9485 (N_9485,N_8848,N_8522);
or U9486 (N_9486,N_8798,N_8644);
and U9487 (N_9487,N_8999,N_8717);
xnor U9488 (N_9488,N_8582,N_8859);
xnor U9489 (N_9489,N_8608,N_8945);
nor U9490 (N_9490,N_8868,N_8639);
nor U9491 (N_9491,N_8974,N_8706);
nand U9492 (N_9492,N_8791,N_8875);
nor U9493 (N_9493,N_8754,N_8804);
and U9494 (N_9494,N_8711,N_8936);
nand U9495 (N_9495,N_8948,N_8875);
or U9496 (N_9496,N_8794,N_8779);
xnor U9497 (N_9497,N_8628,N_8724);
nor U9498 (N_9498,N_8759,N_8903);
nor U9499 (N_9499,N_8547,N_8549);
xnor U9500 (N_9500,N_9054,N_9246);
nand U9501 (N_9501,N_9446,N_9236);
xor U9502 (N_9502,N_9448,N_9279);
nor U9503 (N_9503,N_9186,N_9007);
xor U9504 (N_9504,N_9076,N_9103);
nand U9505 (N_9505,N_9419,N_9318);
nor U9506 (N_9506,N_9127,N_9343);
and U9507 (N_9507,N_9220,N_9250);
and U9508 (N_9508,N_9276,N_9474);
nor U9509 (N_9509,N_9301,N_9353);
nand U9510 (N_9510,N_9471,N_9026);
nor U9511 (N_9511,N_9036,N_9041);
xor U9512 (N_9512,N_9392,N_9191);
nor U9513 (N_9513,N_9348,N_9135);
and U9514 (N_9514,N_9452,N_9477);
nor U9515 (N_9515,N_9299,N_9153);
and U9516 (N_9516,N_9057,N_9126);
nand U9517 (N_9517,N_9045,N_9199);
xnor U9518 (N_9518,N_9174,N_9238);
or U9519 (N_9519,N_9274,N_9495);
xnor U9520 (N_9520,N_9275,N_9244);
nor U9521 (N_9521,N_9034,N_9481);
nor U9522 (N_9522,N_9398,N_9366);
nand U9523 (N_9523,N_9150,N_9214);
or U9524 (N_9524,N_9418,N_9483);
nand U9525 (N_9525,N_9050,N_9493);
or U9526 (N_9526,N_9308,N_9297);
xnor U9527 (N_9527,N_9396,N_9202);
or U9528 (N_9528,N_9109,N_9394);
xor U9529 (N_9529,N_9372,N_9125);
or U9530 (N_9530,N_9385,N_9027);
nand U9531 (N_9531,N_9256,N_9155);
nor U9532 (N_9532,N_9283,N_9375);
nor U9533 (N_9533,N_9435,N_9384);
or U9534 (N_9534,N_9380,N_9492);
and U9535 (N_9535,N_9140,N_9075);
nand U9536 (N_9536,N_9273,N_9223);
or U9537 (N_9537,N_9179,N_9387);
xnor U9538 (N_9538,N_9367,N_9429);
or U9539 (N_9539,N_9200,N_9347);
and U9540 (N_9540,N_9205,N_9116);
xnor U9541 (N_9541,N_9403,N_9177);
xor U9542 (N_9542,N_9431,N_9123);
nand U9543 (N_9543,N_9413,N_9369);
and U9544 (N_9544,N_9132,N_9120);
xnor U9545 (N_9545,N_9163,N_9440);
or U9546 (N_9546,N_9156,N_9022);
xnor U9547 (N_9547,N_9356,N_9194);
nand U9548 (N_9548,N_9263,N_9342);
xor U9549 (N_9549,N_9059,N_9016);
and U9550 (N_9550,N_9300,N_9410);
nor U9551 (N_9551,N_9290,N_9173);
nand U9552 (N_9552,N_9455,N_9399);
or U9553 (N_9553,N_9241,N_9104);
nor U9554 (N_9554,N_9305,N_9011);
nand U9555 (N_9555,N_9061,N_9361);
nand U9556 (N_9556,N_9249,N_9000);
nor U9557 (N_9557,N_9428,N_9306);
nand U9558 (N_9558,N_9425,N_9260);
and U9559 (N_9559,N_9043,N_9340);
xnor U9560 (N_9560,N_9024,N_9251);
xor U9561 (N_9561,N_9234,N_9439);
or U9562 (N_9562,N_9469,N_9136);
xnor U9563 (N_9563,N_9409,N_9258);
xor U9564 (N_9564,N_9467,N_9110);
and U9565 (N_9565,N_9459,N_9006);
nor U9566 (N_9566,N_9063,N_9437);
or U9567 (N_9567,N_9229,N_9151);
and U9568 (N_9568,N_9257,N_9119);
and U9569 (N_9569,N_9154,N_9188);
nor U9570 (N_9570,N_9096,N_9037);
and U9571 (N_9571,N_9230,N_9423);
and U9572 (N_9572,N_9389,N_9111);
xor U9573 (N_9573,N_9053,N_9030);
nor U9574 (N_9574,N_9331,N_9021);
nand U9575 (N_9575,N_9039,N_9082);
or U9576 (N_9576,N_9064,N_9161);
and U9577 (N_9577,N_9268,N_9292);
or U9578 (N_9578,N_9081,N_9303);
xnor U9579 (N_9579,N_9206,N_9350);
and U9580 (N_9580,N_9192,N_9001);
and U9581 (N_9581,N_9470,N_9355);
or U9582 (N_9582,N_9204,N_9227);
and U9583 (N_9583,N_9298,N_9121);
and U9584 (N_9584,N_9092,N_9464);
nand U9585 (N_9585,N_9134,N_9231);
and U9586 (N_9586,N_9487,N_9073);
xor U9587 (N_9587,N_9383,N_9406);
nor U9588 (N_9588,N_9371,N_9052);
or U9589 (N_9589,N_9145,N_9089);
and U9590 (N_9590,N_9472,N_9216);
or U9591 (N_9591,N_9334,N_9449);
xor U9592 (N_9592,N_9479,N_9405);
or U9593 (N_9593,N_9040,N_9072);
or U9594 (N_9594,N_9408,N_9046);
or U9595 (N_9595,N_9243,N_9093);
xnor U9596 (N_9596,N_9203,N_9014);
or U9597 (N_9597,N_9322,N_9259);
or U9598 (N_9598,N_9391,N_9166);
xor U9599 (N_9599,N_9208,N_9284);
and U9600 (N_9600,N_9232,N_9210);
nand U9601 (N_9601,N_9265,N_9165);
xor U9602 (N_9602,N_9183,N_9363);
or U9603 (N_9603,N_9222,N_9182);
and U9604 (N_9604,N_9071,N_9098);
or U9605 (N_9605,N_9485,N_9262);
nand U9606 (N_9606,N_9176,N_9484);
or U9607 (N_9607,N_9444,N_9038);
and U9608 (N_9608,N_9476,N_9247);
nand U9609 (N_9609,N_9003,N_9328);
nand U9610 (N_9610,N_9456,N_9441);
nor U9611 (N_9611,N_9108,N_9240);
and U9612 (N_9612,N_9196,N_9271);
xor U9613 (N_9613,N_9058,N_9160);
or U9614 (N_9614,N_9253,N_9360);
or U9615 (N_9615,N_9304,N_9048);
nand U9616 (N_9616,N_9146,N_9281);
or U9617 (N_9617,N_9379,N_9242);
or U9618 (N_9618,N_9499,N_9029);
or U9619 (N_9619,N_9087,N_9143);
xnor U9620 (N_9620,N_9115,N_9008);
nand U9621 (N_9621,N_9338,N_9184);
and U9622 (N_9622,N_9175,N_9218);
and U9623 (N_9623,N_9417,N_9002);
nor U9624 (N_9624,N_9323,N_9377);
and U9625 (N_9625,N_9239,N_9497);
and U9626 (N_9626,N_9368,N_9460);
nand U9627 (N_9627,N_9498,N_9131);
xor U9628 (N_9628,N_9287,N_9224);
nand U9629 (N_9629,N_9023,N_9374);
nor U9630 (N_9630,N_9434,N_9051);
nand U9631 (N_9631,N_9412,N_9211);
nor U9632 (N_9632,N_9349,N_9101);
and U9633 (N_9633,N_9212,N_9312);
nand U9634 (N_9634,N_9294,N_9221);
and U9635 (N_9635,N_9404,N_9067);
nor U9636 (N_9636,N_9245,N_9461);
xnor U9637 (N_9637,N_9422,N_9285);
nand U9638 (N_9638,N_9463,N_9482);
nand U9639 (N_9639,N_9069,N_9209);
nor U9640 (N_9640,N_9124,N_9376);
xnor U9641 (N_9641,N_9009,N_9272);
nor U9642 (N_9642,N_9167,N_9139);
nor U9643 (N_9643,N_9373,N_9468);
nand U9644 (N_9644,N_9074,N_9491);
nand U9645 (N_9645,N_9102,N_9226);
nor U9646 (N_9646,N_9118,N_9085);
nand U9647 (N_9647,N_9317,N_9270);
or U9648 (N_9648,N_9443,N_9195);
nor U9649 (N_9649,N_9364,N_9496);
and U9650 (N_9650,N_9099,N_9266);
and U9651 (N_9651,N_9321,N_9237);
or U9652 (N_9652,N_9277,N_9433);
and U9653 (N_9653,N_9316,N_9062);
and U9654 (N_9654,N_9033,N_9445);
nand U9655 (N_9655,N_9390,N_9187);
xor U9656 (N_9656,N_9269,N_9019);
and U9657 (N_9657,N_9295,N_9083);
nor U9658 (N_9658,N_9382,N_9447);
or U9659 (N_9659,N_9086,N_9055);
or U9660 (N_9660,N_9314,N_9480);
nand U9661 (N_9661,N_9193,N_9381);
nand U9662 (N_9662,N_9010,N_9351);
nand U9663 (N_9663,N_9473,N_9138);
nand U9664 (N_9664,N_9032,N_9235);
nor U9665 (N_9665,N_9329,N_9286);
xor U9666 (N_9666,N_9130,N_9152);
nand U9667 (N_9667,N_9198,N_9133);
and U9668 (N_9668,N_9171,N_9293);
nand U9669 (N_9669,N_9261,N_9311);
or U9670 (N_9670,N_9004,N_9420);
nand U9671 (N_9671,N_9401,N_9219);
xor U9672 (N_9672,N_9201,N_9185);
xor U9673 (N_9673,N_9147,N_9105);
nor U9674 (N_9674,N_9025,N_9189);
or U9675 (N_9675,N_9432,N_9325);
nand U9676 (N_9676,N_9065,N_9013);
xor U9677 (N_9677,N_9370,N_9042);
nand U9678 (N_9678,N_9309,N_9319);
and U9679 (N_9679,N_9289,N_9264);
nand U9680 (N_9680,N_9352,N_9088);
and U9681 (N_9681,N_9158,N_9337);
and U9682 (N_9682,N_9346,N_9397);
and U9683 (N_9683,N_9015,N_9068);
nor U9684 (N_9684,N_9386,N_9020);
nand U9685 (N_9685,N_9159,N_9248);
and U9686 (N_9686,N_9017,N_9144);
and U9687 (N_9687,N_9056,N_9291);
xnor U9688 (N_9688,N_9333,N_9066);
xnor U9689 (N_9689,N_9424,N_9097);
nor U9690 (N_9690,N_9453,N_9117);
or U9691 (N_9691,N_9326,N_9078);
nor U9692 (N_9692,N_9426,N_9378);
xnor U9693 (N_9693,N_9012,N_9458);
or U9694 (N_9694,N_9114,N_9267);
and U9695 (N_9695,N_9466,N_9489);
or U9696 (N_9696,N_9047,N_9451);
nor U9697 (N_9697,N_9336,N_9148);
or U9698 (N_9698,N_9169,N_9207);
and U9699 (N_9699,N_9213,N_9197);
xnor U9700 (N_9700,N_9107,N_9462);
xnor U9701 (N_9701,N_9049,N_9044);
and U9702 (N_9702,N_9427,N_9307);
xnor U9703 (N_9703,N_9157,N_9180);
nand U9704 (N_9704,N_9494,N_9341);
nand U9705 (N_9705,N_9129,N_9320);
nor U9706 (N_9706,N_9407,N_9090);
nor U9707 (N_9707,N_9288,N_9415);
xor U9708 (N_9708,N_9091,N_9488);
and U9709 (N_9709,N_9280,N_9028);
and U9710 (N_9710,N_9365,N_9490);
nor U9711 (N_9711,N_9168,N_9438);
nand U9712 (N_9712,N_9411,N_9100);
or U9713 (N_9713,N_9457,N_9388);
and U9714 (N_9714,N_9079,N_9310);
nor U9715 (N_9715,N_9475,N_9122);
nor U9716 (N_9716,N_9345,N_9486);
nor U9717 (N_9717,N_9077,N_9454);
nor U9718 (N_9718,N_9255,N_9181);
or U9719 (N_9719,N_9302,N_9225);
nand U9720 (N_9720,N_9170,N_9339);
or U9721 (N_9721,N_9142,N_9402);
nand U9722 (N_9722,N_9335,N_9436);
nor U9723 (N_9723,N_9416,N_9358);
nor U9724 (N_9724,N_9282,N_9296);
and U9725 (N_9725,N_9113,N_9094);
nand U9726 (N_9726,N_9313,N_9106);
and U9727 (N_9727,N_9031,N_9395);
or U9728 (N_9728,N_9450,N_9095);
or U9729 (N_9729,N_9344,N_9162);
or U9730 (N_9730,N_9215,N_9362);
nor U9731 (N_9731,N_9330,N_9332);
nor U9732 (N_9732,N_9278,N_9252);
or U9733 (N_9733,N_9400,N_9359);
xor U9734 (N_9734,N_9112,N_9233);
xnor U9735 (N_9735,N_9018,N_9164);
xor U9736 (N_9736,N_9430,N_9254);
and U9737 (N_9737,N_9190,N_9357);
or U9738 (N_9738,N_9217,N_9414);
nand U9739 (N_9739,N_9478,N_9324);
or U9740 (N_9740,N_9315,N_9228);
and U9741 (N_9741,N_9060,N_9141);
or U9742 (N_9742,N_9421,N_9128);
or U9743 (N_9743,N_9172,N_9178);
nor U9744 (N_9744,N_9080,N_9035);
xor U9745 (N_9745,N_9393,N_9005);
nand U9746 (N_9746,N_9442,N_9070);
nor U9747 (N_9747,N_9149,N_9354);
xnor U9748 (N_9748,N_9465,N_9084);
nand U9749 (N_9749,N_9327,N_9137);
nand U9750 (N_9750,N_9435,N_9468);
nor U9751 (N_9751,N_9199,N_9077);
and U9752 (N_9752,N_9290,N_9048);
and U9753 (N_9753,N_9413,N_9184);
nand U9754 (N_9754,N_9272,N_9106);
nand U9755 (N_9755,N_9144,N_9125);
nand U9756 (N_9756,N_9162,N_9327);
and U9757 (N_9757,N_9290,N_9480);
nor U9758 (N_9758,N_9274,N_9209);
or U9759 (N_9759,N_9295,N_9355);
nand U9760 (N_9760,N_9108,N_9415);
nor U9761 (N_9761,N_9351,N_9318);
nor U9762 (N_9762,N_9051,N_9281);
and U9763 (N_9763,N_9257,N_9085);
and U9764 (N_9764,N_9366,N_9247);
xnor U9765 (N_9765,N_9278,N_9160);
nor U9766 (N_9766,N_9077,N_9097);
nand U9767 (N_9767,N_9335,N_9222);
nand U9768 (N_9768,N_9048,N_9237);
and U9769 (N_9769,N_9490,N_9321);
nand U9770 (N_9770,N_9352,N_9295);
and U9771 (N_9771,N_9064,N_9381);
nor U9772 (N_9772,N_9152,N_9343);
nand U9773 (N_9773,N_9084,N_9207);
nor U9774 (N_9774,N_9178,N_9166);
nand U9775 (N_9775,N_9361,N_9327);
or U9776 (N_9776,N_9179,N_9290);
nand U9777 (N_9777,N_9307,N_9333);
and U9778 (N_9778,N_9397,N_9461);
and U9779 (N_9779,N_9223,N_9161);
nand U9780 (N_9780,N_9298,N_9328);
nor U9781 (N_9781,N_9341,N_9120);
xnor U9782 (N_9782,N_9335,N_9307);
and U9783 (N_9783,N_9320,N_9312);
and U9784 (N_9784,N_9260,N_9314);
or U9785 (N_9785,N_9181,N_9236);
or U9786 (N_9786,N_9101,N_9437);
nand U9787 (N_9787,N_9002,N_9411);
nor U9788 (N_9788,N_9056,N_9282);
nand U9789 (N_9789,N_9382,N_9359);
or U9790 (N_9790,N_9215,N_9272);
xor U9791 (N_9791,N_9063,N_9271);
or U9792 (N_9792,N_9012,N_9181);
nor U9793 (N_9793,N_9191,N_9304);
nor U9794 (N_9794,N_9181,N_9049);
nor U9795 (N_9795,N_9022,N_9274);
nor U9796 (N_9796,N_9302,N_9233);
xor U9797 (N_9797,N_9018,N_9225);
nor U9798 (N_9798,N_9315,N_9312);
or U9799 (N_9799,N_9451,N_9303);
nand U9800 (N_9800,N_9466,N_9210);
and U9801 (N_9801,N_9456,N_9339);
and U9802 (N_9802,N_9367,N_9241);
xor U9803 (N_9803,N_9308,N_9435);
xnor U9804 (N_9804,N_9386,N_9397);
nand U9805 (N_9805,N_9235,N_9355);
or U9806 (N_9806,N_9094,N_9290);
or U9807 (N_9807,N_9163,N_9355);
and U9808 (N_9808,N_9073,N_9388);
and U9809 (N_9809,N_9289,N_9303);
or U9810 (N_9810,N_9120,N_9333);
nor U9811 (N_9811,N_9273,N_9338);
and U9812 (N_9812,N_9157,N_9249);
and U9813 (N_9813,N_9213,N_9499);
or U9814 (N_9814,N_9376,N_9248);
and U9815 (N_9815,N_9113,N_9219);
nand U9816 (N_9816,N_9106,N_9343);
xnor U9817 (N_9817,N_9195,N_9077);
nor U9818 (N_9818,N_9289,N_9075);
nand U9819 (N_9819,N_9256,N_9230);
or U9820 (N_9820,N_9001,N_9127);
and U9821 (N_9821,N_9115,N_9458);
nor U9822 (N_9822,N_9011,N_9343);
xnor U9823 (N_9823,N_9262,N_9125);
nor U9824 (N_9824,N_9162,N_9155);
or U9825 (N_9825,N_9466,N_9457);
nor U9826 (N_9826,N_9367,N_9326);
and U9827 (N_9827,N_9103,N_9131);
xor U9828 (N_9828,N_9325,N_9317);
nand U9829 (N_9829,N_9346,N_9327);
nor U9830 (N_9830,N_9115,N_9045);
nor U9831 (N_9831,N_9308,N_9065);
nand U9832 (N_9832,N_9234,N_9426);
nand U9833 (N_9833,N_9071,N_9312);
or U9834 (N_9834,N_9258,N_9400);
and U9835 (N_9835,N_9274,N_9275);
and U9836 (N_9836,N_9266,N_9459);
nor U9837 (N_9837,N_9187,N_9037);
or U9838 (N_9838,N_9495,N_9124);
or U9839 (N_9839,N_9092,N_9018);
nand U9840 (N_9840,N_9348,N_9076);
nor U9841 (N_9841,N_9378,N_9185);
nand U9842 (N_9842,N_9409,N_9160);
nand U9843 (N_9843,N_9281,N_9222);
or U9844 (N_9844,N_9006,N_9316);
xnor U9845 (N_9845,N_9075,N_9373);
nand U9846 (N_9846,N_9375,N_9213);
or U9847 (N_9847,N_9374,N_9437);
nand U9848 (N_9848,N_9183,N_9466);
and U9849 (N_9849,N_9156,N_9208);
and U9850 (N_9850,N_9322,N_9173);
nand U9851 (N_9851,N_9174,N_9425);
nand U9852 (N_9852,N_9186,N_9432);
nor U9853 (N_9853,N_9284,N_9224);
or U9854 (N_9854,N_9314,N_9377);
nor U9855 (N_9855,N_9122,N_9278);
nor U9856 (N_9856,N_9440,N_9210);
nor U9857 (N_9857,N_9356,N_9146);
or U9858 (N_9858,N_9335,N_9011);
nor U9859 (N_9859,N_9198,N_9467);
or U9860 (N_9860,N_9407,N_9368);
and U9861 (N_9861,N_9235,N_9095);
and U9862 (N_9862,N_9189,N_9470);
or U9863 (N_9863,N_9074,N_9043);
or U9864 (N_9864,N_9018,N_9171);
and U9865 (N_9865,N_9428,N_9051);
and U9866 (N_9866,N_9201,N_9306);
nor U9867 (N_9867,N_9407,N_9371);
or U9868 (N_9868,N_9147,N_9486);
xnor U9869 (N_9869,N_9374,N_9227);
and U9870 (N_9870,N_9010,N_9148);
xor U9871 (N_9871,N_9277,N_9142);
nand U9872 (N_9872,N_9337,N_9304);
and U9873 (N_9873,N_9124,N_9451);
and U9874 (N_9874,N_9087,N_9006);
nand U9875 (N_9875,N_9059,N_9117);
nor U9876 (N_9876,N_9453,N_9186);
and U9877 (N_9877,N_9458,N_9384);
nand U9878 (N_9878,N_9302,N_9310);
nor U9879 (N_9879,N_9246,N_9254);
xnor U9880 (N_9880,N_9221,N_9441);
nand U9881 (N_9881,N_9018,N_9404);
xnor U9882 (N_9882,N_9252,N_9076);
or U9883 (N_9883,N_9057,N_9184);
nand U9884 (N_9884,N_9268,N_9322);
nor U9885 (N_9885,N_9098,N_9276);
or U9886 (N_9886,N_9476,N_9166);
or U9887 (N_9887,N_9109,N_9371);
xnor U9888 (N_9888,N_9431,N_9299);
or U9889 (N_9889,N_9093,N_9270);
or U9890 (N_9890,N_9166,N_9165);
and U9891 (N_9891,N_9402,N_9306);
and U9892 (N_9892,N_9224,N_9197);
xnor U9893 (N_9893,N_9013,N_9315);
nor U9894 (N_9894,N_9312,N_9133);
or U9895 (N_9895,N_9316,N_9288);
xor U9896 (N_9896,N_9472,N_9253);
nand U9897 (N_9897,N_9489,N_9371);
nand U9898 (N_9898,N_9363,N_9165);
nor U9899 (N_9899,N_9441,N_9377);
or U9900 (N_9900,N_9184,N_9472);
nand U9901 (N_9901,N_9414,N_9331);
nor U9902 (N_9902,N_9084,N_9037);
or U9903 (N_9903,N_9187,N_9391);
and U9904 (N_9904,N_9026,N_9453);
xnor U9905 (N_9905,N_9248,N_9216);
xnor U9906 (N_9906,N_9306,N_9336);
or U9907 (N_9907,N_9309,N_9249);
or U9908 (N_9908,N_9342,N_9128);
or U9909 (N_9909,N_9263,N_9151);
nor U9910 (N_9910,N_9064,N_9451);
xor U9911 (N_9911,N_9003,N_9172);
nand U9912 (N_9912,N_9468,N_9131);
or U9913 (N_9913,N_9458,N_9179);
nand U9914 (N_9914,N_9259,N_9056);
nand U9915 (N_9915,N_9116,N_9446);
and U9916 (N_9916,N_9063,N_9126);
nand U9917 (N_9917,N_9022,N_9251);
or U9918 (N_9918,N_9465,N_9118);
nor U9919 (N_9919,N_9434,N_9308);
or U9920 (N_9920,N_9062,N_9325);
or U9921 (N_9921,N_9039,N_9106);
nand U9922 (N_9922,N_9497,N_9443);
nand U9923 (N_9923,N_9182,N_9392);
or U9924 (N_9924,N_9424,N_9409);
or U9925 (N_9925,N_9149,N_9029);
nand U9926 (N_9926,N_9362,N_9481);
nand U9927 (N_9927,N_9452,N_9290);
xor U9928 (N_9928,N_9430,N_9472);
nor U9929 (N_9929,N_9063,N_9173);
nor U9930 (N_9930,N_9396,N_9226);
nor U9931 (N_9931,N_9209,N_9020);
or U9932 (N_9932,N_9247,N_9171);
xnor U9933 (N_9933,N_9340,N_9476);
nand U9934 (N_9934,N_9398,N_9129);
nor U9935 (N_9935,N_9336,N_9440);
nand U9936 (N_9936,N_9334,N_9244);
nor U9937 (N_9937,N_9399,N_9159);
and U9938 (N_9938,N_9096,N_9102);
or U9939 (N_9939,N_9094,N_9324);
xnor U9940 (N_9940,N_9422,N_9205);
nand U9941 (N_9941,N_9073,N_9392);
nand U9942 (N_9942,N_9096,N_9373);
or U9943 (N_9943,N_9155,N_9482);
or U9944 (N_9944,N_9416,N_9164);
nand U9945 (N_9945,N_9251,N_9093);
nand U9946 (N_9946,N_9232,N_9096);
and U9947 (N_9947,N_9443,N_9423);
nor U9948 (N_9948,N_9172,N_9050);
and U9949 (N_9949,N_9157,N_9310);
nor U9950 (N_9950,N_9261,N_9304);
xor U9951 (N_9951,N_9320,N_9059);
xor U9952 (N_9952,N_9285,N_9274);
and U9953 (N_9953,N_9155,N_9176);
or U9954 (N_9954,N_9143,N_9270);
or U9955 (N_9955,N_9378,N_9473);
or U9956 (N_9956,N_9222,N_9073);
nor U9957 (N_9957,N_9447,N_9469);
or U9958 (N_9958,N_9474,N_9493);
nor U9959 (N_9959,N_9374,N_9243);
xor U9960 (N_9960,N_9478,N_9187);
xor U9961 (N_9961,N_9301,N_9166);
xnor U9962 (N_9962,N_9435,N_9333);
xor U9963 (N_9963,N_9121,N_9273);
or U9964 (N_9964,N_9380,N_9469);
nand U9965 (N_9965,N_9369,N_9325);
nor U9966 (N_9966,N_9197,N_9066);
nand U9967 (N_9967,N_9354,N_9445);
or U9968 (N_9968,N_9112,N_9212);
nand U9969 (N_9969,N_9074,N_9203);
nand U9970 (N_9970,N_9058,N_9386);
xnor U9971 (N_9971,N_9495,N_9169);
nand U9972 (N_9972,N_9173,N_9340);
xor U9973 (N_9973,N_9257,N_9456);
and U9974 (N_9974,N_9064,N_9048);
nor U9975 (N_9975,N_9102,N_9051);
or U9976 (N_9976,N_9388,N_9434);
or U9977 (N_9977,N_9458,N_9371);
or U9978 (N_9978,N_9085,N_9100);
or U9979 (N_9979,N_9139,N_9341);
nor U9980 (N_9980,N_9106,N_9056);
xnor U9981 (N_9981,N_9476,N_9379);
xnor U9982 (N_9982,N_9421,N_9069);
nand U9983 (N_9983,N_9052,N_9047);
nand U9984 (N_9984,N_9100,N_9277);
or U9985 (N_9985,N_9486,N_9475);
xor U9986 (N_9986,N_9228,N_9160);
xnor U9987 (N_9987,N_9198,N_9007);
nand U9988 (N_9988,N_9389,N_9357);
xor U9989 (N_9989,N_9415,N_9065);
and U9990 (N_9990,N_9308,N_9244);
or U9991 (N_9991,N_9061,N_9311);
nor U9992 (N_9992,N_9238,N_9066);
or U9993 (N_9993,N_9383,N_9169);
and U9994 (N_9994,N_9082,N_9125);
xor U9995 (N_9995,N_9288,N_9462);
and U9996 (N_9996,N_9352,N_9196);
or U9997 (N_9997,N_9006,N_9115);
or U9998 (N_9998,N_9236,N_9143);
or U9999 (N_9999,N_9258,N_9072);
or U10000 (N_10000,N_9718,N_9581);
nand U10001 (N_10001,N_9604,N_9828);
nand U10002 (N_10002,N_9606,N_9960);
or U10003 (N_10003,N_9788,N_9862);
nor U10004 (N_10004,N_9775,N_9845);
xnor U10005 (N_10005,N_9638,N_9934);
nor U10006 (N_10006,N_9946,N_9688);
nand U10007 (N_10007,N_9897,N_9774);
nand U10008 (N_10008,N_9745,N_9961);
or U10009 (N_10009,N_9559,N_9735);
and U10010 (N_10010,N_9628,N_9858);
and U10011 (N_10011,N_9590,N_9920);
nor U10012 (N_10012,N_9928,N_9723);
nand U10013 (N_10013,N_9556,N_9754);
and U10014 (N_10014,N_9864,N_9511);
nor U10015 (N_10015,N_9903,N_9986);
nor U10016 (N_10016,N_9943,N_9913);
or U10017 (N_10017,N_9938,N_9531);
and U10018 (N_10018,N_9616,N_9999);
xnor U10019 (N_10019,N_9551,N_9653);
and U10020 (N_10020,N_9572,N_9975);
and U10021 (N_10021,N_9921,N_9573);
nor U10022 (N_10022,N_9620,N_9841);
xnor U10023 (N_10023,N_9996,N_9524);
or U10024 (N_10024,N_9885,N_9831);
xor U10025 (N_10025,N_9984,N_9500);
nor U10026 (N_10026,N_9945,N_9583);
xor U10027 (N_10027,N_9591,N_9839);
xnor U10028 (N_10028,N_9801,N_9981);
or U10029 (N_10029,N_9566,N_9567);
and U10030 (N_10030,N_9576,N_9546);
xnor U10031 (N_10031,N_9923,N_9682);
nand U10032 (N_10032,N_9674,N_9692);
or U10033 (N_10033,N_9679,N_9689);
and U10034 (N_10034,N_9894,N_9976);
or U10035 (N_10035,N_9748,N_9643);
nand U10036 (N_10036,N_9677,N_9635);
nand U10037 (N_10037,N_9870,N_9891);
and U10038 (N_10038,N_9985,N_9770);
or U10039 (N_10039,N_9633,N_9807);
or U10040 (N_10040,N_9800,N_9790);
or U10041 (N_10041,N_9697,N_9716);
nor U10042 (N_10042,N_9826,N_9869);
and U10043 (N_10043,N_9930,N_9969);
nand U10044 (N_10044,N_9545,N_9597);
nor U10045 (N_10045,N_9860,N_9505);
nand U10046 (N_10046,N_9655,N_9552);
xor U10047 (N_10047,N_9872,N_9530);
and U10048 (N_10048,N_9783,N_9816);
xnor U10049 (N_10049,N_9776,N_9974);
nor U10050 (N_10050,N_9519,N_9699);
nand U10051 (N_10051,N_9773,N_9861);
and U10052 (N_10052,N_9721,N_9792);
nand U10053 (N_10053,N_9678,N_9970);
xor U10054 (N_10054,N_9939,N_9892);
xnor U10055 (N_10055,N_9514,N_9710);
nor U10056 (N_10056,N_9998,N_9611);
and U10057 (N_10057,N_9520,N_9602);
or U10058 (N_10058,N_9877,N_9762);
or U10059 (N_10059,N_9899,N_9886);
or U10060 (N_10060,N_9512,N_9694);
nand U10061 (N_10061,N_9854,N_9925);
or U10062 (N_10062,N_9900,N_9501);
xnor U10063 (N_10063,N_9742,N_9997);
xnor U10064 (N_10064,N_9702,N_9879);
or U10065 (N_10065,N_9508,N_9901);
or U10066 (N_10066,N_9931,N_9905);
and U10067 (N_10067,N_9914,N_9673);
nor U10068 (N_10068,N_9561,N_9593);
nand U10069 (N_10069,N_9560,N_9589);
nor U10070 (N_10070,N_9663,N_9875);
and U10071 (N_10071,N_9607,N_9781);
xnor U10072 (N_10072,N_9982,N_9918);
nand U10073 (N_10073,N_9952,N_9936);
and U10074 (N_10074,N_9506,N_9640);
xor U10075 (N_10075,N_9672,N_9850);
nand U10076 (N_10076,N_9786,N_9648);
nor U10077 (N_10077,N_9764,N_9851);
nor U10078 (N_10078,N_9769,N_9907);
nor U10079 (N_10079,N_9932,N_9812);
xor U10080 (N_10080,N_9765,N_9883);
and U10081 (N_10081,N_9782,N_9987);
or U10082 (N_10082,N_9726,N_9634);
or U10083 (N_10083,N_9779,N_9789);
nor U10084 (N_10084,N_9941,N_9804);
nor U10085 (N_10085,N_9691,N_9594);
or U10086 (N_10086,N_9617,N_9915);
nor U10087 (N_10087,N_9637,N_9836);
nor U10088 (N_10088,N_9950,N_9859);
xnor U10089 (N_10089,N_9881,N_9740);
nor U10090 (N_10090,N_9784,N_9584);
or U10091 (N_10091,N_9761,N_9542);
and U10092 (N_10092,N_9728,N_9507);
nor U10093 (N_10093,N_9738,N_9618);
xnor U10094 (N_10094,N_9980,N_9675);
and U10095 (N_10095,N_9805,N_9629);
or U10096 (N_10096,N_9527,N_9878);
xnor U10097 (N_10097,N_9821,N_9563);
or U10098 (N_10098,N_9568,N_9731);
or U10099 (N_10099,N_9739,N_9825);
nand U10100 (N_10100,N_9808,N_9562);
nand U10101 (N_10101,N_9684,N_9598);
nand U10102 (N_10102,N_9971,N_9513);
and U10103 (N_10103,N_9570,N_9955);
and U10104 (N_10104,N_9964,N_9515);
and U10105 (N_10105,N_9548,N_9746);
nand U10106 (N_10106,N_9664,N_9579);
or U10107 (N_10107,N_9652,N_9614);
or U10108 (N_10108,N_9772,N_9822);
and U10109 (N_10109,N_9743,N_9715);
xnor U10110 (N_10110,N_9911,N_9809);
nand U10111 (N_10111,N_9734,N_9622);
nand U10112 (N_10112,N_9700,N_9787);
or U10113 (N_10113,N_9994,N_9698);
nand U10114 (N_10114,N_9844,N_9681);
nand U10115 (N_10115,N_9709,N_9797);
and U10116 (N_10116,N_9922,N_9829);
nand U10117 (N_10117,N_9833,N_9924);
nor U10118 (N_10118,N_9532,N_9649);
nand U10119 (N_10119,N_9719,N_9575);
xnor U10120 (N_10120,N_9693,N_9904);
nor U10121 (N_10121,N_9937,N_9749);
nand U10122 (N_10122,N_9510,N_9588);
nor U10123 (N_10123,N_9957,N_9895);
xor U10124 (N_10124,N_9951,N_9780);
nand U10125 (N_10125,N_9671,N_9956);
nand U10126 (N_10126,N_9529,N_9686);
xor U10127 (N_10127,N_9565,N_9866);
xnor U10128 (N_10128,N_9503,N_9701);
nor U10129 (N_10129,N_9820,N_9599);
xnor U10130 (N_10130,N_9755,N_9760);
nor U10131 (N_10131,N_9838,N_9680);
nand U10132 (N_10132,N_9763,N_9636);
xor U10133 (N_10133,N_9523,N_9889);
nand U10134 (N_10134,N_9587,N_9944);
xor U10135 (N_10135,N_9962,N_9535);
or U10136 (N_10136,N_9849,N_9502);
xor U10137 (N_10137,N_9848,N_9509);
or U10138 (N_10138,N_9978,N_9558);
xnor U10139 (N_10139,N_9990,N_9717);
and U10140 (N_10140,N_9544,N_9725);
nand U10141 (N_10141,N_9830,N_9537);
or U10142 (N_10142,N_9720,N_9909);
or U10143 (N_10143,N_9847,N_9857);
xor U10144 (N_10144,N_9627,N_9757);
and U10145 (N_10145,N_9753,N_9906);
xor U10146 (N_10146,N_9890,N_9557);
nor U10147 (N_10147,N_9536,N_9707);
nand U10148 (N_10148,N_9522,N_9654);
nand U10149 (N_10149,N_9690,N_9708);
and U10150 (N_10150,N_9736,N_9626);
nand U10151 (N_10151,N_9660,N_9840);
xnor U10152 (N_10152,N_9540,N_9935);
xnor U10153 (N_10153,N_9865,N_9887);
xnor U10154 (N_10154,N_9714,N_9641);
and U10155 (N_10155,N_9744,N_9882);
xor U10156 (N_10156,N_9703,N_9791);
nor U10157 (N_10157,N_9796,N_9646);
nor U10158 (N_10158,N_9521,N_9767);
xnor U10159 (N_10159,N_9819,N_9824);
xor U10160 (N_10160,N_9871,N_9968);
xnor U10161 (N_10161,N_9948,N_9582);
and U10162 (N_10162,N_9912,N_9547);
nor U10163 (N_10163,N_9518,N_9837);
nor U10164 (N_10164,N_9880,N_9624);
nor U10165 (N_10165,N_9670,N_9733);
nor U10166 (N_10166,N_9983,N_9534);
or U10167 (N_10167,N_9724,N_9873);
nand U10168 (N_10168,N_9741,N_9541);
and U10169 (N_10169,N_9967,N_9603);
or U10170 (N_10170,N_9798,N_9953);
and U10171 (N_10171,N_9963,N_9580);
nand U10172 (N_10172,N_9926,N_9712);
nor U10173 (N_10173,N_9813,N_9942);
and U10174 (N_10174,N_9933,N_9538);
nand U10175 (N_10175,N_9713,N_9516);
nand U10176 (N_10176,N_9929,N_9751);
nor U10177 (N_10177,N_9595,N_9759);
xnor U10178 (N_10178,N_9596,N_9965);
nand U10179 (N_10179,N_9959,N_9814);
xor U10180 (N_10180,N_9666,N_9668);
nor U10181 (N_10181,N_9947,N_9803);
and U10182 (N_10182,N_9711,N_9658);
or U10183 (N_10183,N_9585,N_9908);
nand U10184 (N_10184,N_9571,N_9729);
nand U10185 (N_10185,N_9631,N_9793);
or U10186 (N_10186,N_9966,N_9855);
or U10187 (N_10187,N_9916,N_9954);
nand U10188 (N_10188,N_9676,N_9706);
nor U10189 (N_10189,N_9528,N_9662);
xnor U10190 (N_10190,N_9632,N_9687);
nand U10191 (N_10191,N_9555,N_9525);
or U10192 (N_10192,N_9569,N_9817);
nand U10193 (N_10193,N_9853,N_9893);
and U10194 (N_10194,N_9704,N_9564);
and U10195 (N_10195,N_9910,N_9645);
nand U10196 (N_10196,N_9543,N_9550);
or U10197 (N_10197,N_9806,N_9876);
or U10198 (N_10198,N_9988,N_9644);
xor U10199 (N_10199,N_9667,N_9539);
xnor U10200 (N_10200,N_9730,N_9823);
or U10201 (N_10201,N_9651,N_9517);
xnor U10202 (N_10202,N_9642,N_9610);
and U10203 (N_10203,N_9669,N_9834);
nand U10204 (N_10204,N_9665,N_9615);
nand U10205 (N_10205,N_9608,N_9752);
or U10206 (N_10206,N_9868,N_9613);
or U10207 (N_10207,N_9577,N_9991);
xor U10208 (N_10208,N_9972,N_9795);
and U10209 (N_10209,N_9843,N_9600);
xor U10210 (N_10210,N_9810,N_9768);
or U10211 (N_10211,N_9919,N_9578);
and U10212 (N_10212,N_9874,N_9777);
xnor U10213 (N_10213,N_9949,N_9695);
xor U10214 (N_10214,N_9902,N_9995);
nor U10215 (N_10215,N_9758,N_9846);
xor U10216 (N_10216,N_9794,N_9835);
or U10217 (N_10217,N_9778,N_9827);
and U10218 (N_10218,N_9549,N_9917);
nand U10219 (N_10219,N_9621,N_9732);
and U10220 (N_10220,N_9940,N_9605);
xnor U10221 (N_10221,N_9771,N_9722);
nand U10222 (N_10222,N_9685,N_9601);
or U10223 (N_10223,N_9657,N_9619);
nor U10224 (N_10224,N_9842,N_9747);
or U10225 (N_10225,N_9737,N_9533);
xor U10226 (N_10226,N_9553,N_9630);
nor U10227 (N_10227,N_9727,N_9609);
and U10228 (N_10228,N_9639,N_9592);
or U10229 (N_10229,N_9574,N_9647);
nor U10230 (N_10230,N_9683,N_9993);
or U10231 (N_10231,N_9656,N_9661);
and U10232 (N_10232,N_9811,N_9815);
nand U10233 (N_10233,N_9586,N_9989);
or U10234 (N_10234,N_9554,N_9659);
or U10235 (N_10235,N_9856,N_9888);
or U10236 (N_10236,N_9696,N_9852);
nand U10237 (N_10237,N_9785,N_9863);
nand U10238 (N_10238,N_9504,N_9973);
xnor U10239 (N_10239,N_9958,N_9750);
nor U10240 (N_10240,N_9927,N_9884);
nand U10241 (N_10241,N_9650,N_9756);
xor U10242 (N_10242,N_9799,N_9992);
xnor U10243 (N_10243,N_9867,N_9979);
nor U10244 (N_10244,N_9705,N_9818);
and U10245 (N_10245,N_9623,N_9766);
nand U10246 (N_10246,N_9898,N_9625);
xor U10247 (N_10247,N_9896,N_9977);
and U10248 (N_10248,N_9832,N_9802);
nor U10249 (N_10249,N_9612,N_9526);
xnor U10250 (N_10250,N_9759,N_9508);
nand U10251 (N_10251,N_9513,N_9753);
and U10252 (N_10252,N_9838,N_9633);
nand U10253 (N_10253,N_9781,N_9815);
nand U10254 (N_10254,N_9872,N_9967);
nand U10255 (N_10255,N_9658,N_9580);
nand U10256 (N_10256,N_9810,N_9650);
nor U10257 (N_10257,N_9823,N_9905);
nor U10258 (N_10258,N_9752,N_9994);
nand U10259 (N_10259,N_9925,N_9966);
nor U10260 (N_10260,N_9927,N_9746);
nor U10261 (N_10261,N_9873,N_9695);
or U10262 (N_10262,N_9845,N_9726);
and U10263 (N_10263,N_9625,N_9992);
and U10264 (N_10264,N_9885,N_9511);
or U10265 (N_10265,N_9994,N_9607);
or U10266 (N_10266,N_9831,N_9680);
or U10267 (N_10267,N_9937,N_9824);
xnor U10268 (N_10268,N_9721,N_9847);
nand U10269 (N_10269,N_9688,N_9593);
nor U10270 (N_10270,N_9603,N_9687);
and U10271 (N_10271,N_9817,N_9637);
nand U10272 (N_10272,N_9501,N_9908);
and U10273 (N_10273,N_9787,N_9942);
nand U10274 (N_10274,N_9716,N_9624);
xor U10275 (N_10275,N_9934,N_9740);
or U10276 (N_10276,N_9903,N_9781);
xor U10277 (N_10277,N_9976,N_9662);
nor U10278 (N_10278,N_9931,N_9551);
nand U10279 (N_10279,N_9751,N_9994);
and U10280 (N_10280,N_9899,N_9975);
or U10281 (N_10281,N_9774,N_9806);
nor U10282 (N_10282,N_9768,N_9795);
nor U10283 (N_10283,N_9843,N_9645);
or U10284 (N_10284,N_9776,N_9604);
nor U10285 (N_10285,N_9865,N_9823);
and U10286 (N_10286,N_9949,N_9657);
xnor U10287 (N_10287,N_9717,N_9979);
nor U10288 (N_10288,N_9866,N_9622);
nand U10289 (N_10289,N_9527,N_9658);
nor U10290 (N_10290,N_9706,N_9758);
xor U10291 (N_10291,N_9895,N_9756);
nor U10292 (N_10292,N_9912,N_9813);
nor U10293 (N_10293,N_9867,N_9636);
or U10294 (N_10294,N_9974,N_9703);
and U10295 (N_10295,N_9779,N_9521);
nor U10296 (N_10296,N_9718,N_9592);
or U10297 (N_10297,N_9535,N_9595);
nor U10298 (N_10298,N_9983,N_9825);
xor U10299 (N_10299,N_9761,N_9867);
and U10300 (N_10300,N_9554,N_9776);
nand U10301 (N_10301,N_9942,N_9886);
or U10302 (N_10302,N_9925,N_9980);
or U10303 (N_10303,N_9614,N_9528);
or U10304 (N_10304,N_9785,N_9800);
nand U10305 (N_10305,N_9753,N_9688);
and U10306 (N_10306,N_9792,N_9918);
and U10307 (N_10307,N_9927,N_9948);
xor U10308 (N_10308,N_9607,N_9512);
nand U10309 (N_10309,N_9533,N_9988);
nor U10310 (N_10310,N_9867,N_9823);
and U10311 (N_10311,N_9775,N_9990);
or U10312 (N_10312,N_9985,N_9570);
nand U10313 (N_10313,N_9618,N_9601);
nand U10314 (N_10314,N_9601,N_9937);
xnor U10315 (N_10315,N_9910,N_9914);
and U10316 (N_10316,N_9604,N_9824);
nand U10317 (N_10317,N_9530,N_9762);
nand U10318 (N_10318,N_9705,N_9577);
nor U10319 (N_10319,N_9519,N_9620);
or U10320 (N_10320,N_9779,N_9964);
and U10321 (N_10321,N_9976,N_9810);
xor U10322 (N_10322,N_9973,N_9605);
or U10323 (N_10323,N_9543,N_9741);
and U10324 (N_10324,N_9989,N_9610);
and U10325 (N_10325,N_9946,N_9817);
and U10326 (N_10326,N_9923,N_9750);
and U10327 (N_10327,N_9861,N_9648);
and U10328 (N_10328,N_9791,N_9884);
nor U10329 (N_10329,N_9887,N_9940);
xor U10330 (N_10330,N_9944,N_9931);
nor U10331 (N_10331,N_9652,N_9756);
or U10332 (N_10332,N_9556,N_9781);
nor U10333 (N_10333,N_9697,N_9662);
nor U10334 (N_10334,N_9856,N_9931);
or U10335 (N_10335,N_9702,N_9636);
nor U10336 (N_10336,N_9551,N_9700);
xor U10337 (N_10337,N_9661,N_9620);
nand U10338 (N_10338,N_9809,N_9538);
nand U10339 (N_10339,N_9945,N_9968);
nand U10340 (N_10340,N_9773,N_9816);
nand U10341 (N_10341,N_9891,N_9878);
nand U10342 (N_10342,N_9568,N_9648);
nor U10343 (N_10343,N_9532,N_9761);
nor U10344 (N_10344,N_9805,N_9784);
and U10345 (N_10345,N_9570,N_9742);
xor U10346 (N_10346,N_9613,N_9869);
nor U10347 (N_10347,N_9704,N_9659);
and U10348 (N_10348,N_9617,N_9789);
or U10349 (N_10349,N_9945,N_9639);
nor U10350 (N_10350,N_9696,N_9992);
nand U10351 (N_10351,N_9821,N_9608);
and U10352 (N_10352,N_9698,N_9611);
and U10353 (N_10353,N_9984,N_9583);
xnor U10354 (N_10354,N_9986,N_9670);
xnor U10355 (N_10355,N_9822,N_9948);
and U10356 (N_10356,N_9571,N_9817);
or U10357 (N_10357,N_9865,N_9959);
or U10358 (N_10358,N_9705,N_9990);
nand U10359 (N_10359,N_9557,N_9856);
nand U10360 (N_10360,N_9574,N_9819);
nand U10361 (N_10361,N_9711,N_9632);
nand U10362 (N_10362,N_9894,N_9873);
nor U10363 (N_10363,N_9877,N_9848);
and U10364 (N_10364,N_9635,N_9566);
or U10365 (N_10365,N_9790,N_9534);
nor U10366 (N_10366,N_9828,N_9958);
or U10367 (N_10367,N_9934,N_9989);
nor U10368 (N_10368,N_9582,N_9524);
and U10369 (N_10369,N_9596,N_9695);
and U10370 (N_10370,N_9781,N_9609);
nand U10371 (N_10371,N_9506,N_9783);
xor U10372 (N_10372,N_9756,N_9610);
and U10373 (N_10373,N_9794,N_9976);
and U10374 (N_10374,N_9881,N_9865);
xor U10375 (N_10375,N_9698,N_9742);
nor U10376 (N_10376,N_9590,N_9899);
and U10377 (N_10377,N_9791,N_9934);
nor U10378 (N_10378,N_9740,N_9677);
or U10379 (N_10379,N_9597,N_9840);
nand U10380 (N_10380,N_9911,N_9849);
and U10381 (N_10381,N_9993,N_9898);
and U10382 (N_10382,N_9646,N_9877);
nand U10383 (N_10383,N_9578,N_9551);
nor U10384 (N_10384,N_9874,N_9930);
or U10385 (N_10385,N_9925,N_9674);
nand U10386 (N_10386,N_9519,N_9904);
nand U10387 (N_10387,N_9670,N_9894);
nand U10388 (N_10388,N_9593,N_9923);
or U10389 (N_10389,N_9895,N_9516);
or U10390 (N_10390,N_9794,N_9782);
nand U10391 (N_10391,N_9775,N_9587);
or U10392 (N_10392,N_9670,N_9579);
and U10393 (N_10393,N_9829,N_9675);
and U10394 (N_10394,N_9632,N_9883);
nand U10395 (N_10395,N_9816,N_9826);
nand U10396 (N_10396,N_9927,N_9853);
or U10397 (N_10397,N_9591,N_9675);
nand U10398 (N_10398,N_9664,N_9561);
xnor U10399 (N_10399,N_9959,N_9549);
and U10400 (N_10400,N_9793,N_9933);
nor U10401 (N_10401,N_9789,N_9767);
xnor U10402 (N_10402,N_9926,N_9789);
nor U10403 (N_10403,N_9710,N_9694);
nor U10404 (N_10404,N_9981,N_9836);
nand U10405 (N_10405,N_9686,N_9917);
xnor U10406 (N_10406,N_9989,N_9753);
xnor U10407 (N_10407,N_9524,N_9544);
and U10408 (N_10408,N_9895,N_9540);
xor U10409 (N_10409,N_9501,N_9734);
xnor U10410 (N_10410,N_9967,N_9862);
and U10411 (N_10411,N_9544,N_9929);
and U10412 (N_10412,N_9561,N_9727);
and U10413 (N_10413,N_9997,N_9996);
nand U10414 (N_10414,N_9678,N_9967);
nand U10415 (N_10415,N_9903,N_9512);
and U10416 (N_10416,N_9516,N_9700);
xor U10417 (N_10417,N_9587,N_9741);
and U10418 (N_10418,N_9896,N_9598);
nand U10419 (N_10419,N_9936,N_9522);
nand U10420 (N_10420,N_9910,N_9945);
and U10421 (N_10421,N_9855,N_9978);
nand U10422 (N_10422,N_9554,N_9860);
nand U10423 (N_10423,N_9502,N_9965);
or U10424 (N_10424,N_9780,N_9910);
xor U10425 (N_10425,N_9917,N_9605);
nor U10426 (N_10426,N_9997,N_9543);
nor U10427 (N_10427,N_9839,N_9917);
nand U10428 (N_10428,N_9944,N_9536);
or U10429 (N_10429,N_9858,N_9503);
xor U10430 (N_10430,N_9636,N_9671);
and U10431 (N_10431,N_9890,N_9728);
or U10432 (N_10432,N_9776,N_9692);
and U10433 (N_10433,N_9642,N_9535);
or U10434 (N_10434,N_9777,N_9519);
nand U10435 (N_10435,N_9695,N_9918);
nand U10436 (N_10436,N_9833,N_9708);
or U10437 (N_10437,N_9585,N_9926);
and U10438 (N_10438,N_9904,N_9768);
nand U10439 (N_10439,N_9747,N_9959);
xnor U10440 (N_10440,N_9613,N_9648);
xor U10441 (N_10441,N_9869,N_9637);
nor U10442 (N_10442,N_9552,N_9575);
or U10443 (N_10443,N_9756,N_9937);
and U10444 (N_10444,N_9642,N_9567);
and U10445 (N_10445,N_9694,N_9567);
xor U10446 (N_10446,N_9700,N_9531);
nand U10447 (N_10447,N_9942,N_9533);
nor U10448 (N_10448,N_9742,N_9809);
and U10449 (N_10449,N_9542,N_9632);
nand U10450 (N_10450,N_9927,N_9529);
xor U10451 (N_10451,N_9676,N_9703);
and U10452 (N_10452,N_9503,N_9699);
xnor U10453 (N_10453,N_9965,N_9998);
or U10454 (N_10454,N_9589,N_9636);
nor U10455 (N_10455,N_9837,N_9817);
nor U10456 (N_10456,N_9734,N_9830);
or U10457 (N_10457,N_9524,N_9563);
xnor U10458 (N_10458,N_9733,N_9565);
or U10459 (N_10459,N_9982,N_9664);
nand U10460 (N_10460,N_9940,N_9929);
or U10461 (N_10461,N_9957,N_9879);
nand U10462 (N_10462,N_9721,N_9875);
and U10463 (N_10463,N_9965,N_9733);
or U10464 (N_10464,N_9784,N_9555);
nor U10465 (N_10465,N_9579,N_9589);
and U10466 (N_10466,N_9723,N_9965);
xnor U10467 (N_10467,N_9784,N_9682);
nor U10468 (N_10468,N_9725,N_9582);
and U10469 (N_10469,N_9678,N_9698);
and U10470 (N_10470,N_9819,N_9669);
nor U10471 (N_10471,N_9934,N_9500);
xnor U10472 (N_10472,N_9839,N_9718);
nor U10473 (N_10473,N_9958,N_9911);
nor U10474 (N_10474,N_9515,N_9544);
or U10475 (N_10475,N_9840,N_9609);
nand U10476 (N_10476,N_9735,N_9914);
or U10477 (N_10477,N_9857,N_9529);
nor U10478 (N_10478,N_9927,N_9509);
or U10479 (N_10479,N_9917,N_9895);
xor U10480 (N_10480,N_9965,N_9541);
nor U10481 (N_10481,N_9813,N_9826);
and U10482 (N_10482,N_9796,N_9805);
nor U10483 (N_10483,N_9990,N_9759);
or U10484 (N_10484,N_9733,N_9660);
nand U10485 (N_10485,N_9533,N_9981);
and U10486 (N_10486,N_9976,N_9816);
and U10487 (N_10487,N_9598,N_9789);
nor U10488 (N_10488,N_9766,N_9934);
or U10489 (N_10489,N_9615,N_9627);
and U10490 (N_10490,N_9575,N_9737);
and U10491 (N_10491,N_9746,N_9598);
nor U10492 (N_10492,N_9507,N_9838);
nor U10493 (N_10493,N_9560,N_9707);
and U10494 (N_10494,N_9582,N_9631);
and U10495 (N_10495,N_9884,N_9869);
nor U10496 (N_10496,N_9937,N_9620);
nand U10497 (N_10497,N_9782,N_9982);
or U10498 (N_10498,N_9907,N_9946);
nand U10499 (N_10499,N_9639,N_9559);
nor U10500 (N_10500,N_10277,N_10055);
xnor U10501 (N_10501,N_10409,N_10246);
and U10502 (N_10502,N_10083,N_10245);
xnor U10503 (N_10503,N_10155,N_10071);
nor U10504 (N_10504,N_10313,N_10173);
nand U10505 (N_10505,N_10294,N_10367);
xnor U10506 (N_10506,N_10188,N_10331);
nand U10507 (N_10507,N_10230,N_10272);
and U10508 (N_10508,N_10453,N_10225);
nor U10509 (N_10509,N_10199,N_10201);
xor U10510 (N_10510,N_10027,N_10168);
and U10511 (N_10511,N_10326,N_10039);
nand U10512 (N_10512,N_10337,N_10397);
nor U10513 (N_10513,N_10308,N_10011);
nor U10514 (N_10514,N_10218,N_10260);
and U10515 (N_10515,N_10033,N_10469);
and U10516 (N_10516,N_10498,N_10170);
or U10517 (N_10517,N_10390,N_10096);
nand U10518 (N_10518,N_10169,N_10175);
nand U10519 (N_10519,N_10328,N_10043);
or U10520 (N_10520,N_10004,N_10388);
xnor U10521 (N_10521,N_10040,N_10322);
and U10522 (N_10522,N_10148,N_10319);
or U10523 (N_10523,N_10354,N_10456);
and U10524 (N_10524,N_10248,N_10419);
nand U10525 (N_10525,N_10266,N_10053);
nand U10526 (N_10526,N_10344,N_10285);
nand U10527 (N_10527,N_10365,N_10242);
or U10528 (N_10528,N_10025,N_10446);
or U10529 (N_10529,N_10428,N_10420);
nor U10530 (N_10530,N_10416,N_10452);
xnor U10531 (N_10531,N_10396,N_10299);
nor U10532 (N_10532,N_10210,N_10433);
or U10533 (N_10533,N_10253,N_10327);
and U10534 (N_10534,N_10022,N_10069);
nand U10535 (N_10535,N_10220,N_10182);
xor U10536 (N_10536,N_10256,N_10394);
nand U10537 (N_10537,N_10012,N_10321);
and U10538 (N_10538,N_10198,N_10186);
xor U10539 (N_10539,N_10250,N_10343);
nor U10540 (N_10540,N_10228,N_10400);
nand U10541 (N_10541,N_10197,N_10429);
nand U10542 (N_10542,N_10282,N_10368);
or U10543 (N_10543,N_10317,N_10235);
nand U10544 (N_10544,N_10271,N_10203);
nand U10545 (N_10545,N_10481,N_10221);
and U10546 (N_10546,N_10492,N_10443);
nor U10547 (N_10547,N_10373,N_10112);
nand U10548 (N_10548,N_10440,N_10095);
and U10549 (N_10549,N_10142,N_10496);
and U10550 (N_10550,N_10130,N_10007);
nor U10551 (N_10551,N_10163,N_10264);
nand U10552 (N_10552,N_10167,N_10144);
and U10553 (N_10553,N_10067,N_10426);
or U10554 (N_10554,N_10063,N_10160);
xnor U10555 (N_10555,N_10061,N_10105);
xor U10556 (N_10556,N_10068,N_10091);
xnor U10557 (N_10557,N_10399,N_10474);
nand U10558 (N_10558,N_10306,N_10263);
and U10559 (N_10559,N_10042,N_10140);
nor U10560 (N_10560,N_10449,N_10280);
nand U10561 (N_10561,N_10234,N_10392);
and U10562 (N_10562,N_10251,N_10414);
xnor U10563 (N_10563,N_10060,N_10329);
and U10564 (N_10564,N_10072,N_10323);
and U10565 (N_10565,N_10276,N_10239);
nand U10566 (N_10566,N_10307,N_10471);
and U10567 (N_10567,N_10187,N_10301);
xor U10568 (N_10568,N_10442,N_10461);
nand U10569 (N_10569,N_10048,N_10017);
or U10570 (N_10570,N_10283,N_10162);
and U10571 (N_10571,N_10257,N_10006);
and U10572 (N_10572,N_10190,N_10270);
or U10573 (N_10573,N_10171,N_10044);
nand U10574 (N_10574,N_10172,N_10448);
and U10575 (N_10575,N_10062,N_10389);
xor U10576 (N_10576,N_10114,N_10491);
xnor U10577 (N_10577,N_10485,N_10057);
nor U10578 (N_10578,N_10108,N_10240);
xor U10579 (N_10579,N_10085,N_10339);
and U10580 (N_10580,N_10384,N_10193);
nor U10581 (N_10581,N_10066,N_10434);
nand U10582 (N_10582,N_10413,N_10084);
and U10583 (N_10583,N_10181,N_10178);
and U10584 (N_10584,N_10191,N_10097);
nor U10585 (N_10585,N_10064,N_10179);
and U10586 (N_10586,N_10134,N_10138);
or U10587 (N_10587,N_10415,N_10425);
or U10588 (N_10588,N_10213,N_10423);
xnor U10589 (N_10589,N_10195,N_10212);
xor U10590 (N_10590,N_10151,N_10458);
or U10591 (N_10591,N_10295,N_10079);
nor U10592 (N_10592,N_10102,N_10204);
or U10593 (N_10593,N_10098,N_10335);
or U10594 (N_10594,N_10466,N_10075);
and U10595 (N_10595,N_10464,N_10441);
xor U10596 (N_10596,N_10359,N_10347);
and U10597 (N_10597,N_10303,N_10013);
xor U10598 (N_10598,N_10003,N_10459);
nand U10599 (N_10599,N_10194,N_10244);
nor U10600 (N_10600,N_10137,N_10473);
and U10601 (N_10601,N_10412,N_10383);
and U10602 (N_10602,N_10174,N_10482);
and U10603 (N_10603,N_10126,N_10046);
and U10604 (N_10604,N_10334,N_10393);
or U10605 (N_10605,N_10268,N_10348);
nor U10606 (N_10606,N_10312,N_10031);
and U10607 (N_10607,N_10372,N_10341);
xor U10608 (N_10608,N_10052,N_10118);
nor U10609 (N_10609,N_10088,N_10408);
nor U10610 (N_10610,N_10462,N_10350);
xor U10611 (N_10611,N_10176,N_10345);
or U10612 (N_10612,N_10093,N_10333);
xor U10613 (N_10613,N_10038,N_10028);
or U10614 (N_10614,N_10477,N_10106);
or U10615 (N_10615,N_10216,N_10379);
or U10616 (N_10616,N_10121,N_10489);
xor U10617 (N_10617,N_10499,N_10437);
nand U10618 (N_10618,N_10460,N_10478);
xnor U10619 (N_10619,N_10450,N_10024);
nor U10620 (N_10620,N_10119,N_10382);
nor U10621 (N_10621,N_10374,N_10128);
and U10622 (N_10622,N_10479,N_10315);
and U10623 (N_10623,N_10249,N_10153);
xnor U10624 (N_10624,N_10135,N_10364);
and U10625 (N_10625,N_10385,N_10122);
nor U10626 (N_10626,N_10073,N_10349);
xnor U10627 (N_10627,N_10184,N_10161);
nand U10628 (N_10628,N_10418,N_10497);
nor U10629 (N_10629,N_10158,N_10451);
and U10630 (N_10630,N_10465,N_10141);
nor U10631 (N_10631,N_10094,N_10275);
or U10632 (N_10632,N_10332,N_10092);
nand U10633 (N_10633,N_10431,N_10115);
xnor U10634 (N_10634,N_10300,N_10304);
or U10635 (N_10635,N_10457,N_10136);
xnor U10636 (N_10636,N_10355,N_10041);
nand U10637 (N_10637,N_10487,N_10480);
xnor U10638 (N_10638,N_10254,N_10021);
or U10639 (N_10639,N_10056,N_10340);
nand U10640 (N_10640,N_10346,N_10010);
nand U10641 (N_10641,N_10445,N_10410);
and U10642 (N_10642,N_10087,N_10356);
and U10643 (N_10643,N_10082,N_10147);
nand U10644 (N_10644,N_10018,N_10157);
xnor U10645 (N_10645,N_10164,N_10192);
or U10646 (N_10646,N_10086,N_10180);
nor U10647 (N_10647,N_10290,N_10261);
or U10648 (N_10648,N_10404,N_10016);
and U10649 (N_10649,N_10269,N_10302);
xnor U10650 (N_10650,N_10034,N_10320);
and U10651 (N_10651,N_10424,N_10402);
and U10652 (N_10652,N_10131,N_10101);
and U10653 (N_10653,N_10380,N_10165);
xnor U10654 (N_10654,N_10223,N_10472);
and U10655 (N_10655,N_10037,N_10077);
xor U10656 (N_10656,N_10232,N_10117);
nor U10657 (N_10657,N_10065,N_10375);
and U10658 (N_10658,N_10455,N_10387);
and U10659 (N_10659,N_10475,N_10361);
and U10660 (N_10660,N_10298,N_10316);
xor U10661 (N_10661,N_10336,N_10403);
nor U10662 (N_10662,N_10495,N_10377);
xor U10663 (N_10663,N_10243,N_10120);
or U10664 (N_10664,N_10338,N_10274);
nand U10665 (N_10665,N_10314,N_10351);
nand U10666 (N_10666,N_10454,N_10233);
nor U10667 (N_10667,N_10376,N_10211);
xnor U10668 (N_10668,N_10405,N_10227);
nand U10669 (N_10669,N_10255,N_10159);
nand U10670 (N_10670,N_10435,N_10058);
nand U10671 (N_10671,N_10287,N_10100);
and U10672 (N_10672,N_10305,N_10262);
nor U10673 (N_10673,N_10116,N_10342);
xor U10674 (N_10674,N_10353,N_10047);
or U10675 (N_10675,N_10008,N_10422);
nor U10676 (N_10676,N_10045,N_10133);
xnor U10677 (N_10677,N_10395,N_10059);
nand U10678 (N_10678,N_10296,N_10439);
or U10679 (N_10679,N_10463,N_10050);
nand U10680 (N_10680,N_10154,N_10123);
nand U10681 (N_10681,N_10113,N_10090);
nand U10682 (N_10682,N_10398,N_10378);
xor U10683 (N_10683,N_10486,N_10430);
or U10684 (N_10684,N_10224,N_10156);
nor U10685 (N_10685,N_10222,N_10483);
nand U10686 (N_10686,N_10076,N_10104);
xnor U10687 (N_10687,N_10209,N_10109);
and U10688 (N_10688,N_10129,N_10371);
or U10689 (N_10689,N_10166,N_10318);
nand U10690 (N_10690,N_10330,N_10000);
nor U10691 (N_10691,N_10411,N_10447);
or U10692 (N_10692,N_10089,N_10177);
xnor U10693 (N_10693,N_10436,N_10081);
and U10694 (N_10694,N_10247,N_10202);
xor U10695 (N_10695,N_10444,N_10488);
nand U10696 (N_10696,N_10152,N_10014);
xor U10697 (N_10697,N_10196,N_10421);
and U10698 (N_10698,N_10309,N_10107);
or U10699 (N_10699,N_10265,N_10470);
or U10700 (N_10700,N_10019,N_10110);
xnor U10701 (N_10701,N_10362,N_10205);
xor U10702 (N_10702,N_10183,N_10310);
xor U10703 (N_10703,N_10292,N_10284);
nor U10704 (N_10704,N_10207,N_10074);
xor U10705 (N_10705,N_10078,N_10150);
nor U10706 (N_10706,N_10001,N_10200);
nand U10707 (N_10707,N_10381,N_10149);
and U10708 (N_10708,N_10124,N_10029);
and U10709 (N_10709,N_10417,N_10139);
nand U10710 (N_10710,N_10311,N_10281);
nor U10711 (N_10711,N_10357,N_10009);
and U10712 (N_10712,N_10229,N_10267);
and U10713 (N_10713,N_10325,N_10427);
and U10714 (N_10714,N_10206,N_10238);
or U10715 (N_10715,N_10070,N_10370);
xor U10716 (N_10716,N_10406,N_10363);
and U10717 (N_10717,N_10468,N_10020);
nor U10718 (N_10718,N_10125,N_10476);
xnor U10719 (N_10719,N_10493,N_10217);
nor U10720 (N_10720,N_10484,N_10236);
xnor U10721 (N_10721,N_10185,N_10103);
nor U10722 (N_10722,N_10438,N_10286);
and U10723 (N_10723,N_10189,N_10111);
or U10724 (N_10724,N_10054,N_10002);
nand U10725 (N_10725,N_10352,N_10005);
nor U10726 (N_10726,N_10231,N_10401);
and U10727 (N_10727,N_10490,N_10226);
nor U10728 (N_10728,N_10143,N_10051);
or U10729 (N_10729,N_10132,N_10215);
and U10730 (N_10730,N_10369,N_10015);
or U10731 (N_10731,N_10288,N_10360);
xor U10732 (N_10732,N_10035,N_10324);
xor U10733 (N_10733,N_10049,N_10279);
and U10734 (N_10734,N_10023,N_10259);
and U10735 (N_10735,N_10291,N_10391);
or U10736 (N_10736,N_10258,N_10026);
xnor U10737 (N_10737,N_10030,N_10146);
nand U10738 (N_10738,N_10032,N_10273);
or U10739 (N_10739,N_10214,N_10219);
nand U10740 (N_10740,N_10366,N_10080);
or U10741 (N_10741,N_10252,N_10208);
xnor U10742 (N_10742,N_10293,N_10145);
nor U10743 (N_10743,N_10467,N_10386);
nand U10744 (N_10744,N_10127,N_10297);
nor U10745 (N_10745,N_10289,N_10407);
nand U10746 (N_10746,N_10278,N_10432);
nand U10747 (N_10747,N_10099,N_10358);
nand U10748 (N_10748,N_10494,N_10237);
and U10749 (N_10749,N_10036,N_10241);
or U10750 (N_10750,N_10293,N_10113);
nor U10751 (N_10751,N_10256,N_10038);
or U10752 (N_10752,N_10386,N_10475);
nand U10753 (N_10753,N_10273,N_10433);
and U10754 (N_10754,N_10382,N_10053);
or U10755 (N_10755,N_10060,N_10347);
or U10756 (N_10756,N_10040,N_10036);
xor U10757 (N_10757,N_10221,N_10499);
nand U10758 (N_10758,N_10451,N_10072);
nor U10759 (N_10759,N_10020,N_10051);
and U10760 (N_10760,N_10231,N_10015);
xnor U10761 (N_10761,N_10475,N_10062);
xnor U10762 (N_10762,N_10497,N_10073);
nand U10763 (N_10763,N_10147,N_10218);
xor U10764 (N_10764,N_10172,N_10306);
nor U10765 (N_10765,N_10113,N_10356);
and U10766 (N_10766,N_10447,N_10093);
nor U10767 (N_10767,N_10014,N_10357);
nand U10768 (N_10768,N_10100,N_10302);
xor U10769 (N_10769,N_10014,N_10266);
nor U10770 (N_10770,N_10212,N_10088);
nor U10771 (N_10771,N_10351,N_10438);
or U10772 (N_10772,N_10129,N_10290);
nand U10773 (N_10773,N_10388,N_10059);
nor U10774 (N_10774,N_10187,N_10383);
nand U10775 (N_10775,N_10240,N_10493);
or U10776 (N_10776,N_10236,N_10237);
nor U10777 (N_10777,N_10338,N_10049);
nand U10778 (N_10778,N_10117,N_10306);
or U10779 (N_10779,N_10294,N_10361);
nor U10780 (N_10780,N_10154,N_10084);
nand U10781 (N_10781,N_10278,N_10347);
and U10782 (N_10782,N_10369,N_10220);
nor U10783 (N_10783,N_10479,N_10245);
and U10784 (N_10784,N_10045,N_10268);
xnor U10785 (N_10785,N_10341,N_10408);
and U10786 (N_10786,N_10031,N_10242);
xnor U10787 (N_10787,N_10316,N_10485);
or U10788 (N_10788,N_10006,N_10078);
xnor U10789 (N_10789,N_10363,N_10223);
and U10790 (N_10790,N_10489,N_10075);
or U10791 (N_10791,N_10022,N_10213);
nor U10792 (N_10792,N_10229,N_10453);
nand U10793 (N_10793,N_10262,N_10499);
or U10794 (N_10794,N_10343,N_10238);
nor U10795 (N_10795,N_10076,N_10496);
nor U10796 (N_10796,N_10110,N_10398);
nand U10797 (N_10797,N_10424,N_10141);
nand U10798 (N_10798,N_10497,N_10478);
or U10799 (N_10799,N_10014,N_10286);
nor U10800 (N_10800,N_10217,N_10195);
or U10801 (N_10801,N_10429,N_10302);
or U10802 (N_10802,N_10213,N_10408);
and U10803 (N_10803,N_10135,N_10376);
nor U10804 (N_10804,N_10339,N_10136);
nor U10805 (N_10805,N_10237,N_10028);
nor U10806 (N_10806,N_10491,N_10417);
nor U10807 (N_10807,N_10026,N_10224);
nor U10808 (N_10808,N_10233,N_10274);
or U10809 (N_10809,N_10015,N_10442);
nor U10810 (N_10810,N_10311,N_10286);
nand U10811 (N_10811,N_10378,N_10469);
nand U10812 (N_10812,N_10369,N_10147);
xor U10813 (N_10813,N_10346,N_10024);
and U10814 (N_10814,N_10300,N_10134);
xnor U10815 (N_10815,N_10486,N_10261);
xnor U10816 (N_10816,N_10036,N_10446);
and U10817 (N_10817,N_10437,N_10173);
or U10818 (N_10818,N_10147,N_10310);
nand U10819 (N_10819,N_10187,N_10273);
and U10820 (N_10820,N_10303,N_10435);
nand U10821 (N_10821,N_10131,N_10240);
nor U10822 (N_10822,N_10163,N_10182);
xnor U10823 (N_10823,N_10075,N_10355);
and U10824 (N_10824,N_10095,N_10190);
nand U10825 (N_10825,N_10230,N_10322);
and U10826 (N_10826,N_10453,N_10115);
and U10827 (N_10827,N_10484,N_10172);
nand U10828 (N_10828,N_10054,N_10124);
or U10829 (N_10829,N_10268,N_10247);
xor U10830 (N_10830,N_10256,N_10212);
nor U10831 (N_10831,N_10179,N_10284);
and U10832 (N_10832,N_10229,N_10228);
or U10833 (N_10833,N_10383,N_10351);
nor U10834 (N_10834,N_10178,N_10284);
nand U10835 (N_10835,N_10289,N_10395);
nor U10836 (N_10836,N_10390,N_10309);
or U10837 (N_10837,N_10364,N_10078);
nor U10838 (N_10838,N_10035,N_10351);
or U10839 (N_10839,N_10025,N_10292);
nor U10840 (N_10840,N_10099,N_10449);
nor U10841 (N_10841,N_10143,N_10103);
and U10842 (N_10842,N_10271,N_10057);
xnor U10843 (N_10843,N_10248,N_10247);
nand U10844 (N_10844,N_10302,N_10416);
nand U10845 (N_10845,N_10416,N_10159);
nand U10846 (N_10846,N_10305,N_10356);
xor U10847 (N_10847,N_10180,N_10037);
nand U10848 (N_10848,N_10204,N_10035);
xnor U10849 (N_10849,N_10416,N_10360);
xnor U10850 (N_10850,N_10499,N_10100);
or U10851 (N_10851,N_10474,N_10234);
nand U10852 (N_10852,N_10223,N_10471);
nand U10853 (N_10853,N_10399,N_10122);
nand U10854 (N_10854,N_10462,N_10128);
nand U10855 (N_10855,N_10130,N_10013);
or U10856 (N_10856,N_10158,N_10404);
nand U10857 (N_10857,N_10291,N_10207);
and U10858 (N_10858,N_10433,N_10141);
nand U10859 (N_10859,N_10281,N_10430);
nand U10860 (N_10860,N_10131,N_10485);
nor U10861 (N_10861,N_10133,N_10347);
nand U10862 (N_10862,N_10234,N_10061);
xor U10863 (N_10863,N_10353,N_10272);
nand U10864 (N_10864,N_10276,N_10372);
xnor U10865 (N_10865,N_10467,N_10137);
or U10866 (N_10866,N_10188,N_10490);
nand U10867 (N_10867,N_10186,N_10095);
or U10868 (N_10868,N_10099,N_10096);
and U10869 (N_10869,N_10093,N_10186);
nor U10870 (N_10870,N_10490,N_10100);
nor U10871 (N_10871,N_10499,N_10337);
nor U10872 (N_10872,N_10424,N_10435);
nor U10873 (N_10873,N_10291,N_10234);
xnor U10874 (N_10874,N_10112,N_10319);
or U10875 (N_10875,N_10260,N_10244);
and U10876 (N_10876,N_10136,N_10294);
xnor U10877 (N_10877,N_10452,N_10309);
and U10878 (N_10878,N_10083,N_10182);
nor U10879 (N_10879,N_10400,N_10439);
and U10880 (N_10880,N_10414,N_10136);
or U10881 (N_10881,N_10456,N_10453);
or U10882 (N_10882,N_10488,N_10206);
and U10883 (N_10883,N_10209,N_10186);
and U10884 (N_10884,N_10073,N_10209);
or U10885 (N_10885,N_10096,N_10243);
nor U10886 (N_10886,N_10161,N_10320);
xnor U10887 (N_10887,N_10492,N_10095);
and U10888 (N_10888,N_10486,N_10384);
xor U10889 (N_10889,N_10043,N_10325);
nand U10890 (N_10890,N_10301,N_10312);
xnor U10891 (N_10891,N_10063,N_10238);
nor U10892 (N_10892,N_10326,N_10198);
and U10893 (N_10893,N_10312,N_10114);
and U10894 (N_10894,N_10127,N_10155);
xnor U10895 (N_10895,N_10220,N_10088);
nor U10896 (N_10896,N_10196,N_10239);
or U10897 (N_10897,N_10090,N_10144);
and U10898 (N_10898,N_10121,N_10346);
or U10899 (N_10899,N_10488,N_10235);
or U10900 (N_10900,N_10131,N_10130);
and U10901 (N_10901,N_10349,N_10412);
or U10902 (N_10902,N_10395,N_10082);
xnor U10903 (N_10903,N_10460,N_10442);
xor U10904 (N_10904,N_10014,N_10132);
nor U10905 (N_10905,N_10191,N_10357);
nand U10906 (N_10906,N_10335,N_10167);
or U10907 (N_10907,N_10134,N_10007);
xnor U10908 (N_10908,N_10185,N_10344);
and U10909 (N_10909,N_10366,N_10133);
and U10910 (N_10910,N_10459,N_10254);
nand U10911 (N_10911,N_10267,N_10184);
nand U10912 (N_10912,N_10086,N_10321);
nand U10913 (N_10913,N_10116,N_10233);
xor U10914 (N_10914,N_10299,N_10132);
nor U10915 (N_10915,N_10411,N_10446);
nand U10916 (N_10916,N_10341,N_10095);
xnor U10917 (N_10917,N_10265,N_10309);
xor U10918 (N_10918,N_10273,N_10455);
nand U10919 (N_10919,N_10476,N_10305);
nor U10920 (N_10920,N_10042,N_10426);
nor U10921 (N_10921,N_10124,N_10050);
or U10922 (N_10922,N_10167,N_10399);
nor U10923 (N_10923,N_10379,N_10173);
nor U10924 (N_10924,N_10464,N_10418);
nor U10925 (N_10925,N_10386,N_10275);
nor U10926 (N_10926,N_10395,N_10178);
xor U10927 (N_10927,N_10372,N_10310);
nor U10928 (N_10928,N_10230,N_10067);
nor U10929 (N_10929,N_10064,N_10319);
and U10930 (N_10930,N_10103,N_10264);
and U10931 (N_10931,N_10092,N_10351);
and U10932 (N_10932,N_10290,N_10134);
or U10933 (N_10933,N_10340,N_10075);
nand U10934 (N_10934,N_10233,N_10498);
or U10935 (N_10935,N_10197,N_10359);
or U10936 (N_10936,N_10375,N_10027);
xnor U10937 (N_10937,N_10433,N_10476);
nand U10938 (N_10938,N_10409,N_10027);
and U10939 (N_10939,N_10048,N_10036);
or U10940 (N_10940,N_10364,N_10459);
or U10941 (N_10941,N_10420,N_10252);
and U10942 (N_10942,N_10002,N_10156);
xor U10943 (N_10943,N_10369,N_10233);
or U10944 (N_10944,N_10149,N_10221);
xnor U10945 (N_10945,N_10037,N_10306);
xnor U10946 (N_10946,N_10196,N_10158);
nand U10947 (N_10947,N_10155,N_10409);
xnor U10948 (N_10948,N_10097,N_10120);
and U10949 (N_10949,N_10212,N_10171);
nand U10950 (N_10950,N_10266,N_10396);
or U10951 (N_10951,N_10127,N_10016);
and U10952 (N_10952,N_10055,N_10069);
xor U10953 (N_10953,N_10278,N_10489);
and U10954 (N_10954,N_10429,N_10453);
or U10955 (N_10955,N_10160,N_10429);
or U10956 (N_10956,N_10403,N_10025);
xor U10957 (N_10957,N_10224,N_10358);
nor U10958 (N_10958,N_10171,N_10375);
nor U10959 (N_10959,N_10494,N_10340);
and U10960 (N_10960,N_10492,N_10197);
nor U10961 (N_10961,N_10321,N_10091);
or U10962 (N_10962,N_10079,N_10214);
nand U10963 (N_10963,N_10389,N_10064);
and U10964 (N_10964,N_10276,N_10403);
nor U10965 (N_10965,N_10367,N_10441);
nand U10966 (N_10966,N_10453,N_10359);
nand U10967 (N_10967,N_10301,N_10371);
and U10968 (N_10968,N_10157,N_10124);
nor U10969 (N_10969,N_10368,N_10283);
and U10970 (N_10970,N_10032,N_10468);
and U10971 (N_10971,N_10245,N_10269);
nand U10972 (N_10972,N_10311,N_10256);
and U10973 (N_10973,N_10345,N_10462);
xnor U10974 (N_10974,N_10320,N_10177);
nor U10975 (N_10975,N_10345,N_10295);
xnor U10976 (N_10976,N_10226,N_10123);
nand U10977 (N_10977,N_10308,N_10396);
and U10978 (N_10978,N_10480,N_10180);
or U10979 (N_10979,N_10098,N_10001);
or U10980 (N_10980,N_10079,N_10150);
nand U10981 (N_10981,N_10412,N_10469);
or U10982 (N_10982,N_10115,N_10081);
nand U10983 (N_10983,N_10226,N_10339);
or U10984 (N_10984,N_10156,N_10185);
nand U10985 (N_10985,N_10343,N_10373);
nand U10986 (N_10986,N_10401,N_10305);
or U10987 (N_10987,N_10389,N_10255);
or U10988 (N_10988,N_10141,N_10328);
or U10989 (N_10989,N_10016,N_10230);
or U10990 (N_10990,N_10308,N_10105);
nand U10991 (N_10991,N_10302,N_10347);
and U10992 (N_10992,N_10384,N_10396);
nor U10993 (N_10993,N_10091,N_10443);
nand U10994 (N_10994,N_10487,N_10027);
and U10995 (N_10995,N_10029,N_10401);
and U10996 (N_10996,N_10317,N_10132);
xnor U10997 (N_10997,N_10098,N_10094);
nand U10998 (N_10998,N_10321,N_10214);
nand U10999 (N_10999,N_10485,N_10345);
nand U11000 (N_11000,N_10952,N_10854);
or U11001 (N_11001,N_10721,N_10928);
and U11002 (N_11002,N_10543,N_10531);
nand U11003 (N_11003,N_10724,N_10768);
or U11004 (N_11004,N_10930,N_10949);
and U11005 (N_11005,N_10612,N_10986);
and U11006 (N_11006,N_10801,N_10894);
xor U11007 (N_11007,N_10882,N_10916);
xnor U11008 (N_11008,N_10876,N_10954);
nand U11009 (N_11009,N_10814,N_10793);
or U11010 (N_11010,N_10702,N_10656);
and U11011 (N_11011,N_10686,N_10792);
and U11012 (N_11012,N_10820,N_10956);
xnor U11013 (N_11013,N_10781,N_10697);
xor U11014 (N_11014,N_10677,N_10587);
nor U11015 (N_11015,N_10964,N_10770);
xnor U11016 (N_11016,N_10753,N_10861);
and U11017 (N_11017,N_10520,N_10623);
or U11018 (N_11018,N_10878,N_10761);
nand U11019 (N_11019,N_10832,N_10633);
nor U11020 (N_11020,N_10659,N_10936);
and U11021 (N_11021,N_10555,N_10553);
or U11022 (N_11022,N_10855,N_10707);
or U11023 (N_11023,N_10926,N_10608);
xor U11024 (N_11024,N_10980,N_10698);
nor U11025 (N_11025,N_10643,N_10767);
xnor U11026 (N_11026,N_10618,N_10764);
xor U11027 (N_11027,N_10534,N_10929);
nand U11028 (N_11028,N_10504,N_10819);
or U11029 (N_11029,N_10763,N_10756);
nor U11030 (N_11030,N_10765,N_10525);
nor U11031 (N_11031,N_10701,N_10849);
nand U11032 (N_11032,N_10691,N_10652);
or U11033 (N_11033,N_10584,N_10937);
nand U11034 (N_11034,N_10889,N_10911);
nand U11035 (N_11035,N_10913,N_10734);
nor U11036 (N_11036,N_10902,N_10635);
or U11037 (N_11037,N_10944,N_10884);
or U11038 (N_11038,N_10711,N_10542);
nand U11039 (N_11039,N_10751,N_10963);
nor U11040 (N_11040,N_10544,N_10737);
or U11041 (N_11041,N_10897,N_10715);
and U11042 (N_11042,N_10741,N_10971);
or U11043 (N_11043,N_10506,N_10708);
xor U11044 (N_11044,N_10616,N_10984);
nor U11045 (N_11045,N_10727,N_10901);
nor U11046 (N_11046,N_10967,N_10887);
or U11047 (N_11047,N_10851,N_10719);
nand U11048 (N_11048,N_10529,N_10747);
and U11049 (N_11049,N_10716,N_10759);
or U11050 (N_11050,N_10582,N_10805);
or U11051 (N_11051,N_10508,N_10824);
and U11052 (N_11052,N_10807,N_10953);
or U11053 (N_11053,N_10717,N_10994);
or U11054 (N_11054,N_10596,N_10591);
nand U11055 (N_11055,N_10562,N_10692);
nor U11056 (N_11056,N_10675,N_10650);
nor U11057 (N_11057,N_10774,N_10921);
nor U11058 (N_11058,N_10558,N_10512);
and U11059 (N_11059,N_10748,N_10546);
nor U11060 (N_11060,N_10837,N_10772);
or U11061 (N_11061,N_10996,N_10527);
xnor U11062 (N_11062,N_10760,N_10752);
nor U11063 (N_11063,N_10779,N_10771);
xnor U11064 (N_11064,N_10989,N_10755);
nand U11065 (N_11065,N_10905,N_10658);
nor U11066 (N_11066,N_10922,N_10950);
nor U11067 (N_11067,N_10890,N_10979);
or U11068 (N_11068,N_10733,N_10518);
xor U11069 (N_11069,N_10836,N_10990);
nand U11070 (N_11070,N_10668,N_10862);
xor U11071 (N_11071,N_10821,N_10679);
and U11072 (N_11072,N_10640,N_10706);
nand U11073 (N_11073,N_10941,N_10674);
xnor U11074 (N_11074,N_10648,N_10881);
or U11075 (N_11075,N_10540,N_10636);
nand U11076 (N_11076,N_10829,N_10647);
or U11077 (N_11077,N_10903,N_10704);
or U11078 (N_11078,N_10682,N_10627);
nor U11079 (N_11079,N_10830,N_10871);
nor U11080 (N_11080,N_10723,N_10597);
and U11081 (N_11081,N_10784,N_10539);
xnor U11082 (N_11082,N_10939,N_10766);
nand U11083 (N_11083,N_10530,N_10580);
or U11084 (N_11084,N_10965,N_10680);
nand U11085 (N_11085,N_10695,N_10599);
or U11086 (N_11086,N_10908,N_10883);
xor U11087 (N_11087,N_10607,N_10578);
and U11088 (N_11088,N_10978,N_10517);
nor U11089 (N_11089,N_10893,N_10728);
xnor U11090 (N_11090,N_10735,N_10725);
nor U11091 (N_11091,N_10545,N_10505);
nor U11092 (N_11092,N_10946,N_10993);
and U11093 (N_11093,N_10997,N_10565);
nand U11094 (N_11094,N_10948,N_10856);
xor U11095 (N_11095,N_10892,N_10914);
nand U11096 (N_11096,N_10615,N_10718);
nor U11097 (N_11097,N_10880,N_10696);
nand U11098 (N_11098,N_10931,N_10904);
or U11099 (N_11099,N_10834,N_10590);
nand U11100 (N_11100,N_10681,N_10804);
nor U11101 (N_11101,N_10572,N_10588);
and U11102 (N_11102,N_10577,N_10865);
and U11103 (N_11103,N_10667,N_10657);
or U11104 (N_11104,N_10649,N_10822);
or U11105 (N_11105,N_10869,N_10844);
nor U11106 (N_11106,N_10958,N_10620);
nand U11107 (N_11107,N_10644,N_10502);
and U11108 (N_11108,N_10800,N_10547);
and U11109 (N_11109,N_10666,N_10528);
and U11110 (N_11110,N_10524,N_10859);
or U11111 (N_11111,N_10569,N_10875);
and U11112 (N_11112,N_10817,N_10624);
xnor U11113 (N_11113,N_10799,N_10726);
xor U11114 (N_11114,N_10564,N_10561);
nor U11115 (N_11115,N_10977,N_10815);
nand U11116 (N_11116,N_10919,N_10754);
xor U11117 (N_11117,N_10720,N_10813);
nand U11118 (N_11118,N_10576,N_10992);
nand U11119 (N_11119,N_10773,N_10942);
and U11120 (N_11120,N_10983,N_10513);
nor U11121 (N_11121,N_10809,N_10567);
nand U11122 (N_11122,N_10791,N_10823);
or U11123 (N_11123,N_10522,N_10709);
and U11124 (N_11124,N_10787,N_10568);
nand U11125 (N_11125,N_10974,N_10617);
or U11126 (N_11126,N_10563,N_10625);
nand U11127 (N_11127,N_10628,N_10973);
nor U11128 (N_11128,N_10705,N_10629);
nand U11129 (N_11129,N_10541,N_10847);
xnor U11130 (N_11130,N_10743,N_10637);
xnor U11131 (N_11131,N_10619,N_10808);
xnor U11132 (N_11132,N_10828,N_10742);
nor U11133 (N_11133,N_10879,N_10598);
and U11134 (N_11134,N_10966,N_10998);
nor U11135 (N_11135,N_10671,N_10550);
and U11136 (N_11136,N_10662,N_10841);
and U11137 (N_11137,N_10672,N_10673);
nand U11138 (N_11138,N_10579,N_10638);
xnor U11139 (N_11139,N_10712,N_10669);
or U11140 (N_11140,N_10961,N_10898);
or U11141 (N_11141,N_10864,N_10573);
nor U11142 (N_11142,N_10777,N_10778);
or U11143 (N_11143,N_10639,N_10571);
xor U11144 (N_11144,N_10559,N_10714);
nor U11145 (N_11145,N_10603,N_10503);
xnor U11146 (N_11146,N_10873,N_10918);
xor U11147 (N_11147,N_10651,N_10654);
nand U11148 (N_11148,N_10910,N_10661);
and U11149 (N_11149,N_10899,N_10613);
nand U11150 (N_11150,N_10798,N_10907);
xor U11151 (N_11151,N_10835,N_10885);
xnor U11152 (N_11152,N_10703,N_10968);
xor U11153 (N_11153,N_10626,N_10976);
or U11154 (N_11154,N_10827,N_10886);
and U11155 (N_11155,N_10776,N_10631);
and U11156 (N_11156,N_10653,N_10501);
or U11157 (N_11157,N_10860,N_10690);
nor U11158 (N_11158,N_10664,N_10985);
or U11159 (N_11159,N_10663,N_10786);
and U11160 (N_11160,N_10858,N_10532);
xor U11161 (N_11161,N_10678,N_10556);
or U11162 (N_11162,N_10951,N_10866);
and U11163 (N_11163,N_10806,N_10925);
and U11164 (N_11164,N_10593,N_10700);
xor U11165 (N_11165,N_10960,N_10995);
xnor U11166 (N_11166,N_10857,N_10895);
xnor U11167 (N_11167,N_10660,N_10802);
nor U11168 (N_11168,N_10526,N_10785);
xor U11169 (N_11169,N_10611,N_10872);
nand U11170 (N_11170,N_10610,N_10509);
and U11171 (N_11171,N_10670,N_10699);
nand U11172 (N_11172,N_10840,N_10609);
xor U11173 (N_11173,N_10811,N_10812);
or U11174 (N_11174,N_10548,N_10917);
or U11175 (N_11175,N_10516,N_10713);
and U11176 (N_11176,N_10583,N_10622);
nand U11177 (N_11177,N_10825,N_10888);
or U11178 (N_11178,N_10537,N_10988);
and U11179 (N_11179,N_10843,N_10975);
and U11180 (N_11180,N_10630,N_10646);
nor U11181 (N_11181,N_10987,N_10645);
and U11182 (N_11182,N_10621,N_10632);
nand U11183 (N_11183,N_10775,N_10589);
nand U11184 (N_11184,N_10554,N_10955);
nand U11185 (N_11185,N_10736,N_10938);
nor U11186 (N_11186,N_10693,N_10685);
nor U11187 (N_11187,N_10586,N_10769);
xor U11188 (N_11188,N_10957,N_10924);
or U11189 (N_11189,N_10790,N_10981);
nor U11190 (N_11190,N_10536,N_10818);
and U11191 (N_11191,N_10551,N_10896);
or U11192 (N_11192,N_10797,N_10581);
nor U11193 (N_11193,N_10744,N_10684);
and U11194 (N_11194,N_10933,N_10810);
nor U11195 (N_11195,N_10557,N_10687);
or U11196 (N_11196,N_10959,N_10874);
nor U11197 (N_11197,N_10838,N_10740);
and U11198 (N_11198,N_10634,N_10970);
nand U11199 (N_11199,N_10982,N_10729);
nor U11200 (N_11200,N_10732,N_10906);
nand U11201 (N_11201,N_10604,N_10521);
and U11202 (N_11202,N_10782,N_10831);
nand U11203 (N_11203,N_10566,N_10915);
nand U11204 (N_11204,N_10602,N_10605);
nor U11205 (N_11205,N_10940,N_10738);
nor U11206 (N_11206,N_10794,N_10523);
nor U11207 (N_11207,N_10511,N_10688);
and U11208 (N_11208,N_10826,N_10780);
nand U11209 (N_11209,N_10574,N_10947);
and U11210 (N_11210,N_10932,N_10507);
nor U11211 (N_11211,N_10991,N_10758);
nand U11212 (N_11212,N_10642,N_10935);
and U11213 (N_11213,N_10962,N_10515);
or U11214 (N_11214,N_10789,N_10592);
and U11215 (N_11215,N_10722,N_10842);
or U11216 (N_11216,N_10870,N_10676);
nand U11217 (N_11217,N_10909,N_10969);
or U11218 (N_11218,N_10655,N_10848);
nor U11219 (N_11219,N_10912,N_10923);
or U11220 (N_11220,N_10746,N_10900);
nor U11221 (N_11221,N_10783,N_10560);
nor U11222 (N_11222,N_10595,N_10852);
nor U11223 (N_11223,N_10549,N_10500);
or U11224 (N_11224,N_10514,N_10749);
or U11225 (N_11225,N_10510,N_10877);
or U11226 (N_11226,N_10750,N_10730);
nor U11227 (N_11227,N_10868,N_10999);
and U11228 (N_11228,N_10585,N_10575);
xnor U11229 (N_11229,N_10614,N_10533);
xor U11230 (N_11230,N_10538,N_10891);
or U11231 (N_11231,N_10945,N_10594);
or U11232 (N_11232,N_10745,N_10739);
nand U11233 (N_11233,N_10846,N_10535);
nand U11234 (N_11234,N_10710,N_10853);
nor U11235 (N_11235,N_10803,N_10665);
nor U11236 (N_11236,N_10788,N_10762);
xor U11237 (N_11237,N_10683,N_10796);
nand U11238 (N_11238,N_10833,N_10845);
nor U11239 (N_11239,N_10606,N_10972);
nand U11240 (N_11240,N_10795,N_10863);
and U11241 (N_11241,N_10601,N_10600);
nand U11242 (N_11242,N_10694,N_10920);
and U11243 (N_11243,N_10757,N_10641);
xor U11244 (N_11244,N_10927,N_10816);
xor U11245 (N_11245,N_10570,N_10552);
xor U11246 (N_11246,N_10731,N_10943);
or U11247 (N_11247,N_10519,N_10689);
nand U11248 (N_11248,N_10934,N_10850);
or U11249 (N_11249,N_10867,N_10839);
and U11250 (N_11250,N_10678,N_10633);
or U11251 (N_11251,N_10755,N_10507);
nand U11252 (N_11252,N_10537,N_10692);
or U11253 (N_11253,N_10616,N_10575);
nor U11254 (N_11254,N_10715,N_10731);
nand U11255 (N_11255,N_10738,N_10825);
nand U11256 (N_11256,N_10571,N_10690);
xnor U11257 (N_11257,N_10849,N_10602);
xnor U11258 (N_11258,N_10618,N_10838);
xnor U11259 (N_11259,N_10527,N_10998);
nor U11260 (N_11260,N_10702,N_10770);
nand U11261 (N_11261,N_10715,N_10608);
or U11262 (N_11262,N_10718,N_10532);
nand U11263 (N_11263,N_10716,N_10907);
xor U11264 (N_11264,N_10934,N_10608);
or U11265 (N_11265,N_10958,N_10587);
nor U11266 (N_11266,N_10744,N_10842);
nor U11267 (N_11267,N_10796,N_10819);
nor U11268 (N_11268,N_10817,N_10725);
xor U11269 (N_11269,N_10990,N_10590);
or U11270 (N_11270,N_10618,N_10517);
xnor U11271 (N_11271,N_10833,N_10834);
or U11272 (N_11272,N_10702,N_10854);
or U11273 (N_11273,N_10627,N_10583);
and U11274 (N_11274,N_10965,N_10894);
xnor U11275 (N_11275,N_10785,N_10783);
and U11276 (N_11276,N_10525,N_10560);
xnor U11277 (N_11277,N_10754,N_10824);
xnor U11278 (N_11278,N_10621,N_10892);
xor U11279 (N_11279,N_10776,N_10723);
and U11280 (N_11280,N_10579,N_10680);
nor U11281 (N_11281,N_10885,N_10943);
or U11282 (N_11282,N_10872,N_10617);
and U11283 (N_11283,N_10800,N_10676);
or U11284 (N_11284,N_10979,N_10853);
nand U11285 (N_11285,N_10724,N_10591);
nor U11286 (N_11286,N_10849,N_10997);
or U11287 (N_11287,N_10607,N_10921);
nand U11288 (N_11288,N_10602,N_10698);
and U11289 (N_11289,N_10779,N_10950);
nand U11290 (N_11290,N_10808,N_10660);
nor U11291 (N_11291,N_10625,N_10566);
xor U11292 (N_11292,N_10743,N_10571);
and U11293 (N_11293,N_10667,N_10550);
xnor U11294 (N_11294,N_10753,N_10835);
and U11295 (N_11295,N_10526,N_10764);
xnor U11296 (N_11296,N_10961,N_10950);
xnor U11297 (N_11297,N_10572,N_10656);
and U11298 (N_11298,N_10591,N_10548);
nor U11299 (N_11299,N_10669,N_10905);
or U11300 (N_11300,N_10961,N_10888);
or U11301 (N_11301,N_10801,N_10766);
nand U11302 (N_11302,N_10725,N_10736);
nand U11303 (N_11303,N_10848,N_10798);
or U11304 (N_11304,N_10700,N_10958);
nor U11305 (N_11305,N_10568,N_10653);
xor U11306 (N_11306,N_10791,N_10543);
nor U11307 (N_11307,N_10931,N_10950);
and U11308 (N_11308,N_10576,N_10583);
nand U11309 (N_11309,N_10999,N_10923);
or U11310 (N_11310,N_10666,N_10984);
nand U11311 (N_11311,N_10874,N_10692);
or U11312 (N_11312,N_10762,N_10790);
nor U11313 (N_11313,N_10510,N_10682);
or U11314 (N_11314,N_10535,N_10519);
xnor U11315 (N_11315,N_10715,N_10974);
xor U11316 (N_11316,N_10586,N_10975);
nand U11317 (N_11317,N_10698,N_10529);
nand U11318 (N_11318,N_10638,N_10930);
and U11319 (N_11319,N_10627,N_10615);
nor U11320 (N_11320,N_10634,N_10784);
or U11321 (N_11321,N_10740,N_10757);
nand U11322 (N_11322,N_10866,N_10693);
and U11323 (N_11323,N_10775,N_10877);
or U11324 (N_11324,N_10785,N_10841);
or U11325 (N_11325,N_10699,N_10983);
nand U11326 (N_11326,N_10783,N_10966);
xor U11327 (N_11327,N_10509,N_10918);
xnor U11328 (N_11328,N_10962,N_10703);
or U11329 (N_11329,N_10825,N_10689);
or U11330 (N_11330,N_10986,N_10631);
nand U11331 (N_11331,N_10834,N_10714);
nor U11332 (N_11332,N_10952,N_10540);
or U11333 (N_11333,N_10981,N_10789);
nand U11334 (N_11334,N_10570,N_10860);
xor U11335 (N_11335,N_10670,N_10540);
nor U11336 (N_11336,N_10613,N_10744);
nand U11337 (N_11337,N_10923,N_10598);
or U11338 (N_11338,N_10848,N_10565);
nand U11339 (N_11339,N_10554,N_10902);
xnor U11340 (N_11340,N_10691,N_10523);
and U11341 (N_11341,N_10867,N_10739);
and U11342 (N_11342,N_10745,N_10556);
nand U11343 (N_11343,N_10627,N_10711);
xor U11344 (N_11344,N_10683,N_10755);
or U11345 (N_11345,N_10966,N_10952);
nor U11346 (N_11346,N_10571,N_10803);
or U11347 (N_11347,N_10859,N_10727);
or U11348 (N_11348,N_10574,N_10658);
nand U11349 (N_11349,N_10830,N_10831);
xnor U11350 (N_11350,N_10513,N_10832);
xor U11351 (N_11351,N_10883,N_10693);
xor U11352 (N_11352,N_10694,N_10683);
and U11353 (N_11353,N_10754,N_10833);
nor U11354 (N_11354,N_10790,N_10661);
and U11355 (N_11355,N_10517,N_10859);
nand U11356 (N_11356,N_10766,N_10759);
nand U11357 (N_11357,N_10708,N_10623);
nand U11358 (N_11358,N_10641,N_10952);
and U11359 (N_11359,N_10850,N_10836);
and U11360 (N_11360,N_10965,N_10972);
or U11361 (N_11361,N_10855,N_10595);
nor U11362 (N_11362,N_10511,N_10906);
or U11363 (N_11363,N_10819,N_10961);
xnor U11364 (N_11364,N_10886,N_10845);
xnor U11365 (N_11365,N_10547,N_10976);
xnor U11366 (N_11366,N_10727,N_10842);
or U11367 (N_11367,N_10561,N_10853);
nor U11368 (N_11368,N_10906,N_10679);
xnor U11369 (N_11369,N_10561,N_10992);
nand U11370 (N_11370,N_10897,N_10570);
and U11371 (N_11371,N_10532,N_10775);
nand U11372 (N_11372,N_10894,N_10821);
or U11373 (N_11373,N_10966,N_10857);
nand U11374 (N_11374,N_10935,N_10709);
and U11375 (N_11375,N_10846,N_10845);
and U11376 (N_11376,N_10880,N_10815);
xor U11377 (N_11377,N_10589,N_10855);
xnor U11378 (N_11378,N_10984,N_10577);
nand U11379 (N_11379,N_10818,N_10956);
and U11380 (N_11380,N_10545,N_10526);
or U11381 (N_11381,N_10785,N_10958);
xor U11382 (N_11382,N_10906,N_10878);
nand U11383 (N_11383,N_10833,N_10922);
nand U11384 (N_11384,N_10649,N_10570);
xor U11385 (N_11385,N_10926,N_10819);
xor U11386 (N_11386,N_10908,N_10777);
xor U11387 (N_11387,N_10595,N_10770);
nor U11388 (N_11388,N_10815,N_10969);
and U11389 (N_11389,N_10966,N_10536);
nor U11390 (N_11390,N_10946,N_10585);
nor U11391 (N_11391,N_10928,N_10600);
xnor U11392 (N_11392,N_10729,N_10540);
or U11393 (N_11393,N_10712,N_10564);
and U11394 (N_11394,N_10555,N_10899);
and U11395 (N_11395,N_10554,N_10563);
and U11396 (N_11396,N_10994,N_10881);
nor U11397 (N_11397,N_10703,N_10835);
or U11398 (N_11398,N_10596,N_10947);
or U11399 (N_11399,N_10896,N_10724);
xor U11400 (N_11400,N_10943,N_10899);
or U11401 (N_11401,N_10524,N_10500);
nand U11402 (N_11402,N_10798,N_10692);
nor U11403 (N_11403,N_10776,N_10908);
nor U11404 (N_11404,N_10788,N_10662);
nand U11405 (N_11405,N_10720,N_10525);
and U11406 (N_11406,N_10649,N_10774);
xor U11407 (N_11407,N_10698,N_10664);
or U11408 (N_11408,N_10966,N_10853);
or U11409 (N_11409,N_10643,N_10746);
xor U11410 (N_11410,N_10951,N_10921);
xnor U11411 (N_11411,N_10709,N_10714);
xnor U11412 (N_11412,N_10741,N_10966);
or U11413 (N_11413,N_10681,N_10506);
nor U11414 (N_11414,N_10859,N_10841);
nand U11415 (N_11415,N_10776,N_10963);
xor U11416 (N_11416,N_10730,N_10503);
and U11417 (N_11417,N_10971,N_10579);
xnor U11418 (N_11418,N_10982,N_10856);
xnor U11419 (N_11419,N_10758,N_10597);
nand U11420 (N_11420,N_10834,N_10928);
and U11421 (N_11421,N_10688,N_10650);
or U11422 (N_11422,N_10648,N_10999);
nor U11423 (N_11423,N_10792,N_10932);
or U11424 (N_11424,N_10776,N_10533);
nand U11425 (N_11425,N_10844,N_10914);
nand U11426 (N_11426,N_10915,N_10659);
and U11427 (N_11427,N_10790,N_10692);
xnor U11428 (N_11428,N_10775,N_10921);
xnor U11429 (N_11429,N_10743,N_10649);
nor U11430 (N_11430,N_10970,N_10544);
nand U11431 (N_11431,N_10646,N_10671);
and U11432 (N_11432,N_10995,N_10612);
nor U11433 (N_11433,N_10542,N_10660);
and U11434 (N_11434,N_10666,N_10615);
nand U11435 (N_11435,N_10676,N_10825);
nor U11436 (N_11436,N_10886,N_10854);
xnor U11437 (N_11437,N_10783,N_10515);
and U11438 (N_11438,N_10611,N_10898);
xor U11439 (N_11439,N_10772,N_10608);
nand U11440 (N_11440,N_10536,N_10606);
nor U11441 (N_11441,N_10827,N_10546);
nor U11442 (N_11442,N_10580,N_10924);
and U11443 (N_11443,N_10597,N_10922);
or U11444 (N_11444,N_10563,N_10635);
nor U11445 (N_11445,N_10583,N_10619);
and U11446 (N_11446,N_10737,N_10534);
nor U11447 (N_11447,N_10847,N_10522);
or U11448 (N_11448,N_10570,N_10848);
nand U11449 (N_11449,N_10871,N_10552);
nor U11450 (N_11450,N_10951,N_10689);
nand U11451 (N_11451,N_10828,N_10521);
or U11452 (N_11452,N_10632,N_10830);
or U11453 (N_11453,N_10534,N_10641);
or U11454 (N_11454,N_10983,N_10559);
or U11455 (N_11455,N_10585,N_10706);
or U11456 (N_11456,N_10975,N_10537);
and U11457 (N_11457,N_10543,N_10573);
xnor U11458 (N_11458,N_10661,N_10797);
xnor U11459 (N_11459,N_10690,N_10586);
or U11460 (N_11460,N_10814,N_10502);
or U11461 (N_11461,N_10620,N_10798);
and U11462 (N_11462,N_10983,N_10537);
or U11463 (N_11463,N_10924,N_10903);
nand U11464 (N_11464,N_10914,N_10871);
nand U11465 (N_11465,N_10797,N_10988);
xor U11466 (N_11466,N_10782,N_10673);
nor U11467 (N_11467,N_10961,N_10767);
nor U11468 (N_11468,N_10631,N_10815);
xnor U11469 (N_11469,N_10877,N_10836);
xnor U11470 (N_11470,N_10898,N_10687);
or U11471 (N_11471,N_10519,N_10715);
or U11472 (N_11472,N_10519,N_10769);
nor U11473 (N_11473,N_10685,N_10790);
nor U11474 (N_11474,N_10716,N_10604);
nor U11475 (N_11475,N_10722,N_10608);
or U11476 (N_11476,N_10871,N_10592);
xor U11477 (N_11477,N_10558,N_10658);
xor U11478 (N_11478,N_10983,N_10694);
nand U11479 (N_11479,N_10788,N_10697);
nor U11480 (N_11480,N_10538,N_10922);
xor U11481 (N_11481,N_10564,N_10831);
xnor U11482 (N_11482,N_10604,N_10813);
nor U11483 (N_11483,N_10606,N_10860);
xnor U11484 (N_11484,N_10620,N_10876);
nand U11485 (N_11485,N_10650,N_10958);
or U11486 (N_11486,N_10703,N_10931);
nand U11487 (N_11487,N_10508,N_10974);
nand U11488 (N_11488,N_10879,N_10840);
nand U11489 (N_11489,N_10595,N_10884);
nand U11490 (N_11490,N_10888,N_10817);
or U11491 (N_11491,N_10533,N_10688);
and U11492 (N_11492,N_10549,N_10947);
xnor U11493 (N_11493,N_10832,N_10753);
nor U11494 (N_11494,N_10702,N_10775);
nand U11495 (N_11495,N_10715,N_10564);
nand U11496 (N_11496,N_10922,N_10834);
nand U11497 (N_11497,N_10992,N_10921);
and U11498 (N_11498,N_10875,N_10880);
nand U11499 (N_11499,N_10954,N_10624);
xor U11500 (N_11500,N_11408,N_11300);
nand U11501 (N_11501,N_11069,N_11080);
or U11502 (N_11502,N_11227,N_11200);
nor U11503 (N_11503,N_11269,N_11073);
nand U11504 (N_11504,N_11291,N_11384);
nand U11505 (N_11505,N_11127,N_11093);
nand U11506 (N_11506,N_11433,N_11455);
nor U11507 (N_11507,N_11293,N_11456);
nor U11508 (N_11508,N_11321,N_11358);
and U11509 (N_11509,N_11474,N_11364);
or U11510 (N_11510,N_11397,N_11454);
and U11511 (N_11511,N_11261,N_11079);
or U11512 (N_11512,N_11221,N_11239);
or U11513 (N_11513,N_11262,N_11411);
or U11514 (N_11514,N_11085,N_11062);
nand U11515 (N_11515,N_11307,N_11277);
or U11516 (N_11516,N_11238,N_11254);
and U11517 (N_11517,N_11362,N_11296);
xor U11518 (N_11518,N_11025,N_11136);
xnor U11519 (N_11519,N_11383,N_11045);
nor U11520 (N_11520,N_11459,N_11491);
nand U11521 (N_11521,N_11305,N_11142);
xor U11522 (N_11522,N_11424,N_11382);
and U11523 (N_11523,N_11441,N_11077);
xnor U11524 (N_11524,N_11047,N_11048);
xnor U11525 (N_11525,N_11482,N_11286);
nor U11526 (N_11526,N_11438,N_11041);
xnor U11527 (N_11527,N_11376,N_11074);
and U11528 (N_11528,N_11309,N_11216);
xor U11529 (N_11529,N_11499,N_11380);
nor U11530 (N_11530,N_11193,N_11161);
nand U11531 (N_11531,N_11479,N_11000);
nor U11532 (N_11532,N_11234,N_11138);
nand U11533 (N_11533,N_11445,N_11325);
nor U11534 (N_11534,N_11072,N_11117);
and U11535 (N_11535,N_11279,N_11163);
and U11536 (N_11536,N_11367,N_11091);
nand U11537 (N_11537,N_11355,N_11425);
or U11538 (N_11538,N_11147,N_11359);
nor U11539 (N_11539,N_11273,N_11026);
or U11540 (N_11540,N_11164,N_11437);
or U11541 (N_11541,N_11449,N_11348);
or U11542 (N_11542,N_11143,N_11100);
nor U11543 (N_11543,N_11420,N_11385);
nand U11544 (N_11544,N_11417,N_11229);
and U11545 (N_11545,N_11061,N_11341);
and U11546 (N_11546,N_11212,N_11190);
and U11547 (N_11547,N_11219,N_11034);
or U11548 (N_11548,N_11146,N_11336);
nor U11549 (N_11549,N_11210,N_11166);
or U11550 (N_11550,N_11196,N_11337);
xor U11551 (N_11551,N_11263,N_11480);
or U11552 (N_11552,N_11063,N_11485);
or U11553 (N_11553,N_11160,N_11360);
nor U11554 (N_11554,N_11105,N_11460);
or U11555 (N_11555,N_11418,N_11039);
nor U11556 (N_11556,N_11198,N_11295);
nand U11557 (N_11557,N_11129,N_11225);
and U11558 (N_11558,N_11241,N_11096);
or U11559 (N_11559,N_11173,N_11447);
nor U11560 (N_11560,N_11444,N_11066);
nand U11561 (N_11561,N_11352,N_11020);
or U11562 (N_11562,N_11017,N_11010);
or U11563 (N_11563,N_11270,N_11426);
or U11564 (N_11564,N_11398,N_11451);
nor U11565 (N_11565,N_11400,N_11320);
nor U11566 (N_11566,N_11012,N_11244);
xor U11567 (N_11567,N_11172,N_11230);
nand U11568 (N_11568,N_11457,N_11349);
and U11569 (N_11569,N_11265,N_11264);
xnor U11570 (N_11570,N_11016,N_11285);
and U11571 (N_11571,N_11443,N_11235);
nand U11572 (N_11572,N_11363,N_11381);
or U11573 (N_11573,N_11391,N_11248);
nor U11574 (N_11574,N_11046,N_11332);
nor U11575 (N_11575,N_11159,N_11361);
nand U11576 (N_11576,N_11306,N_11316);
or U11577 (N_11577,N_11188,N_11366);
and U11578 (N_11578,N_11287,N_11171);
or U11579 (N_11579,N_11333,N_11289);
nor U11580 (N_11580,N_11496,N_11175);
and U11581 (N_11581,N_11351,N_11168);
and U11582 (N_11582,N_11106,N_11197);
or U11583 (N_11583,N_11110,N_11257);
and U11584 (N_11584,N_11242,N_11226);
and U11585 (N_11585,N_11431,N_11386);
and U11586 (N_11586,N_11374,N_11467);
xnor U11587 (N_11587,N_11463,N_11109);
and U11588 (N_11588,N_11402,N_11466);
or U11589 (N_11589,N_11208,N_11205);
and U11590 (N_11590,N_11429,N_11089);
or U11591 (N_11591,N_11038,N_11258);
or U11592 (N_11592,N_11094,N_11092);
and U11593 (N_11593,N_11036,N_11489);
or U11594 (N_11594,N_11014,N_11005);
xnor U11595 (N_11595,N_11323,N_11314);
or U11596 (N_11596,N_11107,N_11001);
or U11597 (N_11597,N_11324,N_11217);
nand U11598 (N_11598,N_11345,N_11086);
nor U11599 (N_11599,N_11412,N_11276);
xor U11600 (N_11600,N_11165,N_11095);
and U11601 (N_11601,N_11232,N_11145);
nor U11602 (N_11602,N_11315,N_11275);
xor U11603 (N_11603,N_11243,N_11344);
and U11604 (N_11604,N_11178,N_11253);
and U11605 (N_11605,N_11202,N_11013);
or U11606 (N_11606,N_11153,N_11023);
or U11607 (N_11607,N_11044,N_11304);
xor U11608 (N_11608,N_11192,N_11357);
nor U11609 (N_11609,N_11082,N_11207);
xor U11610 (N_11610,N_11169,N_11354);
and U11611 (N_11611,N_11119,N_11476);
nor U11612 (N_11612,N_11284,N_11492);
xnor U11613 (N_11613,N_11432,N_11167);
or U11614 (N_11614,N_11008,N_11179);
nand U11615 (N_11615,N_11204,N_11250);
xnor U11616 (N_11616,N_11430,N_11422);
xnor U11617 (N_11617,N_11111,N_11003);
and U11618 (N_11618,N_11371,N_11292);
and U11619 (N_11619,N_11246,N_11401);
nand U11620 (N_11620,N_11319,N_11311);
xnor U11621 (N_11621,N_11368,N_11231);
and U11622 (N_11622,N_11483,N_11203);
and U11623 (N_11623,N_11272,N_11099);
and U11624 (N_11624,N_11134,N_11211);
or U11625 (N_11625,N_11191,N_11399);
or U11626 (N_11626,N_11011,N_11084);
or U11627 (N_11627,N_11006,N_11435);
nor U11628 (N_11628,N_11494,N_11007);
xnor U11629 (N_11629,N_11313,N_11312);
xnor U11630 (N_11630,N_11021,N_11245);
nand U11631 (N_11631,N_11365,N_11050);
xor U11632 (N_11632,N_11141,N_11439);
and U11633 (N_11633,N_11068,N_11132);
nand U11634 (N_11634,N_11475,N_11108);
nor U11635 (N_11635,N_11133,N_11199);
nand U11636 (N_11636,N_11298,N_11278);
nor U11637 (N_11637,N_11326,N_11156);
or U11638 (N_11638,N_11124,N_11121);
and U11639 (N_11639,N_11015,N_11347);
and U11640 (N_11640,N_11461,N_11416);
xor U11641 (N_11641,N_11423,N_11233);
and U11642 (N_11642,N_11301,N_11083);
or U11643 (N_11643,N_11081,N_11481);
and U11644 (N_11644,N_11209,N_11058);
xnor U11645 (N_11645,N_11247,N_11155);
and U11646 (N_11646,N_11356,N_11495);
xnor U11647 (N_11647,N_11053,N_11267);
nand U11648 (N_11648,N_11260,N_11327);
nor U11649 (N_11649,N_11059,N_11158);
and U11650 (N_11650,N_11440,N_11448);
and U11651 (N_11651,N_11149,N_11252);
nor U11652 (N_11652,N_11223,N_11157);
nand U11653 (N_11653,N_11116,N_11497);
xnor U11654 (N_11654,N_11335,N_11213);
nor U11655 (N_11655,N_11101,N_11150);
xnor U11656 (N_11656,N_11346,N_11215);
and U11657 (N_11657,N_11472,N_11281);
and U11658 (N_11658,N_11427,N_11464);
and U11659 (N_11659,N_11070,N_11122);
nand U11660 (N_11660,N_11088,N_11282);
and U11661 (N_11661,N_11120,N_11436);
xnor U11662 (N_11662,N_11274,N_11404);
and U11663 (N_11663,N_11259,N_11283);
nand U11664 (N_11664,N_11033,N_11130);
nor U11665 (N_11665,N_11471,N_11114);
or U11666 (N_11666,N_11477,N_11318);
xnor U11667 (N_11667,N_11140,N_11268);
xor U11668 (N_11668,N_11465,N_11104);
xor U11669 (N_11669,N_11330,N_11018);
or U11670 (N_11670,N_11378,N_11372);
nor U11671 (N_11671,N_11396,N_11115);
or U11672 (N_11672,N_11060,N_11137);
nand U11673 (N_11673,N_11322,N_11189);
nand U11674 (N_11674,N_11098,N_11043);
or U11675 (N_11675,N_11035,N_11240);
nand U11676 (N_11676,N_11118,N_11071);
nor U11677 (N_11677,N_11487,N_11389);
nand U11678 (N_11678,N_11303,N_11373);
nand U11679 (N_11679,N_11469,N_11182);
or U11680 (N_11680,N_11379,N_11388);
or U11681 (N_11681,N_11220,N_11369);
xnor U11682 (N_11682,N_11375,N_11128);
xor U11683 (N_11683,N_11031,N_11177);
nor U11684 (N_11684,N_11452,N_11097);
and U11685 (N_11685,N_11251,N_11290);
nand U11686 (N_11686,N_11176,N_11317);
and U11687 (N_11687,N_11377,N_11308);
or U11688 (N_11688,N_11394,N_11414);
nor U11689 (N_11689,N_11334,N_11249);
nor U11690 (N_11690,N_11078,N_11022);
or U11691 (N_11691,N_11112,N_11299);
and U11692 (N_11692,N_11442,N_11067);
or U11693 (N_11693,N_11029,N_11343);
and U11694 (N_11694,N_11478,N_11113);
nand U11695 (N_11695,N_11470,N_11037);
nor U11696 (N_11696,N_11131,N_11194);
xnor U11697 (N_11697,N_11294,N_11331);
nor U11698 (N_11698,N_11135,N_11009);
or U11699 (N_11699,N_11144,N_11090);
and U11700 (N_11700,N_11087,N_11236);
nor U11701 (N_11701,N_11419,N_11490);
xnor U11702 (N_11702,N_11181,N_11288);
nor U11703 (N_11703,N_11187,N_11255);
nor U11704 (N_11704,N_11103,N_11206);
nor U11705 (N_11705,N_11409,N_11390);
nand U11706 (N_11706,N_11473,N_11428);
and U11707 (N_11707,N_11370,N_11201);
nor U11708 (N_11708,N_11004,N_11353);
or U11709 (N_11709,N_11102,N_11126);
or U11710 (N_11710,N_11055,N_11056);
nor U11711 (N_11711,N_11302,N_11256);
xor U11712 (N_11712,N_11338,N_11493);
nand U11713 (N_11713,N_11027,N_11051);
or U11714 (N_11714,N_11453,N_11075);
xnor U11715 (N_11715,N_11329,N_11183);
or U11716 (N_11716,N_11148,N_11415);
nor U11717 (N_11717,N_11151,N_11019);
and U11718 (N_11718,N_11057,N_11076);
or U11719 (N_11719,N_11468,N_11123);
nor U11720 (N_11720,N_11065,N_11186);
or U11721 (N_11721,N_11350,N_11486);
or U11722 (N_11722,N_11450,N_11214);
xor U11723 (N_11723,N_11174,N_11328);
and U11724 (N_11724,N_11340,N_11185);
and U11725 (N_11725,N_11405,N_11152);
nand U11726 (N_11726,N_11154,N_11002);
and U11727 (N_11727,N_11064,N_11406);
and U11728 (N_11728,N_11170,N_11054);
or U11729 (N_11729,N_11024,N_11032);
or U11730 (N_11730,N_11042,N_11271);
xnor U11731 (N_11731,N_11180,N_11446);
nor U11732 (N_11732,N_11434,N_11028);
or U11733 (N_11733,N_11413,N_11218);
and U11734 (N_11734,N_11339,N_11297);
nor U11735 (N_11735,N_11421,N_11403);
nor U11736 (N_11736,N_11228,N_11458);
nor U11737 (N_11737,N_11462,N_11125);
and U11738 (N_11738,N_11342,N_11387);
xnor U11739 (N_11739,N_11049,N_11237);
nand U11740 (N_11740,N_11224,N_11410);
or U11741 (N_11741,N_11040,N_11266);
xnor U11742 (N_11742,N_11052,N_11395);
nand U11743 (N_11743,N_11162,N_11310);
xnor U11744 (N_11744,N_11393,N_11030);
or U11745 (N_11745,N_11280,N_11139);
nor U11746 (N_11746,N_11392,N_11222);
or U11747 (N_11747,N_11184,N_11195);
and U11748 (N_11748,N_11488,N_11407);
xnor U11749 (N_11749,N_11498,N_11484);
nor U11750 (N_11750,N_11072,N_11010);
nor U11751 (N_11751,N_11142,N_11091);
nand U11752 (N_11752,N_11431,N_11485);
nor U11753 (N_11753,N_11187,N_11088);
nand U11754 (N_11754,N_11012,N_11230);
nand U11755 (N_11755,N_11155,N_11018);
nand U11756 (N_11756,N_11120,N_11209);
nor U11757 (N_11757,N_11142,N_11422);
or U11758 (N_11758,N_11135,N_11084);
xor U11759 (N_11759,N_11137,N_11159);
xor U11760 (N_11760,N_11388,N_11073);
or U11761 (N_11761,N_11144,N_11493);
or U11762 (N_11762,N_11322,N_11330);
nor U11763 (N_11763,N_11025,N_11011);
xor U11764 (N_11764,N_11490,N_11027);
nor U11765 (N_11765,N_11038,N_11140);
or U11766 (N_11766,N_11375,N_11242);
and U11767 (N_11767,N_11193,N_11218);
nand U11768 (N_11768,N_11113,N_11134);
or U11769 (N_11769,N_11317,N_11310);
or U11770 (N_11770,N_11365,N_11026);
nand U11771 (N_11771,N_11397,N_11244);
nand U11772 (N_11772,N_11354,N_11152);
nor U11773 (N_11773,N_11462,N_11032);
nor U11774 (N_11774,N_11216,N_11490);
xor U11775 (N_11775,N_11208,N_11429);
and U11776 (N_11776,N_11088,N_11232);
nor U11777 (N_11777,N_11004,N_11282);
xnor U11778 (N_11778,N_11022,N_11373);
nand U11779 (N_11779,N_11196,N_11181);
xor U11780 (N_11780,N_11156,N_11158);
and U11781 (N_11781,N_11304,N_11263);
nand U11782 (N_11782,N_11433,N_11434);
or U11783 (N_11783,N_11323,N_11122);
and U11784 (N_11784,N_11088,N_11330);
nor U11785 (N_11785,N_11326,N_11080);
nor U11786 (N_11786,N_11303,N_11228);
or U11787 (N_11787,N_11078,N_11332);
nor U11788 (N_11788,N_11165,N_11496);
and U11789 (N_11789,N_11419,N_11113);
nand U11790 (N_11790,N_11460,N_11380);
or U11791 (N_11791,N_11288,N_11295);
or U11792 (N_11792,N_11294,N_11479);
or U11793 (N_11793,N_11176,N_11265);
and U11794 (N_11794,N_11331,N_11348);
nor U11795 (N_11795,N_11489,N_11105);
nand U11796 (N_11796,N_11090,N_11121);
nor U11797 (N_11797,N_11298,N_11075);
xor U11798 (N_11798,N_11448,N_11299);
and U11799 (N_11799,N_11214,N_11213);
and U11800 (N_11800,N_11013,N_11426);
nor U11801 (N_11801,N_11242,N_11382);
nor U11802 (N_11802,N_11037,N_11347);
xor U11803 (N_11803,N_11053,N_11387);
nand U11804 (N_11804,N_11307,N_11330);
and U11805 (N_11805,N_11080,N_11472);
xnor U11806 (N_11806,N_11062,N_11445);
nand U11807 (N_11807,N_11411,N_11166);
nor U11808 (N_11808,N_11175,N_11381);
and U11809 (N_11809,N_11284,N_11241);
nand U11810 (N_11810,N_11202,N_11029);
and U11811 (N_11811,N_11289,N_11389);
nor U11812 (N_11812,N_11168,N_11043);
and U11813 (N_11813,N_11257,N_11289);
and U11814 (N_11814,N_11459,N_11174);
nand U11815 (N_11815,N_11057,N_11175);
nor U11816 (N_11816,N_11226,N_11498);
nor U11817 (N_11817,N_11318,N_11437);
nand U11818 (N_11818,N_11288,N_11419);
nor U11819 (N_11819,N_11473,N_11108);
nor U11820 (N_11820,N_11014,N_11001);
nor U11821 (N_11821,N_11453,N_11057);
nand U11822 (N_11822,N_11178,N_11328);
xnor U11823 (N_11823,N_11331,N_11360);
nand U11824 (N_11824,N_11011,N_11364);
nand U11825 (N_11825,N_11161,N_11022);
nor U11826 (N_11826,N_11136,N_11314);
xor U11827 (N_11827,N_11442,N_11448);
nand U11828 (N_11828,N_11100,N_11240);
xnor U11829 (N_11829,N_11199,N_11340);
and U11830 (N_11830,N_11158,N_11159);
xor U11831 (N_11831,N_11054,N_11010);
or U11832 (N_11832,N_11205,N_11378);
or U11833 (N_11833,N_11483,N_11284);
nor U11834 (N_11834,N_11449,N_11051);
nor U11835 (N_11835,N_11060,N_11450);
nor U11836 (N_11836,N_11327,N_11042);
and U11837 (N_11837,N_11419,N_11213);
xnor U11838 (N_11838,N_11488,N_11188);
or U11839 (N_11839,N_11403,N_11054);
and U11840 (N_11840,N_11272,N_11305);
xnor U11841 (N_11841,N_11322,N_11147);
or U11842 (N_11842,N_11021,N_11013);
nor U11843 (N_11843,N_11491,N_11001);
nand U11844 (N_11844,N_11271,N_11232);
nand U11845 (N_11845,N_11355,N_11030);
nand U11846 (N_11846,N_11013,N_11397);
nor U11847 (N_11847,N_11119,N_11379);
or U11848 (N_11848,N_11242,N_11039);
nor U11849 (N_11849,N_11074,N_11445);
or U11850 (N_11850,N_11292,N_11394);
or U11851 (N_11851,N_11384,N_11352);
or U11852 (N_11852,N_11391,N_11015);
or U11853 (N_11853,N_11226,N_11467);
xor U11854 (N_11854,N_11258,N_11014);
nand U11855 (N_11855,N_11092,N_11459);
nand U11856 (N_11856,N_11435,N_11094);
or U11857 (N_11857,N_11324,N_11035);
nor U11858 (N_11858,N_11322,N_11433);
or U11859 (N_11859,N_11332,N_11238);
xor U11860 (N_11860,N_11227,N_11309);
xnor U11861 (N_11861,N_11322,N_11313);
nand U11862 (N_11862,N_11112,N_11071);
nor U11863 (N_11863,N_11426,N_11174);
or U11864 (N_11864,N_11146,N_11253);
nand U11865 (N_11865,N_11410,N_11036);
nand U11866 (N_11866,N_11114,N_11238);
nand U11867 (N_11867,N_11270,N_11179);
nand U11868 (N_11868,N_11272,N_11156);
xnor U11869 (N_11869,N_11110,N_11363);
and U11870 (N_11870,N_11451,N_11386);
or U11871 (N_11871,N_11015,N_11379);
nor U11872 (N_11872,N_11367,N_11290);
xor U11873 (N_11873,N_11385,N_11036);
and U11874 (N_11874,N_11270,N_11358);
nand U11875 (N_11875,N_11213,N_11026);
xor U11876 (N_11876,N_11370,N_11434);
nand U11877 (N_11877,N_11312,N_11045);
nand U11878 (N_11878,N_11382,N_11482);
xnor U11879 (N_11879,N_11216,N_11253);
and U11880 (N_11880,N_11266,N_11260);
xor U11881 (N_11881,N_11453,N_11331);
and U11882 (N_11882,N_11253,N_11498);
xnor U11883 (N_11883,N_11164,N_11447);
xnor U11884 (N_11884,N_11478,N_11397);
xnor U11885 (N_11885,N_11484,N_11417);
xnor U11886 (N_11886,N_11011,N_11095);
xnor U11887 (N_11887,N_11350,N_11106);
xor U11888 (N_11888,N_11115,N_11374);
nand U11889 (N_11889,N_11195,N_11213);
nor U11890 (N_11890,N_11322,N_11373);
xnor U11891 (N_11891,N_11036,N_11026);
nand U11892 (N_11892,N_11266,N_11129);
and U11893 (N_11893,N_11356,N_11445);
nand U11894 (N_11894,N_11424,N_11155);
xnor U11895 (N_11895,N_11286,N_11423);
nor U11896 (N_11896,N_11226,N_11091);
nand U11897 (N_11897,N_11237,N_11397);
xnor U11898 (N_11898,N_11000,N_11344);
or U11899 (N_11899,N_11172,N_11218);
or U11900 (N_11900,N_11208,N_11049);
or U11901 (N_11901,N_11096,N_11225);
or U11902 (N_11902,N_11445,N_11160);
or U11903 (N_11903,N_11142,N_11113);
nand U11904 (N_11904,N_11378,N_11142);
xnor U11905 (N_11905,N_11351,N_11035);
or U11906 (N_11906,N_11361,N_11394);
nand U11907 (N_11907,N_11298,N_11246);
nand U11908 (N_11908,N_11169,N_11496);
xnor U11909 (N_11909,N_11017,N_11109);
and U11910 (N_11910,N_11192,N_11394);
and U11911 (N_11911,N_11207,N_11128);
or U11912 (N_11912,N_11333,N_11109);
xnor U11913 (N_11913,N_11248,N_11089);
or U11914 (N_11914,N_11452,N_11212);
nor U11915 (N_11915,N_11137,N_11224);
or U11916 (N_11916,N_11355,N_11001);
and U11917 (N_11917,N_11134,N_11337);
nand U11918 (N_11918,N_11074,N_11416);
and U11919 (N_11919,N_11294,N_11033);
xnor U11920 (N_11920,N_11372,N_11233);
xor U11921 (N_11921,N_11324,N_11255);
nor U11922 (N_11922,N_11171,N_11020);
nand U11923 (N_11923,N_11054,N_11198);
nand U11924 (N_11924,N_11028,N_11338);
xor U11925 (N_11925,N_11005,N_11373);
and U11926 (N_11926,N_11488,N_11376);
or U11927 (N_11927,N_11275,N_11288);
nor U11928 (N_11928,N_11290,N_11193);
nand U11929 (N_11929,N_11338,N_11389);
nor U11930 (N_11930,N_11481,N_11318);
xor U11931 (N_11931,N_11161,N_11353);
nand U11932 (N_11932,N_11489,N_11259);
and U11933 (N_11933,N_11266,N_11360);
nor U11934 (N_11934,N_11447,N_11118);
nor U11935 (N_11935,N_11152,N_11404);
nand U11936 (N_11936,N_11461,N_11125);
xnor U11937 (N_11937,N_11040,N_11051);
and U11938 (N_11938,N_11111,N_11456);
nand U11939 (N_11939,N_11297,N_11184);
or U11940 (N_11940,N_11047,N_11035);
and U11941 (N_11941,N_11245,N_11066);
or U11942 (N_11942,N_11377,N_11423);
and U11943 (N_11943,N_11449,N_11426);
nand U11944 (N_11944,N_11387,N_11009);
or U11945 (N_11945,N_11311,N_11236);
nor U11946 (N_11946,N_11199,N_11338);
nor U11947 (N_11947,N_11052,N_11224);
xor U11948 (N_11948,N_11395,N_11098);
nor U11949 (N_11949,N_11391,N_11335);
nor U11950 (N_11950,N_11003,N_11282);
or U11951 (N_11951,N_11348,N_11306);
xor U11952 (N_11952,N_11177,N_11033);
and U11953 (N_11953,N_11371,N_11454);
nor U11954 (N_11954,N_11094,N_11409);
xnor U11955 (N_11955,N_11021,N_11390);
and U11956 (N_11956,N_11236,N_11156);
or U11957 (N_11957,N_11129,N_11316);
and U11958 (N_11958,N_11069,N_11286);
xor U11959 (N_11959,N_11391,N_11343);
or U11960 (N_11960,N_11279,N_11392);
and U11961 (N_11961,N_11423,N_11082);
nor U11962 (N_11962,N_11046,N_11486);
or U11963 (N_11963,N_11158,N_11313);
nand U11964 (N_11964,N_11371,N_11030);
and U11965 (N_11965,N_11472,N_11101);
and U11966 (N_11966,N_11015,N_11206);
nor U11967 (N_11967,N_11213,N_11263);
or U11968 (N_11968,N_11021,N_11172);
and U11969 (N_11969,N_11145,N_11170);
nand U11970 (N_11970,N_11359,N_11048);
xor U11971 (N_11971,N_11358,N_11181);
xor U11972 (N_11972,N_11185,N_11415);
xnor U11973 (N_11973,N_11064,N_11358);
nor U11974 (N_11974,N_11460,N_11476);
nor U11975 (N_11975,N_11390,N_11349);
or U11976 (N_11976,N_11033,N_11049);
or U11977 (N_11977,N_11376,N_11068);
nand U11978 (N_11978,N_11121,N_11476);
nor U11979 (N_11979,N_11163,N_11479);
xor U11980 (N_11980,N_11406,N_11273);
nand U11981 (N_11981,N_11245,N_11283);
or U11982 (N_11982,N_11083,N_11295);
and U11983 (N_11983,N_11494,N_11246);
nand U11984 (N_11984,N_11447,N_11320);
and U11985 (N_11985,N_11448,N_11328);
xnor U11986 (N_11986,N_11316,N_11158);
nand U11987 (N_11987,N_11014,N_11245);
and U11988 (N_11988,N_11105,N_11309);
nor U11989 (N_11989,N_11077,N_11407);
nor U11990 (N_11990,N_11076,N_11301);
and U11991 (N_11991,N_11047,N_11213);
or U11992 (N_11992,N_11240,N_11304);
nand U11993 (N_11993,N_11422,N_11381);
and U11994 (N_11994,N_11389,N_11290);
nand U11995 (N_11995,N_11118,N_11135);
and U11996 (N_11996,N_11324,N_11172);
xor U11997 (N_11997,N_11359,N_11320);
nor U11998 (N_11998,N_11292,N_11297);
nor U11999 (N_11999,N_11373,N_11284);
or U12000 (N_12000,N_11740,N_11604);
or U12001 (N_12001,N_11592,N_11571);
and U12002 (N_12002,N_11936,N_11515);
and U12003 (N_12003,N_11827,N_11676);
nor U12004 (N_12004,N_11645,N_11682);
nor U12005 (N_12005,N_11999,N_11848);
and U12006 (N_12006,N_11883,N_11823);
xnor U12007 (N_12007,N_11739,N_11991);
xor U12008 (N_12008,N_11754,N_11553);
nor U12009 (N_12009,N_11766,N_11889);
nand U12010 (N_12010,N_11967,N_11620);
nand U12011 (N_12011,N_11598,N_11583);
or U12012 (N_12012,N_11954,N_11965);
nand U12013 (N_12013,N_11862,N_11916);
xor U12014 (N_12014,N_11536,N_11810);
and U12015 (N_12015,N_11556,N_11863);
nor U12016 (N_12016,N_11730,N_11542);
xnor U12017 (N_12017,N_11885,N_11517);
nand U12018 (N_12018,N_11993,N_11792);
xor U12019 (N_12019,N_11656,N_11821);
or U12020 (N_12020,N_11910,N_11623);
xor U12021 (N_12021,N_11669,N_11909);
xnor U12022 (N_12022,N_11752,N_11962);
or U12023 (N_12023,N_11973,N_11717);
or U12024 (N_12024,N_11902,N_11537);
nor U12025 (N_12025,N_11933,N_11950);
or U12026 (N_12026,N_11624,N_11778);
nand U12027 (N_12027,N_11619,N_11771);
nand U12028 (N_12028,N_11968,N_11648);
nor U12029 (N_12029,N_11704,N_11622);
nor U12030 (N_12030,N_11797,N_11731);
xnor U12031 (N_12031,N_11798,N_11837);
and U12032 (N_12032,N_11805,N_11928);
nor U12033 (N_12033,N_11599,N_11690);
nor U12034 (N_12034,N_11728,N_11847);
nor U12035 (N_12035,N_11667,N_11943);
nand U12036 (N_12036,N_11759,N_11737);
xnor U12037 (N_12037,N_11666,N_11784);
nand U12038 (N_12038,N_11813,N_11744);
nand U12039 (N_12039,N_11932,N_11998);
or U12040 (N_12040,N_11660,N_11977);
nor U12041 (N_12041,N_11531,N_11650);
and U12042 (N_12042,N_11939,N_11670);
xnor U12043 (N_12043,N_11736,N_11819);
xnor U12044 (N_12044,N_11538,N_11637);
xnor U12045 (N_12045,N_11567,N_11591);
or U12046 (N_12046,N_11795,N_11985);
nor U12047 (N_12047,N_11868,N_11516);
nand U12048 (N_12048,N_11816,N_11698);
or U12049 (N_12049,N_11716,N_11590);
and U12050 (N_12050,N_11651,N_11755);
nor U12051 (N_12051,N_11643,N_11652);
and U12052 (N_12052,N_11842,N_11647);
nor U12053 (N_12053,N_11694,N_11904);
nor U12054 (N_12054,N_11680,N_11509);
nand U12055 (N_12055,N_11812,N_11629);
nor U12056 (N_12056,N_11763,N_11701);
nor U12057 (N_12057,N_11794,N_11958);
nand U12058 (N_12058,N_11979,N_11709);
and U12059 (N_12059,N_11757,N_11760);
and U12060 (N_12060,N_11636,N_11508);
xnor U12061 (N_12061,N_11844,N_11984);
and U12062 (N_12062,N_11549,N_11743);
nor U12063 (N_12063,N_11751,N_11606);
or U12064 (N_12064,N_11955,N_11836);
xnor U12065 (N_12065,N_11513,N_11864);
nor U12066 (N_12066,N_11918,N_11673);
and U12067 (N_12067,N_11887,N_11773);
or U12068 (N_12068,N_11859,N_11746);
xor U12069 (N_12069,N_11775,N_11870);
xor U12070 (N_12070,N_11603,N_11845);
xnor U12071 (N_12071,N_11996,N_11687);
xor U12072 (N_12072,N_11785,N_11614);
and U12073 (N_12073,N_11693,N_11634);
xnor U12074 (N_12074,N_11725,N_11576);
and U12075 (N_12075,N_11846,N_11663);
or U12076 (N_12076,N_11871,N_11877);
or U12077 (N_12077,N_11559,N_11723);
nand U12078 (N_12078,N_11500,N_11920);
and U12079 (N_12079,N_11702,N_11849);
or U12080 (N_12080,N_11609,N_11897);
nor U12081 (N_12081,N_11899,N_11886);
or U12082 (N_12082,N_11511,N_11807);
xor U12083 (N_12083,N_11913,N_11679);
or U12084 (N_12084,N_11712,N_11817);
and U12085 (N_12085,N_11681,N_11608);
xnor U12086 (N_12086,N_11654,N_11952);
and U12087 (N_12087,N_11653,N_11944);
nand U12088 (N_12088,N_11878,N_11640);
and U12089 (N_12089,N_11986,N_11708);
nand U12090 (N_12090,N_11523,N_11957);
or U12091 (N_12091,N_11724,N_11808);
nor U12092 (N_12092,N_11930,N_11856);
or U12093 (N_12093,N_11529,N_11796);
nor U12094 (N_12094,N_11664,N_11830);
nand U12095 (N_12095,N_11748,N_11940);
xnor U12096 (N_12096,N_11722,N_11615);
or U12097 (N_12097,N_11988,N_11564);
nand U12098 (N_12098,N_11526,N_11860);
xnor U12099 (N_12099,N_11533,N_11658);
xor U12100 (N_12100,N_11747,N_11544);
or U12101 (N_12101,N_11926,N_11970);
or U12102 (N_12102,N_11600,N_11700);
xnor U12103 (N_12103,N_11912,N_11601);
nor U12104 (N_12104,N_11927,N_11554);
and U12105 (N_12105,N_11602,N_11732);
or U12106 (N_12106,N_11937,N_11616);
or U12107 (N_12107,N_11978,N_11678);
nor U12108 (N_12108,N_11688,N_11857);
nand U12109 (N_12109,N_11689,N_11677);
nand U12110 (N_12110,N_11776,N_11947);
nand U12111 (N_12111,N_11911,N_11834);
nor U12112 (N_12112,N_11990,N_11506);
and U12113 (N_12113,N_11777,N_11512);
nor U12114 (N_12114,N_11642,N_11545);
nor U12115 (N_12115,N_11815,N_11605);
xnor U12116 (N_12116,N_11575,N_11803);
and U12117 (N_12117,N_11518,N_11983);
and U12118 (N_12118,N_11935,N_11586);
and U12119 (N_12119,N_11853,N_11980);
xor U12120 (N_12120,N_11535,N_11555);
xor U12121 (N_12121,N_11800,N_11665);
nand U12122 (N_12122,N_11649,N_11662);
xor U12123 (N_12123,N_11668,N_11753);
and U12124 (N_12124,N_11595,N_11633);
and U12125 (N_12125,N_11691,N_11675);
or U12126 (N_12126,N_11729,N_11561);
nor U12127 (N_12127,N_11560,N_11908);
and U12128 (N_12128,N_11964,N_11971);
nand U12129 (N_12129,N_11593,N_11657);
nor U12130 (N_12130,N_11987,N_11925);
and U12131 (N_12131,N_11949,N_11762);
nor U12132 (N_12132,N_11894,N_11696);
xnor U12133 (N_12133,N_11901,N_11749);
or U12134 (N_12134,N_11788,N_11541);
nand U12135 (N_12135,N_11635,N_11626);
nor U12136 (N_12136,N_11697,N_11850);
nor U12137 (N_12137,N_11764,N_11934);
nor U12138 (N_12138,N_11822,N_11630);
or U12139 (N_12139,N_11825,N_11532);
nor U12140 (N_12140,N_11644,N_11770);
xnor U12141 (N_12141,N_11869,N_11976);
and U12142 (N_12142,N_11574,N_11876);
xnor U12143 (N_12143,N_11915,N_11809);
or U12144 (N_12144,N_11966,N_11563);
and U12145 (N_12145,N_11997,N_11631);
or U12146 (N_12146,N_11782,N_11922);
nand U12147 (N_12147,N_11896,N_11941);
nor U12148 (N_12148,N_11893,N_11588);
or U12149 (N_12149,N_11641,N_11946);
or U12150 (N_12150,N_11585,N_11741);
or U12151 (N_12151,N_11914,N_11613);
nand U12152 (N_12152,N_11761,N_11982);
xor U12153 (N_12153,N_11921,N_11738);
xnor U12154 (N_12154,N_11562,N_11661);
or U12155 (N_12155,N_11875,N_11811);
nor U12156 (N_12156,N_11907,N_11838);
or U12157 (N_12157,N_11750,N_11992);
or U12158 (N_12158,N_11519,N_11557);
xnor U12159 (N_12159,N_11975,N_11938);
nand U12160 (N_12160,N_11715,N_11745);
nand U12161 (N_12161,N_11948,N_11981);
xnor U12162 (N_12162,N_11628,N_11565);
and U12163 (N_12163,N_11772,N_11727);
and U12164 (N_12164,N_11799,N_11735);
nand U12165 (N_12165,N_11801,N_11706);
or U12166 (N_12166,N_11956,N_11524);
or U12167 (N_12167,N_11521,N_11610);
and U12168 (N_12168,N_11787,N_11852);
xor U12169 (N_12169,N_11843,N_11632);
nand U12170 (N_12170,N_11995,N_11572);
xnor U12171 (N_12171,N_11802,N_11703);
or U12172 (N_12172,N_11833,N_11924);
or U12173 (N_12173,N_11683,N_11734);
and U12174 (N_12174,N_11530,N_11768);
nand U12175 (N_12175,N_11959,N_11726);
nor U12176 (N_12176,N_11550,N_11905);
or U12177 (N_12177,N_11969,N_11573);
or U12178 (N_12178,N_11758,N_11718);
or U12179 (N_12179,N_11655,N_11522);
xor U12180 (N_12180,N_11820,N_11818);
nand U12181 (N_12181,N_11510,N_11791);
and U12182 (N_12182,N_11612,N_11552);
or U12183 (N_12183,N_11919,N_11742);
nor U12184 (N_12184,N_11617,N_11534);
and U12185 (N_12185,N_11994,N_11890);
nand U12186 (N_12186,N_11793,N_11923);
nand U12187 (N_12187,N_11929,N_11504);
nor U12188 (N_12188,N_11597,N_11826);
nor U12189 (N_12189,N_11774,N_11547);
or U12190 (N_12190,N_11972,N_11874);
nor U12191 (N_12191,N_11780,N_11814);
xnor U12192 (N_12192,N_11607,N_11866);
nand U12193 (N_12193,N_11721,N_11945);
nand U12194 (N_12194,N_11960,N_11942);
nor U12195 (N_12195,N_11895,N_11841);
and U12196 (N_12196,N_11539,N_11618);
and U12197 (N_12197,N_11828,N_11882);
nand U12198 (N_12198,N_11543,N_11646);
nand U12199 (N_12199,N_11711,N_11756);
nor U12200 (N_12200,N_11831,N_11900);
xor U12201 (N_12201,N_11596,N_11570);
and U12202 (N_12202,N_11625,N_11580);
nand U12203 (N_12203,N_11963,N_11581);
and U12204 (N_12204,N_11527,N_11507);
nor U12205 (N_12205,N_11769,N_11551);
xor U12206 (N_12206,N_11525,N_11790);
and U12207 (N_12207,N_11733,N_11783);
or U12208 (N_12208,N_11514,N_11858);
nor U12209 (N_12209,N_11638,N_11873);
nor U12210 (N_12210,N_11824,N_11705);
nor U12211 (N_12211,N_11579,N_11587);
nor U12212 (N_12212,N_11851,N_11906);
and U12213 (N_12213,N_11714,N_11854);
nor U12214 (N_12214,N_11898,N_11707);
or U12215 (N_12215,N_11710,N_11781);
nand U12216 (N_12216,N_11582,N_11953);
xor U12217 (N_12217,N_11888,N_11502);
or U12218 (N_12218,N_11686,N_11713);
and U12219 (N_12219,N_11584,N_11884);
or U12220 (N_12220,N_11594,N_11855);
or U12221 (N_12221,N_11589,N_11867);
and U12222 (N_12222,N_11558,N_11505);
nand U12223 (N_12223,N_11577,N_11872);
nor U12224 (N_12224,N_11892,N_11684);
xnor U12225 (N_12225,N_11720,N_11528);
nor U12226 (N_12226,N_11659,N_11840);
nand U12227 (N_12227,N_11779,N_11503);
xnor U12228 (N_12228,N_11765,N_11829);
and U12229 (N_12229,N_11695,N_11520);
nand U12230 (N_12230,N_11578,N_11839);
xor U12231 (N_12231,N_11917,N_11789);
nand U12232 (N_12232,N_11672,N_11767);
xor U12233 (N_12233,N_11692,N_11611);
or U12234 (N_12234,N_11566,N_11951);
xor U12235 (N_12235,N_11546,N_11699);
xor U12236 (N_12236,N_11639,N_11989);
or U12237 (N_12237,N_11548,N_11903);
nor U12238 (N_12238,N_11627,N_11880);
or U12239 (N_12239,N_11879,N_11804);
and U12240 (N_12240,N_11568,N_11806);
xor U12241 (N_12241,N_11674,N_11961);
xnor U12242 (N_12242,N_11540,N_11786);
xnor U12243 (N_12243,N_11891,N_11861);
xor U12244 (N_12244,N_11719,N_11974);
nor U12245 (N_12245,N_11865,N_11835);
xnor U12246 (N_12246,N_11569,N_11881);
nand U12247 (N_12247,N_11931,N_11621);
xor U12248 (N_12248,N_11671,N_11501);
nor U12249 (N_12249,N_11685,N_11832);
and U12250 (N_12250,N_11996,N_11539);
xnor U12251 (N_12251,N_11576,N_11545);
nor U12252 (N_12252,N_11707,N_11704);
or U12253 (N_12253,N_11512,N_11714);
or U12254 (N_12254,N_11554,N_11854);
nor U12255 (N_12255,N_11866,N_11685);
or U12256 (N_12256,N_11725,N_11760);
nand U12257 (N_12257,N_11624,N_11586);
nor U12258 (N_12258,N_11875,N_11987);
nand U12259 (N_12259,N_11689,N_11656);
nor U12260 (N_12260,N_11527,N_11765);
nor U12261 (N_12261,N_11818,N_11935);
or U12262 (N_12262,N_11554,N_11977);
nand U12263 (N_12263,N_11712,N_11982);
nor U12264 (N_12264,N_11864,N_11520);
and U12265 (N_12265,N_11734,N_11925);
and U12266 (N_12266,N_11756,N_11586);
nand U12267 (N_12267,N_11932,N_11609);
xnor U12268 (N_12268,N_11847,N_11549);
and U12269 (N_12269,N_11953,N_11946);
nor U12270 (N_12270,N_11718,N_11759);
or U12271 (N_12271,N_11911,N_11764);
nand U12272 (N_12272,N_11583,N_11934);
or U12273 (N_12273,N_11746,N_11909);
nor U12274 (N_12274,N_11899,N_11746);
xnor U12275 (N_12275,N_11707,N_11765);
nor U12276 (N_12276,N_11837,N_11856);
nand U12277 (N_12277,N_11845,N_11866);
and U12278 (N_12278,N_11975,N_11959);
nand U12279 (N_12279,N_11763,N_11780);
nor U12280 (N_12280,N_11737,N_11960);
and U12281 (N_12281,N_11703,N_11549);
nand U12282 (N_12282,N_11734,N_11915);
xor U12283 (N_12283,N_11684,N_11989);
or U12284 (N_12284,N_11778,N_11599);
nand U12285 (N_12285,N_11810,N_11719);
and U12286 (N_12286,N_11577,N_11602);
and U12287 (N_12287,N_11539,N_11655);
nor U12288 (N_12288,N_11679,N_11980);
nand U12289 (N_12289,N_11566,N_11761);
nor U12290 (N_12290,N_11507,N_11677);
xnor U12291 (N_12291,N_11682,N_11553);
nand U12292 (N_12292,N_11718,N_11648);
and U12293 (N_12293,N_11867,N_11615);
or U12294 (N_12294,N_11600,N_11871);
xor U12295 (N_12295,N_11793,N_11859);
xnor U12296 (N_12296,N_11682,N_11777);
or U12297 (N_12297,N_11803,N_11655);
nand U12298 (N_12298,N_11607,N_11829);
and U12299 (N_12299,N_11888,N_11510);
or U12300 (N_12300,N_11626,N_11930);
and U12301 (N_12301,N_11826,N_11659);
and U12302 (N_12302,N_11500,N_11855);
or U12303 (N_12303,N_11816,N_11837);
nor U12304 (N_12304,N_11524,N_11949);
or U12305 (N_12305,N_11597,N_11596);
and U12306 (N_12306,N_11543,N_11542);
xor U12307 (N_12307,N_11822,N_11525);
or U12308 (N_12308,N_11652,N_11948);
nand U12309 (N_12309,N_11924,N_11902);
xor U12310 (N_12310,N_11637,N_11784);
nor U12311 (N_12311,N_11662,N_11541);
xnor U12312 (N_12312,N_11561,N_11920);
or U12313 (N_12313,N_11752,N_11805);
xor U12314 (N_12314,N_11956,N_11591);
and U12315 (N_12315,N_11657,N_11800);
nor U12316 (N_12316,N_11527,N_11868);
nand U12317 (N_12317,N_11654,N_11622);
xor U12318 (N_12318,N_11784,N_11697);
nand U12319 (N_12319,N_11599,N_11741);
xnor U12320 (N_12320,N_11981,N_11767);
nand U12321 (N_12321,N_11986,N_11644);
xnor U12322 (N_12322,N_11612,N_11907);
nand U12323 (N_12323,N_11509,N_11916);
xor U12324 (N_12324,N_11516,N_11541);
xor U12325 (N_12325,N_11640,N_11660);
xnor U12326 (N_12326,N_11534,N_11585);
and U12327 (N_12327,N_11826,N_11647);
or U12328 (N_12328,N_11669,N_11834);
or U12329 (N_12329,N_11782,N_11623);
nor U12330 (N_12330,N_11714,N_11822);
nor U12331 (N_12331,N_11924,N_11669);
nor U12332 (N_12332,N_11817,N_11883);
xnor U12333 (N_12333,N_11934,N_11526);
nand U12334 (N_12334,N_11710,N_11532);
nand U12335 (N_12335,N_11571,N_11560);
or U12336 (N_12336,N_11751,N_11906);
or U12337 (N_12337,N_11576,N_11748);
and U12338 (N_12338,N_11560,N_11569);
and U12339 (N_12339,N_11726,N_11962);
nand U12340 (N_12340,N_11897,N_11785);
xor U12341 (N_12341,N_11872,N_11957);
or U12342 (N_12342,N_11831,N_11889);
nor U12343 (N_12343,N_11973,N_11931);
and U12344 (N_12344,N_11770,N_11937);
nor U12345 (N_12345,N_11574,N_11575);
nor U12346 (N_12346,N_11943,N_11949);
xnor U12347 (N_12347,N_11634,N_11993);
nor U12348 (N_12348,N_11528,N_11813);
or U12349 (N_12349,N_11702,N_11892);
and U12350 (N_12350,N_11655,N_11790);
or U12351 (N_12351,N_11506,N_11914);
nor U12352 (N_12352,N_11693,N_11604);
nor U12353 (N_12353,N_11920,N_11841);
nor U12354 (N_12354,N_11790,N_11637);
or U12355 (N_12355,N_11638,N_11999);
xor U12356 (N_12356,N_11708,N_11682);
xnor U12357 (N_12357,N_11526,N_11838);
and U12358 (N_12358,N_11979,N_11743);
nand U12359 (N_12359,N_11594,N_11758);
nor U12360 (N_12360,N_11616,N_11954);
and U12361 (N_12361,N_11910,N_11921);
xnor U12362 (N_12362,N_11750,N_11588);
nand U12363 (N_12363,N_11551,N_11973);
xor U12364 (N_12364,N_11710,N_11521);
nand U12365 (N_12365,N_11684,N_11596);
or U12366 (N_12366,N_11697,N_11978);
nand U12367 (N_12367,N_11569,N_11791);
nand U12368 (N_12368,N_11571,N_11833);
or U12369 (N_12369,N_11837,N_11700);
xor U12370 (N_12370,N_11648,N_11760);
or U12371 (N_12371,N_11642,N_11500);
xnor U12372 (N_12372,N_11911,N_11541);
or U12373 (N_12373,N_11879,N_11587);
nand U12374 (N_12374,N_11790,N_11731);
nand U12375 (N_12375,N_11912,N_11933);
and U12376 (N_12376,N_11673,N_11787);
nand U12377 (N_12377,N_11733,N_11544);
and U12378 (N_12378,N_11640,N_11914);
xor U12379 (N_12379,N_11674,N_11856);
nor U12380 (N_12380,N_11810,N_11677);
nor U12381 (N_12381,N_11796,N_11701);
nor U12382 (N_12382,N_11950,N_11554);
xor U12383 (N_12383,N_11759,N_11684);
or U12384 (N_12384,N_11867,N_11894);
or U12385 (N_12385,N_11529,N_11916);
nor U12386 (N_12386,N_11966,N_11904);
nand U12387 (N_12387,N_11958,N_11620);
xor U12388 (N_12388,N_11656,N_11717);
nand U12389 (N_12389,N_11805,N_11595);
xnor U12390 (N_12390,N_11698,N_11639);
xor U12391 (N_12391,N_11887,N_11863);
nor U12392 (N_12392,N_11686,N_11733);
nand U12393 (N_12393,N_11959,N_11904);
nor U12394 (N_12394,N_11522,N_11846);
nand U12395 (N_12395,N_11689,N_11737);
nor U12396 (N_12396,N_11705,N_11649);
xor U12397 (N_12397,N_11539,N_11729);
xnor U12398 (N_12398,N_11664,N_11808);
nor U12399 (N_12399,N_11634,N_11500);
xnor U12400 (N_12400,N_11585,N_11974);
xor U12401 (N_12401,N_11866,N_11581);
and U12402 (N_12402,N_11639,N_11501);
xnor U12403 (N_12403,N_11663,N_11939);
and U12404 (N_12404,N_11531,N_11779);
or U12405 (N_12405,N_11616,N_11855);
and U12406 (N_12406,N_11628,N_11907);
nand U12407 (N_12407,N_11579,N_11616);
or U12408 (N_12408,N_11912,N_11749);
and U12409 (N_12409,N_11566,N_11721);
nor U12410 (N_12410,N_11659,N_11870);
nor U12411 (N_12411,N_11663,N_11712);
nor U12412 (N_12412,N_11779,N_11660);
xnor U12413 (N_12413,N_11540,N_11690);
and U12414 (N_12414,N_11606,N_11708);
nand U12415 (N_12415,N_11673,N_11595);
and U12416 (N_12416,N_11685,N_11701);
nor U12417 (N_12417,N_11627,N_11958);
or U12418 (N_12418,N_11784,N_11762);
nor U12419 (N_12419,N_11531,N_11987);
or U12420 (N_12420,N_11517,N_11608);
or U12421 (N_12421,N_11912,N_11890);
nor U12422 (N_12422,N_11856,N_11605);
or U12423 (N_12423,N_11509,N_11644);
nand U12424 (N_12424,N_11750,N_11548);
or U12425 (N_12425,N_11601,N_11619);
or U12426 (N_12426,N_11875,N_11625);
nor U12427 (N_12427,N_11633,N_11580);
nor U12428 (N_12428,N_11911,N_11613);
or U12429 (N_12429,N_11549,N_11933);
nand U12430 (N_12430,N_11752,N_11693);
nor U12431 (N_12431,N_11970,N_11922);
nor U12432 (N_12432,N_11849,N_11658);
xor U12433 (N_12433,N_11754,N_11670);
or U12434 (N_12434,N_11521,N_11988);
xnor U12435 (N_12435,N_11977,N_11566);
nand U12436 (N_12436,N_11814,N_11957);
or U12437 (N_12437,N_11683,N_11870);
and U12438 (N_12438,N_11745,N_11584);
xnor U12439 (N_12439,N_11896,N_11663);
or U12440 (N_12440,N_11982,N_11814);
nor U12441 (N_12441,N_11840,N_11899);
nand U12442 (N_12442,N_11685,N_11534);
nand U12443 (N_12443,N_11500,N_11877);
and U12444 (N_12444,N_11767,N_11721);
or U12445 (N_12445,N_11584,N_11633);
nand U12446 (N_12446,N_11699,N_11598);
nand U12447 (N_12447,N_11814,N_11998);
nor U12448 (N_12448,N_11823,N_11748);
and U12449 (N_12449,N_11714,N_11693);
and U12450 (N_12450,N_11602,N_11628);
nor U12451 (N_12451,N_11783,N_11953);
xnor U12452 (N_12452,N_11997,N_11917);
nand U12453 (N_12453,N_11584,N_11892);
xnor U12454 (N_12454,N_11978,N_11593);
xnor U12455 (N_12455,N_11816,N_11619);
nor U12456 (N_12456,N_11811,N_11886);
nor U12457 (N_12457,N_11787,N_11724);
nor U12458 (N_12458,N_11897,N_11576);
and U12459 (N_12459,N_11935,N_11940);
nor U12460 (N_12460,N_11901,N_11991);
xor U12461 (N_12461,N_11871,N_11763);
nand U12462 (N_12462,N_11922,N_11967);
xnor U12463 (N_12463,N_11715,N_11890);
xor U12464 (N_12464,N_11746,N_11556);
nor U12465 (N_12465,N_11927,N_11581);
xor U12466 (N_12466,N_11795,N_11568);
xor U12467 (N_12467,N_11604,N_11648);
and U12468 (N_12468,N_11959,N_11999);
nor U12469 (N_12469,N_11819,N_11669);
and U12470 (N_12470,N_11991,N_11558);
nand U12471 (N_12471,N_11561,N_11713);
or U12472 (N_12472,N_11961,N_11822);
or U12473 (N_12473,N_11537,N_11824);
and U12474 (N_12474,N_11721,N_11580);
nor U12475 (N_12475,N_11959,N_11961);
nor U12476 (N_12476,N_11936,N_11804);
nand U12477 (N_12477,N_11920,N_11702);
xor U12478 (N_12478,N_11846,N_11939);
xnor U12479 (N_12479,N_11828,N_11637);
nand U12480 (N_12480,N_11563,N_11877);
or U12481 (N_12481,N_11792,N_11723);
xor U12482 (N_12482,N_11580,N_11714);
or U12483 (N_12483,N_11926,N_11824);
xnor U12484 (N_12484,N_11523,N_11569);
nand U12485 (N_12485,N_11724,N_11968);
nor U12486 (N_12486,N_11937,N_11777);
nand U12487 (N_12487,N_11830,N_11683);
or U12488 (N_12488,N_11515,N_11983);
nand U12489 (N_12489,N_11785,N_11535);
nand U12490 (N_12490,N_11884,N_11834);
xor U12491 (N_12491,N_11500,N_11678);
nor U12492 (N_12492,N_11905,N_11922);
and U12493 (N_12493,N_11971,N_11750);
and U12494 (N_12494,N_11801,N_11859);
nor U12495 (N_12495,N_11517,N_11876);
xor U12496 (N_12496,N_11522,N_11804);
nand U12497 (N_12497,N_11854,N_11978);
nand U12498 (N_12498,N_11588,N_11640);
or U12499 (N_12499,N_11883,N_11769);
xnor U12500 (N_12500,N_12195,N_12308);
xnor U12501 (N_12501,N_12234,N_12456);
or U12502 (N_12502,N_12087,N_12417);
nor U12503 (N_12503,N_12472,N_12215);
nor U12504 (N_12504,N_12477,N_12198);
nor U12505 (N_12505,N_12411,N_12406);
xor U12506 (N_12506,N_12491,N_12225);
or U12507 (N_12507,N_12250,N_12400);
xnor U12508 (N_12508,N_12105,N_12189);
and U12509 (N_12509,N_12233,N_12331);
or U12510 (N_12510,N_12364,N_12210);
or U12511 (N_12511,N_12144,N_12296);
nor U12512 (N_12512,N_12078,N_12330);
xor U12513 (N_12513,N_12414,N_12151);
xnor U12514 (N_12514,N_12407,N_12214);
or U12515 (N_12515,N_12249,N_12449);
or U12516 (N_12516,N_12377,N_12138);
and U12517 (N_12517,N_12060,N_12357);
xnor U12518 (N_12518,N_12262,N_12081);
xor U12519 (N_12519,N_12488,N_12036);
nor U12520 (N_12520,N_12143,N_12030);
or U12521 (N_12521,N_12485,N_12427);
nand U12522 (N_12522,N_12346,N_12358);
nand U12523 (N_12523,N_12177,N_12146);
nor U12524 (N_12524,N_12162,N_12051);
nand U12525 (N_12525,N_12307,N_12026);
and U12526 (N_12526,N_12267,N_12447);
and U12527 (N_12527,N_12245,N_12293);
and U12528 (N_12528,N_12123,N_12479);
and U12529 (N_12529,N_12113,N_12220);
or U12530 (N_12530,N_12286,N_12199);
xnor U12531 (N_12531,N_12154,N_12408);
or U12532 (N_12532,N_12440,N_12203);
and U12533 (N_12533,N_12202,N_12473);
and U12534 (N_12534,N_12284,N_12058);
and U12535 (N_12535,N_12270,N_12254);
and U12536 (N_12536,N_12363,N_12366);
xor U12537 (N_12537,N_12148,N_12335);
and U12538 (N_12538,N_12027,N_12108);
nor U12539 (N_12539,N_12495,N_12333);
or U12540 (N_12540,N_12006,N_12188);
nand U12541 (N_12541,N_12150,N_12106);
xnor U12542 (N_12542,N_12290,N_12423);
nand U12543 (N_12543,N_12176,N_12094);
xor U12544 (N_12544,N_12178,N_12183);
nor U12545 (N_12545,N_12111,N_12314);
and U12546 (N_12546,N_12185,N_12297);
nor U12547 (N_12547,N_12458,N_12071);
or U12548 (N_12548,N_12023,N_12080);
and U12549 (N_12549,N_12224,N_12247);
xor U12550 (N_12550,N_12464,N_12374);
nor U12551 (N_12551,N_12015,N_12244);
nand U12552 (N_12552,N_12315,N_12466);
nor U12553 (N_12553,N_12044,N_12226);
nor U12554 (N_12554,N_12276,N_12496);
or U12555 (N_12555,N_12391,N_12003);
and U12556 (N_12556,N_12371,N_12076);
nand U12557 (N_12557,N_12069,N_12103);
or U12558 (N_12558,N_12375,N_12347);
and U12559 (N_12559,N_12031,N_12370);
nor U12560 (N_12560,N_12342,N_12461);
nor U12561 (N_12561,N_12300,N_12119);
and U12562 (N_12562,N_12000,N_12088);
or U12563 (N_12563,N_12145,N_12127);
nand U12564 (N_12564,N_12237,N_12193);
or U12565 (N_12565,N_12478,N_12101);
or U12566 (N_12566,N_12043,N_12431);
and U12567 (N_12567,N_12022,N_12380);
or U12568 (N_12568,N_12499,N_12317);
and U12569 (N_12569,N_12355,N_12465);
nor U12570 (N_12570,N_12186,N_12446);
and U12571 (N_12571,N_12173,N_12344);
or U12572 (N_12572,N_12033,N_12450);
and U12573 (N_12573,N_12329,N_12426);
and U12574 (N_12574,N_12054,N_12309);
and U12575 (N_12575,N_12378,N_12131);
or U12576 (N_12576,N_12057,N_12028);
nand U12577 (N_12577,N_12050,N_12348);
and U12578 (N_12578,N_12480,N_12448);
nand U12579 (N_12579,N_12278,N_12048);
nor U12580 (N_12580,N_12045,N_12134);
nand U12581 (N_12581,N_12139,N_12126);
or U12582 (N_12582,N_12142,N_12194);
nor U12583 (N_12583,N_12065,N_12025);
nor U12584 (N_12584,N_12170,N_12291);
or U12585 (N_12585,N_12201,N_12271);
nand U12586 (N_12586,N_12320,N_12042);
nor U12587 (N_12587,N_12420,N_12181);
and U12588 (N_12588,N_12248,N_12133);
xnor U12589 (N_12589,N_12405,N_12090);
or U12590 (N_12590,N_12155,N_12086);
nor U12591 (N_12591,N_12191,N_12008);
nand U12592 (N_12592,N_12147,N_12040);
xnor U12593 (N_12593,N_12260,N_12324);
nor U12594 (N_12594,N_12056,N_12102);
xor U12595 (N_12595,N_12373,N_12356);
xor U12596 (N_12596,N_12457,N_12012);
nor U12597 (N_12597,N_12402,N_12152);
nand U12598 (N_12598,N_12116,N_12157);
or U12599 (N_12599,N_12269,N_12428);
or U12600 (N_12600,N_12137,N_12359);
and U12601 (N_12601,N_12082,N_12014);
xor U12602 (N_12602,N_12483,N_12268);
nand U12603 (N_12603,N_12239,N_12149);
xnor U12604 (N_12604,N_12338,N_12024);
and U12605 (N_12605,N_12002,N_12068);
or U12606 (N_12606,N_12436,N_12107);
nor U12607 (N_12607,N_12172,N_12334);
nand U12608 (N_12608,N_12416,N_12301);
nor U12609 (N_12609,N_12403,N_12174);
nand U12610 (N_12610,N_12386,N_12265);
xnor U12611 (N_12611,N_12390,N_12441);
xor U12612 (N_12612,N_12322,N_12093);
nor U12613 (N_12613,N_12122,N_12232);
or U12614 (N_12614,N_12099,N_12445);
nand U12615 (N_12615,N_12396,N_12295);
and U12616 (N_12616,N_12264,N_12392);
and U12617 (N_12617,N_12498,N_12156);
nor U12618 (N_12618,N_12326,N_12494);
nor U12619 (N_12619,N_12135,N_12029);
nor U12620 (N_12620,N_12312,N_12055);
xnor U12621 (N_12621,N_12001,N_12217);
nand U12622 (N_12622,N_12236,N_12437);
nor U12623 (N_12623,N_12316,N_12251);
xnor U12624 (N_12624,N_12339,N_12223);
xor U12625 (N_12625,N_12351,N_12281);
or U12626 (N_12626,N_12257,N_12327);
or U12627 (N_12627,N_12365,N_12298);
nor U12628 (N_12628,N_12319,N_12109);
nand U12629 (N_12629,N_12362,N_12490);
nand U12630 (N_12630,N_12360,N_12323);
nor U12631 (N_12631,N_12263,N_12182);
and U12632 (N_12632,N_12282,N_12100);
nand U12633 (N_12633,N_12397,N_12171);
nand U12634 (N_12634,N_12034,N_12321);
or U12635 (N_12635,N_12429,N_12104);
nor U12636 (N_12636,N_12067,N_12388);
xnor U12637 (N_12637,N_12372,N_12433);
and U12638 (N_12638,N_12279,N_12114);
xor U12639 (N_12639,N_12368,N_12482);
or U12640 (N_12640,N_12453,N_12179);
xor U12641 (N_12641,N_12240,N_12350);
nor U12642 (N_12642,N_12163,N_12016);
xor U12643 (N_12643,N_12164,N_12394);
nand U12644 (N_12644,N_12175,N_12092);
nand U12645 (N_12645,N_12196,N_12169);
nor U12646 (N_12646,N_12439,N_12084);
xnor U12647 (N_12647,N_12454,N_12294);
xnor U12648 (N_12648,N_12011,N_12241);
nand U12649 (N_12649,N_12010,N_12197);
and U12650 (N_12650,N_12097,N_12325);
or U12651 (N_12651,N_12077,N_12066);
nor U12652 (N_12652,N_12393,N_12277);
or U12653 (N_12653,N_12207,N_12021);
or U12654 (N_12654,N_12306,N_12367);
xnor U12655 (N_12655,N_12128,N_12412);
nand U12656 (N_12656,N_12005,N_12253);
or U12657 (N_12657,N_12049,N_12337);
nand U12658 (N_12658,N_12047,N_12349);
nand U12659 (N_12659,N_12098,N_12418);
nand U12660 (N_12660,N_12444,N_12039);
or U12661 (N_12661,N_12211,N_12118);
xnor U12662 (N_12662,N_12395,N_12242);
nor U12663 (N_12663,N_12352,N_12041);
xor U12664 (N_12664,N_12474,N_12061);
xnor U12665 (N_12665,N_12341,N_12310);
nor U12666 (N_12666,N_12385,N_12227);
and U12667 (N_12667,N_12129,N_12208);
or U12668 (N_12668,N_12354,N_12432);
or U12669 (N_12669,N_12259,N_12046);
nor U12670 (N_12670,N_12460,N_12059);
and U12671 (N_12671,N_12074,N_12415);
nand U12672 (N_12672,N_12140,N_12110);
and U12673 (N_12673,N_12289,N_12180);
nor U12674 (N_12674,N_12261,N_12213);
and U12675 (N_12675,N_12379,N_12165);
xnor U12676 (N_12676,N_12421,N_12062);
nor U12677 (N_12677,N_12381,N_12486);
xor U12678 (N_12678,N_12459,N_12332);
xnor U12679 (N_12679,N_12443,N_12343);
nand U12680 (N_12680,N_12302,N_12303);
xor U12681 (N_12681,N_12455,N_12299);
nor U12682 (N_12682,N_12075,N_12422);
or U12683 (N_12683,N_12019,N_12409);
nand U12684 (N_12684,N_12125,N_12166);
nand U12685 (N_12685,N_12216,N_12463);
xor U12686 (N_12686,N_12384,N_12221);
nor U12687 (N_12687,N_12252,N_12401);
nor U12688 (N_12688,N_12283,N_12340);
nor U12689 (N_12689,N_12492,N_12287);
and U12690 (N_12690,N_12089,N_12229);
nand U12691 (N_12691,N_12212,N_12266);
nor U12692 (N_12692,N_12072,N_12153);
and U12693 (N_12693,N_12246,N_12305);
or U12694 (N_12694,N_12487,N_12288);
nand U12695 (N_12695,N_12243,N_12132);
or U12696 (N_12696,N_12083,N_12079);
nand U12697 (N_12697,N_12425,N_12064);
nor U12698 (N_12698,N_12256,N_12235);
or U12699 (N_12699,N_12070,N_12184);
or U12700 (N_12700,N_12004,N_12318);
xor U12701 (N_12701,N_12468,N_12493);
nand U12702 (N_12702,N_12419,N_12020);
nor U12703 (N_12703,N_12389,N_12387);
nand U12704 (N_12704,N_12311,N_12255);
nor U12705 (N_12705,N_12369,N_12467);
or U12706 (N_12706,N_12209,N_12274);
xor U12707 (N_12707,N_12238,N_12353);
and U12708 (N_12708,N_12190,N_12345);
xor U12709 (N_12709,N_12438,N_12413);
nor U12710 (N_12710,N_12091,N_12073);
nor U12711 (N_12711,N_12410,N_12398);
and U12712 (N_12712,N_12037,N_12361);
xnor U12713 (N_12713,N_12452,N_12471);
and U12714 (N_12714,N_12130,N_12095);
and U12715 (N_12715,N_12497,N_12328);
xnor U12716 (N_12716,N_12218,N_12204);
and U12717 (N_12717,N_12292,N_12435);
nand U12718 (N_12718,N_12117,N_12304);
or U12719 (N_12719,N_12469,N_12200);
nand U12720 (N_12720,N_12481,N_12115);
nand U12721 (N_12721,N_12285,N_12205);
and U12722 (N_12722,N_12404,N_12007);
or U12723 (N_12723,N_12032,N_12160);
nor U12724 (N_12724,N_12124,N_12484);
xnor U12725 (N_12725,N_12038,N_12489);
nor U12726 (N_12726,N_12275,N_12336);
or U12727 (N_12727,N_12442,N_12168);
nand U12728 (N_12728,N_12112,N_12085);
nand U12729 (N_12729,N_12136,N_12273);
and U12730 (N_12730,N_12192,N_12376);
xor U12731 (N_12731,N_12159,N_12158);
nor U12732 (N_12732,N_12230,N_12399);
nand U12733 (N_12733,N_12017,N_12475);
and U12734 (N_12734,N_12272,N_12161);
xor U12735 (N_12735,N_12383,N_12141);
nand U12736 (N_12736,N_12009,N_12219);
and U12737 (N_12737,N_12052,N_12222);
xor U12738 (N_12738,N_12053,N_12063);
xor U12739 (N_12739,N_12382,N_12228);
nor U12740 (N_12740,N_12035,N_12187);
nor U12741 (N_12741,N_12462,N_12434);
xnor U12742 (N_12742,N_12018,N_12096);
xor U12743 (N_12743,N_12424,N_12430);
nor U12744 (N_12744,N_12470,N_12280);
nand U12745 (N_12745,N_12476,N_12120);
nor U12746 (N_12746,N_12258,N_12231);
nand U12747 (N_12747,N_12313,N_12167);
and U12748 (N_12748,N_12451,N_12206);
nor U12749 (N_12749,N_12013,N_12121);
or U12750 (N_12750,N_12056,N_12270);
nor U12751 (N_12751,N_12029,N_12136);
nand U12752 (N_12752,N_12352,N_12233);
nand U12753 (N_12753,N_12122,N_12144);
nor U12754 (N_12754,N_12364,N_12201);
or U12755 (N_12755,N_12255,N_12309);
nand U12756 (N_12756,N_12073,N_12397);
xor U12757 (N_12757,N_12381,N_12390);
xnor U12758 (N_12758,N_12190,N_12330);
xnor U12759 (N_12759,N_12463,N_12243);
nand U12760 (N_12760,N_12231,N_12031);
or U12761 (N_12761,N_12044,N_12431);
xnor U12762 (N_12762,N_12160,N_12235);
nor U12763 (N_12763,N_12300,N_12387);
xnor U12764 (N_12764,N_12462,N_12124);
nand U12765 (N_12765,N_12118,N_12116);
nand U12766 (N_12766,N_12337,N_12063);
xnor U12767 (N_12767,N_12458,N_12485);
nor U12768 (N_12768,N_12311,N_12268);
xor U12769 (N_12769,N_12387,N_12125);
xor U12770 (N_12770,N_12248,N_12138);
or U12771 (N_12771,N_12252,N_12419);
or U12772 (N_12772,N_12271,N_12224);
nor U12773 (N_12773,N_12139,N_12027);
and U12774 (N_12774,N_12374,N_12080);
xor U12775 (N_12775,N_12032,N_12107);
nand U12776 (N_12776,N_12176,N_12345);
or U12777 (N_12777,N_12255,N_12385);
or U12778 (N_12778,N_12344,N_12258);
or U12779 (N_12779,N_12026,N_12266);
nand U12780 (N_12780,N_12021,N_12087);
or U12781 (N_12781,N_12451,N_12473);
nor U12782 (N_12782,N_12440,N_12358);
or U12783 (N_12783,N_12481,N_12124);
nand U12784 (N_12784,N_12267,N_12420);
and U12785 (N_12785,N_12059,N_12374);
nor U12786 (N_12786,N_12165,N_12281);
nand U12787 (N_12787,N_12079,N_12332);
nor U12788 (N_12788,N_12474,N_12448);
nand U12789 (N_12789,N_12210,N_12209);
xnor U12790 (N_12790,N_12049,N_12113);
or U12791 (N_12791,N_12337,N_12244);
and U12792 (N_12792,N_12093,N_12461);
nor U12793 (N_12793,N_12273,N_12375);
nor U12794 (N_12794,N_12078,N_12112);
and U12795 (N_12795,N_12239,N_12338);
and U12796 (N_12796,N_12356,N_12233);
or U12797 (N_12797,N_12218,N_12086);
and U12798 (N_12798,N_12145,N_12263);
nand U12799 (N_12799,N_12141,N_12283);
xnor U12800 (N_12800,N_12487,N_12321);
and U12801 (N_12801,N_12170,N_12000);
nor U12802 (N_12802,N_12096,N_12424);
xnor U12803 (N_12803,N_12472,N_12204);
or U12804 (N_12804,N_12118,N_12020);
nand U12805 (N_12805,N_12066,N_12456);
or U12806 (N_12806,N_12487,N_12380);
or U12807 (N_12807,N_12000,N_12215);
nand U12808 (N_12808,N_12442,N_12286);
xor U12809 (N_12809,N_12059,N_12270);
nor U12810 (N_12810,N_12296,N_12333);
xor U12811 (N_12811,N_12042,N_12039);
nor U12812 (N_12812,N_12014,N_12017);
and U12813 (N_12813,N_12061,N_12459);
and U12814 (N_12814,N_12468,N_12435);
nand U12815 (N_12815,N_12408,N_12351);
nor U12816 (N_12816,N_12458,N_12187);
and U12817 (N_12817,N_12427,N_12439);
xnor U12818 (N_12818,N_12230,N_12118);
nand U12819 (N_12819,N_12003,N_12355);
xnor U12820 (N_12820,N_12268,N_12394);
or U12821 (N_12821,N_12132,N_12246);
nor U12822 (N_12822,N_12290,N_12277);
xor U12823 (N_12823,N_12411,N_12414);
xor U12824 (N_12824,N_12402,N_12251);
or U12825 (N_12825,N_12465,N_12157);
nand U12826 (N_12826,N_12465,N_12090);
nor U12827 (N_12827,N_12373,N_12361);
and U12828 (N_12828,N_12296,N_12466);
xnor U12829 (N_12829,N_12130,N_12194);
xor U12830 (N_12830,N_12385,N_12055);
nor U12831 (N_12831,N_12101,N_12296);
xor U12832 (N_12832,N_12037,N_12283);
and U12833 (N_12833,N_12116,N_12186);
nor U12834 (N_12834,N_12099,N_12214);
nor U12835 (N_12835,N_12044,N_12191);
nand U12836 (N_12836,N_12403,N_12078);
and U12837 (N_12837,N_12150,N_12146);
or U12838 (N_12838,N_12092,N_12286);
nand U12839 (N_12839,N_12343,N_12229);
xnor U12840 (N_12840,N_12313,N_12066);
and U12841 (N_12841,N_12491,N_12423);
and U12842 (N_12842,N_12435,N_12463);
and U12843 (N_12843,N_12158,N_12213);
and U12844 (N_12844,N_12285,N_12094);
nor U12845 (N_12845,N_12025,N_12469);
nand U12846 (N_12846,N_12109,N_12217);
or U12847 (N_12847,N_12076,N_12405);
xor U12848 (N_12848,N_12278,N_12423);
and U12849 (N_12849,N_12482,N_12075);
nand U12850 (N_12850,N_12119,N_12283);
nor U12851 (N_12851,N_12416,N_12220);
nor U12852 (N_12852,N_12191,N_12268);
nand U12853 (N_12853,N_12156,N_12225);
nor U12854 (N_12854,N_12307,N_12148);
and U12855 (N_12855,N_12096,N_12420);
or U12856 (N_12856,N_12299,N_12104);
xor U12857 (N_12857,N_12423,N_12064);
nand U12858 (N_12858,N_12028,N_12068);
or U12859 (N_12859,N_12114,N_12167);
nand U12860 (N_12860,N_12027,N_12372);
and U12861 (N_12861,N_12135,N_12305);
or U12862 (N_12862,N_12036,N_12254);
xnor U12863 (N_12863,N_12479,N_12006);
or U12864 (N_12864,N_12001,N_12119);
xor U12865 (N_12865,N_12447,N_12404);
or U12866 (N_12866,N_12490,N_12443);
or U12867 (N_12867,N_12214,N_12421);
xor U12868 (N_12868,N_12021,N_12093);
and U12869 (N_12869,N_12368,N_12146);
nand U12870 (N_12870,N_12393,N_12420);
or U12871 (N_12871,N_12346,N_12231);
nor U12872 (N_12872,N_12406,N_12028);
nand U12873 (N_12873,N_12300,N_12176);
xnor U12874 (N_12874,N_12486,N_12306);
or U12875 (N_12875,N_12169,N_12372);
and U12876 (N_12876,N_12083,N_12353);
or U12877 (N_12877,N_12258,N_12105);
nand U12878 (N_12878,N_12178,N_12214);
nand U12879 (N_12879,N_12422,N_12111);
nor U12880 (N_12880,N_12172,N_12054);
nand U12881 (N_12881,N_12187,N_12331);
xnor U12882 (N_12882,N_12215,N_12470);
nor U12883 (N_12883,N_12046,N_12036);
nand U12884 (N_12884,N_12355,N_12125);
nand U12885 (N_12885,N_12228,N_12197);
nand U12886 (N_12886,N_12136,N_12256);
nor U12887 (N_12887,N_12066,N_12397);
nand U12888 (N_12888,N_12219,N_12097);
nor U12889 (N_12889,N_12145,N_12105);
and U12890 (N_12890,N_12033,N_12185);
xnor U12891 (N_12891,N_12315,N_12018);
and U12892 (N_12892,N_12478,N_12334);
or U12893 (N_12893,N_12058,N_12365);
xnor U12894 (N_12894,N_12142,N_12352);
or U12895 (N_12895,N_12353,N_12478);
xnor U12896 (N_12896,N_12220,N_12204);
nand U12897 (N_12897,N_12263,N_12344);
nand U12898 (N_12898,N_12366,N_12192);
nand U12899 (N_12899,N_12348,N_12415);
and U12900 (N_12900,N_12128,N_12391);
xnor U12901 (N_12901,N_12168,N_12454);
nand U12902 (N_12902,N_12009,N_12105);
nand U12903 (N_12903,N_12101,N_12147);
or U12904 (N_12904,N_12348,N_12059);
and U12905 (N_12905,N_12413,N_12206);
xnor U12906 (N_12906,N_12098,N_12172);
or U12907 (N_12907,N_12117,N_12003);
nand U12908 (N_12908,N_12108,N_12123);
or U12909 (N_12909,N_12011,N_12402);
nand U12910 (N_12910,N_12076,N_12236);
and U12911 (N_12911,N_12119,N_12142);
xnor U12912 (N_12912,N_12406,N_12031);
xnor U12913 (N_12913,N_12226,N_12452);
xor U12914 (N_12914,N_12079,N_12419);
nand U12915 (N_12915,N_12480,N_12396);
nor U12916 (N_12916,N_12240,N_12241);
xnor U12917 (N_12917,N_12454,N_12332);
nor U12918 (N_12918,N_12477,N_12003);
or U12919 (N_12919,N_12237,N_12119);
nor U12920 (N_12920,N_12204,N_12482);
and U12921 (N_12921,N_12454,N_12408);
xor U12922 (N_12922,N_12106,N_12039);
nor U12923 (N_12923,N_12381,N_12259);
nor U12924 (N_12924,N_12245,N_12341);
nand U12925 (N_12925,N_12408,N_12303);
nand U12926 (N_12926,N_12405,N_12030);
xnor U12927 (N_12927,N_12185,N_12199);
nor U12928 (N_12928,N_12165,N_12468);
nor U12929 (N_12929,N_12069,N_12238);
xnor U12930 (N_12930,N_12155,N_12232);
xnor U12931 (N_12931,N_12141,N_12451);
nor U12932 (N_12932,N_12262,N_12379);
or U12933 (N_12933,N_12239,N_12075);
nor U12934 (N_12934,N_12362,N_12059);
and U12935 (N_12935,N_12484,N_12092);
and U12936 (N_12936,N_12070,N_12320);
nand U12937 (N_12937,N_12111,N_12151);
nor U12938 (N_12938,N_12146,N_12431);
nand U12939 (N_12939,N_12289,N_12388);
or U12940 (N_12940,N_12184,N_12055);
xnor U12941 (N_12941,N_12432,N_12171);
xnor U12942 (N_12942,N_12250,N_12130);
and U12943 (N_12943,N_12306,N_12439);
nand U12944 (N_12944,N_12217,N_12063);
nand U12945 (N_12945,N_12021,N_12480);
or U12946 (N_12946,N_12380,N_12179);
or U12947 (N_12947,N_12217,N_12266);
xor U12948 (N_12948,N_12244,N_12418);
xnor U12949 (N_12949,N_12037,N_12387);
or U12950 (N_12950,N_12459,N_12194);
or U12951 (N_12951,N_12344,N_12332);
and U12952 (N_12952,N_12073,N_12076);
or U12953 (N_12953,N_12132,N_12076);
or U12954 (N_12954,N_12106,N_12171);
xor U12955 (N_12955,N_12448,N_12187);
nor U12956 (N_12956,N_12090,N_12378);
or U12957 (N_12957,N_12241,N_12149);
and U12958 (N_12958,N_12131,N_12215);
xnor U12959 (N_12959,N_12002,N_12079);
and U12960 (N_12960,N_12385,N_12365);
nand U12961 (N_12961,N_12275,N_12312);
nor U12962 (N_12962,N_12026,N_12351);
nand U12963 (N_12963,N_12114,N_12283);
xor U12964 (N_12964,N_12472,N_12340);
or U12965 (N_12965,N_12387,N_12483);
xnor U12966 (N_12966,N_12222,N_12340);
xnor U12967 (N_12967,N_12360,N_12381);
nand U12968 (N_12968,N_12404,N_12168);
nand U12969 (N_12969,N_12260,N_12210);
and U12970 (N_12970,N_12347,N_12212);
nand U12971 (N_12971,N_12092,N_12202);
xnor U12972 (N_12972,N_12295,N_12453);
nor U12973 (N_12973,N_12452,N_12173);
nand U12974 (N_12974,N_12149,N_12046);
nor U12975 (N_12975,N_12010,N_12432);
nor U12976 (N_12976,N_12227,N_12105);
nor U12977 (N_12977,N_12095,N_12126);
nor U12978 (N_12978,N_12473,N_12416);
xor U12979 (N_12979,N_12388,N_12284);
nand U12980 (N_12980,N_12397,N_12365);
nor U12981 (N_12981,N_12077,N_12279);
nand U12982 (N_12982,N_12066,N_12315);
nor U12983 (N_12983,N_12426,N_12105);
and U12984 (N_12984,N_12219,N_12405);
nor U12985 (N_12985,N_12002,N_12034);
and U12986 (N_12986,N_12467,N_12250);
nor U12987 (N_12987,N_12368,N_12453);
nand U12988 (N_12988,N_12303,N_12249);
nand U12989 (N_12989,N_12495,N_12188);
and U12990 (N_12990,N_12152,N_12495);
nand U12991 (N_12991,N_12432,N_12378);
xor U12992 (N_12992,N_12172,N_12217);
xnor U12993 (N_12993,N_12032,N_12339);
or U12994 (N_12994,N_12157,N_12019);
or U12995 (N_12995,N_12270,N_12214);
xnor U12996 (N_12996,N_12315,N_12352);
and U12997 (N_12997,N_12172,N_12496);
and U12998 (N_12998,N_12319,N_12425);
or U12999 (N_12999,N_12391,N_12353);
nand U13000 (N_13000,N_12981,N_12532);
nand U13001 (N_13001,N_12903,N_12553);
nor U13002 (N_13002,N_12504,N_12699);
xor U13003 (N_13003,N_12618,N_12865);
nor U13004 (N_13004,N_12871,N_12772);
xnor U13005 (N_13005,N_12637,N_12831);
or U13006 (N_13006,N_12956,N_12842);
nor U13007 (N_13007,N_12507,N_12920);
nor U13008 (N_13008,N_12967,N_12513);
xnor U13009 (N_13009,N_12774,N_12694);
or U13010 (N_13010,N_12990,N_12812);
and U13011 (N_13011,N_12782,N_12900);
xor U13012 (N_13012,N_12551,N_12785);
nand U13013 (N_13013,N_12888,N_12586);
nand U13014 (N_13014,N_12718,N_12789);
nor U13015 (N_13015,N_12826,N_12672);
or U13016 (N_13016,N_12550,N_12657);
nand U13017 (N_13017,N_12554,N_12670);
and U13018 (N_13018,N_12603,N_12620);
or U13019 (N_13019,N_12750,N_12829);
or U13020 (N_13020,N_12910,N_12567);
and U13021 (N_13021,N_12897,N_12992);
or U13022 (N_13022,N_12945,N_12678);
xor U13023 (N_13023,N_12837,N_12748);
and U13024 (N_13024,N_12839,N_12998);
or U13025 (N_13025,N_12723,N_12921);
nor U13026 (N_13026,N_12914,N_12960);
xnor U13027 (N_13027,N_12760,N_12957);
nor U13028 (N_13028,N_12629,N_12882);
or U13029 (N_13029,N_12576,N_12597);
and U13030 (N_13030,N_12798,N_12705);
xor U13031 (N_13031,N_12820,N_12793);
nor U13032 (N_13032,N_12850,N_12607);
and U13033 (N_13033,N_12704,N_12674);
nor U13034 (N_13034,N_12982,N_12630);
xor U13035 (N_13035,N_12893,N_12941);
or U13036 (N_13036,N_12765,N_12936);
xor U13037 (N_13037,N_12885,N_12622);
and U13038 (N_13038,N_12777,N_12632);
nand U13039 (N_13039,N_12980,N_12677);
nor U13040 (N_13040,N_12841,N_12985);
nor U13041 (N_13041,N_12883,N_12728);
nor U13042 (N_13042,N_12948,N_12844);
xnor U13043 (N_13043,N_12743,N_12825);
and U13044 (N_13044,N_12868,N_12827);
xnor U13045 (N_13045,N_12911,N_12977);
and U13046 (N_13046,N_12619,N_12764);
and U13047 (N_13047,N_12819,N_12509);
or U13048 (N_13048,N_12573,N_12621);
and U13049 (N_13049,N_12665,N_12526);
xnor U13050 (N_13050,N_12984,N_12878);
or U13051 (N_13051,N_12915,N_12738);
nand U13052 (N_13052,N_12582,N_12849);
or U13053 (N_13053,N_12611,N_12780);
and U13054 (N_13054,N_12500,N_12845);
nand U13055 (N_13055,N_12909,N_12881);
nor U13056 (N_13056,N_12527,N_12668);
and U13057 (N_13057,N_12733,N_12864);
and U13058 (N_13058,N_12763,N_12684);
and U13059 (N_13059,N_12523,N_12828);
and U13060 (N_13060,N_12719,N_12861);
xnor U13061 (N_13061,N_12902,N_12688);
xnor U13062 (N_13062,N_12856,N_12848);
nand U13063 (N_13063,N_12735,N_12536);
nor U13064 (N_13064,N_12519,N_12824);
xnor U13065 (N_13065,N_12886,N_12924);
and U13066 (N_13066,N_12997,N_12737);
or U13067 (N_13067,N_12862,N_12912);
xor U13068 (N_13068,N_12725,N_12769);
or U13069 (N_13069,N_12524,N_12716);
and U13070 (N_13070,N_12867,N_12757);
and U13071 (N_13071,N_12649,N_12510);
and U13072 (N_13072,N_12580,N_12836);
xor U13073 (N_13073,N_12802,N_12773);
or U13074 (N_13074,N_12592,N_12788);
nor U13075 (N_13075,N_12559,N_12961);
xor U13076 (N_13076,N_12821,N_12575);
or U13077 (N_13077,N_12690,N_12934);
or U13078 (N_13078,N_12648,N_12685);
and U13079 (N_13079,N_12853,N_12574);
xor U13080 (N_13080,N_12954,N_12969);
nand U13081 (N_13081,N_12606,N_12561);
nand U13082 (N_13082,N_12917,N_12535);
and U13083 (N_13083,N_12778,N_12986);
xnor U13084 (N_13084,N_12754,N_12762);
nand U13085 (N_13085,N_12680,N_12963);
nand U13086 (N_13086,N_12692,N_12758);
and U13087 (N_13087,N_12614,N_12811);
nand U13088 (N_13088,N_12974,N_12999);
nor U13089 (N_13089,N_12726,N_12759);
nand U13090 (N_13090,N_12833,N_12993);
nor U13091 (N_13091,N_12698,N_12816);
nor U13092 (N_13092,N_12939,N_12894);
or U13093 (N_13093,N_12506,N_12892);
nor U13094 (N_13094,N_12585,N_12695);
and U13095 (N_13095,N_12708,N_12971);
nor U13096 (N_13096,N_12741,N_12783);
nand U13097 (N_13097,N_12988,N_12615);
xnor U13098 (N_13098,N_12562,N_12807);
nand U13099 (N_13099,N_12919,N_12715);
and U13100 (N_13100,N_12563,N_12639);
xor U13101 (N_13101,N_12751,N_12656);
or U13102 (N_13102,N_12702,N_12959);
nor U13103 (N_13103,N_12840,N_12756);
xnor U13104 (N_13104,N_12505,N_12681);
or U13105 (N_13105,N_12556,N_12873);
or U13106 (N_13106,N_12687,N_12608);
nand U13107 (N_13107,N_12935,N_12682);
or U13108 (N_13108,N_12642,N_12929);
or U13109 (N_13109,N_12635,N_12846);
nor U13110 (N_13110,N_12636,N_12647);
or U13111 (N_13111,N_12875,N_12626);
xnor U13112 (N_13112,N_12791,N_12858);
and U13113 (N_13113,N_12666,N_12801);
or U13114 (N_13114,N_12720,N_12518);
and U13115 (N_13115,N_12852,N_12706);
xnor U13116 (N_13116,N_12926,N_12591);
or U13117 (N_13117,N_12517,N_12970);
nand U13118 (N_13118,N_12928,N_12638);
nand U13119 (N_13119,N_12860,N_12631);
nor U13120 (N_13120,N_12516,N_12533);
nor U13121 (N_13121,N_12528,N_12958);
and U13122 (N_13122,N_12525,N_12923);
and U13123 (N_13123,N_12755,N_12729);
or U13124 (N_13124,N_12799,N_12584);
or U13125 (N_13125,N_12673,N_12805);
xnor U13126 (N_13126,N_12529,N_12855);
nor U13127 (N_13127,N_12601,N_12627);
nor U13128 (N_13128,N_12596,N_12796);
or U13129 (N_13129,N_12545,N_12641);
and U13130 (N_13130,N_12835,N_12895);
xor U13131 (N_13131,N_12818,N_12650);
or U13132 (N_13132,N_12968,N_12918);
or U13133 (N_13133,N_12595,N_12538);
nand U13134 (N_13134,N_12579,N_12691);
nand U13135 (N_13135,N_12625,N_12710);
nand U13136 (N_13136,N_12887,N_12823);
and U13137 (N_13137,N_12697,N_12880);
and U13138 (N_13138,N_12612,N_12983);
xor U13139 (N_13139,N_12966,N_12730);
xnor U13140 (N_13140,N_12976,N_12962);
xor U13141 (N_13141,N_12570,N_12989);
and U13142 (N_13142,N_12790,N_12740);
and U13143 (N_13143,N_12520,N_12943);
xor U13144 (N_13144,N_12834,N_12944);
nand U13145 (N_13145,N_12515,N_12600);
and U13146 (N_13146,N_12775,N_12731);
nand U13147 (N_13147,N_12664,N_12714);
and U13148 (N_13148,N_12501,N_12599);
or U13149 (N_13149,N_12671,N_12727);
and U13150 (N_13150,N_12663,N_12899);
and U13151 (N_13151,N_12544,N_12761);
or U13152 (N_13152,N_12593,N_12679);
xor U13153 (N_13153,N_12991,N_12587);
xor U13154 (N_13154,N_12891,N_12749);
and U13155 (N_13155,N_12616,N_12797);
nor U13156 (N_13156,N_12511,N_12675);
nor U13157 (N_13157,N_12667,N_12514);
nand U13158 (N_13158,N_12925,N_12572);
nor U13159 (N_13159,N_12508,N_12734);
nor U13160 (N_13160,N_12598,N_12901);
nand U13161 (N_13161,N_12537,N_12541);
xor U13162 (N_13162,N_12589,N_12847);
or U13163 (N_13163,N_12571,N_12542);
nor U13164 (N_13164,N_12813,N_12905);
xor U13165 (N_13165,N_12930,N_12549);
or U13166 (N_13166,N_12686,N_12744);
and U13167 (N_13167,N_12776,N_12870);
nand U13168 (N_13168,N_12569,N_12683);
nand U13169 (N_13169,N_12978,N_12916);
or U13170 (N_13170,N_12908,N_12784);
nand U13171 (N_13171,N_12721,N_12953);
nand U13172 (N_13172,N_12605,N_12712);
or U13173 (N_13173,N_12724,N_12651);
or U13174 (N_13174,N_12800,N_12947);
xor U13175 (N_13175,N_12717,N_12661);
or U13176 (N_13176,N_12964,N_12932);
xnor U13177 (N_13177,N_12907,N_12940);
nand U13178 (N_13178,N_12808,N_12530);
nand U13179 (N_13179,N_12972,N_12604);
nor U13180 (N_13180,N_12779,N_12951);
nand U13181 (N_13181,N_12560,N_12857);
xor U13182 (N_13182,N_12781,N_12889);
or U13183 (N_13183,N_12872,N_12624);
and U13184 (N_13184,N_12874,N_12931);
nand U13185 (N_13185,N_12747,N_12746);
xnor U13186 (N_13186,N_12927,N_12568);
nand U13187 (N_13187,N_12806,N_12906);
nor U13188 (N_13188,N_12884,N_12896);
nor U13189 (N_13189,N_12736,N_12644);
and U13190 (N_13190,N_12803,N_12768);
or U13191 (N_13191,N_12946,N_12659);
nor U13192 (N_13192,N_12742,N_12832);
nor U13193 (N_13193,N_12555,N_12890);
or U13194 (N_13194,N_12794,N_12658);
nand U13195 (N_13195,N_12922,N_12534);
nor U13196 (N_13196,N_12830,N_12531);
nor U13197 (N_13197,N_12843,N_12558);
or U13198 (N_13198,N_12937,N_12609);
nand U13199 (N_13199,N_12552,N_12942);
or U13200 (N_13200,N_12546,N_12689);
or U13201 (N_13201,N_12594,N_12696);
or U13202 (N_13202,N_12711,N_12652);
and U13203 (N_13203,N_12628,N_12640);
xor U13204 (N_13204,N_12952,N_12822);
xnor U13205 (N_13205,N_12617,N_12660);
xor U13206 (N_13206,N_12804,N_12613);
nand U13207 (N_13207,N_12950,N_12877);
or U13208 (N_13208,N_12786,N_12577);
nor U13209 (N_13209,N_12522,N_12540);
or U13210 (N_13210,N_12787,N_12566);
nor U13211 (N_13211,N_12987,N_12578);
nor U13212 (N_13212,N_12913,N_12869);
nand U13213 (N_13213,N_12753,N_12610);
nand U13214 (N_13214,N_12645,N_12866);
and U13215 (N_13215,N_12732,N_12810);
and U13216 (N_13216,N_12633,N_12838);
nand U13217 (N_13217,N_12996,N_12770);
nor U13218 (N_13218,N_12979,N_12709);
nor U13219 (N_13219,N_12851,N_12512);
nand U13220 (N_13220,N_12557,N_12933);
xor U13221 (N_13221,N_12854,N_12564);
or U13222 (N_13222,N_12703,N_12814);
xnor U13223 (N_13223,N_12634,N_12539);
xnor U13224 (N_13224,N_12548,N_12655);
and U13225 (N_13225,N_12713,N_12521);
xnor U13226 (N_13226,N_12503,N_12973);
xor U13227 (N_13227,N_12662,N_12771);
nor U13228 (N_13228,N_12879,N_12792);
nand U13229 (N_13229,N_12739,N_12547);
nor U13230 (N_13230,N_12669,N_12817);
nor U13231 (N_13231,N_12722,N_12646);
nand U13232 (N_13232,N_12904,N_12745);
nand U13233 (N_13233,N_12949,N_12653);
nor U13234 (N_13234,N_12654,N_12767);
xor U13235 (N_13235,N_12995,N_12752);
nor U13236 (N_13236,N_12898,N_12766);
nand U13237 (N_13237,N_12965,N_12955);
and U13238 (N_13238,N_12590,N_12602);
nor U13239 (N_13239,N_12859,N_12809);
or U13240 (N_13240,N_12583,N_12938);
or U13241 (N_13241,N_12700,N_12994);
and U13242 (N_13242,N_12795,N_12588);
xnor U13243 (N_13243,N_12623,N_12643);
and U13244 (N_13244,N_12701,N_12565);
and U13245 (N_13245,N_12975,N_12815);
and U13246 (N_13246,N_12581,N_12693);
or U13247 (N_13247,N_12707,N_12876);
nand U13248 (N_13248,N_12863,N_12676);
nand U13249 (N_13249,N_12543,N_12502);
nor U13250 (N_13250,N_12974,N_12532);
or U13251 (N_13251,N_12646,N_12503);
xor U13252 (N_13252,N_12596,N_12523);
xor U13253 (N_13253,N_12981,N_12839);
nor U13254 (N_13254,N_12830,N_12666);
or U13255 (N_13255,N_12886,N_12687);
xnor U13256 (N_13256,N_12560,N_12730);
xor U13257 (N_13257,N_12870,N_12533);
or U13258 (N_13258,N_12905,N_12715);
or U13259 (N_13259,N_12841,N_12992);
and U13260 (N_13260,N_12735,N_12608);
nor U13261 (N_13261,N_12600,N_12854);
xor U13262 (N_13262,N_12815,N_12760);
nand U13263 (N_13263,N_12777,N_12928);
and U13264 (N_13264,N_12647,N_12524);
xor U13265 (N_13265,N_12527,N_12872);
xnor U13266 (N_13266,N_12646,N_12710);
nand U13267 (N_13267,N_12527,N_12512);
nor U13268 (N_13268,N_12566,N_12622);
nand U13269 (N_13269,N_12647,N_12709);
nor U13270 (N_13270,N_12576,N_12773);
or U13271 (N_13271,N_12936,N_12945);
or U13272 (N_13272,N_12536,N_12633);
xnor U13273 (N_13273,N_12792,N_12828);
nor U13274 (N_13274,N_12721,N_12519);
xnor U13275 (N_13275,N_12710,N_12551);
or U13276 (N_13276,N_12796,N_12767);
or U13277 (N_13277,N_12608,N_12680);
or U13278 (N_13278,N_12745,N_12551);
nand U13279 (N_13279,N_12663,N_12582);
nand U13280 (N_13280,N_12915,N_12726);
nor U13281 (N_13281,N_12724,N_12835);
xor U13282 (N_13282,N_12762,N_12613);
nand U13283 (N_13283,N_12596,N_12950);
nand U13284 (N_13284,N_12776,N_12788);
xnor U13285 (N_13285,N_12801,N_12849);
nand U13286 (N_13286,N_12619,N_12637);
and U13287 (N_13287,N_12613,N_12784);
nand U13288 (N_13288,N_12575,N_12721);
xor U13289 (N_13289,N_12668,N_12877);
and U13290 (N_13290,N_12956,N_12751);
and U13291 (N_13291,N_12571,N_12681);
or U13292 (N_13292,N_12753,N_12671);
nor U13293 (N_13293,N_12993,N_12946);
nor U13294 (N_13294,N_12899,N_12811);
nor U13295 (N_13295,N_12785,N_12639);
and U13296 (N_13296,N_12744,N_12831);
nor U13297 (N_13297,N_12998,N_12531);
xor U13298 (N_13298,N_12688,N_12532);
xnor U13299 (N_13299,N_12739,N_12579);
and U13300 (N_13300,N_12587,N_12722);
or U13301 (N_13301,N_12725,N_12993);
nand U13302 (N_13302,N_12816,N_12787);
nand U13303 (N_13303,N_12529,N_12669);
nand U13304 (N_13304,N_12633,N_12689);
nor U13305 (N_13305,N_12753,N_12763);
xnor U13306 (N_13306,N_12702,N_12571);
or U13307 (N_13307,N_12860,N_12975);
or U13308 (N_13308,N_12692,N_12705);
and U13309 (N_13309,N_12671,N_12639);
nand U13310 (N_13310,N_12586,N_12571);
nor U13311 (N_13311,N_12924,N_12893);
and U13312 (N_13312,N_12759,N_12624);
or U13313 (N_13313,N_12547,N_12973);
xnor U13314 (N_13314,N_12756,N_12707);
or U13315 (N_13315,N_12832,N_12537);
and U13316 (N_13316,N_12812,N_12976);
nand U13317 (N_13317,N_12833,N_12942);
or U13318 (N_13318,N_12846,N_12829);
or U13319 (N_13319,N_12615,N_12558);
or U13320 (N_13320,N_12707,N_12632);
nor U13321 (N_13321,N_12925,N_12591);
nand U13322 (N_13322,N_12748,N_12890);
nor U13323 (N_13323,N_12869,N_12612);
or U13324 (N_13324,N_12806,N_12620);
and U13325 (N_13325,N_12667,N_12572);
and U13326 (N_13326,N_12677,N_12860);
or U13327 (N_13327,N_12611,N_12542);
nand U13328 (N_13328,N_12654,N_12796);
xor U13329 (N_13329,N_12508,N_12677);
xnor U13330 (N_13330,N_12762,N_12769);
xnor U13331 (N_13331,N_12670,N_12714);
xor U13332 (N_13332,N_12652,N_12915);
nor U13333 (N_13333,N_12965,N_12792);
nand U13334 (N_13334,N_12538,N_12924);
and U13335 (N_13335,N_12710,N_12523);
nor U13336 (N_13336,N_12844,N_12987);
nor U13337 (N_13337,N_12533,N_12632);
and U13338 (N_13338,N_12808,N_12524);
or U13339 (N_13339,N_12633,N_12808);
nand U13340 (N_13340,N_12932,N_12626);
nand U13341 (N_13341,N_12849,N_12700);
or U13342 (N_13342,N_12621,N_12577);
nor U13343 (N_13343,N_12544,N_12775);
nor U13344 (N_13344,N_12859,N_12690);
or U13345 (N_13345,N_12793,N_12901);
nand U13346 (N_13346,N_12782,N_12996);
nor U13347 (N_13347,N_12580,N_12837);
nand U13348 (N_13348,N_12858,N_12752);
nand U13349 (N_13349,N_12968,N_12520);
nor U13350 (N_13350,N_12819,N_12751);
and U13351 (N_13351,N_12989,N_12592);
xnor U13352 (N_13352,N_12663,N_12666);
or U13353 (N_13353,N_12794,N_12808);
and U13354 (N_13354,N_12717,N_12711);
and U13355 (N_13355,N_12526,N_12869);
xnor U13356 (N_13356,N_12691,N_12525);
nor U13357 (N_13357,N_12547,N_12677);
nor U13358 (N_13358,N_12667,N_12849);
xor U13359 (N_13359,N_12680,N_12503);
or U13360 (N_13360,N_12706,N_12660);
nor U13361 (N_13361,N_12742,N_12802);
and U13362 (N_13362,N_12543,N_12541);
and U13363 (N_13363,N_12548,N_12751);
or U13364 (N_13364,N_12612,N_12776);
or U13365 (N_13365,N_12740,N_12771);
nor U13366 (N_13366,N_12672,N_12706);
and U13367 (N_13367,N_12788,N_12855);
or U13368 (N_13368,N_12928,N_12867);
xnor U13369 (N_13369,N_12836,N_12941);
or U13370 (N_13370,N_12835,N_12515);
or U13371 (N_13371,N_12733,N_12625);
and U13372 (N_13372,N_12912,N_12516);
or U13373 (N_13373,N_12763,N_12715);
or U13374 (N_13374,N_12833,N_12790);
xnor U13375 (N_13375,N_12658,N_12880);
and U13376 (N_13376,N_12526,N_12893);
or U13377 (N_13377,N_12895,N_12960);
xnor U13378 (N_13378,N_12832,N_12503);
nand U13379 (N_13379,N_12890,N_12738);
and U13380 (N_13380,N_12959,N_12547);
nand U13381 (N_13381,N_12772,N_12830);
nor U13382 (N_13382,N_12969,N_12717);
or U13383 (N_13383,N_12953,N_12718);
and U13384 (N_13384,N_12565,N_12860);
or U13385 (N_13385,N_12985,N_12689);
nor U13386 (N_13386,N_12998,N_12791);
and U13387 (N_13387,N_12740,N_12970);
or U13388 (N_13388,N_12913,N_12564);
or U13389 (N_13389,N_12632,N_12713);
xor U13390 (N_13390,N_12543,N_12589);
xor U13391 (N_13391,N_12590,N_12739);
xnor U13392 (N_13392,N_12582,N_12951);
or U13393 (N_13393,N_12818,N_12507);
nor U13394 (N_13394,N_12610,N_12611);
and U13395 (N_13395,N_12790,N_12931);
nor U13396 (N_13396,N_12895,N_12657);
nor U13397 (N_13397,N_12663,N_12966);
nand U13398 (N_13398,N_12647,N_12526);
nor U13399 (N_13399,N_12785,N_12557);
and U13400 (N_13400,N_12807,N_12671);
nand U13401 (N_13401,N_12909,N_12649);
nand U13402 (N_13402,N_12646,N_12811);
nand U13403 (N_13403,N_12615,N_12961);
and U13404 (N_13404,N_12983,N_12695);
nand U13405 (N_13405,N_12789,N_12667);
nor U13406 (N_13406,N_12988,N_12778);
and U13407 (N_13407,N_12728,N_12545);
nor U13408 (N_13408,N_12896,N_12573);
or U13409 (N_13409,N_12920,N_12777);
xor U13410 (N_13410,N_12756,N_12892);
xnor U13411 (N_13411,N_12868,N_12965);
xor U13412 (N_13412,N_12894,N_12643);
nor U13413 (N_13413,N_12837,N_12855);
nor U13414 (N_13414,N_12631,N_12822);
xor U13415 (N_13415,N_12758,N_12536);
nand U13416 (N_13416,N_12659,N_12557);
or U13417 (N_13417,N_12849,N_12741);
nor U13418 (N_13418,N_12635,N_12830);
nor U13419 (N_13419,N_12953,N_12797);
and U13420 (N_13420,N_12833,N_12947);
or U13421 (N_13421,N_12995,N_12571);
nor U13422 (N_13422,N_12568,N_12519);
xor U13423 (N_13423,N_12933,N_12795);
xor U13424 (N_13424,N_12534,N_12732);
or U13425 (N_13425,N_12778,N_12589);
or U13426 (N_13426,N_12766,N_12660);
xnor U13427 (N_13427,N_12931,N_12743);
nand U13428 (N_13428,N_12602,N_12518);
or U13429 (N_13429,N_12853,N_12695);
nand U13430 (N_13430,N_12719,N_12507);
nand U13431 (N_13431,N_12709,N_12571);
and U13432 (N_13432,N_12770,N_12622);
nand U13433 (N_13433,N_12987,N_12646);
and U13434 (N_13434,N_12957,N_12617);
or U13435 (N_13435,N_12765,N_12911);
or U13436 (N_13436,N_12740,N_12845);
nand U13437 (N_13437,N_12584,N_12748);
nor U13438 (N_13438,N_12998,N_12950);
xor U13439 (N_13439,N_12952,N_12802);
nand U13440 (N_13440,N_12957,N_12846);
or U13441 (N_13441,N_12898,N_12595);
xnor U13442 (N_13442,N_12602,N_12977);
nand U13443 (N_13443,N_12822,N_12678);
xnor U13444 (N_13444,N_12619,N_12646);
or U13445 (N_13445,N_12725,N_12698);
nor U13446 (N_13446,N_12894,N_12786);
xor U13447 (N_13447,N_12928,N_12548);
or U13448 (N_13448,N_12763,N_12822);
nor U13449 (N_13449,N_12938,N_12701);
xnor U13450 (N_13450,N_12662,N_12618);
nor U13451 (N_13451,N_12775,N_12866);
and U13452 (N_13452,N_12971,N_12944);
nor U13453 (N_13453,N_12558,N_12886);
and U13454 (N_13454,N_12619,N_12743);
nand U13455 (N_13455,N_12879,N_12823);
nor U13456 (N_13456,N_12545,N_12599);
or U13457 (N_13457,N_12909,N_12615);
xnor U13458 (N_13458,N_12677,N_12930);
nand U13459 (N_13459,N_12677,N_12846);
xor U13460 (N_13460,N_12580,N_12855);
xor U13461 (N_13461,N_12924,N_12509);
nand U13462 (N_13462,N_12761,N_12591);
xor U13463 (N_13463,N_12652,N_12736);
or U13464 (N_13464,N_12959,N_12919);
and U13465 (N_13465,N_12800,N_12974);
or U13466 (N_13466,N_12599,N_12967);
nor U13467 (N_13467,N_12942,N_12771);
nand U13468 (N_13468,N_12773,N_12783);
or U13469 (N_13469,N_12851,N_12690);
nand U13470 (N_13470,N_12662,N_12745);
nor U13471 (N_13471,N_12984,N_12988);
xor U13472 (N_13472,N_12717,N_12771);
and U13473 (N_13473,N_12810,N_12792);
xnor U13474 (N_13474,N_12712,N_12508);
and U13475 (N_13475,N_12690,N_12548);
nand U13476 (N_13476,N_12951,N_12552);
nand U13477 (N_13477,N_12669,N_12678);
and U13478 (N_13478,N_12876,N_12746);
and U13479 (N_13479,N_12520,N_12635);
nor U13480 (N_13480,N_12505,N_12716);
nand U13481 (N_13481,N_12718,N_12913);
nand U13482 (N_13482,N_12896,N_12855);
nand U13483 (N_13483,N_12966,N_12853);
and U13484 (N_13484,N_12552,N_12523);
nor U13485 (N_13485,N_12864,N_12539);
nor U13486 (N_13486,N_12563,N_12620);
or U13487 (N_13487,N_12759,N_12630);
and U13488 (N_13488,N_12831,N_12693);
nor U13489 (N_13489,N_12778,N_12993);
and U13490 (N_13490,N_12663,N_12641);
or U13491 (N_13491,N_12612,N_12696);
xnor U13492 (N_13492,N_12739,N_12763);
nor U13493 (N_13493,N_12761,N_12613);
nand U13494 (N_13494,N_12887,N_12924);
nand U13495 (N_13495,N_12617,N_12598);
xnor U13496 (N_13496,N_12755,N_12658);
xnor U13497 (N_13497,N_12920,N_12764);
xnor U13498 (N_13498,N_12563,N_12855);
xnor U13499 (N_13499,N_12801,N_12507);
and U13500 (N_13500,N_13421,N_13489);
nand U13501 (N_13501,N_13416,N_13232);
and U13502 (N_13502,N_13316,N_13236);
nand U13503 (N_13503,N_13053,N_13064);
or U13504 (N_13504,N_13363,N_13433);
nor U13505 (N_13505,N_13076,N_13481);
nor U13506 (N_13506,N_13307,N_13122);
nor U13507 (N_13507,N_13067,N_13080);
or U13508 (N_13508,N_13235,N_13256);
xor U13509 (N_13509,N_13482,N_13066);
nor U13510 (N_13510,N_13400,N_13218);
xor U13511 (N_13511,N_13277,N_13303);
nand U13512 (N_13512,N_13128,N_13021);
nand U13513 (N_13513,N_13180,N_13099);
xnor U13514 (N_13514,N_13007,N_13205);
and U13515 (N_13515,N_13188,N_13000);
or U13516 (N_13516,N_13127,N_13250);
nand U13517 (N_13517,N_13019,N_13257);
nor U13518 (N_13518,N_13274,N_13030);
nor U13519 (N_13519,N_13430,N_13210);
or U13520 (N_13520,N_13005,N_13137);
or U13521 (N_13521,N_13154,N_13417);
and U13522 (N_13522,N_13260,N_13097);
xnor U13523 (N_13523,N_13114,N_13008);
nor U13524 (N_13524,N_13141,N_13254);
xor U13525 (N_13525,N_13468,N_13471);
xnor U13526 (N_13526,N_13388,N_13462);
nor U13527 (N_13527,N_13176,N_13085);
nor U13528 (N_13528,N_13365,N_13090);
and U13529 (N_13529,N_13164,N_13442);
and U13530 (N_13530,N_13144,N_13006);
or U13531 (N_13531,N_13174,N_13337);
nand U13532 (N_13532,N_13033,N_13161);
nor U13533 (N_13533,N_13116,N_13084);
xor U13534 (N_13534,N_13278,N_13439);
xnor U13535 (N_13535,N_13310,N_13179);
or U13536 (N_13536,N_13271,N_13317);
nor U13537 (N_13537,N_13418,N_13025);
and U13538 (N_13538,N_13301,N_13420);
and U13539 (N_13539,N_13268,N_13057);
xor U13540 (N_13540,N_13318,N_13121);
and U13541 (N_13541,N_13238,N_13491);
nand U13542 (N_13542,N_13496,N_13044);
or U13543 (N_13543,N_13294,N_13389);
xnor U13544 (N_13544,N_13133,N_13426);
and U13545 (N_13545,N_13447,N_13159);
xor U13546 (N_13546,N_13204,N_13039);
nor U13547 (N_13547,N_13275,N_13492);
xnor U13548 (N_13548,N_13403,N_13158);
or U13549 (N_13549,N_13056,N_13060);
and U13550 (N_13550,N_13225,N_13153);
xor U13551 (N_13551,N_13020,N_13049);
and U13552 (N_13552,N_13495,N_13217);
and U13553 (N_13553,N_13279,N_13356);
nor U13554 (N_13554,N_13382,N_13304);
xor U13555 (N_13555,N_13408,N_13051);
and U13556 (N_13556,N_13074,N_13374);
xnor U13557 (N_13557,N_13096,N_13211);
and U13558 (N_13558,N_13390,N_13229);
and U13559 (N_13559,N_13401,N_13034);
or U13560 (N_13560,N_13119,N_13379);
or U13561 (N_13561,N_13483,N_13252);
xnor U13562 (N_13562,N_13348,N_13415);
nand U13563 (N_13563,N_13023,N_13264);
xor U13564 (N_13564,N_13293,N_13283);
or U13565 (N_13565,N_13267,N_13460);
and U13566 (N_13566,N_13166,N_13290);
nand U13567 (N_13567,N_13367,N_13227);
and U13568 (N_13568,N_13427,N_13100);
nor U13569 (N_13569,N_13387,N_13436);
xnor U13570 (N_13570,N_13340,N_13344);
and U13571 (N_13571,N_13322,N_13215);
or U13572 (N_13572,N_13075,N_13043);
and U13573 (N_13573,N_13380,N_13109);
or U13574 (N_13574,N_13332,N_13308);
nor U13575 (N_13575,N_13172,N_13297);
and U13576 (N_13576,N_13086,N_13150);
or U13577 (N_13577,N_13376,N_13269);
nor U13578 (N_13578,N_13151,N_13233);
or U13579 (N_13579,N_13364,N_13328);
or U13580 (N_13580,N_13313,N_13031);
nand U13581 (N_13581,N_13476,N_13018);
xor U13582 (N_13582,N_13148,N_13146);
nand U13583 (N_13583,N_13342,N_13063);
or U13584 (N_13584,N_13231,N_13410);
nor U13585 (N_13585,N_13455,N_13047);
or U13586 (N_13586,N_13435,N_13406);
nand U13587 (N_13587,N_13444,N_13357);
and U13588 (N_13588,N_13014,N_13163);
and U13589 (N_13589,N_13138,N_13177);
nand U13590 (N_13590,N_13372,N_13386);
nand U13591 (N_13591,N_13486,N_13145);
and U13592 (N_13592,N_13123,N_13032);
and U13593 (N_13593,N_13465,N_13355);
xor U13594 (N_13594,N_13399,N_13253);
and U13595 (N_13595,N_13477,N_13350);
and U13596 (N_13596,N_13396,N_13368);
xor U13597 (N_13597,N_13326,N_13152);
and U13598 (N_13598,N_13422,N_13338);
nand U13599 (N_13599,N_13445,N_13249);
and U13600 (N_13600,N_13234,N_13016);
and U13601 (N_13601,N_13300,N_13201);
and U13602 (N_13602,N_13036,N_13089);
and U13603 (N_13603,N_13011,N_13200);
nand U13604 (N_13604,N_13393,N_13289);
and U13605 (N_13605,N_13391,N_13354);
nor U13606 (N_13606,N_13054,N_13149);
nor U13607 (N_13607,N_13309,N_13402);
nand U13608 (N_13608,N_13070,N_13347);
or U13609 (N_13609,N_13432,N_13125);
and U13610 (N_13610,N_13115,N_13212);
or U13611 (N_13611,N_13171,N_13194);
xnor U13612 (N_13612,N_13377,N_13078);
or U13613 (N_13613,N_13245,N_13373);
nand U13614 (N_13614,N_13286,N_13384);
nand U13615 (N_13615,N_13027,N_13330);
or U13616 (N_13616,N_13088,N_13428);
or U13617 (N_13617,N_13339,N_13366);
nand U13618 (N_13618,N_13052,N_13110);
or U13619 (N_13619,N_13198,N_13098);
nand U13620 (N_13620,N_13459,N_13397);
xor U13621 (N_13621,N_13108,N_13320);
nor U13622 (N_13622,N_13083,N_13265);
and U13623 (N_13623,N_13130,N_13321);
nand U13624 (N_13624,N_13038,N_13493);
and U13625 (N_13625,N_13228,N_13454);
and U13626 (N_13626,N_13017,N_13139);
or U13627 (N_13627,N_13395,N_13223);
nand U13628 (N_13628,N_13434,N_13214);
xnor U13629 (N_13629,N_13040,N_13494);
and U13630 (N_13630,N_13118,N_13453);
nor U13631 (N_13631,N_13336,N_13192);
and U13632 (N_13632,N_13319,N_13069);
and U13633 (N_13633,N_13299,N_13143);
xor U13634 (N_13634,N_13282,N_13498);
and U13635 (N_13635,N_13461,N_13246);
nor U13636 (N_13636,N_13302,N_13015);
nor U13637 (N_13637,N_13203,N_13315);
and U13638 (N_13638,N_13375,N_13305);
and U13639 (N_13639,N_13202,N_13082);
nor U13640 (N_13640,N_13136,N_13323);
nand U13641 (N_13641,N_13222,N_13142);
xor U13642 (N_13642,N_13026,N_13472);
nand U13643 (N_13643,N_13412,N_13487);
and U13644 (N_13644,N_13276,N_13263);
or U13645 (N_13645,N_13117,N_13104);
and U13646 (N_13646,N_13213,N_13475);
and U13647 (N_13647,N_13425,N_13126);
or U13648 (N_13648,N_13243,N_13424);
nor U13649 (N_13649,N_13371,N_13079);
xor U13650 (N_13650,N_13423,N_13346);
or U13651 (N_13651,N_13295,N_13009);
and U13652 (N_13652,N_13247,N_13189);
nor U13653 (N_13653,N_13361,N_13167);
nand U13654 (N_13654,N_13285,N_13292);
and U13655 (N_13655,N_13370,N_13062);
nand U13656 (N_13656,N_13258,N_13112);
nand U13657 (N_13657,N_13353,N_13010);
xnor U13658 (N_13658,N_13147,N_13464);
and U13659 (N_13659,N_13178,N_13497);
nor U13660 (N_13660,N_13446,N_13093);
or U13661 (N_13661,N_13207,N_13002);
nor U13662 (N_13662,N_13242,N_13448);
or U13663 (N_13663,N_13102,N_13383);
xnor U13664 (N_13664,N_13065,N_13441);
nand U13665 (N_13665,N_13480,N_13484);
and U13666 (N_13666,N_13124,N_13129);
or U13667 (N_13667,N_13029,N_13012);
nand U13668 (N_13668,N_13187,N_13071);
nand U13669 (N_13669,N_13132,N_13022);
xor U13670 (N_13670,N_13013,N_13091);
or U13671 (N_13671,N_13061,N_13473);
nor U13672 (N_13672,N_13429,N_13081);
and U13673 (N_13673,N_13345,N_13329);
or U13674 (N_13674,N_13437,N_13284);
xnor U13675 (N_13675,N_13073,N_13479);
and U13676 (N_13676,N_13381,N_13255);
nor U13677 (N_13677,N_13281,N_13199);
or U13678 (N_13678,N_13259,N_13398);
or U13679 (N_13679,N_13162,N_13248);
nand U13680 (N_13680,N_13237,N_13343);
nand U13681 (N_13681,N_13131,N_13358);
or U13682 (N_13682,N_13298,N_13490);
and U13683 (N_13683,N_13443,N_13287);
or U13684 (N_13684,N_13270,N_13160);
xnor U13685 (N_13685,N_13107,N_13120);
nand U13686 (N_13686,N_13157,N_13470);
nand U13687 (N_13687,N_13488,N_13431);
nand U13688 (N_13688,N_13226,N_13469);
nand U13689 (N_13689,N_13195,N_13452);
nand U13690 (N_13690,N_13466,N_13208);
nand U13691 (N_13691,N_13186,N_13048);
xnor U13692 (N_13692,N_13059,N_13407);
or U13693 (N_13693,N_13334,N_13156);
xnor U13694 (N_13694,N_13306,N_13113);
and U13695 (N_13695,N_13405,N_13001);
xor U13696 (N_13696,N_13419,N_13457);
nand U13697 (N_13697,N_13003,N_13272);
nor U13698 (N_13698,N_13209,N_13134);
nor U13699 (N_13699,N_13037,N_13499);
nand U13700 (N_13700,N_13467,N_13335);
xnor U13701 (N_13701,N_13224,N_13450);
xnor U13702 (N_13702,N_13411,N_13280);
or U13703 (N_13703,N_13392,N_13463);
nor U13704 (N_13704,N_13474,N_13193);
and U13705 (N_13705,N_13378,N_13312);
and U13706 (N_13706,N_13165,N_13413);
xor U13707 (N_13707,N_13058,N_13333);
nor U13708 (N_13708,N_13101,N_13055);
and U13709 (N_13709,N_13291,N_13414);
nand U13710 (N_13710,N_13095,N_13028);
and U13711 (N_13711,N_13311,N_13077);
or U13712 (N_13712,N_13216,N_13197);
or U13713 (N_13713,N_13351,N_13169);
nor U13714 (N_13714,N_13325,N_13103);
nand U13715 (N_13715,N_13106,N_13349);
nor U13716 (N_13716,N_13324,N_13087);
and U13717 (N_13717,N_13362,N_13296);
nor U13718 (N_13718,N_13045,N_13266);
nor U13719 (N_13719,N_13105,N_13182);
and U13720 (N_13720,N_13314,N_13241);
xor U13721 (N_13721,N_13394,N_13220);
or U13722 (N_13722,N_13206,N_13240);
xor U13723 (N_13723,N_13183,N_13331);
xor U13724 (N_13724,N_13181,N_13185);
or U13725 (N_13725,N_13341,N_13404);
xor U13726 (N_13726,N_13004,N_13478);
xnor U13727 (N_13727,N_13173,N_13170);
xor U13728 (N_13728,N_13359,N_13244);
and U13729 (N_13729,N_13327,N_13438);
or U13730 (N_13730,N_13094,N_13369);
xor U13731 (N_13731,N_13440,N_13042);
and U13732 (N_13732,N_13135,N_13262);
nor U13733 (N_13733,N_13092,N_13352);
nand U13734 (N_13734,N_13024,N_13168);
nor U13735 (N_13735,N_13458,N_13111);
nand U13736 (N_13736,N_13449,N_13261);
xnor U13737 (N_13737,N_13190,N_13251);
or U13738 (N_13738,N_13196,N_13219);
and U13739 (N_13739,N_13046,N_13230);
nand U13740 (N_13740,N_13385,N_13155);
or U13741 (N_13741,N_13485,N_13451);
nand U13742 (N_13742,N_13041,N_13221);
nor U13743 (N_13743,N_13456,N_13273);
or U13744 (N_13744,N_13191,N_13239);
and U13745 (N_13745,N_13175,N_13288);
and U13746 (N_13746,N_13409,N_13360);
and U13747 (N_13747,N_13184,N_13050);
xor U13748 (N_13748,N_13035,N_13068);
and U13749 (N_13749,N_13072,N_13140);
nand U13750 (N_13750,N_13228,N_13238);
and U13751 (N_13751,N_13026,N_13392);
nand U13752 (N_13752,N_13101,N_13094);
nor U13753 (N_13753,N_13311,N_13225);
nor U13754 (N_13754,N_13440,N_13050);
nand U13755 (N_13755,N_13083,N_13158);
and U13756 (N_13756,N_13407,N_13388);
and U13757 (N_13757,N_13004,N_13279);
or U13758 (N_13758,N_13483,N_13247);
and U13759 (N_13759,N_13222,N_13093);
nand U13760 (N_13760,N_13027,N_13205);
and U13761 (N_13761,N_13317,N_13302);
nor U13762 (N_13762,N_13074,N_13184);
nand U13763 (N_13763,N_13324,N_13343);
or U13764 (N_13764,N_13429,N_13431);
xnor U13765 (N_13765,N_13034,N_13379);
nor U13766 (N_13766,N_13080,N_13254);
nand U13767 (N_13767,N_13478,N_13038);
nand U13768 (N_13768,N_13253,N_13431);
nand U13769 (N_13769,N_13025,N_13055);
and U13770 (N_13770,N_13385,N_13070);
nor U13771 (N_13771,N_13265,N_13353);
or U13772 (N_13772,N_13487,N_13041);
and U13773 (N_13773,N_13366,N_13234);
and U13774 (N_13774,N_13340,N_13117);
nor U13775 (N_13775,N_13426,N_13224);
nor U13776 (N_13776,N_13241,N_13088);
or U13777 (N_13777,N_13369,N_13346);
nand U13778 (N_13778,N_13457,N_13331);
and U13779 (N_13779,N_13406,N_13099);
and U13780 (N_13780,N_13264,N_13416);
xnor U13781 (N_13781,N_13176,N_13242);
nor U13782 (N_13782,N_13380,N_13143);
xnor U13783 (N_13783,N_13428,N_13386);
nor U13784 (N_13784,N_13050,N_13436);
and U13785 (N_13785,N_13246,N_13176);
nand U13786 (N_13786,N_13451,N_13004);
xor U13787 (N_13787,N_13057,N_13223);
xnor U13788 (N_13788,N_13251,N_13024);
xnor U13789 (N_13789,N_13251,N_13423);
nand U13790 (N_13790,N_13495,N_13403);
xor U13791 (N_13791,N_13382,N_13034);
nor U13792 (N_13792,N_13240,N_13344);
and U13793 (N_13793,N_13066,N_13275);
nor U13794 (N_13794,N_13209,N_13083);
or U13795 (N_13795,N_13306,N_13446);
nand U13796 (N_13796,N_13125,N_13045);
and U13797 (N_13797,N_13289,N_13435);
nand U13798 (N_13798,N_13180,N_13114);
nand U13799 (N_13799,N_13383,N_13226);
or U13800 (N_13800,N_13033,N_13024);
and U13801 (N_13801,N_13235,N_13133);
and U13802 (N_13802,N_13196,N_13485);
nor U13803 (N_13803,N_13445,N_13105);
nor U13804 (N_13804,N_13128,N_13462);
or U13805 (N_13805,N_13036,N_13163);
or U13806 (N_13806,N_13088,N_13167);
nand U13807 (N_13807,N_13032,N_13163);
xnor U13808 (N_13808,N_13170,N_13460);
nor U13809 (N_13809,N_13363,N_13106);
nor U13810 (N_13810,N_13401,N_13451);
nand U13811 (N_13811,N_13466,N_13113);
and U13812 (N_13812,N_13295,N_13086);
or U13813 (N_13813,N_13256,N_13371);
xor U13814 (N_13814,N_13469,N_13141);
and U13815 (N_13815,N_13146,N_13462);
nand U13816 (N_13816,N_13472,N_13180);
or U13817 (N_13817,N_13387,N_13112);
and U13818 (N_13818,N_13314,N_13083);
nor U13819 (N_13819,N_13423,N_13096);
xnor U13820 (N_13820,N_13083,N_13197);
nor U13821 (N_13821,N_13022,N_13030);
nand U13822 (N_13822,N_13040,N_13124);
and U13823 (N_13823,N_13381,N_13002);
and U13824 (N_13824,N_13288,N_13493);
xor U13825 (N_13825,N_13137,N_13104);
and U13826 (N_13826,N_13078,N_13181);
nor U13827 (N_13827,N_13408,N_13305);
xnor U13828 (N_13828,N_13464,N_13363);
or U13829 (N_13829,N_13062,N_13051);
nor U13830 (N_13830,N_13330,N_13224);
xor U13831 (N_13831,N_13099,N_13326);
nand U13832 (N_13832,N_13441,N_13009);
or U13833 (N_13833,N_13455,N_13218);
nand U13834 (N_13834,N_13441,N_13004);
xor U13835 (N_13835,N_13131,N_13081);
or U13836 (N_13836,N_13322,N_13098);
and U13837 (N_13837,N_13427,N_13405);
nor U13838 (N_13838,N_13163,N_13489);
and U13839 (N_13839,N_13212,N_13492);
nand U13840 (N_13840,N_13066,N_13311);
or U13841 (N_13841,N_13028,N_13258);
nor U13842 (N_13842,N_13411,N_13072);
xnor U13843 (N_13843,N_13082,N_13298);
or U13844 (N_13844,N_13428,N_13352);
or U13845 (N_13845,N_13171,N_13448);
nand U13846 (N_13846,N_13468,N_13042);
nor U13847 (N_13847,N_13221,N_13209);
nand U13848 (N_13848,N_13160,N_13387);
nor U13849 (N_13849,N_13328,N_13283);
nand U13850 (N_13850,N_13287,N_13377);
and U13851 (N_13851,N_13471,N_13329);
or U13852 (N_13852,N_13278,N_13093);
and U13853 (N_13853,N_13477,N_13386);
nor U13854 (N_13854,N_13032,N_13139);
or U13855 (N_13855,N_13382,N_13255);
or U13856 (N_13856,N_13490,N_13198);
xnor U13857 (N_13857,N_13154,N_13348);
and U13858 (N_13858,N_13242,N_13335);
xnor U13859 (N_13859,N_13089,N_13063);
nand U13860 (N_13860,N_13112,N_13142);
nand U13861 (N_13861,N_13007,N_13170);
nand U13862 (N_13862,N_13165,N_13466);
and U13863 (N_13863,N_13118,N_13010);
nand U13864 (N_13864,N_13294,N_13371);
xnor U13865 (N_13865,N_13110,N_13289);
and U13866 (N_13866,N_13068,N_13415);
and U13867 (N_13867,N_13437,N_13039);
or U13868 (N_13868,N_13286,N_13196);
or U13869 (N_13869,N_13026,N_13432);
or U13870 (N_13870,N_13165,N_13305);
nand U13871 (N_13871,N_13280,N_13028);
or U13872 (N_13872,N_13199,N_13496);
and U13873 (N_13873,N_13229,N_13054);
or U13874 (N_13874,N_13066,N_13087);
nand U13875 (N_13875,N_13225,N_13124);
nor U13876 (N_13876,N_13319,N_13267);
nand U13877 (N_13877,N_13183,N_13444);
nor U13878 (N_13878,N_13435,N_13019);
or U13879 (N_13879,N_13022,N_13434);
nand U13880 (N_13880,N_13052,N_13450);
or U13881 (N_13881,N_13367,N_13264);
xor U13882 (N_13882,N_13115,N_13012);
xnor U13883 (N_13883,N_13070,N_13283);
xnor U13884 (N_13884,N_13232,N_13300);
or U13885 (N_13885,N_13274,N_13459);
or U13886 (N_13886,N_13167,N_13285);
and U13887 (N_13887,N_13032,N_13054);
and U13888 (N_13888,N_13477,N_13299);
nor U13889 (N_13889,N_13253,N_13494);
nor U13890 (N_13890,N_13046,N_13323);
nand U13891 (N_13891,N_13050,N_13276);
xnor U13892 (N_13892,N_13014,N_13251);
nor U13893 (N_13893,N_13042,N_13169);
or U13894 (N_13894,N_13396,N_13023);
or U13895 (N_13895,N_13210,N_13033);
and U13896 (N_13896,N_13042,N_13230);
nor U13897 (N_13897,N_13261,N_13087);
nor U13898 (N_13898,N_13234,N_13015);
xor U13899 (N_13899,N_13407,N_13473);
or U13900 (N_13900,N_13382,N_13201);
nand U13901 (N_13901,N_13028,N_13212);
nand U13902 (N_13902,N_13141,N_13207);
nand U13903 (N_13903,N_13314,N_13353);
nand U13904 (N_13904,N_13409,N_13008);
nor U13905 (N_13905,N_13301,N_13021);
nand U13906 (N_13906,N_13205,N_13294);
or U13907 (N_13907,N_13488,N_13250);
nand U13908 (N_13908,N_13000,N_13483);
nand U13909 (N_13909,N_13076,N_13150);
and U13910 (N_13910,N_13238,N_13442);
xnor U13911 (N_13911,N_13162,N_13367);
nand U13912 (N_13912,N_13168,N_13331);
nand U13913 (N_13913,N_13043,N_13182);
nor U13914 (N_13914,N_13056,N_13157);
nor U13915 (N_13915,N_13202,N_13105);
and U13916 (N_13916,N_13012,N_13161);
or U13917 (N_13917,N_13108,N_13216);
or U13918 (N_13918,N_13225,N_13396);
xor U13919 (N_13919,N_13336,N_13154);
xor U13920 (N_13920,N_13478,N_13212);
nand U13921 (N_13921,N_13296,N_13087);
nand U13922 (N_13922,N_13066,N_13211);
and U13923 (N_13923,N_13228,N_13292);
nor U13924 (N_13924,N_13400,N_13459);
nor U13925 (N_13925,N_13056,N_13430);
xor U13926 (N_13926,N_13272,N_13101);
xor U13927 (N_13927,N_13417,N_13447);
and U13928 (N_13928,N_13396,N_13034);
or U13929 (N_13929,N_13044,N_13250);
and U13930 (N_13930,N_13178,N_13087);
nand U13931 (N_13931,N_13228,N_13264);
nor U13932 (N_13932,N_13222,N_13006);
nor U13933 (N_13933,N_13087,N_13312);
nor U13934 (N_13934,N_13394,N_13051);
nand U13935 (N_13935,N_13239,N_13235);
xor U13936 (N_13936,N_13419,N_13078);
or U13937 (N_13937,N_13478,N_13048);
nand U13938 (N_13938,N_13077,N_13137);
xor U13939 (N_13939,N_13246,N_13335);
nor U13940 (N_13940,N_13236,N_13357);
and U13941 (N_13941,N_13366,N_13368);
and U13942 (N_13942,N_13167,N_13405);
nor U13943 (N_13943,N_13286,N_13335);
xor U13944 (N_13944,N_13292,N_13210);
xnor U13945 (N_13945,N_13187,N_13042);
nand U13946 (N_13946,N_13167,N_13115);
xnor U13947 (N_13947,N_13433,N_13249);
and U13948 (N_13948,N_13402,N_13056);
or U13949 (N_13949,N_13213,N_13286);
xnor U13950 (N_13950,N_13485,N_13300);
and U13951 (N_13951,N_13133,N_13266);
nor U13952 (N_13952,N_13181,N_13321);
nor U13953 (N_13953,N_13327,N_13494);
and U13954 (N_13954,N_13100,N_13073);
and U13955 (N_13955,N_13377,N_13013);
nor U13956 (N_13956,N_13477,N_13383);
and U13957 (N_13957,N_13145,N_13344);
nand U13958 (N_13958,N_13270,N_13361);
nand U13959 (N_13959,N_13489,N_13115);
and U13960 (N_13960,N_13125,N_13235);
nor U13961 (N_13961,N_13146,N_13493);
or U13962 (N_13962,N_13189,N_13296);
or U13963 (N_13963,N_13104,N_13143);
xor U13964 (N_13964,N_13000,N_13485);
nand U13965 (N_13965,N_13496,N_13209);
and U13966 (N_13966,N_13227,N_13080);
nand U13967 (N_13967,N_13400,N_13267);
nor U13968 (N_13968,N_13276,N_13429);
nand U13969 (N_13969,N_13316,N_13224);
xnor U13970 (N_13970,N_13265,N_13392);
xnor U13971 (N_13971,N_13007,N_13402);
nand U13972 (N_13972,N_13042,N_13330);
and U13973 (N_13973,N_13497,N_13195);
xnor U13974 (N_13974,N_13305,N_13236);
and U13975 (N_13975,N_13189,N_13374);
nand U13976 (N_13976,N_13031,N_13370);
nor U13977 (N_13977,N_13418,N_13469);
or U13978 (N_13978,N_13429,N_13069);
or U13979 (N_13979,N_13037,N_13498);
nand U13980 (N_13980,N_13414,N_13313);
nor U13981 (N_13981,N_13127,N_13287);
or U13982 (N_13982,N_13187,N_13325);
and U13983 (N_13983,N_13472,N_13488);
or U13984 (N_13984,N_13303,N_13422);
or U13985 (N_13985,N_13272,N_13251);
nand U13986 (N_13986,N_13059,N_13284);
nor U13987 (N_13987,N_13433,N_13209);
xnor U13988 (N_13988,N_13071,N_13003);
or U13989 (N_13989,N_13373,N_13042);
or U13990 (N_13990,N_13025,N_13290);
nand U13991 (N_13991,N_13441,N_13488);
nand U13992 (N_13992,N_13332,N_13224);
nor U13993 (N_13993,N_13071,N_13402);
or U13994 (N_13994,N_13399,N_13114);
or U13995 (N_13995,N_13433,N_13296);
or U13996 (N_13996,N_13466,N_13051);
and U13997 (N_13997,N_13432,N_13350);
xnor U13998 (N_13998,N_13267,N_13487);
nand U13999 (N_13999,N_13095,N_13470);
nor U14000 (N_14000,N_13580,N_13690);
nand U14001 (N_14001,N_13950,N_13696);
and U14002 (N_14002,N_13832,N_13612);
nor U14003 (N_14003,N_13531,N_13662);
xor U14004 (N_14004,N_13562,N_13740);
or U14005 (N_14005,N_13719,N_13659);
or U14006 (N_14006,N_13536,N_13835);
or U14007 (N_14007,N_13958,N_13547);
nor U14008 (N_14008,N_13848,N_13882);
and U14009 (N_14009,N_13657,N_13729);
or U14010 (N_14010,N_13801,N_13620);
and U14011 (N_14011,N_13557,N_13791);
nand U14012 (N_14012,N_13626,N_13676);
nor U14013 (N_14013,N_13826,N_13649);
and U14014 (N_14014,N_13522,N_13820);
or U14015 (N_14015,N_13936,N_13877);
xnor U14016 (N_14016,N_13955,N_13571);
nand U14017 (N_14017,N_13900,N_13831);
nor U14018 (N_14018,N_13697,N_13583);
and U14019 (N_14019,N_13504,N_13737);
and U14020 (N_14020,N_13681,N_13703);
or U14021 (N_14021,N_13718,N_13741);
xnor U14022 (N_14022,N_13714,N_13810);
and U14023 (N_14023,N_13734,N_13559);
nand U14024 (N_14024,N_13691,N_13969);
or U14025 (N_14025,N_13869,N_13646);
or U14026 (N_14026,N_13995,N_13596);
or U14027 (N_14027,N_13710,N_13767);
and U14028 (N_14028,N_13605,N_13518);
or U14029 (N_14029,N_13752,N_13813);
and U14030 (N_14030,N_13927,N_13806);
nor U14031 (N_14031,N_13725,N_13683);
xnor U14032 (N_14032,N_13787,N_13949);
or U14033 (N_14033,N_13852,N_13985);
nand U14034 (N_14034,N_13759,N_13713);
nor U14035 (N_14035,N_13712,N_13903);
or U14036 (N_14036,N_13513,N_13598);
or U14037 (N_14037,N_13622,N_13753);
nor U14038 (N_14038,N_13867,N_13977);
nand U14039 (N_14039,N_13802,N_13998);
nor U14040 (N_14040,N_13883,N_13669);
xnor U14041 (N_14041,N_13749,N_13613);
xor U14042 (N_14042,N_13763,N_13823);
nand U14043 (N_14043,N_13671,N_13754);
nor U14044 (N_14044,N_13644,N_13542);
nor U14045 (N_14045,N_13785,N_13871);
or U14046 (N_14046,N_13680,N_13979);
nand U14047 (N_14047,N_13567,N_13807);
or U14048 (N_14048,N_13684,N_13630);
and U14049 (N_14049,N_13606,N_13940);
or U14050 (N_14050,N_13842,N_13670);
or U14051 (N_14051,N_13973,N_13610);
and U14052 (N_14052,N_13677,N_13849);
and U14053 (N_14053,N_13821,N_13739);
and U14054 (N_14054,N_13730,N_13541);
or U14055 (N_14055,N_13993,N_13937);
and U14056 (N_14056,N_13561,N_13830);
xnor U14057 (N_14057,N_13614,N_13885);
and U14058 (N_14058,N_13588,N_13625);
or U14059 (N_14059,N_13535,N_13576);
xor U14060 (N_14060,N_13500,N_13627);
and U14061 (N_14061,N_13653,N_13912);
and U14062 (N_14062,N_13575,N_13716);
or U14063 (N_14063,N_13947,N_13794);
or U14064 (N_14064,N_13892,N_13584);
and U14065 (N_14065,N_13896,N_13976);
xor U14066 (N_14066,N_13984,N_13824);
nor U14067 (N_14067,N_13724,N_13827);
nand U14068 (N_14068,N_13895,N_13796);
nor U14069 (N_14069,N_13861,N_13915);
nand U14070 (N_14070,N_13743,N_13774);
or U14071 (N_14071,N_13768,N_13881);
nor U14072 (N_14072,N_13540,N_13582);
xnor U14073 (N_14073,N_13530,N_13616);
nor U14074 (N_14074,N_13579,N_13551);
or U14075 (N_14075,N_13964,N_13890);
xor U14076 (N_14076,N_13901,N_13524);
nor U14077 (N_14077,N_13589,N_13933);
and U14078 (N_14078,N_13889,N_13856);
xnor U14079 (N_14079,N_13899,N_13760);
or U14080 (N_14080,N_13814,N_13917);
nor U14081 (N_14081,N_13640,N_13845);
or U14082 (N_14082,N_13790,N_13516);
xnor U14083 (N_14083,N_13980,N_13968);
xor U14084 (N_14084,N_13502,N_13913);
xor U14085 (N_14085,N_13988,N_13641);
xnor U14086 (N_14086,N_13747,N_13593);
or U14087 (N_14087,N_13688,N_13778);
and U14088 (N_14088,N_13506,N_13943);
nor U14089 (N_14089,N_13986,N_13717);
nand U14090 (N_14090,N_13898,N_13772);
nor U14091 (N_14091,N_13991,N_13636);
xnor U14092 (N_14092,N_13639,N_13928);
nand U14093 (N_14093,N_13581,N_13971);
and U14094 (N_14094,N_13954,N_13565);
or U14095 (N_14095,N_13634,N_13672);
nor U14096 (N_14096,N_13544,N_13638);
xor U14097 (N_14097,N_13577,N_13800);
nand U14098 (N_14098,N_13833,N_13545);
nor U14099 (N_14099,N_13843,N_13891);
or U14100 (N_14100,N_13929,N_13918);
and U14101 (N_14101,N_13909,N_13548);
nor U14102 (N_14102,N_13893,N_13678);
nand U14103 (N_14103,N_13699,N_13533);
or U14104 (N_14104,N_13837,N_13698);
nand U14105 (N_14105,N_13797,N_13897);
nand U14106 (N_14106,N_13687,N_13878);
nor U14107 (N_14107,N_13569,N_13799);
and U14108 (N_14108,N_13910,N_13534);
xor U14109 (N_14109,N_13628,N_13925);
and U14110 (N_14110,N_13758,N_13857);
xnor U14111 (N_14111,N_13674,N_13864);
nor U14112 (N_14112,N_13963,N_13686);
or U14113 (N_14113,N_13709,N_13553);
and U14114 (N_14114,N_13563,N_13959);
or U14115 (N_14115,N_13961,N_13818);
or U14116 (N_14116,N_13609,N_13967);
nor U14117 (N_14117,N_13668,N_13834);
and U14118 (N_14118,N_13602,N_13815);
nor U14119 (N_14119,N_13994,N_13956);
xnor U14120 (N_14120,N_13789,N_13860);
xnor U14121 (N_14121,N_13523,N_13769);
or U14122 (N_14122,N_13804,N_13507);
xor U14123 (N_14123,N_13922,N_13989);
or U14124 (N_14124,N_13706,N_13761);
nand U14125 (N_14125,N_13786,N_13597);
and U14126 (N_14126,N_13733,N_13855);
xnor U14127 (N_14127,N_13951,N_13920);
nor U14128 (N_14128,N_13766,N_13708);
or U14129 (N_14129,N_13735,N_13750);
and U14130 (N_14130,N_13811,N_13930);
or U14131 (N_14131,N_13911,N_13679);
and U14132 (N_14132,N_13650,N_13519);
or U14133 (N_14133,N_13600,N_13720);
nand U14134 (N_14134,N_13742,N_13643);
and U14135 (N_14135,N_13608,N_13793);
nor U14136 (N_14136,N_13721,N_13983);
or U14137 (N_14137,N_13965,N_13603);
and U14138 (N_14138,N_13923,N_13558);
or U14139 (N_14139,N_13746,N_13525);
xor U14140 (N_14140,N_13623,N_13512);
nor U14141 (N_14141,N_13654,N_13941);
nor U14142 (N_14142,N_13874,N_13660);
or U14143 (N_14143,N_13744,N_13945);
or U14144 (N_14144,N_13722,N_13546);
nor U14145 (N_14145,N_13919,N_13550);
and U14146 (N_14146,N_13745,N_13887);
nand U14147 (N_14147,N_13798,N_13817);
nand U14148 (N_14148,N_13854,N_13585);
xnor U14149 (N_14149,N_13549,N_13664);
and U14150 (N_14150,N_13829,N_13972);
nand U14151 (N_14151,N_13607,N_13702);
xnor U14152 (N_14152,N_13942,N_13731);
nand U14153 (N_14153,N_13776,N_13999);
nand U14154 (N_14154,N_13902,N_13946);
xnor U14155 (N_14155,N_13554,N_13858);
nand U14156 (N_14156,N_13701,N_13822);
nor U14157 (N_14157,N_13665,N_13884);
nor U14158 (N_14158,N_13953,N_13651);
or U14159 (N_14159,N_13652,N_13894);
or U14160 (N_14160,N_13962,N_13886);
or U14161 (N_14161,N_13591,N_13592);
or U14162 (N_14162,N_13921,N_13604);
and U14163 (N_14163,N_13944,N_13594);
nor U14164 (N_14164,N_13990,N_13632);
nand U14165 (N_14165,N_13635,N_13952);
or U14166 (N_14166,N_13538,N_13556);
xnor U14167 (N_14167,N_13624,N_13700);
nand U14168 (N_14168,N_13847,N_13841);
nor U14169 (N_14169,N_13779,N_13570);
xnor U14170 (N_14170,N_13783,N_13511);
nand U14171 (N_14171,N_13738,N_13875);
nand U14172 (N_14172,N_13808,N_13532);
nor U14173 (N_14173,N_13528,N_13693);
nor U14174 (N_14174,N_13595,N_13906);
or U14175 (N_14175,N_13888,N_13846);
xor U14176 (N_14176,N_13865,N_13501);
nor U14177 (N_14177,N_13658,N_13982);
and U14178 (N_14178,N_13568,N_13552);
and U14179 (N_14179,N_13788,N_13844);
xor U14180 (N_14180,N_13764,N_13819);
nor U14181 (N_14181,N_13924,N_13862);
nand U14182 (N_14182,N_13715,N_13876);
or U14183 (N_14183,N_13615,N_13560);
nor U14184 (N_14184,N_13656,N_13880);
and U14185 (N_14185,N_13859,N_13838);
xor U14186 (N_14186,N_13939,N_13762);
xnor U14187 (N_14187,N_13637,N_13723);
nand U14188 (N_14188,N_13966,N_13618);
or U14189 (N_14189,N_13932,N_13564);
nand U14190 (N_14190,N_13572,N_13689);
or U14191 (N_14191,N_13780,N_13851);
and U14192 (N_14192,N_13773,N_13514);
or U14193 (N_14193,N_13825,N_13647);
and U14194 (N_14194,N_13732,N_13704);
nor U14195 (N_14195,N_13621,N_13601);
xor U14196 (N_14196,N_13926,N_13836);
nand U14197 (N_14197,N_13795,N_13587);
nor U14198 (N_14198,N_13711,N_13782);
or U14199 (N_14199,N_13960,N_13775);
nor U14200 (N_14200,N_13685,N_13997);
nor U14201 (N_14201,N_13992,N_13777);
and U14202 (N_14202,N_13853,N_13505);
or U14203 (N_14203,N_13840,N_13539);
or U14204 (N_14204,N_13996,N_13629);
and U14205 (N_14205,N_13537,N_13934);
and U14206 (N_14206,N_13633,N_13515);
nor U14207 (N_14207,N_13916,N_13663);
nand U14208 (N_14208,N_13978,N_13908);
and U14209 (N_14209,N_13520,N_13736);
xor U14210 (N_14210,N_13529,N_13682);
nor U14211 (N_14211,N_13673,N_13757);
nand U14212 (N_14212,N_13509,N_13642);
nor U14213 (N_14213,N_13508,N_13948);
nor U14214 (N_14214,N_13599,N_13879);
and U14215 (N_14215,N_13905,N_13648);
and U14216 (N_14216,N_13617,N_13667);
or U14217 (N_14217,N_13974,N_13527);
and U14218 (N_14218,N_13694,N_13850);
nand U14219 (N_14219,N_13931,N_13770);
nor U14220 (N_14220,N_13792,N_13816);
or U14221 (N_14221,N_13503,N_13521);
xor U14222 (N_14222,N_13866,N_13828);
nor U14223 (N_14223,N_13870,N_13765);
nand U14224 (N_14224,N_13987,N_13755);
nand U14225 (N_14225,N_13873,N_13872);
nor U14226 (N_14226,N_13981,N_13543);
nor U14227 (N_14227,N_13590,N_13611);
nand U14228 (N_14228,N_13812,N_13661);
xnor U14229 (N_14229,N_13868,N_13707);
nand U14230 (N_14230,N_13573,N_13631);
nor U14231 (N_14231,N_13695,N_13957);
nor U14232 (N_14232,N_13526,N_13784);
xnor U14233 (N_14233,N_13619,N_13510);
and U14234 (N_14234,N_13578,N_13938);
xnor U14235 (N_14235,N_13809,N_13803);
nand U14236 (N_14236,N_13655,N_13839);
or U14237 (N_14237,N_13645,N_13975);
nand U14238 (N_14238,N_13692,N_13675);
or U14239 (N_14239,N_13756,N_13805);
nand U14240 (N_14240,N_13781,N_13727);
and U14241 (N_14241,N_13935,N_13863);
nor U14242 (N_14242,N_13728,N_13705);
or U14243 (N_14243,N_13751,N_13748);
nor U14244 (N_14244,N_13904,N_13914);
nand U14245 (N_14245,N_13517,N_13907);
or U14246 (N_14246,N_13666,N_13726);
nor U14247 (N_14247,N_13566,N_13970);
nor U14248 (N_14248,N_13586,N_13574);
nor U14249 (N_14249,N_13555,N_13771);
xor U14250 (N_14250,N_13601,N_13668);
and U14251 (N_14251,N_13817,N_13593);
nor U14252 (N_14252,N_13934,N_13673);
and U14253 (N_14253,N_13508,N_13828);
xnor U14254 (N_14254,N_13521,N_13653);
xnor U14255 (N_14255,N_13883,N_13641);
or U14256 (N_14256,N_13603,N_13749);
or U14257 (N_14257,N_13782,N_13666);
xor U14258 (N_14258,N_13542,N_13967);
and U14259 (N_14259,N_13831,N_13710);
or U14260 (N_14260,N_13610,N_13902);
nor U14261 (N_14261,N_13927,N_13660);
or U14262 (N_14262,N_13600,N_13654);
or U14263 (N_14263,N_13904,N_13748);
xnor U14264 (N_14264,N_13600,N_13966);
or U14265 (N_14265,N_13973,N_13844);
xor U14266 (N_14266,N_13978,N_13551);
and U14267 (N_14267,N_13868,N_13768);
nand U14268 (N_14268,N_13777,N_13873);
or U14269 (N_14269,N_13572,N_13749);
nand U14270 (N_14270,N_13756,N_13936);
xor U14271 (N_14271,N_13964,N_13955);
and U14272 (N_14272,N_13581,N_13746);
or U14273 (N_14273,N_13810,N_13977);
xnor U14274 (N_14274,N_13690,N_13707);
nor U14275 (N_14275,N_13567,N_13766);
nand U14276 (N_14276,N_13868,N_13627);
or U14277 (N_14277,N_13589,N_13697);
or U14278 (N_14278,N_13772,N_13906);
nor U14279 (N_14279,N_13947,N_13537);
or U14280 (N_14280,N_13605,N_13896);
xnor U14281 (N_14281,N_13706,N_13651);
and U14282 (N_14282,N_13979,N_13992);
xnor U14283 (N_14283,N_13573,N_13952);
nor U14284 (N_14284,N_13863,N_13737);
nor U14285 (N_14285,N_13934,N_13936);
xnor U14286 (N_14286,N_13758,N_13601);
nor U14287 (N_14287,N_13593,N_13939);
nor U14288 (N_14288,N_13885,N_13554);
xor U14289 (N_14289,N_13595,N_13997);
nand U14290 (N_14290,N_13536,N_13738);
nor U14291 (N_14291,N_13920,N_13849);
and U14292 (N_14292,N_13772,N_13886);
and U14293 (N_14293,N_13677,N_13886);
nand U14294 (N_14294,N_13822,N_13612);
or U14295 (N_14295,N_13507,N_13919);
xnor U14296 (N_14296,N_13578,N_13638);
nor U14297 (N_14297,N_13635,N_13663);
or U14298 (N_14298,N_13740,N_13731);
nor U14299 (N_14299,N_13689,N_13628);
and U14300 (N_14300,N_13547,N_13515);
or U14301 (N_14301,N_13937,N_13555);
nor U14302 (N_14302,N_13818,N_13628);
and U14303 (N_14303,N_13523,N_13518);
nor U14304 (N_14304,N_13543,N_13994);
nor U14305 (N_14305,N_13867,N_13682);
nand U14306 (N_14306,N_13949,N_13506);
nand U14307 (N_14307,N_13655,N_13988);
nand U14308 (N_14308,N_13513,N_13571);
and U14309 (N_14309,N_13881,N_13795);
and U14310 (N_14310,N_13893,N_13756);
xor U14311 (N_14311,N_13887,N_13693);
nor U14312 (N_14312,N_13846,N_13568);
nand U14313 (N_14313,N_13832,N_13769);
and U14314 (N_14314,N_13770,N_13754);
nand U14315 (N_14315,N_13720,N_13761);
and U14316 (N_14316,N_13588,N_13660);
xor U14317 (N_14317,N_13886,N_13592);
and U14318 (N_14318,N_13863,N_13553);
nand U14319 (N_14319,N_13750,N_13700);
nand U14320 (N_14320,N_13780,N_13910);
xor U14321 (N_14321,N_13989,N_13522);
nor U14322 (N_14322,N_13965,N_13941);
or U14323 (N_14323,N_13892,N_13672);
and U14324 (N_14324,N_13790,N_13855);
nor U14325 (N_14325,N_13715,N_13843);
or U14326 (N_14326,N_13919,N_13636);
nor U14327 (N_14327,N_13684,N_13871);
and U14328 (N_14328,N_13934,N_13878);
or U14329 (N_14329,N_13928,N_13680);
xor U14330 (N_14330,N_13975,N_13919);
nor U14331 (N_14331,N_13779,N_13587);
or U14332 (N_14332,N_13938,N_13895);
xor U14333 (N_14333,N_13881,N_13843);
xor U14334 (N_14334,N_13749,N_13912);
nand U14335 (N_14335,N_13977,N_13695);
xor U14336 (N_14336,N_13849,N_13927);
xor U14337 (N_14337,N_13848,N_13651);
nor U14338 (N_14338,N_13913,N_13817);
nor U14339 (N_14339,N_13748,N_13640);
nand U14340 (N_14340,N_13863,N_13512);
nand U14341 (N_14341,N_13643,N_13557);
xnor U14342 (N_14342,N_13855,N_13768);
and U14343 (N_14343,N_13967,N_13863);
nand U14344 (N_14344,N_13515,N_13821);
nand U14345 (N_14345,N_13799,N_13646);
xor U14346 (N_14346,N_13566,N_13972);
or U14347 (N_14347,N_13513,N_13706);
or U14348 (N_14348,N_13655,N_13651);
and U14349 (N_14349,N_13911,N_13893);
and U14350 (N_14350,N_13783,N_13587);
nor U14351 (N_14351,N_13671,N_13801);
nand U14352 (N_14352,N_13631,N_13968);
xnor U14353 (N_14353,N_13985,N_13901);
xor U14354 (N_14354,N_13721,N_13835);
or U14355 (N_14355,N_13856,N_13754);
nand U14356 (N_14356,N_13541,N_13956);
or U14357 (N_14357,N_13818,N_13763);
nor U14358 (N_14358,N_13638,N_13640);
and U14359 (N_14359,N_13728,N_13518);
xnor U14360 (N_14360,N_13960,N_13644);
nand U14361 (N_14361,N_13597,N_13892);
and U14362 (N_14362,N_13630,N_13837);
nor U14363 (N_14363,N_13537,N_13786);
xnor U14364 (N_14364,N_13916,N_13633);
nor U14365 (N_14365,N_13514,N_13615);
nor U14366 (N_14366,N_13709,N_13566);
nand U14367 (N_14367,N_13697,N_13529);
and U14368 (N_14368,N_13826,N_13928);
xor U14369 (N_14369,N_13657,N_13707);
nand U14370 (N_14370,N_13582,N_13624);
or U14371 (N_14371,N_13511,N_13533);
and U14372 (N_14372,N_13930,N_13714);
nand U14373 (N_14373,N_13549,N_13539);
and U14374 (N_14374,N_13976,N_13870);
xor U14375 (N_14375,N_13596,N_13708);
nor U14376 (N_14376,N_13793,N_13657);
and U14377 (N_14377,N_13535,N_13998);
xnor U14378 (N_14378,N_13739,N_13850);
and U14379 (N_14379,N_13526,N_13592);
and U14380 (N_14380,N_13533,N_13629);
or U14381 (N_14381,N_13619,N_13938);
nor U14382 (N_14382,N_13813,N_13666);
nor U14383 (N_14383,N_13880,N_13511);
and U14384 (N_14384,N_13569,N_13647);
nand U14385 (N_14385,N_13799,N_13966);
nor U14386 (N_14386,N_13506,N_13881);
and U14387 (N_14387,N_13747,N_13963);
and U14388 (N_14388,N_13655,N_13739);
and U14389 (N_14389,N_13903,N_13594);
and U14390 (N_14390,N_13783,N_13991);
nand U14391 (N_14391,N_13867,N_13841);
nand U14392 (N_14392,N_13683,N_13786);
nand U14393 (N_14393,N_13583,N_13652);
and U14394 (N_14394,N_13539,N_13779);
xnor U14395 (N_14395,N_13829,N_13999);
nor U14396 (N_14396,N_13704,N_13607);
and U14397 (N_14397,N_13975,N_13549);
or U14398 (N_14398,N_13962,N_13510);
and U14399 (N_14399,N_13866,N_13720);
nand U14400 (N_14400,N_13772,N_13850);
and U14401 (N_14401,N_13943,N_13746);
xnor U14402 (N_14402,N_13634,N_13894);
or U14403 (N_14403,N_13952,N_13616);
nand U14404 (N_14404,N_13892,N_13819);
nand U14405 (N_14405,N_13801,N_13698);
nand U14406 (N_14406,N_13516,N_13561);
and U14407 (N_14407,N_13804,N_13869);
nor U14408 (N_14408,N_13974,N_13823);
nor U14409 (N_14409,N_13661,N_13787);
and U14410 (N_14410,N_13809,N_13541);
or U14411 (N_14411,N_13866,N_13990);
xor U14412 (N_14412,N_13762,N_13843);
xnor U14413 (N_14413,N_13775,N_13851);
or U14414 (N_14414,N_13606,N_13699);
nor U14415 (N_14415,N_13625,N_13667);
nand U14416 (N_14416,N_13704,N_13726);
nor U14417 (N_14417,N_13770,N_13557);
nor U14418 (N_14418,N_13966,N_13767);
or U14419 (N_14419,N_13873,N_13693);
nor U14420 (N_14420,N_13835,N_13512);
nor U14421 (N_14421,N_13743,N_13762);
xnor U14422 (N_14422,N_13792,N_13566);
xnor U14423 (N_14423,N_13598,N_13720);
nor U14424 (N_14424,N_13649,N_13900);
xor U14425 (N_14425,N_13563,N_13582);
xnor U14426 (N_14426,N_13501,N_13741);
nand U14427 (N_14427,N_13616,N_13524);
nor U14428 (N_14428,N_13958,N_13657);
xnor U14429 (N_14429,N_13725,N_13907);
or U14430 (N_14430,N_13911,N_13588);
xnor U14431 (N_14431,N_13782,N_13678);
nand U14432 (N_14432,N_13584,N_13616);
nor U14433 (N_14433,N_13889,N_13825);
xor U14434 (N_14434,N_13670,N_13837);
or U14435 (N_14435,N_13519,N_13765);
or U14436 (N_14436,N_13824,N_13656);
nor U14437 (N_14437,N_13703,N_13665);
nor U14438 (N_14438,N_13614,N_13977);
and U14439 (N_14439,N_13621,N_13881);
and U14440 (N_14440,N_13961,N_13955);
xor U14441 (N_14441,N_13860,N_13802);
nor U14442 (N_14442,N_13910,N_13977);
nand U14443 (N_14443,N_13890,N_13948);
and U14444 (N_14444,N_13976,N_13993);
nor U14445 (N_14445,N_13525,N_13758);
nor U14446 (N_14446,N_13986,N_13935);
nor U14447 (N_14447,N_13900,N_13865);
nor U14448 (N_14448,N_13824,N_13698);
nand U14449 (N_14449,N_13577,N_13544);
and U14450 (N_14450,N_13567,N_13921);
or U14451 (N_14451,N_13745,N_13610);
nor U14452 (N_14452,N_13700,N_13618);
and U14453 (N_14453,N_13609,N_13957);
xnor U14454 (N_14454,N_13528,N_13744);
nor U14455 (N_14455,N_13849,N_13815);
nor U14456 (N_14456,N_13714,N_13916);
nor U14457 (N_14457,N_13979,N_13713);
nor U14458 (N_14458,N_13777,N_13852);
nor U14459 (N_14459,N_13869,N_13993);
nand U14460 (N_14460,N_13825,N_13947);
and U14461 (N_14461,N_13669,N_13944);
nand U14462 (N_14462,N_13644,N_13817);
or U14463 (N_14463,N_13815,N_13501);
and U14464 (N_14464,N_13715,N_13747);
or U14465 (N_14465,N_13769,N_13655);
nand U14466 (N_14466,N_13842,N_13533);
xor U14467 (N_14467,N_13840,N_13510);
and U14468 (N_14468,N_13724,N_13840);
nand U14469 (N_14469,N_13576,N_13743);
nor U14470 (N_14470,N_13565,N_13882);
and U14471 (N_14471,N_13700,N_13927);
nor U14472 (N_14472,N_13936,N_13588);
xnor U14473 (N_14473,N_13867,N_13665);
xor U14474 (N_14474,N_13625,N_13763);
nand U14475 (N_14475,N_13826,N_13944);
nor U14476 (N_14476,N_13769,N_13585);
or U14477 (N_14477,N_13988,N_13781);
xor U14478 (N_14478,N_13660,N_13985);
xor U14479 (N_14479,N_13659,N_13791);
and U14480 (N_14480,N_13534,N_13521);
nor U14481 (N_14481,N_13808,N_13662);
nor U14482 (N_14482,N_13865,N_13776);
xor U14483 (N_14483,N_13530,N_13568);
or U14484 (N_14484,N_13614,N_13656);
nand U14485 (N_14485,N_13996,N_13846);
or U14486 (N_14486,N_13838,N_13812);
xor U14487 (N_14487,N_13536,N_13930);
or U14488 (N_14488,N_13974,N_13998);
nor U14489 (N_14489,N_13701,N_13885);
nor U14490 (N_14490,N_13628,N_13756);
xor U14491 (N_14491,N_13666,N_13728);
nor U14492 (N_14492,N_13531,N_13854);
nand U14493 (N_14493,N_13707,N_13750);
nand U14494 (N_14494,N_13504,N_13923);
or U14495 (N_14495,N_13806,N_13561);
and U14496 (N_14496,N_13943,N_13600);
and U14497 (N_14497,N_13869,N_13582);
nand U14498 (N_14498,N_13701,N_13696);
nor U14499 (N_14499,N_13519,N_13626);
nor U14500 (N_14500,N_14129,N_14148);
and U14501 (N_14501,N_14239,N_14086);
xor U14502 (N_14502,N_14370,N_14394);
nor U14503 (N_14503,N_14065,N_14125);
xnor U14504 (N_14504,N_14448,N_14126);
or U14505 (N_14505,N_14099,N_14090);
and U14506 (N_14506,N_14103,N_14180);
xnor U14507 (N_14507,N_14313,N_14211);
nand U14508 (N_14508,N_14135,N_14317);
xnor U14509 (N_14509,N_14410,N_14253);
or U14510 (N_14510,N_14344,N_14234);
xnor U14511 (N_14511,N_14462,N_14481);
xnor U14512 (N_14512,N_14142,N_14031);
or U14513 (N_14513,N_14266,N_14063);
nor U14514 (N_14514,N_14433,N_14392);
nor U14515 (N_14515,N_14096,N_14223);
nand U14516 (N_14516,N_14451,N_14300);
nor U14517 (N_14517,N_14443,N_14101);
xnor U14518 (N_14518,N_14442,N_14175);
nand U14519 (N_14519,N_14262,N_14062);
xor U14520 (N_14520,N_14081,N_14035);
xor U14521 (N_14521,N_14112,N_14469);
nand U14522 (N_14522,N_14042,N_14116);
and U14523 (N_14523,N_14309,N_14140);
xor U14524 (N_14524,N_14236,N_14267);
or U14525 (N_14525,N_14075,N_14215);
or U14526 (N_14526,N_14359,N_14438);
or U14527 (N_14527,N_14078,N_14431);
or U14528 (N_14528,N_14289,N_14486);
and U14529 (N_14529,N_14018,N_14165);
xor U14530 (N_14530,N_14196,N_14318);
xnor U14531 (N_14531,N_14014,N_14154);
and U14532 (N_14532,N_14004,N_14480);
nor U14533 (N_14533,N_14237,N_14200);
xor U14534 (N_14534,N_14232,N_14415);
nor U14535 (N_14535,N_14437,N_14388);
or U14536 (N_14536,N_14386,N_14320);
and U14537 (N_14537,N_14263,N_14383);
and U14538 (N_14538,N_14221,N_14464);
nand U14539 (N_14539,N_14463,N_14212);
xor U14540 (N_14540,N_14285,N_14074);
nand U14541 (N_14541,N_14173,N_14294);
nand U14542 (N_14542,N_14270,N_14174);
xor U14543 (N_14543,N_14029,N_14070);
and U14544 (N_14544,N_14187,N_14498);
or U14545 (N_14545,N_14179,N_14241);
or U14546 (N_14546,N_14189,N_14322);
xnor U14547 (N_14547,N_14380,N_14046);
nor U14548 (N_14548,N_14355,N_14152);
xnor U14549 (N_14549,N_14155,N_14444);
xnor U14550 (N_14550,N_14115,N_14254);
xor U14551 (N_14551,N_14319,N_14087);
or U14552 (N_14552,N_14199,N_14238);
or U14553 (N_14553,N_14349,N_14177);
nand U14554 (N_14554,N_14325,N_14250);
or U14555 (N_14555,N_14417,N_14166);
or U14556 (N_14556,N_14231,N_14176);
or U14557 (N_14557,N_14290,N_14001);
xor U14558 (N_14558,N_14378,N_14160);
nand U14559 (N_14559,N_14235,N_14037);
or U14560 (N_14560,N_14472,N_14182);
xor U14561 (N_14561,N_14039,N_14033);
nor U14562 (N_14562,N_14424,N_14406);
nor U14563 (N_14563,N_14495,N_14242);
nor U14564 (N_14564,N_14120,N_14222);
nand U14565 (N_14565,N_14207,N_14399);
and U14566 (N_14566,N_14002,N_14402);
xnor U14567 (N_14567,N_14150,N_14181);
nor U14568 (N_14568,N_14168,N_14186);
nand U14569 (N_14569,N_14038,N_14157);
nand U14570 (N_14570,N_14192,N_14401);
nor U14571 (N_14571,N_14418,N_14027);
nor U14572 (N_14572,N_14413,N_14365);
xor U14573 (N_14573,N_14416,N_14047);
and U14574 (N_14574,N_14275,N_14356);
nor U14575 (N_14575,N_14283,N_14434);
or U14576 (N_14576,N_14217,N_14379);
nor U14577 (N_14577,N_14229,N_14023);
nor U14578 (N_14578,N_14298,N_14385);
nand U14579 (N_14579,N_14350,N_14430);
and U14580 (N_14580,N_14393,N_14473);
nor U14581 (N_14581,N_14206,N_14408);
or U14582 (N_14582,N_14375,N_14137);
nor U14583 (N_14583,N_14389,N_14381);
nor U14584 (N_14584,N_14366,N_14012);
and U14585 (N_14585,N_14219,N_14195);
nand U14586 (N_14586,N_14303,N_14308);
and U14587 (N_14587,N_14427,N_14147);
nor U14588 (N_14588,N_14045,N_14151);
nand U14589 (N_14589,N_14017,N_14387);
xnor U14590 (N_14590,N_14497,N_14460);
and U14591 (N_14591,N_14056,N_14414);
xnor U14592 (N_14592,N_14162,N_14185);
or U14593 (N_14593,N_14257,N_14288);
or U14594 (N_14594,N_14404,N_14139);
or U14595 (N_14595,N_14272,N_14423);
or U14596 (N_14596,N_14227,N_14209);
nor U14597 (N_14597,N_14026,N_14407);
nor U14598 (N_14598,N_14145,N_14247);
and U14599 (N_14599,N_14055,N_14293);
nand U14600 (N_14600,N_14198,N_14025);
nand U14601 (N_14601,N_14493,N_14226);
xor U14602 (N_14602,N_14178,N_14419);
or U14603 (N_14603,N_14061,N_14456);
or U14604 (N_14604,N_14021,N_14422);
or U14605 (N_14605,N_14453,N_14119);
and U14606 (N_14606,N_14452,N_14287);
xor U14607 (N_14607,N_14088,N_14102);
nand U14608 (N_14608,N_14377,N_14138);
nor U14609 (N_14609,N_14032,N_14073);
or U14610 (N_14610,N_14468,N_14396);
and U14611 (N_14611,N_14008,N_14341);
nor U14612 (N_14612,N_14307,N_14425);
or U14613 (N_14613,N_14244,N_14020);
and U14614 (N_14614,N_14302,N_14123);
and U14615 (N_14615,N_14084,N_14091);
nor U14616 (N_14616,N_14041,N_14278);
or U14617 (N_14617,N_14197,N_14083);
or U14618 (N_14618,N_14048,N_14144);
or U14619 (N_14619,N_14076,N_14305);
and U14620 (N_14620,N_14265,N_14492);
nand U14621 (N_14621,N_14457,N_14213);
or U14622 (N_14622,N_14465,N_14240);
and U14623 (N_14623,N_14286,N_14216);
nor U14624 (N_14624,N_14301,N_14328);
nand U14625 (N_14625,N_14333,N_14225);
or U14626 (N_14626,N_14490,N_14246);
and U14627 (N_14627,N_14011,N_14329);
and U14628 (N_14628,N_14339,N_14024);
or U14629 (N_14629,N_14342,N_14489);
and U14630 (N_14630,N_14436,N_14447);
nand U14631 (N_14631,N_14391,N_14057);
nand U14632 (N_14632,N_14113,N_14013);
nand U14633 (N_14633,N_14255,N_14141);
nand U14634 (N_14634,N_14233,N_14044);
nand U14635 (N_14635,N_14475,N_14440);
nor U14636 (N_14636,N_14243,N_14069);
or U14637 (N_14637,N_14282,N_14450);
nand U14638 (N_14638,N_14337,N_14170);
xor U14639 (N_14639,N_14327,N_14276);
or U14640 (N_14640,N_14454,N_14347);
xnor U14641 (N_14641,N_14260,N_14340);
nand U14642 (N_14642,N_14172,N_14161);
xor U14643 (N_14643,N_14346,N_14252);
and U14644 (N_14644,N_14127,N_14398);
xnor U14645 (N_14645,N_14251,N_14296);
or U14646 (N_14646,N_14368,N_14336);
xnor U14647 (N_14647,N_14249,N_14171);
xor U14648 (N_14648,N_14095,N_14133);
or U14649 (N_14649,N_14034,N_14000);
nor U14650 (N_14650,N_14132,N_14374);
and U14651 (N_14651,N_14203,N_14299);
nand U14652 (N_14652,N_14040,N_14268);
xnor U14653 (N_14653,N_14482,N_14077);
and U14654 (N_14654,N_14036,N_14367);
xor U14655 (N_14655,N_14357,N_14376);
nand U14656 (N_14656,N_14403,N_14130);
or U14657 (N_14657,N_14228,N_14369);
or U14658 (N_14658,N_14390,N_14284);
nor U14659 (N_14659,N_14353,N_14466);
or U14660 (N_14660,N_14100,N_14358);
xnor U14661 (N_14661,N_14131,N_14261);
and U14662 (N_14662,N_14054,N_14459);
and U14663 (N_14663,N_14190,N_14109);
or U14664 (N_14664,N_14167,N_14446);
nor U14665 (N_14665,N_14354,N_14068);
and U14666 (N_14666,N_14019,N_14499);
nor U14667 (N_14667,N_14277,N_14258);
xnor U14668 (N_14668,N_14106,N_14271);
nor U14669 (N_14669,N_14264,N_14193);
and U14670 (N_14670,N_14467,N_14124);
nor U14671 (N_14671,N_14146,N_14121);
xor U14672 (N_14672,N_14134,N_14089);
nor U14673 (N_14673,N_14051,N_14210);
xor U14674 (N_14674,N_14052,N_14316);
nor U14675 (N_14675,N_14050,N_14028);
or U14676 (N_14676,N_14435,N_14111);
and U14677 (N_14677,N_14487,N_14094);
xnor U14678 (N_14678,N_14085,N_14332);
nand U14679 (N_14679,N_14364,N_14312);
and U14680 (N_14680,N_14156,N_14164);
xnor U14681 (N_14681,N_14071,N_14292);
nand U14682 (N_14682,N_14483,N_14194);
or U14683 (N_14683,N_14478,N_14330);
or U14684 (N_14684,N_14420,N_14280);
and U14685 (N_14685,N_14371,N_14471);
xor U14686 (N_14686,N_14494,N_14479);
or U14687 (N_14687,N_14248,N_14496);
and U14688 (N_14688,N_14455,N_14345);
or U14689 (N_14689,N_14022,N_14159);
or U14690 (N_14690,N_14143,N_14449);
nand U14691 (N_14691,N_14006,N_14400);
xor U14692 (N_14692,N_14432,N_14397);
and U14693 (N_14693,N_14058,N_14184);
and U14694 (N_14694,N_14352,N_14461);
or U14695 (N_14695,N_14291,N_14007);
nand U14696 (N_14696,N_14439,N_14049);
nand U14697 (N_14697,N_14441,N_14043);
nor U14698 (N_14698,N_14477,N_14351);
nand U14699 (N_14699,N_14191,N_14384);
and U14700 (N_14700,N_14362,N_14323);
nor U14701 (N_14701,N_14488,N_14183);
nor U14702 (N_14702,N_14421,N_14343);
and U14703 (N_14703,N_14411,N_14079);
xor U14704 (N_14704,N_14279,N_14335);
xor U14705 (N_14705,N_14016,N_14220);
or U14706 (N_14706,N_14169,N_14098);
or U14707 (N_14707,N_14338,N_14348);
xor U14708 (N_14708,N_14128,N_14395);
xor U14709 (N_14709,N_14218,N_14458);
and U14710 (N_14710,N_14314,N_14256);
and U14711 (N_14711,N_14163,N_14015);
and U14712 (N_14712,N_14136,N_14245);
nand U14713 (N_14713,N_14110,N_14188);
nand U14714 (N_14714,N_14093,N_14426);
and U14715 (N_14715,N_14202,N_14067);
nor U14716 (N_14716,N_14274,N_14310);
nand U14717 (N_14717,N_14297,N_14412);
or U14718 (N_14718,N_14114,N_14484);
nor U14719 (N_14719,N_14470,N_14010);
or U14720 (N_14720,N_14108,N_14273);
and U14721 (N_14721,N_14360,N_14214);
and U14722 (N_14722,N_14072,N_14104);
nor U14723 (N_14723,N_14372,N_14429);
xnor U14724 (N_14724,N_14122,N_14476);
and U14725 (N_14725,N_14009,N_14409);
or U14726 (N_14726,N_14334,N_14311);
nor U14727 (N_14727,N_14053,N_14059);
xor U14728 (N_14728,N_14201,N_14281);
xnor U14729 (N_14729,N_14030,N_14080);
and U14730 (N_14730,N_14158,N_14097);
and U14731 (N_14731,N_14208,N_14205);
and U14732 (N_14732,N_14149,N_14117);
or U14733 (N_14733,N_14321,N_14230);
and U14734 (N_14734,N_14005,N_14361);
or U14735 (N_14735,N_14092,N_14306);
xor U14736 (N_14736,N_14382,N_14204);
or U14737 (N_14737,N_14373,N_14224);
or U14738 (N_14738,N_14153,N_14295);
nor U14739 (N_14739,N_14445,N_14485);
nand U14740 (N_14740,N_14304,N_14474);
xor U14741 (N_14741,N_14269,N_14105);
nor U14742 (N_14742,N_14066,N_14118);
or U14743 (N_14743,N_14326,N_14315);
nand U14744 (N_14744,N_14491,N_14003);
nand U14745 (N_14745,N_14064,N_14060);
nand U14746 (N_14746,N_14107,N_14324);
xnor U14747 (N_14747,N_14331,N_14363);
nor U14748 (N_14748,N_14259,N_14405);
nor U14749 (N_14749,N_14428,N_14082);
nor U14750 (N_14750,N_14199,N_14339);
xnor U14751 (N_14751,N_14029,N_14352);
xor U14752 (N_14752,N_14224,N_14276);
xor U14753 (N_14753,N_14115,N_14195);
nor U14754 (N_14754,N_14298,N_14215);
or U14755 (N_14755,N_14203,N_14389);
and U14756 (N_14756,N_14186,N_14089);
nand U14757 (N_14757,N_14194,N_14095);
and U14758 (N_14758,N_14465,N_14316);
nor U14759 (N_14759,N_14312,N_14217);
and U14760 (N_14760,N_14440,N_14178);
nor U14761 (N_14761,N_14397,N_14045);
nor U14762 (N_14762,N_14495,N_14271);
or U14763 (N_14763,N_14097,N_14024);
and U14764 (N_14764,N_14159,N_14125);
and U14765 (N_14765,N_14343,N_14388);
and U14766 (N_14766,N_14304,N_14076);
xnor U14767 (N_14767,N_14433,N_14445);
nand U14768 (N_14768,N_14458,N_14167);
or U14769 (N_14769,N_14378,N_14105);
and U14770 (N_14770,N_14445,N_14390);
nor U14771 (N_14771,N_14349,N_14260);
and U14772 (N_14772,N_14177,N_14089);
or U14773 (N_14773,N_14089,N_14189);
nor U14774 (N_14774,N_14319,N_14137);
nand U14775 (N_14775,N_14307,N_14123);
xor U14776 (N_14776,N_14069,N_14221);
nor U14777 (N_14777,N_14072,N_14416);
nor U14778 (N_14778,N_14302,N_14019);
xnor U14779 (N_14779,N_14463,N_14211);
nor U14780 (N_14780,N_14250,N_14398);
nor U14781 (N_14781,N_14475,N_14109);
nor U14782 (N_14782,N_14171,N_14192);
xnor U14783 (N_14783,N_14106,N_14047);
nor U14784 (N_14784,N_14078,N_14223);
and U14785 (N_14785,N_14263,N_14378);
and U14786 (N_14786,N_14148,N_14336);
and U14787 (N_14787,N_14447,N_14438);
xnor U14788 (N_14788,N_14440,N_14136);
or U14789 (N_14789,N_14264,N_14459);
or U14790 (N_14790,N_14341,N_14243);
and U14791 (N_14791,N_14242,N_14116);
and U14792 (N_14792,N_14091,N_14499);
nand U14793 (N_14793,N_14370,N_14184);
nand U14794 (N_14794,N_14310,N_14476);
nand U14795 (N_14795,N_14499,N_14227);
nand U14796 (N_14796,N_14306,N_14444);
and U14797 (N_14797,N_14099,N_14140);
and U14798 (N_14798,N_14041,N_14449);
nor U14799 (N_14799,N_14190,N_14421);
and U14800 (N_14800,N_14467,N_14367);
xnor U14801 (N_14801,N_14042,N_14433);
nor U14802 (N_14802,N_14450,N_14401);
xor U14803 (N_14803,N_14494,N_14069);
or U14804 (N_14804,N_14034,N_14411);
xnor U14805 (N_14805,N_14454,N_14149);
xnor U14806 (N_14806,N_14312,N_14435);
and U14807 (N_14807,N_14130,N_14262);
or U14808 (N_14808,N_14389,N_14418);
nand U14809 (N_14809,N_14157,N_14119);
nand U14810 (N_14810,N_14232,N_14487);
xnor U14811 (N_14811,N_14089,N_14398);
nand U14812 (N_14812,N_14212,N_14021);
and U14813 (N_14813,N_14271,N_14124);
and U14814 (N_14814,N_14299,N_14102);
or U14815 (N_14815,N_14089,N_14196);
nand U14816 (N_14816,N_14176,N_14364);
nand U14817 (N_14817,N_14012,N_14443);
or U14818 (N_14818,N_14054,N_14029);
nor U14819 (N_14819,N_14118,N_14491);
and U14820 (N_14820,N_14179,N_14362);
or U14821 (N_14821,N_14424,N_14065);
nor U14822 (N_14822,N_14180,N_14205);
nand U14823 (N_14823,N_14288,N_14181);
and U14824 (N_14824,N_14195,N_14448);
or U14825 (N_14825,N_14439,N_14176);
xor U14826 (N_14826,N_14478,N_14096);
nor U14827 (N_14827,N_14042,N_14299);
and U14828 (N_14828,N_14442,N_14145);
xnor U14829 (N_14829,N_14013,N_14123);
xnor U14830 (N_14830,N_14261,N_14055);
or U14831 (N_14831,N_14410,N_14183);
nor U14832 (N_14832,N_14474,N_14091);
or U14833 (N_14833,N_14471,N_14472);
xnor U14834 (N_14834,N_14363,N_14122);
nand U14835 (N_14835,N_14496,N_14017);
and U14836 (N_14836,N_14188,N_14286);
or U14837 (N_14837,N_14296,N_14138);
or U14838 (N_14838,N_14083,N_14142);
nor U14839 (N_14839,N_14373,N_14258);
or U14840 (N_14840,N_14131,N_14356);
and U14841 (N_14841,N_14391,N_14095);
nor U14842 (N_14842,N_14440,N_14100);
and U14843 (N_14843,N_14493,N_14092);
and U14844 (N_14844,N_14127,N_14154);
and U14845 (N_14845,N_14113,N_14293);
xnor U14846 (N_14846,N_14355,N_14197);
nor U14847 (N_14847,N_14246,N_14320);
xor U14848 (N_14848,N_14131,N_14461);
nand U14849 (N_14849,N_14493,N_14309);
nor U14850 (N_14850,N_14477,N_14427);
nand U14851 (N_14851,N_14039,N_14402);
nor U14852 (N_14852,N_14224,N_14364);
nand U14853 (N_14853,N_14498,N_14472);
xnor U14854 (N_14854,N_14041,N_14400);
or U14855 (N_14855,N_14196,N_14364);
xnor U14856 (N_14856,N_14363,N_14111);
or U14857 (N_14857,N_14012,N_14218);
nand U14858 (N_14858,N_14329,N_14061);
nand U14859 (N_14859,N_14224,N_14086);
xnor U14860 (N_14860,N_14147,N_14093);
nor U14861 (N_14861,N_14033,N_14253);
or U14862 (N_14862,N_14271,N_14410);
xnor U14863 (N_14863,N_14032,N_14046);
nand U14864 (N_14864,N_14257,N_14248);
nand U14865 (N_14865,N_14322,N_14094);
xor U14866 (N_14866,N_14411,N_14027);
and U14867 (N_14867,N_14091,N_14367);
or U14868 (N_14868,N_14018,N_14186);
and U14869 (N_14869,N_14203,N_14168);
and U14870 (N_14870,N_14181,N_14127);
or U14871 (N_14871,N_14276,N_14331);
nand U14872 (N_14872,N_14295,N_14186);
nand U14873 (N_14873,N_14060,N_14083);
or U14874 (N_14874,N_14414,N_14130);
nor U14875 (N_14875,N_14340,N_14493);
xnor U14876 (N_14876,N_14211,N_14476);
xnor U14877 (N_14877,N_14347,N_14238);
or U14878 (N_14878,N_14342,N_14442);
and U14879 (N_14879,N_14473,N_14384);
or U14880 (N_14880,N_14394,N_14000);
nor U14881 (N_14881,N_14423,N_14016);
nor U14882 (N_14882,N_14184,N_14125);
nand U14883 (N_14883,N_14037,N_14287);
and U14884 (N_14884,N_14251,N_14199);
nor U14885 (N_14885,N_14260,N_14300);
nand U14886 (N_14886,N_14172,N_14271);
or U14887 (N_14887,N_14220,N_14062);
nand U14888 (N_14888,N_14499,N_14102);
and U14889 (N_14889,N_14393,N_14437);
nor U14890 (N_14890,N_14140,N_14069);
nand U14891 (N_14891,N_14181,N_14114);
nand U14892 (N_14892,N_14341,N_14348);
and U14893 (N_14893,N_14169,N_14146);
nor U14894 (N_14894,N_14400,N_14150);
nor U14895 (N_14895,N_14026,N_14067);
or U14896 (N_14896,N_14480,N_14199);
and U14897 (N_14897,N_14171,N_14048);
or U14898 (N_14898,N_14056,N_14267);
xor U14899 (N_14899,N_14344,N_14429);
nand U14900 (N_14900,N_14210,N_14377);
and U14901 (N_14901,N_14021,N_14490);
and U14902 (N_14902,N_14353,N_14383);
nand U14903 (N_14903,N_14484,N_14401);
xnor U14904 (N_14904,N_14477,N_14116);
xnor U14905 (N_14905,N_14053,N_14450);
nand U14906 (N_14906,N_14377,N_14419);
xnor U14907 (N_14907,N_14450,N_14272);
nor U14908 (N_14908,N_14455,N_14229);
and U14909 (N_14909,N_14460,N_14033);
nor U14910 (N_14910,N_14203,N_14154);
nand U14911 (N_14911,N_14380,N_14323);
xnor U14912 (N_14912,N_14157,N_14252);
or U14913 (N_14913,N_14471,N_14450);
nor U14914 (N_14914,N_14188,N_14033);
and U14915 (N_14915,N_14401,N_14448);
nand U14916 (N_14916,N_14077,N_14299);
xnor U14917 (N_14917,N_14444,N_14473);
xnor U14918 (N_14918,N_14097,N_14435);
nand U14919 (N_14919,N_14357,N_14368);
nor U14920 (N_14920,N_14057,N_14353);
xor U14921 (N_14921,N_14373,N_14461);
nor U14922 (N_14922,N_14329,N_14392);
xor U14923 (N_14923,N_14250,N_14447);
and U14924 (N_14924,N_14156,N_14465);
and U14925 (N_14925,N_14374,N_14146);
nand U14926 (N_14926,N_14190,N_14084);
nor U14927 (N_14927,N_14174,N_14398);
nand U14928 (N_14928,N_14118,N_14306);
or U14929 (N_14929,N_14271,N_14076);
nor U14930 (N_14930,N_14322,N_14421);
and U14931 (N_14931,N_14143,N_14248);
xor U14932 (N_14932,N_14053,N_14362);
nor U14933 (N_14933,N_14282,N_14211);
nor U14934 (N_14934,N_14279,N_14211);
xnor U14935 (N_14935,N_14461,N_14244);
or U14936 (N_14936,N_14466,N_14016);
and U14937 (N_14937,N_14469,N_14403);
nor U14938 (N_14938,N_14421,N_14440);
nor U14939 (N_14939,N_14019,N_14136);
xor U14940 (N_14940,N_14035,N_14115);
nand U14941 (N_14941,N_14062,N_14392);
nor U14942 (N_14942,N_14412,N_14428);
nor U14943 (N_14943,N_14183,N_14217);
or U14944 (N_14944,N_14253,N_14291);
nand U14945 (N_14945,N_14034,N_14183);
and U14946 (N_14946,N_14468,N_14392);
and U14947 (N_14947,N_14244,N_14456);
nor U14948 (N_14948,N_14048,N_14186);
or U14949 (N_14949,N_14119,N_14286);
and U14950 (N_14950,N_14407,N_14121);
or U14951 (N_14951,N_14195,N_14192);
and U14952 (N_14952,N_14349,N_14407);
nand U14953 (N_14953,N_14121,N_14355);
and U14954 (N_14954,N_14251,N_14222);
nand U14955 (N_14955,N_14000,N_14397);
and U14956 (N_14956,N_14326,N_14122);
or U14957 (N_14957,N_14024,N_14273);
and U14958 (N_14958,N_14273,N_14132);
nor U14959 (N_14959,N_14082,N_14323);
nand U14960 (N_14960,N_14317,N_14319);
nand U14961 (N_14961,N_14386,N_14223);
nand U14962 (N_14962,N_14243,N_14296);
and U14963 (N_14963,N_14473,N_14260);
xnor U14964 (N_14964,N_14443,N_14132);
or U14965 (N_14965,N_14163,N_14162);
nor U14966 (N_14966,N_14138,N_14431);
or U14967 (N_14967,N_14408,N_14416);
or U14968 (N_14968,N_14189,N_14466);
and U14969 (N_14969,N_14234,N_14115);
or U14970 (N_14970,N_14349,N_14176);
nor U14971 (N_14971,N_14238,N_14325);
xor U14972 (N_14972,N_14401,N_14466);
or U14973 (N_14973,N_14307,N_14099);
xor U14974 (N_14974,N_14457,N_14438);
nand U14975 (N_14975,N_14086,N_14316);
nor U14976 (N_14976,N_14133,N_14123);
nor U14977 (N_14977,N_14497,N_14495);
nand U14978 (N_14978,N_14180,N_14408);
xnor U14979 (N_14979,N_14148,N_14408);
xnor U14980 (N_14980,N_14298,N_14338);
nand U14981 (N_14981,N_14319,N_14219);
and U14982 (N_14982,N_14162,N_14223);
nor U14983 (N_14983,N_14186,N_14143);
and U14984 (N_14984,N_14242,N_14186);
or U14985 (N_14985,N_14296,N_14335);
nand U14986 (N_14986,N_14388,N_14483);
and U14987 (N_14987,N_14315,N_14358);
nand U14988 (N_14988,N_14140,N_14333);
xor U14989 (N_14989,N_14266,N_14274);
nor U14990 (N_14990,N_14459,N_14006);
nor U14991 (N_14991,N_14035,N_14284);
or U14992 (N_14992,N_14397,N_14192);
nor U14993 (N_14993,N_14278,N_14418);
nor U14994 (N_14994,N_14413,N_14077);
or U14995 (N_14995,N_14147,N_14319);
or U14996 (N_14996,N_14365,N_14380);
xnor U14997 (N_14997,N_14081,N_14125);
and U14998 (N_14998,N_14029,N_14447);
or U14999 (N_14999,N_14278,N_14256);
and U15000 (N_15000,N_14665,N_14685);
or U15001 (N_15001,N_14963,N_14738);
nand U15002 (N_15002,N_14777,N_14946);
and U15003 (N_15003,N_14784,N_14915);
or U15004 (N_15004,N_14558,N_14678);
or U15005 (N_15005,N_14856,N_14932);
or U15006 (N_15006,N_14864,N_14965);
or U15007 (N_15007,N_14889,N_14773);
nand U15008 (N_15008,N_14703,N_14522);
xor U15009 (N_15009,N_14511,N_14680);
and U15010 (N_15010,N_14766,N_14536);
xnor U15011 (N_15011,N_14663,N_14636);
nor U15012 (N_15012,N_14579,N_14865);
or U15013 (N_15013,N_14585,N_14602);
xor U15014 (N_15014,N_14978,N_14944);
nor U15015 (N_15015,N_14521,N_14826);
and U15016 (N_15016,N_14917,N_14986);
nand U15017 (N_15017,N_14785,N_14653);
nor U15018 (N_15018,N_14822,N_14976);
nor U15019 (N_15019,N_14689,N_14983);
nand U15020 (N_15020,N_14592,N_14625);
nand U15021 (N_15021,N_14537,N_14567);
and U15022 (N_15022,N_14517,N_14791);
xnor U15023 (N_15023,N_14989,N_14745);
or U15024 (N_15024,N_14500,N_14502);
nor U15025 (N_15025,N_14734,N_14699);
xnor U15026 (N_15026,N_14798,N_14572);
and U15027 (N_15027,N_14939,N_14775);
nand U15028 (N_15028,N_14818,N_14520);
xor U15029 (N_15029,N_14763,N_14878);
or U15030 (N_15030,N_14575,N_14611);
or U15031 (N_15031,N_14613,N_14778);
nor U15032 (N_15032,N_14913,N_14735);
xnor U15033 (N_15033,N_14759,N_14929);
and U15034 (N_15034,N_14597,N_14967);
xnor U15035 (N_15035,N_14987,N_14796);
nor U15036 (N_15036,N_14669,N_14909);
nor U15037 (N_15037,N_14615,N_14606);
nand U15038 (N_15038,N_14790,N_14740);
or U15039 (N_15039,N_14538,N_14524);
nor U15040 (N_15040,N_14860,N_14859);
nand U15041 (N_15041,N_14968,N_14523);
and U15042 (N_15042,N_14687,N_14568);
and U15043 (N_15043,N_14867,N_14662);
xnor U15044 (N_15044,N_14566,N_14846);
or U15045 (N_15045,N_14563,N_14507);
and U15046 (N_15046,N_14619,N_14649);
and U15047 (N_15047,N_14897,N_14719);
and U15048 (N_15048,N_14840,N_14970);
nand U15049 (N_15049,N_14623,N_14927);
nor U15050 (N_15050,N_14684,N_14600);
xor U15051 (N_15051,N_14694,N_14549);
xor U15052 (N_15052,N_14858,N_14701);
or U15053 (N_15053,N_14919,N_14633);
or U15054 (N_15054,N_14945,N_14670);
nand U15055 (N_15055,N_14804,N_14608);
or U15056 (N_15056,N_14937,N_14799);
nor U15057 (N_15057,N_14879,N_14589);
or U15058 (N_15058,N_14988,N_14783);
nand U15059 (N_15059,N_14863,N_14871);
or U15060 (N_15060,N_14727,N_14626);
xnor U15061 (N_15061,N_14949,N_14838);
xnor U15062 (N_15062,N_14995,N_14922);
and U15063 (N_15063,N_14887,N_14627);
nor U15064 (N_15064,N_14621,N_14547);
or U15065 (N_15065,N_14971,N_14555);
nand U15066 (N_15066,N_14749,N_14657);
and U15067 (N_15067,N_14692,N_14630);
and U15068 (N_15068,N_14902,N_14709);
nor U15069 (N_15069,N_14910,N_14730);
xnor U15070 (N_15070,N_14673,N_14705);
nor U15071 (N_15071,N_14837,N_14564);
nor U15072 (N_15072,N_14722,N_14924);
or U15073 (N_15073,N_14543,N_14721);
xor U15074 (N_15074,N_14542,N_14587);
nor U15075 (N_15075,N_14938,N_14647);
and U15076 (N_15076,N_14664,N_14565);
and U15077 (N_15077,N_14757,N_14557);
nand U15078 (N_15078,N_14618,N_14786);
and U15079 (N_15079,N_14569,N_14805);
and U15080 (N_15080,N_14855,N_14961);
nor U15081 (N_15081,N_14831,N_14894);
nor U15082 (N_15082,N_14788,N_14732);
and U15083 (N_15083,N_14953,N_14936);
xor U15084 (N_15084,N_14642,N_14849);
or U15085 (N_15085,N_14612,N_14883);
and U15086 (N_15086,N_14546,N_14548);
and U15087 (N_15087,N_14952,N_14659);
nand U15088 (N_15088,N_14872,N_14529);
or U15089 (N_15089,N_14545,N_14741);
and U15090 (N_15090,N_14898,N_14903);
and U15091 (N_15091,N_14803,N_14646);
xnor U15092 (N_15092,N_14886,N_14984);
or U15093 (N_15093,N_14590,N_14852);
xnor U15094 (N_15094,N_14601,N_14603);
nor U15095 (N_15095,N_14693,N_14880);
nor U15096 (N_15096,N_14885,N_14966);
nor U15097 (N_15097,N_14723,N_14700);
and U15098 (N_15098,N_14931,N_14651);
nand U15099 (N_15099,N_14764,N_14714);
and U15100 (N_15100,N_14586,N_14861);
and U15101 (N_15101,N_14881,N_14999);
nor U15102 (N_15102,N_14682,N_14720);
and U15103 (N_15103,N_14655,N_14577);
or U15104 (N_15104,N_14993,N_14594);
nand U15105 (N_15105,N_14675,N_14526);
xor U15106 (N_15106,N_14528,N_14997);
nor U15107 (N_15107,N_14743,N_14591);
xor U15108 (N_15108,N_14847,N_14827);
nand U15109 (N_15109,N_14906,N_14862);
nor U15110 (N_15110,N_14576,N_14789);
and U15111 (N_15111,N_14553,N_14809);
nand U15112 (N_15112,N_14581,N_14992);
and U15113 (N_15113,N_14930,N_14672);
and U15114 (N_15114,N_14504,N_14940);
xor U15115 (N_15115,N_14656,N_14750);
xor U15116 (N_15116,N_14697,N_14787);
nand U15117 (N_15117,N_14532,N_14969);
xor U15118 (N_15118,N_14641,N_14710);
nor U15119 (N_15119,N_14540,N_14754);
nor U15120 (N_15120,N_14920,N_14531);
xnor U15121 (N_15121,N_14715,N_14893);
or U15122 (N_15122,N_14718,N_14588);
and U15123 (N_15123,N_14560,N_14981);
and U15124 (N_15124,N_14679,N_14661);
or U15125 (N_15125,N_14728,N_14868);
nor U15126 (N_15126,N_14515,N_14503);
nand U15127 (N_15127,N_14559,N_14998);
nor U15128 (N_15128,N_14811,N_14781);
and U15129 (N_15129,N_14921,N_14774);
nor U15130 (N_15130,N_14658,N_14935);
nor U15131 (N_15131,N_14828,N_14683);
nor U15132 (N_15132,N_14794,N_14990);
xnor U15133 (N_15133,N_14731,N_14578);
nor U15134 (N_15134,N_14996,N_14807);
and U15135 (N_15135,N_14900,N_14599);
and U15136 (N_15136,N_14896,N_14985);
nor U15137 (N_15137,N_14533,N_14583);
nand U15138 (N_15138,N_14876,N_14795);
nand U15139 (N_15139,N_14844,N_14725);
nor U15140 (N_15140,N_14635,N_14891);
xnor U15141 (N_15141,N_14681,N_14851);
and U15142 (N_15142,N_14899,N_14857);
xor U15143 (N_15143,N_14737,N_14620);
nand U15144 (N_15144,N_14758,N_14869);
nand U15145 (N_15145,N_14595,N_14593);
or U15146 (N_15146,N_14711,N_14808);
and U15147 (N_15147,N_14810,N_14742);
nor U15148 (N_15148,N_14518,N_14570);
nor U15149 (N_15149,N_14823,N_14982);
nor U15150 (N_15150,N_14842,N_14875);
xnor U15151 (N_15151,N_14839,N_14760);
and U15152 (N_15152,N_14813,N_14519);
and U15153 (N_15153,N_14888,N_14960);
nand U15154 (N_15154,N_14845,N_14918);
xor U15155 (N_15155,N_14671,N_14505);
nand U15156 (N_15156,N_14956,N_14748);
nor U15157 (N_15157,N_14660,N_14776);
nand U15158 (N_15158,N_14510,N_14890);
nor U15159 (N_15159,N_14527,N_14561);
or U15160 (N_15160,N_14668,N_14525);
nand U15161 (N_15161,N_14770,N_14706);
xnor U15162 (N_15162,N_14884,N_14854);
or U15163 (N_15163,N_14580,N_14755);
or U15164 (N_15164,N_14958,N_14729);
or U15165 (N_15165,N_14556,N_14877);
nor U15166 (N_15166,N_14639,N_14991);
nand U15167 (N_15167,N_14512,N_14702);
and U15168 (N_15168,N_14582,N_14780);
and U15169 (N_15169,N_14690,N_14712);
or U15170 (N_15170,N_14610,N_14914);
xor U15171 (N_15171,N_14955,N_14691);
or U15172 (N_15172,N_14850,N_14779);
and U15173 (N_15173,N_14550,N_14977);
or U15174 (N_15174,N_14733,N_14501);
xor U15175 (N_15175,N_14761,N_14716);
nor U15176 (N_15176,N_14830,N_14832);
or U15177 (N_15177,N_14614,N_14950);
nor U15178 (N_15178,N_14629,N_14762);
nand U15179 (N_15179,N_14994,N_14513);
or U15180 (N_15180,N_14751,N_14747);
nand U15181 (N_15181,N_14972,N_14739);
xor U15182 (N_15182,N_14916,N_14874);
nand U15183 (N_15183,N_14695,N_14873);
and U15184 (N_15184,N_14640,N_14508);
nor U15185 (N_15185,N_14605,N_14870);
or U15186 (N_15186,N_14624,N_14704);
or U15187 (N_15187,N_14892,N_14833);
nand U15188 (N_15188,N_14923,N_14698);
nand U15189 (N_15189,N_14713,N_14571);
nand U15190 (N_15190,N_14836,N_14980);
nor U15191 (N_15191,N_14908,N_14825);
and U15192 (N_15192,N_14843,N_14882);
and U15193 (N_15193,N_14707,N_14814);
nand U15194 (N_15194,N_14933,N_14573);
nor U15195 (N_15195,N_14821,N_14973);
nor U15196 (N_15196,N_14650,N_14816);
nor U15197 (N_15197,N_14696,N_14752);
nand U15198 (N_15198,N_14631,N_14954);
or U15199 (N_15199,N_14767,N_14962);
and U15200 (N_15200,N_14552,N_14736);
or U15201 (N_15201,N_14901,N_14688);
and U15202 (N_15202,N_14841,N_14535);
xnor U15203 (N_15203,N_14911,N_14596);
nand U15204 (N_15204,N_14717,N_14514);
or U15205 (N_15205,N_14634,N_14637);
xnor U15206 (N_15206,N_14746,N_14598);
nor U15207 (N_15207,N_14644,N_14643);
or U15208 (N_15208,N_14584,N_14534);
xnor U15209 (N_15209,N_14928,N_14853);
and U15210 (N_15210,N_14943,N_14638);
xnor U15211 (N_15211,N_14934,N_14793);
or U15212 (N_15212,N_14907,N_14632);
and U15213 (N_15213,N_14574,N_14607);
xnor U15214 (N_15214,N_14895,N_14975);
nand U15215 (N_15215,N_14948,N_14771);
or U15216 (N_15216,N_14926,N_14768);
nand U15217 (N_15217,N_14645,N_14516);
and U15218 (N_15218,N_14802,N_14648);
nor U15219 (N_15219,N_14562,N_14905);
or U15220 (N_15220,N_14792,N_14942);
nand U15221 (N_15221,N_14666,N_14753);
nand U15222 (N_15222,N_14951,N_14617);
xor U15223 (N_15223,N_14604,N_14866);
nor U15224 (N_15224,N_14628,N_14551);
xnor U15225 (N_15225,N_14835,N_14801);
nor U15226 (N_15226,N_14765,N_14676);
nand U15227 (N_15227,N_14957,N_14667);
nor U15228 (N_15228,N_14509,N_14654);
xnor U15229 (N_15229,N_14677,N_14769);
xor U15230 (N_15230,N_14756,N_14622);
nor U15231 (N_15231,N_14530,N_14979);
xnor U15232 (N_15232,N_14541,N_14848);
or U15233 (N_15233,N_14708,N_14964);
nor U15234 (N_15234,N_14947,N_14912);
nor U15235 (N_15235,N_14674,N_14925);
or U15236 (N_15236,N_14815,N_14820);
nand U15237 (N_15237,N_14609,N_14772);
xnor U15238 (N_15238,N_14554,N_14834);
or U15239 (N_15239,N_14959,N_14539);
and U15240 (N_15240,N_14652,N_14819);
nand U15241 (N_15241,N_14817,N_14506);
nand U15242 (N_15242,N_14616,N_14941);
and U15243 (N_15243,N_14812,N_14797);
and U15244 (N_15244,N_14829,N_14744);
xnor U15245 (N_15245,N_14724,N_14806);
xor U15246 (N_15246,N_14544,N_14726);
and U15247 (N_15247,N_14974,N_14686);
nor U15248 (N_15248,N_14824,N_14800);
nor U15249 (N_15249,N_14904,N_14782);
xor U15250 (N_15250,N_14909,N_14565);
nand U15251 (N_15251,N_14704,N_14735);
nand U15252 (N_15252,N_14569,N_14791);
or U15253 (N_15253,N_14587,N_14673);
nor U15254 (N_15254,N_14644,N_14691);
xor U15255 (N_15255,N_14580,N_14820);
nand U15256 (N_15256,N_14606,N_14908);
xnor U15257 (N_15257,N_14936,N_14933);
and U15258 (N_15258,N_14966,N_14875);
or U15259 (N_15259,N_14596,N_14978);
and U15260 (N_15260,N_14781,N_14864);
and U15261 (N_15261,N_14714,N_14517);
nand U15262 (N_15262,N_14820,N_14741);
nor U15263 (N_15263,N_14811,N_14500);
xnor U15264 (N_15264,N_14814,N_14939);
nand U15265 (N_15265,N_14577,N_14561);
or U15266 (N_15266,N_14980,N_14603);
and U15267 (N_15267,N_14542,N_14981);
and U15268 (N_15268,N_14849,N_14588);
nor U15269 (N_15269,N_14749,N_14919);
nand U15270 (N_15270,N_14860,N_14572);
and U15271 (N_15271,N_14543,N_14565);
and U15272 (N_15272,N_14943,N_14796);
nor U15273 (N_15273,N_14873,N_14923);
or U15274 (N_15274,N_14689,N_14851);
xor U15275 (N_15275,N_14710,N_14568);
and U15276 (N_15276,N_14595,N_14848);
or U15277 (N_15277,N_14614,N_14833);
xnor U15278 (N_15278,N_14532,N_14681);
or U15279 (N_15279,N_14743,N_14963);
and U15280 (N_15280,N_14522,N_14709);
or U15281 (N_15281,N_14807,N_14777);
and U15282 (N_15282,N_14787,N_14552);
and U15283 (N_15283,N_14861,N_14683);
xor U15284 (N_15284,N_14957,N_14576);
nand U15285 (N_15285,N_14840,N_14542);
nand U15286 (N_15286,N_14644,N_14945);
and U15287 (N_15287,N_14768,N_14856);
xor U15288 (N_15288,N_14564,N_14643);
xnor U15289 (N_15289,N_14999,N_14730);
and U15290 (N_15290,N_14673,N_14858);
and U15291 (N_15291,N_14598,N_14744);
nor U15292 (N_15292,N_14637,N_14788);
and U15293 (N_15293,N_14842,N_14544);
xnor U15294 (N_15294,N_14524,N_14620);
and U15295 (N_15295,N_14531,N_14948);
or U15296 (N_15296,N_14534,N_14869);
or U15297 (N_15297,N_14706,N_14843);
xnor U15298 (N_15298,N_14743,N_14952);
or U15299 (N_15299,N_14890,N_14768);
xnor U15300 (N_15300,N_14736,N_14851);
or U15301 (N_15301,N_14680,N_14991);
or U15302 (N_15302,N_14827,N_14956);
nand U15303 (N_15303,N_14539,N_14708);
or U15304 (N_15304,N_14672,N_14614);
or U15305 (N_15305,N_14556,N_14509);
xnor U15306 (N_15306,N_14620,N_14831);
nand U15307 (N_15307,N_14694,N_14788);
nor U15308 (N_15308,N_14556,N_14946);
nor U15309 (N_15309,N_14590,N_14977);
xnor U15310 (N_15310,N_14892,N_14974);
and U15311 (N_15311,N_14942,N_14904);
nor U15312 (N_15312,N_14947,N_14519);
nor U15313 (N_15313,N_14910,N_14536);
nand U15314 (N_15314,N_14657,N_14931);
nand U15315 (N_15315,N_14762,N_14598);
or U15316 (N_15316,N_14560,N_14979);
nor U15317 (N_15317,N_14678,N_14840);
nor U15318 (N_15318,N_14583,N_14925);
or U15319 (N_15319,N_14715,N_14759);
xnor U15320 (N_15320,N_14566,N_14696);
xor U15321 (N_15321,N_14816,N_14768);
and U15322 (N_15322,N_14741,N_14982);
xor U15323 (N_15323,N_14549,N_14920);
or U15324 (N_15324,N_14948,N_14642);
nor U15325 (N_15325,N_14580,N_14993);
or U15326 (N_15326,N_14923,N_14697);
nor U15327 (N_15327,N_14544,N_14861);
nor U15328 (N_15328,N_14557,N_14814);
and U15329 (N_15329,N_14554,N_14861);
nand U15330 (N_15330,N_14964,N_14719);
xnor U15331 (N_15331,N_14811,N_14995);
xor U15332 (N_15332,N_14541,N_14868);
xnor U15333 (N_15333,N_14772,N_14683);
xnor U15334 (N_15334,N_14727,N_14784);
nand U15335 (N_15335,N_14951,N_14530);
and U15336 (N_15336,N_14618,N_14682);
xor U15337 (N_15337,N_14569,N_14538);
nor U15338 (N_15338,N_14966,N_14925);
nor U15339 (N_15339,N_14882,N_14905);
nand U15340 (N_15340,N_14557,N_14553);
nand U15341 (N_15341,N_14980,N_14778);
nor U15342 (N_15342,N_14530,N_14770);
and U15343 (N_15343,N_14632,N_14773);
nor U15344 (N_15344,N_14603,N_14648);
or U15345 (N_15345,N_14791,N_14939);
nor U15346 (N_15346,N_14920,N_14956);
nor U15347 (N_15347,N_14836,N_14771);
or U15348 (N_15348,N_14911,N_14721);
and U15349 (N_15349,N_14863,N_14686);
or U15350 (N_15350,N_14635,N_14675);
and U15351 (N_15351,N_14791,N_14597);
or U15352 (N_15352,N_14695,N_14709);
or U15353 (N_15353,N_14813,N_14547);
nor U15354 (N_15354,N_14591,N_14960);
nand U15355 (N_15355,N_14522,N_14951);
or U15356 (N_15356,N_14997,N_14713);
or U15357 (N_15357,N_14849,N_14910);
or U15358 (N_15358,N_14551,N_14706);
and U15359 (N_15359,N_14976,N_14837);
nand U15360 (N_15360,N_14545,N_14829);
or U15361 (N_15361,N_14700,N_14704);
xnor U15362 (N_15362,N_14659,N_14825);
or U15363 (N_15363,N_14785,N_14983);
nand U15364 (N_15364,N_14972,N_14613);
or U15365 (N_15365,N_14502,N_14621);
nor U15366 (N_15366,N_14822,N_14893);
xnor U15367 (N_15367,N_14550,N_14960);
or U15368 (N_15368,N_14668,N_14634);
nor U15369 (N_15369,N_14902,N_14854);
and U15370 (N_15370,N_14595,N_14702);
xor U15371 (N_15371,N_14766,N_14802);
nand U15372 (N_15372,N_14975,N_14918);
and U15373 (N_15373,N_14774,N_14907);
and U15374 (N_15374,N_14582,N_14973);
or U15375 (N_15375,N_14773,N_14621);
nor U15376 (N_15376,N_14604,N_14605);
or U15377 (N_15377,N_14571,N_14527);
or U15378 (N_15378,N_14618,N_14993);
nand U15379 (N_15379,N_14551,N_14590);
and U15380 (N_15380,N_14685,N_14927);
nor U15381 (N_15381,N_14613,N_14654);
nor U15382 (N_15382,N_14704,N_14932);
xnor U15383 (N_15383,N_14610,N_14877);
nor U15384 (N_15384,N_14957,N_14501);
nand U15385 (N_15385,N_14993,N_14995);
nor U15386 (N_15386,N_14670,N_14504);
nor U15387 (N_15387,N_14610,N_14879);
xor U15388 (N_15388,N_14826,N_14637);
or U15389 (N_15389,N_14507,N_14889);
and U15390 (N_15390,N_14853,N_14672);
or U15391 (N_15391,N_14718,N_14560);
xor U15392 (N_15392,N_14697,N_14690);
xnor U15393 (N_15393,N_14659,N_14823);
nor U15394 (N_15394,N_14807,N_14834);
and U15395 (N_15395,N_14881,N_14608);
or U15396 (N_15396,N_14636,N_14761);
nand U15397 (N_15397,N_14839,N_14941);
or U15398 (N_15398,N_14963,N_14932);
or U15399 (N_15399,N_14541,N_14947);
and U15400 (N_15400,N_14900,N_14801);
nor U15401 (N_15401,N_14945,N_14614);
nor U15402 (N_15402,N_14711,N_14599);
and U15403 (N_15403,N_14580,N_14581);
xor U15404 (N_15404,N_14778,N_14692);
nor U15405 (N_15405,N_14631,N_14903);
xor U15406 (N_15406,N_14943,N_14519);
nand U15407 (N_15407,N_14763,N_14996);
or U15408 (N_15408,N_14935,N_14707);
or U15409 (N_15409,N_14594,N_14777);
and U15410 (N_15410,N_14777,N_14721);
xor U15411 (N_15411,N_14602,N_14996);
or U15412 (N_15412,N_14646,N_14942);
or U15413 (N_15413,N_14737,N_14606);
nor U15414 (N_15414,N_14717,N_14855);
nand U15415 (N_15415,N_14747,N_14616);
xor U15416 (N_15416,N_14759,N_14724);
xor U15417 (N_15417,N_14541,N_14662);
and U15418 (N_15418,N_14619,N_14737);
or U15419 (N_15419,N_14753,N_14737);
and U15420 (N_15420,N_14517,N_14905);
and U15421 (N_15421,N_14964,N_14507);
and U15422 (N_15422,N_14884,N_14777);
and U15423 (N_15423,N_14813,N_14556);
nand U15424 (N_15424,N_14985,N_14799);
or U15425 (N_15425,N_14731,N_14607);
nand U15426 (N_15426,N_14946,N_14650);
and U15427 (N_15427,N_14702,N_14862);
nand U15428 (N_15428,N_14903,N_14977);
and U15429 (N_15429,N_14777,N_14875);
nand U15430 (N_15430,N_14508,N_14654);
xor U15431 (N_15431,N_14610,N_14905);
nor U15432 (N_15432,N_14890,N_14884);
nand U15433 (N_15433,N_14872,N_14515);
or U15434 (N_15434,N_14716,N_14552);
nand U15435 (N_15435,N_14914,N_14980);
xnor U15436 (N_15436,N_14813,N_14794);
and U15437 (N_15437,N_14581,N_14937);
nor U15438 (N_15438,N_14980,N_14978);
xor U15439 (N_15439,N_14721,N_14540);
or U15440 (N_15440,N_14543,N_14689);
nor U15441 (N_15441,N_14571,N_14648);
nor U15442 (N_15442,N_14707,N_14842);
nand U15443 (N_15443,N_14802,N_14858);
xor U15444 (N_15444,N_14576,N_14797);
nor U15445 (N_15445,N_14603,N_14751);
nor U15446 (N_15446,N_14829,N_14684);
nor U15447 (N_15447,N_14585,N_14730);
or U15448 (N_15448,N_14941,N_14619);
nor U15449 (N_15449,N_14574,N_14950);
and U15450 (N_15450,N_14813,N_14651);
nand U15451 (N_15451,N_14996,N_14677);
and U15452 (N_15452,N_14654,N_14801);
nor U15453 (N_15453,N_14595,N_14920);
nand U15454 (N_15454,N_14506,N_14737);
or U15455 (N_15455,N_14665,N_14963);
and U15456 (N_15456,N_14826,N_14989);
nand U15457 (N_15457,N_14910,N_14620);
xor U15458 (N_15458,N_14611,N_14933);
nand U15459 (N_15459,N_14966,N_14734);
nand U15460 (N_15460,N_14702,N_14592);
or U15461 (N_15461,N_14985,N_14651);
xor U15462 (N_15462,N_14888,N_14882);
nand U15463 (N_15463,N_14524,N_14873);
xor U15464 (N_15464,N_14661,N_14563);
nand U15465 (N_15465,N_14513,N_14805);
or U15466 (N_15466,N_14761,N_14841);
and U15467 (N_15467,N_14976,N_14741);
xor U15468 (N_15468,N_14607,N_14684);
and U15469 (N_15469,N_14725,N_14957);
and U15470 (N_15470,N_14665,N_14502);
or U15471 (N_15471,N_14734,N_14977);
nor U15472 (N_15472,N_14925,N_14880);
nand U15473 (N_15473,N_14747,N_14627);
and U15474 (N_15474,N_14800,N_14838);
or U15475 (N_15475,N_14950,N_14587);
nand U15476 (N_15476,N_14667,N_14599);
nand U15477 (N_15477,N_14523,N_14506);
nor U15478 (N_15478,N_14992,N_14928);
nand U15479 (N_15479,N_14747,N_14685);
and U15480 (N_15480,N_14863,N_14811);
and U15481 (N_15481,N_14965,N_14956);
and U15482 (N_15482,N_14882,N_14959);
and U15483 (N_15483,N_14981,N_14898);
nand U15484 (N_15484,N_14982,N_14522);
or U15485 (N_15485,N_14679,N_14524);
or U15486 (N_15486,N_14760,N_14977);
xnor U15487 (N_15487,N_14638,N_14851);
nor U15488 (N_15488,N_14639,N_14653);
and U15489 (N_15489,N_14540,N_14981);
or U15490 (N_15490,N_14705,N_14691);
xor U15491 (N_15491,N_14885,N_14979);
nand U15492 (N_15492,N_14918,N_14534);
nor U15493 (N_15493,N_14811,N_14864);
and U15494 (N_15494,N_14576,N_14632);
or U15495 (N_15495,N_14654,N_14909);
nand U15496 (N_15496,N_14814,N_14702);
nand U15497 (N_15497,N_14510,N_14683);
xor U15498 (N_15498,N_14734,N_14650);
and U15499 (N_15499,N_14796,N_14532);
nand U15500 (N_15500,N_15432,N_15294);
nand U15501 (N_15501,N_15301,N_15363);
nor U15502 (N_15502,N_15210,N_15118);
xnor U15503 (N_15503,N_15009,N_15473);
or U15504 (N_15504,N_15231,N_15233);
or U15505 (N_15505,N_15139,N_15239);
and U15506 (N_15506,N_15491,N_15217);
xor U15507 (N_15507,N_15218,N_15168);
xor U15508 (N_15508,N_15484,N_15490);
xnor U15509 (N_15509,N_15090,N_15430);
or U15510 (N_15510,N_15185,N_15415);
nor U15511 (N_15511,N_15469,N_15485);
xor U15512 (N_15512,N_15074,N_15425);
xor U15513 (N_15513,N_15482,N_15406);
or U15514 (N_15514,N_15195,N_15014);
xnor U15515 (N_15515,N_15046,N_15329);
and U15516 (N_15516,N_15311,N_15049);
or U15517 (N_15517,N_15006,N_15033);
xnor U15518 (N_15518,N_15022,N_15105);
nor U15519 (N_15519,N_15480,N_15488);
or U15520 (N_15520,N_15366,N_15325);
nand U15521 (N_15521,N_15212,N_15296);
xnor U15522 (N_15522,N_15287,N_15276);
and U15523 (N_15523,N_15242,N_15310);
or U15524 (N_15524,N_15391,N_15302);
or U15525 (N_15525,N_15267,N_15135);
nor U15526 (N_15526,N_15284,N_15131);
nor U15527 (N_15527,N_15037,N_15385);
xnor U15528 (N_15528,N_15171,N_15120);
or U15529 (N_15529,N_15256,N_15424);
or U15530 (N_15530,N_15305,N_15463);
xor U15531 (N_15531,N_15420,N_15334);
xor U15532 (N_15532,N_15353,N_15297);
nor U15533 (N_15533,N_15290,N_15309);
nand U15534 (N_15534,N_15274,N_15140);
xor U15535 (N_15535,N_15020,N_15495);
or U15536 (N_15536,N_15017,N_15204);
or U15537 (N_15537,N_15054,N_15460);
nor U15538 (N_15538,N_15379,N_15184);
nand U15539 (N_15539,N_15253,N_15499);
xor U15540 (N_15540,N_15081,N_15240);
xnor U15541 (N_15541,N_15373,N_15316);
xor U15542 (N_15542,N_15344,N_15498);
nor U15543 (N_15543,N_15221,N_15361);
and U15544 (N_15544,N_15387,N_15359);
nand U15545 (N_15545,N_15393,N_15289);
xor U15546 (N_15546,N_15132,N_15278);
nor U15547 (N_15547,N_15030,N_15021);
and U15548 (N_15548,N_15157,N_15112);
nor U15549 (N_15549,N_15147,N_15101);
nand U15550 (N_15550,N_15328,N_15422);
and U15551 (N_15551,N_15031,N_15234);
nor U15552 (N_15552,N_15412,N_15126);
and U15553 (N_15553,N_15095,N_15360);
and U15554 (N_15554,N_15461,N_15208);
nand U15555 (N_15555,N_15403,N_15201);
nor U15556 (N_15556,N_15409,N_15151);
xnor U15557 (N_15557,N_15048,N_15141);
nand U15558 (N_15558,N_15323,N_15308);
xnor U15559 (N_15559,N_15179,N_15227);
or U15560 (N_15560,N_15032,N_15164);
or U15561 (N_15561,N_15427,N_15117);
nor U15562 (N_15562,N_15451,N_15470);
or U15563 (N_15563,N_15486,N_15069);
or U15564 (N_15564,N_15155,N_15313);
or U15565 (N_15565,N_15189,N_15439);
nand U15566 (N_15566,N_15483,N_15443);
and U15567 (N_15567,N_15119,N_15161);
and U15568 (N_15568,N_15175,N_15199);
nor U15569 (N_15569,N_15459,N_15364);
and U15570 (N_15570,N_15375,N_15073);
nor U15571 (N_15571,N_15288,N_15307);
and U15572 (N_15572,N_15400,N_15114);
and U15573 (N_15573,N_15177,N_15444);
and U15574 (N_15574,N_15371,N_15350);
or U15575 (N_15575,N_15270,N_15153);
nor U15576 (N_15576,N_15023,N_15041);
xor U15577 (N_15577,N_15143,N_15268);
or U15578 (N_15578,N_15417,N_15413);
or U15579 (N_15579,N_15182,N_15015);
nand U15580 (N_15580,N_15396,N_15247);
or U15581 (N_15581,N_15075,N_15008);
nor U15582 (N_15582,N_15216,N_15255);
nand U15583 (N_15583,N_15079,N_15370);
nand U15584 (N_15584,N_15229,N_15293);
and U15585 (N_15585,N_15192,N_15205);
and U15586 (N_15586,N_15181,N_15038);
or U15587 (N_15587,N_15138,N_15213);
xnor U15588 (N_15588,N_15066,N_15133);
or U15589 (N_15589,N_15282,N_15130);
nor U15590 (N_15590,N_15345,N_15176);
or U15591 (N_15591,N_15449,N_15273);
or U15592 (N_15592,N_15367,N_15222);
and U15593 (N_15593,N_15405,N_15466);
or U15594 (N_15594,N_15381,N_15374);
xnor U15595 (N_15595,N_15028,N_15152);
nor U15596 (N_15596,N_15453,N_15283);
nor U15597 (N_15597,N_15437,N_15378);
or U15598 (N_15598,N_15394,N_15340);
nand U15599 (N_15599,N_15025,N_15377);
xor U15600 (N_15600,N_15388,N_15264);
and U15601 (N_15601,N_15355,N_15115);
nor U15602 (N_15602,N_15298,N_15085);
nor U15603 (N_15603,N_15280,N_15261);
and U15604 (N_15604,N_15193,N_15232);
or U15605 (N_15605,N_15144,N_15376);
nor U15606 (N_15606,N_15122,N_15477);
and U15607 (N_15607,N_15129,N_15436);
nand U15608 (N_15608,N_15326,N_15243);
nand U15609 (N_15609,N_15078,N_15224);
nor U15610 (N_15610,N_15097,N_15497);
nor U15611 (N_15611,N_15348,N_15362);
xor U15612 (N_15612,N_15235,N_15404);
nand U15613 (N_15613,N_15162,N_15013);
nor U15614 (N_15614,N_15089,N_15416);
nor U15615 (N_15615,N_15072,N_15435);
and U15616 (N_15616,N_15431,N_15083);
nor U15617 (N_15617,N_15271,N_15172);
xor U15618 (N_15618,N_15277,N_15029);
nor U15619 (N_15619,N_15197,N_15346);
xor U15620 (N_15620,N_15263,N_15244);
xor U15621 (N_15621,N_15158,N_15440);
nor U15622 (N_15622,N_15342,N_15254);
xor U15623 (N_15623,N_15035,N_15382);
nor U15624 (N_15624,N_15266,N_15214);
xor U15625 (N_15625,N_15170,N_15438);
and U15626 (N_15626,N_15225,N_15414);
xor U15627 (N_15627,N_15055,N_15057);
and U15628 (N_15628,N_15341,N_15462);
or U15629 (N_15629,N_15465,N_15246);
or U15630 (N_15630,N_15471,N_15314);
or U15631 (N_15631,N_15352,N_15300);
xnor U15632 (N_15632,N_15110,N_15335);
or U15633 (N_15633,N_15474,N_15230);
nand U15634 (N_15634,N_15318,N_15368);
nand U15635 (N_15635,N_15019,N_15052);
xor U15636 (N_15636,N_15206,N_15076);
nor U15637 (N_15637,N_15312,N_15454);
nand U15638 (N_15638,N_15339,N_15059);
and U15639 (N_15639,N_15433,N_15160);
nand U15640 (N_15640,N_15149,N_15063);
and U15641 (N_15641,N_15040,N_15426);
nand U15642 (N_15642,N_15408,N_15167);
nand U15643 (N_15643,N_15386,N_15262);
xor U15644 (N_15644,N_15343,N_15450);
or U15645 (N_15645,N_15134,N_15183);
or U15646 (N_15646,N_15203,N_15001);
nand U15647 (N_15647,N_15257,N_15445);
nand U15648 (N_15648,N_15292,N_15324);
xor U15649 (N_15649,N_15291,N_15331);
xnor U15650 (N_15650,N_15036,N_15452);
nand U15651 (N_15651,N_15091,N_15489);
xnor U15652 (N_15652,N_15104,N_15142);
and U15653 (N_15653,N_15125,N_15338);
xnor U15654 (N_15654,N_15281,N_15209);
nand U15655 (N_15655,N_15475,N_15173);
nand U15656 (N_15656,N_15137,N_15456);
nand U15657 (N_15657,N_15457,N_15159);
xor U15658 (N_15658,N_15027,N_15447);
or U15659 (N_15659,N_15087,N_15357);
and U15660 (N_15660,N_15188,N_15395);
and U15661 (N_15661,N_15111,N_15082);
and U15662 (N_15662,N_15496,N_15481);
xnor U15663 (N_15663,N_15306,N_15410);
nor U15664 (N_15664,N_15349,N_15051);
and U15665 (N_15665,N_15319,N_15012);
nand U15666 (N_15666,N_15421,N_15102);
nor U15667 (N_15667,N_15100,N_15320);
or U15668 (N_15668,N_15024,N_15042);
nor U15669 (N_15669,N_15016,N_15441);
and U15670 (N_15670,N_15200,N_15211);
xor U15671 (N_15671,N_15047,N_15464);
xor U15672 (N_15672,N_15002,N_15207);
nor U15673 (N_15673,N_15434,N_15322);
or U15674 (N_15674,N_15468,N_15148);
or U15675 (N_15675,N_15194,N_15249);
and U15676 (N_15676,N_15077,N_15004);
and U15677 (N_15677,N_15067,N_15398);
xnor U15678 (N_15678,N_15223,N_15265);
and U15679 (N_15679,N_15169,N_15044);
or U15680 (N_15680,N_15018,N_15248);
nand U15681 (N_15681,N_15237,N_15088);
and U15682 (N_15682,N_15163,N_15180);
xnor U15683 (N_15683,N_15080,N_15071);
nand U15684 (N_15684,N_15198,N_15442);
and U15685 (N_15685,N_15272,N_15401);
xor U15686 (N_15686,N_15258,N_15092);
and U15687 (N_15687,N_15065,N_15056);
and U15688 (N_15688,N_15127,N_15099);
nand U15689 (N_15689,N_15084,N_15252);
nand U15690 (N_15690,N_15113,N_15116);
nor U15691 (N_15691,N_15124,N_15472);
xnor U15692 (N_15692,N_15384,N_15303);
or U15693 (N_15693,N_15446,N_15423);
nand U15694 (N_15694,N_15103,N_15109);
nor U15695 (N_15695,N_15154,N_15236);
nand U15696 (N_15696,N_15150,N_15333);
xnor U15697 (N_15697,N_15251,N_15347);
nand U15698 (N_15698,N_15005,N_15011);
and U15699 (N_15699,N_15245,N_15178);
and U15700 (N_15700,N_15226,N_15156);
or U15701 (N_15701,N_15215,N_15060);
or U15702 (N_15702,N_15478,N_15330);
xor U15703 (N_15703,N_15007,N_15108);
and U15704 (N_15704,N_15238,N_15128);
and U15705 (N_15705,N_15492,N_15166);
nand U15706 (N_15706,N_15279,N_15383);
and U15707 (N_15707,N_15086,N_15402);
nand U15708 (N_15708,N_15250,N_15487);
or U15709 (N_15709,N_15045,N_15190);
or U15710 (N_15710,N_15145,N_15354);
or U15711 (N_15711,N_15098,N_15275);
and U15712 (N_15712,N_15315,N_15321);
nand U15713 (N_15713,N_15399,N_15332);
and U15714 (N_15714,N_15455,N_15053);
nand U15715 (N_15715,N_15070,N_15043);
or U15716 (N_15716,N_15068,N_15380);
and U15717 (N_15717,N_15372,N_15259);
nand U15718 (N_15718,N_15096,N_15479);
nor U15719 (N_15719,N_15365,N_15003);
xnor U15720 (N_15720,N_15062,N_15304);
xnor U15721 (N_15721,N_15407,N_15327);
xnor U15722 (N_15722,N_15269,N_15220);
and U15723 (N_15723,N_15034,N_15026);
and U15724 (N_15724,N_15295,N_15419);
and U15725 (N_15725,N_15146,N_15392);
or U15726 (N_15726,N_15039,N_15121);
nor U15727 (N_15727,N_15390,N_15428);
or U15728 (N_15728,N_15186,N_15093);
nand U15729 (N_15729,N_15336,N_15467);
and U15730 (N_15730,N_15356,N_15094);
or U15731 (N_15731,N_15050,N_15202);
nand U15732 (N_15732,N_15458,N_15286);
nand U15733 (N_15733,N_15397,N_15000);
nand U15734 (N_15734,N_15010,N_15418);
nand U15735 (N_15735,N_15358,N_15260);
nand U15736 (N_15736,N_15241,N_15493);
and U15737 (N_15737,N_15476,N_15369);
xnor U15738 (N_15738,N_15494,N_15429);
or U15739 (N_15739,N_15191,N_15219);
nor U15740 (N_15740,N_15107,N_15123);
nand U15741 (N_15741,N_15165,N_15389);
nand U15742 (N_15742,N_15448,N_15061);
nand U15743 (N_15743,N_15299,N_15337);
nand U15744 (N_15744,N_15174,N_15196);
xnor U15745 (N_15745,N_15187,N_15106);
and U15746 (N_15746,N_15411,N_15351);
or U15747 (N_15747,N_15058,N_15064);
nor U15748 (N_15748,N_15228,N_15317);
nand U15749 (N_15749,N_15285,N_15136);
nor U15750 (N_15750,N_15331,N_15358);
and U15751 (N_15751,N_15179,N_15394);
nand U15752 (N_15752,N_15160,N_15330);
and U15753 (N_15753,N_15487,N_15187);
nor U15754 (N_15754,N_15181,N_15010);
or U15755 (N_15755,N_15323,N_15420);
nand U15756 (N_15756,N_15022,N_15270);
nor U15757 (N_15757,N_15010,N_15234);
xor U15758 (N_15758,N_15128,N_15425);
nor U15759 (N_15759,N_15260,N_15161);
or U15760 (N_15760,N_15269,N_15008);
nand U15761 (N_15761,N_15200,N_15376);
nand U15762 (N_15762,N_15028,N_15229);
nand U15763 (N_15763,N_15267,N_15147);
nor U15764 (N_15764,N_15214,N_15110);
nor U15765 (N_15765,N_15152,N_15358);
or U15766 (N_15766,N_15120,N_15497);
nand U15767 (N_15767,N_15391,N_15240);
or U15768 (N_15768,N_15176,N_15063);
nor U15769 (N_15769,N_15288,N_15053);
or U15770 (N_15770,N_15400,N_15478);
and U15771 (N_15771,N_15329,N_15178);
nor U15772 (N_15772,N_15393,N_15042);
xor U15773 (N_15773,N_15245,N_15417);
nor U15774 (N_15774,N_15346,N_15333);
or U15775 (N_15775,N_15122,N_15113);
nand U15776 (N_15776,N_15229,N_15441);
xnor U15777 (N_15777,N_15409,N_15445);
nand U15778 (N_15778,N_15334,N_15323);
or U15779 (N_15779,N_15075,N_15386);
nand U15780 (N_15780,N_15096,N_15358);
xor U15781 (N_15781,N_15173,N_15491);
xor U15782 (N_15782,N_15130,N_15374);
nand U15783 (N_15783,N_15382,N_15357);
nor U15784 (N_15784,N_15024,N_15178);
nand U15785 (N_15785,N_15382,N_15249);
nand U15786 (N_15786,N_15284,N_15242);
nand U15787 (N_15787,N_15374,N_15196);
xor U15788 (N_15788,N_15251,N_15423);
xnor U15789 (N_15789,N_15453,N_15157);
and U15790 (N_15790,N_15364,N_15439);
and U15791 (N_15791,N_15470,N_15352);
or U15792 (N_15792,N_15166,N_15320);
xor U15793 (N_15793,N_15239,N_15021);
or U15794 (N_15794,N_15158,N_15157);
nor U15795 (N_15795,N_15069,N_15488);
or U15796 (N_15796,N_15458,N_15467);
xor U15797 (N_15797,N_15210,N_15076);
and U15798 (N_15798,N_15037,N_15052);
xor U15799 (N_15799,N_15185,N_15059);
nand U15800 (N_15800,N_15249,N_15380);
nand U15801 (N_15801,N_15412,N_15200);
nand U15802 (N_15802,N_15203,N_15169);
nor U15803 (N_15803,N_15171,N_15387);
xnor U15804 (N_15804,N_15359,N_15255);
and U15805 (N_15805,N_15448,N_15487);
nand U15806 (N_15806,N_15230,N_15137);
and U15807 (N_15807,N_15188,N_15037);
and U15808 (N_15808,N_15486,N_15412);
nor U15809 (N_15809,N_15111,N_15431);
and U15810 (N_15810,N_15214,N_15205);
nand U15811 (N_15811,N_15317,N_15193);
and U15812 (N_15812,N_15049,N_15425);
and U15813 (N_15813,N_15262,N_15096);
xor U15814 (N_15814,N_15333,N_15031);
or U15815 (N_15815,N_15075,N_15190);
and U15816 (N_15816,N_15320,N_15366);
nor U15817 (N_15817,N_15130,N_15078);
nand U15818 (N_15818,N_15098,N_15171);
nand U15819 (N_15819,N_15267,N_15054);
nor U15820 (N_15820,N_15086,N_15420);
nor U15821 (N_15821,N_15142,N_15433);
nor U15822 (N_15822,N_15331,N_15230);
nand U15823 (N_15823,N_15487,N_15333);
nand U15824 (N_15824,N_15195,N_15132);
and U15825 (N_15825,N_15324,N_15163);
or U15826 (N_15826,N_15467,N_15151);
xnor U15827 (N_15827,N_15213,N_15432);
or U15828 (N_15828,N_15321,N_15225);
and U15829 (N_15829,N_15331,N_15380);
xnor U15830 (N_15830,N_15142,N_15268);
xor U15831 (N_15831,N_15032,N_15455);
xor U15832 (N_15832,N_15022,N_15401);
nand U15833 (N_15833,N_15438,N_15252);
nor U15834 (N_15834,N_15042,N_15012);
nor U15835 (N_15835,N_15325,N_15238);
xnor U15836 (N_15836,N_15433,N_15098);
or U15837 (N_15837,N_15129,N_15240);
nand U15838 (N_15838,N_15269,N_15476);
nor U15839 (N_15839,N_15166,N_15030);
xnor U15840 (N_15840,N_15012,N_15343);
or U15841 (N_15841,N_15497,N_15397);
or U15842 (N_15842,N_15403,N_15406);
or U15843 (N_15843,N_15176,N_15396);
nor U15844 (N_15844,N_15094,N_15160);
xor U15845 (N_15845,N_15250,N_15399);
and U15846 (N_15846,N_15383,N_15192);
xnor U15847 (N_15847,N_15066,N_15335);
or U15848 (N_15848,N_15478,N_15098);
or U15849 (N_15849,N_15483,N_15403);
and U15850 (N_15850,N_15047,N_15203);
or U15851 (N_15851,N_15481,N_15003);
nor U15852 (N_15852,N_15211,N_15002);
xor U15853 (N_15853,N_15226,N_15094);
nand U15854 (N_15854,N_15494,N_15217);
nand U15855 (N_15855,N_15449,N_15069);
xnor U15856 (N_15856,N_15445,N_15326);
xor U15857 (N_15857,N_15370,N_15216);
nand U15858 (N_15858,N_15437,N_15185);
and U15859 (N_15859,N_15204,N_15149);
xnor U15860 (N_15860,N_15362,N_15222);
nor U15861 (N_15861,N_15496,N_15169);
nor U15862 (N_15862,N_15090,N_15247);
or U15863 (N_15863,N_15346,N_15163);
and U15864 (N_15864,N_15432,N_15034);
and U15865 (N_15865,N_15038,N_15420);
nor U15866 (N_15866,N_15123,N_15186);
nor U15867 (N_15867,N_15486,N_15000);
nand U15868 (N_15868,N_15195,N_15430);
nand U15869 (N_15869,N_15122,N_15180);
xnor U15870 (N_15870,N_15263,N_15250);
and U15871 (N_15871,N_15447,N_15024);
nand U15872 (N_15872,N_15267,N_15229);
xor U15873 (N_15873,N_15151,N_15217);
or U15874 (N_15874,N_15434,N_15189);
or U15875 (N_15875,N_15185,N_15279);
xor U15876 (N_15876,N_15178,N_15428);
nor U15877 (N_15877,N_15236,N_15092);
xor U15878 (N_15878,N_15053,N_15126);
and U15879 (N_15879,N_15234,N_15201);
and U15880 (N_15880,N_15319,N_15375);
nand U15881 (N_15881,N_15347,N_15056);
nor U15882 (N_15882,N_15227,N_15026);
nor U15883 (N_15883,N_15431,N_15174);
xnor U15884 (N_15884,N_15130,N_15048);
or U15885 (N_15885,N_15042,N_15106);
xor U15886 (N_15886,N_15157,N_15189);
xnor U15887 (N_15887,N_15306,N_15365);
nand U15888 (N_15888,N_15305,N_15320);
nand U15889 (N_15889,N_15336,N_15025);
nor U15890 (N_15890,N_15121,N_15081);
and U15891 (N_15891,N_15111,N_15426);
and U15892 (N_15892,N_15219,N_15012);
or U15893 (N_15893,N_15235,N_15073);
or U15894 (N_15894,N_15357,N_15009);
or U15895 (N_15895,N_15042,N_15092);
nand U15896 (N_15896,N_15323,N_15077);
nand U15897 (N_15897,N_15216,N_15281);
nand U15898 (N_15898,N_15480,N_15434);
nand U15899 (N_15899,N_15294,N_15024);
or U15900 (N_15900,N_15039,N_15228);
nor U15901 (N_15901,N_15222,N_15106);
nand U15902 (N_15902,N_15335,N_15446);
nor U15903 (N_15903,N_15078,N_15335);
and U15904 (N_15904,N_15217,N_15296);
or U15905 (N_15905,N_15266,N_15069);
and U15906 (N_15906,N_15371,N_15084);
nand U15907 (N_15907,N_15045,N_15412);
nor U15908 (N_15908,N_15406,N_15059);
and U15909 (N_15909,N_15264,N_15119);
xor U15910 (N_15910,N_15054,N_15320);
nor U15911 (N_15911,N_15178,N_15157);
nand U15912 (N_15912,N_15269,N_15179);
or U15913 (N_15913,N_15247,N_15318);
and U15914 (N_15914,N_15389,N_15341);
or U15915 (N_15915,N_15039,N_15415);
or U15916 (N_15916,N_15028,N_15356);
and U15917 (N_15917,N_15003,N_15081);
or U15918 (N_15918,N_15190,N_15173);
nor U15919 (N_15919,N_15441,N_15136);
nor U15920 (N_15920,N_15021,N_15281);
xor U15921 (N_15921,N_15159,N_15448);
and U15922 (N_15922,N_15468,N_15004);
and U15923 (N_15923,N_15303,N_15016);
xor U15924 (N_15924,N_15235,N_15462);
nor U15925 (N_15925,N_15388,N_15042);
or U15926 (N_15926,N_15066,N_15421);
xor U15927 (N_15927,N_15381,N_15288);
nand U15928 (N_15928,N_15032,N_15146);
xor U15929 (N_15929,N_15468,N_15452);
nand U15930 (N_15930,N_15037,N_15215);
and U15931 (N_15931,N_15173,N_15342);
and U15932 (N_15932,N_15066,N_15059);
and U15933 (N_15933,N_15000,N_15352);
and U15934 (N_15934,N_15350,N_15489);
and U15935 (N_15935,N_15480,N_15211);
or U15936 (N_15936,N_15024,N_15430);
nor U15937 (N_15937,N_15028,N_15007);
or U15938 (N_15938,N_15130,N_15006);
and U15939 (N_15939,N_15389,N_15243);
nor U15940 (N_15940,N_15166,N_15315);
nand U15941 (N_15941,N_15036,N_15341);
nand U15942 (N_15942,N_15062,N_15485);
xor U15943 (N_15943,N_15349,N_15183);
nand U15944 (N_15944,N_15108,N_15085);
nand U15945 (N_15945,N_15009,N_15244);
nor U15946 (N_15946,N_15484,N_15201);
xnor U15947 (N_15947,N_15463,N_15035);
nand U15948 (N_15948,N_15194,N_15464);
or U15949 (N_15949,N_15262,N_15326);
nand U15950 (N_15950,N_15106,N_15486);
and U15951 (N_15951,N_15483,N_15212);
xor U15952 (N_15952,N_15496,N_15287);
and U15953 (N_15953,N_15090,N_15143);
and U15954 (N_15954,N_15089,N_15140);
and U15955 (N_15955,N_15030,N_15256);
xor U15956 (N_15956,N_15071,N_15008);
nand U15957 (N_15957,N_15146,N_15302);
nand U15958 (N_15958,N_15495,N_15492);
or U15959 (N_15959,N_15402,N_15003);
nand U15960 (N_15960,N_15401,N_15329);
and U15961 (N_15961,N_15006,N_15120);
nor U15962 (N_15962,N_15365,N_15401);
and U15963 (N_15963,N_15150,N_15068);
and U15964 (N_15964,N_15343,N_15289);
and U15965 (N_15965,N_15015,N_15450);
nand U15966 (N_15966,N_15119,N_15329);
and U15967 (N_15967,N_15031,N_15105);
or U15968 (N_15968,N_15301,N_15059);
nand U15969 (N_15969,N_15410,N_15445);
nor U15970 (N_15970,N_15477,N_15229);
nand U15971 (N_15971,N_15114,N_15002);
xnor U15972 (N_15972,N_15333,N_15227);
and U15973 (N_15973,N_15364,N_15146);
xor U15974 (N_15974,N_15325,N_15196);
or U15975 (N_15975,N_15469,N_15163);
and U15976 (N_15976,N_15310,N_15303);
xnor U15977 (N_15977,N_15267,N_15237);
nor U15978 (N_15978,N_15362,N_15467);
nor U15979 (N_15979,N_15101,N_15458);
or U15980 (N_15980,N_15134,N_15175);
nor U15981 (N_15981,N_15407,N_15129);
xnor U15982 (N_15982,N_15091,N_15301);
nor U15983 (N_15983,N_15043,N_15037);
xnor U15984 (N_15984,N_15441,N_15006);
nor U15985 (N_15985,N_15138,N_15083);
and U15986 (N_15986,N_15280,N_15127);
and U15987 (N_15987,N_15376,N_15083);
or U15988 (N_15988,N_15216,N_15221);
nor U15989 (N_15989,N_15491,N_15354);
xnor U15990 (N_15990,N_15253,N_15279);
xnor U15991 (N_15991,N_15110,N_15305);
and U15992 (N_15992,N_15153,N_15204);
nand U15993 (N_15993,N_15177,N_15187);
or U15994 (N_15994,N_15143,N_15186);
xor U15995 (N_15995,N_15007,N_15184);
xnor U15996 (N_15996,N_15314,N_15262);
xor U15997 (N_15997,N_15146,N_15085);
or U15998 (N_15998,N_15479,N_15127);
xnor U15999 (N_15999,N_15395,N_15155);
xor U16000 (N_16000,N_15735,N_15736);
xor U16001 (N_16001,N_15758,N_15563);
nor U16002 (N_16002,N_15623,N_15667);
or U16003 (N_16003,N_15649,N_15504);
nand U16004 (N_16004,N_15966,N_15848);
nand U16005 (N_16005,N_15600,N_15536);
or U16006 (N_16006,N_15689,N_15850);
xor U16007 (N_16007,N_15816,N_15503);
nor U16008 (N_16008,N_15897,N_15602);
and U16009 (N_16009,N_15896,N_15703);
nor U16010 (N_16010,N_15859,N_15585);
xor U16011 (N_16011,N_15944,N_15864);
xnor U16012 (N_16012,N_15755,N_15799);
or U16013 (N_16013,N_15590,N_15734);
or U16014 (N_16014,N_15541,N_15670);
xor U16015 (N_16015,N_15862,N_15930);
nor U16016 (N_16016,N_15962,N_15565);
or U16017 (N_16017,N_15543,N_15673);
xor U16018 (N_16018,N_15837,N_15745);
or U16019 (N_16019,N_15801,N_15681);
xor U16020 (N_16020,N_15947,N_15676);
xor U16021 (N_16021,N_15885,N_15544);
xnor U16022 (N_16022,N_15639,N_15892);
nand U16023 (N_16023,N_15948,N_15883);
and U16024 (N_16024,N_15636,N_15526);
nor U16025 (N_16025,N_15952,N_15683);
nor U16026 (N_16026,N_15942,N_15559);
or U16027 (N_16027,N_15945,N_15956);
nand U16028 (N_16028,N_15672,N_15566);
and U16029 (N_16029,N_15936,N_15800);
xor U16030 (N_16030,N_15542,N_15949);
nand U16031 (N_16031,N_15824,N_15847);
nand U16032 (N_16032,N_15865,N_15695);
or U16033 (N_16033,N_15669,N_15756);
nand U16034 (N_16034,N_15823,N_15931);
and U16035 (N_16035,N_15884,N_15899);
or U16036 (N_16036,N_15518,N_15707);
xnor U16037 (N_16037,N_15723,N_15797);
or U16038 (N_16038,N_15882,N_15785);
or U16039 (N_16039,N_15713,N_15727);
xor U16040 (N_16040,N_15712,N_15902);
nor U16041 (N_16041,N_15693,N_15992);
and U16042 (N_16042,N_15511,N_15665);
nor U16043 (N_16043,N_15732,N_15617);
xnor U16044 (N_16044,N_15510,N_15920);
and U16045 (N_16045,N_15788,N_15980);
xnor U16046 (N_16046,N_15783,N_15622);
nor U16047 (N_16047,N_15711,N_15630);
and U16048 (N_16048,N_15817,N_15972);
nand U16049 (N_16049,N_15808,N_15915);
nor U16050 (N_16050,N_15615,N_15519);
and U16051 (N_16051,N_15933,N_15644);
and U16052 (N_16052,N_15546,N_15964);
xnor U16053 (N_16053,N_15997,N_15626);
xor U16054 (N_16054,N_15989,N_15564);
nand U16055 (N_16055,N_15886,N_15838);
and U16056 (N_16056,N_15918,N_15879);
nand U16057 (N_16057,N_15582,N_15539);
nand U16058 (N_16058,N_15728,N_15715);
or U16059 (N_16059,N_15769,N_15650);
nand U16060 (N_16060,N_15668,N_15509);
and U16061 (N_16061,N_15993,N_15825);
or U16062 (N_16062,N_15963,N_15973);
nand U16063 (N_16063,N_15770,N_15596);
nand U16064 (N_16064,N_15606,N_15985);
or U16065 (N_16065,N_15893,N_15593);
xor U16066 (N_16066,N_15744,N_15528);
and U16067 (N_16067,N_15595,N_15690);
or U16068 (N_16068,N_15950,N_15999);
nand U16069 (N_16069,N_15926,N_15822);
nand U16070 (N_16070,N_15748,N_15740);
nand U16071 (N_16071,N_15567,N_15522);
and U16072 (N_16072,N_15682,N_15759);
nor U16073 (N_16073,N_15905,N_15558);
nor U16074 (N_16074,N_15638,N_15811);
nor U16075 (N_16075,N_15571,N_15877);
or U16076 (N_16076,N_15588,N_15629);
nand U16077 (N_16077,N_15991,N_15773);
xor U16078 (N_16078,N_15984,N_15694);
and U16079 (N_16079,N_15778,N_15798);
xor U16080 (N_16080,N_15535,N_15821);
or U16081 (N_16081,N_15548,N_15718);
nor U16082 (N_16082,N_15873,N_15790);
or U16083 (N_16083,N_15632,N_15538);
nor U16084 (N_16084,N_15965,N_15525);
or U16085 (N_16085,N_15974,N_15851);
nor U16086 (N_16086,N_15531,N_15975);
and U16087 (N_16087,N_15895,N_15730);
or U16088 (N_16088,N_15854,N_15852);
nor U16089 (N_16089,N_15919,N_15516);
nor U16090 (N_16090,N_15842,N_15860);
or U16091 (N_16091,N_15749,N_15866);
nand U16092 (N_16092,N_15994,N_15584);
xnor U16093 (N_16093,N_15805,N_15520);
nor U16094 (N_16094,N_15507,N_15809);
or U16095 (N_16095,N_15738,N_15601);
nor U16096 (N_16096,N_15917,N_15709);
and U16097 (N_16097,N_15943,N_15951);
or U16098 (N_16098,N_15988,N_15908);
xor U16099 (N_16099,N_15954,N_15836);
nor U16100 (N_16100,N_15910,N_15871);
or U16101 (N_16101,N_15796,N_15935);
nor U16102 (N_16102,N_15764,N_15557);
and U16103 (N_16103,N_15870,N_15970);
xor U16104 (N_16104,N_15998,N_15708);
nor U16105 (N_16105,N_15932,N_15686);
and U16106 (N_16106,N_15657,N_15894);
nand U16107 (N_16107,N_15653,N_15841);
nand U16108 (N_16108,N_15849,N_15826);
and U16109 (N_16109,N_15524,N_15628);
xnor U16110 (N_16110,N_15924,N_15643);
or U16111 (N_16111,N_15699,N_15731);
or U16112 (N_16112,N_15634,N_15791);
and U16113 (N_16113,N_15875,N_15663);
or U16114 (N_16114,N_15804,N_15505);
nor U16115 (N_16115,N_15929,N_15726);
and U16116 (N_16116,N_15645,N_15517);
xor U16117 (N_16117,N_15872,N_15530);
nand U16118 (N_16118,N_15500,N_15685);
nor U16119 (N_16119,N_15705,N_15829);
nand U16120 (N_16120,N_15714,N_15587);
nor U16121 (N_16121,N_15780,N_15752);
and U16122 (N_16122,N_15671,N_15716);
nand U16123 (N_16123,N_15552,N_15968);
and U16124 (N_16124,N_15569,N_15662);
xor U16125 (N_16125,N_15922,N_15815);
nor U16126 (N_16126,N_15818,N_15578);
xnor U16127 (N_16127,N_15573,N_15696);
nor U16128 (N_16128,N_15659,N_15513);
xnor U16129 (N_16129,N_15957,N_15574);
nand U16130 (N_16130,N_15627,N_15666);
xnor U16131 (N_16131,N_15688,N_15655);
nor U16132 (N_16132,N_15594,N_15706);
nor U16133 (N_16133,N_15561,N_15807);
xnor U16134 (N_16134,N_15856,N_15534);
nor U16135 (N_16135,N_15928,N_15921);
xnor U16136 (N_16136,N_15604,N_15609);
nor U16137 (N_16137,N_15772,N_15958);
nor U16138 (N_16138,N_15996,N_15853);
and U16139 (N_16139,N_15967,N_15946);
nor U16140 (N_16140,N_15961,N_15674);
nor U16141 (N_16141,N_15656,N_15890);
xor U16142 (N_16142,N_15642,N_15540);
and U16143 (N_16143,N_15802,N_15925);
nand U16144 (N_16144,N_15907,N_15583);
and U16145 (N_16145,N_15913,N_15608);
xnor U16146 (N_16146,N_15679,N_15855);
or U16147 (N_16147,N_15621,N_15635);
or U16148 (N_16148,N_15739,N_15550);
nand U16149 (N_16149,N_15737,N_15750);
nor U16150 (N_16150,N_15664,N_15580);
nor U16151 (N_16151,N_15793,N_15547);
xor U16152 (N_16152,N_15572,N_15983);
xnor U16153 (N_16153,N_15684,N_15955);
nor U16154 (N_16154,N_15888,N_15813);
nor U16155 (N_16155,N_15979,N_15654);
xor U16156 (N_16156,N_15911,N_15831);
and U16157 (N_16157,N_15576,N_15833);
xor U16158 (N_16158,N_15971,N_15903);
nor U16159 (N_16159,N_15721,N_15941);
xnor U16160 (N_16160,N_15819,N_15789);
and U16161 (N_16161,N_15515,N_15687);
xnor U16162 (N_16162,N_15599,N_15768);
or U16163 (N_16163,N_15904,N_15720);
nor U16164 (N_16164,N_15810,N_15845);
xor U16165 (N_16165,N_15710,N_15795);
nand U16166 (N_16166,N_15959,N_15940);
nand U16167 (N_16167,N_15633,N_15733);
nor U16168 (N_16168,N_15803,N_15960);
and U16169 (N_16169,N_15697,N_15631);
xor U16170 (N_16170,N_15719,N_15501);
or U16171 (N_16171,N_15820,N_15906);
xor U16172 (N_16172,N_15767,N_15577);
xnor U16173 (N_16173,N_15867,N_15828);
nor U16174 (N_16174,N_15912,N_15771);
or U16175 (N_16175,N_15830,N_15614);
xnor U16176 (N_16176,N_15660,N_15506);
nand U16177 (N_16177,N_15640,N_15575);
nand U16178 (N_16178,N_15527,N_15598);
and U16179 (N_16179,N_15746,N_15757);
nor U16180 (N_16180,N_15880,N_15637);
and U16181 (N_16181,N_15909,N_15692);
or U16182 (N_16182,N_15874,N_15939);
xnor U16183 (N_16183,N_15981,N_15512);
xor U16184 (N_16184,N_15938,N_15551);
and U16185 (N_16185,N_15900,N_15765);
or U16186 (N_16186,N_15616,N_15610);
nor U16187 (N_16187,N_15556,N_15953);
nand U16188 (N_16188,N_15562,N_15597);
nand U16189 (N_16189,N_15717,N_15763);
nor U16190 (N_16190,N_15658,N_15700);
nand U16191 (N_16191,N_15647,N_15620);
nand U16192 (N_16192,N_15646,N_15781);
or U16193 (N_16193,N_15982,N_15835);
nor U16194 (N_16194,N_15869,N_15704);
nand U16195 (N_16195,N_15995,N_15502);
nand U16196 (N_16196,N_15651,N_15680);
or U16197 (N_16197,N_15747,N_15891);
nand U16198 (N_16198,N_15529,N_15579);
and U16199 (N_16199,N_15914,N_15827);
and U16200 (N_16200,N_15533,N_15612);
and U16201 (N_16201,N_15987,N_15787);
xnor U16202 (N_16202,N_15678,N_15560);
or U16203 (N_16203,N_15916,N_15592);
and U16204 (N_16204,N_15762,N_15898);
nand U16205 (N_16205,N_15545,N_15652);
nor U16206 (N_16206,N_15549,N_15844);
nand U16207 (N_16207,N_15605,N_15889);
or U16208 (N_16208,N_15753,N_15553);
nor U16209 (N_16209,N_15661,N_15832);
nand U16210 (N_16210,N_15701,N_15846);
xor U16211 (N_16211,N_15969,N_15754);
nor U16212 (N_16212,N_15618,N_15834);
and U16213 (N_16213,N_15868,N_15775);
or U16214 (N_16214,N_15514,N_15641);
and U16215 (N_16215,N_15812,N_15570);
nand U16216 (N_16216,N_15779,N_15603);
and U16217 (N_16217,N_15751,N_15766);
or U16218 (N_16218,N_15843,N_15702);
nor U16219 (N_16219,N_15786,N_15839);
nand U16220 (N_16220,N_15977,N_15806);
or U16221 (N_16221,N_15581,N_15976);
nor U16222 (N_16222,N_15613,N_15792);
xor U16223 (N_16223,N_15523,N_15741);
nand U16224 (N_16224,N_15776,N_15881);
nand U16225 (N_16225,N_15923,N_15782);
xnor U16226 (N_16226,N_15857,N_15937);
or U16227 (N_16227,N_15554,N_15777);
nand U16228 (N_16228,N_15624,N_15648);
and U16229 (N_16229,N_15774,N_15761);
nand U16230 (N_16230,N_15840,N_15537);
xnor U16231 (N_16231,N_15927,N_15625);
nor U16232 (N_16232,N_15521,N_15675);
and U16233 (N_16233,N_15725,N_15532);
nand U16234 (N_16234,N_15698,N_15760);
or U16235 (N_16235,N_15722,N_15887);
xnor U16236 (N_16236,N_15611,N_15591);
xor U16237 (N_16237,N_15691,N_15568);
xnor U16238 (N_16238,N_15742,N_15990);
and U16239 (N_16239,N_15555,N_15619);
or U16240 (N_16240,N_15794,N_15724);
nor U16241 (N_16241,N_15861,N_15858);
and U16242 (N_16242,N_15589,N_15677);
or U16243 (N_16243,N_15934,N_15986);
xor U16244 (N_16244,N_15508,N_15814);
and U16245 (N_16245,N_15876,N_15586);
and U16246 (N_16246,N_15863,N_15784);
or U16247 (N_16247,N_15607,N_15901);
or U16248 (N_16248,N_15729,N_15878);
or U16249 (N_16249,N_15978,N_15743);
nor U16250 (N_16250,N_15769,N_15523);
nand U16251 (N_16251,N_15985,N_15749);
nand U16252 (N_16252,N_15986,N_15901);
nand U16253 (N_16253,N_15654,N_15840);
or U16254 (N_16254,N_15502,N_15620);
and U16255 (N_16255,N_15817,N_15653);
nand U16256 (N_16256,N_15526,N_15511);
and U16257 (N_16257,N_15935,N_15956);
or U16258 (N_16258,N_15755,N_15778);
or U16259 (N_16259,N_15984,N_15560);
and U16260 (N_16260,N_15778,N_15886);
or U16261 (N_16261,N_15583,N_15951);
nand U16262 (N_16262,N_15677,N_15719);
and U16263 (N_16263,N_15530,N_15896);
nand U16264 (N_16264,N_15909,N_15838);
nand U16265 (N_16265,N_15865,N_15950);
and U16266 (N_16266,N_15759,N_15926);
or U16267 (N_16267,N_15798,N_15720);
xnor U16268 (N_16268,N_15553,N_15915);
nor U16269 (N_16269,N_15712,N_15849);
xor U16270 (N_16270,N_15683,N_15793);
or U16271 (N_16271,N_15872,N_15854);
xnor U16272 (N_16272,N_15534,N_15861);
and U16273 (N_16273,N_15692,N_15733);
nand U16274 (N_16274,N_15795,N_15673);
and U16275 (N_16275,N_15666,N_15969);
and U16276 (N_16276,N_15714,N_15724);
and U16277 (N_16277,N_15841,N_15961);
nand U16278 (N_16278,N_15722,N_15855);
or U16279 (N_16279,N_15769,N_15521);
nand U16280 (N_16280,N_15755,N_15990);
or U16281 (N_16281,N_15539,N_15585);
nand U16282 (N_16282,N_15664,N_15724);
and U16283 (N_16283,N_15540,N_15755);
nand U16284 (N_16284,N_15833,N_15807);
and U16285 (N_16285,N_15783,N_15957);
nand U16286 (N_16286,N_15768,N_15569);
xnor U16287 (N_16287,N_15618,N_15531);
and U16288 (N_16288,N_15982,N_15836);
or U16289 (N_16289,N_15588,N_15803);
nor U16290 (N_16290,N_15594,N_15882);
xnor U16291 (N_16291,N_15630,N_15675);
xor U16292 (N_16292,N_15907,N_15664);
xnor U16293 (N_16293,N_15713,N_15951);
nand U16294 (N_16294,N_15834,N_15996);
nand U16295 (N_16295,N_15596,N_15617);
or U16296 (N_16296,N_15916,N_15714);
nor U16297 (N_16297,N_15641,N_15668);
and U16298 (N_16298,N_15636,N_15876);
and U16299 (N_16299,N_15734,N_15691);
and U16300 (N_16300,N_15654,N_15699);
and U16301 (N_16301,N_15579,N_15500);
or U16302 (N_16302,N_15984,N_15726);
and U16303 (N_16303,N_15533,N_15536);
nand U16304 (N_16304,N_15747,N_15666);
and U16305 (N_16305,N_15833,N_15818);
or U16306 (N_16306,N_15842,N_15848);
nor U16307 (N_16307,N_15650,N_15542);
and U16308 (N_16308,N_15925,N_15814);
or U16309 (N_16309,N_15550,N_15926);
xnor U16310 (N_16310,N_15543,N_15836);
or U16311 (N_16311,N_15710,N_15650);
or U16312 (N_16312,N_15537,N_15990);
nor U16313 (N_16313,N_15966,N_15685);
or U16314 (N_16314,N_15510,N_15638);
and U16315 (N_16315,N_15985,N_15978);
or U16316 (N_16316,N_15830,N_15551);
nand U16317 (N_16317,N_15924,N_15570);
and U16318 (N_16318,N_15938,N_15607);
or U16319 (N_16319,N_15971,N_15668);
nor U16320 (N_16320,N_15817,N_15926);
xnor U16321 (N_16321,N_15522,N_15883);
xor U16322 (N_16322,N_15519,N_15668);
xor U16323 (N_16323,N_15507,N_15547);
nand U16324 (N_16324,N_15668,N_15654);
nand U16325 (N_16325,N_15861,N_15848);
or U16326 (N_16326,N_15869,N_15855);
xnor U16327 (N_16327,N_15858,N_15984);
or U16328 (N_16328,N_15802,N_15948);
nand U16329 (N_16329,N_15579,N_15619);
nand U16330 (N_16330,N_15833,N_15902);
nor U16331 (N_16331,N_15720,N_15733);
nand U16332 (N_16332,N_15652,N_15867);
nor U16333 (N_16333,N_15852,N_15863);
xor U16334 (N_16334,N_15894,N_15644);
nor U16335 (N_16335,N_15687,N_15920);
and U16336 (N_16336,N_15615,N_15679);
or U16337 (N_16337,N_15982,N_15511);
and U16338 (N_16338,N_15857,N_15725);
nand U16339 (N_16339,N_15760,N_15578);
nand U16340 (N_16340,N_15681,N_15588);
nor U16341 (N_16341,N_15752,N_15699);
and U16342 (N_16342,N_15829,N_15863);
and U16343 (N_16343,N_15830,N_15967);
xor U16344 (N_16344,N_15922,N_15715);
and U16345 (N_16345,N_15586,N_15732);
and U16346 (N_16346,N_15625,N_15830);
nor U16347 (N_16347,N_15812,N_15671);
nor U16348 (N_16348,N_15669,N_15900);
and U16349 (N_16349,N_15841,N_15839);
xnor U16350 (N_16350,N_15862,N_15518);
or U16351 (N_16351,N_15644,N_15937);
nand U16352 (N_16352,N_15987,N_15576);
and U16353 (N_16353,N_15590,N_15639);
xor U16354 (N_16354,N_15674,N_15921);
and U16355 (N_16355,N_15863,N_15759);
or U16356 (N_16356,N_15536,N_15979);
or U16357 (N_16357,N_15562,N_15606);
and U16358 (N_16358,N_15620,N_15742);
or U16359 (N_16359,N_15811,N_15731);
and U16360 (N_16360,N_15621,N_15962);
or U16361 (N_16361,N_15506,N_15517);
xnor U16362 (N_16362,N_15653,N_15688);
xnor U16363 (N_16363,N_15636,N_15692);
nor U16364 (N_16364,N_15610,N_15693);
nor U16365 (N_16365,N_15742,N_15524);
xor U16366 (N_16366,N_15792,N_15917);
or U16367 (N_16367,N_15512,N_15561);
nand U16368 (N_16368,N_15862,N_15607);
or U16369 (N_16369,N_15647,N_15850);
nand U16370 (N_16370,N_15531,N_15729);
or U16371 (N_16371,N_15827,N_15565);
nand U16372 (N_16372,N_15863,N_15765);
or U16373 (N_16373,N_15759,N_15839);
xnor U16374 (N_16374,N_15886,N_15676);
nor U16375 (N_16375,N_15658,N_15751);
and U16376 (N_16376,N_15900,N_15884);
or U16377 (N_16377,N_15680,N_15541);
and U16378 (N_16378,N_15832,N_15586);
xnor U16379 (N_16379,N_15968,N_15582);
or U16380 (N_16380,N_15934,N_15508);
xor U16381 (N_16381,N_15702,N_15603);
nor U16382 (N_16382,N_15987,N_15912);
and U16383 (N_16383,N_15596,N_15915);
nor U16384 (N_16384,N_15686,N_15736);
xor U16385 (N_16385,N_15980,N_15533);
xor U16386 (N_16386,N_15937,N_15537);
or U16387 (N_16387,N_15806,N_15925);
or U16388 (N_16388,N_15863,N_15869);
xnor U16389 (N_16389,N_15845,N_15992);
or U16390 (N_16390,N_15512,N_15700);
nor U16391 (N_16391,N_15773,N_15695);
or U16392 (N_16392,N_15701,N_15503);
and U16393 (N_16393,N_15932,N_15769);
and U16394 (N_16394,N_15591,N_15681);
or U16395 (N_16395,N_15998,N_15626);
and U16396 (N_16396,N_15975,N_15508);
nor U16397 (N_16397,N_15941,N_15899);
or U16398 (N_16398,N_15656,N_15644);
nor U16399 (N_16399,N_15723,N_15805);
or U16400 (N_16400,N_15955,N_15507);
nor U16401 (N_16401,N_15604,N_15555);
xor U16402 (N_16402,N_15586,N_15601);
nor U16403 (N_16403,N_15587,N_15520);
nand U16404 (N_16404,N_15725,N_15740);
nor U16405 (N_16405,N_15985,N_15701);
nor U16406 (N_16406,N_15559,N_15803);
nor U16407 (N_16407,N_15939,N_15780);
xnor U16408 (N_16408,N_15511,N_15828);
and U16409 (N_16409,N_15889,N_15999);
nand U16410 (N_16410,N_15836,N_15813);
nand U16411 (N_16411,N_15623,N_15740);
and U16412 (N_16412,N_15778,N_15968);
and U16413 (N_16413,N_15766,N_15771);
or U16414 (N_16414,N_15797,N_15884);
xor U16415 (N_16415,N_15720,N_15749);
nor U16416 (N_16416,N_15636,N_15585);
and U16417 (N_16417,N_15732,N_15954);
nand U16418 (N_16418,N_15526,N_15543);
or U16419 (N_16419,N_15556,N_15901);
or U16420 (N_16420,N_15651,N_15909);
xnor U16421 (N_16421,N_15566,N_15873);
or U16422 (N_16422,N_15964,N_15524);
xnor U16423 (N_16423,N_15726,N_15861);
xnor U16424 (N_16424,N_15602,N_15561);
nor U16425 (N_16425,N_15976,N_15854);
xnor U16426 (N_16426,N_15701,N_15728);
xnor U16427 (N_16427,N_15858,N_15538);
xnor U16428 (N_16428,N_15529,N_15510);
or U16429 (N_16429,N_15681,N_15941);
and U16430 (N_16430,N_15994,N_15902);
or U16431 (N_16431,N_15960,N_15621);
nand U16432 (N_16432,N_15871,N_15579);
and U16433 (N_16433,N_15817,N_15542);
and U16434 (N_16434,N_15530,N_15875);
nand U16435 (N_16435,N_15532,N_15573);
nand U16436 (N_16436,N_15769,N_15722);
or U16437 (N_16437,N_15574,N_15911);
nand U16438 (N_16438,N_15885,N_15696);
and U16439 (N_16439,N_15629,N_15905);
or U16440 (N_16440,N_15988,N_15800);
xnor U16441 (N_16441,N_15655,N_15907);
or U16442 (N_16442,N_15884,N_15927);
xnor U16443 (N_16443,N_15963,N_15822);
or U16444 (N_16444,N_15753,N_15613);
nor U16445 (N_16445,N_15572,N_15939);
and U16446 (N_16446,N_15515,N_15991);
or U16447 (N_16447,N_15511,N_15541);
nand U16448 (N_16448,N_15883,N_15502);
or U16449 (N_16449,N_15832,N_15973);
and U16450 (N_16450,N_15625,N_15709);
xnor U16451 (N_16451,N_15960,N_15530);
or U16452 (N_16452,N_15586,N_15788);
xor U16453 (N_16453,N_15796,N_15967);
xnor U16454 (N_16454,N_15792,N_15601);
or U16455 (N_16455,N_15845,N_15575);
nor U16456 (N_16456,N_15873,N_15898);
or U16457 (N_16457,N_15729,N_15551);
or U16458 (N_16458,N_15582,N_15505);
nand U16459 (N_16459,N_15601,N_15643);
nand U16460 (N_16460,N_15843,N_15695);
and U16461 (N_16461,N_15847,N_15506);
or U16462 (N_16462,N_15979,N_15565);
or U16463 (N_16463,N_15524,N_15654);
nor U16464 (N_16464,N_15919,N_15909);
and U16465 (N_16465,N_15848,N_15734);
or U16466 (N_16466,N_15898,N_15986);
and U16467 (N_16467,N_15640,N_15809);
nor U16468 (N_16468,N_15724,N_15597);
xnor U16469 (N_16469,N_15652,N_15823);
xor U16470 (N_16470,N_15942,N_15661);
and U16471 (N_16471,N_15762,N_15700);
and U16472 (N_16472,N_15707,N_15803);
and U16473 (N_16473,N_15510,N_15794);
nand U16474 (N_16474,N_15716,N_15873);
nor U16475 (N_16475,N_15921,N_15572);
nand U16476 (N_16476,N_15698,N_15527);
nor U16477 (N_16477,N_15875,N_15768);
or U16478 (N_16478,N_15946,N_15960);
or U16479 (N_16479,N_15573,N_15993);
and U16480 (N_16480,N_15905,N_15782);
or U16481 (N_16481,N_15986,N_15938);
xor U16482 (N_16482,N_15968,N_15575);
nand U16483 (N_16483,N_15914,N_15652);
nor U16484 (N_16484,N_15718,N_15944);
xor U16485 (N_16485,N_15914,N_15518);
nor U16486 (N_16486,N_15595,N_15610);
or U16487 (N_16487,N_15534,N_15781);
xor U16488 (N_16488,N_15862,N_15884);
and U16489 (N_16489,N_15647,N_15993);
nor U16490 (N_16490,N_15755,N_15787);
nand U16491 (N_16491,N_15817,N_15679);
or U16492 (N_16492,N_15929,N_15801);
xnor U16493 (N_16493,N_15703,N_15695);
or U16494 (N_16494,N_15664,N_15795);
nor U16495 (N_16495,N_15618,N_15793);
nor U16496 (N_16496,N_15607,N_15693);
xnor U16497 (N_16497,N_15850,N_15690);
xnor U16498 (N_16498,N_15588,N_15998);
xnor U16499 (N_16499,N_15928,N_15565);
nor U16500 (N_16500,N_16167,N_16331);
or U16501 (N_16501,N_16321,N_16459);
nand U16502 (N_16502,N_16018,N_16009);
and U16503 (N_16503,N_16270,N_16303);
and U16504 (N_16504,N_16186,N_16230);
nor U16505 (N_16505,N_16235,N_16098);
xor U16506 (N_16506,N_16236,N_16240);
and U16507 (N_16507,N_16277,N_16266);
nor U16508 (N_16508,N_16374,N_16182);
and U16509 (N_16509,N_16088,N_16008);
nor U16510 (N_16510,N_16205,N_16347);
or U16511 (N_16511,N_16258,N_16226);
xnor U16512 (N_16512,N_16125,N_16464);
nor U16513 (N_16513,N_16492,N_16245);
nor U16514 (N_16514,N_16308,N_16419);
xnor U16515 (N_16515,N_16070,N_16227);
nand U16516 (N_16516,N_16335,N_16007);
xnor U16517 (N_16517,N_16283,N_16072);
xnor U16518 (N_16518,N_16327,N_16407);
nand U16519 (N_16519,N_16218,N_16472);
nor U16520 (N_16520,N_16267,N_16163);
nor U16521 (N_16521,N_16409,N_16176);
or U16522 (N_16522,N_16121,N_16362);
nand U16523 (N_16523,N_16164,N_16402);
and U16524 (N_16524,N_16463,N_16170);
nand U16525 (N_16525,N_16027,N_16153);
xor U16526 (N_16526,N_16467,N_16032);
nor U16527 (N_16527,N_16221,N_16297);
or U16528 (N_16528,N_16312,N_16006);
nor U16529 (N_16529,N_16063,N_16275);
nand U16530 (N_16530,N_16204,N_16049);
nor U16531 (N_16531,N_16333,N_16002);
or U16532 (N_16532,N_16054,N_16106);
and U16533 (N_16533,N_16260,N_16396);
and U16534 (N_16534,N_16116,N_16271);
nand U16535 (N_16535,N_16013,N_16352);
nand U16536 (N_16536,N_16279,N_16247);
xnor U16537 (N_16537,N_16102,N_16147);
or U16538 (N_16538,N_16250,N_16446);
and U16539 (N_16539,N_16034,N_16484);
nand U16540 (N_16540,N_16497,N_16046);
nand U16541 (N_16541,N_16051,N_16242);
and U16542 (N_16542,N_16315,N_16078);
nand U16543 (N_16543,N_16356,N_16265);
or U16544 (N_16544,N_16138,N_16041);
and U16545 (N_16545,N_16491,N_16365);
xnor U16546 (N_16546,N_16338,N_16089);
nand U16547 (N_16547,N_16152,N_16208);
nand U16548 (N_16548,N_16367,N_16456);
and U16549 (N_16549,N_16068,N_16393);
xnor U16550 (N_16550,N_16418,N_16022);
nor U16551 (N_16551,N_16263,N_16398);
or U16552 (N_16552,N_16177,N_16012);
and U16553 (N_16553,N_16290,N_16423);
and U16554 (N_16554,N_16123,N_16000);
or U16555 (N_16555,N_16129,N_16136);
and U16556 (N_16556,N_16162,N_16376);
or U16557 (N_16557,N_16103,N_16132);
nor U16558 (N_16558,N_16209,N_16118);
xor U16559 (N_16559,N_16028,N_16062);
nor U16560 (N_16560,N_16415,N_16380);
and U16561 (N_16561,N_16206,N_16498);
or U16562 (N_16562,N_16092,N_16035);
xor U16563 (N_16563,N_16053,N_16172);
xnor U16564 (N_16564,N_16391,N_16159);
or U16565 (N_16565,N_16410,N_16499);
nand U16566 (N_16566,N_16495,N_16431);
nand U16567 (N_16567,N_16289,N_16274);
nor U16568 (N_16568,N_16420,N_16453);
nand U16569 (N_16569,N_16366,N_16481);
and U16570 (N_16570,N_16430,N_16069);
xnor U16571 (N_16571,N_16476,N_16071);
xor U16572 (N_16572,N_16417,N_16108);
nand U16573 (N_16573,N_16211,N_16318);
nand U16574 (N_16574,N_16044,N_16451);
nand U16575 (N_16575,N_16440,N_16193);
xnor U16576 (N_16576,N_16201,N_16364);
nor U16577 (N_16577,N_16157,N_16389);
xnor U16578 (N_16578,N_16355,N_16181);
or U16579 (N_16579,N_16300,N_16128);
or U16580 (N_16580,N_16405,N_16220);
nand U16581 (N_16581,N_16319,N_16166);
or U16582 (N_16582,N_16252,N_16349);
or U16583 (N_16583,N_16486,N_16408);
or U16584 (N_16584,N_16056,N_16134);
nand U16585 (N_16585,N_16400,N_16082);
nor U16586 (N_16586,N_16381,N_16229);
or U16587 (N_16587,N_16392,N_16388);
nand U16588 (N_16588,N_16328,N_16048);
xnor U16589 (N_16589,N_16443,N_16097);
and U16590 (N_16590,N_16360,N_16469);
nor U16591 (N_16591,N_16248,N_16199);
or U16592 (N_16592,N_16494,N_16038);
xnor U16593 (N_16593,N_16188,N_16212);
nand U16594 (N_16594,N_16496,N_16363);
or U16595 (N_16595,N_16219,N_16313);
and U16596 (N_16596,N_16004,N_16351);
xor U16597 (N_16597,N_16194,N_16447);
and U16598 (N_16598,N_16401,N_16302);
and U16599 (N_16599,N_16354,N_16042);
nand U16600 (N_16600,N_16026,N_16369);
xor U16601 (N_16601,N_16117,N_16285);
nor U16602 (N_16602,N_16382,N_16168);
or U16603 (N_16603,N_16478,N_16146);
or U16604 (N_16604,N_16251,N_16386);
and U16605 (N_16605,N_16019,N_16175);
and U16606 (N_16606,N_16413,N_16073);
or U16607 (N_16607,N_16210,N_16390);
nor U16608 (N_16608,N_16003,N_16173);
and U16609 (N_16609,N_16133,N_16010);
xnor U16610 (N_16610,N_16406,N_16301);
nor U16611 (N_16611,N_16294,N_16100);
or U16612 (N_16612,N_16341,N_16231);
and U16613 (N_16613,N_16024,N_16436);
xor U16614 (N_16614,N_16334,N_16373);
and U16615 (N_16615,N_16330,N_16130);
or U16616 (N_16616,N_16150,N_16145);
or U16617 (N_16617,N_16115,N_16343);
or U16618 (N_16618,N_16375,N_16259);
or U16619 (N_16619,N_16438,N_16113);
and U16620 (N_16620,N_16021,N_16090);
or U16621 (N_16621,N_16445,N_16482);
and U16622 (N_16622,N_16067,N_16353);
nor U16623 (N_16623,N_16148,N_16262);
xor U16624 (N_16624,N_16404,N_16191);
nand U16625 (N_16625,N_16213,N_16025);
nor U16626 (N_16626,N_16239,N_16087);
nand U16627 (N_16627,N_16298,N_16096);
or U16628 (N_16628,N_16122,N_16377);
xor U16629 (N_16629,N_16269,N_16109);
or U16630 (N_16630,N_16348,N_16457);
nor U16631 (N_16631,N_16387,N_16383);
nor U16632 (N_16632,N_16394,N_16254);
and U16633 (N_16633,N_16340,N_16143);
xnor U16634 (N_16634,N_16075,N_16261);
xnor U16635 (N_16635,N_16095,N_16237);
nand U16636 (N_16636,N_16149,N_16414);
or U16637 (N_16637,N_16358,N_16399);
nor U16638 (N_16638,N_16310,N_16015);
xnor U16639 (N_16639,N_16005,N_16155);
or U16640 (N_16640,N_16344,N_16187);
or U16641 (N_16641,N_16077,N_16085);
nand U16642 (N_16642,N_16161,N_16223);
or U16643 (N_16643,N_16475,N_16485);
nor U16644 (N_16644,N_16299,N_16435);
and U16645 (N_16645,N_16337,N_16238);
and U16646 (N_16646,N_16076,N_16083);
or U16647 (N_16647,N_16370,N_16437);
nor U16648 (N_16648,N_16416,N_16196);
xor U16649 (N_16649,N_16441,N_16342);
xnor U16650 (N_16650,N_16309,N_16105);
nor U16651 (N_16651,N_16452,N_16180);
xnor U16652 (N_16652,N_16139,N_16215);
and U16653 (N_16653,N_16140,N_16224);
and U16654 (N_16654,N_16253,N_16099);
xnor U16655 (N_16655,N_16074,N_16110);
and U16656 (N_16656,N_16178,N_16378);
xnor U16657 (N_16657,N_16061,N_16185);
or U16658 (N_16658,N_16489,N_16306);
nand U16659 (N_16659,N_16124,N_16039);
and U16660 (N_16660,N_16084,N_16473);
xnor U16661 (N_16661,N_16278,N_16086);
xor U16662 (N_16662,N_16477,N_16411);
nor U16663 (N_16663,N_16280,N_16284);
or U16664 (N_16664,N_16059,N_16273);
and U16665 (N_16665,N_16192,N_16169);
nand U16666 (N_16666,N_16058,N_16030);
or U16667 (N_16667,N_16043,N_16322);
nand U16668 (N_16668,N_16001,N_16055);
nor U16669 (N_16669,N_16326,N_16346);
and U16670 (N_16670,N_16428,N_16427);
xnor U16671 (N_16671,N_16144,N_16444);
or U16672 (N_16672,N_16426,N_16281);
xnor U16673 (N_16673,N_16455,N_16357);
nor U16674 (N_16674,N_16060,N_16305);
and U16675 (N_16675,N_16079,N_16243);
or U16676 (N_16676,N_16291,N_16040);
or U16677 (N_16677,N_16127,N_16244);
nor U16678 (N_16678,N_16225,N_16135);
and U16679 (N_16679,N_16307,N_16200);
or U16680 (N_16680,N_16422,N_16372);
xor U16681 (N_16681,N_16222,N_16037);
and U16682 (N_16682,N_16017,N_16432);
and U16683 (N_16683,N_16036,N_16421);
nand U16684 (N_16684,N_16450,N_16470);
nor U16685 (N_16685,N_16429,N_16057);
or U16686 (N_16686,N_16268,N_16490);
and U16687 (N_16687,N_16296,N_16190);
or U16688 (N_16688,N_16462,N_16320);
nor U16689 (N_16689,N_16295,N_16207);
and U16690 (N_16690,N_16233,N_16137);
xnor U16691 (N_16691,N_16126,N_16214);
nand U16692 (N_16692,N_16151,N_16114);
or U16693 (N_16693,N_16276,N_16286);
nand U16694 (N_16694,N_16120,N_16434);
xnor U16695 (N_16695,N_16045,N_16460);
xnor U16696 (N_16696,N_16493,N_16241);
nor U16697 (N_16697,N_16094,N_16292);
or U16698 (N_16698,N_16131,N_16471);
xnor U16699 (N_16699,N_16234,N_16154);
or U16700 (N_16700,N_16016,N_16111);
and U16701 (N_16701,N_16158,N_16112);
or U16702 (N_16702,N_16107,N_16314);
or U16703 (N_16703,N_16316,N_16014);
nand U16704 (N_16704,N_16179,N_16104);
nand U16705 (N_16705,N_16202,N_16332);
and U16706 (N_16706,N_16361,N_16449);
or U16707 (N_16707,N_16119,N_16461);
or U16708 (N_16708,N_16091,N_16439);
nor U16709 (N_16709,N_16256,N_16384);
and U16710 (N_16710,N_16282,N_16198);
xnor U16711 (N_16711,N_16195,N_16011);
nor U16712 (N_16712,N_16228,N_16257);
nand U16713 (N_16713,N_16047,N_16329);
xnor U16714 (N_16714,N_16424,N_16050);
or U16715 (N_16715,N_16156,N_16080);
nand U16716 (N_16716,N_16217,N_16488);
nor U16717 (N_16717,N_16397,N_16336);
xor U16718 (N_16718,N_16317,N_16345);
nor U16719 (N_16719,N_16466,N_16324);
xnor U16720 (N_16720,N_16368,N_16448);
nand U16721 (N_16721,N_16171,N_16165);
xnor U16722 (N_16722,N_16385,N_16197);
nor U16723 (N_16723,N_16183,N_16052);
and U16724 (N_16724,N_16272,N_16474);
and U16725 (N_16725,N_16468,N_16033);
nand U16726 (N_16726,N_16288,N_16189);
nand U16727 (N_16727,N_16425,N_16479);
xor U16728 (N_16728,N_16412,N_16325);
nand U16729 (N_16729,N_16246,N_16184);
nor U16730 (N_16730,N_16031,N_16293);
or U16731 (N_16731,N_16483,N_16304);
xnor U16732 (N_16732,N_16023,N_16174);
nor U16733 (N_16733,N_16264,N_16081);
and U16734 (N_16734,N_16395,N_16287);
nor U16735 (N_16735,N_16066,N_16458);
nand U16736 (N_16736,N_16480,N_16216);
nor U16737 (N_16737,N_16160,N_16065);
or U16738 (N_16738,N_16487,N_16311);
xor U16739 (N_16739,N_16350,N_16101);
xnor U16740 (N_16740,N_16454,N_16403);
and U16741 (N_16741,N_16371,N_16255);
nand U16742 (N_16742,N_16141,N_16020);
nand U16743 (N_16743,N_16064,N_16142);
and U16744 (N_16744,N_16323,N_16029);
xnor U16745 (N_16745,N_16249,N_16359);
or U16746 (N_16746,N_16379,N_16465);
and U16747 (N_16747,N_16339,N_16442);
or U16748 (N_16748,N_16433,N_16203);
xnor U16749 (N_16749,N_16093,N_16232);
and U16750 (N_16750,N_16261,N_16422);
or U16751 (N_16751,N_16236,N_16014);
and U16752 (N_16752,N_16475,N_16265);
nor U16753 (N_16753,N_16180,N_16403);
xor U16754 (N_16754,N_16220,N_16352);
nand U16755 (N_16755,N_16007,N_16175);
nand U16756 (N_16756,N_16246,N_16129);
and U16757 (N_16757,N_16079,N_16405);
xnor U16758 (N_16758,N_16028,N_16321);
and U16759 (N_16759,N_16136,N_16124);
nor U16760 (N_16760,N_16197,N_16356);
or U16761 (N_16761,N_16207,N_16246);
and U16762 (N_16762,N_16299,N_16136);
or U16763 (N_16763,N_16099,N_16174);
or U16764 (N_16764,N_16077,N_16293);
nand U16765 (N_16765,N_16247,N_16363);
xor U16766 (N_16766,N_16233,N_16269);
or U16767 (N_16767,N_16013,N_16391);
or U16768 (N_16768,N_16275,N_16189);
or U16769 (N_16769,N_16346,N_16097);
xor U16770 (N_16770,N_16201,N_16032);
and U16771 (N_16771,N_16442,N_16184);
nand U16772 (N_16772,N_16230,N_16317);
xnor U16773 (N_16773,N_16212,N_16047);
nand U16774 (N_16774,N_16256,N_16347);
nor U16775 (N_16775,N_16087,N_16262);
and U16776 (N_16776,N_16376,N_16173);
nand U16777 (N_16777,N_16084,N_16377);
xor U16778 (N_16778,N_16096,N_16312);
nand U16779 (N_16779,N_16357,N_16416);
xor U16780 (N_16780,N_16112,N_16469);
and U16781 (N_16781,N_16288,N_16091);
and U16782 (N_16782,N_16395,N_16495);
nor U16783 (N_16783,N_16074,N_16399);
nor U16784 (N_16784,N_16390,N_16492);
or U16785 (N_16785,N_16327,N_16395);
nand U16786 (N_16786,N_16164,N_16250);
or U16787 (N_16787,N_16352,N_16341);
or U16788 (N_16788,N_16411,N_16275);
nand U16789 (N_16789,N_16100,N_16027);
nand U16790 (N_16790,N_16032,N_16401);
nor U16791 (N_16791,N_16404,N_16366);
nor U16792 (N_16792,N_16171,N_16184);
nand U16793 (N_16793,N_16199,N_16227);
and U16794 (N_16794,N_16104,N_16259);
and U16795 (N_16795,N_16334,N_16026);
and U16796 (N_16796,N_16185,N_16225);
xnor U16797 (N_16797,N_16138,N_16380);
and U16798 (N_16798,N_16256,N_16135);
xor U16799 (N_16799,N_16334,N_16149);
nand U16800 (N_16800,N_16210,N_16416);
and U16801 (N_16801,N_16045,N_16148);
or U16802 (N_16802,N_16041,N_16047);
and U16803 (N_16803,N_16157,N_16146);
nand U16804 (N_16804,N_16233,N_16001);
nor U16805 (N_16805,N_16139,N_16304);
xor U16806 (N_16806,N_16222,N_16040);
or U16807 (N_16807,N_16299,N_16342);
nor U16808 (N_16808,N_16491,N_16076);
and U16809 (N_16809,N_16031,N_16180);
or U16810 (N_16810,N_16001,N_16356);
nand U16811 (N_16811,N_16155,N_16238);
nor U16812 (N_16812,N_16258,N_16196);
nor U16813 (N_16813,N_16307,N_16148);
and U16814 (N_16814,N_16180,N_16333);
and U16815 (N_16815,N_16115,N_16419);
nand U16816 (N_16816,N_16292,N_16253);
or U16817 (N_16817,N_16207,N_16067);
and U16818 (N_16818,N_16083,N_16073);
nor U16819 (N_16819,N_16226,N_16459);
nand U16820 (N_16820,N_16332,N_16126);
nand U16821 (N_16821,N_16452,N_16453);
nand U16822 (N_16822,N_16149,N_16262);
and U16823 (N_16823,N_16475,N_16169);
nor U16824 (N_16824,N_16113,N_16138);
nor U16825 (N_16825,N_16370,N_16192);
or U16826 (N_16826,N_16439,N_16443);
xor U16827 (N_16827,N_16108,N_16383);
nor U16828 (N_16828,N_16430,N_16126);
and U16829 (N_16829,N_16016,N_16263);
nand U16830 (N_16830,N_16155,N_16054);
or U16831 (N_16831,N_16355,N_16087);
or U16832 (N_16832,N_16218,N_16128);
nor U16833 (N_16833,N_16306,N_16252);
nand U16834 (N_16834,N_16050,N_16381);
or U16835 (N_16835,N_16236,N_16472);
nand U16836 (N_16836,N_16403,N_16054);
or U16837 (N_16837,N_16354,N_16066);
and U16838 (N_16838,N_16195,N_16399);
or U16839 (N_16839,N_16300,N_16211);
nand U16840 (N_16840,N_16213,N_16482);
nor U16841 (N_16841,N_16357,N_16250);
nor U16842 (N_16842,N_16360,N_16438);
nor U16843 (N_16843,N_16064,N_16146);
and U16844 (N_16844,N_16391,N_16144);
and U16845 (N_16845,N_16383,N_16320);
and U16846 (N_16846,N_16333,N_16344);
or U16847 (N_16847,N_16136,N_16150);
or U16848 (N_16848,N_16454,N_16030);
nor U16849 (N_16849,N_16138,N_16470);
and U16850 (N_16850,N_16324,N_16049);
xor U16851 (N_16851,N_16258,N_16152);
nand U16852 (N_16852,N_16412,N_16316);
nand U16853 (N_16853,N_16012,N_16357);
nor U16854 (N_16854,N_16426,N_16483);
xnor U16855 (N_16855,N_16202,N_16340);
and U16856 (N_16856,N_16266,N_16164);
and U16857 (N_16857,N_16475,N_16362);
nand U16858 (N_16858,N_16322,N_16171);
xor U16859 (N_16859,N_16274,N_16298);
or U16860 (N_16860,N_16144,N_16122);
nor U16861 (N_16861,N_16127,N_16234);
or U16862 (N_16862,N_16027,N_16339);
nor U16863 (N_16863,N_16204,N_16248);
nor U16864 (N_16864,N_16339,N_16377);
or U16865 (N_16865,N_16189,N_16270);
or U16866 (N_16866,N_16269,N_16325);
xnor U16867 (N_16867,N_16235,N_16167);
and U16868 (N_16868,N_16336,N_16373);
xnor U16869 (N_16869,N_16450,N_16228);
or U16870 (N_16870,N_16377,N_16313);
and U16871 (N_16871,N_16422,N_16191);
xnor U16872 (N_16872,N_16139,N_16199);
xor U16873 (N_16873,N_16065,N_16353);
and U16874 (N_16874,N_16454,N_16107);
or U16875 (N_16875,N_16353,N_16082);
or U16876 (N_16876,N_16398,N_16407);
nor U16877 (N_16877,N_16084,N_16233);
xnor U16878 (N_16878,N_16456,N_16438);
nor U16879 (N_16879,N_16181,N_16421);
nor U16880 (N_16880,N_16354,N_16051);
xnor U16881 (N_16881,N_16152,N_16302);
and U16882 (N_16882,N_16005,N_16182);
and U16883 (N_16883,N_16127,N_16029);
xor U16884 (N_16884,N_16281,N_16153);
nand U16885 (N_16885,N_16108,N_16452);
nand U16886 (N_16886,N_16325,N_16087);
or U16887 (N_16887,N_16408,N_16391);
and U16888 (N_16888,N_16188,N_16104);
xnor U16889 (N_16889,N_16144,N_16368);
or U16890 (N_16890,N_16250,N_16418);
or U16891 (N_16891,N_16149,N_16221);
nand U16892 (N_16892,N_16404,N_16411);
nor U16893 (N_16893,N_16291,N_16211);
xnor U16894 (N_16894,N_16314,N_16096);
nor U16895 (N_16895,N_16498,N_16323);
nor U16896 (N_16896,N_16212,N_16499);
nand U16897 (N_16897,N_16053,N_16057);
nand U16898 (N_16898,N_16005,N_16067);
nor U16899 (N_16899,N_16068,N_16358);
nand U16900 (N_16900,N_16213,N_16073);
nor U16901 (N_16901,N_16196,N_16108);
nor U16902 (N_16902,N_16283,N_16055);
nand U16903 (N_16903,N_16043,N_16231);
xnor U16904 (N_16904,N_16128,N_16427);
xnor U16905 (N_16905,N_16174,N_16226);
and U16906 (N_16906,N_16058,N_16433);
nor U16907 (N_16907,N_16292,N_16001);
and U16908 (N_16908,N_16380,N_16374);
and U16909 (N_16909,N_16334,N_16262);
and U16910 (N_16910,N_16135,N_16124);
and U16911 (N_16911,N_16009,N_16048);
nand U16912 (N_16912,N_16079,N_16117);
and U16913 (N_16913,N_16054,N_16318);
and U16914 (N_16914,N_16145,N_16315);
nor U16915 (N_16915,N_16349,N_16299);
xor U16916 (N_16916,N_16439,N_16484);
or U16917 (N_16917,N_16323,N_16468);
xor U16918 (N_16918,N_16268,N_16077);
nor U16919 (N_16919,N_16089,N_16476);
nor U16920 (N_16920,N_16223,N_16341);
and U16921 (N_16921,N_16370,N_16391);
xor U16922 (N_16922,N_16341,N_16398);
xor U16923 (N_16923,N_16248,N_16492);
and U16924 (N_16924,N_16278,N_16023);
nor U16925 (N_16925,N_16038,N_16268);
or U16926 (N_16926,N_16238,N_16087);
and U16927 (N_16927,N_16175,N_16137);
xnor U16928 (N_16928,N_16199,N_16377);
nand U16929 (N_16929,N_16327,N_16268);
and U16930 (N_16930,N_16213,N_16071);
or U16931 (N_16931,N_16095,N_16120);
xor U16932 (N_16932,N_16253,N_16071);
or U16933 (N_16933,N_16370,N_16476);
or U16934 (N_16934,N_16263,N_16141);
nand U16935 (N_16935,N_16226,N_16239);
or U16936 (N_16936,N_16491,N_16133);
nand U16937 (N_16937,N_16397,N_16095);
nor U16938 (N_16938,N_16230,N_16146);
nor U16939 (N_16939,N_16375,N_16247);
nor U16940 (N_16940,N_16303,N_16251);
and U16941 (N_16941,N_16322,N_16435);
nand U16942 (N_16942,N_16241,N_16074);
nand U16943 (N_16943,N_16012,N_16037);
and U16944 (N_16944,N_16128,N_16237);
and U16945 (N_16945,N_16440,N_16014);
xor U16946 (N_16946,N_16015,N_16418);
xnor U16947 (N_16947,N_16135,N_16178);
nor U16948 (N_16948,N_16144,N_16022);
and U16949 (N_16949,N_16490,N_16454);
nand U16950 (N_16950,N_16243,N_16337);
xnor U16951 (N_16951,N_16360,N_16315);
xnor U16952 (N_16952,N_16052,N_16114);
nor U16953 (N_16953,N_16445,N_16299);
nor U16954 (N_16954,N_16454,N_16215);
and U16955 (N_16955,N_16360,N_16405);
nor U16956 (N_16956,N_16166,N_16093);
nand U16957 (N_16957,N_16327,N_16149);
xor U16958 (N_16958,N_16232,N_16242);
or U16959 (N_16959,N_16146,N_16169);
and U16960 (N_16960,N_16358,N_16107);
or U16961 (N_16961,N_16375,N_16174);
nand U16962 (N_16962,N_16326,N_16195);
or U16963 (N_16963,N_16341,N_16327);
nand U16964 (N_16964,N_16061,N_16346);
nor U16965 (N_16965,N_16034,N_16330);
or U16966 (N_16966,N_16132,N_16425);
and U16967 (N_16967,N_16394,N_16224);
and U16968 (N_16968,N_16036,N_16372);
and U16969 (N_16969,N_16068,N_16098);
or U16970 (N_16970,N_16058,N_16022);
and U16971 (N_16971,N_16370,N_16104);
and U16972 (N_16972,N_16432,N_16227);
nor U16973 (N_16973,N_16232,N_16216);
nand U16974 (N_16974,N_16081,N_16498);
nor U16975 (N_16975,N_16099,N_16416);
or U16976 (N_16976,N_16416,N_16232);
nor U16977 (N_16977,N_16003,N_16239);
and U16978 (N_16978,N_16394,N_16175);
or U16979 (N_16979,N_16347,N_16496);
nand U16980 (N_16980,N_16115,N_16221);
xor U16981 (N_16981,N_16463,N_16493);
nor U16982 (N_16982,N_16325,N_16265);
or U16983 (N_16983,N_16136,N_16280);
and U16984 (N_16984,N_16241,N_16472);
and U16985 (N_16985,N_16469,N_16426);
and U16986 (N_16986,N_16237,N_16413);
nand U16987 (N_16987,N_16101,N_16347);
xor U16988 (N_16988,N_16411,N_16482);
xnor U16989 (N_16989,N_16437,N_16436);
xnor U16990 (N_16990,N_16323,N_16049);
or U16991 (N_16991,N_16129,N_16270);
or U16992 (N_16992,N_16277,N_16049);
and U16993 (N_16993,N_16024,N_16058);
or U16994 (N_16994,N_16150,N_16109);
nor U16995 (N_16995,N_16229,N_16340);
and U16996 (N_16996,N_16132,N_16283);
nand U16997 (N_16997,N_16087,N_16193);
nand U16998 (N_16998,N_16440,N_16467);
xnor U16999 (N_16999,N_16256,N_16243);
nor U17000 (N_17000,N_16564,N_16749);
xor U17001 (N_17001,N_16980,N_16981);
nand U17002 (N_17002,N_16839,N_16534);
nand U17003 (N_17003,N_16550,N_16668);
and U17004 (N_17004,N_16714,N_16545);
nor U17005 (N_17005,N_16568,N_16913);
nand U17006 (N_17006,N_16645,N_16625);
nor U17007 (N_17007,N_16755,N_16826);
nor U17008 (N_17008,N_16995,N_16794);
nand U17009 (N_17009,N_16976,N_16522);
and U17010 (N_17010,N_16802,N_16742);
nor U17011 (N_17011,N_16660,N_16946);
nand U17012 (N_17012,N_16528,N_16650);
xor U17013 (N_17013,N_16613,N_16789);
nor U17014 (N_17014,N_16822,N_16731);
or U17015 (N_17015,N_16554,N_16932);
and U17016 (N_17016,N_16724,N_16923);
xnor U17017 (N_17017,N_16898,N_16697);
xor U17018 (N_17018,N_16865,N_16909);
xor U17019 (N_17019,N_16986,N_16639);
and U17020 (N_17020,N_16730,N_16886);
xor U17021 (N_17021,N_16566,N_16585);
or U17022 (N_17022,N_16633,N_16962);
nor U17023 (N_17023,N_16837,N_16655);
nor U17024 (N_17024,N_16838,N_16996);
xor U17025 (N_17025,N_16988,N_16944);
xnor U17026 (N_17026,N_16868,N_16629);
or U17027 (N_17027,N_16748,N_16906);
xnor U17028 (N_17028,N_16505,N_16860);
xnor U17029 (N_17029,N_16567,N_16542);
or U17030 (N_17030,N_16527,N_16921);
nor U17031 (N_17031,N_16611,N_16649);
nand U17032 (N_17032,N_16713,N_16679);
and U17033 (N_17033,N_16694,N_16676);
or U17034 (N_17034,N_16840,N_16992);
xor U17035 (N_17035,N_16561,N_16752);
nor U17036 (N_17036,N_16523,N_16994);
nand U17037 (N_17037,N_16776,N_16610);
and U17038 (N_17038,N_16983,N_16847);
and U17039 (N_17039,N_16654,N_16594);
nand U17040 (N_17040,N_16916,N_16619);
xnor U17041 (N_17041,N_16695,N_16598);
xor U17042 (N_17042,N_16774,N_16772);
and U17043 (N_17043,N_16907,N_16854);
xor U17044 (N_17044,N_16795,N_16973);
and U17045 (N_17045,N_16663,N_16920);
or U17046 (N_17046,N_16581,N_16940);
and U17047 (N_17047,N_16929,N_16969);
or U17048 (N_17048,N_16778,N_16669);
or U17049 (N_17049,N_16721,N_16693);
xor U17050 (N_17050,N_16606,N_16856);
nand U17051 (N_17051,N_16820,N_16869);
xor U17052 (N_17052,N_16905,N_16600);
nor U17053 (N_17053,N_16716,N_16531);
nand U17054 (N_17054,N_16555,N_16915);
xnor U17055 (N_17055,N_16756,N_16873);
nor U17056 (N_17056,N_16703,N_16551);
or U17057 (N_17057,N_16532,N_16931);
or U17058 (N_17058,N_16546,N_16958);
nand U17059 (N_17059,N_16949,N_16674);
xor U17060 (N_17060,N_16991,N_16684);
or U17061 (N_17061,N_16500,N_16956);
or U17062 (N_17062,N_16979,N_16841);
or U17063 (N_17063,N_16975,N_16572);
nand U17064 (N_17064,N_16569,N_16623);
nor U17065 (N_17065,N_16607,N_16705);
xor U17066 (N_17066,N_16615,N_16535);
xor U17067 (N_17067,N_16894,N_16603);
or U17068 (N_17068,N_16720,N_16521);
nor U17069 (N_17069,N_16799,N_16953);
xnor U17070 (N_17070,N_16770,N_16791);
nor U17071 (N_17071,N_16543,N_16595);
or U17072 (N_17072,N_16876,N_16782);
nand U17073 (N_17073,N_16833,N_16656);
xor U17074 (N_17074,N_16671,N_16638);
nand U17075 (N_17075,N_16788,N_16941);
xor U17076 (N_17076,N_16664,N_16836);
or U17077 (N_17077,N_16883,N_16516);
and U17078 (N_17078,N_16939,N_16616);
or U17079 (N_17079,N_16580,N_16754);
nand U17080 (N_17080,N_16675,N_16634);
xnor U17081 (N_17081,N_16851,N_16766);
and U17082 (N_17082,N_16740,N_16628);
or U17083 (N_17083,N_16790,N_16526);
and U17084 (N_17084,N_16525,N_16970);
and U17085 (N_17085,N_16942,N_16702);
and U17086 (N_17086,N_16768,N_16621);
and U17087 (N_17087,N_16578,N_16746);
and U17088 (N_17088,N_16699,N_16759);
and U17089 (N_17089,N_16582,N_16643);
or U17090 (N_17090,N_16723,N_16848);
and U17091 (N_17091,N_16618,N_16771);
nand U17092 (N_17092,N_16733,N_16914);
nor U17093 (N_17093,N_16514,N_16792);
nand U17094 (N_17094,N_16753,N_16509);
nor U17095 (N_17095,N_16903,N_16692);
or U17096 (N_17096,N_16571,N_16640);
nor U17097 (N_17097,N_16875,N_16821);
or U17098 (N_17098,N_16857,N_16548);
nand U17099 (N_17099,N_16503,N_16574);
or U17100 (N_17100,N_16501,N_16943);
nand U17101 (N_17101,N_16646,N_16573);
and U17102 (N_17102,N_16722,N_16597);
and U17103 (N_17103,N_16965,N_16729);
nor U17104 (N_17104,N_16918,N_16818);
or U17105 (N_17105,N_16718,N_16626);
and U17106 (N_17106,N_16957,N_16565);
nand U17107 (N_17107,N_16747,N_16576);
or U17108 (N_17108,N_16579,N_16644);
nand U17109 (N_17109,N_16517,N_16888);
or U17110 (N_17110,N_16924,N_16866);
or U17111 (N_17111,N_16937,N_16651);
nand U17112 (N_17112,N_16558,N_16895);
nor U17113 (N_17113,N_16672,N_16709);
nor U17114 (N_17114,N_16764,N_16850);
or U17115 (N_17115,N_16617,N_16959);
or U17116 (N_17116,N_16605,N_16925);
nand U17117 (N_17117,N_16659,N_16648);
xnor U17118 (N_17118,N_16596,N_16750);
or U17119 (N_17119,N_16910,N_16736);
or U17120 (N_17120,N_16584,N_16877);
and U17121 (N_17121,N_16963,N_16817);
nor U17122 (N_17122,N_16518,N_16711);
or U17123 (N_17123,N_16891,N_16536);
nand U17124 (N_17124,N_16867,N_16950);
xnor U17125 (N_17125,N_16680,N_16701);
xnor U17126 (N_17126,N_16880,N_16588);
nor U17127 (N_17127,N_16948,N_16859);
nor U17128 (N_17128,N_16508,N_16583);
nor U17129 (N_17129,N_16539,N_16512);
xnor U17130 (N_17130,N_16696,N_16902);
xor U17131 (N_17131,N_16874,N_16870);
xor U17132 (N_17132,N_16652,N_16587);
or U17133 (N_17133,N_16919,N_16801);
and U17134 (N_17134,N_16636,N_16624);
and U17135 (N_17135,N_16667,N_16954);
xnor U17136 (N_17136,N_16544,N_16602);
or U17137 (N_17137,N_16922,N_16520);
nand U17138 (N_17138,N_16717,N_16510);
nand U17139 (N_17139,N_16642,N_16912);
or U17140 (N_17140,N_16599,N_16845);
and U17141 (N_17141,N_16832,N_16974);
xnor U17142 (N_17142,N_16879,N_16515);
and U17143 (N_17143,N_16783,N_16775);
nand U17144 (N_17144,N_16786,N_16890);
and U17145 (N_17145,N_16553,N_16745);
and U17146 (N_17146,N_16834,N_16966);
nor U17147 (N_17147,N_16604,N_16538);
nor U17148 (N_17148,N_16908,N_16726);
or U17149 (N_17149,N_16853,N_16989);
and U17150 (N_17150,N_16777,N_16530);
or U17151 (N_17151,N_16997,N_16686);
nor U17152 (N_17152,N_16627,N_16511);
or U17153 (N_17153,N_16631,N_16519);
nor U17154 (N_17154,N_16805,N_16936);
nor U17155 (N_17155,N_16739,N_16899);
xnor U17156 (N_17156,N_16773,N_16813);
and U17157 (N_17157,N_16592,N_16562);
nor U17158 (N_17158,N_16762,N_16765);
nand U17159 (N_17159,N_16661,N_16691);
and U17160 (N_17160,N_16677,N_16767);
xnor U17161 (N_17161,N_16964,N_16938);
nand U17162 (N_17162,N_16549,N_16999);
xnor U17163 (N_17163,N_16590,N_16779);
nand U17164 (N_17164,N_16635,N_16657);
or U17165 (N_17165,N_16904,N_16968);
or U17166 (N_17166,N_16985,N_16798);
nand U17167 (N_17167,N_16557,N_16810);
or U17168 (N_17168,N_16710,N_16926);
or U17169 (N_17169,N_16612,N_16744);
or U17170 (N_17170,N_16814,N_16653);
xor U17171 (N_17171,N_16559,N_16601);
nand U17172 (N_17172,N_16529,N_16537);
and U17173 (N_17173,N_16758,N_16734);
xnor U17174 (N_17174,N_16825,N_16751);
and U17175 (N_17175,N_16727,N_16743);
nor U17176 (N_17176,N_16785,N_16872);
xnor U17177 (N_17177,N_16998,N_16861);
xnor U17178 (N_17178,N_16698,N_16900);
xor U17179 (N_17179,N_16708,N_16620);
or U17180 (N_17180,N_16560,N_16862);
nor U17181 (N_17181,N_16960,N_16945);
nand U17182 (N_17182,N_16984,N_16881);
and U17183 (N_17183,N_16556,N_16547);
xnor U17184 (N_17184,N_16673,N_16893);
xor U17185 (N_17185,N_16715,N_16885);
nor U17186 (N_17186,N_16808,N_16504);
and U17187 (N_17187,N_16884,N_16570);
xnor U17188 (N_17188,N_16678,N_16804);
xor U17189 (N_17189,N_16670,N_16955);
xnor U17190 (N_17190,N_16760,N_16972);
nor U17191 (N_17191,N_16816,N_16577);
nor U17192 (N_17192,N_16593,N_16683);
or U17193 (N_17193,N_16971,N_16982);
nand U17194 (N_17194,N_16533,N_16608);
or U17195 (N_17195,N_16685,N_16990);
xnor U17196 (N_17196,N_16892,N_16889);
and U17197 (N_17197,N_16911,N_16540);
and U17198 (N_17198,N_16882,N_16704);
nor U17199 (N_17199,N_16793,N_16666);
and U17200 (N_17200,N_16700,N_16846);
xor U17201 (N_17201,N_16689,N_16812);
or U17202 (N_17202,N_16707,N_16961);
nor U17203 (N_17203,N_16513,N_16896);
nor U17204 (N_17204,N_16614,N_16632);
and U17205 (N_17205,N_16586,N_16687);
xnor U17206 (N_17206,N_16637,N_16927);
nor U17207 (N_17207,N_16987,N_16763);
nand U17208 (N_17208,N_16849,N_16738);
nor U17209 (N_17209,N_16829,N_16855);
nand U17210 (N_17210,N_16928,N_16807);
xor U17211 (N_17211,N_16591,N_16863);
and U17212 (N_17212,N_16934,N_16552);
or U17213 (N_17213,N_16658,N_16780);
or U17214 (N_17214,N_16524,N_16978);
and U17215 (N_17215,N_16815,N_16728);
or U17216 (N_17216,N_16630,N_16622);
xor U17217 (N_17217,N_16800,N_16641);
nor U17218 (N_17218,N_16933,N_16796);
and U17219 (N_17219,N_16811,N_16947);
and U17220 (N_17220,N_16977,N_16741);
nor U17221 (N_17221,N_16831,N_16507);
xnor U17222 (N_17222,N_16842,N_16828);
and U17223 (N_17223,N_16784,N_16662);
and U17224 (N_17224,N_16806,N_16835);
xor U17225 (N_17225,N_16952,N_16609);
nor U17226 (N_17226,N_16563,N_16732);
nor U17227 (N_17227,N_16901,N_16823);
xor U17228 (N_17228,N_16819,N_16706);
and U17229 (N_17229,N_16712,N_16682);
nor U17230 (N_17230,N_16993,N_16852);
or U17231 (N_17231,N_16735,N_16502);
or U17232 (N_17232,N_16844,N_16647);
xnor U17233 (N_17233,N_16864,N_16809);
and U17234 (N_17234,N_16757,N_16930);
and U17235 (N_17235,N_16843,N_16897);
nand U17236 (N_17236,N_16737,N_16917);
nor U17237 (N_17237,N_16589,N_16878);
xnor U17238 (N_17238,N_16830,N_16803);
xnor U17239 (N_17239,N_16824,N_16871);
nand U17240 (N_17240,N_16935,N_16688);
nor U17241 (N_17241,N_16725,N_16951);
xnor U17242 (N_17242,N_16575,N_16681);
or U17243 (N_17243,N_16827,N_16781);
or U17244 (N_17244,N_16967,N_16797);
or U17245 (N_17245,N_16506,N_16719);
and U17246 (N_17246,N_16665,N_16887);
and U17247 (N_17247,N_16769,N_16858);
or U17248 (N_17248,N_16787,N_16690);
and U17249 (N_17249,N_16541,N_16761);
nand U17250 (N_17250,N_16705,N_16755);
nand U17251 (N_17251,N_16646,N_16519);
nor U17252 (N_17252,N_16513,N_16963);
xnor U17253 (N_17253,N_16965,N_16749);
or U17254 (N_17254,N_16756,N_16957);
nor U17255 (N_17255,N_16733,N_16957);
nand U17256 (N_17256,N_16961,N_16728);
xnor U17257 (N_17257,N_16894,N_16758);
nand U17258 (N_17258,N_16519,N_16883);
nand U17259 (N_17259,N_16707,N_16879);
xor U17260 (N_17260,N_16569,N_16980);
and U17261 (N_17261,N_16688,N_16585);
nor U17262 (N_17262,N_16973,N_16658);
nor U17263 (N_17263,N_16985,N_16969);
or U17264 (N_17264,N_16678,N_16906);
or U17265 (N_17265,N_16943,N_16736);
xor U17266 (N_17266,N_16899,N_16702);
and U17267 (N_17267,N_16932,N_16912);
and U17268 (N_17268,N_16618,N_16817);
nor U17269 (N_17269,N_16854,N_16786);
or U17270 (N_17270,N_16757,N_16784);
xnor U17271 (N_17271,N_16516,N_16814);
xnor U17272 (N_17272,N_16796,N_16750);
nand U17273 (N_17273,N_16538,N_16963);
or U17274 (N_17274,N_16818,N_16863);
and U17275 (N_17275,N_16531,N_16876);
xor U17276 (N_17276,N_16678,N_16781);
and U17277 (N_17277,N_16782,N_16964);
xnor U17278 (N_17278,N_16932,N_16705);
nand U17279 (N_17279,N_16712,N_16794);
or U17280 (N_17280,N_16652,N_16933);
and U17281 (N_17281,N_16839,N_16735);
xnor U17282 (N_17282,N_16844,N_16926);
xnor U17283 (N_17283,N_16893,N_16539);
nor U17284 (N_17284,N_16583,N_16847);
xor U17285 (N_17285,N_16715,N_16600);
nand U17286 (N_17286,N_16990,N_16957);
and U17287 (N_17287,N_16965,N_16994);
or U17288 (N_17288,N_16801,N_16618);
nand U17289 (N_17289,N_16507,N_16943);
nand U17290 (N_17290,N_16999,N_16796);
nand U17291 (N_17291,N_16777,N_16774);
nor U17292 (N_17292,N_16969,N_16609);
and U17293 (N_17293,N_16888,N_16817);
xnor U17294 (N_17294,N_16877,N_16750);
or U17295 (N_17295,N_16716,N_16506);
nor U17296 (N_17296,N_16786,N_16954);
xor U17297 (N_17297,N_16973,N_16695);
nor U17298 (N_17298,N_16990,N_16900);
xnor U17299 (N_17299,N_16744,N_16559);
nand U17300 (N_17300,N_16821,N_16927);
nand U17301 (N_17301,N_16510,N_16997);
nor U17302 (N_17302,N_16996,N_16910);
and U17303 (N_17303,N_16886,N_16865);
and U17304 (N_17304,N_16569,N_16901);
or U17305 (N_17305,N_16579,N_16774);
and U17306 (N_17306,N_16998,N_16595);
and U17307 (N_17307,N_16509,N_16747);
or U17308 (N_17308,N_16915,N_16733);
nor U17309 (N_17309,N_16910,N_16971);
nand U17310 (N_17310,N_16892,N_16609);
and U17311 (N_17311,N_16788,N_16961);
nor U17312 (N_17312,N_16769,N_16533);
or U17313 (N_17313,N_16907,N_16934);
nand U17314 (N_17314,N_16981,N_16690);
nand U17315 (N_17315,N_16999,N_16940);
and U17316 (N_17316,N_16623,N_16638);
nor U17317 (N_17317,N_16788,N_16946);
or U17318 (N_17318,N_16803,N_16861);
nor U17319 (N_17319,N_16965,N_16912);
or U17320 (N_17320,N_16922,N_16804);
or U17321 (N_17321,N_16849,N_16532);
nand U17322 (N_17322,N_16968,N_16927);
or U17323 (N_17323,N_16557,N_16566);
or U17324 (N_17324,N_16941,N_16927);
nor U17325 (N_17325,N_16505,N_16589);
xnor U17326 (N_17326,N_16540,N_16527);
and U17327 (N_17327,N_16698,N_16949);
and U17328 (N_17328,N_16743,N_16665);
and U17329 (N_17329,N_16682,N_16978);
nand U17330 (N_17330,N_16671,N_16526);
nor U17331 (N_17331,N_16675,N_16878);
nor U17332 (N_17332,N_16817,N_16941);
xnor U17333 (N_17333,N_16726,N_16552);
or U17334 (N_17334,N_16960,N_16662);
xor U17335 (N_17335,N_16875,N_16678);
nand U17336 (N_17336,N_16646,N_16704);
nand U17337 (N_17337,N_16883,N_16604);
nor U17338 (N_17338,N_16879,N_16560);
or U17339 (N_17339,N_16942,N_16884);
xnor U17340 (N_17340,N_16691,N_16787);
or U17341 (N_17341,N_16620,N_16635);
xnor U17342 (N_17342,N_16992,N_16860);
nor U17343 (N_17343,N_16656,N_16642);
and U17344 (N_17344,N_16547,N_16954);
or U17345 (N_17345,N_16603,N_16663);
or U17346 (N_17346,N_16652,N_16577);
nor U17347 (N_17347,N_16570,N_16772);
or U17348 (N_17348,N_16907,N_16747);
xor U17349 (N_17349,N_16981,N_16889);
nand U17350 (N_17350,N_16555,N_16646);
xnor U17351 (N_17351,N_16878,N_16511);
nand U17352 (N_17352,N_16813,N_16895);
nor U17353 (N_17353,N_16654,N_16970);
nor U17354 (N_17354,N_16667,N_16679);
and U17355 (N_17355,N_16618,N_16831);
or U17356 (N_17356,N_16504,N_16564);
and U17357 (N_17357,N_16626,N_16711);
nand U17358 (N_17358,N_16912,N_16542);
and U17359 (N_17359,N_16510,N_16519);
and U17360 (N_17360,N_16677,N_16515);
xor U17361 (N_17361,N_16645,N_16962);
nand U17362 (N_17362,N_16696,N_16606);
xnor U17363 (N_17363,N_16771,N_16648);
nor U17364 (N_17364,N_16683,N_16882);
or U17365 (N_17365,N_16515,N_16800);
xnor U17366 (N_17366,N_16903,N_16623);
nor U17367 (N_17367,N_16649,N_16701);
and U17368 (N_17368,N_16653,N_16661);
nor U17369 (N_17369,N_16988,N_16858);
or U17370 (N_17370,N_16527,N_16618);
or U17371 (N_17371,N_16512,N_16716);
or U17372 (N_17372,N_16582,N_16509);
and U17373 (N_17373,N_16658,N_16737);
nand U17374 (N_17374,N_16808,N_16684);
nor U17375 (N_17375,N_16629,N_16636);
nor U17376 (N_17376,N_16502,N_16829);
nor U17377 (N_17377,N_16980,N_16667);
or U17378 (N_17378,N_16807,N_16755);
or U17379 (N_17379,N_16946,N_16641);
nor U17380 (N_17380,N_16847,N_16705);
or U17381 (N_17381,N_16525,N_16754);
or U17382 (N_17382,N_16659,N_16854);
or U17383 (N_17383,N_16863,N_16858);
or U17384 (N_17384,N_16678,N_16571);
xnor U17385 (N_17385,N_16681,N_16973);
xnor U17386 (N_17386,N_16967,N_16643);
xnor U17387 (N_17387,N_16668,N_16720);
or U17388 (N_17388,N_16680,N_16885);
or U17389 (N_17389,N_16698,N_16667);
nor U17390 (N_17390,N_16681,N_16844);
and U17391 (N_17391,N_16505,N_16889);
nor U17392 (N_17392,N_16641,N_16728);
or U17393 (N_17393,N_16918,N_16644);
and U17394 (N_17394,N_16764,N_16735);
nand U17395 (N_17395,N_16829,N_16651);
nor U17396 (N_17396,N_16921,N_16916);
xnor U17397 (N_17397,N_16535,N_16894);
and U17398 (N_17398,N_16697,N_16961);
nor U17399 (N_17399,N_16839,N_16640);
nand U17400 (N_17400,N_16592,N_16838);
nor U17401 (N_17401,N_16573,N_16788);
nand U17402 (N_17402,N_16944,N_16940);
xor U17403 (N_17403,N_16650,N_16768);
and U17404 (N_17404,N_16576,N_16648);
nor U17405 (N_17405,N_16501,N_16739);
nand U17406 (N_17406,N_16623,N_16515);
nand U17407 (N_17407,N_16955,N_16900);
nand U17408 (N_17408,N_16914,N_16853);
nor U17409 (N_17409,N_16771,N_16803);
and U17410 (N_17410,N_16672,N_16928);
or U17411 (N_17411,N_16548,N_16865);
or U17412 (N_17412,N_16803,N_16825);
and U17413 (N_17413,N_16720,N_16555);
xnor U17414 (N_17414,N_16724,N_16863);
and U17415 (N_17415,N_16574,N_16680);
nand U17416 (N_17416,N_16712,N_16963);
nand U17417 (N_17417,N_16923,N_16559);
nor U17418 (N_17418,N_16970,N_16537);
or U17419 (N_17419,N_16691,N_16634);
xnor U17420 (N_17420,N_16603,N_16858);
nor U17421 (N_17421,N_16842,N_16682);
xnor U17422 (N_17422,N_16599,N_16941);
xor U17423 (N_17423,N_16613,N_16866);
or U17424 (N_17424,N_16517,N_16526);
nand U17425 (N_17425,N_16642,N_16898);
nor U17426 (N_17426,N_16905,N_16781);
or U17427 (N_17427,N_16918,N_16536);
and U17428 (N_17428,N_16931,N_16652);
and U17429 (N_17429,N_16946,N_16583);
or U17430 (N_17430,N_16579,N_16726);
nand U17431 (N_17431,N_16918,N_16580);
xnor U17432 (N_17432,N_16931,N_16511);
xor U17433 (N_17433,N_16730,N_16789);
xnor U17434 (N_17434,N_16806,N_16520);
and U17435 (N_17435,N_16954,N_16683);
and U17436 (N_17436,N_16999,N_16971);
nor U17437 (N_17437,N_16780,N_16576);
nand U17438 (N_17438,N_16739,N_16875);
or U17439 (N_17439,N_16919,N_16986);
nand U17440 (N_17440,N_16761,N_16571);
nor U17441 (N_17441,N_16584,N_16959);
nor U17442 (N_17442,N_16987,N_16909);
xor U17443 (N_17443,N_16640,N_16975);
nand U17444 (N_17444,N_16798,N_16955);
and U17445 (N_17445,N_16654,N_16531);
nor U17446 (N_17446,N_16900,N_16883);
nor U17447 (N_17447,N_16759,N_16664);
or U17448 (N_17448,N_16703,N_16726);
or U17449 (N_17449,N_16943,N_16921);
nor U17450 (N_17450,N_16541,N_16938);
and U17451 (N_17451,N_16731,N_16938);
nand U17452 (N_17452,N_16964,N_16933);
nand U17453 (N_17453,N_16797,N_16773);
nand U17454 (N_17454,N_16768,N_16769);
xnor U17455 (N_17455,N_16747,N_16952);
nor U17456 (N_17456,N_16727,N_16813);
nor U17457 (N_17457,N_16934,N_16748);
xnor U17458 (N_17458,N_16508,N_16589);
nor U17459 (N_17459,N_16585,N_16842);
xor U17460 (N_17460,N_16720,N_16918);
xnor U17461 (N_17461,N_16903,N_16775);
xnor U17462 (N_17462,N_16812,N_16664);
and U17463 (N_17463,N_16541,N_16538);
nor U17464 (N_17464,N_16768,N_16631);
and U17465 (N_17465,N_16992,N_16766);
nor U17466 (N_17466,N_16984,N_16528);
nand U17467 (N_17467,N_16758,N_16600);
xnor U17468 (N_17468,N_16867,N_16652);
xnor U17469 (N_17469,N_16678,N_16726);
and U17470 (N_17470,N_16504,N_16571);
nor U17471 (N_17471,N_16546,N_16967);
and U17472 (N_17472,N_16942,N_16891);
nand U17473 (N_17473,N_16874,N_16858);
xor U17474 (N_17474,N_16860,N_16696);
xnor U17475 (N_17475,N_16537,N_16603);
nand U17476 (N_17476,N_16994,N_16593);
xnor U17477 (N_17477,N_16632,N_16629);
nand U17478 (N_17478,N_16966,N_16551);
and U17479 (N_17479,N_16685,N_16775);
nor U17480 (N_17480,N_16565,N_16904);
and U17481 (N_17481,N_16673,N_16628);
or U17482 (N_17482,N_16725,N_16826);
or U17483 (N_17483,N_16886,N_16821);
or U17484 (N_17484,N_16884,N_16933);
nor U17485 (N_17485,N_16917,N_16631);
or U17486 (N_17486,N_16933,N_16597);
or U17487 (N_17487,N_16822,N_16775);
and U17488 (N_17488,N_16822,N_16864);
nand U17489 (N_17489,N_16904,N_16570);
xnor U17490 (N_17490,N_16820,N_16847);
or U17491 (N_17491,N_16803,N_16823);
xor U17492 (N_17492,N_16827,N_16815);
nand U17493 (N_17493,N_16731,N_16593);
or U17494 (N_17494,N_16974,N_16947);
nor U17495 (N_17495,N_16821,N_16972);
nand U17496 (N_17496,N_16669,N_16588);
and U17497 (N_17497,N_16557,N_16706);
or U17498 (N_17498,N_16528,N_16772);
or U17499 (N_17499,N_16881,N_16884);
and U17500 (N_17500,N_17325,N_17005);
nor U17501 (N_17501,N_17057,N_17191);
or U17502 (N_17502,N_17400,N_17226);
and U17503 (N_17503,N_17468,N_17122);
or U17504 (N_17504,N_17270,N_17124);
xnor U17505 (N_17505,N_17352,N_17008);
xnor U17506 (N_17506,N_17004,N_17131);
and U17507 (N_17507,N_17480,N_17207);
xnor U17508 (N_17508,N_17332,N_17200);
nor U17509 (N_17509,N_17446,N_17474);
nor U17510 (N_17510,N_17157,N_17436);
nor U17511 (N_17511,N_17060,N_17299);
or U17512 (N_17512,N_17054,N_17027);
or U17513 (N_17513,N_17222,N_17215);
nand U17514 (N_17514,N_17264,N_17421);
or U17515 (N_17515,N_17162,N_17477);
nor U17516 (N_17516,N_17263,N_17188);
xor U17517 (N_17517,N_17497,N_17425);
or U17518 (N_17518,N_17078,N_17063);
nor U17519 (N_17519,N_17096,N_17174);
nand U17520 (N_17520,N_17383,N_17149);
and U17521 (N_17521,N_17449,N_17311);
nor U17522 (N_17522,N_17429,N_17259);
xnor U17523 (N_17523,N_17353,N_17238);
and U17524 (N_17524,N_17049,N_17143);
nor U17525 (N_17525,N_17064,N_17164);
nand U17526 (N_17526,N_17062,N_17097);
and U17527 (N_17527,N_17252,N_17462);
nor U17528 (N_17528,N_17028,N_17220);
nor U17529 (N_17529,N_17190,N_17165);
and U17530 (N_17530,N_17022,N_17184);
nor U17531 (N_17531,N_17050,N_17209);
xnor U17532 (N_17532,N_17350,N_17065);
nand U17533 (N_17533,N_17388,N_17414);
xor U17534 (N_17534,N_17245,N_17045);
and U17535 (N_17535,N_17267,N_17137);
or U17536 (N_17536,N_17309,N_17125);
nor U17537 (N_17537,N_17253,N_17128);
or U17538 (N_17538,N_17195,N_17248);
nor U17539 (N_17539,N_17290,N_17335);
nand U17540 (N_17540,N_17379,N_17079);
and U17541 (N_17541,N_17043,N_17151);
xor U17542 (N_17542,N_17108,N_17336);
xor U17543 (N_17543,N_17288,N_17442);
xor U17544 (N_17544,N_17339,N_17265);
and U17545 (N_17545,N_17107,N_17189);
nand U17546 (N_17546,N_17070,N_17167);
xnor U17547 (N_17547,N_17275,N_17213);
nor U17548 (N_17548,N_17452,N_17084);
nand U17549 (N_17549,N_17235,N_17103);
nor U17550 (N_17550,N_17496,N_17201);
nor U17551 (N_17551,N_17431,N_17277);
nor U17552 (N_17552,N_17306,N_17115);
xnor U17553 (N_17553,N_17021,N_17334);
nand U17554 (N_17554,N_17327,N_17397);
or U17555 (N_17555,N_17017,N_17173);
nor U17556 (N_17556,N_17071,N_17016);
nor U17557 (N_17557,N_17059,N_17111);
or U17558 (N_17558,N_17202,N_17438);
nand U17559 (N_17559,N_17374,N_17018);
and U17560 (N_17560,N_17198,N_17182);
and U17561 (N_17561,N_17396,N_17150);
or U17562 (N_17562,N_17185,N_17241);
xnor U17563 (N_17563,N_17328,N_17029);
xnor U17564 (N_17564,N_17444,N_17205);
nor U17565 (N_17565,N_17003,N_17142);
nand U17566 (N_17566,N_17460,N_17410);
and U17567 (N_17567,N_17356,N_17344);
and U17568 (N_17568,N_17331,N_17192);
nor U17569 (N_17569,N_17387,N_17395);
nand U17570 (N_17570,N_17113,N_17038);
xnor U17571 (N_17571,N_17116,N_17092);
xor U17572 (N_17572,N_17242,N_17489);
nand U17573 (N_17573,N_17441,N_17146);
or U17574 (N_17574,N_17469,N_17066);
nand U17575 (N_17575,N_17020,N_17011);
nor U17576 (N_17576,N_17394,N_17268);
nor U17577 (N_17577,N_17280,N_17240);
nand U17578 (N_17578,N_17037,N_17133);
and U17579 (N_17579,N_17316,N_17117);
nor U17580 (N_17580,N_17281,N_17168);
nor U17581 (N_17581,N_17010,N_17406);
and U17582 (N_17582,N_17499,N_17294);
xor U17583 (N_17583,N_17181,N_17451);
nor U17584 (N_17584,N_17109,N_17119);
xor U17585 (N_17585,N_17278,N_17312);
and U17586 (N_17586,N_17219,N_17361);
xnor U17587 (N_17587,N_17076,N_17083);
or U17588 (N_17588,N_17372,N_17177);
or U17589 (N_17589,N_17385,N_17030);
nor U17590 (N_17590,N_17292,N_17284);
or U17591 (N_17591,N_17376,N_17329);
nor U17592 (N_17592,N_17208,N_17392);
or U17593 (N_17593,N_17416,N_17286);
and U17594 (N_17594,N_17405,N_17251);
xor U17595 (N_17595,N_17390,N_17368);
nand U17596 (N_17596,N_17269,N_17106);
xor U17597 (N_17597,N_17461,N_17206);
xnor U17598 (N_17598,N_17169,N_17012);
or U17599 (N_17599,N_17166,N_17424);
nor U17600 (N_17600,N_17129,N_17458);
xor U17601 (N_17601,N_17330,N_17378);
nor U17602 (N_17602,N_17310,N_17061);
xor U17603 (N_17603,N_17360,N_17298);
xor U17604 (N_17604,N_17254,N_17357);
nand U17605 (N_17605,N_17145,N_17450);
xor U17606 (N_17606,N_17479,N_17121);
or U17607 (N_17607,N_17110,N_17464);
nor U17608 (N_17608,N_17423,N_17171);
nor U17609 (N_17609,N_17428,N_17340);
or U17610 (N_17610,N_17417,N_17026);
nand U17611 (N_17611,N_17052,N_17123);
and U17612 (N_17612,N_17307,N_17354);
nand U17613 (N_17613,N_17419,N_17488);
and U17614 (N_17614,N_17345,N_17170);
nor U17615 (N_17615,N_17302,N_17212);
xor U17616 (N_17616,N_17250,N_17224);
nand U17617 (N_17617,N_17322,N_17147);
nand U17618 (N_17618,N_17039,N_17313);
xnor U17619 (N_17619,N_17051,N_17276);
nand U17620 (N_17620,N_17285,N_17471);
nand U17621 (N_17621,N_17384,N_17291);
xnor U17622 (N_17622,N_17087,N_17440);
or U17623 (N_17623,N_17478,N_17454);
nand U17624 (N_17624,N_17303,N_17093);
xnor U17625 (N_17625,N_17034,N_17375);
nor U17626 (N_17626,N_17035,N_17366);
xnor U17627 (N_17627,N_17148,N_17118);
xnor U17628 (N_17628,N_17348,N_17413);
xor U17629 (N_17629,N_17033,N_17056);
nor U17630 (N_17630,N_17230,N_17180);
or U17631 (N_17631,N_17132,N_17160);
xnor U17632 (N_17632,N_17176,N_17415);
nand U17633 (N_17633,N_17472,N_17355);
xnor U17634 (N_17634,N_17435,N_17102);
or U17635 (N_17635,N_17492,N_17154);
nand U17636 (N_17636,N_17426,N_17156);
xnor U17637 (N_17637,N_17046,N_17297);
and U17638 (N_17638,N_17247,N_17323);
nor U17639 (N_17639,N_17490,N_17283);
nand U17640 (N_17640,N_17495,N_17272);
and U17641 (N_17641,N_17006,N_17483);
or U17642 (N_17642,N_17377,N_17282);
nand U17643 (N_17643,N_17347,N_17214);
and U17644 (N_17644,N_17439,N_17369);
xnor U17645 (N_17645,N_17326,N_17465);
or U17646 (N_17646,N_17130,N_17058);
nand U17647 (N_17647,N_17024,N_17105);
nand U17648 (N_17648,N_17042,N_17085);
nand U17649 (N_17649,N_17186,N_17304);
or U17650 (N_17650,N_17258,N_17041);
xnor U17651 (N_17651,N_17373,N_17262);
and U17652 (N_17652,N_17138,N_17342);
or U17653 (N_17653,N_17141,N_17048);
nand U17654 (N_17654,N_17089,N_17470);
nand U17655 (N_17655,N_17221,N_17296);
or U17656 (N_17656,N_17074,N_17420);
nor U17657 (N_17657,N_17199,N_17475);
nand U17658 (N_17658,N_17203,N_17144);
xnor U17659 (N_17659,N_17498,N_17434);
or U17660 (N_17660,N_17257,N_17244);
nand U17661 (N_17661,N_17314,N_17239);
and U17662 (N_17662,N_17112,N_17104);
nor U17663 (N_17663,N_17289,N_17365);
nand U17664 (N_17664,N_17467,N_17216);
xor U17665 (N_17665,N_17364,N_17228);
and U17666 (N_17666,N_17408,N_17009);
nand U17667 (N_17667,N_17370,N_17000);
and U17668 (N_17668,N_17140,N_17305);
or U17669 (N_17669,N_17015,N_17163);
nor U17670 (N_17670,N_17196,N_17236);
or U17671 (N_17671,N_17274,N_17249);
nand U17672 (N_17672,N_17204,N_17362);
nor U17673 (N_17673,N_17134,N_17403);
nand U17674 (N_17674,N_17098,N_17227);
or U17675 (N_17675,N_17437,N_17308);
nor U17676 (N_17676,N_17175,N_17430);
or U17677 (N_17677,N_17422,N_17100);
and U17678 (N_17678,N_17178,N_17381);
or U17679 (N_17679,N_17346,N_17073);
xor U17680 (N_17680,N_17371,N_17491);
and U17681 (N_17681,N_17023,N_17032);
or U17682 (N_17682,N_17359,N_17279);
nand U17683 (N_17683,N_17389,N_17126);
nor U17684 (N_17684,N_17179,N_17402);
xor U17685 (N_17685,N_17445,N_17211);
or U17686 (N_17686,N_17187,N_17466);
nand U17687 (N_17687,N_17094,N_17481);
and U17688 (N_17688,N_17153,N_17159);
nand U17689 (N_17689,N_17067,N_17194);
or U17690 (N_17690,N_17273,N_17114);
xnor U17691 (N_17691,N_17321,N_17493);
or U17692 (N_17692,N_17231,N_17161);
and U17693 (N_17693,N_17072,N_17456);
or U17694 (N_17694,N_17139,N_17287);
nor U17695 (N_17695,N_17455,N_17031);
or U17696 (N_17696,N_17300,N_17463);
nor U17697 (N_17697,N_17324,N_17301);
xor U17698 (N_17698,N_17053,N_17136);
or U17699 (N_17699,N_17399,N_17197);
and U17700 (N_17700,N_17320,N_17295);
and U17701 (N_17701,N_17081,N_17338);
nand U17702 (N_17702,N_17082,N_17077);
nand U17703 (N_17703,N_17343,N_17172);
xnor U17704 (N_17704,N_17432,N_17255);
nor U17705 (N_17705,N_17486,N_17418);
or U17706 (N_17706,N_17086,N_17101);
nand U17707 (N_17707,N_17473,N_17382);
xnor U17708 (N_17708,N_17341,N_17237);
and U17709 (N_17709,N_17095,N_17256);
nand U17710 (N_17710,N_17152,N_17494);
and U17711 (N_17711,N_17453,N_17261);
xnor U17712 (N_17712,N_17243,N_17229);
and U17713 (N_17713,N_17001,N_17337);
or U17714 (N_17714,N_17223,N_17487);
or U17715 (N_17715,N_17044,N_17409);
xnor U17716 (N_17716,N_17363,N_17019);
nand U17717 (N_17717,N_17358,N_17080);
nor U17718 (N_17718,N_17427,N_17091);
nand U17719 (N_17719,N_17036,N_17391);
xor U17720 (N_17720,N_17349,N_17476);
nor U17721 (N_17721,N_17433,N_17069);
xnor U17722 (N_17722,N_17099,N_17225);
xnor U17723 (N_17723,N_17319,N_17047);
xor U17724 (N_17724,N_17412,N_17443);
or U17725 (N_17725,N_17002,N_17485);
xnor U17726 (N_17726,N_17457,N_17158);
or U17727 (N_17727,N_17386,N_17155);
nand U17728 (N_17728,N_17398,N_17318);
nor U17729 (N_17729,N_17217,N_17448);
nor U17730 (N_17730,N_17401,N_17411);
or U17731 (N_17731,N_17218,N_17260);
nor U17732 (N_17732,N_17090,N_17407);
and U17733 (N_17733,N_17351,N_17135);
xnor U17734 (N_17734,N_17210,N_17484);
or U17735 (N_17735,N_17013,N_17075);
nor U17736 (N_17736,N_17068,N_17233);
or U17737 (N_17737,N_17367,N_17120);
or U17738 (N_17738,N_17127,N_17232);
xor U17739 (N_17739,N_17055,N_17025);
xnor U17740 (N_17740,N_17315,N_17014);
nor U17741 (N_17741,N_17393,N_17447);
and U17742 (N_17742,N_17293,N_17317);
xor U17743 (N_17743,N_17234,N_17183);
and U17744 (N_17744,N_17271,N_17266);
and U17745 (N_17745,N_17088,N_17007);
and U17746 (N_17746,N_17459,N_17040);
or U17747 (N_17747,N_17193,N_17246);
xnor U17748 (N_17748,N_17380,N_17404);
and U17749 (N_17749,N_17333,N_17482);
nand U17750 (N_17750,N_17220,N_17327);
and U17751 (N_17751,N_17238,N_17258);
or U17752 (N_17752,N_17304,N_17328);
nand U17753 (N_17753,N_17177,N_17351);
or U17754 (N_17754,N_17011,N_17307);
or U17755 (N_17755,N_17170,N_17231);
and U17756 (N_17756,N_17438,N_17354);
and U17757 (N_17757,N_17189,N_17180);
and U17758 (N_17758,N_17143,N_17222);
and U17759 (N_17759,N_17485,N_17461);
nor U17760 (N_17760,N_17152,N_17287);
xnor U17761 (N_17761,N_17340,N_17000);
nand U17762 (N_17762,N_17471,N_17099);
or U17763 (N_17763,N_17422,N_17196);
nor U17764 (N_17764,N_17005,N_17312);
nor U17765 (N_17765,N_17185,N_17405);
or U17766 (N_17766,N_17363,N_17012);
nor U17767 (N_17767,N_17134,N_17191);
and U17768 (N_17768,N_17387,N_17254);
nand U17769 (N_17769,N_17245,N_17139);
or U17770 (N_17770,N_17001,N_17096);
xor U17771 (N_17771,N_17371,N_17034);
xnor U17772 (N_17772,N_17074,N_17020);
nor U17773 (N_17773,N_17380,N_17244);
and U17774 (N_17774,N_17218,N_17325);
nor U17775 (N_17775,N_17461,N_17157);
or U17776 (N_17776,N_17278,N_17071);
nor U17777 (N_17777,N_17226,N_17242);
and U17778 (N_17778,N_17440,N_17243);
or U17779 (N_17779,N_17076,N_17426);
or U17780 (N_17780,N_17035,N_17236);
and U17781 (N_17781,N_17002,N_17453);
or U17782 (N_17782,N_17069,N_17011);
nand U17783 (N_17783,N_17177,N_17266);
nor U17784 (N_17784,N_17126,N_17103);
nand U17785 (N_17785,N_17358,N_17224);
and U17786 (N_17786,N_17319,N_17459);
nor U17787 (N_17787,N_17432,N_17424);
and U17788 (N_17788,N_17022,N_17070);
xor U17789 (N_17789,N_17233,N_17370);
nor U17790 (N_17790,N_17245,N_17200);
xor U17791 (N_17791,N_17490,N_17327);
xnor U17792 (N_17792,N_17056,N_17006);
nand U17793 (N_17793,N_17304,N_17181);
and U17794 (N_17794,N_17141,N_17482);
nor U17795 (N_17795,N_17119,N_17468);
and U17796 (N_17796,N_17247,N_17048);
nand U17797 (N_17797,N_17005,N_17145);
or U17798 (N_17798,N_17302,N_17190);
and U17799 (N_17799,N_17168,N_17391);
xor U17800 (N_17800,N_17424,N_17067);
nand U17801 (N_17801,N_17221,N_17002);
and U17802 (N_17802,N_17457,N_17123);
nor U17803 (N_17803,N_17297,N_17320);
nor U17804 (N_17804,N_17180,N_17208);
and U17805 (N_17805,N_17046,N_17274);
or U17806 (N_17806,N_17482,N_17461);
xnor U17807 (N_17807,N_17462,N_17437);
and U17808 (N_17808,N_17322,N_17123);
and U17809 (N_17809,N_17355,N_17312);
xor U17810 (N_17810,N_17443,N_17479);
nand U17811 (N_17811,N_17075,N_17156);
or U17812 (N_17812,N_17497,N_17279);
or U17813 (N_17813,N_17204,N_17062);
and U17814 (N_17814,N_17184,N_17127);
and U17815 (N_17815,N_17018,N_17406);
xnor U17816 (N_17816,N_17479,N_17386);
nand U17817 (N_17817,N_17196,N_17006);
or U17818 (N_17818,N_17495,N_17385);
nand U17819 (N_17819,N_17181,N_17002);
or U17820 (N_17820,N_17312,N_17279);
nor U17821 (N_17821,N_17414,N_17149);
nand U17822 (N_17822,N_17393,N_17102);
and U17823 (N_17823,N_17068,N_17069);
xnor U17824 (N_17824,N_17300,N_17026);
nand U17825 (N_17825,N_17352,N_17351);
and U17826 (N_17826,N_17312,N_17134);
nor U17827 (N_17827,N_17313,N_17053);
nor U17828 (N_17828,N_17380,N_17237);
and U17829 (N_17829,N_17498,N_17424);
and U17830 (N_17830,N_17048,N_17047);
nand U17831 (N_17831,N_17163,N_17178);
nor U17832 (N_17832,N_17382,N_17364);
or U17833 (N_17833,N_17315,N_17395);
nand U17834 (N_17834,N_17183,N_17240);
nor U17835 (N_17835,N_17237,N_17399);
nor U17836 (N_17836,N_17131,N_17172);
or U17837 (N_17837,N_17470,N_17058);
and U17838 (N_17838,N_17102,N_17249);
xnor U17839 (N_17839,N_17409,N_17000);
xnor U17840 (N_17840,N_17410,N_17363);
and U17841 (N_17841,N_17367,N_17290);
and U17842 (N_17842,N_17028,N_17275);
xnor U17843 (N_17843,N_17058,N_17490);
and U17844 (N_17844,N_17475,N_17295);
and U17845 (N_17845,N_17054,N_17377);
and U17846 (N_17846,N_17237,N_17171);
or U17847 (N_17847,N_17337,N_17048);
or U17848 (N_17848,N_17473,N_17414);
or U17849 (N_17849,N_17392,N_17077);
or U17850 (N_17850,N_17398,N_17249);
xor U17851 (N_17851,N_17314,N_17217);
nand U17852 (N_17852,N_17343,N_17210);
or U17853 (N_17853,N_17469,N_17263);
nand U17854 (N_17854,N_17475,N_17368);
and U17855 (N_17855,N_17421,N_17265);
nand U17856 (N_17856,N_17324,N_17371);
or U17857 (N_17857,N_17103,N_17075);
xor U17858 (N_17858,N_17213,N_17496);
nor U17859 (N_17859,N_17190,N_17188);
and U17860 (N_17860,N_17367,N_17496);
nor U17861 (N_17861,N_17372,N_17026);
or U17862 (N_17862,N_17052,N_17332);
nand U17863 (N_17863,N_17079,N_17390);
xor U17864 (N_17864,N_17489,N_17186);
or U17865 (N_17865,N_17293,N_17350);
nand U17866 (N_17866,N_17158,N_17292);
nand U17867 (N_17867,N_17480,N_17375);
or U17868 (N_17868,N_17422,N_17079);
or U17869 (N_17869,N_17451,N_17095);
and U17870 (N_17870,N_17248,N_17021);
and U17871 (N_17871,N_17091,N_17462);
and U17872 (N_17872,N_17406,N_17222);
nor U17873 (N_17873,N_17340,N_17165);
nor U17874 (N_17874,N_17379,N_17017);
or U17875 (N_17875,N_17170,N_17287);
nor U17876 (N_17876,N_17178,N_17128);
xor U17877 (N_17877,N_17124,N_17015);
nor U17878 (N_17878,N_17092,N_17388);
or U17879 (N_17879,N_17377,N_17486);
nor U17880 (N_17880,N_17389,N_17487);
and U17881 (N_17881,N_17394,N_17444);
xnor U17882 (N_17882,N_17298,N_17172);
nor U17883 (N_17883,N_17120,N_17374);
nor U17884 (N_17884,N_17412,N_17499);
xnor U17885 (N_17885,N_17163,N_17371);
nand U17886 (N_17886,N_17342,N_17385);
and U17887 (N_17887,N_17220,N_17011);
xor U17888 (N_17888,N_17492,N_17442);
nor U17889 (N_17889,N_17028,N_17027);
or U17890 (N_17890,N_17412,N_17079);
nor U17891 (N_17891,N_17372,N_17253);
nand U17892 (N_17892,N_17314,N_17199);
and U17893 (N_17893,N_17170,N_17023);
and U17894 (N_17894,N_17467,N_17493);
xnor U17895 (N_17895,N_17388,N_17352);
or U17896 (N_17896,N_17286,N_17418);
nand U17897 (N_17897,N_17229,N_17184);
nand U17898 (N_17898,N_17005,N_17158);
nor U17899 (N_17899,N_17450,N_17358);
and U17900 (N_17900,N_17299,N_17471);
xnor U17901 (N_17901,N_17415,N_17313);
and U17902 (N_17902,N_17391,N_17060);
or U17903 (N_17903,N_17216,N_17206);
or U17904 (N_17904,N_17497,N_17326);
xor U17905 (N_17905,N_17073,N_17169);
nand U17906 (N_17906,N_17261,N_17127);
xor U17907 (N_17907,N_17244,N_17233);
xnor U17908 (N_17908,N_17254,N_17097);
nor U17909 (N_17909,N_17171,N_17080);
nor U17910 (N_17910,N_17122,N_17333);
nand U17911 (N_17911,N_17119,N_17464);
or U17912 (N_17912,N_17013,N_17319);
xor U17913 (N_17913,N_17314,N_17326);
nor U17914 (N_17914,N_17392,N_17144);
nand U17915 (N_17915,N_17491,N_17133);
nor U17916 (N_17916,N_17373,N_17263);
and U17917 (N_17917,N_17454,N_17202);
nor U17918 (N_17918,N_17199,N_17455);
nand U17919 (N_17919,N_17022,N_17369);
or U17920 (N_17920,N_17232,N_17255);
nor U17921 (N_17921,N_17384,N_17399);
xnor U17922 (N_17922,N_17321,N_17234);
xnor U17923 (N_17923,N_17096,N_17395);
or U17924 (N_17924,N_17433,N_17398);
or U17925 (N_17925,N_17176,N_17139);
xor U17926 (N_17926,N_17177,N_17203);
nand U17927 (N_17927,N_17324,N_17420);
nor U17928 (N_17928,N_17058,N_17143);
nand U17929 (N_17929,N_17215,N_17017);
or U17930 (N_17930,N_17435,N_17205);
or U17931 (N_17931,N_17199,N_17005);
nand U17932 (N_17932,N_17421,N_17133);
or U17933 (N_17933,N_17232,N_17058);
and U17934 (N_17934,N_17407,N_17154);
nor U17935 (N_17935,N_17171,N_17072);
and U17936 (N_17936,N_17122,N_17002);
nand U17937 (N_17937,N_17031,N_17189);
nand U17938 (N_17938,N_17148,N_17005);
or U17939 (N_17939,N_17200,N_17282);
nand U17940 (N_17940,N_17338,N_17443);
and U17941 (N_17941,N_17331,N_17433);
nor U17942 (N_17942,N_17343,N_17204);
or U17943 (N_17943,N_17219,N_17470);
xnor U17944 (N_17944,N_17061,N_17367);
nor U17945 (N_17945,N_17451,N_17324);
nor U17946 (N_17946,N_17205,N_17158);
nor U17947 (N_17947,N_17160,N_17087);
nand U17948 (N_17948,N_17349,N_17473);
nand U17949 (N_17949,N_17237,N_17004);
nand U17950 (N_17950,N_17275,N_17344);
or U17951 (N_17951,N_17202,N_17265);
and U17952 (N_17952,N_17322,N_17057);
or U17953 (N_17953,N_17119,N_17408);
or U17954 (N_17954,N_17052,N_17410);
nor U17955 (N_17955,N_17338,N_17240);
nand U17956 (N_17956,N_17421,N_17418);
nor U17957 (N_17957,N_17214,N_17043);
nor U17958 (N_17958,N_17335,N_17026);
nand U17959 (N_17959,N_17045,N_17463);
xor U17960 (N_17960,N_17362,N_17429);
nor U17961 (N_17961,N_17322,N_17024);
or U17962 (N_17962,N_17101,N_17097);
nor U17963 (N_17963,N_17351,N_17087);
and U17964 (N_17964,N_17131,N_17100);
or U17965 (N_17965,N_17100,N_17000);
nand U17966 (N_17966,N_17119,N_17201);
and U17967 (N_17967,N_17373,N_17481);
nor U17968 (N_17968,N_17085,N_17330);
nand U17969 (N_17969,N_17126,N_17460);
nand U17970 (N_17970,N_17490,N_17032);
nor U17971 (N_17971,N_17093,N_17001);
nor U17972 (N_17972,N_17355,N_17457);
and U17973 (N_17973,N_17439,N_17340);
nor U17974 (N_17974,N_17333,N_17045);
xnor U17975 (N_17975,N_17266,N_17052);
and U17976 (N_17976,N_17145,N_17297);
nor U17977 (N_17977,N_17414,N_17441);
nand U17978 (N_17978,N_17319,N_17469);
nor U17979 (N_17979,N_17109,N_17035);
nor U17980 (N_17980,N_17320,N_17342);
nand U17981 (N_17981,N_17413,N_17285);
or U17982 (N_17982,N_17077,N_17104);
and U17983 (N_17983,N_17314,N_17142);
nand U17984 (N_17984,N_17041,N_17218);
or U17985 (N_17985,N_17118,N_17454);
xnor U17986 (N_17986,N_17209,N_17305);
or U17987 (N_17987,N_17386,N_17478);
or U17988 (N_17988,N_17098,N_17350);
and U17989 (N_17989,N_17156,N_17310);
or U17990 (N_17990,N_17155,N_17452);
nor U17991 (N_17991,N_17462,N_17151);
xor U17992 (N_17992,N_17421,N_17293);
or U17993 (N_17993,N_17161,N_17364);
xor U17994 (N_17994,N_17306,N_17193);
nand U17995 (N_17995,N_17253,N_17352);
nor U17996 (N_17996,N_17305,N_17279);
xnor U17997 (N_17997,N_17019,N_17008);
xor U17998 (N_17998,N_17362,N_17098);
xnor U17999 (N_17999,N_17422,N_17291);
and U18000 (N_18000,N_17526,N_17994);
nor U18001 (N_18001,N_17591,N_17594);
and U18002 (N_18002,N_17802,N_17668);
or U18003 (N_18003,N_17933,N_17694);
and U18004 (N_18004,N_17882,N_17809);
nor U18005 (N_18005,N_17761,N_17639);
nor U18006 (N_18006,N_17716,N_17949);
xor U18007 (N_18007,N_17930,N_17601);
and U18008 (N_18008,N_17756,N_17862);
xnor U18009 (N_18009,N_17645,N_17599);
xnor U18010 (N_18010,N_17845,N_17648);
nand U18011 (N_18011,N_17695,N_17530);
or U18012 (N_18012,N_17532,N_17989);
and U18013 (N_18013,N_17813,N_17541);
nand U18014 (N_18014,N_17792,N_17634);
and U18015 (N_18015,N_17707,N_17570);
nor U18016 (N_18016,N_17840,N_17603);
nor U18017 (N_18017,N_17640,N_17647);
or U18018 (N_18018,N_17965,N_17927);
and U18019 (N_18019,N_17614,N_17995);
nand U18020 (N_18020,N_17819,N_17589);
nor U18021 (N_18021,N_17925,N_17698);
and U18022 (N_18022,N_17699,N_17815);
or U18023 (N_18023,N_17774,N_17737);
and U18024 (N_18024,N_17676,N_17944);
xor U18025 (N_18025,N_17818,N_17899);
xnor U18026 (N_18026,N_17666,N_17598);
or U18027 (N_18027,N_17613,N_17763);
nor U18028 (N_18028,N_17664,N_17654);
and U18029 (N_18029,N_17890,N_17606);
or U18030 (N_18030,N_17875,N_17799);
and U18031 (N_18031,N_17857,N_17978);
or U18032 (N_18032,N_17775,N_17896);
xnor U18033 (N_18033,N_17521,N_17936);
nand U18034 (N_18034,N_17754,N_17502);
and U18035 (N_18035,N_17710,N_17827);
nor U18036 (N_18036,N_17977,N_17876);
and U18037 (N_18037,N_17718,N_17981);
and U18038 (N_18038,N_17895,N_17586);
nor U18039 (N_18039,N_17641,N_17773);
and U18040 (N_18040,N_17968,N_17579);
xor U18041 (N_18041,N_17536,N_17672);
nand U18042 (N_18042,N_17758,N_17663);
and U18043 (N_18043,N_17904,N_17905);
nor U18044 (N_18044,N_17538,N_17630);
xnor U18045 (N_18045,N_17726,N_17920);
xnor U18046 (N_18046,N_17826,N_17839);
nand U18047 (N_18047,N_17789,N_17550);
or U18048 (N_18048,N_17797,N_17912);
xnor U18049 (N_18049,N_17720,N_17881);
xnor U18050 (N_18050,N_17516,N_17955);
xnor U18051 (N_18051,N_17546,N_17796);
and U18052 (N_18052,N_17525,N_17506);
nor U18053 (N_18053,N_17612,N_17836);
nand U18054 (N_18054,N_17730,N_17508);
xnor U18055 (N_18055,N_17846,N_17988);
and U18056 (N_18056,N_17787,N_17572);
and U18057 (N_18057,N_17831,N_17644);
nand U18058 (N_18058,N_17868,N_17585);
or U18059 (N_18059,N_17638,N_17558);
xor U18060 (N_18060,N_17766,N_17979);
or U18061 (N_18061,N_17619,N_17709);
and U18062 (N_18062,N_17690,N_17780);
nand U18063 (N_18063,N_17617,N_17629);
nor U18064 (N_18064,N_17514,N_17545);
nand U18065 (N_18065,N_17755,N_17593);
nand U18066 (N_18066,N_17739,N_17531);
nand U18067 (N_18067,N_17941,N_17627);
and U18068 (N_18068,N_17632,N_17960);
or U18069 (N_18069,N_17733,N_17553);
or U18070 (N_18070,N_17624,N_17577);
and U18071 (N_18071,N_17856,N_17623);
nor U18072 (N_18072,N_17682,N_17747);
nor U18073 (N_18073,N_17885,N_17501);
nand U18074 (N_18074,N_17938,N_17542);
or U18075 (N_18075,N_17537,N_17554);
nor U18076 (N_18076,N_17841,N_17829);
xor U18077 (N_18077,N_17575,N_17866);
xnor U18078 (N_18078,N_17520,N_17587);
xnor U18079 (N_18079,N_17633,N_17686);
nor U18080 (N_18080,N_17740,N_17966);
nand U18081 (N_18081,N_17671,N_17584);
nand U18082 (N_18082,N_17736,N_17511);
nand U18083 (N_18083,N_17771,N_17529);
nor U18084 (N_18084,N_17693,N_17565);
or U18085 (N_18085,N_17732,N_17569);
and U18086 (N_18086,N_17679,N_17801);
or U18087 (N_18087,N_17561,N_17580);
or U18088 (N_18088,N_17855,N_17702);
or U18089 (N_18089,N_17642,N_17877);
nand U18090 (N_18090,N_17910,N_17534);
nand U18091 (N_18091,N_17901,N_17967);
nor U18092 (N_18092,N_17604,N_17953);
and U18093 (N_18093,N_17822,N_17971);
and U18094 (N_18094,N_17777,N_17918);
nand U18095 (N_18095,N_17670,N_17873);
or U18096 (N_18096,N_17932,N_17838);
or U18097 (N_18097,N_17849,N_17620);
nor U18098 (N_18098,N_17893,N_17615);
nor U18099 (N_18099,N_17705,N_17800);
nand U18100 (N_18100,N_17986,N_17888);
nor U18101 (N_18101,N_17980,N_17689);
xor U18102 (N_18102,N_17959,N_17505);
or U18103 (N_18103,N_17688,N_17880);
and U18104 (N_18104,N_17749,N_17753);
xor U18105 (N_18105,N_17790,N_17871);
xnor U18106 (N_18106,N_17785,N_17512);
and U18107 (N_18107,N_17782,N_17625);
and U18108 (N_18108,N_17719,N_17869);
or U18109 (N_18109,N_17578,N_17748);
xor U18110 (N_18110,N_17573,N_17608);
or U18111 (N_18111,N_17607,N_17916);
nand U18112 (N_18112,N_17677,N_17651);
or U18113 (N_18113,N_17768,N_17975);
nand U18114 (N_18114,N_17879,N_17729);
nor U18115 (N_18115,N_17543,N_17674);
or U18116 (N_18116,N_17524,N_17778);
and U18117 (N_18117,N_17811,N_17961);
nand U18118 (N_18118,N_17878,N_17795);
xor U18119 (N_18119,N_17513,N_17909);
and U18120 (N_18120,N_17700,N_17807);
xnor U18121 (N_18121,N_17539,N_17596);
nand U18122 (N_18122,N_17982,N_17970);
nand U18123 (N_18123,N_17704,N_17544);
and U18124 (N_18124,N_17557,N_17844);
nor U18125 (N_18125,N_17969,N_17746);
xnor U18126 (N_18126,N_17590,N_17983);
nand U18127 (N_18127,N_17581,N_17507);
and U18128 (N_18128,N_17781,N_17518);
or U18129 (N_18129,N_17911,N_17821);
or U18130 (N_18130,N_17610,N_17687);
nand U18131 (N_18131,N_17742,N_17697);
nand U18132 (N_18132,N_17919,N_17997);
nand U18133 (N_18133,N_17533,N_17931);
nor U18134 (N_18134,N_17667,N_17816);
nand U18135 (N_18135,N_17863,N_17934);
nand U18136 (N_18136,N_17540,N_17952);
or U18137 (N_18137,N_17765,N_17825);
or U18138 (N_18138,N_17947,N_17655);
or U18139 (N_18139,N_17653,N_17680);
and U18140 (N_18140,N_17987,N_17940);
xnor U18141 (N_18141,N_17884,N_17652);
xnor U18142 (N_18142,N_17996,N_17675);
nand U18143 (N_18143,N_17958,N_17650);
xor U18144 (N_18144,N_17552,N_17973);
nand U18145 (N_18145,N_17832,N_17835);
nor U18146 (N_18146,N_17850,N_17741);
nor U18147 (N_18147,N_17762,N_17887);
xor U18148 (N_18148,N_17939,N_17820);
nand U18149 (N_18149,N_17954,N_17658);
nand U18150 (N_18150,N_17523,N_17963);
nand U18151 (N_18151,N_17808,N_17517);
or U18152 (N_18152,N_17728,N_17510);
or U18153 (N_18153,N_17528,N_17990);
xnor U18154 (N_18154,N_17559,N_17837);
nor U18155 (N_18155,N_17784,N_17847);
and U18156 (N_18156,N_17722,N_17595);
or U18157 (N_18157,N_17870,N_17600);
nor U18158 (N_18158,N_17872,N_17571);
nor U18159 (N_18159,N_17555,N_17972);
or U18160 (N_18160,N_17738,N_17928);
or U18161 (N_18161,N_17891,N_17860);
xnor U18162 (N_18162,N_17892,N_17805);
nand U18163 (N_18163,N_17976,N_17929);
or U18164 (N_18164,N_17576,N_17984);
and U18165 (N_18165,N_17854,N_17611);
or U18166 (N_18166,N_17567,N_17556);
nand U18167 (N_18167,N_17894,N_17964);
xor U18168 (N_18168,N_17724,N_17527);
xnor U18169 (N_18169,N_17588,N_17776);
xnor U18170 (N_18170,N_17669,N_17951);
and U18171 (N_18171,N_17662,N_17824);
nand U18172 (N_18172,N_17767,N_17812);
or U18173 (N_18173,N_17685,N_17937);
xnor U18174 (N_18174,N_17605,N_17962);
nor U18175 (N_18175,N_17548,N_17574);
or U18176 (N_18176,N_17999,N_17779);
nand U18177 (N_18177,N_17725,N_17810);
nand U18178 (N_18178,N_17804,N_17743);
nor U18179 (N_18179,N_17752,N_17744);
and U18180 (N_18180,N_17843,N_17865);
or U18181 (N_18181,N_17727,N_17681);
nand U18182 (N_18182,N_17830,N_17745);
nand U18183 (N_18183,N_17957,N_17735);
nor U18184 (N_18184,N_17913,N_17902);
xnor U18185 (N_18185,N_17649,N_17943);
nand U18186 (N_18186,N_17900,N_17564);
nor U18187 (N_18187,N_17769,N_17562);
and U18188 (N_18188,N_17609,N_17833);
nor U18189 (N_18189,N_17519,N_17874);
or U18190 (N_18190,N_17924,N_17906);
nor U18191 (N_18191,N_17621,N_17858);
nor U18192 (N_18192,N_17898,N_17721);
nand U18193 (N_18193,N_17717,N_17848);
nor U18194 (N_18194,N_17656,N_17974);
nor U18195 (N_18195,N_17760,N_17515);
nor U18196 (N_18196,N_17635,N_17903);
nor U18197 (N_18197,N_17713,N_17950);
nand U18198 (N_18198,N_17500,N_17788);
and U18199 (N_18199,N_17915,N_17616);
nand U18200 (N_18200,N_17946,N_17631);
and U18201 (N_18201,N_17683,N_17646);
nor U18202 (N_18202,N_17993,N_17628);
or U18203 (N_18203,N_17568,N_17926);
or U18204 (N_18204,N_17706,N_17908);
and U18205 (N_18205,N_17923,N_17842);
nor U18206 (N_18206,N_17673,N_17886);
or U18207 (N_18207,N_17956,N_17823);
and U18208 (N_18208,N_17907,N_17817);
nand U18209 (N_18209,N_17560,N_17889);
nand U18210 (N_18210,N_17547,N_17897);
nand U18211 (N_18211,N_17509,N_17867);
or U18212 (N_18212,N_17757,N_17791);
and U18213 (N_18213,N_17985,N_17859);
nand U18214 (N_18214,N_17691,N_17659);
nor U18215 (N_18215,N_17992,N_17636);
nor U18216 (N_18216,N_17626,N_17597);
nand U18217 (N_18217,N_17711,N_17715);
and U18218 (N_18218,N_17714,N_17883);
and U18219 (N_18219,N_17917,N_17921);
nor U18220 (N_18220,N_17643,N_17582);
nand U18221 (N_18221,N_17549,N_17914);
xor U18222 (N_18222,N_17551,N_17661);
nor U18223 (N_18223,N_17803,N_17786);
or U18224 (N_18224,N_17814,N_17566);
nor U18225 (N_18225,N_17504,N_17991);
or U18226 (N_18226,N_17563,N_17535);
nand U18227 (N_18227,N_17770,N_17592);
nand U18228 (N_18228,N_17852,N_17783);
and U18229 (N_18229,N_17731,N_17853);
and U18230 (N_18230,N_17750,N_17945);
nand U18231 (N_18231,N_17712,N_17657);
nor U18232 (N_18232,N_17948,N_17751);
xor U18233 (N_18233,N_17922,N_17583);
xor U18234 (N_18234,N_17806,N_17764);
or U18235 (N_18235,N_17703,N_17637);
and U18236 (N_18236,N_17622,N_17692);
and U18237 (N_18237,N_17772,N_17851);
nor U18238 (N_18238,N_17998,N_17522);
nor U18239 (N_18239,N_17864,N_17503);
nand U18240 (N_18240,N_17794,N_17798);
and U18241 (N_18241,N_17723,N_17834);
xnor U18242 (N_18242,N_17793,N_17696);
nand U18243 (N_18243,N_17708,N_17678);
and U18244 (N_18244,N_17701,N_17602);
nand U18245 (N_18245,N_17828,N_17861);
and U18246 (N_18246,N_17684,N_17942);
nor U18247 (N_18247,N_17734,N_17618);
xnor U18248 (N_18248,N_17935,N_17660);
nand U18249 (N_18249,N_17665,N_17759);
nand U18250 (N_18250,N_17701,N_17535);
nor U18251 (N_18251,N_17524,N_17804);
nand U18252 (N_18252,N_17538,N_17946);
xnor U18253 (N_18253,N_17592,N_17714);
or U18254 (N_18254,N_17741,N_17689);
and U18255 (N_18255,N_17527,N_17838);
nand U18256 (N_18256,N_17554,N_17982);
nand U18257 (N_18257,N_17696,N_17856);
and U18258 (N_18258,N_17631,N_17665);
nand U18259 (N_18259,N_17548,N_17957);
or U18260 (N_18260,N_17936,N_17844);
nor U18261 (N_18261,N_17748,N_17616);
nand U18262 (N_18262,N_17554,N_17826);
or U18263 (N_18263,N_17817,N_17756);
nor U18264 (N_18264,N_17861,N_17723);
xor U18265 (N_18265,N_17536,N_17545);
and U18266 (N_18266,N_17783,N_17701);
nor U18267 (N_18267,N_17791,N_17566);
nor U18268 (N_18268,N_17505,N_17864);
xor U18269 (N_18269,N_17517,N_17890);
nand U18270 (N_18270,N_17779,N_17695);
nor U18271 (N_18271,N_17573,N_17888);
xnor U18272 (N_18272,N_17932,N_17757);
nor U18273 (N_18273,N_17810,N_17973);
and U18274 (N_18274,N_17858,N_17905);
nor U18275 (N_18275,N_17600,N_17563);
nor U18276 (N_18276,N_17719,N_17810);
nand U18277 (N_18277,N_17664,N_17788);
or U18278 (N_18278,N_17712,N_17854);
nor U18279 (N_18279,N_17839,N_17565);
and U18280 (N_18280,N_17516,N_17802);
nand U18281 (N_18281,N_17826,N_17803);
or U18282 (N_18282,N_17862,N_17795);
nand U18283 (N_18283,N_17904,N_17519);
nor U18284 (N_18284,N_17656,N_17622);
xor U18285 (N_18285,N_17549,N_17635);
or U18286 (N_18286,N_17647,N_17582);
or U18287 (N_18287,N_17952,N_17701);
nand U18288 (N_18288,N_17906,N_17664);
or U18289 (N_18289,N_17500,N_17732);
nor U18290 (N_18290,N_17594,N_17988);
or U18291 (N_18291,N_17699,N_17720);
and U18292 (N_18292,N_17866,N_17557);
nand U18293 (N_18293,N_17808,N_17737);
or U18294 (N_18294,N_17512,N_17675);
nor U18295 (N_18295,N_17896,N_17819);
and U18296 (N_18296,N_17527,N_17802);
or U18297 (N_18297,N_17788,N_17768);
nand U18298 (N_18298,N_17595,N_17926);
xor U18299 (N_18299,N_17922,N_17720);
or U18300 (N_18300,N_17942,N_17729);
or U18301 (N_18301,N_17970,N_17937);
nor U18302 (N_18302,N_17951,N_17894);
nor U18303 (N_18303,N_17997,N_17939);
or U18304 (N_18304,N_17526,N_17667);
and U18305 (N_18305,N_17938,N_17924);
nand U18306 (N_18306,N_17918,N_17504);
or U18307 (N_18307,N_17935,N_17569);
and U18308 (N_18308,N_17972,N_17908);
or U18309 (N_18309,N_17975,N_17741);
nor U18310 (N_18310,N_17524,N_17593);
nor U18311 (N_18311,N_17948,N_17694);
nor U18312 (N_18312,N_17975,N_17929);
and U18313 (N_18313,N_17676,N_17959);
nor U18314 (N_18314,N_17867,N_17641);
nor U18315 (N_18315,N_17880,N_17704);
or U18316 (N_18316,N_17865,N_17601);
nor U18317 (N_18317,N_17522,N_17796);
nand U18318 (N_18318,N_17763,N_17658);
nor U18319 (N_18319,N_17735,N_17739);
or U18320 (N_18320,N_17954,N_17756);
xor U18321 (N_18321,N_17942,N_17711);
and U18322 (N_18322,N_17890,N_17579);
and U18323 (N_18323,N_17513,N_17869);
nand U18324 (N_18324,N_17501,N_17892);
and U18325 (N_18325,N_17718,N_17702);
and U18326 (N_18326,N_17786,N_17584);
or U18327 (N_18327,N_17709,N_17526);
xor U18328 (N_18328,N_17823,N_17720);
nor U18329 (N_18329,N_17609,N_17557);
and U18330 (N_18330,N_17515,N_17719);
xnor U18331 (N_18331,N_17950,N_17763);
nor U18332 (N_18332,N_17780,N_17919);
nand U18333 (N_18333,N_17548,N_17527);
or U18334 (N_18334,N_17697,N_17858);
and U18335 (N_18335,N_17516,N_17630);
xor U18336 (N_18336,N_17688,N_17776);
or U18337 (N_18337,N_17568,N_17542);
or U18338 (N_18338,N_17945,N_17701);
nand U18339 (N_18339,N_17659,N_17753);
nor U18340 (N_18340,N_17553,N_17966);
nor U18341 (N_18341,N_17840,N_17503);
nor U18342 (N_18342,N_17971,N_17904);
and U18343 (N_18343,N_17820,N_17993);
xor U18344 (N_18344,N_17554,N_17510);
xor U18345 (N_18345,N_17923,N_17732);
nor U18346 (N_18346,N_17598,N_17810);
nor U18347 (N_18347,N_17808,N_17665);
or U18348 (N_18348,N_17521,N_17610);
or U18349 (N_18349,N_17928,N_17702);
nor U18350 (N_18350,N_17845,N_17544);
and U18351 (N_18351,N_17986,N_17776);
and U18352 (N_18352,N_17755,N_17802);
nand U18353 (N_18353,N_17617,N_17926);
xnor U18354 (N_18354,N_17610,N_17791);
nand U18355 (N_18355,N_17566,N_17556);
nor U18356 (N_18356,N_17567,N_17546);
nor U18357 (N_18357,N_17555,N_17980);
xnor U18358 (N_18358,N_17628,N_17915);
and U18359 (N_18359,N_17617,N_17535);
nor U18360 (N_18360,N_17828,N_17532);
nand U18361 (N_18361,N_17911,N_17597);
or U18362 (N_18362,N_17542,N_17596);
and U18363 (N_18363,N_17857,N_17940);
or U18364 (N_18364,N_17848,N_17926);
nor U18365 (N_18365,N_17919,N_17938);
xnor U18366 (N_18366,N_17958,N_17981);
xnor U18367 (N_18367,N_17753,N_17697);
nor U18368 (N_18368,N_17570,N_17525);
xnor U18369 (N_18369,N_17986,N_17562);
and U18370 (N_18370,N_17995,N_17717);
and U18371 (N_18371,N_17595,N_17830);
xnor U18372 (N_18372,N_17855,N_17715);
or U18373 (N_18373,N_17987,N_17693);
xnor U18374 (N_18374,N_17964,N_17524);
and U18375 (N_18375,N_17818,N_17798);
nand U18376 (N_18376,N_17979,N_17963);
xnor U18377 (N_18377,N_17624,N_17705);
xnor U18378 (N_18378,N_17893,N_17530);
nand U18379 (N_18379,N_17605,N_17564);
and U18380 (N_18380,N_17674,N_17612);
or U18381 (N_18381,N_17565,N_17775);
nor U18382 (N_18382,N_17862,N_17902);
and U18383 (N_18383,N_17587,N_17845);
or U18384 (N_18384,N_17587,N_17854);
or U18385 (N_18385,N_17530,N_17616);
nor U18386 (N_18386,N_17502,N_17717);
nor U18387 (N_18387,N_17819,N_17617);
nor U18388 (N_18388,N_17974,N_17930);
or U18389 (N_18389,N_17542,N_17570);
nor U18390 (N_18390,N_17781,N_17589);
nor U18391 (N_18391,N_17998,N_17679);
nand U18392 (N_18392,N_17958,N_17671);
nor U18393 (N_18393,N_17964,N_17638);
nor U18394 (N_18394,N_17582,N_17692);
and U18395 (N_18395,N_17573,N_17577);
nand U18396 (N_18396,N_17877,N_17543);
nand U18397 (N_18397,N_17972,N_17504);
or U18398 (N_18398,N_17751,N_17847);
nor U18399 (N_18399,N_17888,N_17600);
xor U18400 (N_18400,N_17872,N_17916);
xnor U18401 (N_18401,N_17728,N_17600);
xor U18402 (N_18402,N_17742,N_17718);
nor U18403 (N_18403,N_17579,N_17845);
xnor U18404 (N_18404,N_17633,N_17571);
nor U18405 (N_18405,N_17658,N_17593);
nor U18406 (N_18406,N_17669,N_17975);
nor U18407 (N_18407,N_17928,N_17931);
nand U18408 (N_18408,N_17739,N_17663);
nand U18409 (N_18409,N_17688,N_17740);
xor U18410 (N_18410,N_17621,N_17951);
xor U18411 (N_18411,N_17614,N_17864);
or U18412 (N_18412,N_17875,N_17646);
nor U18413 (N_18413,N_17890,N_17870);
xor U18414 (N_18414,N_17553,N_17538);
nand U18415 (N_18415,N_17777,N_17510);
or U18416 (N_18416,N_17701,N_17555);
xnor U18417 (N_18417,N_17915,N_17881);
xor U18418 (N_18418,N_17540,N_17615);
or U18419 (N_18419,N_17725,N_17611);
nor U18420 (N_18420,N_17599,N_17783);
or U18421 (N_18421,N_17826,N_17745);
or U18422 (N_18422,N_17906,N_17784);
and U18423 (N_18423,N_17918,N_17751);
and U18424 (N_18424,N_17557,N_17645);
xor U18425 (N_18425,N_17857,N_17854);
nor U18426 (N_18426,N_17527,N_17511);
nor U18427 (N_18427,N_17823,N_17643);
xor U18428 (N_18428,N_17877,N_17869);
and U18429 (N_18429,N_17616,N_17617);
xnor U18430 (N_18430,N_17667,N_17831);
xor U18431 (N_18431,N_17611,N_17652);
nand U18432 (N_18432,N_17894,N_17953);
nor U18433 (N_18433,N_17511,N_17641);
nand U18434 (N_18434,N_17646,N_17578);
nor U18435 (N_18435,N_17881,N_17858);
xnor U18436 (N_18436,N_17697,N_17520);
nand U18437 (N_18437,N_17896,N_17516);
nor U18438 (N_18438,N_17573,N_17635);
or U18439 (N_18439,N_17962,N_17644);
nand U18440 (N_18440,N_17609,N_17979);
nand U18441 (N_18441,N_17872,N_17574);
nor U18442 (N_18442,N_17859,N_17532);
or U18443 (N_18443,N_17538,N_17818);
xor U18444 (N_18444,N_17644,N_17898);
xnor U18445 (N_18445,N_17802,N_17563);
or U18446 (N_18446,N_17546,N_17539);
nor U18447 (N_18447,N_17647,N_17933);
xor U18448 (N_18448,N_17989,N_17971);
or U18449 (N_18449,N_17796,N_17904);
or U18450 (N_18450,N_17868,N_17864);
xnor U18451 (N_18451,N_17642,N_17649);
nor U18452 (N_18452,N_17819,N_17912);
nand U18453 (N_18453,N_17777,N_17578);
and U18454 (N_18454,N_17738,N_17790);
nand U18455 (N_18455,N_17654,N_17636);
xnor U18456 (N_18456,N_17797,N_17562);
nand U18457 (N_18457,N_17585,N_17960);
or U18458 (N_18458,N_17748,N_17520);
nand U18459 (N_18459,N_17835,N_17720);
xor U18460 (N_18460,N_17597,N_17929);
xnor U18461 (N_18461,N_17714,N_17737);
xnor U18462 (N_18462,N_17594,N_17720);
and U18463 (N_18463,N_17828,N_17964);
and U18464 (N_18464,N_17693,N_17612);
nand U18465 (N_18465,N_17690,N_17515);
xnor U18466 (N_18466,N_17719,N_17600);
nor U18467 (N_18467,N_17663,N_17731);
or U18468 (N_18468,N_17643,N_17939);
or U18469 (N_18469,N_17937,N_17950);
nand U18470 (N_18470,N_17947,N_17871);
and U18471 (N_18471,N_17962,N_17588);
xnor U18472 (N_18472,N_17704,N_17667);
nand U18473 (N_18473,N_17717,N_17778);
xnor U18474 (N_18474,N_17515,N_17837);
nor U18475 (N_18475,N_17767,N_17824);
and U18476 (N_18476,N_17787,N_17540);
xnor U18477 (N_18477,N_17815,N_17781);
and U18478 (N_18478,N_17735,N_17882);
nand U18479 (N_18479,N_17665,N_17721);
xnor U18480 (N_18480,N_17913,N_17746);
nand U18481 (N_18481,N_17868,N_17537);
nor U18482 (N_18482,N_17513,N_17878);
nor U18483 (N_18483,N_17666,N_17718);
xnor U18484 (N_18484,N_17687,N_17671);
nand U18485 (N_18485,N_17802,N_17783);
nand U18486 (N_18486,N_17774,N_17743);
xor U18487 (N_18487,N_17760,N_17539);
nor U18488 (N_18488,N_17863,N_17730);
nand U18489 (N_18489,N_17851,N_17548);
nor U18490 (N_18490,N_17931,N_17506);
and U18491 (N_18491,N_17618,N_17750);
xor U18492 (N_18492,N_17986,N_17599);
xnor U18493 (N_18493,N_17709,N_17656);
and U18494 (N_18494,N_17920,N_17618);
nor U18495 (N_18495,N_17959,N_17669);
nor U18496 (N_18496,N_17868,N_17506);
or U18497 (N_18497,N_17534,N_17651);
xnor U18498 (N_18498,N_17978,N_17763);
or U18499 (N_18499,N_17817,N_17547);
nor U18500 (N_18500,N_18021,N_18400);
nand U18501 (N_18501,N_18161,N_18132);
xnor U18502 (N_18502,N_18305,N_18251);
nand U18503 (N_18503,N_18091,N_18254);
xnor U18504 (N_18504,N_18367,N_18278);
xor U18505 (N_18505,N_18435,N_18436);
xnor U18506 (N_18506,N_18343,N_18123);
xor U18507 (N_18507,N_18065,N_18330);
nor U18508 (N_18508,N_18474,N_18110);
and U18509 (N_18509,N_18419,N_18147);
or U18510 (N_18510,N_18046,N_18177);
xnor U18511 (N_18511,N_18024,N_18019);
and U18512 (N_18512,N_18433,N_18472);
and U18513 (N_18513,N_18141,N_18238);
and U18514 (N_18514,N_18361,N_18095);
and U18515 (N_18515,N_18009,N_18338);
or U18516 (N_18516,N_18350,N_18039);
xor U18517 (N_18517,N_18490,N_18062);
and U18518 (N_18518,N_18405,N_18285);
nand U18519 (N_18519,N_18037,N_18340);
nand U18520 (N_18520,N_18003,N_18239);
or U18521 (N_18521,N_18189,N_18026);
and U18522 (N_18522,N_18374,N_18449);
and U18523 (N_18523,N_18059,N_18210);
or U18524 (N_18524,N_18319,N_18315);
nand U18525 (N_18525,N_18455,N_18415);
nor U18526 (N_18526,N_18420,N_18223);
or U18527 (N_18527,N_18067,N_18380);
nand U18528 (N_18528,N_18001,N_18148);
nand U18529 (N_18529,N_18035,N_18480);
xor U18530 (N_18530,N_18297,N_18152);
and U18531 (N_18531,N_18324,N_18334);
or U18532 (N_18532,N_18481,N_18401);
or U18533 (N_18533,N_18450,N_18145);
nand U18534 (N_18534,N_18103,N_18393);
xor U18535 (N_18535,N_18206,N_18234);
nor U18536 (N_18536,N_18235,N_18366);
nand U18537 (N_18537,N_18335,N_18448);
or U18538 (N_18538,N_18329,N_18248);
and U18539 (N_18539,N_18004,N_18006);
nand U18540 (N_18540,N_18398,N_18341);
or U18541 (N_18541,N_18317,N_18016);
nor U18542 (N_18542,N_18089,N_18201);
nand U18543 (N_18543,N_18042,N_18224);
nor U18544 (N_18544,N_18121,N_18051);
nand U18545 (N_18545,N_18243,N_18069);
and U18546 (N_18546,N_18176,N_18404);
and U18547 (N_18547,N_18390,N_18137);
or U18548 (N_18548,N_18286,N_18219);
xor U18549 (N_18549,N_18063,N_18339);
xnor U18550 (N_18550,N_18300,N_18395);
and U18551 (N_18551,N_18074,N_18055);
and U18552 (N_18552,N_18231,N_18421);
nand U18553 (N_18553,N_18213,N_18038);
and U18554 (N_18554,N_18183,N_18031);
nor U18555 (N_18555,N_18119,N_18475);
nor U18556 (N_18556,N_18295,N_18032);
and U18557 (N_18557,N_18205,N_18386);
or U18558 (N_18558,N_18198,N_18108);
xor U18559 (N_18559,N_18075,N_18427);
nand U18560 (N_18560,N_18258,N_18222);
and U18561 (N_18561,N_18247,N_18263);
nand U18562 (N_18562,N_18154,N_18406);
and U18563 (N_18563,N_18098,N_18166);
xor U18564 (N_18564,N_18259,N_18458);
nor U18565 (N_18565,N_18129,N_18280);
nand U18566 (N_18566,N_18272,N_18376);
nor U18567 (N_18567,N_18167,N_18347);
xor U18568 (N_18568,N_18498,N_18159);
xnor U18569 (N_18569,N_18471,N_18113);
and U18570 (N_18570,N_18131,N_18264);
or U18571 (N_18571,N_18208,N_18283);
nor U18572 (N_18572,N_18365,N_18105);
nor U18573 (N_18573,N_18076,N_18482);
and U18574 (N_18574,N_18096,N_18168);
nand U18575 (N_18575,N_18157,N_18479);
nor U18576 (N_18576,N_18146,N_18342);
nor U18577 (N_18577,N_18382,N_18158);
nor U18578 (N_18578,N_18190,N_18097);
nand U18579 (N_18579,N_18269,N_18426);
and U18580 (N_18580,N_18478,N_18446);
and U18581 (N_18581,N_18171,N_18277);
nand U18582 (N_18582,N_18495,N_18261);
and U18583 (N_18583,N_18291,N_18072);
nand U18584 (N_18584,N_18360,N_18165);
or U18585 (N_18585,N_18402,N_18211);
or U18586 (N_18586,N_18422,N_18413);
xor U18587 (N_18587,N_18106,N_18028);
nand U18588 (N_18588,N_18044,N_18452);
and U18589 (N_18589,N_18348,N_18034);
or U18590 (N_18590,N_18179,N_18346);
xnor U18591 (N_18591,N_18468,N_18104);
or U18592 (N_18592,N_18194,N_18271);
and U18593 (N_18593,N_18461,N_18212);
xnor U18594 (N_18594,N_18425,N_18227);
nor U18595 (N_18595,N_18333,N_18134);
and U18596 (N_18596,N_18188,N_18394);
nand U18597 (N_18597,N_18181,N_18417);
and U18598 (N_18598,N_18195,N_18388);
nand U18599 (N_18599,N_18245,N_18185);
xor U18600 (N_18600,N_18193,N_18163);
xor U18601 (N_18601,N_18088,N_18312);
nand U18602 (N_18602,N_18497,N_18048);
nor U18603 (N_18603,N_18356,N_18276);
nand U18604 (N_18604,N_18443,N_18151);
or U18605 (N_18605,N_18303,N_18407);
nor U18606 (N_18606,N_18012,N_18217);
nand U18607 (N_18607,N_18030,N_18116);
nand U18608 (N_18608,N_18070,N_18220);
nand U18609 (N_18609,N_18473,N_18029);
nand U18610 (N_18610,N_18314,N_18225);
or U18611 (N_18611,N_18383,N_18424);
xor U18612 (N_18612,N_18444,N_18066);
xnor U18613 (N_18613,N_18270,N_18127);
xor U18614 (N_18614,N_18307,N_18204);
nand U18615 (N_18615,N_18375,N_18470);
nor U18616 (N_18616,N_18354,N_18392);
nor U18617 (N_18617,N_18087,N_18249);
xnor U18618 (N_18618,N_18318,N_18228);
xor U18619 (N_18619,N_18438,N_18336);
nor U18620 (N_18620,N_18408,N_18310);
or U18621 (N_18621,N_18302,N_18207);
or U18622 (N_18622,N_18050,N_18064);
nand U18623 (N_18623,N_18491,N_18149);
xor U18624 (N_18624,N_18080,N_18494);
xor U18625 (N_18625,N_18369,N_18410);
xnor U18626 (N_18626,N_18320,N_18174);
xnor U18627 (N_18627,N_18477,N_18061);
or U18628 (N_18628,N_18265,N_18214);
xor U18629 (N_18629,N_18483,N_18237);
and U18630 (N_18630,N_18043,N_18102);
and U18631 (N_18631,N_18484,N_18010);
nand U18632 (N_18632,N_18018,N_18308);
or U18633 (N_18633,N_18298,N_18118);
or U18634 (N_18634,N_18184,N_18378);
nor U18635 (N_18635,N_18349,N_18486);
nand U18636 (N_18636,N_18294,N_18372);
nand U18637 (N_18637,N_18057,N_18371);
or U18638 (N_18638,N_18133,N_18156);
and U18639 (N_18639,N_18230,N_18391);
nor U18640 (N_18640,N_18496,N_18049);
or U18641 (N_18641,N_18439,N_18288);
and U18642 (N_18642,N_18462,N_18411);
and U18643 (N_18643,N_18164,N_18309);
and U18644 (N_18644,N_18142,N_18437);
nand U18645 (N_18645,N_18327,N_18197);
nand U18646 (N_18646,N_18052,N_18240);
or U18647 (N_18647,N_18389,N_18418);
nor U18648 (N_18648,N_18453,N_18290);
or U18649 (N_18649,N_18492,N_18456);
nand U18650 (N_18650,N_18100,N_18445);
or U18651 (N_18651,N_18172,N_18144);
nor U18652 (N_18652,N_18083,N_18301);
xor U18653 (N_18653,N_18200,N_18430);
nand U18654 (N_18654,N_18429,N_18381);
nor U18655 (N_18655,N_18191,N_18005);
nor U18656 (N_18656,N_18364,N_18092);
and U18657 (N_18657,N_18460,N_18221);
nand U18658 (N_18658,N_18284,N_18485);
nand U18659 (N_18659,N_18428,N_18373);
or U18660 (N_18660,N_18126,N_18178);
nand U18661 (N_18661,N_18466,N_18322);
or U18662 (N_18662,N_18325,N_18332);
nand U18663 (N_18663,N_18111,N_18299);
xnor U18664 (N_18664,N_18273,N_18275);
and U18665 (N_18665,N_18447,N_18357);
or U18666 (N_18666,N_18099,N_18112);
xor U18667 (N_18667,N_18125,N_18022);
xor U18668 (N_18668,N_18316,N_18090);
and U18669 (N_18669,N_18250,N_18465);
nor U18670 (N_18670,N_18107,N_18232);
or U18671 (N_18671,N_18115,N_18236);
nor U18672 (N_18672,N_18441,N_18027);
and U18673 (N_18673,N_18467,N_18081);
nand U18674 (N_18674,N_18182,N_18377);
nor U18675 (N_18675,N_18345,N_18011);
and U18676 (N_18676,N_18464,N_18252);
or U18677 (N_18677,N_18122,N_18139);
xor U18678 (N_18678,N_18257,N_18186);
and U18679 (N_18679,N_18060,N_18084);
xor U18680 (N_18680,N_18442,N_18101);
nand U18681 (N_18681,N_18033,N_18082);
and U18682 (N_18682,N_18279,N_18397);
nor U18683 (N_18683,N_18135,N_18323);
or U18684 (N_18684,N_18241,N_18017);
and U18685 (N_18685,N_18457,N_18109);
nand U18686 (N_18686,N_18169,N_18114);
nor U18687 (N_18687,N_18313,N_18399);
or U18688 (N_18688,N_18140,N_18244);
or U18689 (N_18689,N_18013,N_18358);
or U18690 (N_18690,N_18352,N_18306);
or U18691 (N_18691,N_18362,N_18054);
xnor U18692 (N_18692,N_18047,N_18267);
and U18693 (N_18693,N_18476,N_18431);
or U18694 (N_18694,N_18218,N_18370);
nand U18695 (N_18695,N_18138,N_18053);
nor U18696 (N_18696,N_18488,N_18153);
nor U18697 (N_18697,N_18233,N_18384);
nor U18698 (N_18698,N_18155,N_18175);
or U18699 (N_18699,N_18094,N_18409);
or U18700 (N_18700,N_18293,N_18085);
xor U18701 (N_18701,N_18454,N_18368);
nor U18702 (N_18702,N_18423,N_18120);
xnor U18703 (N_18703,N_18268,N_18403);
xnor U18704 (N_18704,N_18432,N_18292);
and U18705 (N_18705,N_18150,N_18266);
xor U18706 (N_18706,N_18321,N_18199);
nand U18707 (N_18707,N_18287,N_18469);
and U18708 (N_18708,N_18160,N_18187);
or U18709 (N_18709,N_18058,N_18173);
xnor U18710 (N_18710,N_18256,N_18353);
or U18711 (N_18711,N_18162,N_18451);
xor U18712 (N_18712,N_18337,N_18086);
or U18713 (N_18713,N_18056,N_18304);
nor U18714 (N_18714,N_18229,N_18203);
xor U18715 (N_18715,N_18008,N_18412);
nand U18716 (N_18716,N_18282,N_18296);
nor U18717 (N_18717,N_18385,N_18202);
and U18718 (N_18718,N_18260,N_18209);
nor U18719 (N_18719,N_18192,N_18071);
or U18720 (N_18720,N_18093,N_18344);
nor U18721 (N_18721,N_18216,N_18196);
nor U18722 (N_18722,N_18242,N_18117);
nor U18723 (N_18723,N_18226,N_18020);
nand U18724 (N_18724,N_18493,N_18079);
and U18725 (N_18725,N_18328,N_18036);
xnor U18726 (N_18726,N_18459,N_18170);
and U18727 (N_18727,N_18014,N_18414);
and U18728 (N_18728,N_18487,N_18463);
nand U18729 (N_18729,N_18387,N_18274);
nand U18730 (N_18730,N_18180,N_18253);
or U18731 (N_18731,N_18434,N_18040);
xnor U18732 (N_18732,N_18041,N_18068);
nor U18733 (N_18733,N_18363,N_18078);
or U18734 (N_18734,N_18326,N_18281);
and U18735 (N_18735,N_18379,N_18025);
or U18736 (N_18736,N_18311,N_18499);
or U18737 (N_18737,N_18396,N_18215);
or U18738 (N_18738,N_18073,N_18262);
or U18739 (N_18739,N_18489,N_18355);
xor U18740 (N_18740,N_18015,N_18124);
or U18741 (N_18741,N_18023,N_18128);
and U18742 (N_18742,N_18255,N_18000);
nand U18743 (N_18743,N_18440,N_18289);
nor U18744 (N_18744,N_18359,N_18416);
and U18745 (N_18745,N_18136,N_18045);
and U18746 (N_18746,N_18246,N_18130);
or U18747 (N_18747,N_18002,N_18007);
nor U18748 (N_18748,N_18331,N_18351);
and U18749 (N_18749,N_18077,N_18143);
nand U18750 (N_18750,N_18103,N_18324);
nor U18751 (N_18751,N_18057,N_18091);
or U18752 (N_18752,N_18412,N_18387);
and U18753 (N_18753,N_18251,N_18276);
or U18754 (N_18754,N_18107,N_18052);
or U18755 (N_18755,N_18112,N_18170);
or U18756 (N_18756,N_18109,N_18246);
and U18757 (N_18757,N_18487,N_18366);
xnor U18758 (N_18758,N_18010,N_18057);
and U18759 (N_18759,N_18071,N_18440);
or U18760 (N_18760,N_18421,N_18360);
nand U18761 (N_18761,N_18190,N_18495);
xnor U18762 (N_18762,N_18087,N_18364);
nor U18763 (N_18763,N_18413,N_18174);
or U18764 (N_18764,N_18461,N_18375);
xor U18765 (N_18765,N_18106,N_18454);
xor U18766 (N_18766,N_18452,N_18444);
xor U18767 (N_18767,N_18325,N_18125);
nand U18768 (N_18768,N_18365,N_18443);
nor U18769 (N_18769,N_18099,N_18376);
nor U18770 (N_18770,N_18498,N_18351);
xor U18771 (N_18771,N_18191,N_18349);
or U18772 (N_18772,N_18360,N_18454);
nor U18773 (N_18773,N_18380,N_18048);
nand U18774 (N_18774,N_18258,N_18330);
nand U18775 (N_18775,N_18356,N_18432);
nor U18776 (N_18776,N_18477,N_18205);
nand U18777 (N_18777,N_18363,N_18170);
nand U18778 (N_18778,N_18025,N_18156);
nor U18779 (N_18779,N_18430,N_18217);
nor U18780 (N_18780,N_18122,N_18323);
and U18781 (N_18781,N_18427,N_18355);
xor U18782 (N_18782,N_18087,N_18165);
or U18783 (N_18783,N_18360,N_18475);
xnor U18784 (N_18784,N_18087,N_18142);
xor U18785 (N_18785,N_18033,N_18447);
or U18786 (N_18786,N_18315,N_18196);
and U18787 (N_18787,N_18055,N_18279);
and U18788 (N_18788,N_18119,N_18217);
or U18789 (N_18789,N_18188,N_18027);
and U18790 (N_18790,N_18162,N_18144);
and U18791 (N_18791,N_18174,N_18302);
nor U18792 (N_18792,N_18423,N_18380);
xnor U18793 (N_18793,N_18035,N_18151);
nand U18794 (N_18794,N_18062,N_18370);
and U18795 (N_18795,N_18011,N_18452);
xor U18796 (N_18796,N_18248,N_18155);
nor U18797 (N_18797,N_18293,N_18412);
nor U18798 (N_18798,N_18010,N_18127);
xnor U18799 (N_18799,N_18218,N_18418);
nand U18800 (N_18800,N_18285,N_18328);
xor U18801 (N_18801,N_18363,N_18266);
and U18802 (N_18802,N_18168,N_18039);
nor U18803 (N_18803,N_18490,N_18392);
xor U18804 (N_18804,N_18412,N_18269);
nand U18805 (N_18805,N_18325,N_18209);
nor U18806 (N_18806,N_18083,N_18370);
nand U18807 (N_18807,N_18359,N_18070);
and U18808 (N_18808,N_18304,N_18431);
or U18809 (N_18809,N_18397,N_18057);
or U18810 (N_18810,N_18331,N_18099);
nor U18811 (N_18811,N_18145,N_18172);
or U18812 (N_18812,N_18108,N_18361);
xnor U18813 (N_18813,N_18335,N_18480);
nor U18814 (N_18814,N_18256,N_18202);
nand U18815 (N_18815,N_18296,N_18000);
xor U18816 (N_18816,N_18089,N_18197);
nor U18817 (N_18817,N_18257,N_18275);
or U18818 (N_18818,N_18380,N_18256);
and U18819 (N_18819,N_18262,N_18256);
nor U18820 (N_18820,N_18468,N_18264);
xor U18821 (N_18821,N_18132,N_18006);
and U18822 (N_18822,N_18401,N_18277);
nor U18823 (N_18823,N_18247,N_18475);
xnor U18824 (N_18824,N_18351,N_18089);
nand U18825 (N_18825,N_18442,N_18335);
nand U18826 (N_18826,N_18208,N_18251);
xnor U18827 (N_18827,N_18046,N_18431);
nor U18828 (N_18828,N_18235,N_18435);
nand U18829 (N_18829,N_18136,N_18145);
xnor U18830 (N_18830,N_18462,N_18019);
and U18831 (N_18831,N_18136,N_18079);
and U18832 (N_18832,N_18299,N_18195);
or U18833 (N_18833,N_18400,N_18293);
nand U18834 (N_18834,N_18130,N_18420);
and U18835 (N_18835,N_18083,N_18135);
and U18836 (N_18836,N_18411,N_18070);
nand U18837 (N_18837,N_18058,N_18017);
xnor U18838 (N_18838,N_18010,N_18170);
or U18839 (N_18839,N_18108,N_18058);
xnor U18840 (N_18840,N_18455,N_18294);
xor U18841 (N_18841,N_18270,N_18130);
or U18842 (N_18842,N_18053,N_18035);
xor U18843 (N_18843,N_18457,N_18160);
nand U18844 (N_18844,N_18030,N_18287);
or U18845 (N_18845,N_18479,N_18350);
and U18846 (N_18846,N_18193,N_18289);
nand U18847 (N_18847,N_18122,N_18433);
nand U18848 (N_18848,N_18380,N_18167);
nand U18849 (N_18849,N_18309,N_18386);
nor U18850 (N_18850,N_18412,N_18330);
nor U18851 (N_18851,N_18495,N_18149);
or U18852 (N_18852,N_18435,N_18132);
nor U18853 (N_18853,N_18347,N_18106);
nand U18854 (N_18854,N_18365,N_18051);
and U18855 (N_18855,N_18005,N_18038);
or U18856 (N_18856,N_18194,N_18402);
nand U18857 (N_18857,N_18480,N_18404);
or U18858 (N_18858,N_18374,N_18444);
nand U18859 (N_18859,N_18423,N_18457);
nand U18860 (N_18860,N_18272,N_18315);
xnor U18861 (N_18861,N_18129,N_18100);
nand U18862 (N_18862,N_18247,N_18005);
nand U18863 (N_18863,N_18492,N_18265);
and U18864 (N_18864,N_18400,N_18228);
xnor U18865 (N_18865,N_18122,N_18385);
or U18866 (N_18866,N_18447,N_18263);
or U18867 (N_18867,N_18473,N_18404);
nand U18868 (N_18868,N_18331,N_18460);
and U18869 (N_18869,N_18208,N_18483);
xor U18870 (N_18870,N_18443,N_18012);
or U18871 (N_18871,N_18242,N_18294);
nand U18872 (N_18872,N_18466,N_18282);
or U18873 (N_18873,N_18254,N_18416);
nor U18874 (N_18874,N_18462,N_18143);
nand U18875 (N_18875,N_18324,N_18340);
nor U18876 (N_18876,N_18273,N_18405);
and U18877 (N_18877,N_18018,N_18181);
nand U18878 (N_18878,N_18148,N_18379);
nand U18879 (N_18879,N_18120,N_18297);
and U18880 (N_18880,N_18354,N_18008);
and U18881 (N_18881,N_18249,N_18438);
nand U18882 (N_18882,N_18102,N_18073);
and U18883 (N_18883,N_18425,N_18118);
and U18884 (N_18884,N_18215,N_18293);
nor U18885 (N_18885,N_18227,N_18474);
and U18886 (N_18886,N_18269,N_18251);
xor U18887 (N_18887,N_18343,N_18423);
xnor U18888 (N_18888,N_18268,N_18111);
or U18889 (N_18889,N_18145,N_18221);
xnor U18890 (N_18890,N_18068,N_18095);
nor U18891 (N_18891,N_18366,N_18192);
nand U18892 (N_18892,N_18041,N_18000);
and U18893 (N_18893,N_18467,N_18054);
or U18894 (N_18894,N_18412,N_18415);
and U18895 (N_18895,N_18071,N_18187);
and U18896 (N_18896,N_18061,N_18378);
and U18897 (N_18897,N_18145,N_18019);
xor U18898 (N_18898,N_18338,N_18216);
nor U18899 (N_18899,N_18249,N_18219);
xor U18900 (N_18900,N_18353,N_18460);
xor U18901 (N_18901,N_18280,N_18348);
and U18902 (N_18902,N_18278,N_18409);
and U18903 (N_18903,N_18329,N_18298);
nor U18904 (N_18904,N_18200,N_18127);
nand U18905 (N_18905,N_18467,N_18211);
xor U18906 (N_18906,N_18035,N_18079);
or U18907 (N_18907,N_18286,N_18198);
nand U18908 (N_18908,N_18413,N_18095);
xnor U18909 (N_18909,N_18021,N_18458);
nor U18910 (N_18910,N_18334,N_18244);
and U18911 (N_18911,N_18127,N_18404);
xor U18912 (N_18912,N_18209,N_18036);
or U18913 (N_18913,N_18298,N_18192);
or U18914 (N_18914,N_18048,N_18263);
and U18915 (N_18915,N_18308,N_18419);
and U18916 (N_18916,N_18255,N_18248);
or U18917 (N_18917,N_18379,N_18437);
xnor U18918 (N_18918,N_18299,N_18047);
nor U18919 (N_18919,N_18203,N_18092);
and U18920 (N_18920,N_18137,N_18202);
or U18921 (N_18921,N_18406,N_18112);
nand U18922 (N_18922,N_18184,N_18422);
xor U18923 (N_18923,N_18171,N_18449);
xnor U18924 (N_18924,N_18290,N_18266);
nor U18925 (N_18925,N_18060,N_18307);
or U18926 (N_18926,N_18097,N_18053);
nor U18927 (N_18927,N_18105,N_18395);
and U18928 (N_18928,N_18262,N_18340);
nor U18929 (N_18929,N_18423,N_18024);
or U18930 (N_18930,N_18009,N_18285);
and U18931 (N_18931,N_18448,N_18243);
nor U18932 (N_18932,N_18330,N_18186);
nand U18933 (N_18933,N_18462,N_18447);
and U18934 (N_18934,N_18401,N_18278);
nand U18935 (N_18935,N_18105,N_18317);
or U18936 (N_18936,N_18130,N_18179);
nand U18937 (N_18937,N_18127,N_18222);
nor U18938 (N_18938,N_18237,N_18092);
nand U18939 (N_18939,N_18428,N_18398);
or U18940 (N_18940,N_18306,N_18304);
nand U18941 (N_18941,N_18383,N_18397);
xnor U18942 (N_18942,N_18405,N_18128);
nand U18943 (N_18943,N_18472,N_18222);
xor U18944 (N_18944,N_18004,N_18170);
nand U18945 (N_18945,N_18017,N_18240);
or U18946 (N_18946,N_18201,N_18118);
xor U18947 (N_18947,N_18117,N_18400);
nor U18948 (N_18948,N_18104,N_18249);
nand U18949 (N_18949,N_18480,N_18076);
xnor U18950 (N_18950,N_18287,N_18456);
nand U18951 (N_18951,N_18321,N_18159);
nand U18952 (N_18952,N_18156,N_18486);
or U18953 (N_18953,N_18385,N_18417);
nand U18954 (N_18954,N_18371,N_18378);
or U18955 (N_18955,N_18114,N_18388);
or U18956 (N_18956,N_18488,N_18393);
or U18957 (N_18957,N_18244,N_18040);
or U18958 (N_18958,N_18059,N_18053);
xor U18959 (N_18959,N_18427,N_18112);
and U18960 (N_18960,N_18026,N_18447);
nor U18961 (N_18961,N_18341,N_18483);
xor U18962 (N_18962,N_18428,N_18140);
nand U18963 (N_18963,N_18046,N_18209);
and U18964 (N_18964,N_18419,N_18107);
or U18965 (N_18965,N_18071,N_18197);
xor U18966 (N_18966,N_18303,N_18112);
xor U18967 (N_18967,N_18480,N_18478);
xnor U18968 (N_18968,N_18062,N_18116);
and U18969 (N_18969,N_18018,N_18482);
nand U18970 (N_18970,N_18146,N_18267);
or U18971 (N_18971,N_18124,N_18487);
or U18972 (N_18972,N_18299,N_18043);
and U18973 (N_18973,N_18024,N_18266);
and U18974 (N_18974,N_18004,N_18244);
xnor U18975 (N_18975,N_18489,N_18496);
xnor U18976 (N_18976,N_18037,N_18040);
nand U18977 (N_18977,N_18166,N_18265);
and U18978 (N_18978,N_18206,N_18434);
or U18979 (N_18979,N_18128,N_18050);
nand U18980 (N_18980,N_18273,N_18055);
and U18981 (N_18981,N_18171,N_18447);
and U18982 (N_18982,N_18313,N_18273);
and U18983 (N_18983,N_18352,N_18224);
xnor U18984 (N_18984,N_18449,N_18152);
nand U18985 (N_18985,N_18330,N_18324);
xnor U18986 (N_18986,N_18006,N_18073);
or U18987 (N_18987,N_18080,N_18204);
and U18988 (N_18988,N_18069,N_18456);
xor U18989 (N_18989,N_18260,N_18284);
or U18990 (N_18990,N_18107,N_18403);
and U18991 (N_18991,N_18320,N_18182);
nor U18992 (N_18992,N_18302,N_18216);
xor U18993 (N_18993,N_18003,N_18092);
and U18994 (N_18994,N_18095,N_18113);
nand U18995 (N_18995,N_18219,N_18109);
nor U18996 (N_18996,N_18117,N_18031);
xnor U18997 (N_18997,N_18009,N_18430);
nor U18998 (N_18998,N_18294,N_18063);
nor U18999 (N_18999,N_18045,N_18143);
nand U19000 (N_19000,N_18788,N_18831);
nor U19001 (N_19001,N_18514,N_18961);
nor U19002 (N_19002,N_18992,N_18977);
or U19003 (N_19003,N_18872,N_18569);
or U19004 (N_19004,N_18882,N_18713);
and U19005 (N_19005,N_18669,N_18628);
xnor U19006 (N_19006,N_18832,N_18829);
nand U19007 (N_19007,N_18976,N_18627);
nand U19008 (N_19008,N_18813,N_18674);
nand U19009 (N_19009,N_18880,N_18658);
xnor U19010 (N_19010,N_18620,N_18906);
and U19011 (N_19011,N_18915,N_18913);
or U19012 (N_19012,N_18608,N_18954);
xnor U19013 (N_19013,N_18546,N_18556);
xnor U19014 (N_19014,N_18517,N_18667);
and U19015 (N_19015,N_18771,N_18607);
nand U19016 (N_19016,N_18874,N_18663);
nand U19017 (N_19017,N_18951,N_18903);
xor U19018 (N_19018,N_18854,N_18626);
xor U19019 (N_19019,N_18821,N_18591);
or U19020 (N_19020,N_18834,N_18726);
nor U19021 (N_19021,N_18935,N_18602);
or U19022 (N_19022,N_18752,N_18792);
or U19023 (N_19023,N_18579,N_18531);
or U19024 (N_19024,N_18775,N_18745);
xor U19025 (N_19025,N_18601,N_18853);
or U19026 (N_19026,N_18810,N_18852);
nor U19027 (N_19027,N_18860,N_18805);
or U19028 (N_19028,N_18555,N_18549);
nand U19029 (N_19029,N_18523,N_18635);
nand U19030 (N_19030,N_18707,N_18962);
and U19031 (N_19031,N_18868,N_18532);
nand U19032 (N_19032,N_18550,N_18947);
nand U19033 (N_19033,N_18747,N_18789);
and U19034 (N_19034,N_18925,N_18917);
nand U19035 (N_19035,N_18650,N_18864);
nand U19036 (N_19036,N_18583,N_18916);
nand U19037 (N_19037,N_18898,N_18883);
nor U19038 (N_19038,N_18763,N_18630);
nand U19039 (N_19039,N_18993,N_18575);
or U19040 (N_19040,N_18536,N_18886);
xor U19041 (N_19041,N_18758,N_18899);
xnor U19042 (N_19042,N_18670,N_18735);
nor U19043 (N_19043,N_18595,N_18980);
xnor U19044 (N_19044,N_18599,N_18557);
or U19045 (N_19045,N_18999,N_18772);
nand U19046 (N_19046,N_18900,N_18818);
xor U19047 (N_19047,N_18957,N_18969);
and U19048 (N_19048,N_18732,N_18625);
or U19049 (N_19049,N_18875,N_18610);
or U19050 (N_19050,N_18580,N_18837);
nor U19051 (N_19051,N_18901,N_18764);
xnor U19052 (N_19052,N_18553,N_18985);
and U19053 (N_19053,N_18811,N_18799);
or U19054 (N_19054,N_18582,N_18940);
nand U19055 (N_19055,N_18982,N_18693);
nor U19056 (N_19056,N_18702,N_18933);
nand U19057 (N_19057,N_18688,N_18604);
nor U19058 (N_19058,N_18912,N_18621);
and U19059 (N_19059,N_18928,N_18681);
xnor U19060 (N_19060,N_18790,N_18807);
and U19061 (N_19061,N_18718,N_18785);
or U19062 (N_19062,N_18716,N_18644);
or U19063 (N_19063,N_18664,N_18887);
and U19064 (N_19064,N_18585,N_18709);
xnor U19065 (N_19065,N_18861,N_18510);
xnor U19066 (N_19066,N_18544,N_18683);
or U19067 (N_19067,N_18939,N_18565);
nand U19068 (N_19068,N_18808,N_18629);
nand U19069 (N_19069,N_18509,N_18761);
nor U19070 (N_19070,N_18522,N_18938);
xor U19071 (N_19071,N_18835,N_18960);
nor U19072 (N_19072,N_18855,N_18513);
xnor U19073 (N_19073,N_18678,N_18572);
xnor U19074 (N_19074,N_18816,N_18826);
xor U19075 (N_19075,N_18934,N_18979);
nand U19076 (N_19076,N_18742,N_18843);
and U19077 (N_19077,N_18526,N_18698);
or U19078 (N_19078,N_18654,N_18609);
or U19079 (N_19079,N_18779,N_18998);
nor U19080 (N_19080,N_18701,N_18756);
or U19081 (N_19081,N_18668,N_18974);
nand U19082 (N_19082,N_18511,N_18639);
nor U19083 (N_19083,N_18722,N_18566);
and U19084 (N_19084,N_18520,N_18770);
or U19085 (N_19085,N_18944,N_18636);
nand U19086 (N_19086,N_18721,N_18729);
and U19087 (N_19087,N_18649,N_18840);
nor U19088 (N_19088,N_18795,N_18867);
or U19089 (N_19089,N_18802,N_18577);
xor U19090 (N_19090,N_18652,N_18885);
xor U19091 (N_19091,N_18727,N_18893);
or U19092 (N_19092,N_18749,N_18551);
or U19093 (N_19093,N_18911,N_18907);
nor U19094 (N_19094,N_18945,N_18989);
and U19095 (N_19095,N_18878,N_18733);
nand U19096 (N_19096,N_18830,N_18598);
nor U19097 (N_19097,N_18528,N_18997);
xnor U19098 (N_19098,N_18755,N_18844);
or U19099 (N_19099,N_18869,N_18936);
xnor U19100 (N_19100,N_18593,N_18919);
nor U19101 (N_19101,N_18995,N_18814);
nand U19102 (N_19102,N_18508,N_18615);
nor U19103 (N_19103,N_18684,N_18967);
nand U19104 (N_19104,N_18923,N_18632);
nor U19105 (N_19105,N_18804,N_18502);
xnor U19106 (N_19106,N_18687,N_18700);
nor U19107 (N_19107,N_18952,N_18503);
nand U19108 (N_19108,N_18803,N_18791);
and U19109 (N_19109,N_18847,N_18894);
nand U19110 (N_19110,N_18856,N_18827);
nand U19111 (N_19111,N_18798,N_18611);
xor U19112 (N_19112,N_18578,N_18706);
nand U19113 (N_19113,N_18760,N_18736);
nor U19114 (N_19114,N_18889,N_18981);
nand U19115 (N_19115,N_18955,N_18676);
and U19116 (N_19116,N_18638,N_18527);
and U19117 (N_19117,N_18746,N_18783);
nor U19118 (N_19118,N_18589,N_18504);
nand U19119 (N_19119,N_18571,N_18624);
xnor U19120 (N_19120,N_18581,N_18806);
nor U19121 (N_19121,N_18765,N_18574);
nor U19122 (N_19122,N_18970,N_18622);
xnor U19123 (N_19123,N_18708,N_18588);
or U19124 (N_19124,N_18710,N_18542);
and U19125 (N_19125,N_18680,N_18535);
xor U19126 (N_19126,N_18929,N_18930);
nand U19127 (N_19127,N_18846,N_18948);
and U19128 (N_19128,N_18812,N_18543);
or U19129 (N_19129,N_18988,N_18618);
nand U19130 (N_19130,N_18876,N_18741);
nand U19131 (N_19131,N_18796,N_18673);
nor U19132 (N_19132,N_18540,N_18932);
nand U19133 (N_19133,N_18659,N_18686);
nor U19134 (N_19134,N_18605,N_18506);
or U19135 (N_19135,N_18822,N_18538);
and U19136 (N_19136,N_18515,N_18877);
nor U19137 (N_19137,N_18922,N_18845);
and U19138 (N_19138,N_18753,N_18768);
or U19139 (N_19139,N_18613,N_18897);
xnor U19140 (N_19140,N_18776,N_18920);
and U19141 (N_19141,N_18634,N_18778);
nand U19142 (N_19142,N_18672,N_18567);
and U19143 (N_19143,N_18773,N_18524);
nand U19144 (N_19144,N_18757,N_18914);
nand U19145 (N_19145,N_18507,N_18850);
and U19146 (N_19146,N_18744,N_18541);
or U19147 (N_19147,N_18560,N_18941);
or U19148 (N_19148,N_18576,N_18682);
nor U19149 (N_19149,N_18884,N_18691);
nand U19150 (N_19150,N_18724,N_18539);
and U19151 (N_19151,N_18623,N_18817);
nand U19152 (N_19152,N_18642,N_18751);
and U19153 (N_19153,N_18963,N_18848);
and U19154 (N_19154,N_18612,N_18921);
and U19155 (N_19155,N_18660,N_18740);
xor U19156 (N_19156,N_18743,N_18694);
xor U19157 (N_19157,N_18833,N_18987);
nor U19158 (N_19158,N_18501,N_18841);
and U19159 (N_19159,N_18533,N_18679);
nand U19160 (N_19160,N_18782,N_18849);
and U19161 (N_19161,N_18759,N_18866);
nor U19162 (N_19162,N_18685,N_18748);
nand U19163 (N_19163,N_18728,N_18704);
or U19164 (N_19164,N_18570,N_18797);
nor U19165 (N_19165,N_18534,N_18888);
nand U19166 (N_19166,N_18881,N_18675);
and U19167 (N_19167,N_18950,N_18586);
nor U19168 (N_19168,N_18842,N_18926);
xor U19169 (N_19169,N_18892,N_18971);
nor U19170 (N_19170,N_18953,N_18645);
nor U19171 (N_19171,N_18737,N_18879);
xor U19172 (N_19172,N_18958,N_18870);
or U19173 (N_19173,N_18712,N_18548);
or U19174 (N_19174,N_18851,N_18895);
nor U19175 (N_19175,N_18859,N_18653);
and U19176 (N_19176,N_18697,N_18978);
nand U19177 (N_19177,N_18774,N_18552);
or U19178 (N_19178,N_18873,N_18937);
and U19179 (N_19179,N_18717,N_18705);
and U19180 (N_19180,N_18631,N_18619);
xor U19181 (N_19181,N_18656,N_18890);
and U19182 (N_19182,N_18564,N_18643);
xor U19183 (N_19183,N_18828,N_18975);
nor U19184 (N_19184,N_18908,N_18857);
or U19185 (N_19185,N_18924,N_18910);
or U19186 (N_19186,N_18730,N_18714);
nor U19187 (N_19187,N_18616,N_18902);
and U19188 (N_19188,N_18784,N_18562);
or U19189 (N_19189,N_18597,N_18633);
or U19190 (N_19190,N_18786,N_18594);
or U19191 (N_19191,N_18767,N_18862);
or U19192 (N_19192,N_18972,N_18896);
and U19193 (N_19193,N_18500,N_18968);
xnor U19194 (N_19194,N_18655,N_18647);
xnor U19195 (N_19195,N_18777,N_18991);
nor U19196 (N_19196,N_18815,N_18587);
or U19197 (N_19197,N_18769,N_18545);
and U19198 (N_19198,N_18561,N_18927);
nor U19199 (N_19199,N_18909,N_18819);
and U19200 (N_19200,N_18603,N_18606);
or U19201 (N_19201,N_18711,N_18671);
nand U19202 (N_19202,N_18525,N_18512);
and U19203 (N_19203,N_18568,N_18648);
and U19204 (N_19204,N_18738,N_18600);
and U19205 (N_19205,N_18690,N_18946);
xnor U19206 (N_19206,N_18666,N_18838);
or U19207 (N_19207,N_18554,N_18518);
xnor U19208 (N_19208,N_18662,N_18965);
or U19209 (N_19209,N_18699,N_18537);
or U19210 (N_19210,N_18596,N_18959);
nand U19211 (N_19211,N_18665,N_18590);
nand U19212 (N_19212,N_18530,N_18731);
and U19213 (N_19213,N_18966,N_18996);
xor U19214 (N_19214,N_18956,N_18592);
nor U19215 (N_19215,N_18904,N_18719);
nor U19216 (N_19216,N_18505,N_18794);
or U19217 (N_19217,N_18547,N_18984);
xor U19218 (N_19218,N_18725,N_18766);
and U19219 (N_19219,N_18865,N_18825);
nand U19220 (N_19220,N_18820,N_18931);
nor U19221 (N_19221,N_18780,N_18871);
xnor U19222 (N_19222,N_18836,N_18646);
or U19223 (N_19223,N_18703,N_18824);
or U19224 (N_19224,N_18762,N_18516);
nand U19225 (N_19225,N_18734,N_18529);
or U19226 (N_19226,N_18823,N_18715);
or U19227 (N_19227,N_18614,N_18781);
nand U19228 (N_19228,N_18750,N_18793);
xor U19229 (N_19229,N_18990,N_18640);
nand U19230 (N_19230,N_18994,N_18573);
or U19231 (N_19231,N_18986,N_18809);
xnor U19232 (N_19232,N_18964,N_18787);
xnor U19233 (N_19233,N_18973,N_18918);
nor U19234 (N_19234,N_18720,N_18695);
xnor U19235 (N_19235,N_18863,N_18739);
nor U19236 (N_19236,N_18858,N_18651);
nor U19237 (N_19237,N_18641,N_18559);
and U19238 (N_19238,N_18942,N_18521);
or U19239 (N_19239,N_18949,N_18563);
and U19240 (N_19240,N_18696,N_18905);
and U19241 (N_19241,N_18723,N_18617);
nor U19242 (N_19242,N_18519,N_18801);
nand U19243 (N_19243,N_18661,N_18657);
nor U19244 (N_19244,N_18558,N_18637);
xnor U19245 (N_19245,N_18689,N_18677);
and U19246 (N_19246,N_18943,N_18983);
nand U19247 (N_19247,N_18891,N_18800);
or U19248 (N_19248,N_18584,N_18754);
and U19249 (N_19249,N_18839,N_18692);
or U19250 (N_19250,N_18815,N_18772);
nor U19251 (N_19251,N_18591,N_18943);
xnor U19252 (N_19252,N_18606,N_18514);
nor U19253 (N_19253,N_18592,N_18815);
and U19254 (N_19254,N_18509,N_18965);
nor U19255 (N_19255,N_18931,N_18537);
nand U19256 (N_19256,N_18535,N_18537);
nand U19257 (N_19257,N_18898,N_18686);
and U19258 (N_19258,N_18512,N_18757);
nand U19259 (N_19259,N_18668,N_18521);
and U19260 (N_19260,N_18996,N_18906);
nand U19261 (N_19261,N_18757,N_18819);
or U19262 (N_19262,N_18552,N_18620);
nand U19263 (N_19263,N_18534,N_18833);
and U19264 (N_19264,N_18595,N_18658);
nand U19265 (N_19265,N_18814,N_18671);
nand U19266 (N_19266,N_18945,N_18583);
or U19267 (N_19267,N_18844,N_18876);
nand U19268 (N_19268,N_18547,N_18542);
or U19269 (N_19269,N_18797,N_18596);
xnor U19270 (N_19270,N_18707,N_18765);
nor U19271 (N_19271,N_18626,N_18597);
nor U19272 (N_19272,N_18659,N_18842);
nand U19273 (N_19273,N_18798,N_18801);
xor U19274 (N_19274,N_18919,N_18543);
nand U19275 (N_19275,N_18795,N_18615);
and U19276 (N_19276,N_18748,N_18899);
or U19277 (N_19277,N_18705,N_18904);
xor U19278 (N_19278,N_18867,N_18536);
nor U19279 (N_19279,N_18513,N_18529);
xor U19280 (N_19280,N_18984,N_18669);
nor U19281 (N_19281,N_18665,N_18743);
or U19282 (N_19282,N_18810,N_18561);
or U19283 (N_19283,N_18542,N_18502);
or U19284 (N_19284,N_18804,N_18874);
and U19285 (N_19285,N_18778,N_18503);
and U19286 (N_19286,N_18592,N_18934);
xnor U19287 (N_19287,N_18982,N_18639);
or U19288 (N_19288,N_18544,N_18565);
nand U19289 (N_19289,N_18772,N_18654);
nor U19290 (N_19290,N_18879,N_18921);
xnor U19291 (N_19291,N_18808,N_18919);
and U19292 (N_19292,N_18647,N_18601);
or U19293 (N_19293,N_18836,N_18995);
nor U19294 (N_19294,N_18985,N_18571);
nor U19295 (N_19295,N_18545,N_18514);
xnor U19296 (N_19296,N_18558,N_18795);
or U19297 (N_19297,N_18926,N_18561);
nand U19298 (N_19298,N_18705,N_18757);
nand U19299 (N_19299,N_18696,N_18560);
and U19300 (N_19300,N_18918,N_18986);
nand U19301 (N_19301,N_18867,N_18809);
nor U19302 (N_19302,N_18595,N_18984);
and U19303 (N_19303,N_18978,N_18996);
nand U19304 (N_19304,N_18851,N_18523);
nor U19305 (N_19305,N_18948,N_18523);
nand U19306 (N_19306,N_18595,N_18787);
and U19307 (N_19307,N_18597,N_18954);
or U19308 (N_19308,N_18817,N_18936);
or U19309 (N_19309,N_18786,N_18898);
or U19310 (N_19310,N_18698,N_18971);
nand U19311 (N_19311,N_18934,N_18581);
nor U19312 (N_19312,N_18731,N_18776);
nor U19313 (N_19313,N_18743,N_18575);
or U19314 (N_19314,N_18747,N_18637);
nor U19315 (N_19315,N_18570,N_18650);
xnor U19316 (N_19316,N_18685,N_18647);
and U19317 (N_19317,N_18827,N_18957);
or U19318 (N_19318,N_18927,N_18677);
nor U19319 (N_19319,N_18935,N_18897);
xor U19320 (N_19320,N_18500,N_18877);
or U19321 (N_19321,N_18656,N_18927);
and U19322 (N_19322,N_18651,N_18539);
xor U19323 (N_19323,N_18771,N_18709);
and U19324 (N_19324,N_18611,N_18776);
nor U19325 (N_19325,N_18804,N_18980);
or U19326 (N_19326,N_18513,N_18669);
nand U19327 (N_19327,N_18501,N_18859);
and U19328 (N_19328,N_18618,N_18763);
nor U19329 (N_19329,N_18673,N_18552);
nor U19330 (N_19330,N_18603,N_18643);
or U19331 (N_19331,N_18944,N_18885);
xor U19332 (N_19332,N_18550,N_18712);
nand U19333 (N_19333,N_18664,N_18677);
xor U19334 (N_19334,N_18657,N_18813);
or U19335 (N_19335,N_18639,N_18520);
and U19336 (N_19336,N_18590,N_18761);
xor U19337 (N_19337,N_18650,N_18723);
xnor U19338 (N_19338,N_18963,N_18581);
and U19339 (N_19339,N_18804,N_18865);
xor U19340 (N_19340,N_18510,N_18765);
or U19341 (N_19341,N_18659,N_18827);
nand U19342 (N_19342,N_18724,N_18821);
xnor U19343 (N_19343,N_18513,N_18545);
or U19344 (N_19344,N_18604,N_18683);
nand U19345 (N_19345,N_18914,N_18886);
xor U19346 (N_19346,N_18912,N_18850);
nor U19347 (N_19347,N_18680,N_18851);
nor U19348 (N_19348,N_18680,N_18540);
nand U19349 (N_19349,N_18800,N_18755);
nor U19350 (N_19350,N_18506,N_18845);
nor U19351 (N_19351,N_18663,N_18889);
nor U19352 (N_19352,N_18683,N_18771);
xor U19353 (N_19353,N_18814,N_18616);
nand U19354 (N_19354,N_18976,N_18665);
nand U19355 (N_19355,N_18905,N_18774);
nor U19356 (N_19356,N_18997,N_18890);
or U19357 (N_19357,N_18829,N_18719);
and U19358 (N_19358,N_18901,N_18829);
xor U19359 (N_19359,N_18668,N_18877);
xnor U19360 (N_19360,N_18658,N_18500);
nor U19361 (N_19361,N_18746,N_18688);
nand U19362 (N_19362,N_18695,N_18629);
and U19363 (N_19363,N_18842,N_18748);
nand U19364 (N_19364,N_18730,N_18622);
nand U19365 (N_19365,N_18640,N_18980);
xnor U19366 (N_19366,N_18550,N_18993);
nand U19367 (N_19367,N_18689,N_18664);
and U19368 (N_19368,N_18978,N_18769);
xor U19369 (N_19369,N_18599,N_18555);
and U19370 (N_19370,N_18986,N_18690);
or U19371 (N_19371,N_18659,N_18840);
and U19372 (N_19372,N_18917,N_18568);
nor U19373 (N_19373,N_18590,N_18699);
nand U19374 (N_19374,N_18513,N_18917);
xor U19375 (N_19375,N_18532,N_18641);
nor U19376 (N_19376,N_18925,N_18822);
or U19377 (N_19377,N_18665,N_18795);
nor U19378 (N_19378,N_18533,N_18538);
xnor U19379 (N_19379,N_18869,N_18691);
or U19380 (N_19380,N_18526,N_18702);
nor U19381 (N_19381,N_18994,N_18895);
or U19382 (N_19382,N_18589,N_18736);
and U19383 (N_19383,N_18906,N_18961);
or U19384 (N_19384,N_18580,N_18925);
or U19385 (N_19385,N_18823,N_18643);
nand U19386 (N_19386,N_18630,N_18533);
nand U19387 (N_19387,N_18668,N_18816);
xor U19388 (N_19388,N_18676,N_18878);
nor U19389 (N_19389,N_18924,N_18755);
nor U19390 (N_19390,N_18523,N_18751);
and U19391 (N_19391,N_18820,N_18923);
or U19392 (N_19392,N_18947,N_18508);
or U19393 (N_19393,N_18625,N_18592);
and U19394 (N_19394,N_18894,N_18726);
nand U19395 (N_19395,N_18897,N_18833);
or U19396 (N_19396,N_18982,N_18515);
nand U19397 (N_19397,N_18897,N_18534);
nand U19398 (N_19398,N_18534,N_18975);
and U19399 (N_19399,N_18982,N_18827);
or U19400 (N_19400,N_18566,N_18931);
and U19401 (N_19401,N_18981,N_18918);
and U19402 (N_19402,N_18553,N_18587);
or U19403 (N_19403,N_18919,N_18560);
xor U19404 (N_19404,N_18616,N_18632);
or U19405 (N_19405,N_18936,N_18852);
nand U19406 (N_19406,N_18961,N_18875);
nor U19407 (N_19407,N_18653,N_18983);
xor U19408 (N_19408,N_18991,N_18676);
xor U19409 (N_19409,N_18781,N_18825);
xnor U19410 (N_19410,N_18713,N_18760);
and U19411 (N_19411,N_18668,N_18651);
and U19412 (N_19412,N_18549,N_18863);
nand U19413 (N_19413,N_18574,N_18701);
or U19414 (N_19414,N_18535,N_18541);
nor U19415 (N_19415,N_18571,N_18609);
nand U19416 (N_19416,N_18938,N_18849);
xor U19417 (N_19417,N_18722,N_18747);
or U19418 (N_19418,N_18523,N_18872);
nand U19419 (N_19419,N_18917,N_18762);
and U19420 (N_19420,N_18973,N_18871);
and U19421 (N_19421,N_18670,N_18625);
and U19422 (N_19422,N_18958,N_18824);
nand U19423 (N_19423,N_18779,N_18604);
nand U19424 (N_19424,N_18634,N_18867);
or U19425 (N_19425,N_18533,N_18544);
nor U19426 (N_19426,N_18706,N_18798);
xor U19427 (N_19427,N_18865,N_18916);
and U19428 (N_19428,N_18524,N_18586);
or U19429 (N_19429,N_18541,N_18878);
xnor U19430 (N_19430,N_18788,N_18754);
nand U19431 (N_19431,N_18792,N_18652);
xor U19432 (N_19432,N_18953,N_18557);
xnor U19433 (N_19433,N_18982,N_18921);
nand U19434 (N_19434,N_18567,N_18670);
nand U19435 (N_19435,N_18557,N_18526);
nor U19436 (N_19436,N_18861,N_18814);
nor U19437 (N_19437,N_18880,N_18943);
or U19438 (N_19438,N_18843,N_18548);
or U19439 (N_19439,N_18771,N_18747);
nand U19440 (N_19440,N_18665,N_18820);
or U19441 (N_19441,N_18827,N_18675);
nor U19442 (N_19442,N_18794,N_18641);
nand U19443 (N_19443,N_18745,N_18853);
or U19444 (N_19444,N_18675,N_18992);
or U19445 (N_19445,N_18830,N_18539);
xor U19446 (N_19446,N_18772,N_18652);
and U19447 (N_19447,N_18931,N_18904);
or U19448 (N_19448,N_18927,N_18761);
xnor U19449 (N_19449,N_18583,N_18873);
nor U19450 (N_19450,N_18979,N_18858);
and U19451 (N_19451,N_18868,N_18668);
nor U19452 (N_19452,N_18796,N_18679);
nor U19453 (N_19453,N_18756,N_18629);
nand U19454 (N_19454,N_18632,N_18794);
or U19455 (N_19455,N_18967,N_18572);
or U19456 (N_19456,N_18643,N_18757);
xnor U19457 (N_19457,N_18994,N_18633);
or U19458 (N_19458,N_18817,N_18931);
or U19459 (N_19459,N_18744,N_18546);
xor U19460 (N_19460,N_18678,N_18705);
or U19461 (N_19461,N_18827,N_18837);
or U19462 (N_19462,N_18742,N_18880);
and U19463 (N_19463,N_18976,N_18532);
xnor U19464 (N_19464,N_18976,N_18737);
nand U19465 (N_19465,N_18557,N_18715);
xnor U19466 (N_19466,N_18717,N_18698);
and U19467 (N_19467,N_18828,N_18538);
xor U19468 (N_19468,N_18778,N_18748);
nor U19469 (N_19469,N_18529,N_18939);
and U19470 (N_19470,N_18861,N_18657);
or U19471 (N_19471,N_18948,N_18534);
and U19472 (N_19472,N_18770,N_18771);
or U19473 (N_19473,N_18606,N_18504);
nand U19474 (N_19474,N_18556,N_18791);
nor U19475 (N_19475,N_18953,N_18651);
nor U19476 (N_19476,N_18635,N_18700);
or U19477 (N_19477,N_18900,N_18509);
or U19478 (N_19478,N_18802,N_18933);
and U19479 (N_19479,N_18710,N_18594);
or U19480 (N_19480,N_18854,N_18597);
xnor U19481 (N_19481,N_18858,N_18530);
xor U19482 (N_19482,N_18709,N_18545);
nand U19483 (N_19483,N_18590,N_18960);
or U19484 (N_19484,N_18951,N_18935);
nor U19485 (N_19485,N_18825,N_18587);
nor U19486 (N_19486,N_18834,N_18839);
or U19487 (N_19487,N_18981,N_18868);
nor U19488 (N_19488,N_18949,N_18955);
and U19489 (N_19489,N_18705,N_18575);
and U19490 (N_19490,N_18593,N_18841);
or U19491 (N_19491,N_18874,N_18946);
or U19492 (N_19492,N_18936,N_18919);
xor U19493 (N_19493,N_18957,N_18693);
or U19494 (N_19494,N_18843,N_18641);
nand U19495 (N_19495,N_18530,N_18914);
or U19496 (N_19496,N_18527,N_18528);
or U19497 (N_19497,N_18937,N_18788);
xor U19498 (N_19498,N_18854,N_18524);
xor U19499 (N_19499,N_18994,N_18710);
xnor U19500 (N_19500,N_19363,N_19259);
xor U19501 (N_19501,N_19273,N_19257);
nor U19502 (N_19502,N_19166,N_19222);
nor U19503 (N_19503,N_19148,N_19024);
xor U19504 (N_19504,N_19250,N_19214);
xnor U19505 (N_19505,N_19204,N_19489);
nor U19506 (N_19506,N_19415,N_19416);
nor U19507 (N_19507,N_19288,N_19099);
nor U19508 (N_19508,N_19106,N_19201);
or U19509 (N_19509,N_19015,N_19296);
xor U19510 (N_19510,N_19134,N_19058);
or U19511 (N_19511,N_19388,N_19062);
and U19512 (N_19512,N_19269,N_19498);
or U19513 (N_19513,N_19030,N_19367);
or U19514 (N_19514,N_19037,N_19258);
nand U19515 (N_19515,N_19235,N_19104);
nor U19516 (N_19516,N_19292,N_19084);
and U19517 (N_19517,N_19274,N_19365);
nor U19518 (N_19518,N_19179,N_19494);
nand U19519 (N_19519,N_19353,N_19404);
or U19520 (N_19520,N_19120,N_19387);
or U19521 (N_19521,N_19013,N_19185);
and U19522 (N_19522,N_19420,N_19176);
xnor U19523 (N_19523,N_19069,N_19169);
nor U19524 (N_19524,N_19117,N_19244);
or U19525 (N_19525,N_19121,N_19209);
xor U19526 (N_19526,N_19054,N_19101);
and U19527 (N_19527,N_19380,N_19397);
or U19528 (N_19528,N_19364,N_19177);
xor U19529 (N_19529,N_19391,N_19399);
or U19530 (N_19530,N_19187,N_19394);
nand U19531 (N_19531,N_19412,N_19402);
xnor U19532 (N_19532,N_19163,N_19303);
nor U19533 (N_19533,N_19432,N_19389);
xnor U19534 (N_19534,N_19170,N_19252);
nor U19535 (N_19535,N_19261,N_19354);
nand U19536 (N_19536,N_19322,N_19267);
nand U19537 (N_19537,N_19345,N_19211);
nor U19538 (N_19538,N_19039,N_19038);
xnor U19539 (N_19539,N_19338,N_19183);
nand U19540 (N_19540,N_19255,N_19167);
xnor U19541 (N_19541,N_19196,N_19295);
and U19542 (N_19542,N_19074,N_19301);
or U19543 (N_19543,N_19458,N_19475);
nor U19544 (N_19544,N_19012,N_19279);
and U19545 (N_19545,N_19122,N_19119);
or U19546 (N_19546,N_19061,N_19236);
nand U19547 (N_19547,N_19348,N_19092);
nand U19548 (N_19548,N_19063,N_19499);
xor U19549 (N_19549,N_19493,N_19290);
nand U19550 (N_19550,N_19421,N_19194);
and U19551 (N_19551,N_19327,N_19492);
or U19552 (N_19552,N_19316,N_19103);
xnor U19553 (N_19553,N_19243,N_19145);
nand U19554 (N_19554,N_19151,N_19060);
or U19555 (N_19555,N_19464,N_19487);
or U19556 (N_19556,N_19359,N_19133);
xnor U19557 (N_19557,N_19197,N_19232);
xor U19558 (N_19558,N_19112,N_19278);
nor U19559 (N_19559,N_19118,N_19337);
and U19560 (N_19560,N_19124,N_19025);
nor U19561 (N_19561,N_19346,N_19116);
or U19562 (N_19562,N_19158,N_19430);
or U19563 (N_19563,N_19254,N_19020);
nor U19564 (N_19564,N_19484,N_19126);
nor U19565 (N_19565,N_19351,N_19154);
and U19566 (N_19566,N_19050,N_19335);
nor U19567 (N_19567,N_19272,N_19263);
nor U19568 (N_19568,N_19479,N_19083);
nor U19569 (N_19569,N_19444,N_19073);
xor U19570 (N_19570,N_19468,N_19419);
and U19571 (N_19571,N_19390,N_19241);
and U19572 (N_19572,N_19311,N_19052);
nor U19573 (N_19573,N_19018,N_19182);
xor U19574 (N_19574,N_19178,N_19193);
xor U19575 (N_19575,N_19071,N_19300);
nand U19576 (N_19576,N_19482,N_19195);
xnor U19577 (N_19577,N_19008,N_19028);
or U19578 (N_19578,N_19342,N_19481);
nor U19579 (N_19579,N_19023,N_19281);
nor U19580 (N_19580,N_19417,N_19109);
nor U19581 (N_19581,N_19105,N_19141);
nand U19582 (N_19582,N_19143,N_19299);
and U19583 (N_19583,N_19051,N_19010);
nand U19584 (N_19584,N_19239,N_19245);
or U19585 (N_19585,N_19005,N_19251);
and U19586 (N_19586,N_19307,N_19040);
nor U19587 (N_19587,N_19032,N_19089);
xnor U19588 (N_19588,N_19072,N_19057);
nor U19589 (N_19589,N_19159,N_19473);
xor U19590 (N_19590,N_19205,N_19107);
and U19591 (N_19591,N_19045,N_19344);
xnor U19592 (N_19592,N_19217,N_19441);
nand U19593 (N_19593,N_19293,N_19006);
and U19594 (N_19594,N_19375,N_19044);
nor U19595 (N_19595,N_19377,N_19142);
nor U19596 (N_19596,N_19082,N_19139);
or U19597 (N_19597,N_19004,N_19264);
nor U19598 (N_19598,N_19123,N_19437);
nor U19599 (N_19599,N_19445,N_19047);
and U19600 (N_19600,N_19396,N_19407);
or U19601 (N_19601,N_19488,N_19280);
or U19602 (N_19602,N_19036,N_19406);
or U19603 (N_19603,N_19312,N_19393);
nor U19604 (N_19604,N_19284,N_19373);
xor U19605 (N_19605,N_19248,N_19450);
nor U19606 (N_19606,N_19231,N_19276);
xor U19607 (N_19607,N_19137,N_19426);
nor U19608 (N_19608,N_19080,N_19224);
nand U19609 (N_19609,N_19483,N_19368);
or U19610 (N_19610,N_19305,N_19331);
nor U19611 (N_19611,N_19277,N_19165);
xnor U19612 (N_19612,N_19429,N_19199);
and U19613 (N_19613,N_19433,N_19285);
xor U19614 (N_19614,N_19340,N_19059);
nor U19615 (N_19615,N_19233,N_19302);
or U19616 (N_19616,N_19027,N_19424);
nor U19617 (N_19617,N_19097,N_19026);
and U19618 (N_19618,N_19144,N_19435);
nor U19619 (N_19619,N_19265,N_19210);
and U19620 (N_19620,N_19094,N_19153);
xor U19621 (N_19621,N_19164,N_19086);
and U19622 (N_19622,N_19381,N_19398);
xnor U19623 (N_19623,N_19212,N_19078);
nand U19624 (N_19624,N_19070,N_19455);
xor U19625 (N_19625,N_19392,N_19275);
or U19626 (N_19626,N_19230,N_19218);
xor U19627 (N_19627,N_19135,N_19262);
nand U19628 (N_19628,N_19496,N_19081);
nor U19629 (N_19629,N_19332,N_19349);
xor U19630 (N_19630,N_19422,N_19095);
xor U19631 (N_19631,N_19019,N_19405);
and U19632 (N_19632,N_19253,N_19403);
nor U19633 (N_19633,N_19000,N_19480);
xnor U19634 (N_19634,N_19439,N_19477);
and U19635 (N_19635,N_19298,N_19333);
nand U19636 (N_19636,N_19127,N_19465);
nand U19637 (N_19637,N_19449,N_19049);
nand U19638 (N_19638,N_19219,N_19223);
and U19639 (N_19639,N_19411,N_19234);
and U19640 (N_19640,N_19457,N_19181);
nand U19641 (N_19641,N_19221,N_19075);
xor U19642 (N_19642,N_19310,N_19129);
or U19643 (N_19643,N_19068,N_19090);
nor U19644 (N_19644,N_19022,N_19096);
or U19645 (N_19645,N_19246,N_19461);
nand U19646 (N_19646,N_19323,N_19011);
nor U19647 (N_19647,N_19400,N_19472);
nand U19648 (N_19648,N_19270,N_19329);
or U19649 (N_19649,N_19352,N_19066);
and U19650 (N_19650,N_19016,N_19238);
nor U19651 (N_19651,N_19171,N_19256);
nor U19652 (N_19652,N_19056,N_19172);
nor U19653 (N_19653,N_19240,N_19002);
and U19654 (N_19654,N_19319,N_19079);
and U19655 (N_19655,N_19087,N_19309);
nor U19656 (N_19656,N_19456,N_19366);
and U19657 (N_19657,N_19091,N_19410);
nor U19658 (N_19658,N_19418,N_19428);
nand U19659 (N_19659,N_19085,N_19125);
xor U19660 (N_19660,N_19438,N_19371);
xnor U19661 (N_19661,N_19014,N_19485);
or U19662 (N_19662,N_19341,N_19283);
xor U19663 (N_19663,N_19017,N_19053);
or U19664 (N_19664,N_19361,N_19155);
nand U19665 (N_19665,N_19495,N_19471);
or U19666 (N_19666,N_19128,N_19132);
and U19667 (N_19667,N_19088,N_19093);
and U19668 (N_19668,N_19156,N_19491);
and U19669 (N_19669,N_19157,N_19451);
nand U19670 (N_19670,N_19136,N_19436);
nor U19671 (N_19671,N_19478,N_19043);
nand U19672 (N_19672,N_19378,N_19476);
nor U19673 (N_19673,N_19304,N_19454);
and U19674 (N_19674,N_19102,N_19131);
or U19675 (N_19675,N_19356,N_19174);
and U19676 (N_19676,N_19490,N_19379);
nor U19677 (N_19677,N_19330,N_19100);
or U19678 (N_19678,N_19313,N_19374);
and U19679 (N_19679,N_19370,N_19110);
and U19680 (N_19680,N_19162,N_19328);
or U19681 (N_19681,N_19149,N_19431);
nor U19682 (N_19682,N_19453,N_19462);
nor U19683 (N_19683,N_19202,N_19188);
xor U19684 (N_19684,N_19152,N_19065);
and U19685 (N_19685,N_19376,N_19076);
xnor U19686 (N_19686,N_19042,N_19460);
xor U19687 (N_19687,N_19320,N_19306);
xnor U19688 (N_19688,N_19160,N_19334);
nor U19689 (N_19689,N_19098,N_19360);
or U19690 (N_19690,N_19466,N_19297);
nand U19691 (N_19691,N_19048,N_19180);
xnor U19692 (N_19692,N_19409,N_19446);
xor U19693 (N_19693,N_19140,N_19147);
and U19694 (N_19694,N_19497,N_19318);
and U19695 (N_19695,N_19200,N_19486);
nor U19696 (N_19696,N_19384,N_19347);
and U19697 (N_19697,N_19247,N_19452);
or U19698 (N_19698,N_19003,N_19358);
and U19699 (N_19699,N_19186,N_19175);
nand U19700 (N_19700,N_19443,N_19146);
and U19701 (N_19701,N_19463,N_19034);
nor U19702 (N_19702,N_19350,N_19077);
nand U19703 (N_19703,N_19369,N_19041);
or U19704 (N_19704,N_19440,N_19216);
nor U19705 (N_19705,N_19326,N_19161);
nand U19706 (N_19706,N_19386,N_19138);
xnor U19707 (N_19707,N_19260,N_19286);
xnor U19708 (N_19708,N_19268,N_19294);
nor U19709 (N_19709,N_19173,N_19064);
nor U19710 (N_19710,N_19324,N_19021);
xnor U19711 (N_19711,N_19242,N_19325);
or U19712 (N_19712,N_19282,N_19215);
xor U19713 (N_19713,N_19434,N_19067);
xnor U19714 (N_19714,N_19108,N_19395);
nor U19715 (N_19715,N_19442,N_19111);
nand U19716 (N_19716,N_19029,N_19469);
and U19717 (N_19717,N_19362,N_19423);
and U19718 (N_19718,N_19208,N_19321);
and U19719 (N_19719,N_19425,N_19237);
or U19720 (N_19720,N_19168,N_19249);
xnor U19721 (N_19721,N_19383,N_19206);
nand U19722 (N_19722,N_19291,N_19467);
or U19723 (N_19723,N_19317,N_19227);
and U19724 (N_19724,N_19336,N_19459);
and U19725 (N_19725,N_19007,N_19308);
or U19726 (N_19726,N_19355,N_19220);
xor U19727 (N_19727,N_19009,N_19427);
xor U19728 (N_19728,N_19314,N_19474);
nor U19729 (N_19729,N_19192,N_19184);
or U19730 (N_19730,N_19191,N_19001);
or U19731 (N_19731,N_19343,N_19289);
and U19732 (N_19732,N_19113,N_19150);
or U19733 (N_19733,N_19115,N_19385);
xor U19734 (N_19734,N_19413,N_19266);
xor U19735 (N_19735,N_19315,N_19189);
nor U19736 (N_19736,N_19198,N_19046);
or U19737 (N_19737,N_19225,N_19190);
nand U19738 (N_19738,N_19033,N_19372);
or U19739 (N_19739,N_19408,N_19414);
nor U19740 (N_19740,N_19031,N_19401);
and U19741 (N_19741,N_19229,N_19382);
nor U19742 (N_19742,N_19207,N_19357);
nand U19743 (N_19743,N_19339,N_19228);
or U19744 (N_19744,N_19470,N_19203);
xnor U19745 (N_19745,N_19130,N_19114);
nor U19746 (N_19746,N_19447,N_19448);
xor U19747 (N_19747,N_19055,N_19035);
and U19748 (N_19748,N_19226,N_19287);
or U19749 (N_19749,N_19213,N_19271);
nor U19750 (N_19750,N_19133,N_19207);
nand U19751 (N_19751,N_19117,N_19464);
nor U19752 (N_19752,N_19281,N_19296);
nor U19753 (N_19753,N_19479,N_19234);
and U19754 (N_19754,N_19053,N_19013);
and U19755 (N_19755,N_19428,N_19443);
xor U19756 (N_19756,N_19214,N_19035);
nand U19757 (N_19757,N_19144,N_19356);
nand U19758 (N_19758,N_19290,N_19417);
xor U19759 (N_19759,N_19060,N_19025);
or U19760 (N_19760,N_19255,N_19391);
or U19761 (N_19761,N_19168,N_19163);
and U19762 (N_19762,N_19442,N_19286);
nor U19763 (N_19763,N_19188,N_19441);
and U19764 (N_19764,N_19143,N_19425);
and U19765 (N_19765,N_19061,N_19427);
xor U19766 (N_19766,N_19292,N_19270);
nor U19767 (N_19767,N_19435,N_19182);
or U19768 (N_19768,N_19160,N_19150);
or U19769 (N_19769,N_19090,N_19003);
nand U19770 (N_19770,N_19141,N_19271);
nor U19771 (N_19771,N_19222,N_19113);
xor U19772 (N_19772,N_19358,N_19486);
xnor U19773 (N_19773,N_19154,N_19426);
nand U19774 (N_19774,N_19235,N_19438);
xor U19775 (N_19775,N_19270,N_19454);
xnor U19776 (N_19776,N_19018,N_19200);
nand U19777 (N_19777,N_19340,N_19165);
nand U19778 (N_19778,N_19097,N_19153);
or U19779 (N_19779,N_19024,N_19405);
and U19780 (N_19780,N_19496,N_19149);
and U19781 (N_19781,N_19119,N_19412);
nor U19782 (N_19782,N_19040,N_19173);
nor U19783 (N_19783,N_19203,N_19103);
and U19784 (N_19784,N_19428,N_19131);
nor U19785 (N_19785,N_19378,N_19093);
xnor U19786 (N_19786,N_19131,N_19229);
nor U19787 (N_19787,N_19286,N_19299);
xor U19788 (N_19788,N_19288,N_19491);
nor U19789 (N_19789,N_19232,N_19417);
and U19790 (N_19790,N_19202,N_19440);
nor U19791 (N_19791,N_19434,N_19150);
xnor U19792 (N_19792,N_19357,N_19020);
nor U19793 (N_19793,N_19071,N_19382);
xor U19794 (N_19794,N_19133,N_19433);
nand U19795 (N_19795,N_19419,N_19286);
and U19796 (N_19796,N_19353,N_19096);
xnor U19797 (N_19797,N_19471,N_19240);
or U19798 (N_19798,N_19405,N_19147);
nor U19799 (N_19799,N_19069,N_19223);
or U19800 (N_19800,N_19400,N_19245);
nand U19801 (N_19801,N_19357,N_19426);
nand U19802 (N_19802,N_19452,N_19004);
nand U19803 (N_19803,N_19494,N_19072);
nand U19804 (N_19804,N_19082,N_19286);
xor U19805 (N_19805,N_19060,N_19122);
and U19806 (N_19806,N_19373,N_19065);
or U19807 (N_19807,N_19436,N_19314);
nand U19808 (N_19808,N_19487,N_19444);
or U19809 (N_19809,N_19331,N_19003);
nor U19810 (N_19810,N_19091,N_19457);
nand U19811 (N_19811,N_19338,N_19456);
nand U19812 (N_19812,N_19212,N_19391);
or U19813 (N_19813,N_19275,N_19039);
xor U19814 (N_19814,N_19179,N_19015);
nor U19815 (N_19815,N_19044,N_19126);
nand U19816 (N_19816,N_19110,N_19234);
and U19817 (N_19817,N_19407,N_19202);
and U19818 (N_19818,N_19140,N_19380);
or U19819 (N_19819,N_19339,N_19409);
and U19820 (N_19820,N_19132,N_19332);
or U19821 (N_19821,N_19464,N_19062);
xor U19822 (N_19822,N_19015,N_19418);
nor U19823 (N_19823,N_19286,N_19028);
or U19824 (N_19824,N_19274,N_19313);
xor U19825 (N_19825,N_19479,N_19298);
and U19826 (N_19826,N_19499,N_19133);
or U19827 (N_19827,N_19334,N_19072);
or U19828 (N_19828,N_19356,N_19449);
or U19829 (N_19829,N_19403,N_19281);
or U19830 (N_19830,N_19181,N_19251);
or U19831 (N_19831,N_19321,N_19102);
xnor U19832 (N_19832,N_19068,N_19254);
nor U19833 (N_19833,N_19135,N_19202);
nand U19834 (N_19834,N_19271,N_19263);
xnor U19835 (N_19835,N_19357,N_19412);
and U19836 (N_19836,N_19473,N_19244);
nor U19837 (N_19837,N_19066,N_19316);
nand U19838 (N_19838,N_19225,N_19387);
xnor U19839 (N_19839,N_19433,N_19309);
or U19840 (N_19840,N_19163,N_19006);
xor U19841 (N_19841,N_19088,N_19112);
nor U19842 (N_19842,N_19305,N_19472);
nor U19843 (N_19843,N_19424,N_19113);
xor U19844 (N_19844,N_19216,N_19268);
xor U19845 (N_19845,N_19103,N_19235);
or U19846 (N_19846,N_19351,N_19256);
nand U19847 (N_19847,N_19325,N_19112);
nor U19848 (N_19848,N_19273,N_19075);
xor U19849 (N_19849,N_19174,N_19260);
and U19850 (N_19850,N_19126,N_19012);
nor U19851 (N_19851,N_19140,N_19385);
nor U19852 (N_19852,N_19059,N_19386);
or U19853 (N_19853,N_19458,N_19444);
nand U19854 (N_19854,N_19314,N_19211);
or U19855 (N_19855,N_19229,N_19077);
xor U19856 (N_19856,N_19080,N_19070);
or U19857 (N_19857,N_19365,N_19450);
or U19858 (N_19858,N_19349,N_19480);
nor U19859 (N_19859,N_19204,N_19105);
xor U19860 (N_19860,N_19021,N_19081);
nand U19861 (N_19861,N_19262,N_19173);
nor U19862 (N_19862,N_19059,N_19431);
nand U19863 (N_19863,N_19026,N_19131);
nor U19864 (N_19864,N_19374,N_19007);
nor U19865 (N_19865,N_19419,N_19233);
nor U19866 (N_19866,N_19085,N_19276);
nor U19867 (N_19867,N_19408,N_19044);
xnor U19868 (N_19868,N_19266,N_19164);
nand U19869 (N_19869,N_19214,N_19205);
or U19870 (N_19870,N_19109,N_19262);
or U19871 (N_19871,N_19357,N_19127);
xnor U19872 (N_19872,N_19439,N_19072);
nor U19873 (N_19873,N_19330,N_19392);
nor U19874 (N_19874,N_19240,N_19234);
and U19875 (N_19875,N_19375,N_19497);
nand U19876 (N_19876,N_19367,N_19414);
nor U19877 (N_19877,N_19221,N_19471);
xor U19878 (N_19878,N_19459,N_19198);
and U19879 (N_19879,N_19260,N_19191);
or U19880 (N_19880,N_19104,N_19273);
nand U19881 (N_19881,N_19038,N_19298);
or U19882 (N_19882,N_19448,N_19089);
or U19883 (N_19883,N_19432,N_19411);
nand U19884 (N_19884,N_19081,N_19288);
or U19885 (N_19885,N_19477,N_19191);
xor U19886 (N_19886,N_19260,N_19497);
or U19887 (N_19887,N_19313,N_19217);
nand U19888 (N_19888,N_19055,N_19008);
and U19889 (N_19889,N_19496,N_19085);
nor U19890 (N_19890,N_19223,N_19312);
nor U19891 (N_19891,N_19179,N_19067);
or U19892 (N_19892,N_19119,N_19243);
nand U19893 (N_19893,N_19179,N_19375);
or U19894 (N_19894,N_19115,N_19009);
nand U19895 (N_19895,N_19265,N_19236);
xor U19896 (N_19896,N_19470,N_19159);
xor U19897 (N_19897,N_19037,N_19466);
and U19898 (N_19898,N_19363,N_19218);
and U19899 (N_19899,N_19011,N_19375);
xnor U19900 (N_19900,N_19068,N_19491);
nor U19901 (N_19901,N_19258,N_19315);
xor U19902 (N_19902,N_19440,N_19014);
or U19903 (N_19903,N_19196,N_19143);
or U19904 (N_19904,N_19339,N_19395);
nand U19905 (N_19905,N_19210,N_19096);
nand U19906 (N_19906,N_19264,N_19116);
nor U19907 (N_19907,N_19134,N_19167);
nand U19908 (N_19908,N_19164,N_19220);
nand U19909 (N_19909,N_19137,N_19473);
and U19910 (N_19910,N_19245,N_19243);
nand U19911 (N_19911,N_19297,N_19008);
xor U19912 (N_19912,N_19222,N_19051);
xnor U19913 (N_19913,N_19331,N_19208);
xor U19914 (N_19914,N_19461,N_19088);
xor U19915 (N_19915,N_19366,N_19058);
xor U19916 (N_19916,N_19062,N_19272);
and U19917 (N_19917,N_19469,N_19454);
nor U19918 (N_19918,N_19222,N_19392);
nor U19919 (N_19919,N_19359,N_19002);
nor U19920 (N_19920,N_19323,N_19369);
nor U19921 (N_19921,N_19104,N_19234);
nand U19922 (N_19922,N_19203,N_19163);
or U19923 (N_19923,N_19325,N_19149);
nor U19924 (N_19924,N_19358,N_19078);
nor U19925 (N_19925,N_19002,N_19155);
and U19926 (N_19926,N_19115,N_19204);
nor U19927 (N_19927,N_19014,N_19448);
nand U19928 (N_19928,N_19222,N_19104);
nand U19929 (N_19929,N_19488,N_19036);
xnor U19930 (N_19930,N_19402,N_19000);
nand U19931 (N_19931,N_19389,N_19050);
nor U19932 (N_19932,N_19102,N_19106);
xor U19933 (N_19933,N_19428,N_19464);
nand U19934 (N_19934,N_19476,N_19087);
nand U19935 (N_19935,N_19035,N_19229);
nor U19936 (N_19936,N_19148,N_19459);
nand U19937 (N_19937,N_19311,N_19264);
nor U19938 (N_19938,N_19343,N_19287);
and U19939 (N_19939,N_19307,N_19464);
xnor U19940 (N_19940,N_19164,N_19423);
nor U19941 (N_19941,N_19122,N_19493);
xnor U19942 (N_19942,N_19137,N_19200);
and U19943 (N_19943,N_19320,N_19199);
or U19944 (N_19944,N_19490,N_19212);
nand U19945 (N_19945,N_19277,N_19075);
and U19946 (N_19946,N_19060,N_19435);
and U19947 (N_19947,N_19288,N_19110);
and U19948 (N_19948,N_19172,N_19265);
or U19949 (N_19949,N_19429,N_19137);
nand U19950 (N_19950,N_19241,N_19426);
and U19951 (N_19951,N_19221,N_19377);
xnor U19952 (N_19952,N_19161,N_19331);
nor U19953 (N_19953,N_19491,N_19350);
xor U19954 (N_19954,N_19033,N_19011);
or U19955 (N_19955,N_19219,N_19246);
nand U19956 (N_19956,N_19439,N_19013);
and U19957 (N_19957,N_19036,N_19136);
and U19958 (N_19958,N_19062,N_19081);
or U19959 (N_19959,N_19479,N_19193);
xnor U19960 (N_19960,N_19059,N_19442);
or U19961 (N_19961,N_19492,N_19483);
and U19962 (N_19962,N_19479,N_19492);
nor U19963 (N_19963,N_19365,N_19488);
nor U19964 (N_19964,N_19454,N_19307);
and U19965 (N_19965,N_19204,N_19416);
or U19966 (N_19966,N_19263,N_19039);
or U19967 (N_19967,N_19431,N_19411);
nor U19968 (N_19968,N_19344,N_19308);
nand U19969 (N_19969,N_19143,N_19122);
xor U19970 (N_19970,N_19120,N_19083);
nor U19971 (N_19971,N_19049,N_19179);
or U19972 (N_19972,N_19062,N_19216);
and U19973 (N_19973,N_19017,N_19403);
nor U19974 (N_19974,N_19177,N_19395);
nand U19975 (N_19975,N_19369,N_19318);
nand U19976 (N_19976,N_19363,N_19334);
xnor U19977 (N_19977,N_19478,N_19092);
and U19978 (N_19978,N_19414,N_19264);
or U19979 (N_19979,N_19183,N_19318);
and U19980 (N_19980,N_19004,N_19275);
xor U19981 (N_19981,N_19056,N_19418);
and U19982 (N_19982,N_19136,N_19087);
xor U19983 (N_19983,N_19054,N_19035);
and U19984 (N_19984,N_19354,N_19232);
nand U19985 (N_19985,N_19342,N_19059);
nor U19986 (N_19986,N_19059,N_19029);
nand U19987 (N_19987,N_19106,N_19020);
and U19988 (N_19988,N_19059,N_19306);
xor U19989 (N_19989,N_19161,N_19481);
nor U19990 (N_19990,N_19051,N_19041);
or U19991 (N_19991,N_19334,N_19045);
xnor U19992 (N_19992,N_19029,N_19462);
xnor U19993 (N_19993,N_19156,N_19030);
or U19994 (N_19994,N_19361,N_19446);
nor U19995 (N_19995,N_19181,N_19046);
and U19996 (N_19996,N_19471,N_19287);
nor U19997 (N_19997,N_19463,N_19096);
nor U19998 (N_19998,N_19436,N_19218);
nor U19999 (N_19999,N_19071,N_19234);
nor U20000 (N_20000,N_19828,N_19925);
or U20001 (N_20001,N_19788,N_19558);
or U20002 (N_20002,N_19520,N_19934);
or U20003 (N_20003,N_19849,N_19709);
and U20004 (N_20004,N_19635,N_19726);
or U20005 (N_20005,N_19852,N_19620);
and U20006 (N_20006,N_19910,N_19835);
nor U20007 (N_20007,N_19814,N_19880);
xor U20008 (N_20008,N_19525,N_19713);
nor U20009 (N_20009,N_19649,N_19899);
and U20010 (N_20010,N_19924,N_19837);
nor U20011 (N_20011,N_19956,N_19686);
xnor U20012 (N_20012,N_19907,N_19903);
nand U20013 (N_20013,N_19871,N_19563);
nor U20014 (N_20014,N_19808,N_19574);
nor U20015 (N_20015,N_19592,N_19509);
nand U20016 (N_20016,N_19840,N_19610);
or U20017 (N_20017,N_19973,N_19549);
and U20018 (N_20018,N_19969,N_19733);
and U20019 (N_20019,N_19851,N_19653);
nand U20020 (N_20020,N_19571,N_19751);
or U20021 (N_20021,N_19701,N_19506);
and U20022 (N_20022,N_19916,N_19881);
and U20023 (N_20023,N_19514,N_19942);
nor U20024 (N_20024,N_19995,N_19984);
or U20025 (N_20025,N_19669,N_19583);
xor U20026 (N_20026,N_19988,N_19636);
nand U20027 (N_20027,N_19890,N_19914);
xor U20028 (N_20028,N_19845,N_19820);
nor U20029 (N_20029,N_19867,N_19927);
nand U20030 (N_20030,N_19508,N_19959);
nor U20031 (N_20031,N_19770,N_19875);
nand U20032 (N_20032,N_19750,N_19690);
or U20033 (N_20033,N_19576,N_19797);
nor U20034 (N_20034,N_19812,N_19947);
xnor U20035 (N_20035,N_19609,N_19803);
and U20036 (N_20036,N_19911,N_19912);
and U20037 (N_20037,N_19585,N_19985);
nor U20038 (N_20038,N_19843,N_19938);
xnor U20039 (N_20039,N_19930,N_19975);
and U20040 (N_20040,N_19554,N_19968);
xor U20041 (N_20041,N_19760,N_19996);
nor U20042 (N_20042,N_19602,N_19965);
xor U20043 (N_20043,N_19889,N_19815);
or U20044 (N_20044,N_19736,N_19562);
or U20045 (N_20045,N_19891,N_19601);
nor U20046 (N_20046,N_19801,N_19778);
or U20047 (N_20047,N_19958,N_19948);
nand U20048 (N_20048,N_19595,N_19672);
xnor U20049 (N_20049,N_19680,N_19901);
and U20050 (N_20050,N_19710,N_19747);
nor U20051 (N_20051,N_19668,N_19557);
xor U20052 (N_20052,N_19687,N_19898);
or U20053 (N_20053,N_19749,N_19839);
or U20054 (N_20054,N_19630,N_19842);
and U20055 (N_20055,N_19704,N_19847);
xnor U20056 (N_20056,N_19765,N_19708);
and U20057 (N_20057,N_19722,N_19882);
nor U20058 (N_20058,N_19699,N_19949);
and U20059 (N_20059,N_19874,N_19718);
xor U20060 (N_20060,N_19634,N_19950);
nand U20061 (N_20061,N_19999,N_19553);
and U20062 (N_20062,N_19759,N_19757);
xor U20063 (N_20063,N_19724,N_19646);
and U20064 (N_20064,N_19945,N_19922);
xnor U20065 (N_20065,N_19537,N_19795);
nor U20066 (N_20066,N_19737,N_19863);
or U20067 (N_20067,N_19829,N_19512);
nand U20068 (N_20068,N_19594,N_19769);
and U20069 (N_20069,N_19569,N_19859);
nand U20070 (N_20070,N_19885,N_19982);
nand U20071 (N_20071,N_19918,N_19732);
and U20072 (N_20072,N_19648,N_19540);
and U20073 (N_20073,N_19887,N_19626);
xor U20074 (N_20074,N_19864,N_19692);
xnor U20075 (N_20075,N_19857,N_19575);
or U20076 (N_20076,N_19846,N_19748);
nor U20077 (N_20077,N_19834,N_19696);
and U20078 (N_20078,N_19972,N_19979);
nand U20079 (N_20079,N_19772,N_19745);
and U20080 (N_20080,N_19678,N_19742);
nor U20081 (N_20081,N_19931,N_19593);
or U20082 (N_20082,N_19976,N_19675);
and U20083 (N_20083,N_19654,N_19667);
xor U20084 (N_20084,N_19856,N_19831);
or U20085 (N_20085,N_19767,N_19937);
nand U20086 (N_20086,N_19728,N_19622);
or U20087 (N_20087,N_19762,N_19673);
xnor U20088 (N_20088,N_19717,N_19621);
nor U20089 (N_20089,N_19816,N_19682);
xor U20090 (N_20090,N_19544,N_19596);
xnor U20091 (N_20091,N_19700,N_19502);
nor U20092 (N_20092,N_19735,N_19894);
xnor U20093 (N_20093,N_19702,N_19993);
or U20094 (N_20094,N_19613,N_19866);
nor U20095 (N_20095,N_19739,N_19651);
nor U20096 (N_20096,N_19813,N_19522);
nand U20097 (N_20097,N_19543,N_19555);
xor U20098 (N_20098,N_19510,N_19637);
nor U20099 (N_20099,N_19752,N_19986);
and U20100 (N_20100,N_19598,N_19560);
or U20101 (N_20101,N_19695,N_19793);
and U20102 (N_20102,N_19868,N_19940);
and U20103 (N_20103,N_19679,N_19774);
nor U20104 (N_20104,N_19643,N_19865);
or U20105 (N_20105,N_19943,N_19923);
nor U20106 (N_20106,N_19779,N_19853);
xor U20107 (N_20107,N_19967,N_19548);
nand U20108 (N_20108,N_19565,N_19906);
or U20109 (N_20109,N_19507,N_19960);
or U20110 (N_20110,N_19823,N_19581);
nand U20111 (N_20111,N_19974,N_19902);
xor U20112 (N_20112,N_19661,N_19504);
nand U20113 (N_20113,N_19784,N_19604);
and U20114 (N_20114,N_19542,N_19663);
nand U20115 (N_20115,N_19693,N_19719);
nor U20116 (N_20116,N_19633,N_19670);
nor U20117 (N_20117,N_19536,N_19981);
and U20118 (N_20118,N_19624,N_19939);
nand U20119 (N_20119,N_19792,N_19721);
or U20120 (N_20120,N_19546,N_19773);
nand U20121 (N_20121,N_19926,N_19952);
xor U20122 (N_20122,N_19676,N_19954);
xor U20123 (N_20123,N_19659,N_19564);
nor U20124 (N_20124,N_19935,N_19917);
nor U20125 (N_20125,N_19505,N_19753);
nor U20126 (N_20126,N_19664,N_19720);
or U20127 (N_20127,N_19612,N_19511);
nand U20128 (N_20128,N_19928,N_19987);
xor U20129 (N_20129,N_19531,N_19919);
xnor U20130 (N_20130,N_19878,N_19545);
nand U20131 (N_20131,N_19639,N_19578);
nor U20132 (N_20132,N_19821,N_19627);
nor U20133 (N_20133,N_19798,N_19755);
or U20134 (N_20134,N_19730,N_19645);
nor U20135 (N_20135,N_19833,N_19660);
nand U20136 (N_20136,N_19589,N_19962);
xor U20137 (N_20137,N_19777,N_19892);
and U20138 (N_20138,N_19811,N_19799);
xor U20139 (N_20139,N_19688,N_19744);
and U20140 (N_20140,N_19825,N_19883);
and U20141 (N_20141,N_19703,N_19625);
and U20142 (N_20142,N_19523,N_19838);
or U20143 (N_20143,N_19666,N_19603);
or U20144 (N_20144,N_19805,N_19638);
xnor U20145 (N_20145,N_19991,N_19599);
nor U20146 (N_20146,N_19587,N_19832);
nor U20147 (N_20147,N_19944,N_19617);
xor U20148 (N_20148,N_19964,N_19781);
nand U20149 (N_20149,N_19607,N_19684);
nor U20150 (N_20150,N_19641,N_19980);
nor U20151 (N_20151,N_19656,N_19989);
nand U20152 (N_20152,N_19776,N_19904);
nor U20153 (N_20153,N_19715,N_19992);
and U20154 (N_20154,N_19802,N_19909);
or U20155 (N_20155,N_19674,N_19539);
xor U20156 (N_20156,N_19528,N_19614);
or U20157 (N_20157,N_19888,N_19824);
and U20158 (N_20158,N_19970,N_19963);
or U20159 (N_20159,N_19997,N_19933);
xor U20160 (N_20160,N_19579,N_19941);
nor U20161 (N_20161,N_19896,N_19810);
nand U20162 (N_20162,N_19794,N_19771);
nor U20163 (N_20163,N_19761,N_19615);
and U20164 (N_20164,N_19550,N_19628);
or U20165 (N_20165,N_19527,N_19605);
or U20166 (N_20166,N_19725,N_19644);
nor U20167 (N_20167,N_19913,N_19915);
and U20168 (N_20168,N_19862,N_19681);
nor U20169 (N_20169,N_19920,N_19559);
and U20170 (N_20170,N_19652,N_19848);
or U20171 (N_20171,N_19691,N_19590);
and U20172 (N_20172,N_19642,N_19501);
nor U20173 (N_20173,N_19905,N_19657);
or U20174 (N_20174,N_19712,N_19796);
xor U20175 (N_20175,N_19500,N_19729);
and U20176 (N_20176,N_19978,N_19809);
and U20177 (N_20177,N_19876,N_19530);
nor U20178 (N_20178,N_19606,N_19618);
nor U20179 (N_20179,N_19854,N_19764);
nor U20180 (N_20180,N_19597,N_19631);
xnor U20181 (N_20181,N_19754,N_19870);
xnor U20182 (N_20182,N_19588,N_19685);
nand U20183 (N_20183,N_19850,N_19577);
nor U20184 (N_20184,N_19671,N_19541);
and U20185 (N_20185,N_19766,N_19932);
xor U20186 (N_20186,N_19727,N_19705);
nand U20187 (N_20187,N_19689,N_19716);
or U20188 (N_20188,N_19584,N_19547);
or U20189 (N_20189,N_19619,N_19858);
nor U20190 (N_20190,N_19783,N_19785);
or U20191 (N_20191,N_19807,N_19731);
nand U20192 (N_20192,N_19780,N_19658);
nand U20193 (N_20193,N_19647,N_19826);
and U20194 (N_20194,N_19786,N_19782);
or U20195 (N_20195,N_19591,N_19743);
and U20196 (N_20196,N_19741,N_19921);
or U20197 (N_20197,N_19532,N_19860);
nor U20198 (N_20198,N_19697,N_19830);
xor U20199 (N_20199,N_19971,N_19568);
or U20200 (N_20200,N_19534,N_19819);
or U20201 (N_20201,N_19841,N_19998);
xnor U20202 (N_20202,N_19650,N_19869);
and U20203 (N_20203,N_19977,N_19763);
nand U20204 (N_20204,N_19711,N_19655);
nand U20205 (N_20205,N_19877,N_19608);
nand U20206 (N_20206,N_19526,N_19518);
and U20207 (N_20207,N_19775,N_19519);
and U20208 (N_20208,N_19677,N_19817);
and U20209 (N_20209,N_19662,N_19758);
or U20210 (N_20210,N_19698,N_19804);
xor U20211 (N_20211,N_19535,N_19929);
or U20212 (N_20212,N_19768,N_19879);
and U20213 (N_20213,N_19836,N_19517);
xnor U20214 (N_20214,N_19953,N_19503);
and U20215 (N_20215,N_19600,N_19827);
nand U20216 (N_20216,N_19893,N_19990);
xnor U20217 (N_20217,N_19861,N_19582);
xnor U20218 (N_20218,N_19818,N_19665);
nor U20219 (N_20219,N_19886,N_19936);
or U20220 (N_20220,N_19966,N_19533);
and U20221 (N_20221,N_19900,N_19586);
or U20222 (N_20222,N_19640,N_19897);
nor U20223 (N_20223,N_19567,N_19552);
nor U20224 (N_20224,N_19683,N_19895);
nand U20225 (N_20225,N_19551,N_19872);
and U20226 (N_20226,N_19951,N_19791);
nand U20227 (N_20227,N_19994,N_19707);
and U20228 (N_20228,N_19787,N_19515);
nor U20229 (N_20229,N_19844,N_19623);
or U20230 (N_20230,N_19572,N_19873);
xor U20231 (N_20231,N_19516,N_19955);
or U20232 (N_20232,N_19740,N_19790);
and U20233 (N_20233,N_19694,N_19908);
nand U20234 (N_20234,N_19822,N_19957);
and U20235 (N_20235,N_19756,N_19961);
nor U20236 (N_20236,N_19538,N_19946);
and U20237 (N_20237,N_19570,N_19734);
and U20238 (N_20238,N_19561,N_19806);
nand U20239 (N_20239,N_19746,N_19580);
and U20240 (N_20240,N_19521,N_19629);
and U20241 (N_20241,N_19855,N_19983);
xor U20242 (N_20242,N_19789,N_19524);
nor U20243 (N_20243,N_19738,N_19723);
or U20244 (N_20244,N_19513,N_19616);
nand U20245 (N_20245,N_19573,N_19556);
nor U20246 (N_20246,N_19714,N_19529);
or U20247 (N_20247,N_19611,N_19800);
nor U20248 (N_20248,N_19632,N_19706);
nor U20249 (N_20249,N_19566,N_19884);
xor U20250 (N_20250,N_19649,N_19607);
xnor U20251 (N_20251,N_19551,N_19716);
and U20252 (N_20252,N_19546,N_19830);
xnor U20253 (N_20253,N_19665,N_19538);
nor U20254 (N_20254,N_19626,N_19786);
or U20255 (N_20255,N_19577,N_19954);
xor U20256 (N_20256,N_19518,N_19843);
and U20257 (N_20257,N_19993,N_19937);
xnor U20258 (N_20258,N_19772,N_19545);
or U20259 (N_20259,N_19609,N_19577);
xor U20260 (N_20260,N_19710,N_19735);
nand U20261 (N_20261,N_19953,N_19516);
and U20262 (N_20262,N_19801,N_19873);
nor U20263 (N_20263,N_19957,N_19557);
nand U20264 (N_20264,N_19525,N_19587);
and U20265 (N_20265,N_19660,N_19630);
and U20266 (N_20266,N_19682,N_19688);
and U20267 (N_20267,N_19503,N_19785);
nand U20268 (N_20268,N_19617,N_19968);
nor U20269 (N_20269,N_19725,N_19928);
xnor U20270 (N_20270,N_19696,N_19871);
nor U20271 (N_20271,N_19932,N_19892);
nor U20272 (N_20272,N_19744,N_19888);
and U20273 (N_20273,N_19831,N_19676);
nor U20274 (N_20274,N_19729,N_19984);
nor U20275 (N_20275,N_19674,N_19533);
xor U20276 (N_20276,N_19979,N_19906);
nor U20277 (N_20277,N_19758,N_19707);
nand U20278 (N_20278,N_19525,N_19911);
or U20279 (N_20279,N_19927,N_19820);
nand U20280 (N_20280,N_19513,N_19968);
nand U20281 (N_20281,N_19535,N_19670);
nor U20282 (N_20282,N_19724,N_19968);
xnor U20283 (N_20283,N_19818,N_19867);
xor U20284 (N_20284,N_19930,N_19855);
nor U20285 (N_20285,N_19681,N_19769);
or U20286 (N_20286,N_19906,N_19552);
or U20287 (N_20287,N_19776,N_19819);
or U20288 (N_20288,N_19875,N_19656);
nand U20289 (N_20289,N_19617,N_19611);
or U20290 (N_20290,N_19981,N_19779);
and U20291 (N_20291,N_19508,N_19528);
xnor U20292 (N_20292,N_19949,N_19702);
nor U20293 (N_20293,N_19648,N_19877);
nor U20294 (N_20294,N_19724,N_19894);
and U20295 (N_20295,N_19877,N_19942);
nor U20296 (N_20296,N_19810,N_19989);
nor U20297 (N_20297,N_19658,N_19533);
or U20298 (N_20298,N_19612,N_19943);
and U20299 (N_20299,N_19973,N_19969);
nand U20300 (N_20300,N_19960,N_19608);
or U20301 (N_20301,N_19885,N_19791);
nand U20302 (N_20302,N_19769,N_19654);
nand U20303 (N_20303,N_19640,N_19705);
xnor U20304 (N_20304,N_19680,N_19830);
and U20305 (N_20305,N_19880,N_19746);
or U20306 (N_20306,N_19542,N_19959);
nor U20307 (N_20307,N_19972,N_19532);
and U20308 (N_20308,N_19935,N_19908);
and U20309 (N_20309,N_19906,N_19690);
xor U20310 (N_20310,N_19584,N_19538);
or U20311 (N_20311,N_19545,N_19903);
xnor U20312 (N_20312,N_19933,N_19705);
and U20313 (N_20313,N_19830,N_19688);
and U20314 (N_20314,N_19905,N_19835);
nor U20315 (N_20315,N_19966,N_19739);
and U20316 (N_20316,N_19921,N_19640);
and U20317 (N_20317,N_19950,N_19819);
nand U20318 (N_20318,N_19904,N_19768);
nand U20319 (N_20319,N_19720,N_19919);
nor U20320 (N_20320,N_19840,N_19544);
or U20321 (N_20321,N_19906,N_19776);
xnor U20322 (N_20322,N_19817,N_19761);
nand U20323 (N_20323,N_19534,N_19905);
nand U20324 (N_20324,N_19917,N_19969);
xor U20325 (N_20325,N_19982,N_19518);
xor U20326 (N_20326,N_19568,N_19727);
and U20327 (N_20327,N_19716,N_19968);
xor U20328 (N_20328,N_19502,N_19812);
xnor U20329 (N_20329,N_19686,N_19570);
and U20330 (N_20330,N_19796,N_19784);
or U20331 (N_20331,N_19926,N_19747);
or U20332 (N_20332,N_19734,N_19667);
or U20333 (N_20333,N_19660,N_19998);
nand U20334 (N_20334,N_19999,N_19566);
nor U20335 (N_20335,N_19987,N_19539);
and U20336 (N_20336,N_19615,N_19543);
or U20337 (N_20337,N_19620,N_19930);
and U20338 (N_20338,N_19743,N_19707);
nand U20339 (N_20339,N_19778,N_19851);
nor U20340 (N_20340,N_19531,N_19633);
xor U20341 (N_20341,N_19558,N_19640);
or U20342 (N_20342,N_19551,N_19909);
nand U20343 (N_20343,N_19627,N_19907);
nor U20344 (N_20344,N_19944,N_19739);
nor U20345 (N_20345,N_19957,N_19708);
nor U20346 (N_20346,N_19818,N_19574);
nand U20347 (N_20347,N_19730,N_19831);
nand U20348 (N_20348,N_19737,N_19749);
nand U20349 (N_20349,N_19765,N_19693);
nand U20350 (N_20350,N_19556,N_19848);
or U20351 (N_20351,N_19505,N_19604);
xor U20352 (N_20352,N_19751,N_19661);
nor U20353 (N_20353,N_19526,N_19725);
or U20354 (N_20354,N_19535,N_19896);
xor U20355 (N_20355,N_19909,N_19948);
xor U20356 (N_20356,N_19583,N_19529);
nor U20357 (N_20357,N_19808,N_19999);
or U20358 (N_20358,N_19637,N_19746);
nor U20359 (N_20359,N_19727,N_19776);
and U20360 (N_20360,N_19970,N_19825);
nand U20361 (N_20361,N_19958,N_19590);
or U20362 (N_20362,N_19724,N_19977);
nor U20363 (N_20363,N_19872,N_19552);
xor U20364 (N_20364,N_19781,N_19604);
nor U20365 (N_20365,N_19583,N_19846);
or U20366 (N_20366,N_19585,N_19877);
nor U20367 (N_20367,N_19966,N_19718);
or U20368 (N_20368,N_19805,N_19572);
nor U20369 (N_20369,N_19682,N_19742);
nand U20370 (N_20370,N_19521,N_19796);
xor U20371 (N_20371,N_19850,N_19907);
nand U20372 (N_20372,N_19637,N_19568);
nand U20373 (N_20373,N_19545,N_19715);
and U20374 (N_20374,N_19677,N_19548);
and U20375 (N_20375,N_19888,N_19874);
nor U20376 (N_20376,N_19661,N_19862);
and U20377 (N_20377,N_19965,N_19871);
and U20378 (N_20378,N_19803,N_19928);
nand U20379 (N_20379,N_19679,N_19806);
xnor U20380 (N_20380,N_19978,N_19503);
xnor U20381 (N_20381,N_19693,N_19570);
and U20382 (N_20382,N_19801,N_19646);
and U20383 (N_20383,N_19729,N_19957);
nand U20384 (N_20384,N_19541,N_19591);
or U20385 (N_20385,N_19925,N_19593);
or U20386 (N_20386,N_19628,N_19884);
nand U20387 (N_20387,N_19848,N_19575);
and U20388 (N_20388,N_19820,N_19538);
nand U20389 (N_20389,N_19946,N_19884);
or U20390 (N_20390,N_19632,N_19790);
and U20391 (N_20391,N_19909,N_19973);
nand U20392 (N_20392,N_19788,N_19776);
or U20393 (N_20393,N_19575,N_19883);
and U20394 (N_20394,N_19666,N_19842);
nor U20395 (N_20395,N_19981,N_19892);
nor U20396 (N_20396,N_19751,N_19875);
nand U20397 (N_20397,N_19818,N_19507);
xnor U20398 (N_20398,N_19794,N_19933);
nand U20399 (N_20399,N_19512,N_19851);
and U20400 (N_20400,N_19718,N_19724);
xnor U20401 (N_20401,N_19769,N_19575);
nand U20402 (N_20402,N_19501,N_19590);
nor U20403 (N_20403,N_19929,N_19952);
xor U20404 (N_20404,N_19839,N_19698);
xor U20405 (N_20405,N_19837,N_19532);
and U20406 (N_20406,N_19646,N_19859);
or U20407 (N_20407,N_19508,N_19570);
nand U20408 (N_20408,N_19848,N_19800);
nor U20409 (N_20409,N_19983,N_19922);
nand U20410 (N_20410,N_19627,N_19617);
xnor U20411 (N_20411,N_19813,N_19739);
nand U20412 (N_20412,N_19536,N_19998);
or U20413 (N_20413,N_19768,N_19837);
and U20414 (N_20414,N_19855,N_19638);
and U20415 (N_20415,N_19808,N_19939);
xnor U20416 (N_20416,N_19811,N_19821);
nand U20417 (N_20417,N_19701,N_19688);
xor U20418 (N_20418,N_19619,N_19580);
nor U20419 (N_20419,N_19970,N_19956);
xor U20420 (N_20420,N_19829,N_19997);
nor U20421 (N_20421,N_19716,N_19999);
nor U20422 (N_20422,N_19885,N_19890);
and U20423 (N_20423,N_19714,N_19838);
or U20424 (N_20424,N_19621,N_19789);
or U20425 (N_20425,N_19519,N_19947);
and U20426 (N_20426,N_19595,N_19910);
or U20427 (N_20427,N_19836,N_19973);
xnor U20428 (N_20428,N_19992,N_19668);
nand U20429 (N_20429,N_19695,N_19642);
nor U20430 (N_20430,N_19595,N_19887);
xnor U20431 (N_20431,N_19515,N_19643);
nand U20432 (N_20432,N_19867,N_19722);
and U20433 (N_20433,N_19625,N_19645);
and U20434 (N_20434,N_19505,N_19671);
or U20435 (N_20435,N_19708,N_19702);
and U20436 (N_20436,N_19923,N_19659);
and U20437 (N_20437,N_19795,N_19598);
or U20438 (N_20438,N_19727,N_19915);
or U20439 (N_20439,N_19890,N_19728);
or U20440 (N_20440,N_19686,N_19940);
nand U20441 (N_20441,N_19994,N_19521);
nand U20442 (N_20442,N_19656,N_19525);
or U20443 (N_20443,N_19718,N_19693);
and U20444 (N_20444,N_19905,N_19776);
or U20445 (N_20445,N_19814,N_19568);
and U20446 (N_20446,N_19972,N_19599);
nor U20447 (N_20447,N_19903,N_19984);
nand U20448 (N_20448,N_19655,N_19855);
xor U20449 (N_20449,N_19917,N_19587);
nor U20450 (N_20450,N_19942,N_19532);
nand U20451 (N_20451,N_19594,N_19702);
and U20452 (N_20452,N_19514,N_19606);
nor U20453 (N_20453,N_19733,N_19713);
nor U20454 (N_20454,N_19745,N_19716);
xor U20455 (N_20455,N_19539,N_19581);
nor U20456 (N_20456,N_19713,N_19896);
and U20457 (N_20457,N_19944,N_19724);
nor U20458 (N_20458,N_19839,N_19853);
xnor U20459 (N_20459,N_19636,N_19939);
nor U20460 (N_20460,N_19953,N_19832);
nor U20461 (N_20461,N_19596,N_19672);
and U20462 (N_20462,N_19500,N_19512);
xor U20463 (N_20463,N_19926,N_19642);
nor U20464 (N_20464,N_19543,N_19648);
xor U20465 (N_20465,N_19777,N_19689);
nand U20466 (N_20466,N_19769,N_19729);
xor U20467 (N_20467,N_19627,N_19502);
nor U20468 (N_20468,N_19958,N_19537);
nand U20469 (N_20469,N_19718,N_19648);
nand U20470 (N_20470,N_19808,N_19799);
nand U20471 (N_20471,N_19790,N_19810);
or U20472 (N_20472,N_19836,N_19861);
nand U20473 (N_20473,N_19709,N_19636);
or U20474 (N_20474,N_19788,N_19616);
xnor U20475 (N_20475,N_19500,N_19896);
xor U20476 (N_20476,N_19731,N_19662);
or U20477 (N_20477,N_19858,N_19880);
nand U20478 (N_20478,N_19758,N_19988);
nor U20479 (N_20479,N_19750,N_19609);
xor U20480 (N_20480,N_19725,N_19950);
nor U20481 (N_20481,N_19976,N_19583);
or U20482 (N_20482,N_19994,N_19701);
nor U20483 (N_20483,N_19628,N_19773);
xnor U20484 (N_20484,N_19797,N_19964);
or U20485 (N_20485,N_19894,N_19605);
and U20486 (N_20486,N_19636,N_19711);
nor U20487 (N_20487,N_19932,N_19685);
xor U20488 (N_20488,N_19812,N_19715);
and U20489 (N_20489,N_19822,N_19571);
and U20490 (N_20490,N_19649,N_19523);
xnor U20491 (N_20491,N_19519,N_19761);
xor U20492 (N_20492,N_19565,N_19755);
nor U20493 (N_20493,N_19810,N_19768);
nor U20494 (N_20494,N_19796,N_19589);
and U20495 (N_20495,N_19595,N_19881);
or U20496 (N_20496,N_19971,N_19584);
or U20497 (N_20497,N_19508,N_19817);
nor U20498 (N_20498,N_19961,N_19998);
nand U20499 (N_20499,N_19653,N_19658);
nand U20500 (N_20500,N_20010,N_20339);
xor U20501 (N_20501,N_20314,N_20490);
nor U20502 (N_20502,N_20057,N_20203);
nand U20503 (N_20503,N_20414,N_20014);
xnor U20504 (N_20504,N_20267,N_20037);
nand U20505 (N_20505,N_20047,N_20016);
and U20506 (N_20506,N_20297,N_20146);
or U20507 (N_20507,N_20184,N_20123);
nor U20508 (N_20508,N_20201,N_20159);
xnor U20509 (N_20509,N_20138,N_20394);
nand U20510 (N_20510,N_20245,N_20217);
xor U20511 (N_20511,N_20038,N_20074);
nor U20512 (N_20512,N_20359,N_20418);
or U20513 (N_20513,N_20457,N_20369);
or U20514 (N_20514,N_20006,N_20335);
xor U20515 (N_20515,N_20287,N_20374);
nor U20516 (N_20516,N_20273,N_20404);
nor U20517 (N_20517,N_20298,N_20009);
or U20518 (N_20518,N_20222,N_20248);
xor U20519 (N_20519,N_20432,N_20232);
nand U20520 (N_20520,N_20086,N_20459);
xnor U20521 (N_20521,N_20475,N_20401);
or U20522 (N_20522,N_20283,N_20258);
xor U20523 (N_20523,N_20356,N_20393);
or U20524 (N_20524,N_20063,N_20148);
nand U20525 (N_20525,N_20228,N_20041);
xor U20526 (N_20526,N_20291,N_20377);
nand U20527 (N_20527,N_20301,N_20387);
or U20528 (N_20528,N_20033,N_20462);
or U20529 (N_20529,N_20397,N_20115);
nand U20530 (N_20530,N_20199,N_20149);
xor U20531 (N_20531,N_20425,N_20350);
or U20532 (N_20532,N_20464,N_20077);
or U20533 (N_20533,N_20482,N_20155);
xor U20534 (N_20534,N_20214,N_20048);
xor U20535 (N_20535,N_20271,N_20489);
nor U20536 (N_20536,N_20160,N_20323);
or U20537 (N_20537,N_20054,N_20238);
or U20538 (N_20538,N_20315,N_20352);
and U20539 (N_20539,N_20223,N_20304);
or U20540 (N_20540,N_20257,N_20171);
or U20541 (N_20541,N_20461,N_20428);
nor U20542 (N_20542,N_20151,N_20341);
or U20543 (N_20543,N_20126,N_20376);
or U20544 (N_20544,N_20039,N_20474);
nand U20545 (N_20545,N_20353,N_20140);
and U20546 (N_20546,N_20130,N_20012);
or U20547 (N_20547,N_20247,N_20485);
xor U20548 (N_20548,N_20429,N_20479);
nor U20549 (N_20549,N_20473,N_20196);
nand U20550 (N_20550,N_20208,N_20124);
nand U20551 (N_20551,N_20221,N_20026);
or U20552 (N_20552,N_20436,N_20231);
nand U20553 (N_20553,N_20233,N_20426);
nand U20554 (N_20554,N_20185,N_20051);
nor U20555 (N_20555,N_20164,N_20225);
or U20556 (N_20556,N_20205,N_20325);
nand U20557 (N_20557,N_20040,N_20005);
nor U20558 (N_20558,N_20491,N_20191);
and U20559 (N_20559,N_20193,N_20253);
or U20560 (N_20560,N_20072,N_20498);
xor U20561 (N_20561,N_20405,N_20286);
nor U20562 (N_20562,N_20101,N_20194);
nor U20563 (N_20563,N_20117,N_20168);
nor U20564 (N_20564,N_20268,N_20343);
nor U20565 (N_20565,N_20493,N_20161);
or U20566 (N_20566,N_20105,N_20224);
nand U20567 (N_20567,N_20295,N_20227);
nor U20568 (N_20568,N_20034,N_20406);
nand U20569 (N_20569,N_20109,N_20319);
xor U20570 (N_20570,N_20088,N_20477);
nor U20571 (N_20571,N_20239,N_20007);
and U20572 (N_20572,N_20183,N_20282);
and U20573 (N_20573,N_20158,N_20066);
nand U20574 (N_20574,N_20480,N_20293);
nor U20575 (N_20575,N_20334,N_20053);
and U20576 (N_20576,N_20311,N_20338);
xor U20577 (N_20577,N_20154,N_20241);
xor U20578 (N_20578,N_20081,N_20032);
or U20579 (N_20579,N_20269,N_20178);
xnor U20580 (N_20580,N_20444,N_20035);
and U20581 (N_20581,N_20305,N_20455);
and U20582 (N_20582,N_20372,N_20058);
nand U20583 (N_20583,N_20112,N_20244);
nor U20584 (N_20584,N_20450,N_20270);
or U20585 (N_20585,N_20478,N_20492);
xor U20586 (N_20586,N_20379,N_20254);
and U20587 (N_20587,N_20437,N_20195);
or U20588 (N_20588,N_20467,N_20162);
nor U20589 (N_20589,N_20496,N_20389);
and U20590 (N_20590,N_20210,N_20095);
xor U20591 (N_20591,N_20261,N_20192);
nor U20592 (N_20592,N_20133,N_20013);
nor U20593 (N_20593,N_20055,N_20336);
nor U20594 (N_20594,N_20454,N_20441);
nor U20595 (N_20595,N_20136,N_20288);
nand U20596 (N_20596,N_20187,N_20327);
and U20597 (N_20597,N_20422,N_20345);
xnor U20598 (N_20598,N_20218,N_20307);
or U20599 (N_20599,N_20220,N_20022);
nor U20600 (N_20600,N_20069,N_20383);
and U20601 (N_20601,N_20344,N_20243);
nand U20602 (N_20602,N_20141,N_20078);
nand U20603 (N_20603,N_20279,N_20188);
xor U20604 (N_20604,N_20104,N_20110);
and U20605 (N_20605,N_20263,N_20127);
and U20606 (N_20606,N_20303,N_20285);
nor U20607 (N_20607,N_20177,N_20278);
xor U20608 (N_20608,N_20476,N_20116);
and U20609 (N_20609,N_20329,N_20020);
nor U20610 (N_20610,N_20424,N_20302);
or U20611 (N_20611,N_20294,N_20173);
nand U20612 (N_20612,N_20407,N_20371);
nand U20613 (N_20613,N_20355,N_20103);
xnor U20614 (N_20614,N_20060,N_20309);
or U20615 (N_20615,N_20023,N_20075);
xor U20616 (N_20616,N_20202,N_20453);
or U20617 (N_20617,N_20167,N_20310);
or U20618 (N_20618,N_20018,N_20318);
nor U20619 (N_20619,N_20392,N_20114);
nor U20620 (N_20620,N_20403,N_20382);
or U20621 (N_20621,N_20251,N_20071);
or U20622 (N_20622,N_20118,N_20120);
xnor U20623 (N_20623,N_20246,N_20331);
xnor U20624 (N_20624,N_20347,N_20050);
or U20625 (N_20625,N_20460,N_20409);
xor U20626 (N_20626,N_20153,N_20157);
nand U20627 (N_20627,N_20434,N_20396);
and U20628 (N_20628,N_20456,N_20084);
nand U20629 (N_20629,N_20156,N_20135);
xnor U20630 (N_20630,N_20240,N_20272);
and U20631 (N_20631,N_20198,N_20024);
nand U20632 (N_20632,N_20229,N_20209);
xnor U20633 (N_20633,N_20447,N_20385);
and U20634 (N_20634,N_20259,N_20096);
xor U20635 (N_20635,N_20300,N_20342);
xor U20636 (N_20636,N_20332,N_20427);
and U20637 (N_20637,N_20408,N_20235);
or U20638 (N_20638,N_20122,N_20179);
or U20639 (N_20639,N_20090,N_20200);
or U20640 (N_20640,N_20445,N_20367);
nor U20641 (N_20641,N_20398,N_20150);
xor U20642 (N_20642,N_20333,N_20093);
or U20643 (N_20643,N_20264,N_20180);
nand U20644 (N_20644,N_20438,N_20337);
and U20645 (N_20645,N_20145,N_20175);
or U20646 (N_20646,N_20381,N_20322);
xnor U20647 (N_20647,N_20349,N_20487);
or U20648 (N_20648,N_20068,N_20139);
and U20649 (N_20649,N_20423,N_20365);
and U20650 (N_20650,N_20181,N_20119);
and U20651 (N_20651,N_20049,N_20000);
and U20652 (N_20652,N_20292,N_20419);
nor U20653 (N_20653,N_20137,N_20413);
and U20654 (N_20654,N_20215,N_20388);
xnor U20655 (N_20655,N_20417,N_20076);
nand U20656 (N_20656,N_20172,N_20001);
nor U20657 (N_20657,N_20308,N_20025);
nor U20658 (N_20658,N_20121,N_20097);
xnor U20659 (N_20659,N_20028,N_20091);
and U20660 (N_20660,N_20165,N_20497);
nand U20661 (N_20661,N_20363,N_20439);
and U20662 (N_20662,N_20087,N_20340);
or U20663 (N_20663,N_20316,N_20062);
or U20664 (N_20664,N_20463,N_20312);
and U20665 (N_20665,N_20242,N_20236);
or U20666 (N_20666,N_20470,N_20364);
or U20667 (N_20667,N_20197,N_20380);
and U20668 (N_20668,N_20163,N_20395);
or U20669 (N_20669,N_20237,N_20330);
and U20670 (N_20670,N_20290,N_20390);
nor U20671 (N_20671,N_20174,N_20266);
xnor U20672 (N_20672,N_20361,N_20129);
nand U20673 (N_20673,N_20354,N_20368);
nor U20674 (N_20674,N_20391,N_20275);
nor U20675 (N_20675,N_20362,N_20465);
and U20676 (N_20676,N_20435,N_20052);
xnor U20677 (N_20677,N_20065,N_20080);
and U20678 (N_20678,N_20134,N_20042);
or U20679 (N_20679,N_20113,N_20299);
nor U20680 (N_20680,N_20471,N_20384);
and U20681 (N_20681,N_20002,N_20262);
xnor U20682 (N_20682,N_20255,N_20143);
nand U20683 (N_20683,N_20466,N_20256);
nor U20684 (N_20684,N_20061,N_20206);
xnor U20685 (N_20685,N_20250,N_20416);
nor U20686 (N_20686,N_20044,N_20082);
nor U20687 (N_20687,N_20015,N_20265);
nor U20688 (N_20688,N_20415,N_20189);
or U20689 (N_20689,N_20375,N_20452);
nor U20690 (N_20690,N_20274,N_20211);
and U20691 (N_20691,N_20313,N_20442);
nand U20692 (N_20692,N_20226,N_20411);
or U20693 (N_20693,N_20469,N_20433);
nand U20694 (N_20694,N_20486,N_20449);
and U20695 (N_20695,N_20128,N_20070);
nand U20696 (N_20696,N_20351,N_20169);
xor U20697 (N_20697,N_20111,N_20089);
xor U20698 (N_20698,N_20213,N_20030);
nor U20699 (N_20699,N_20458,N_20495);
or U20700 (N_20700,N_20166,N_20421);
nor U20701 (N_20701,N_20410,N_20046);
nor U20702 (N_20702,N_20289,N_20402);
and U20703 (N_20703,N_20207,N_20276);
nand U20704 (N_20704,N_20008,N_20031);
or U20705 (N_20705,N_20125,N_20219);
nor U20706 (N_20706,N_20399,N_20147);
xor U20707 (N_20707,N_20190,N_20431);
nor U20708 (N_20708,N_20446,N_20073);
and U20709 (N_20709,N_20317,N_20412);
and U20710 (N_20710,N_20059,N_20027);
nor U20711 (N_20711,N_20100,N_20281);
xor U20712 (N_20712,N_20108,N_20320);
or U20713 (N_20713,N_20131,N_20306);
nand U20714 (N_20714,N_20420,N_20083);
and U20715 (N_20715,N_20106,N_20249);
and U20716 (N_20716,N_20366,N_20252);
and U20717 (N_20717,N_20045,N_20216);
and U20718 (N_20718,N_20186,N_20321);
xor U20719 (N_20719,N_20011,N_20326);
xnor U20720 (N_20720,N_20484,N_20176);
or U20721 (N_20721,N_20358,N_20378);
nor U20722 (N_20722,N_20182,N_20152);
xor U20723 (N_20723,N_20021,N_20067);
or U20724 (N_20724,N_20260,N_20277);
and U20725 (N_20725,N_20346,N_20004);
nor U20726 (N_20726,N_20056,N_20373);
or U20727 (N_20727,N_20284,N_20017);
xnor U20728 (N_20728,N_20079,N_20234);
xor U20729 (N_20729,N_20440,N_20102);
nand U20730 (N_20730,N_20094,N_20144);
xor U20731 (N_20731,N_20488,N_20036);
and U20732 (N_20732,N_20280,N_20451);
nor U20733 (N_20733,N_20107,N_20212);
nor U20734 (N_20734,N_20483,N_20092);
and U20735 (N_20735,N_20142,N_20443);
nand U20736 (N_20736,N_20132,N_20085);
or U20737 (N_20737,N_20468,N_20472);
or U20738 (N_20738,N_20370,N_20230);
and U20739 (N_20739,N_20019,N_20360);
nand U20740 (N_20740,N_20043,N_20430);
or U20741 (N_20741,N_20029,N_20170);
nand U20742 (N_20742,N_20064,N_20448);
nand U20743 (N_20743,N_20204,N_20400);
nor U20744 (N_20744,N_20328,N_20357);
or U20745 (N_20745,N_20494,N_20348);
nor U20746 (N_20746,N_20098,N_20386);
and U20747 (N_20747,N_20296,N_20099);
or U20748 (N_20748,N_20481,N_20003);
nand U20749 (N_20749,N_20324,N_20499);
or U20750 (N_20750,N_20031,N_20412);
xor U20751 (N_20751,N_20328,N_20228);
and U20752 (N_20752,N_20226,N_20076);
nand U20753 (N_20753,N_20385,N_20365);
nand U20754 (N_20754,N_20419,N_20353);
and U20755 (N_20755,N_20258,N_20035);
nor U20756 (N_20756,N_20431,N_20039);
or U20757 (N_20757,N_20195,N_20094);
nand U20758 (N_20758,N_20402,N_20290);
or U20759 (N_20759,N_20177,N_20154);
or U20760 (N_20760,N_20286,N_20276);
nand U20761 (N_20761,N_20458,N_20056);
nand U20762 (N_20762,N_20027,N_20428);
nor U20763 (N_20763,N_20185,N_20030);
and U20764 (N_20764,N_20045,N_20354);
and U20765 (N_20765,N_20225,N_20059);
or U20766 (N_20766,N_20326,N_20007);
xnor U20767 (N_20767,N_20318,N_20326);
nor U20768 (N_20768,N_20140,N_20069);
nor U20769 (N_20769,N_20465,N_20346);
or U20770 (N_20770,N_20115,N_20000);
or U20771 (N_20771,N_20448,N_20161);
nand U20772 (N_20772,N_20464,N_20461);
or U20773 (N_20773,N_20260,N_20443);
and U20774 (N_20774,N_20296,N_20453);
nand U20775 (N_20775,N_20234,N_20028);
and U20776 (N_20776,N_20187,N_20261);
nor U20777 (N_20777,N_20194,N_20148);
nand U20778 (N_20778,N_20004,N_20329);
xor U20779 (N_20779,N_20298,N_20413);
or U20780 (N_20780,N_20279,N_20341);
nor U20781 (N_20781,N_20445,N_20180);
and U20782 (N_20782,N_20073,N_20447);
and U20783 (N_20783,N_20017,N_20313);
nor U20784 (N_20784,N_20141,N_20454);
or U20785 (N_20785,N_20413,N_20387);
or U20786 (N_20786,N_20094,N_20423);
and U20787 (N_20787,N_20254,N_20423);
nand U20788 (N_20788,N_20003,N_20286);
nor U20789 (N_20789,N_20409,N_20283);
or U20790 (N_20790,N_20446,N_20153);
nor U20791 (N_20791,N_20228,N_20101);
nor U20792 (N_20792,N_20208,N_20048);
nand U20793 (N_20793,N_20052,N_20050);
nor U20794 (N_20794,N_20221,N_20042);
nand U20795 (N_20795,N_20450,N_20218);
nand U20796 (N_20796,N_20352,N_20089);
xor U20797 (N_20797,N_20158,N_20313);
nor U20798 (N_20798,N_20073,N_20127);
nand U20799 (N_20799,N_20021,N_20310);
nor U20800 (N_20800,N_20331,N_20129);
and U20801 (N_20801,N_20031,N_20457);
nor U20802 (N_20802,N_20275,N_20454);
and U20803 (N_20803,N_20062,N_20296);
and U20804 (N_20804,N_20191,N_20042);
or U20805 (N_20805,N_20167,N_20268);
xor U20806 (N_20806,N_20358,N_20217);
nor U20807 (N_20807,N_20164,N_20173);
xor U20808 (N_20808,N_20477,N_20466);
nor U20809 (N_20809,N_20212,N_20384);
or U20810 (N_20810,N_20186,N_20205);
or U20811 (N_20811,N_20179,N_20380);
nand U20812 (N_20812,N_20484,N_20231);
nand U20813 (N_20813,N_20078,N_20106);
nand U20814 (N_20814,N_20008,N_20479);
xor U20815 (N_20815,N_20072,N_20112);
and U20816 (N_20816,N_20367,N_20328);
nand U20817 (N_20817,N_20014,N_20419);
nor U20818 (N_20818,N_20333,N_20325);
or U20819 (N_20819,N_20158,N_20023);
nor U20820 (N_20820,N_20251,N_20051);
and U20821 (N_20821,N_20490,N_20288);
or U20822 (N_20822,N_20101,N_20410);
xnor U20823 (N_20823,N_20198,N_20205);
and U20824 (N_20824,N_20022,N_20316);
and U20825 (N_20825,N_20260,N_20242);
and U20826 (N_20826,N_20493,N_20019);
xnor U20827 (N_20827,N_20108,N_20028);
or U20828 (N_20828,N_20141,N_20321);
or U20829 (N_20829,N_20310,N_20384);
or U20830 (N_20830,N_20409,N_20466);
or U20831 (N_20831,N_20474,N_20400);
and U20832 (N_20832,N_20032,N_20396);
nand U20833 (N_20833,N_20271,N_20108);
nand U20834 (N_20834,N_20456,N_20211);
nand U20835 (N_20835,N_20201,N_20267);
nor U20836 (N_20836,N_20247,N_20452);
and U20837 (N_20837,N_20178,N_20056);
nand U20838 (N_20838,N_20280,N_20460);
or U20839 (N_20839,N_20180,N_20259);
xnor U20840 (N_20840,N_20128,N_20469);
nand U20841 (N_20841,N_20049,N_20003);
nand U20842 (N_20842,N_20284,N_20148);
xor U20843 (N_20843,N_20035,N_20368);
and U20844 (N_20844,N_20111,N_20393);
or U20845 (N_20845,N_20335,N_20478);
nor U20846 (N_20846,N_20342,N_20140);
xor U20847 (N_20847,N_20301,N_20076);
and U20848 (N_20848,N_20280,N_20471);
or U20849 (N_20849,N_20138,N_20075);
nand U20850 (N_20850,N_20428,N_20441);
nand U20851 (N_20851,N_20344,N_20115);
nand U20852 (N_20852,N_20059,N_20313);
or U20853 (N_20853,N_20076,N_20268);
xor U20854 (N_20854,N_20262,N_20407);
and U20855 (N_20855,N_20176,N_20253);
nor U20856 (N_20856,N_20226,N_20123);
nor U20857 (N_20857,N_20080,N_20293);
xnor U20858 (N_20858,N_20288,N_20191);
nor U20859 (N_20859,N_20126,N_20300);
xor U20860 (N_20860,N_20136,N_20314);
xor U20861 (N_20861,N_20189,N_20068);
or U20862 (N_20862,N_20452,N_20382);
xor U20863 (N_20863,N_20390,N_20312);
nor U20864 (N_20864,N_20172,N_20275);
or U20865 (N_20865,N_20107,N_20269);
nor U20866 (N_20866,N_20308,N_20215);
xnor U20867 (N_20867,N_20160,N_20368);
nand U20868 (N_20868,N_20011,N_20199);
nand U20869 (N_20869,N_20018,N_20429);
or U20870 (N_20870,N_20131,N_20317);
nor U20871 (N_20871,N_20456,N_20185);
xnor U20872 (N_20872,N_20374,N_20080);
and U20873 (N_20873,N_20103,N_20417);
nor U20874 (N_20874,N_20348,N_20322);
or U20875 (N_20875,N_20409,N_20023);
or U20876 (N_20876,N_20017,N_20183);
and U20877 (N_20877,N_20005,N_20083);
nand U20878 (N_20878,N_20158,N_20437);
nor U20879 (N_20879,N_20354,N_20334);
or U20880 (N_20880,N_20212,N_20073);
nor U20881 (N_20881,N_20105,N_20125);
xnor U20882 (N_20882,N_20424,N_20017);
and U20883 (N_20883,N_20433,N_20094);
xnor U20884 (N_20884,N_20458,N_20004);
nand U20885 (N_20885,N_20349,N_20370);
nand U20886 (N_20886,N_20189,N_20157);
and U20887 (N_20887,N_20311,N_20453);
nor U20888 (N_20888,N_20058,N_20477);
nand U20889 (N_20889,N_20214,N_20210);
and U20890 (N_20890,N_20445,N_20439);
nand U20891 (N_20891,N_20119,N_20070);
xor U20892 (N_20892,N_20283,N_20082);
xnor U20893 (N_20893,N_20473,N_20466);
xnor U20894 (N_20894,N_20437,N_20291);
nor U20895 (N_20895,N_20286,N_20355);
or U20896 (N_20896,N_20260,N_20028);
xnor U20897 (N_20897,N_20045,N_20167);
or U20898 (N_20898,N_20309,N_20139);
xnor U20899 (N_20899,N_20297,N_20428);
nor U20900 (N_20900,N_20245,N_20122);
and U20901 (N_20901,N_20467,N_20364);
or U20902 (N_20902,N_20482,N_20120);
nor U20903 (N_20903,N_20301,N_20411);
or U20904 (N_20904,N_20233,N_20052);
xor U20905 (N_20905,N_20072,N_20085);
nand U20906 (N_20906,N_20101,N_20407);
nand U20907 (N_20907,N_20167,N_20273);
nor U20908 (N_20908,N_20407,N_20300);
or U20909 (N_20909,N_20354,N_20459);
and U20910 (N_20910,N_20237,N_20462);
or U20911 (N_20911,N_20309,N_20407);
nand U20912 (N_20912,N_20371,N_20195);
and U20913 (N_20913,N_20399,N_20388);
and U20914 (N_20914,N_20370,N_20356);
and U20915 (N_20915,N_20162,N_20003);
or U20916 (N_20916,N_20377,N_20024);
or U20917 (N_20917,N_20078,N_20032);
xnor U20918 (N_20918,N_20036,N_20120);
and U20919 (N_20919,N_20036,N_20281);
nand U20920 (N_20920,N_20015,N_20492);
nor U20921 (N_20921,N_20324,N_20259);
or U20922 (N_20922,N_20275,N_20165);
nand U20923 (N_20923,N_20259,N_20045);
and U20924 (N_20924,N_20150,N_20051);
nand U20925 (N_20925,N_20340,N_20277);
nand U20926 (N_20926,N_20065,N_20292);
nand U20927 (N_20927,N_20294,N_20457);
xor U20928 (N_20928,N_20221,N_20267);
nor U20929 (N_20929,N_20086,N_20005);
nor U20930 (N_20930,N_20392,N_20414);
or U20931 (N_20931,N_20028,N_20451);
or U20932 (N_20932,N_20068,N_20452);
or U20933 (N_20933,N_20208,N_20272);
nand U20934 (N_20934,N_20268,N_20273);
or U20935 (N_20935,N_20002,N_20123);
and U20936 (N_20936,N_20447,N_20212);
xor U20937 (N_20937,N_20209,N_20332);
or U20938 (N_20938,N_20129,N_20442);
xnor U20939 (N_20939,N_20135,N_20289);
nor U20940 (N_20940,N_20278,N_20074);
or U20941 (N_20941,N_20142,N_20086);
and U20942 (N_20942,N_20099,N_20193);
or U20943 (N_20943,N_20028,N_20084);
nor U20944 (N_20944,N_20255,N_20297);
xnor U20945 (N_20945,N_20102,N_20002);
and U20946 (N_20946,N_20455,N_20373);
nand U20947 (N_20947,N_20378,N_20275);
xnor U20948 (N_20948,N_20207,N_20386);
nor U20949 (N_20949,N_20393,N_20462);
and U20950 (N_20950,N_20026,N_20080);
nor U20951 (N_20951,N_20177,N_20112);
nand U20952 (N_20952,N_20343,N_20452);
xnor U20953 (N_20953,N_20449,N_20464);
xor U20954 (N_20954,N_20009,N_20080);
nor U20955 (N_20955,N_20285,N_20362);
nor U20956 (N_20956,N_20007,N_20224);
nand U20957 (N_20957,N_20046,N_20367);
or U20958 (N_20958,N_20007,N_20156);
or U20959 (N_20959,N_20465,N_20147);
or U20960 (N_20960,N_20107,N_20135);
nor U20961 (N_20961,N_20125,N_20129);
xor U20962 (N_20962,N_20140,N_20197);
xnor U20963 (N_20963,N_20484,N_20012);
nand U20964 (N_20964,N_20385,N_20361);
nor U20965 (N_20965,N_20429,N_20085);
nor U20966 (N_20966,N_20335,N_20169);
or U20967 (N_20967,N_20186,N_20124);
xor U20968 (N_20968,N_20017,N_20486);
or U20969 (N_20969,N_20097,N_20054);
or U20970 (N_20970,N_20032,N_20458);
or U20971 (N_20971,N_20358,N_20298);
nand U20972 (N_20972,N_20137,N_20028);
or U20973 (N_20973,N_20089,N_20373);
or U20974 (N_20974,N_20110,N_20323);
xnor U20975 (N_20975,N_20342,N_20147);
xor U20976 (N_20976,N_20230,N_20302);
nor U20977 (N_20977,N_20236,N_20100);
xnor U20978 (N_20978,N_20203,N_20093);
nor U20979 (N_20979,N_20358,N_20240);
and U20980 (N_20980,N_20107,N_20307);
nand U20981 (N_20981,N_20248,N_20169);
nand U20982 (N_20982,N_20055,N_20051);
nand U20983 (N_20983,N_20312,N_20343);
and U20984 (N_20984,N_20078,N_20203);
and U20985 (N_20985,N_20268,N_20092);
or U20986 (N_20986,N_20120,N_20350);
or U20987 (N_20987,N_20156,N_20222);
nand U20988 (N_20988,N_20191,N_20206);
xnor U20989 (N_20989,N_20397,N_20223);
nor U20990 (N_20990,N_20295,N_20443);
and U20991 (N_20991,N_20258,N_20297);
xnor U20992 (N_20992,N_20247,N_20416);
and U20993 (N_20993,N_20420,N_20246);
nor U20994 (N_20994,N_20428,N_20345);
xnor U20995 (N_20995,N_20276,N_20362);
or U20996 (N_20996,N_20201,N_20098);
xor U20997 (N_20997,N_20083,N_20464);
or U20998 (N_20998,N_20029,N_20228);
xnor U20999 (N_20999,N_20393,N_20338);
nand U21000 (N_21000,N_20841,N_20984);
xor U21001 (N_21001,N_20670,N_20934);
xor U21002 (N_21002,N_20528,N_20625);
and U21003 (N_21003,N_20777,N_20734);
nand U21004 (N_21004,N_20909,N_20659);
xnor U21005 (N_21005,N_20719,N_20683);
nor U21006 (N_21006,N_20970,N_20703);
nand U21007 (N_21007,N_20839,N_20940);
and U21008 (N_21008,N_20722,N_20891);
nand U21009 (N_21009,N_20557,N_20791);
nand U21010 (N_21010,N_20564,N_20926);
or U21011 (N_21011,N_20827,N_20952);
nor U21012 (N_21012,N_20639,N_20662);
nor U21013 (N_21013,N_20716,N_20942);
nor U21014 (N_21014,N_20559,N_20663);
nor U21015 (N_21015,N_20938,N_20987);
nand U21016 (N_21016,N_20798,N_20968);
nor U21017 (N_21017,N_20994,N_20515);
and U21018 (N_21018,N_20961,N_20573);
nand U21019 (N_21019,N_20972,N_20910);
nand U21020 (N_21020,N_20580,N_20503);
and U21021 (N_21021,N_20854,N_20561);
xnor U21022 (N_21022,N_20989,N_20999);
nor U21023 (N_21023,N_20852,N_20792);
nand U21024 (N_21024,N_20634,N_20983);
and U21025 (N_21025,N_20894,N_20523);
or U21026 (N_21026,N_20607,N_20705);
xor U21027 (N_21027,N_20697,N_20500);
or U21028 (N_21028,N_20700,N_20554);
nor U21029 (N_21029,N_20981,N_20600);
nand U21030 (N_21030,N_20933,N_20855);
xnor U21031 (N_21031,N_20743,N_20847);
nand U21032 (N_21032,N_20589,N_20951);
or U21033 (N_21033,N_20566,N_20982);
nand U21034 (N_21034,N_20714,N_20737);
xnor U21035 (N_21035,N_20995,N_20651);
and U21036 (N_21036,N_20755,N_20797);
and U21037 (N_21037,N_20794,N_20789);
or U21038 (N_21038,N_20832,N_20635);
or U21039 (N_21039,N_20907,N_20867);
nor U21040 (N_21040,N_20885,N_20581);
or U21041 (N_21041,N_20537,N_20686);
or U21042 (N_21042,N_20658,N_20930);
xor U21043 (N_21043,N_20502,N_20807);
nor U21044 (N_21044,N_20853,N_20936);
xnor U21045 (N_21045,N_20617,N_20753);
xor U21046 (N_21046,N_20920,N_20610);
nand U21047 (N_21047,N_20598,N_20612);
nor U21048 (N_21048,N_20766,N_20547);
xnor U21049 (N_21049,N_20908,N_20551);
or U21050 (N_21050,N_20601,N_20943);
nand U21051 (N_21051,N_20979,N_20870);
or U21052 (N_21052,N_20991,N_20747);
and U21053 (N_21053,N_20882,N_20988);
xor U21054 (N_21054,N_20896,N_20849);
or U21055 (N_21055,N_20819,N_20821);
and U21056 (N_21056,N_20919,N_20548);
and U21057 (N_21057,N_20965,N_20895);
nand U21058 (N_21058,N_20623,N_20869);
and U21059 (N_21059,N_20680,N_20518);
and U21060 (N_21060,N_20558,N_20775);
and U21061 (N_21061,N_20825,N_20699);
xor U21062 (N_21062,N_20615,N_20517);
and U21063 (N_21063,N_20893,N_20715);
nand U21064 (N_21064,N_20721,N_20770);
nand U21065 (N_21065,N_20980,N_20949);
and U21066 (N_21066,N_20552,N_20532);
or U21067 (N_21067,N_20521,N_20652);
xor U21068 (N_21068,N_20871,N_20897);
and U21069 (N_21069,N_20831,N_20687);
xor U21070 (N_21070,N_20866,N_20509);
nand U21071 (N_21071,N_20993,N_20595);
and U21072 (N_21072,N_20728,N_20860);
nand U21073 (N_21073,N_20813,N_20768);
nor U21074 (N_21074,N_20875,N_20591);
and U21075 (N_21075,N_20778,N_20932);
and U21076 (N_21076,N_20585,N_20750);
xnor U21077 (N_21077,N_20837,N_20584);
nand U21078 (N_21078,N_20536,N_20742);
or U21079 (N_21079,N_20929,N_20917);
nor U21080 (N_21080,N_20850,N_20935);
xor U21081 (N_21081,N_20643,N_20784);
nand U21082 (N_21082,N_20619,N_20783);
nand U21083 (N_21083,N_20726,N_20709);
and U21084 (N_21084,N_20960,N_20512);
and U21085 (N_21085,N_20824,N_20758);
or U21086 (N_21086,N_20710,N_20818);
nand U21087 (N_21087,N_20539,N_20641);
or U21088 (N_21088,N_20801,N_20673);
and U21089 (N_21089,N_20906,N_20959);
or U21090 (N_21090,N_20859,N_20508);
or U21091 (N_21091,N_20505,N_20796);
or U21092 (N_21092,N_20803,N_20542);
nor U21093 (N_21093,N_20540,N_20974);
xnor U21094 (N_21094,N_20717,N_20514);
nor U21095 (N_21095,N_20749,N_20513);
and U21096 (N_21096,N_20773,N_20937);
and U21097 (N_21097,N_20668,N_20681);
or U21098 (N_21098,N_20614,N_20820);
nor U21099 (N_21099,N_20953,N_20605);
nand U21100 (N_21100,N_20571,N_20724);
nor U21101 (N_21101,N_20956,N_20975);
nand U21102 (N_21102,N_20918,N_20772);
or U21103 (N_21103,N_20708,N_20622);
nor U21104 (N_21104,N_20568,N_20701);
xnor U21105 (N_21105,N_20694,N_20613);
or U21106 (N_21106,N_20915,N_20712);
xnor U21107 (N_21107,N_20696,N_20881);
and U21108 (N_21108,N_20997,N_20851);
or U21109 (N_21109,N_20744,N_20575);
xnor U21110 (N_21110,N_20901,N_20780);
nand U21111 (N_21111,N_20624,N_20690);
or U21112 (N_21112,N_20550,N_20762);
or U21113 (N_21113,N_20544,N_20977);
nand U21114 (N_21114,N_20606,N_20725);
and U21115 (N_21115,N_20525,N_20732);
or U21116 (N_21116,N_20657,N_20998);
xnor U21117 (N_21117,N_20948,N_20654);
nor U21118 (N_21118,N_20966,N_20964);
or U21119 (N_21119,N_20609,N_20834);
nor U21120 (N_21120,N_20905,N_20805);
xor U21121 (N_21121,N_20769,N_20620);
nor U21122 (N_21122,N_20863,N_20611);
and U21123 (N_21123,N_20817,N_20782);
nand U21124 (N_21124,N_20946,N_20592);
nor U21125 (N_21125,N_20857,N_20602);
nor U21126 (N_21126,N_20793,N_20745);
xnor U21127 (N_21127,N_20648,N_20752);
and U21128 (N_21128,N_20692,N_20858);
and U21129 (N_21129,N_20604,N_20939);
and U21130 (N_21130,N_20771,N_20608);
xnor U21131 (N_21131,N_20815,N_20963);
nor U21132 (N_21132,N_20636,N_20921);
or U21133 (N_21133,N_20923,N_20947);
nand U21134 (N_21134,N_20653,N_20671);
nand U21135 (N_21135,N_20883,N_20957);
xor U21136 (N_21136,N_20836,N_20637);
xor U21137 (N_21137,N_20674,N_20931);
xor U21138 (N_21138,N_20877,N_20814);
and U21139 (N_21139,N_20914,N_20578);
nand U21140 (N_21140,N_20546,N_20629);
and U21141 (N_21141,N_20644,N_20695);
nor U21142 (N_21142,N_20757,N_20520);
and U21143 (N_21143,N_20735,N_20844);
nor U21144 (N_21144,N_20835,N_20976);
xor U21145 (N_21145,N_20626,N_20678);
nor U21146 (N_21146,N_20675,N_20543);
nand U21147 (N_21147,N_20685,N_20810);
xor U21148 (N_21148,N_20565,N_20524);
nand U21149 (N_21149,N_20630,N_20656);
xor U21150 (N_21150,N_20779,N_20872);
or U21151 (N_21151,N_20638,N_20927);
or U21152 (N_21152,N_20698,N_20787);
nor U21153 (N_21153,N_20822,N_20902);
nor U21154 (N_21154,N_20913,N_20527);
nand U21155 (N_21155,N_20996,N_20603);
or U21156 (N_21156,N_20761,N_20774);
and U21157 (N_21157,N_20799,N_20838);
or U21158 (N_21158,N_20868,N_20884);
and U21159 (N_21159,N_20655,N_20567);
nor U21160 (N_21160,N_20616,N_20873);
nor U21161 (N_21161,N_20765,N_20900);
and U21162 (N_21162,N_20516,N_20806);
xnor U21163 (N_21163,N_20583,N_20950);
or U21164 (N_21164,N_20955,N_20553);
nor U21165 (N_21165,N_20978,N_20519);
and U21166 (N_21166,N_20691,N_20945);
xnor U21167 (N_21167,N_20865,N_20647);
and U21168 (N_21168,N_20706,N_20862);
and U21169 (N_21169,N_20941,N_20577);
or U21170 (N_21170,N_20534,N_20985);
nor U21171 (N_21171,N_20723,N_20800);
and U21172 (N_21172,N_20861,N_20666);
and U21173 (N_21173,N_20899,N_20535);
xnor U21174 (N_21174,N_20590,N_20848);
nor U21175 (N_21175,N_20594,N_20618);
and U21176 (N_21176,N_20597,N_20530);
nand U21177 (N_21177,N_20642,N_20628);
nand U21178 (N_21178,N_20828,N_20533);
nand U21179 (N_21179,N_20621,N_20510);
nor U21180 (N_21180,N_20730,N_20746);
xnor U21181 (N_21181,N_20788,N_20511);
nand U21182 (N_21182,N_20785,N_20888);
nand U21183 (N_21183,N_20627,N_20763);
or U21184 (N_21184,N_20645,N_20556);
xor U21185 (N_21185,N_20689,N_20713);
nor U21186 (N_21186,N_20633,N_20596);
or U21187 (N_21187,N_20661,N_20588);
xor U21188 (N_21188,N_20579,N_20593);
nor U21189 (N_21189,N_20632,N_20912);
xor U21190 (N_21190,N_20876,N_20846);
and U21191 (N_21191,N_20676,N_20576);
nand U21192 (N_21192,N_20973,N_20986);
and U21193 (N_21193,N_20741,N_20808);
xor U21194 (N_21194,N_20954,N_20925);
or U21195 (N_21195,N_20679,N_20887);
xnor U21196 (N_21196,N_20572,N_20754);
nand U21197 (N_21197,N_20856,N_20504);
xnor U21198 (N_21198,N_20879,N_20677);
or U21199 (N_21199,N_20830,N_20911);
and U21200 (N_21200,N_20971,N_20751);
nand U21201 (N_21201,N_20992,N_20874);
and U21202 (N_21202,N_20560,N_20760);
or U21203 (N_21203,N_20812,N_20727);
nor U21204 (N_21204,N_20693,N_20702);
and U21205 (N_21205,N_20833,N_20506);
nand U21206 (N_21206,N_20878,N_20748);
and U21207 (N_21207,N_20843,N_20649);
xnor U21208 (N_21208,N_20664,N_20507);
or U21209 (N_21209,N_20924,N_20574);
or U21210 (N_21210,N_20587,N_20903);
and U21211 (N_21211,N_20672,N_20707);
nand U21212 (N_21212,N_20667,N_20786);
and U21213 (N_21213,N_20809,N_20684);
nor U21214 (N_21214,N_20682,N_20570);
or U21215 (N_21215,N_20890,N_20916);
or U21216 (N_21216,N_20545,N_20549);
xor U21217 (N_21217,N_20880,N_20740);
or U21218 (N_21218,N_20767,N_20711);
xnor U21219 (N_21219,N_20733,N_20736);
or U21220 (N_21220,N_20764,N_20898);
or U21221 (N_21221,N_20718,N_20660);
nand U21222 (N_21222,N_20776,N_20811);
xnor U21223 (N_21223,N_20720,N_20738);
and U21224 (N_21224,N_20795,N_20665);
or U21225 (N_21225,N_20631,N_20790);
and U21226 (N_21226,N_20704,N_20688);
nor U21227 (N_21227,N_20845,N_20967);
and U21228 (N_21228,N_20729,N_20640);
nor U21229 (N_21229,N_20759,N_20646);
or U21230 (N_21230,N_20840,N_20526);
and U21231 (N_21231,N_20731,N_20886);
or U21232 (N_21232,N_20944,N_20563);
nand U21233 (N_21233,N_20781,N_20756);
xor U21234 (N_21234,N_20531,N_20555);
nor U21235 (N_21235,N_20928,N_20842);
nor U21236 (N_21236,N_20599,N_20541);
or U21237 (N_21237,N_20892,N_20802);
or U21238 (N_21238,N_20969,N_20826);
and U21239 (N_21239,N_20829,N_20669);
or U21240 (N_21240,N_20922,N_20501);
or U21241 (N_21241,N_20958,N_20522);
or U21242 (N_21242,N_20889,N_20562);
or U21243 (N_21243,N_20823,N_20569);
and U21244 (N_21244,N_20864,N_20650);
nand U21245 (N_21245,N_20538,N_20739);
nand U21246 (N_21246,N_20816,N_20904);
xor U21247 (N_21247,N_20586,N_20529);
or U21248 (N_21248,N_20962,N_20804);
nor U21249 (N_21249,N_20582,N_20990);
nand U21250 (N_21250,N_20532,N_20519);
and U21251 (N_21251,N_20914,N_20853);
nor U21252 (N_21252,N_20790,N_20982);
nand U21253 (N_21253,N_20874,N_20868);
xor U21254 (N_21254,N_20760,N_20926);
and U21255 (N_21255,N_20716,N_20881);
nand U21256 (N_21256,N_20889,N_20665);
and U21257 (N_21257,N_20791,N_20951);
or U21258 (N_21258,N_20791,N_20970);
nand U21259 (N_21259,N_20830,N_20663);
xnor U21260 (N_21260,N_20784,N_20947);
nor U21261 (N_21261,N_20588,N_20675);
or U21262 (N_21262,N_20619,N_20659);
nor U21263 (N_21263,N_20529,N_20837);
nand U21264 (N_21264,N_20619,N_20868);
and U21265 (N_21265,N_20623,N_20709);
nor U21266 (N_21266,N_20619,N_20835);
xnor U21267 (N_21267,N_20850,N_20602);
nand U21268 (N_21268,N_20617,N_20766);
xnor U21269 (N_21269,N_20599,N_20767);
or U21270 (N_21270,N_20653,N_20577);
or U21271 (N_21271,N_20827,N_20687);
nand U21272 (N_21272,N_20822,N_20903);
xnor U21273 (N_21273,N_20752,N_20651);
and U21274 (N_21274,N_20686,N_20669);
or U21275 (N_21275,N_20561,N_20760);
or U21276 (N_21276,N_20857,N_20583);
nand U21277 (N_21277,N_20738,N_20617);
xnor U21278 (N_21278,N_20755,N_20585);
and U21279 (N_21279,N_20679,N_20907);
and U21280 (N_21280,N_20823,N_20852);
or U21281 (N_21281,N_20631,N_20828);
nand U21282 (N_21282,N_20926,N_20520);
xnor U21283 (N_21283,N_20940,N_20784);
nand U21284 (N_21284,N_20871,N_20607);
and U21285 (N_21285,N_20718,N_20699);
nand U21286 (N_21286,N_20513,N_20715);
or U21287 (N_21287,N_20775,N_20961);
xnor U21288 (N_21288,N_20811,N_20802);
or U21289 (N_21289,N_20667,N_20614);
nor U21290 (N_21290,N_20649,N_20937);
xnor U21291 (N_21291,N_20521,N_20708);
nand U21292 (N_21292,N_20586,N_20673);
xor U21293 (N_21293,N_20574,N_20586);
nand U21294 (N_21294,N_20589,N_20929);
and U21295 (N_21295,N_20710,N_20666);
xor U21296 (N_21296,N_20551,N_20956);
or U21297 (N_21297,N_20881,N_20870);
and U21298 (N_21298,N_20729,N_20625);
or U21299 (N_21299,N_20750,N_20765);
nor U21300 (N_21300,N_20982,N_20695);
or U21301 (N_21301,N_20734,N_20543);
nor U21302 (N_21302,N_20978,N_20860);
and U21303 (N_21303,N_20680,N_20921);
or U21304 (N_21304,N_20744,N_20922);
or U21305 (N_21305,N_20785,N_20848);
or U21306 (N_21306,N_20676,N_20795);
nor U21307 (N_21307,N_20861,N_20885);
or U21308 (N_21308,N_20916,N_20900);
nor U21309 (N_21309,N_20958,N_20977);
xor U21310 (N_21310,N_20628,N_20865);
nor U21311 (N_21311,N_20808,N_20627);
nand U21312 (N_21312,N_20647,N_20791);
nand U21313 (N_21313,N_20606,N_20966);
or U21314 (N_21314,N_20776,N_20672);
xnor U21315 (N_21315,N_20865,N_20837);
or U21316 (N_21316,N_20832,N_20631);
and U21317 (N_21317,N_20844,N_20757);
and U21318 (N_21318,N_20622,N_20631);
xnor U21319 (N_21319,N_20859,N_20876);
xnor U21320 (N_21320,N_20794,N_20807);
or U21321 (N_21321,N_20848,N_20514);
xnor U21322 (N_21322,N_20862,N_20682);
nand U21323 (N_21323,N_20725,N_20855);
or U21324 (N_21324,N_20972,N_20992);
and U21325 (N_21325,N_20733,N_20944);
nand U21326 (N_21326,N_20860,N_20529);
and U21327 (N_21327,N_20650,N_20918);
or U21328 (N_21328,N_20709,N_20838);
and U21329 (N_21329,N_20778,N_20717);
and U21330 (N_21330,N_20604,N_20956);
nor U21331 (N_21331,N_20777,N_20607);
nor U21332 (N_21332,N_20685,N_20795);
xnor U21333 (N_21333,N_20728,N_20523);
xnor U21334 (N_21334,N_20573,N_20748);
xnor U21335 (N_21335,N_20803,N_20760);
nand U21336 (N_21336,N_20764,N_20548);
or U21337 (N_21337,N_20888,N_20843);
and U21338 (N_21338,N_20898,N_20891);
xnor U21339 (N_21339,N_20968,N_20762);
nor U21340 (N_21340,N_20930,N_20724);
and U21341 (N_21341,N_20692,N_20671);
nand U21342 (N_21342,N_20689,N_20853);
or U21343 (N_21343,N_20844,N_20622);
nor U21344 (N_21344,N_20635,N_20690);
and U21345 (N_21345,N_20854,N_20967);
and U21346 (N_21346,N_20628,N_20513);
nor U21347 (N_21347,N_20526,N_20630);
xnor U21348 (N_21348,N_20660,N_20844);
nor U21349 (N_21349,N_20793,N_20538);
nor U21350 (N_21350,N_20757,N_20758);
xnor U21351 (N_21351,N_20769,N_20995);
xor U21352 (N_21352,N_20719,N_20720);
and U21353 (N_21353,N_20984,N_20950);
nor U21354 (N_21354,N_20657,N_20557);
xnor U21355 (N_21355,N_20747,N_20556);
or U21356 (N_21356,N_20873,N_20940);
xor U21357 (N_21357,N_20597,N_20819);
nand U21358 (N_21358,N_20576,N_20832);
nand U21359 (N_21359,N_20633,N_20770);
or U21360 (N_21360,N_20745,N_20633);
nand U21361 (N_21361,N_20505,N_20868);
nor U21362 (N_21362,N_20958,N_20694);
nor U21363 (N_21363,N_20558,N_20910);
or U21364 (N_21364,N_20815,N_20590);
nor U21365 (N_21365,N_20718,N_20789);
xnor U21366 (N_21366,N_20549,N_20609);
or U21367 (N_21367,N_20778,N_20532);
xor U21368 (N_21368,N_20957,N_20582);
xnor U21369 (N_21369,N_20992,N_20996);
xnor U21370 (N_21370,N_20974,N_20976);
xor U21371 (N_21371,N_20579,N_20974);
nand U21372 (N_21372,N_20719,N_20562);
and U21373 (N_21373,N_20961,N_20520);
and U21374 (N_21374,N_20861,N_20572);
or U21375 (N_21375,N_20869,N_20766);
or U21376 (N_21376,N_20576,N_20972);
and U21377 (N_21377,N_20628,N_20966);
or U21378 (N_21378,N_20993,N_20533);
and U21379 (N_21379,N_20603,N_20881);
and U21380 (N_21380,N_20931,N_20710);
and U21381 (N_21381,N_20533,N_20535);
or U21382 (N_21382,N_20537,N_20798);
nand U21383 (N_21383,N_20754,N_20542);
nand U21384 (N_21384,N_20979,N_20643);
nor U21385 (N_21385,N_20631,N_20769);
nand U21386 (N_21386,N_20728,N_20559);
or U21387 (N_21387,N_20931,N_20978);
nand U21388 (N_21388,N_20658,N_20995);
xnor U21389 (N_21389,N_20755,N_20806);
xor U21390 (N_21390,N_20868,N_20974);
nand U21391 (N_21391,N_20780,N_20626);
and U21392 (N_21392,N_20896,N_20830);
xor U21393 (N_21393,N_20908,N_20929);
and U21394 (N_21394,N_20741,N_20886);
or U21395 (N_21395,N_20879,N_20535);
xnor U21396 (N_21396,N_20828,N_20660);
or U21397 (N_21397,N_20689,N_20673);
or U21398 (N_21398,N_20985,N_20852);
or U21399 (N_21399,N_20857,N_20682);
xnor U21400 (N_21400,N_20802,N_20617);
and U21401 (N_21401,N_20905,N_20850);
or U21402 (N_21402,N_20599,N_20829);
or U21403 (N_21403,N_20854,N_20638);
and U21404 (N_21404,N_20652,N_20971);
or U21405 (N_21405,N_20759,N_20628);
xnor U21406 (N_21406,N_20601,N_20857);
nor U21407 (N_21407,N_20559,N_20800);
or U21408 (N_21408,N_20539,N_20606);
xor U21409 (N_21409,N_20850,N_20640);
and U21410 (N_21410,N_20666,N_20607);
nand U21411 (N_21411,N_20533,N_20583);
xnor U21412 (N_21412,N_20993,N_20941);
nand U21413 (N_21413,N_20517,N_20777);
xnor U21414 (N_21414,N_20540,N_20938);
nand U21415 (N_21415,N_20540,N_20929);
xor U21416 (N_21416,N_20541,N_20831);
xnor U21417 (N_21417,N_20923,N_20823);
or U21418 (N_21418,N_20661,N_20548);
nor U21419 (N_21419,N_20850,N_20552);
xnor U21420 (N_21420,N_20620,N_20747);
nand U21421 (N_21421,N_20671,N_20939);
xor U21422 (N_21422,N_20747,N_20536);
and U21423 (N_21423,N_20741,N_20598);
nor U21424 (N_21424,N_20557,N_20992);
or U21425 (N_21425,N_20761,N_20620);
nor U21426 (N_21426,N_20945,N_20722);
nor U21427 (N_21427,N_20714,N_20938);
nor U21428 (N_21428,N_20661,N_20659);
and U21429 (N_21429,N_20763,N_20830);
and U21430 (N_21430,N_20813,N_20958);
and U21431 (N_21431,N_20724,N_20996);
xnor U21432 (N_21432,N_20550,N_20504);
xor U21433 (N_21433,N_20852,N_20805);
and U21434 (N_21434,N_20661,N_20766);
xnor U21435 (N_21435,N_20831,N_20503);
and U21436 (N_21436,N_20671,N_20500);
xor U21437 (N_21437,N_20906,N_20642);
nor U21438 (N_21438,N_20841,N_20736);
nand U21439 (N_21439,N_20517,N_20671);
xor U21440 (N_21440,N_20575,N_20756);
nor U21441 (N_21441,N_20669,N_20594);
xnor U21442 (N_21442,N_20652,N_20998);
nor U21443 (N_21443,N_20589,N_20844);
or U21444 (N_21444,N_20793,N_20915);
nand U21445 (N_21445,N_20751,N_20966);
xor U21446 (N_21446,N_20603,N_20859);
xor U21447 (N_21447,N_20545,N_20610);
nand U21448 (N_21448,N_20696,N_20582);
xor U21449 (N_21449,N_20546,N_20849);
xnor U21450 (N_21450,N_20569,N_20557);
and U21451 (N_21451,N_20536,N_20728);
and U21452 (N_21452,N_20656,N_20673);
nor U21453 (N_21453,N_20517,N_20592);
nor U21454 (N_21454,N_20736,N_20958);
xor U21455 (N_21455,N_20500,N_20925);
nand U21456 (N_21456,N_20815,N_20747);
xnor U21457 (N_21457,N_20946,N_20860);
and U21458 (N_21458,N_20721,N_20554);
and U21459 (N_21459,N_20981,N_20532);
nand U21460 (N_21460,N_20953,N_20869);
nand U21461 (N_21461,N_20500,N_20585);
and U21462 (N_21462,N_20628,N_20547);
nand U21463 (N_21463,N_20925,N_20562);
nor U21464 (N_21464,N_20536,N_20953);
xnor U21465 (N_21465,N_20626,N_20675);
nand U21466 (N_21466,N_20677,N_20570);
and U21467 (N_21467,N_20777,N_20520);
and U21468 (N_21468,N_20679,N_20587);
nor U21469 (N_21469,N_20619,N_20839);
or U21470 (N_21470,N_20594,N_20967);
and U21471 (N_21471,N_20942,N_20707);
xor U21472 (N_21472,N_20684,N_20519);
or U21473 (N_21473,N_20927,N_20511);
nor U21474 (N_21474,N_20764,N_20760);
xnor U21475 (N_21475,N_20943,N_20893);
nand U21476 (N_21476,N_20504,N_20668);
nand U21477 (N_21477,N_20927,N_20639);
nand U21478 (N_21478,N_20769,N_20749);
nor U21479 (N_21479,N_20740,N_20979);
and U21480 (N_21480,N_20955,N_20933);
nor U21481 (N_21481,N_20692,N_20801);
nor U21482 (N_21482,N_20605,N_20522);
nor U21483 (N_21483,N_20963,N_20581);
nor U21484 (N_21484,N_20983,N_20985);
nand U21485 (N_21485,N_20829,N_20631);
or U21486 (N_21486,N_20572,N_20512);
or U21487 (N_21487,N_20600,N_20592);
and U21488 (N_21488,N_20951,N_20605);
nand U21489 (N_21489,N_20611,N_20519);
or U21490 (N_21490,N_20771,N_20900);
or U21491 (N_21491,N_20792,N_20568);
nor U21492 (N_21492,N_20695,N_20780);
xor U21493 (N_21493,N_20783,N_20656);
and U21494 (N_21494,N_20782,N_20928);
nand U21495 (N_21495,N_20992,N_20678);
nor U21496 (N_21496,N_20534,N_20628);
nand U21497 (N_21497,N_20997,N_20872);
or U21498 (N_21498,N_20852,N_20681);
or U21499 (N_21499,N_20902,N_20516);
and U21500 (N_21500,N_21472,N_21384);
nand U21501 (N_21501,N_21376,N_21297);
xor U21502 (N_21502,N_21150,N_21071);
or U21503 (N_21503,N_21331,N_21054);
and U21504 (N_21504,N_21091,N_21353);
nor U21505 (N_21505,N_21455,N_21327);
or U21506 (N_21506,N_21029,N_21214);
nand U21507 (N_21507,N_21474,N_21027);
nor U21508 (N_21508,N_21227,N_21436);
nor U21509 (N_21509,N_21460,N_21388);
and U21510 (N_21510,N_21125,N_21269);
or U21511 (N_21511,N_21032,N_21058);
and U21512 (N_21512,N_21082,N_21239);
nor U21513 (N_21513,N_21184,N_21172);
xor U21514 (N_21514,N_21129,N_21347);
or U21515 (N_21515,N_21086,N_21392);
or U21516 (N_21516,N_21034,N_21256);
and U21517 (N_21517,N_21352,N_21015);
xnor U21518 (N_21518,N_21064,N_21275);
or U21519 (N_21519,N_21025,N_21461);
and U21520 (N_21520,N_21076,N_21263);
or U21521 (N_21521,N_21037,N_21469);
nor U21522 (N_21522,N_21398,N_21238);
xor U21523 (N_21523,N_21145,N_21024);
xor U21524 (N_21524,N_21278,N_21133);
xor U21525 (N_21525,N_21268,N_21247);
nand U21526 (N_21526,N_21201,N_21063);
nor U21527 (N_21527,N_21118,N_21336);
nor U21528 (N_21528,N_21020,N_21323);
and U21529 (N_21529,N_21276,N_21042);
nand U21530 (N_21530,N_21023,N_21121);
or U21531 (N_21531,N_21369,N_21223);
or U21532 (N_21532,N_21229,N_21138);
nand U21533 (N_21533,N_21390,N_21218);
or U21534 (N_21534,N_21070,N_21136);
or U21535 (N_21535,N_21094,N_21226);
nand U21536 (N_21536,N_21394,N_21132);
and U21537 (N_21537,N_21333,N_21093);
and U21538 (N_21538,N_21252,N_21154);
or U21539 (N_21539,N_21308,N_21135);
and U21540 (N_21540,N_21065,N_21210);
or U21541 (N_21541,N_21350,N_21111);
xnor U21542 (N_21542,N_21199,N_21096);
xor U21543 (N_21543,N_21232,N_21446);
nor U21544 (N_21544,N_21311,N_21113);
xor U21545 (N_21545,N_21485,N_21495);
and U21546 (N_21546,N_21442,N_21028);
xor U21547 (N_21547,N_21470,N_21321);
or U21548 (N_21548,N_21147,N_21072);
nand U21549 (N_21549,N_21157,N_21477);
and U21550 (N_21550,N_21481,N_21457);
or U21551 (N_21551,N_21441,N_21193);
and U21552 (N_21552,N_21494,N_21045);
nor U21553 (N_21553,N_21168,N_21440);
or U21554 (N_21554,N_21013,N_21270);
nor U21555 (N_21555,N_21379,N_21224);
xnor U21556 (N_21556,N_21438,N_21162);
and U21557 (N_21557,N_21406,N_21416);
nor U21558 (N_21558,N_21351,N_21274);
nand U21559 (N_21559,N_21397,N_21453);
xnor U21560 (N_21560,N_21487,N_21359);
or U21561 (N_21561,N_21001,N_21435);
and U21562 (N_21562,N_21332,N_21185);
and U21563 (N_21563,N_21366,N_21383);
or U21564 (N_21564,N_21476,N_21281);
nand U21565 (N_21565,N_21097,N_21213);
nand U21566 (N_21566,N_21099,N_21326);
or U21567 (N_21567,N_21445,N_21217);
and U21568 (N_21568,N_21468,N_21279);
and U21569 (N_21569,N_21000,N_21221);
and U21570 (N_21570,N_21466,N_21048);
xor U21571 (N_21571,N_21095,N_21044);
or U21572 (N_21572,N_21148,N_21035);
nand U21573 (N_21573,N_21374,N_21335);
nand U21574 (N_21574,N_21262,N_21200);
nand U21575 (N_21575,N_21038,N_21292);
nor U21576 (N_21576,N_21191,N_21273);
nor U21577 (N_21577,N_21315,N_21041);
xor U21578 (N_21578,N_21115,N_21235);
and U21579 (N_21579,N_21219,N_21016);
nor U21580 (N_21580,N_21426,N_21146);
or U21581 (N_21581,N_21299,N_21073);
or U21582 (N_21582,N_21380,N_21152);
and U21583 (N_21583,N_21117,N_21074);
and U21584 (N_21584,N_21459,N_21451);
and U21585 (N_21585,N_21040,N_21225);
xnor U21586 (N_21586,N_21230,N_21030);
nand U21587 (N_21587,N_21008,N_21497);
nor U21588 (N_21588,N_21414,N_21370);
or U21589 (N_21589,N_21019,N_21300);
or U21590 (N_21590,N_21362,N_21081);
and U21591 (N_21591,N_21202,N_21182);
nand U21592 (N_21592,N_21309,N_21189);
nand U21593 (N_21593,N_21410,N_21429);
and U21594 (N_21594,N_21005,N_21106);
or U21595 (N_21595,N_21478,N_21314);
xor U21596 (N_21596,N_21052,N_21491);
xor U21597 (N_21597,N_21346,N_21365);
xnor U21598 (N_21598,N_21204,N_21062);
and U21599 (N_21599,N_21198,N_21180);
nor U21600 (N_21600,N_21284,N_21395);
or U21601 (N_21601,N_21004,N_21192);
nand U21602 (N_21602,N_21434,N_21285);
and U21603 (N_21603,N_21294,N_21128);
nor U21604 (N_21604,N_21183,N_21264);
and U21605 (N_21605,N_21250,N_21055);
nor U21606 (N_21606,N_21006,N_21194);
nand U21607 (N_21607,N_21405,N_21156);
nand U21608 (N_21608,N_21293,N_21197);
or U21609 (N_21609,N_21389,N_21069);
nor U21610 (N_21610,N_21159,N_21059);
and U21611 (N_21611,N_21344,N_21216);
nor U21612 (N_21612,N_21266,N_21039);
xor U21613 (N_21613,N_21211,N_21240);
nand U21614 (N_21614,N_21473,N_21153);
nor U21615 (N_21615,N_21448,N_21258);
xnor U21616 (N_21616,N_21155,N_21367);
xor U21617 (N_21617,N_21399,N_21131);
or U21618 (N_21618,N_21303,N_21482);
and U21619 (N_21619,N_21080,N_21017);
and U21620 (N_21620,N_21393,N_21100);
xnor U21621 (N_21621,N_21291,N_21430);
or U21622 (N_21622,N_21026,N_21375);
and U21623 (N_21623,N_21396,N_21205);
or U21624 (N_21624,N_21431,N_21361);
nor U21625 (N_21625,N_21167,N_21415);
nor U21626 (N_21626,N_21400,N_21496);
nand U21627 (N_21627,N_21464,N_21174);
nand U21628 (N_21628,N_21207,N_21498);
nor U21629 (N_21629,N_21186,N_21358);
nand U21630 (N_21630,N_21348,N_21134);
nor U21631 (N_21631,N_21089,N_21165);
or U21632 (N_21632,N_21137,N_21046);
and U21633 (N_21633,N_21319,N_21068);
or U21634 (N_21634,N_21112,N_21212);
or U21635 (N_21635,N_21088,N_21283);
nand U21636 (N_21636,N_21480,N_21043);
nand U21637 (N_21637,N_21463,N_21007);
nor U21638 (N_21638,N_21003,N_21298);
xnor U21639 (N_21639,N_21231,N_21458);
or U21640 (N_21640,N_21011,N_21077);
and U21641 (N_21641,N_21424,N_21439);
and U21642 (N_21642,N_21098,N_21161);
xnor U21643 (N_21643,N_21103,N_21364);
and U21644 (N_21644,N_21176,N_21404);
nor U21645 (N_21645,N_21413,N_21411);
or U21646 (N_21646,N_21060,N_21363);
and U21647 (N_21647,N_21475,N_21310);
or U21648 (N_21648,N_21142,N_21158);
or U21649 (N_21649,N_21143,N_21493);
and U21650 (N_21650,N_21306,N_21325);
xor U21651 (N_21651,N_21206,N_21181);
or U21652 (N_21652,N_21305,N_21010);
nand U21653 (N_21653,N_21289,N_21151);
and U21654 (N_21654,N_21109,N_21377);
and U21655 (N_21655,N_21382,N_21343);
nor U21656 (N_21656,N_21368,N_21130);
nand U21657 (N_21657,N_21149,N_21160);
nor U21658 (N_21658,N_21021,N_21251);
or U21659 (N_21659,N_21433,N_21342);
xnor U21660 (N_21660,N_21124,N_21237);
xor U21661 (N_21661,N_21102,N_21360);
or U21662 (N_21662,N_21108,N_21313);
and U21663 (N_21663,N_21277,N_21012);
nor U21664 (N_21664,N_21177,N_21421);
nand U21665 (N_21665,N_21107,N_21418);
or U21666 (N_21666,N_21033,N_21338);
or U21667 (N_21667,N_21356,N_21340);
or U21668 (N_21668,N_21244,N_21403);
and U21669 (N_21669,N_21241,N_21328);
or U21670 (N_21670,N_21373,N_21220);
nor U21671 (N_21671,N_21419,N_21320);
nor U21672 (N_21672,N_21170,N_21190);
xor U21673 (N_21673,N_21428,N_21049);
xnor U21674 (N_21674,N_21272,N_21246);
nand U21675 (N_21675,N_21391,N_21349);
xor U21676 (N_21676,N_21345,N_21144);
and U21677 (N_21677,N_21215,N_21022);
nor U21678 (N_21678,N_21339,N_21423);
or U21679 (N_21679,N_21208,N_21127);
nand U21680 (N_21680,N_21228,N_21322);
nor U21681 (N_21681,N_21222,N_21452);
and U21682 (N_21682,N_21465,N_21499);
and U21683 (N_21683,N_21265,N_21486);
or U21684 (N_21684,N_21260,N_21178);
and U21685 (N_21685,N_21280,N_21420);
nor U21686 (N_21686,N_21188,N_21409);
xnor U21687 (N_21687,N_21408,N_21267);
nor U21688 (N_21688,N_21120,N_21286);
xor U21689 (N_21689,N_21454,N_21209);
xor U21690 (N_21690,N_21372,N_21075);
nand U21691 (N_21691,N_21341,N_21123);
nor U21692 (N_21692,N_21317,N_21047);
or U21693 (N_21693,N_21355,N_21371);
or U21694 (N_21694,N_21248,N_21479);
xnor U21695 (N_21695,N_21381,N_21490);
and U21696 (N_21696,N_21101,N_21387);
or U21697 (N_21697,N_21053,N_21078);
or U21698 (N_21698,N_21014,N_21432);
or U21699 (N_21699,N_21259,N_21304);
nand U21700 (N_21700,N_21085,N_21324);
nor U21701 (N_21701,N_21056,N_21116);
nor U21702 (N_21702,N_21233,N_21295);
nor U21703 (N_21703,N_21083,N_21234);
xnor U21704 (N_21704,N_21057,N_21119);
and U21705 (N_21705,N_21316,N_21171);
and U21706 (N_21706,N_21422,N_21122);
nand U21707 (N_21707,N_21031,N_21492);
nor U21708 (N_21708,N_21447,N_21412);
xnor U21709 (N_21709,N_21079,N_21456);
nor U21710 (N_21710,N_21386,N_21253);
nor U21711 (N_21711,N_21141,N_21483);
or U21712 (N_21712,N_21066,N_21163);
or U21713 (N_21713,N_21126,N_21402);
nor U21714 (N_21714,N_21307,N_21245);
nand U21715 (N_21715,N_21484,N_21301);
or U21716 (N_21716,N_21449,N_21257);
or U21717 (N_21717,N_21051,N_21318);
or U21718 (N_21718,N_21087,N_21092);
and U21719 (N_21719,N_21255,N_21407);
and U21720 (N_21720,N_21288,N_21337);
nor U21721 (N_21721,N_21471,N_21282);
and U21722 (N_21722,N_21385,N_21243);
xnor U21723 (N_21723,N_21140,N_21090);
nand U21724 (N_21724,N_21290,N_21249);
or U21725 (N_21725,N_21067,N_21203);
nand U21726 (N_21726,N_21061,N_21462);
nand U21727 (N_21727,N_21009,N_21236);
and U21728 (N_21728,N_21254,N_21179);
and U21729 (N_21729,N_21139,N_21488);
nand U21730 (N_21730,N_21357,N_21302);
or U21731 (N_21731,N_21105,N_21271);
and U21732 (N_21732,N_21401,N_21467);
and U21733 (N_21733,N_21169,N_21334);
or U21734 (N_21734,N_21450,N_21444);
nand U21735 (N_21735,N_21175,N_21018);
xor U21736 (N_21736,N_21443,N_21166);
nor U21737 (N_21737,N_21417,N_21002);
or U21738 (N_21738,N_21261,N_21287);
xor U21739 (N_21739,N_21354,N_21427);
or U21740 (N_21740,N_21084,N_21110);
nor U21741 (N_21741,N_21164,N_21187);
nor U21742 (N_21742,N_21329,N_21425);
nand U21743 (N_21743,N_21173,N_21114);
or U21744 (N_21744,N_21296,N_21312);
or U21745 (N_21745,N_21036,N_21196);
and U21746 (N_21746,N_21437,N_21242);
xor U21747 (N_21747,N_21050,N_21195);
nand U21748 (N_21748,N_21104,N_21330);
and U21749 (N_21749,N_21489,N_21378);
nand U21750 (N_21750,N_21158,N_21183);
nand U21751 (N_21751,N_21398,N_21189);
or U21752 (N_21752,N_21486,N_21423);
nor U21753 (N_21753,N_21430,N_21362);
and U21754 (N_21754,N_21241,N_21221);
xor U21755 (N_21755,N_21296,N_21309);
or U21756 (N_21756,N_21485,N_21077);
nand U21757 (N_21757,N_21206,N_21019);
nor U21758 (N_21758,N_21279,N_21165);
nand U21759 (N_21759,N_21057,N_21094);
or U21760 (N_21760,N_21057,N_21101);
or U21761 (N_21761,N_21224,N_21364);
or U21762 (N_21762,N_21056,N_21335);
nand U21763 (N_21763,N_21450,N_21132);
and U21764 (N_21764,N_21349,N_21312);
nand U21765 (N_21765,N_21489,N_21160);
xor U21766 (N_21766,N_21454,N_21345);
and U21767 (N_21767,N_21345,N_21434);
xnor U21768 (N_21768,N_21162,N_21279);
nor U21769 (N_21769,N_21164,N_21434);
nor U21770 (N_21770,N_21125,N_21105);
xor U21771 (N_21771,N_21287,N_21202);
nor U21772 (N_21772,N_21236,N_21233);
or U21773 (N_21773,N_21096,N_21001);
and U21774 (N_21774,N_21034,N_21368);
nand U21775 (N_21775,N_21050,N_21266);
xnor U21776 (N_21776,N_21486,N_21080);
nand U21777 (N_21777,N_21249,N_21114);
nand U21778 (N_21778,N_21095,N_21388);
xnor U21779 (N_21779,N_21329,N_21114);
xor U21780 (N_21780,N_21448,N_21184);
and U21781 (N_21781,N_21369,N_21287);
nand U21782 (N_21782,N_21090,N_21023);
and U21783 (N_21783,N_21334,N_21331);
xnor U21784 (N_21784,N_21435,N_21467);
xor U21785 (N_21785,N_21472,N_21346);
nand U21786 (N_21786,N_21073,N_21254);
or U21787 (N_21787,N_21235,N_21200);
nand U21788 (N_21788,N_21444,N_21166);
or U21789 (N_21789,N_21378,N_21231);
nand U21790 (N_21790,N_21179,N_21076);
or U21791 (N_21791,N_21450,N_21324);
nor U21792 (N_21792,N_21099,N_21429);
nand U21793 (N_21793,N_21496,N_21480);
or U21794 (N_21794,N_21162,N_21499);
nor U21795 (N_21795,N_21274,N_21146);
or U21796 (N_21796,N_21227,N_21025);
or U21797 (N_21797,N_21424,N_21025);
and U21798 (N_21798,N_21448,N_21408);
nand U21799 (N_21799,N_21050,N_21357);
nor U21800 (N_21800,N_21298,N_21060);
and U21801 (N_21801,N_21211,N_21051);
nand U21802 (N_21802,N_21358,N_21245);
nor U21803 (N_21803,N_21125,N_21119);
nand U21804 (N_21804,N_21012,N_21323);
or U21805 (N_21805,N_21347,N_21459);
nand U21806 (N_21806,N_21147,N_21276);
nand U21807 (N_21807,N_21325,N_21224);
or U21808 (N_21808,N_21499,N_21295);
nor U21809 (N_21809,N_21231,N_21408);
nor U21810 (N_21810,N_21309,N_21456);
nand U21811 (N_21811,N_21297,N_21069);
nand U21812 (N_21812,N_21447,N_21206);
and U21813 (N_21813,N_21097,N_21449);
and U21814 (N_21814,N_21251,N_21477);
nor U21815 (N_21815,N_21096,N_21131);
or U21816 (N_21816,N_21362,N_21441);
xor U21817 (N_21817,N_21169,N_21104);
xor U21818 (N_21818,N_21405,N_21491);
or U21819 (N_21819,N_21169,N_21305);
xnor U21820 (N_21820,N_21482,N_21083);
xor U21821 (N_21821,N_21323,N_21044);
and U21822 (N_21822,N_21370,N_21126);
nand U21823 (N_21823,N_21079,N_21029);
nand U21824 (N_21824,N_21475,N_21243);
xnor U21825 (N_21825,N_21450,N_21246);
nand U21826 (N_21826,N_21385,N_21427);
nand U21827 (N_21827,N_21204,N_21213);
xnor U21828 (N_21828,N_21156,N_21372);
and U21829 (N_21829,N_21464,N_21291);
xnor U21830 (N_21830,N_21376,N_21019);
and U21831 (N_21831,N_21335,N_21434);
nor U21832 (N_21832,N_21104,N_21052);
nand U21833 (N_21833,N_21215,N_21287);
and U21834 (N_21834,N_21092,N_21433);
nand U21835 (N_21835,N_21468,N_21426);
nor U21836 (N_21836,N_21043,N_21389);
nor U21837 (N_21837,N_21085,N_21205);
nand U21838 (N_21838,N_21242,N_21355);
and U21839 (N_21839,N_21058,N_21402);
nor U21840 (N_21840,N_21398,N_21165);
or U21841 (N_21841,N_21391,N_21357);
xor U21842 (N_21842,N_21193,N_21387);
or U21843 (N_21843,N_21091,N_21386);
or U21844 (N_21844,N_21202,N_21402);
and U21845 (N_21845,N_21173,N_21232);
nor U21846 (N_21846,N_21467,N_21020);
xnor U21847 (N_21847,N_21379,N_21065);
xor U21848 (N_21848,N_21303,N_21254);
nand U21849 (N_21849,N_21386,N_21247);
nor U21850 (N_21850,N_21396,N_21338);
and U21851 (N_21851,N_21355,N_21099);
xor U21852 (N_21852,N_21271,N_21485);
nand U21853 (N_21853,N_21209,N_21297);
or U21854 (N_21854,N_21283,N_21398);
nor U21855 (N_21855,N_21223,N_21429);
nor U21856 (N_21856,N_21010,N_21061);
or U21857 (N_21857,N_21335,N_21156);
nor U21858 (N_21858,N_21226,N_21033);
nand U21859 (N_21859,N_21461,N_21118);
and U21860 (N_21860,N_21021,N_21171);
xnor U21861 (N_21861,N_21103,N_21007);
or U21862 (N_21862,N_21363,N_21437);
nor U21863 (N_21863,N_21194,N_21036);
xnor U21864 (N_21864,N_21481,N_21409);
xnor U21865 (N_21865,N_21365,N_21034);
or U21866 (N_21866,N_21062,N_21290);
or U21867 (N_21867,N_21010,N_21145);
nand U21868 (N_21868,N_21361,N_21374);
nand U21869 (N_21869,N_21128,N_21183);
nor U21870 (N_21870,N_21208,N_21214);
or U21871 (N_21871,N_21127,N_21298);
nand U21872 (N_21872,N_21189,N_21201);
nor U21873 (N_21873,N_21318,N_21444);
or U21874 (N_21874,N_21156,N_21388);
or U21875 (N_21875,N_21416,N_21274);
xor U21876 (N_21876,N_21415,N_21200);
nand U21877 (N_21877,N_21219,N_21275);
or U21878 (N_21878,N_21236,N_21047);
or U21879 (N_21879,N_21394,N_21129);
nand U21880 (N_21880,N_21129,N_21273);
xor U21881 (N_21881,N_21148,N_21093);
xor U21882 (N_21882,N_21068,N_21151);
xnor U21883 (N_21883,N_21316,N_21134);
xnor U21884 (N_21884,N_21409,N_21045);
and U21885 (N_21885,N_21005,N_21338);
xnor U21886 (N_21886,N_21081,N_21131);
nand U21887 (N_21887,N_21386,N_21269);
nand U21888 (N_21888,N_21144,N_21089);
xnor U21889 (N_21889,N_21011,N_21135);
nand U21890 (N_21890,N_21078,N_21433);
nand U21891 (N_21891,N_21277,N_21278);
nor U21892 (N_21892,N_21210,N_21334);
and U21893 (N_21893,N_21329,N_21028);
xor U21894 (N_21894,N_21415,N_21078);
or U21895 (N_21895,N_21179,N_21222);
or U21896 (N_21896,N_21321,N_21345);
and U21897 (N_21897,N_21457,N_21315);
nand U21898 (N_21898,N_21420,N_21263);
nor U21899 (N_21899,N_21141,N_21009);
xor U21900 (N_21900,N_21369,N_21356);
nand U21901 (N_21901,N_21363,N_21129);
nor U21902 (N_21902,N_21083,N_21378);
xnor U21903 (N_21903,N_21325,N_21387);
nor U21904 (N_21904,N_21196,N_21084);
and U21905 (N_21905,N_21307,N_21323);
and U21906 (N_21906,N_21240,N_21258);
and U21907 (N_21907,N_21273,N_21474);
xnor U21908 (N_21908,N_21151,N_21021);
and U21909 (N_21909,N_21445,N_21470);
and U21910 (N_21910,N_21119,N_21293);
nand U21911 (N_21911,N_21207,N_21126);
nor U21912 (N_21912,N_21087,N_21295);
xnor U21913 (N_21913,N_21321,N_21136);
nor U21914 (N_21914,N_21080,N_21200);
or U21915 (N_21915,N_21296,N_21107);
nand U21916 (N_21916,N_21423,N_21391);
xnor U21917 (N_21917,N_21265,N_21247);
nand U21918 (N_21918,N_21141,N_21374);
and U21919 (N_21919,N_21148,N_21256);
nor U21920 (N_21920,N_21201,N_21007);
and U21921 (N_21921,N_21124,N_21231);
xnor U21922 (N_21922,N_21125,N_21048);
and U21923 (N_21923,N_21263,N_21429);
or U21924 (N_21924,N_21109,N_21310);
or U21925 (N_21925,N_21331,N_21417);
xor U21926 (N_21926,N_21210,N_21155);
xor U21927 (N_21927,N_21297,N_21180);
or U21928 (N_21928,N_21199,N_21141);
nand U21929 (N_21929,N_21403,N_21194);
xor U21930 (N_21930,N_21424,N_21088);
nand U21931 (N_21931,N_21472,N_21014);
or U21932 (N_21932,N_21162,N_21096);
xnor U21933 (N_21933,N_21120,N_21100);
and U21934 (N_21934,N_21476,N_21357);
or U21935 (N_21935,N_21469,N_21391);
xor U21936 (N_21936,N_21420,N_21258);
and U21937 (N_21937,N_21476,N_21449);
nand U21938 (N_21938,N_21140,N_21158);
or U21939 (N_21939,N_21145,N_21127);
and U21940 (N_21940,N_21274,N_21386);
xnor U21941 (N_21941,N_21455,N_21257);
nor U21942 (N_21942,N_21004,N_21297);
or U21943 (N_21943,N_21130,N_21311);
or U21944 (N_21944,N_21197,N_21186);
xor U21945 (N_21945,N_21437,N_21191);
or U21946 (N_21946,N_21366,N_21099);
and U21947 (N_21947,N_21196,N_21427);
or U21948 (N_21948,N_21466,N_21054);
xnor U21949 (N_21949,N_21164,N_21212);
nor U21950 (N_21950,N_21181,N_21007);
or U21951 (N_21951,N_21374,N_21245);
nor U21952 (N_21952,N_21195,N_21081);
nand U21953 (N_21953,N_21238,N_21438);
and U21954 (N_21954,N_21246,N_21421);
nand U21955 (N_21955,N_21211,N_21107);
xnor U21956 (N_21956,N_21344,N_21394);
nand U21957 (N_21957,N_21328,N_21013);
nand U21958 (N_21958,N_21438,N_21111);
nand U21959 (N_21959,N_21390,N_21182);
nor U21960 (N_21960,N_21149,N_21405);
or U21961 (N_21961,N_21271,N_21036);
and U21962 (N_21962,N_21272,N_21178);
xnor U21963 (N_21963,N_21436,N_21119);
and U21964 (N_21964,N_21034,N_21249);
or U21965 (N_21965,N_21491,N_21012);
or U21966 (N_21966,N_21025,N_21195);
and U21967 (N_21967,N_21310,N_21466);
or U21968 (N_21968,N_21338,N_21089);
nand U21969 (N_21969,N_21374,N_21429);
and U21970 (N_21970,N_21056,N_21372);
or U21971 (N_21971,N_21209,N_21139);
or U21972 (N_21972,N_21333,N_21424);
or U21973 (N_21973,N_21231,N_21318);
xor U21974 (N_21974,N_21382,N_21045);
nor U21975 (N_21975,N_21276,N_21260);
or U21976 (N_21976,N_21431,N_21111);
nor U21977 (N_21977,N_21242,N_21170);
or U21978 (N_21978,N_21348,N_21230);
nor U21979 (N_21979,N_21159,N_21119);
xor U21980 (N_21980,N_21398,N_21272);
or U21981 (N_21981,N_21056,N_21289);
xor U21982 (N_21982,N_21080,N_21292);
xnor U21983 (N_21983,N_21079,N_21253);
nand U21984 (N_21984,N_21296,N_21165);
or U21985 (N_21985,N_21022,N_21117);
nand U21986 (N_21986,N_21199,N_21409);
and U21987 (N_21987,N_21008,N_21316);
nand U21988 (N_21988,N_21014,N_21440);
xor U21989 (N_21989,N_21351,N_21273);
and U21990 (N_21990,N_21265,N_21307);
xnor U21991 (N_21991,N_21296,N_21109);
xor U21992 (N_21992,N_21198,N_21478);
or U21993 (N_21993,N_21269,N_21132);
and U21994 (N_21994,N_21408,N_21018);
nor U21995 (N_21995,N_21094,N_21434);
and U21996 (N_21996,N_21158,N_21029);
nor U21997 (N_21997,N_21258,N_21083);
or U21998 (N_21998,N_21413,N_21018);
or U21999 (N_21999,N_21407,N_21061);
or U22000 (N_22000,N_21597,N_21673);
nand U22001 (N_22001,N_21697,N_21713);
or U22002 (N_22002,N_21779,N_21830);
xor U22003 (N_22003,N_21881,N_21503);
or U22004 (N_22004,N_21658,N_21685);
nor U22005 (N_22005,N_21801,N_21898);
and U22006 (N_22006,N_21901,N_21880);
or U22007 (N_22007,N_21680,N_21646);
nand U22008 (N_22008,N_21927,N_21986);
nand U22009 (N_22009,N_21660,N_21719);
xnor U22010 (N_22010,N_21859,N_21698);
nand U22011 (N_22011,N_21607,N_21797);
or U22012 (N_22012,N_21774,N_21521);
nor U22013 (N_22013,N_21670,N_21605);
nor U22014 (N_22014,N_21993,N_21688);
or U22015 (N_22015,N_21835,N_21930);
or U22016 (N_22016,N_21904,N_21924);
or U22017 (N_22017,N_21582,N_21967);
nor U22018 (N_22018,N_21731,N_21662);
nor U22019 (N_22019,N_21960,N_21592);
nand U22020 (N_22020,N_21946,N_21523);
or U22021 (N_22021,N_21739,N_21598);
nor U22022 (N_22022,N_21542,N_21971);
and U22023 (N_22023,N_21763,N_21515);
or U22024 (N_22024,N_21558,N_21847);
and U22025 (N_22025,N_21601,N_21970);
and U22026 (N_22026,N_21926,N_21997);
nor U22027 (N_22027,N_21985,N_21989);
nor U22028 (N_22028,N_21629,N_21596);
or U22029 (N_22029,N_21613,N_21788);
or U22030 (N_22030,N_21691,N_21868);
nor U22031 (N_22031,N_21715,N_21900);
nor U22032 (N_22032,N_21866,N_21925);
xor U22033 (N_22033,N_21699,N_21812);
and U22034 (N_22034,N_21931,N_21943);
nand U22035 (N_22035,N_21841,N_21965);
nand U22036 (N_22036,N_21617,N_21722);
nand U22037 (N_22037,N_21517,N_21548);
nand U22038 (N_22038,N_21909,N_21837);
and U22039 (N_22039,N_21727,N_21700);
xor U22040 (N_22040,N_21689,N_21753);
and U22041 (N_22041,N_21953,N_21831);
and U22042 (N_22042,N_21978,N_21981);
or U22043 (N_22043,N_21832,N_21638);
nor U22044 (N_22044,N_21569,N_21583);
nand U22045 (N_22045,N_21720,N_21649);
nand U22046 (N_22046,N_21518,N_21822);
and U22047 (N_22047,N_21612,N_21661);
and U22048 (N_22048,N_21975,N_21892);
and U22049 (N_22049,N_21908,N_21854);
xnor U22050 (N_22050,N_21765,N_21508);
nor U22051 (N_22051,N_21815,N_21556);
and U22052 (N_22052,N_21844,N_21546);
and U22053 (N_22053,N_21737,N_21532);
or U22054 (N_22054,N_21734,N_21846);
xnor U22055 (N_22055,N_21555,N_21852);
nor U22056 (N_22056,N_21879,N_21684);
and U22057 (N_22057,N_21600,N_21857);
nor U22058 (N_22058,N_21936,N_21510);
and U22059 (N_22059,N_21762,N_21787);
nand U22060 (N_22060,N_21544,N_21608);
xnor U22061 (N_22061,N_21921,N_21690);
nor U22062 (N_22062,N_21827,N_21705);
and U22063 (N_22063,N_21826,N_21703);
nand U22064 (N_22064,N_21587,N_21526);
nand U22065 (N_22065,N_21833,N_21954);
nand U22066 (N_22066,N_21778,N_21724);
nor U22067 (N_22067,N_21780,N_21864);
xor U22068 (N_22068,N_21919,N_21792);
nand U22069 (N_22069,N_21584,N_21655);
or U22070 (N_22070,N_21748,N_21545);
xor U22071 (N_22071,N_21906,N_21987);
nand U22072 (N_22072,N_21956,N_21781);
nor U22073 (N_22073,N_21502,N_21885);
xnor U22074 (N_22074,N_21648,N_21603);
nand U22075 (N_22075,N_21593,N_21917);
nor U22076 (N_22076,N_21741,N_21652);
xnor U22077 (N_22077,N_21524,N_21594);
or U22078 (N_22078,N_21610,N_21541);
xor U22079 (N_22079,N_21902,N_21512);
nor U22080 (N_22080,N_21863,N_21687);
or U22081 (N_22081,N_21893,N_21566);
and U22082 (N_22082,N_21990,N_21630);
nor U22083 (N_22083,N_21775,N_21800);
nor U22084 (N_22084,N_21530,N_21760);
or U22085 (N_22085,N_21851,N_21643);
nand U22086 (N_22086,N_21769,N_21855);
nor U22087 (N_22087,N_21790,N_21692);
or U22088 (N_22088,N_21972,N_21935);
xnor U22089 (N_22089,N_21567,N_21820);
nor U22090 (N_22090,N_21750,N_21573);
xor U22091 (N_22091,N_21883,N_21791);
xor U22092 (N_22092,N_21782,N_21554);
or U22093 (N_22093,N_21614,N_21562);
or U22094 (N_22094,N_21811,N_21907);
nor U22095 (N_22095,N_21942,N_21723);
nand U22096 (N_22096,N_21807,N_21568);
xnor U22097 (N_22097,N_21860,N_21611);
nand U22098 (N_22098,N_21821,N_21983);
nand U22099 (N_22099,N_21585,N_21736);
or U22100 (N_22100,N_21706,N_21520);
nor U22101 (N_22101,N_21913,N_21957);
nand U22102 (N_22102,N_21572,N_21945);
or U22103 (N_22103,N_21561,N_21547);
nor U22104 (N_22104,N_21626,N_21529);
and U22105 (N_22105,N_21798,N_21606);
or U22106 (N_22106,N_21549,N_21633);
nor U22107 (N_22107,N_21962,N_21828);
xor U22108 (N_22108,N_21964,N_21789);
nor U22109 (N_22109,N_21783,N_21726);
and U22110 (N_22110,N_21513,N_21669);
nand U22111 (N_22111,N_21755,N_21533);
nor U22112 (N_22112,N_21838,N_21966);
or U22113 (N_22113,N_21850,N_21730);
or U22114 (N_22114,N_21668,N_21628);
xor U22115 (N_22115,N_21522,N_21514);
xor U22116 (N_22116,N_21525,N_21616);
nor U22117 (N_22117,N_21708,N_21624);
or U22118 (N_22118,N_21580,N_21988);
nor U22119 (N_22119,N_21707,N_21756);
or U22120 (N_22120,N_21777,N_21785);
or U22121 (N_22121,N_21682,N_21874);
nor U22122 (N_22122,N_21559,N_21905);
and U22123 (N_22123,N_21922,N_21923);
xnor U22124 (N_22124,N_21938,N_21933);
or U22125 (N_22125,N_21805,N_21581);
and U22126 (N_22126,N_21876,N_21656);
xnor U22127 (N_22127,N_21560,N_21823);
nor U22128 (N_22128,N_21910,N_21887);
nor U22129 (N_22129,N_21916,N_21886);
xor U22130 (N_22130,N_21976,N_21504);
xor U22131 (N_22131,N_21570,N_21709);
nor U22132 (N_22132,N_21959,N_21712);
and U22133 (N_22133,N_21637,N_21511);
and U22134 (N_22134,N_21528,N_21507);
xnor U22135 (N_22135,N_21675,N_21767);
and U22136 (N_22136,N_21540,N_21784);
or U22137 (N_22137,N_21872,N_21998);
or U22138 (N_22138,N_21856,N_21527);
and U22139 (N_22139,N_21602,N_21799);
and U22140 (N_22140,N_21758,N_21721);
and U22141 (N_22141,N_21576,N_21625);
nand U22142 (N_22142,N_21818,N_21834);
or U22143 (N_22143,N_21615,N_21825);
and U22144 (N_22144,N_21672,N_21751);
xnor U22145 (N_22145,N_21944,N_21579);
xnor U22146 (N_22146,N_21961,N_21819);
nor U22147 (N_22147,N_21686,N_21744);
nand U22148 (N_22148,N_21659,N_21947);
and U22149 (N_22149,N_21589,N_21786);
xor U22150 (N_22150,N_21873,N_21539);
and U22151 (N_22151,N_21796,N_21551);
xnor U22152 (N_22152,N_21870,N_21500);
nor U22153 (N_22153,N_21577,N_21996);
or U22154 (N_22154,N_21557,N_21553);
nand U22155 (N_22155,N_21563,N_21537);
and U22156 (N_22156,N_21969,N_21729);
and U22157 (N_22157,N_21928,N_21757);
or U22158 (N_22158,N_21701,N_21814);
nor U22159 (N_22159,N_21621,N_21861);
nor U22160 (N_22160,N_21694,N_21695);
xnor U22161 (N_22161,N_21754,N_21644);
nand U22162 (N_22162,N_21746,N_21733);
nor U22163 (N_22163,N_21677,N_21620);
xnor U22164 (N_22164,N_21939,N_21586);
or U22165 (N_22165,N_21806,N_21968);
xor U22166 (N_22166,N_21932,N_21915);
or U22167 (N_22167,N_21505,N_21647);
or U22168 (N_22168,N_21952,N_21536);
xor U22169 (N_22169,N_21764,N_21889);
nand U22170 (N_22170,N_21671,N_21631);
xor U22171 (N_22171,N_21808,N_21534);
nand U22172 (N_22172,N_21666,N_21979);
nor U22173 (N_22173,N_21711,N_21848);
nor U22174 (N_22174,N_21725,N_21619);
xnor U22175 (N_22175,N_21949,N_21575);
xor U22176 (N_22176,N_21578,N_21871);
or U22177 (N_22177,N_21552,N_21749);
nor U22178 (N_22178,N_21977,N_21604);
and U22179 (N_22179,N_21982,N_21609);
nand U22180 (N_22180,N_21716,N_21667);
xnor U22181 (N_22181,N_21941,N_21535);
nand U22182 (N_22182,N_21678,N_21664);
nand U22183 (N_22183,N_21911,N_21743);
and U22184 (N_22184,N_21738,N_21999);
or U22185 (N_22185,N_21980,N_21842);
nor U22186 (N_22186,N_21693,N_21795);
nand U22187 (N_22187,N_21803,N_21653);
nor U22188 (N_22188,N_21651,N_21897);
and U22189 (N_22189,N_21802,N_21766);
and U22190 (N_22190,N_21877,N_21895);
or U22191 (N_22191,N_21955,N_21702);
nand U22192 (N_22192,N_21934,N_21650);
nand U22193 (N_22193,N_21696,N_21878);
or U22194 (N_22194,N_21940,N_21618);
and U22195 (N_22195,N_21890,N_21824);
nor U22196 (N_22196,N_21588,N_21858);
and U22197 (N_22197,N_21595,N_21676);
nor U22198 (N_22198,N_21809,N_21564);
xnor U22199 (N_22199,N_21679,N_21645);
nor U22200 (N_22200,N_21742,N_21654);
nand U22201 (N_22201,N_21718,N_21710);
xnor U22202 (N_22202,N_21565,N_21770);
or U22203 (N_22203,N_21963,N_21912);
xnor U22204 (N_22204,N_21973,N_21531);
or U22205 (N_22205,N_21994,N_21732);
nand U22206 (N_22206,N_21867,N_21639);
nand U22207 (N_22207,N_21817,N_21836);
nand U22208 (N_22208,N_21899,N_21903);
nand U22209 (N_22209,N_21914,N_21918);
or U22210 (N_22210,N_21622,N_21761);
and U22211 (N_22211,N_21829,N_21896);
nor U22212 (N_22212,N_21632,N_21634);
xnor U22213 (N_22213,N_21804,N_21853);
and U22214 (N_22214,N_21665,N_21888);
xor U22215 (N_22215,N_21704,N_21640);
nand U22216 (N_22216,N_21538,N_21813);
and U22217 (N_22217,N_21843,N_21891);
nor U22218 (N_22218,N_21862,N_21717);
nand U22219 (N_22219,N_21506,N_21840);
and U22220 (N_22220,N_21635,N_21974);
nand U22221 (N_22221,N_21550,N_21776);
and U22222 (N_22222,N_21958,N_21752);
nand U22223 (N_22223,N_21623,N_21948);
or U22224 (N_22224,N_21992,N_21772);
and U22225 (N_22225,N_21773,N_21516);
and U22226 (N_22226,N_21728,N_21683);
nor U22227 (N_22227,N_21951,N_21875);
or U22228 (N_22228,N_21884,N_21571);
or U22229 (N_22229,N_21663,N_21794);
and U22230 (N_22230,N_21681,N_21995);
nand U22231 (N_22231,N_21501,N_21740);
nand U22232 (N_22232,N_21747,N_21519);
xor U22233 (N_22233,N_21735,N_21590);
nor U22234 (N_22234,N_21845,N_21627);
or U22235 (N_22235,N_21849,N_21950);
and U22236 (N_22236,N_21865,N_21816);
nor U22237 (N_22237,N_21929,N_21810);
nor U22238 (N_22238,N_21636,N_21839);
or U22239 (N_22239,N_21882,N_21937);
and U22240 (N_22240,N_21674,N_21714);
or U22241 (N_22241,N_21768,N_21869);
nor U22242 (N_22242,N_21771,N_21641);
xor U22243 (N_22243,N_21745,N_21759);
or U22244 (N_22244,N_21793,N_21984);
nor U22245 (N_22245,N_21657,N_21642);
and U22246 (N_22246,N_21894,N_21543);
nand U22247 (N_22247,N_21591,N_21574);
nor U22248 (N_22248,N_21920,N_21509);
or U22249 (N_22249,N_21991,N_21599);
xor U22250 (N_22250,N_21535,N_21679);
nor U22251 (N_22251,N_21819,N_21966);
or U22252 (N_22252,N_21522,N_21892);
or U22253 (N_22253,N_21522,N_21871);
or U22254 (N_22254,N_21868,N_21545);
nand U22255 (N_22255,N_21509,N_21563);
nand U22256 (N_22256,N_21892,N_21595);
nand U22257 (N_22257,N_21807,N_21662);
xor U22258 (N_22258,N_21944,N_21699);
or U22259 (N_22259,N_21600,N_21791);
nand U22260 (N_22260,N_21911,N_21736);
or U22261 (N_22261,N_21730,N_21715);
and U22262 (N_22262,N_21523,N_21561);
and U22263 (N_22263,N_21627,N_21772);
or U22264 (N_22264,N_21772,N_21831);
nor U22265 (N_22265,N_21823,N_21802);
or U22266 (N_22266,N_21765,N_21721);
nor U22267 (N_22267,N_21642,N_21678);
nor U22268 (N_22268,N_21836,N_21691);
nor U22269 (N_22269,N_21757,N_21887);
xnor U22270 (N_22270,N_21992,N_21950);
nand U22271 (N_22271,N_21640,N_21826);
nor U22272 (N_22272,N_21910,N_21698);
or U22273 (N_22273,N_21727,N_21857);
nor U22274 (N_22274,N_21545,N_21804);
nor U22275 (N_22275,N_21779,N_21732);
xor U22276 (N_22276,N_21675,N_21831);
and U22277 (N_22277,N_21681,N_21845);
nand U22278 (N_22278,N_21938,N_21533);
nor U22279 (N_22279,N_21722,N_21601);
or U22280 (N_22280,N_21516,N_21735);
or U22281 (N_22281,N_21634,N_21528);
xnor U22282 (N_22282,N_21600,N_21698);
or U22283 (N_22283,N_21534,N_21930);
or U22284 (N_22284,N_21751,N_21704);
or U22285 (N_22285,N_21628,N_21971);
and U22286 (N_22286,N_21903,N_21919);
xnor U22287 (N_22287,N_21831,N_21771);
nor U22288 (N_22288,N_21691,N_21591);
xnor U22289 (N_22289,N_21882,N_21964);
nand U22290 (N_22290,N_21723,N_21989);
or U22291 (N_22291,N_21953,N_21650);
xnor U22292 (N_22292,N_21971,N_21560);
or U22293 (N_22293,N_21557,N_21904);
xor U22294 (N_22294,N_21668,N_21823);
and U22295 (N_22295,N_21756,N_21540);
nand U22296 (N_22296,N_21658,N_21903);
or U22297 (N_22297,N_21911,N_21543);
nor U22298 (N_22298,N_21715,N_21523);
or U22299 (N_22299,N_21992,N_21958);
and U22300 (N_22300,N_21769,N_21878);
nor U22301 (N_22301,N_21973,N_21566);
and U22302 (N_22302,N_21657,N_21952);
nand U22303 (N_22303,N_21863,N_21971);
and U22304 (N_22304,N_21884,N_21511);
and U22305 (N_22305,N_21546,N_21803);
or U22306 (N_22306,N_21623,N_21650);
nor U22307 (N_22307,N_21556,N_21666);
and U22308 (N_22308,N_21524,N_21805);
or U22309 (N_22309,N_21651,N_21988);
and U22310 (N_22310,N_21598,N_21529);
or U22311 (N_22311,N_21539,N_21702);
and U22312 (N_22312,N_21705,N_21653);
xor U22313 (N_22313,N_21573,N_21602);
xor U22314 (N_22314,N_21792,N_21655);
xnor U22315 (N_22315,N_21998,N_21666);
xnor U22316 (N_22316,N_21632,N_21504);
and U22317 (N_22317,N_21542,N_21864);
and U22318 (N_22318,N_21742,N_21741);
xnor U22319 (N_22319,N_21749,N_21940);
nand U22320 (N_22320,N_21754,N_21598);
or U22321 (N_22321,N_21622,N_21888);
and U22322 (N_22322,N_21886,N_21540);
xor U22323 (N_22323,N_21695,N_21678);
xor U22324 (N_22324,N_21968,N_21988);
and U22325 (N_22325,N_21686,N_21561);
and U22326 (N_22326,N_21956,N_21851);
nor U22327 (N_22327,N_21633,N_21670);
nand U22328 (N_22328,N_21984,N_21698);
nand U22329 (N_22329,N_21970,N_21931);
nor U22330 (N_22330,N_21704,N_21969);
xnor U22331 (N_22331,N_21555,N_21902);
xor U22332 (N_22332,N_21527,N_21939);
nor U22333 (N_22333,N_21938,N_21921);
nand U22334 (N_22334,N_21549,N_21514);
nand U22335 (N_22335,N_21977,N_21976);
xnor U22336 (N_22336,N_21841,N_21770);
and U22337 (N_22337,N_21914,N_21662);
and U22338 (N_22338,N_21716,N_21592);
nand U22339 (N_22339,N_21733,N_21646);
nand U22340 (N_22340,N_21774,N_21550);
and U22341 (N_22341,N_21552,N_21828);
nor U22342 (N_22342,N_21545,N_21986);
or U22343 (N_22343,N_21529,N_21769);
and U22344 (N_22344,N_21508,N_21612);
and U22345 (N_22345,N_21554,N_21564);
nand U22346 (N_22346,N_21520,N_21709);
nor U22347 (N_22347,N_21500,N_21896);
nand U22348 (N_22348,N_21564,N_21608);
and U22349 (N_22349,N_21990,N_21913);
nand U22350 (N_22350,N_21814,N_21661);
nor U22351 (N_22351,N_21712,N_21545);
nor U22352 (N_22352,N_21882,N_21668);
nand U22353 (N_22353,N_21520,N_21826);
and U22354 (N_22354,N_21931,N_21984);
xnor U22355 (N_22355,N_21599,N_21817);
or U22356 (N_22356,N_21617,N_21621);
xor U22357 (N_22357,N_21696,N_21824);
xor U22358 (N_22358,N_21801,N_21798);
nor U22359 (N_22359,N_21517,N_21617);
nand U22360 (N_22360,N_21981,N_21789);
and U22361 (N_22361,N_21647,N_21951);
nor U22362 (N_22362,N_21600,N_21972);
and U22363 (N_22363,N_21965,N_21894);
nand U22364 (N_22364,N_21505,N_21965);
nor U22365 (N_22365,N_21760,N_21914);
nor U22366 (N_22366,N_21967,N_21819);
xor U22367 (N_22367,N_21671,N_21657);
nor U22368 (N_22368,N_21686,N_21877);
xor U22369 (N_22369,N_21550,N_21951);
xor U22370 (N_22370,N_21902,N_21972);
xor U22371 (N_22371,N_21975,N_21703);
xnor U22372 (N_22372,N_21644,N_21536);
xnor U22373 (N_22373,N_21514,N_21720);
or U22374 (N_22374,N_21542,N_21694);
nand U22375 (N_22375,N_21793,N_21981);
and U22376 (N_22376,N_21624,N_21536);
and U22377 (N_22377,N_21692,N_21885);
xnor U22378 (N_22378,N_21538,N_21571);
or U22379 (N_22379,N_21548,N_21864);
xor U22380 (N_22380,N_21959,N_21534);
nor U22381 (N_22381,N_21962,N_21787);
and U22382 (N_22382,N_21984,N_21591);
or U22383 (N_22383,N_21518,N_21634);
xor U22384 (N_22384,N_21884,N_21669);
and U22385 (N_22385,N_21656,N_21823);
nor U22386 (N_22386,N_21913,N_21972);
nand U22387 (N_22387,N_21851,N_21612);
and U22388 (N_22388,N_21912,N_21573);
or U22389 (N_22389,N_21862,N_21819);
nor U22390 (N_22390,N_21541,N_21501);
or U22391 (N_22391,N_21503,N_21551);
nor U22392 (N_22392,N_21723,N_21598);
or U22393 (N_22393,N_21936,N_21662);
nor U22394 (N_22394,N_21516,N_21704);
and U22395 (N_22395,N_21523,N_21648);
or U22396 (N_22396,N_21583,N_21912);
nand U22397 (N_22397,N_21962,N_21535);
nor U22398 (N_22398,N_21869,N_21999);
and U22399 (N_22399,N_21883,N_21729);
xnor U22400 (N_22400,N_21715,N_21904);
or U22401 (N_22401,N_21538,N_21753);
xnor U22402 (N_22402,N_21838,N_21689);
or U22403 (N_22403,N_21763,N_21709);
nand U22404 (N_22404,N_21706,N_21701);
xor U22405 (N_22405,N_21803,N_21853);
xnor U22406 (N_22406,N_21966,N_21887);
and U22407 (N_22407,N_21520,N_21639);
nor U22408 (N_22408,N_21966,N_21916);
xor U22409 (N_22409,N_21560,N_21960);
nor U22410 (N_22410,N_21675,N_21883);
and U22411 (N_22411,N_21919,N_21699);
or U22412 (N_22412,N_21989,N_21917);
xnor U22413 (N_22413,N_21768,N_21932);
or U22414 (N_22414,N_21654,N_21993);
xnor U22415 (N_22415,N_21825,N_21512);
xor U22416 (N_22416,N_21815,N_21693);
xor U22417 (N_22417,N_21740,N_21847);
nor U22418 (N_22418,N_21893,N_21654);
xnor U22419 (N_22419,N_21776,N_21912);
nor U22420 (N_22420,N_21727,N_21787);
nand U22421 (N_22421,N_21578,N_21766);
and U22422 (N_22422,N_21541,N_21511);
or U22423 (N_22423,N_21912,N_21702);
and U22424 (N_22424,N_21882,N_21722);
and U22425 (N_22425,N_21824,N_21522);
and U22426 (N_22426,N_21951,N_21833);
xor U22427 (N_22427,N_21767,N_21833);
xnor U22428 (N_22428,N_21878,N_21764);
xnor U22429 (N_22429,N_21622,N_21604);
nor U22430 (N_22430,N_21595,N_21941);
xor U22431 (N_22431,N_21665,N_21549);
and U22432 (N_22432,N_21841,N_21760);
nor U22433 (N_22433,N_21539,N_21940);
nand U22434 (N_22434,N_21875,N_21551);
xnor U22435 (N_22435,N_21922,N_21799);
nor U22436 (N_22436,N_21652,N_21545);
xnor U22437 (N_22437,N_21571,N_21894);
xor U22438 (N_22438,N_21936,N_21742);
and U22439 (N_22439,N_21842,N_21939);
or U22440 (N_22440,N_21523,N_21594);
or U22441 (N_22441,N_21786,N_21511);
xnor U22442 (N_22442,N_21908,N_21544);
xor U22443 (N_22443,N_21538,N_21876);
xor U22444 (N_22444,N_21646,N_21983);
or U22445 (N_22445,N_21650,N_21648);
or U22446 (N_22446,N_21730,N_21888);
xnor U22447 (N_22447,N_21695,N_21784);
and U22448 (N_22448,N_21856,N_21605);
and U22449 (N_22449,N_21732,N_21648);
or U22450 (N_22450,N_21774,N_21845);
and U22451 (N_22451,N_21558,N_21743);
and U22452 (N_22452,N_21627,N_21656);
nand U22453 (N_22453,N_21814,N_21587);
or U22454 (N_22454,N_21809,N_21520);
nor U22455 (N_22455,N_21605,N_21995);
nand U22456 (N_22456,N_21960,N_21721);
nor U22457 (N_22457,N_21546,N_21882);
and U22458 (N_22458,N_21638,N_21887);
nor U22459 (N_22459,N_21575,N_21519);
nor U22460 (N_22460,N_21653,N_21688);
and U22461 (N_22461,N_21926,N_21773);
and U22462 (N_22462,N_21861,N_21608);
and U22463 (N_22463,N_21567,N_21704);
and U22464 (N_22464,N_21686,N_21954);
or U22465 (N_22465,N_21720,N_21749);
or U22466 (N_22466,N_21949,N_21518);
xnor U22467 (N_22467,N_21616,N_21613);
nor U22468 (N_22468,N_21866,N_21771);
nor U22469 (N_22469,N_21818,N_21870);
nand U22470 (N_22470,N_21748,N_21916);
xnor U22471 (N_22471,N_21587,N_21957);
xnor U22472 (N_22472,N_21549,N_21924);
or U22473 (N_22473,N_21923,N_21907);
and U22474 (N_22474,N_21544,N_21789);
xor U22475 (N_22475,N_21531,N_21944);
xor U22476 (N_22476,N_21936,N_21972);
or U22477 (N_22477,N_21518,N_21919);
nor U22478 (N_22478,N_21569,N_21780);
and U22479 (N_22479,N_21835,N_21547);
nor U22480 (N_22480,N_21849,N_21931);
nor U22481 (N_22481,N_21910,N_21748);
nor U22482 (N_22482,N_21946,N_21624);
nand U22483 (N_22483,N_21819,N_21806);
or U22484 (N_22484,N_21729,N_21721);
nor U22485 (N_22485,N_21633,N_21580);
nor U22486 (N_22486,N_21543,N_21690);
xnor U22487 (N_22487,N_21572,N_21874);
nand U22488 (N_22488,N_21875,N_21859);
and U22489 (N_22489,N_21508,N_21504);
xnor U22490 (N_22490,N_21633,N_21822);
xor U22491 (N_22491,N_21630,N_21799);
xor U22492 (N_22492,N_21672,N_21777);
nand U22493 (N_22493,N_21912,N_21681);
nand U22494 (N_22494,N_21596,N_21755);
xnor U22495 (N_22495,N_21814,N_21728);
xnor U22496 (N_22496,N_21732,N_21909);
xnor U22497 (N_22497,N_21625,N_21519);
nor U22498 (N_22498,N_21962,N_21686);
xnor U22499 (N_22499,N_21672,N_21522);
xnor U22500 (N_22500,N_22491,N_22237);
xor U22501 (N_22501,N_22444,N_22140);
and U22502 (N_22502,N_22210,N_22246);
xor U22503 (N_22503,N_22313,N_22471);
nand U22504 (N_22504,N_22350,N_22042);
or U22505 (N_22505,N_22255,N_22121);
nand U22506 (N_22506,N_22302,N_22467);
xnor U22507 (N_22507,N_22122,N_22410);
nor U22508 (N_22508,N_22059,N_22175);
and U22509 (N_22509,N_22331,N_22016);
nand U22510 (N_22510,N_22440,N_22184);
nand U22511 (N_22511,N_22002,N_22182);
and U22512 (N_22512,N_22137,N_22238);
nand U22513 (N_22513,N_22080,N_22063);
xor U22514 (N_22514,N_22213,N_22144);
xnor U22515 (N_22515,N_22096,N_22229);
and U22516 (N_22516,N_22011,N_22161);
nand U22517 (N_22517,N_22085,N_22020);
xor U22518 (N_22518,N_22435,N_22256);
xor U22519 (N_22519,N_22266,N_22226);
or U22520 (N_22520,N_22239,N_22363);
nand U22521 (N_22521,N_22103,N_22318);
and U22522 (N_22522,N_22214,N_22132);
xnor U22523 (N_22523,N_22118,N_22336);
nand U22524 (N_22524,N_22249,N_22048);
xnor U22525 (N_22525,N_22022,N_22480);
and U22526 (N_22526,N_22233,N_22324);
and U22527 (N_22527,N_22101,N_22352);
nor U22528 (N_22528,N_22450,N_22338);
nor U22529 (N_22529,N_22337,N_22291);
xnor U22530 (N_22530,N_22040,N_22117);
or U22531 (N_22531,N_22031,N_22333);
or U22532 (N_22532,N_22236,N_22369);
and U22533 (N_22533,N_22160,N_22299);
nor U22534 (N_22534,N_22403,N_22304);
xnor U22535 (N_22535,N_22455,N_22407);
or U22536 (N_22536,N_22207,N_22286);
and U22537 (N_22537,N_22176,N_22008);
xor U22538 (N_22538,N_22125,N_22279);
nand U22539 (N_22539,N_22376,N_22190);
xnor U22540 (N_22540,N_22128,N_22457);
or U22541 (N_22541,N_22405,N_22078);
nand U22542 (N_22542,N_22469,N_22409);
and U22543 (N_22543,N_22033,N_22007);
nand U22544 (N_22544,N_22472,N_22201);
xnor U22545 (N_22545,N_22342,N_22018);
and U22546 (N_22546,N_22120,N_22251);
xnor U22547 (N_22547,N_22146,N_22025);
xor U22548 (N_22548,N_22221,N_22116);
nand U22549 (N_22549,N_22058,N_22478);
xnor U22550 (N_22550,N_22258,N_22327);
and U22551 (N_22551,N_22298,N_22242);
and U22552 (N_22552,N_22306,N_22164);
xnor U22553 (N_22553,N_22278,N_22465);
nor U22554 (N_22554,N_22408,N_22382);
or U22555 (N_22555,N_22322,N_22325);
and U22556 (N_22556,N_22473,N_22060);
xnor U22557 (N_22557,N_22432,N_22428);
xor U22558 (N_22558,N_22070,N_22170);
or U22559 (N_22559,N_22191,N_22395);
and U22560 (N_22560,N_22202,N_22030);
or U22561 (N_22561,N_22394,N_22415);
and U22562 (N_22562,N_22267,N_22458);
and U22563 (N_22563,N_22314,N_22454);
nor U22564 (N_22564,N_22464,N_22406);
nand U22565 (N_22565,N_22390,N_22490);
nor U22566 (N_22566,N_22339,N_22094);
nor U22567 (N_22567,N_22418,N_22481);
and U22568 (N_22568,N_22487,N_22452);
or U22569 (N_22569,N_22069,N_22218);
xor U22570 (N_22570,N_22013,N_22067);
xor U22571 (N_22571,N_22381,N_22429);
and U22572 (N_22572,N_22173,N_22163);
nor U22573 (N_22573,N_22451,N_22054);
xnor U22574 (N_22574,N_22206,N_22447);
and U22575 (N_22575,N_22316,N_22353);
nand U22576 (N_22576,N_22149,N_22272);
nand U22577 (N_22577,N_22086,N_22220);
xnor U22578 (N_22578,N_22398,N_22466);
nor U22579 (N_22579,N_22035,N_22127);
xnor U22580 (N_22580,N_22050,N_22416);
xor U22581 (N_22581,N_22228,N_22459);
nand U22582 (N_22582,N_22097,N_22276);
nand U22583 (N_22583,N_22106,N_22104);
xnor U22584 (N_22584,N_22355,N_22215);
nand U22585 (N_22585,N_22311,N_22270);
xor U22586 (N_22586,N_22372,N_22178);
xnor U22587 (N_22587,N_22148,N_22212);
nand U22588 (N_22588,N_22391,N_22289);
or U22589 (N_22589,N_22377,N_22165);
nor U22590 (N_22590,N_22371,N_22187);
and U22591 (N_22591,N_22283,N_22043);
and U22592 (N_22592,N_22066,N_22129);
or U22593 (N_22593,N_22168,N_22188);
xnor U22594 (N_22594,N_22496,N_22095);
xor U22595 (N_22595,N_22326,N_22105);
nor U22596 (N_22596,N_22001,N_22098);
xnor U22597 (N_22597,N_22413,N_22345);
or U22598 (N_22598,N_22474,N_22053);
or U22599 (N_22599,N_22365,N_22281);
nor U22600 (N_22600,N_22378,N_22360);
xor U22601 (N_22601,N_22023,N_22072);
nand U22602 (N_22602,N_22028,N_22052);
and U22603 (N_22603,N_22358,N_22319);
nand U22604 (N_22604,N_22074,N_22453);
or U22605 (N_22605,N_22423,N_22292);
nor U22606 (N_22606,N_22064,N_22047);
nand U22607 (N_22607,N_22290,N_22483);
or U22608 (N_22608,N_22077,N_22056);
nor U22609 (N_22609,N_22456,N_22385);
or U22610 (N_22610,N_22169,N_22351);
nor U22611 (N_22611,N_22075,N_22208);
and U22612 (N_22612,N_22262,N_22424);
nor U22613 (N_22613,N_22192,N_22356);
nor U22614 (N_22614,N_22426,N_22373);
nor U22615 (N_22615,N_22115,N_22235);
nand U22616 (N_22616,N_22183,N_22384);
nand U22617 (N_22617,N_22330,N_22359);
nor U22618 (N_22618,N_22089,N_22216);
or U22619 (N_22619,N_22126,N_22323);
and U22620 (N_22620,N_22261,N_22166);
xnor U22621 (N_22621,N_22332,N_22019);
and U22622 (N_22622,N_22108,N_22422);
nor U22623 (N_22623,N_22032,N_22366);
or U22624 (N_22624,N_22257,N_22172);
or U22625 (N_22625,N_22123,N_22189);
xor U22626 (N_22626,N_22181,N_22341);
xnor U22627 (N_22627,N_22203,N_22073);
and U22628 (N_22628,N_22107,N_22375);
nor U22629 (N_22629,N_22484,N_22434);
and U22630 (N_22630,N_22263,N_22162);
nand U22631 (N_22631,N_22209,N_22492);
nand U22632 (N_22632,N_22329,N_22026);
and U22633 (N_22633,N_22293,N_22417);
or U22634 (N_22634,N_22370,N_22393);
and U22635 (N_22635,N_22227,N_22388);
nor U22636 (N_22636,N_22100,N_22017);
xor U22637 (N_22637,N_22138,N_22294);
nor U22638 (N_22638,N_22486,N_22046);
xnor U22639 (N_22639,N_22079,N_22461);
nor U22640 (N_22640,N_22158,N_22240);
xor U22641 (N_22641,N_22380,N_22437);
and U22642 (N_22642,N_22133,N_22335);
and U22643 (N_22643,N_22055,N_22036);
nor U22644 (N_22644,N_22065,N_22130);
or U22645 (N_22645,N_22387,N_22143);
xor U22646 (N_22646,N_22156,N_22194);
xnor U22647 (N_22647,N_22248,N_22153);
xor U22648 (N_22648,N_22280,N_22463);
xnor U22649 (N_22649,N_22124,N_22147);
xor U22650 (N_22650,N_22245,N_22044);
and U22651 (N_22651,N_22199,N_22051);
nor U22652 (N_22652,N_22421,N_22347);
and U22653 (N_22653,N_22092,N_22296);
and U22654 (N_22654,N_22307,N_22139);
or U22655 (N_22655,N_22441,N_22038);
nand U22656 (N_22656,N_22468,N_22389);
or U22657 (N_22657,N_22346,N_22400);
or U22658 (N_22658,N_22275,N_22135);
xor U22659 (N_22659,N_22099,N_22195);
and U22660 (N_22660,N_22334,N_22340);
or U22661 (N_22661,N_22386,N_22232);
nor U22662 (N_22662,N_22068,N_22301);
nand U22663 (N_22663,N_22430,N_22110);
nand U22664 (N_22664,N_22009,N_22269);
nand U22665 (N_22665,N_22476,N_22443);
nand U22666 (N_22666,N_22273,N_22475);
xor U22667 (N_22667,N_22489,N_22439);
xor U22668 (N_22668,N_22010,N_22320);
nor U22669 (N_22669,N_22303,N_22284);
xnor U22670 (N_22670,N_22024,N_22446);
nand U22671 (N_22671,N_22401,N_22062);
nand U22672 (N_22672,N_22177,N_22211);
and U22673 (N_22673,N_22493,N_22297);
xor U22674 (N_22674,N_22196,N_22253);
nand U22675 (N_22675,N_22193,N_22374);
xnor U22676 (N_22676,N_22057,N_22436);
xnor U22677 (N_22677,N_22109,N_22392);
xnor U22678 (N_22678,N_22462,N_22477);
xnor U22679 (N_22679,N_22084,N_22343);
and U22680 (N_22680,N_22448,N_22287);
nand U22681 (N_22681,N_22223,N_22159);
and U22682 (N_22682,N_22015,N_22309);
nand U22683 (N_22683,N_22234,N_22041);
and U22684 (N_22684,N_22268,N_22495);
and U22685 (N_22685,N_22250,N_22300);
or U22686 (N_22686,N_22399,N_22145);
or U22687 (N_22687,N_22154,N_22005);
and U22688 (N_22688,N_22167,N_22321);
xnor U22689 (N_22689,N_22397,N_22197);
xor U22690 (N_22690,N_22244,N_22241);
or U22691 (N_22691,N_22282,N_22349);
nor U22692 (N_22692,N_22368,N_22499);
xor U22693 (N_22693,N_22119,N_22076);
or U22694 (N_22694,N_22243,N_22252);
xor U22695 (N_22695,N_22090,N_22083);
nor U22696 (N_22696,N_22419,N_22151);
nor U22697 (N_22697,N_22264,N_22141);
nor U22698 (N_22698,N_22479,N_22488);
nor U22699 (N_22699,N_22029,N_22003);
nand U22700 (N_22700,N_22362,N_22171);
or U22701 (N_22701,N_22111,N_22412);
or U22702 (N_22702,N_22305,N_22112);
or U22703 (N_22703,N_22498,N_22039);
or U22704 (N_22704,N_22222,N_22271);
nor U22705 (N_22705,N_22285,N_22259);
nor U22706 (N_22706,N_22012,N_22460);
and U22707 (N_22707,N_22087,N_22470);
nand U22708 (N_22708,N_22217,N_22354);
nand U22709 (N_22709,N_22186,N_22091);
nand U22710 (N_22710,N_22006,N_22344);
nor U22711 (N_22711,N_22425,N_22225);
nor U22712 (N_22712,N_22420,N_22404);
nor U22713 (N_22713,N_22247,N_22000);
nor U22714 (N_22714,N_22411,N_22482);
nand U22715 (N_22715,N_22082,N_22402);
xnor U22716 (N_22716,N_22204,N_22142);
or U22717 (N_22717,N_22260,N_22383);
nand U22718 (N_22718,N_22157,N_22317);
nor U22719 (N_22719,N_22364,N_22004);
nand U22720 (N_22720,N_22494,N_22180);
xor U22721 (N_22721,N_22071,N_22131);
and U22722 (N_22722,N_22061,N_22308);
xnor U22723 (N_22723,N_22045,N_22136);
nand U22724 (N_22724,N_22328,N_22155);
and U22725 (N_22725,N_22113,N_22088);
nor U22726 (N_22726,N_22205,N_22014);
nor U22727 (N_22727,N_22485,N_22231);
and U22728 (N_22728,N_22134,N_22150);
xor U22729 (N_22729,N_22093,N_22312);
xnor U22730 (N_22730,N_22174,N_22396);
nand U22731 (N_22731,N_22361,N_22152);
nor U22732 (N_22732,N_22021,N_22442);
and U22733 (N_22733,N_22219,N_22367);
nand U22734 (N_22734,N_22295,N_22274);
or U22735 (N_22735,N_22265,N_22224);
and U22736 (N_22736,N_22497,N_22081);
nand U22737 (N_22737,N_22310,N_22049);
xnor U22738 (N_22738,N_22427,N_22414);
nor U22739 (N_22739,N_22198,N_22431);
nor U22740 (N_22740,N_22102,N_22254);
xor U22741 (N_22741,N_22438,N_22449);
nand U22742 (N_22742,N_22037,N_22230);
xor U22743 (N_22743,N_22034,N_22288);
or U22744 (N_22744,N_22185,N_22114);
nand U22745 (N_22745,N_22433,N_22179);
xnor U22746 (N_22746,N_22348,N_22200);
nand U22747 (N_22747,N_22445,N_22277);
nand U22748 (N_22748,N_22027,N_22379);
nand U22749 (N_22749,N_22357,N_22315);
nor U22750 (N_22750,N_22242,N_22135);
xor U22751 (N_22751,N_22129,N_22279);
and U22752 (N_22752,N_22205,N_22357);
nor U22753 (N_22753,N_22462,N_22287);
xnor U22754 (N_22754,N_22322,N_22267);
xor U22755 (N_22755,N_22425,N_22001);
nand U22756 (N_22756,N_22437,N_22215);
or U22757 (N_22757,N_22005,N_22478);
nor U22758 (N_22758,N_22055,N_22370);
and U22759 (N_22759,N_22407,N_22209);
or U22760 (N_22760,N_22345,N_22126);
or U22761 (N_22761,N_22170,N_22136);
and U22762 (N_22762,N_22354,N_22182);
or U22763 (N_22763,N_22454,N_22001);
nor U22764 (N_22764,N_22005,N_22088);
nor U22765 (N_22765,N_22163,N_22422);
nor U22766 (N_22766,N_22240,N_22437);
or U22767 (N_22767,N_22090,N_22192);
xor U22768 (N_22768,N_22374,N_22356);
nand U22769 (N_22769,N_22190,N_22321);
and U22770 (N_22770,N_22254,N_22318);
xnor U22771 (N_22771,N_22449,N_22124);
nor U22772 (N_22772,N_22149,N_22321);
and U22773 (N_22773,N_22065,N_22334);
or U22774 (N_22774,N_22401,N_22128);
nand U22775 (N_22775,N_22145,N_22090);
and U22776 (N_22776,N_22076,N_22413);
nand U22777 (N_22777,N_22316,N_22212);
nand U22778 (N_22778,N_22450,N_22451);
and U22779 (N_22779,N_22206,N_22220);
or U22780 (N_22780,N_22189,N_22269);
xnor U22781 (N_22781,N_22255,N_22182);
xor U22782 (N_22782,N_22202,N_22293);
nand U22783 (N_22783,N_22354,N_22174);
nor U22784 (N_22784,N_22341,N_22361);
nand U22785 (N_22785,N_22087,N_22415);
nand U22786 (N_22786,N_22266,N_22462);
nor U22787 (N_22787,N_22170,N_22418);
nand U22788 (N_22788,N_22193,N_22202);
nand U22789 (N_22789,N_22402,N_22043);
or U22790 (N_22790,N_22119,N_22138);
and U22791 (N_22791,N_22158,N_22043);
xor U22792 (N_22792,N_22084,N_22239);
and U22793 (N_22793,N_22185,N_22108);
nor U22794 (N_22794,N_22118,N_22487);
or U22795 (N_22795,N_22038,N_22020);
xor U22796 (N_22796,N_22261,N_22079);
nand U22797 (N_22797,N_22490,N_22084);
and U22798 (N_22798,N_22017,N_22257);
and U22799 (N_22799,N_22372,N_22336);
nor U22800 (N_22800,N_22178,N_22008);
nand U22801 (N_22801,N_22160,N_22325);
nand U22802 (N_22802,N_22310,N_22332);
nand U22803 (N_22803,N_22043,N_22274);
nor U22804 (N_22804,N_22429,N_22302);
or U22805 (N_22805,N_22178,N_22460);
nor U22806 (N_22806,N_22133,N_22306);
nor U22807 (N_22807,N_22180,N_22114);
and U22808 (N_22808,N_22323,N_22310);
or U22809 (N_22809,N_22208,N_22255);
nor U22810 (N_22810,N_22484,N_22091);
and U22811 (N_22811,N_22008,N_22063);
nor U22812 (N_22812,N_22169,N_22126);
nand U22813 (N_22813,N_22381,N_22069);
and U22814 (N_22814,N_22367,N_22484);
or U22815 (N_22815,N_22117,N_22358);
or U22816 (N_22816,N_22146,N_22331);
xor U22817 (N_22817,N_22272,N_22357);
or U22818 (N_22818,N_22027,N_22206);
nor U22819 (N_22819,N_22262,N_22103);
xor U22820 (N_22820,N_22486,N_22411);
nor U22821 (N_22821,N_22243,N_22281);
xor U22822 (N_22822,N_22186,N_22004);
nand U22823 (N_22823,N_22157,N_22417);
nor U22824 (N_22824,N_22277,N_22324);
and U22825 (N_22825,N_22459,N_22219);
and U22826 (N_22826,N_22275,N_22291);
xor U22827 (N_22827,N_22331,N_22319);
nor U22828 (N_22828,N_22119,N_22299);
or U22829 (N_22829,N_22392,N_22220);
or U22830 (N_22830,N_22422,N_22462);
nor U22831 (N_22831,N_22073,N_22003);
or U22832 (N_22832,N_22081,N_22038);
xnor U22833 (N_22833,N_22172,N_22245);
nand U22834 (N_22834,N_22426,N_22040);
nor U22835 (N_22835,N_22266,N_22293);
or U22836 (N_22836,N_22107,N_22059);
or U22837 (N_22837,N_22441,N_22286);
nor U22838 (N_22838,N_22110,N_22001);
nor U22839 (N_22839,N_22133,N_22024);
and U22840 (N_22840,N_22262,N_22336);
xnor U22841 (N_22841,N_22124,N_22222);
or U22842 (N_22842,N_22086,N_22043);
xor U22843 (N_22843,N_22440,N_22333);
and U22844 (N_22844,N_22499,N_22184);
nor U22845 (N_22845,N_22233,N_22155);
nand U22846 (N_22846,N_22007,N_22401);
and U22847 (N_22847,N_22024,N_22072);
nor U22848 (N_22848,N_22232,N_22289);
nor U22849 (N_22849,N_22168,N_22172);
nor U22850 (N_22850,N_22474,N_22108);
and U22851 (N_22851,N_22413,N_22191);
nor U22852 (N_22852,N_22001,N_22012);
or U22853 (N_22853,N_22033,N_22048);
nor U22854 (N_22854,N_22169,N_22321);
xnor U22855 (N_22855,N_22156,N_22452);
nand U22856 (N_22856,N_22322,N_22185);
xnor U22857 (N_22857,N_22176,N_22060);
xnor U22858 (N_22858,N_22014,N_22240);
xnor U22859 (N_22859,N_22388,N_22204);
xnor U22860 (N_22860,N_22161,N_22207);
nor U22861 (N_22861,N_22476,N_22106);
nand U22862 (N_22862,N_22334,N_22077);
xor U22863 (N_22863,N_22135,N_22353);
nand U22864 (N_22864,N_22262,N_22330);
nor U22865 (N_22865,N_22196,N_22413);
nor U22866 (N_22866,N_22433,N_22094);
or U22867 (N_22867,N_22058,N_22422);
nand U22868 (N_22868,N_22134,N_22137);
or U22869 (N_22869,N_22481,N_22366);
and U22870 (N_22870,N_22443,N_22052);
xnor U22871 (N_22871,N_22080,N_22056);
xnor U22872 (N_22872,N_22054,N_22222);
or U22873 (N_22873,N_22175,N_22298);
nand U22874 (N_22874,N_22092,N_22361);
and U22875 (N_22875,N_22064,N_22129);
xor U22876 (N_22876,N_22325,N_22174);
nor U22877 (N_22877,N_22483,N_22311);
xor U22878 (N_22878,N_22088,N_22219);
and U22879 (N_22879,N_22449,N_22058);
or U22880 (N_22880,N_22003,N_22002);
nand U22881 (N_22881,N_22199,N_22333);
and U22882 (N_22882,N_22071,N_22105);
and U22883 (N_22883,N_22041,N_22206);
xnor U22884 (N_22884,N_22127,N_22449);
nand U22885 (N_22885,N_22138,N_22357);
nand U22886 (N_22886,N_22120,N_22100);
xnor U22887 (N_22887,N_22012,N_22410);
nor U22888 (N_22888,N_22478,N_22182);
or U22889 (N_22889,N_22066,N_22085);
xor U22890 (N_22890,N_22058,N_22221);
or U22891 (N_22891,N_22380,N_22042);
or U22892 (N_22892,N_22419,N_22311);
xnor U22893 (N_22893,N_22296,N_22051);
nor U22894 (N_22894,N_22299,N_22445);
or U22895 (N_22895,N_22488,N_22493);
nand U22896 (N_22896,N_22170,N_22496);
nand U22897 (N_22897,N_22473,N_22179);
xnor U22898 (N_22898,N_22485,N_22048);
or U22899 (N_22899,N_22332,N_22385);
or U22900 (N_22900,N_22099,N_22330);
and U22901 (N_22901,N_22281,N_22479);
or U22902 (N_22902,N_22318,N_22359);
and U22903 (N_22903,N_22498,N_22418);
or U22904 (N_22904,N_22252,N_22080);
nand U22905 (N_22905,N_22278,N_22158);
xor U22906 (N_22906,N_22057,N_22156);
or U22907 (N_22907,N_22360,N_22245);
or U22908 (N_22908,N_22298,N_22121);
and U22909 (N_22909,N_22018,N_22133);
and U22910 (N_22910,N_22065,N_22273);
xor U22911 (N_22911,N_22018,N_22138);
nor U22912 (N_22912,N_22029,N_22109);
xor U22913 (N_22913,N_22032,N_22148);
xor U22914 (N_22914,N_22152,N_22397);
nand U22915 (N_22915,N_22071,N_22487);
nor U22916 (N_22916,N_22122,N_22288);
or U22917 (N_22917,N_22041,N_22157);
xor U22918 (N_22918,N_22226,N_22125);
or U22919 (N_22919,N_22497,N_22290);
xnor U22920 (N_22920,N_22335,N_22437);
xor U22921 (N_22921,N_22374,N_22259);
nand U22922 (N_22922,N_22454,N_22341);
nand U22923 (N_22923,N_22261,N_22433);
xnor U22924 (N_22924,N_22330,N_22317);
and U22925 (N_22925,N_22452,N_22200);
xor U22926 (N_22926,N_22190,N_22346);
and U22927 (N_22927,N_22341,N_22364);
nand U22928 (N_22928,N_22244,N_22221);
nor U22929 (N_22929,N_22202,N_22239);
nand U22930 (N_22930,N_22074,N_22212);
xor U22931 (N_22931,N_22201,N_22231);
or U22932 (N_22932,N_22029,N_22184);
nor U22933 (N_22933,N_22334,N_22037);
xnor U22934 (N_22934,N_22426,N_22277);
xnor U22935 (N_22935,N_22027,N_22357);
and U22936 (N_22936,N_22033,N_22022);
and U22937 (N_22937,N_22059,N_22291);
nor U22938 (N_22938,N_22348,N_22437);
nor U22939 (N_22939,N_22191,N_22187);
xor U22940 (N_22940,N_22475,N_22454);
or U22941 (N_22941,N_22229,N_22058);
or U22942 (N_22942,N_22245,N_22190);
and U22943 (N_22943,N_22106,N_22277);
nor U22944 (N_22944,N_22165,N_22196);
and U22945 (N_22945,N_22486,N_22218);
or U22946 (N_22946,N_22036,N_22015);
nor U22947 (N_22947,N_22348,N_22284);
or U22948 (N_22948,N_22359,N_22339);
xnor U22949 (N_22949,N_22311,N_22444);
xnor U22950 (N_22950,N_22209,N_22342);
or U22951 (N_22951,N_22309,N_22224);
and U22952 (N_22952,N_22189,N_22156);
and U22953 (N_22953,N_22136,N_22154);
or U22954 (N_22954,N_22057,N_22100);
nand U22955 (N_22955,N_22462,N_22066);
and U22956 (N_22956,N_22126,N_22331);
nor U22957 (N_22957,N_22436,N_22107);
or U22958 (N_22958,N_22224,N_22212);
and U22959 (N_22959,N_22330,N_22009);
nand U22960 (N_22960,N_22184,N_22084);
xor U22961 (N_22961,N_22193,N_22496);
and U22962 (N_22962,N_22356,N_22321);
or U22963 (N_22963,N_22287,N_22193);
nand U22964 (N_22964,N_22345,N_22219);
or U22965 (N_22965,N_22496,N_22008);
nor U22966 (N_22966,N_22281,N_22411);
nor U22967 (N_22967,N_22465,N_22378);
and U22968 (N_22968,N_22067,N_22334);
or U22969 (N_22969,N_22049,N_22090);
or U22970 (N_22970,N_22124,N_22215);
nand U22971 (N_22971,N_22182,N_22310);
or U22972 (N_22972,N_22208,N_22448);
and U22973 (N_22973,N_22100,N_22042);
or U22974 (N_22974,N_22208,N_22436);
xor U22975 (N_22975,N_22441,N_22081);
and U22976 (N_22976,N_22374,N_22077);
nor U22977 (N_22977,N_22197,N_22376);
xnor U22978 (N_22978,N_22365,N_22303);
or U22979 (N_22979,N_22182,N_22269);
nand U22980 (N_22980,N_22235,N_22103);
nand U22981 (N_22981,N_22182,N_22240);
or U22982 (N_22982,N_22228,N_22005);
or U22983 (N_22983,N_22055,N_22353);
or U22984 (N_22984,N_22114,N_22497);
or U22985 (N_22985,N_22191,N_22097);
and U22986 (N_22986,N_22135,N_22383);
nand U22987 (N_22987,N_22216,N_22096);
nand U22988 (N_22988,N_22189,N_22209);
xor U22989 (N_22989,N_22147,N_22200);
and U22990 (N_22990,N_22461,N_22106);
and U22991 (N_22991,N_22422,N_22350);
and U22992 (N_22992,N_22238,N_22437);
nand U22993 (N_22993,N_22252,N_22402);
nor U22994 (N_22994,N_22130,N_22448);
nand U22995 (N_22995,N_22216,N_22148);
and U22996 (N_22996,N_22072,N_22236);
nand U22997 (N_22997,N_22264,N_22280);
nand U22998 (N_22998,N_22023,N_22231);
xnor U22999 (N_22999,N_22165,N_22232);
nand U23000 (N_23000,N_22912,N_22997);
nand U23001 (N_23001,N_22546,N_22878);
xnor U23002 (N_23002,N_22974,N_22867);
nor U23003 (N_23003,N_22693,N_22925);
and U23004 (N_23004,N_22580,N_22574);
and U23005 (N_23005,N_22554,N_22705);
xor U23006 (N_23006,N_22835,N_22948);
nand U23007 (N_23007,N_22916,N_22853);
or U23008 (N_23008,N_22504,N_22551);
nor U23009 (N_23009,N_22647,N_22501);
xnor U23010 (N_23010,N_22825,N_22720);
xnor U23011 (N_23011,N_22964,N_22619);
nand U23012 (N_23012,N_22671,N_22783);
xor U23013 (N_23013,N_22814,N_22793);
nor U23014 (N_23014,N_22957,N_22821);
xor U23015 (N_23015,N_22659,N_22928);
nor U23016 (N_23016,N_22588,N_22585);
and U23017 (N_23017,N_22566,N_22518);
and U23018 (N_23018,N_22533,N_22941);
and U23019 (N_23019,N_22852,N_22782);
or U23020 (N_23020,N_22900,N_22700);
nor U23021 (N_23021,N_22876,N_22984);
and U23022 (N_23022,N_22594,N_22718);
xnor U23023 (N_23023,N_22911,N_22988);
xor U23024 (N_23024,N_22775,N_22759);
or U23025 (N_23025,N_22810,N_22990);
xor U23026 (N_23026,N_22528,N_22622);
nand U23027 (N_23027,N_22956,N_22638);
and U23028 (N_23028,N_22550,N_22966);
nand U23029 (N_23029,N_22584,N_22532);
nand U23030 (N_23030,N_22939,N_22895);
and U23031 (N_23031,N_22781,N_22751);
nand U23032 (N_23032,N_22500,N_22543);
and U23033 (N_23033,N_22592,N_22747);
xnor U23034 (N_23034,N_22962,N_22861);
nor U23035 (N_23035,N_22943,N_22901);
and U23036 (N_23036,N_22667,N_22732);
xor U23037 (N_23037,N_22573,N_22885);
and U23038 (N_23038,N_22934,N_22965);
and U23039 (N_23039,N_22762,N_22818);
or U23040 (N_23040,N_22691,N_22576);
or U23041 (N_23041,N_22797,N_22665);
and U23042 (N_23042,N_22578,N_22581);
nand U23043 (N_23043,N_22661,N_22973);
or U23044 (N_23044,N_22505,N_22800);
nand U23045 (N_23045,N_22709,N_22772);
nand U23046 (N_23046,N_22807,N_22830);
or U23047 (N_23047,N_22906,N_22519);
xor U23048 (N_23048,N_22557,N_22664);
nand U23049 (N_23049,N_22841,N_22669);
or U23050 (N_23050,N_22789,N_22947);
and U23051 (N_23051,N_22828,N_22752);
and U23052 (N_23052,N_22648,N_22560);
nor U23053 (N_23053,N_22866,N_22535);
nor U23054 (N_23054,N_22676,N_22612);
or U23055 (N_23055,N_22981,N_22549);
or U23056 (N_23056,N_22844,N_22827);
or U23057 (N_23057,N_22963,N_22597);
nor U23058 (N_23058,N_22982,N_22614);
nor U23059 (N_23059,N_22708,N_22863);
and U23060 (N_23060,N_22564,N_22608);
and U23061 (N_23061,N_22858,N_22544);
nor U23062 (N_23062,N_22923,N_22625);
or U23063 (N_23063,N_22960,N_22513);
nand U23064 (N_23064,N_22673,N_22817);
xnor U23065 (N_23065,N_22552,N_22542);
nor U23066 (N_23066,N_22675,N_22570);
and U23067 (N_23067,N_22530,N_22763);
and U23068 (N_23068,N_22954,N_22712);
or U23069 (N_23069,N_22711,N_22780);
nand U23070 (N_23070,N_22694,N_22833);
or U23071 (N_23071,N_22740,N_22680);
nand U23072 (N_23072,N_22908,N_22804);
nor U23073 (N_23073,N_22650,N_22688);
nor U23074 (N_23074,N_22904,N_22596);
nand U23075 (N_23075,N_22522,N_22998);
or U23076 (N_23076,N_22803,N_22989);
nor U23077 (N_23077,N_22586,N_22644);
and U23078 (N_23078,N_22887,N_22690);
and U23079 (N_23079,N_22764,N_22639);
nor U23080 (N_23080,N_22593,N_22826);
nor U23081 (N_23081,N_22565,N_22508);
and U23082 (N_23082,N_22702,N_22869);
and U23083 (N_23083,N_22822,N_22643);
xnor U23084 (N_23084,N_22641,N_22628);
nor U23085 (N_23085,N_22521,N_22698);
or U23086 (N_23086,N_22598,N_22506);
xnor U23087 (N_23087,N_22791,N_22829);
nand U23088 (N_23088,N_22539,N_22972);
or U23089 (N_23089,N_22657,N_22819);
nor U23090 (N_23090,N_22716,N_22894);
xor U23091 (N_23091,N_22811,N_22813);
or U23092 (N_23092,N_22556,N_22976);
nor U23093 (N_23093,N_22746,N_22798);
or U23094 (N_23094,N_22699,N_22953);
nand U23095 (N_23095,N_22995,N_22651);
nand U23096 (N_23096,N_22996,N_22731);
nand U23097 (N_23097,N_22986,N_22874);
xnor U23098 (N_23098,N_22607,N_22859);
or U23099 (N_23099,N_22662,N_22606);
xnor U23100 (N_23100,N_22864,N_22517);
xnor U23101 (N_23101,N_22575,N_22590);
xor U23102 (N_23102,N_22926,N_22843);
nor U23103 (N_23103,N_22815,N_22725);
and U23104 (N_23104,N_22541,N_22758);
or U23105 (N_23105,N_22971,N_22748);
xnor U23106 (N_23106,N_22631,N_22761);
xor U23107 (N_23107,N_22896,N_22778);
nand U23108 (N_23108,N_22735,N_22886);
or U23109 (N_23109,N_22786,N_22857);
or U23110 (N_23110,N_22950,N_22978);
xnor U23111 (N_23111,N_22790,N_22892);
or U23112 (N_23112,N_22794,N_22801);
or U23113 (N_23113,N_22890,N_22738);
xor U23114 (N_23114,N_22872,N_22701);
xnor U23115 (N_23115,N_22837,N_22579);
nand U23116 (N_23116,N_22572,N_22724);
and U23117 (N_23117,N_22930,N_22524);
nand U23118 (N_23118,N_22511,N_22634);
nor U23119 (N_23119,N_22577,N_22681);
nand U23120 (N_23120,N_22654,N_22558);
or U23121 (N_23121,N_22929,N_22666);
nor U23122 (N_23122,N_22734,N_22591);
and U23123 (N_23123,N_22601,N_22999);
nor U23124 (N_23124,N_22773,N_22697);
nand U23125 (N_23125,N_22921,N_22567);
nor U23126 (N_23126,N_22683,N_22526);
nand U23127 (N_23127,N_22940,N_22985);
nand U23128 (N_23128,N_22931,N_22714);
and U23129 (N_23129,N_22975,N_22561);
and U23130 (N_23130,N_22722,N_22868);
and U23131 (N_23131,N_22674,N_22873);
xnor U23132 (N_23132,N_22820,N_22952);
and U23133 (N_23133,N_22726,N_22704);
nor U23134 (N_23134,N_22706,N_22727);
or U23135 (N_23135,N_22935,N_22686);
or U23136 (N_23136,N_22563,N_22958);
nand U23137 (N_23137,N_22776,N_22509);
xor U23138 (N_23138,N_22766,N_22503);
or U23139 (N_23139,N_22888,N_22587);
nand U23140 (N_23140,N_22792,N_22627);
xor U23141 (N_23141,N_22715,N_22919);
and U23142 (N_23142,N_22512,N_22768);
nor U23143 (N_23143,N_22692,N_22583);
or U23144 (N_23144,N_22562,N_22805);
nor U23145 (N_23145,N_22707,N_22905);
or U23146 (N_23146,N_22653,N_22932);
nand U23147 (N_23147,N_22721,N_22605);
nand U23148 (N_23148,N_22632,N_22992);
or U23149 (N_23149,N_22514,N_22668);
xor U23150 (N_23150,N_22696,N_22754);
or U23151 (N_23151,N_22553,N_22689);
and U23152 (N_23152,N_22969,N_22603);
nand U23153 (N_23153,N_22831,N_22760);
and U23154 (N_23154,N_22617,N_22865);
or U23155 (N_23155,N_22540,N_22796);
xnor U23156 (N_23156,N_22523,N_22944);
or U23157 (N_23157,N_22879,N_22610);
and U23158 (N_23158,N_22942,N_22640);
or U23159 (N_23159,N_22660,N_22949);
and U23160 (N_23160,N_22951,N_22870);
or U23161 (N_23161,N_22795,N_22595);
nor U23162 (N_23162,N_22757,N_22891);
nand U23163 (N_23163,N_22955,N_22623);
nor U23164 (N_23164,N_22626,N_22678);
and U23165 (N_23165,N_22645,N_22710);
or U23166 (N_23166,N_22967,N_22538);
and U23167 (N_23167,N_22679,N_22907);
or U23168 (N_23168,N_22621,N_22624);
nor U23169 (N_23169,N_22730,N_22862);
nand U23170 (N_23170,N_22615,N_22629);
or U23171 (N_23171,N_22860,N_22658);
xor U23172 (N_23172,N_22770,N_22832);
or U23173 (N_23173,N_22914,N_22924);
nand U23174 (N_23174,N_22824,N_22808);
nand U23175 (N_23175,N_22779,N_22893);
nand U23176 (N_23176,N_22785,N_22784);
nand U23177 (N_23177,N_22520,N_22600);
xor U23178 (N_23178,N_22685,N_22806);
xnor U23179 (N_23179,N_22946,N_22655);
and U23180 (N_23180,N_22980,N_22510);
nand U23181 (N_23181,N_22915,N_22717);
nor U23182 (N_23182,N_22589,N_22515);
xor U23183 (N_23183,N_22756,N_22882);
and U23184 (N_23184,N_22719,N_22670);
or U23185 (N_23185,N_22850,N_22910);
and U23186 (N_23186,N_22637,N_22902);
nand U23187 (N_23187,N_22855,N_22527);
and U23188 (N_23188,N_22582,N_22611);
or U23189 (N_23189,N_22548,N_22846);
nand U23190 (N_23190,N_22968,N_22695);
or U23191 (N_23191,N_22994,N_22753);
and U23192 (N_23192,N_22788,N_22672);
xor U23193 (N_23193,N_22507,N_22729);
and U23194 (N_23194,N_22502,N_22677);
or U23195 (N_23195,N_22845,N_22875);
nand U23196 (N_23196,N_22630,N_22884);
or U23197 (N_23197,N_22802,N_22568);
nor U23198 (N_23198,N_22534,N_22613);
or U23199 (N_23199,N_22927,N_22849);
nand U23200 (N_23200,N_22703,N_22903);
xnor U23201 (N_23201,N_22713,N_22663);
nor U23202 (N_23202,N_22842,N_22733);
nor U23203 (N_23203,N_22938,N_22744);
nor U23204 (N_23204,N_22959,N_22602);
xor U23205 (N_23205,N_22774,N_22871);
xnor U23206 (N_23206,N_22616,N_22979);
or U23207 (N_23207,N_22749,N_22609);
xor U23208 (N_23208,N_22991,N_22883);
nand U23209 (N_23209,N_22987,N_22765);
and U23210 (N_23210,N_22977,N_22741);
nor U23211 (N_23211,N_22620,N_22652);
nor U23212 (N_23212,N_22656,N_22769);
or U23213 (N_23213,N_22880,N_22687);
nor U23214 (N_23214,N_22569,N_22646);
xor U23215 (N_23215,N_22684,N_22633);
xnor U23216 (N_23216,N_22516,N_22537);
and U23217 (N_23217,N_22728,N_22599);
or U23218 (N_23218,N_22742,N_22983);
xor U23219 (N_23219,N_22937,N_22636);
and U23220 (N_23220,N_22897,N_22745);
nand U23221 (N_23221,N_22559,N_22851);
xnor U23222 (N_23222,N_22961,N_22816);
or U23223 (N_23223,N_22823,N_22529);
or U23224 (N_23224,N_22854,N_22933);
xor U23225 (N_23225,N_22531,N_22881);
nor U23226 (N_23226,N_22970,N_22918);
xor U23227 (N_23227,N_22877,N_22834);
and U23228 (N_23228,N_22723,N_22856);
or U23229 (N_23229,N_22649,N_22889);
nand U23230 (N_23230,N_22767,N_22922);
nor U23231 (N_23231,N_22555,N_22799);
xnor U23232 (N_23232,N_22840,N_22743);
xor U23233 (N_23233,N_22787,N_22809);
nor U23234 (N_23234,N_22898,N_22736);
nor U23235 (N_23235,N_22777,N_22755);
nand U23236 (N_23236,N_22604,N_22571);
or U23237 (N_23237,N_22737,N_22771);
xor U23238 (N_23238,N_22917,N_22525);
nand U23239 (N_23239,N_22635,N_22545);
and U23240 (N_23240,N_22836,N_22913);
nor U23241 (N_23241,N_22750,N_22812);
or U23242 (N_23242,N_22920,N_22739);
xor U23243 (N_23243,N_22642,N_22682);
nand U23244 (N_23244,N_22899,N_22945);
nor U23245 (N_23245,N_22618,N_22847);
xor U23246 (N_23246,N_22536,N_22839);
nand U23247 (N_23247,N_22909,N_22547);
nor U23248 (N_23248,N_22993,N_22848);
or U23249 (N_23249,N_22838,N_22936);
and U23250 (N_23250,N_22746,N_22968);
and U23251 (N_23251,N_22789,N_22650);
and U23252 (N_23252,N_22540,N_22589);
nand U23253 (N_23253,N_22857,N_22879);
and U23254 (N_23254,N_22856,N_22626);
nand U23255 (N_23255,N_22809,N_22640);
nor U23256 (N_23256,N_22658,N_22871);
and U23257 (N_23257,N_22868,N_22979);
and U23258 (N_23258,N_22852,N_22655);
nor U23259 (N_23259,N_22714,N_22987);
and U23260 (N_23260,N_22557,N_22565);
and U23261 (N_23261,N_22908,N_22712);
or U23262 (N_23262,N_22642,N_22706);
or U23263 (N_23263,N_22612,N_22773);
xor U23264 (N_23264,N_22684,N_22982);
nand U23265 (N_23265,N_22938,N_22694);
or U23266 (N_23266,N_22899,N_22935);
nand U23267 (N_23267,N_22882,N_22834);
and U23268 (N_23268,N_22536,N_22851);
and U23269 (N_23269,N_22951,N_22660);
xnor U23270 (N_23270,N_22552,N_22651);
xnor U23271 (N_23271,N_22659,N_22706);
nor U23272 (N_23272,N_22797,N_22641);
and U23273 (N_23273,N_22853,N_22811);
nand U23274 (N_23274,N_22988,N_22614);
xor U23275 (N_23275,N_22743,N_22597);
or U23276 (N_23276,N_22719,N_22795);
nand U23277 (N_23277,N_22606,N_22524);
or U23278 (N_23278,N_22892,N_22885);
and U23279 (N_23279,N_22971,N_22701);
and U23280 (N_23280,N_22613,N_22847);
or U23281 (N_23281,N_22947,N_22862);
and U23282 (N_23282,N_22984,N_22555);
nand U23283 (N_23283,N_22849,N_22988);
and U23284 (N_23284,N_22846,N_22912);
xor U23285 (N_23285,N_22741,N_22678);
or U23286 (N_23286,N_22728,N_22981);
nand U23287 (N_23287,N_22604,N_22659);
xor U23288 (N_23288,N_22892,N_22565);
nand U23289 (N_23289,N_22551,N_22637);
and U23290 (N_23290,N_22926,N_22697);
and U23291 (N_23291,N_22879,N_22902);
xor U23292 (N_23292,N_22761,N_22805);
and U23293 (N_23293,N_22912,N_22628);
and U23294 (N_23294,N_22987,N_22640);
nand U23295 (N_23295,N_22719,N_22702);
nand U23296 (N_23296,N_22737,N_22964);
xnor U23297 (N_23297,N_22563,N_22686);
nor U23298 (N_23298,N_22831,N_22624);
xor U23299 (N_23299,N_22515,N_22590);
nand U23300 (N_23300,N_22898,N_22520);
nand U23301 (N_23301,N_22551,N_22550);
nor U23302 (N_23302,N_22683,N_22719);
nor U23303 (N_23303,N_22725,N_22688);
xnor U23304 (N_23304,N_22696,N_22641);
xor U23305 (N_23305,N_22927,N_22763);
nor U23306 (N_23306,N_22570,N_22532);
and U23307 (N_23307,N_22854,N_22878);
nor U23308 (N_23308,N_22560,N_22834);
xnor U23309 (N_23309,N_22784,N_22715);
nor U23310 (N_23310,N_22700,N_22949);
or U23311 (N_23311,N_22721,N_22574);
and U23312 (N_23312,N_22814,N_22985);
xor U23313 (N_23313,N_22564,N_22908);
nor U23314 (N_23314,N_22844,N_22842);
nor U23315 (N_23315,N_22648,N_22632);
nand U23316 (N_23316,N_22960,N_22883);
and U23317 (N_23317,N_22718,N_22831);
nand U23318 (N_23318,N_22769,N_22621);
nand U23319 (N_23319,N_22584,N_22845);
or U23320 (N_23320,N_22959,N_22640);
nor U23321 (N_23321,N_22562,N_22837);
nor U23322 (N_23322,N_22520,N_22612);
or U23323 (N_23323,N_22665,N_22910);
nand U23324 (N_23324,N_22752,N_22917);
and U23325 (N_23325,N_22523,N_22797);
nand U23326 (N_23326,N_22748,N_22623);
and U23327 (N_23327,N_22772,N_22597);
or U23328 (N_23328,N_22976,N_22672);
nand U23329 (N_23329,N_22910,N_22730);
xnor U23330 (N_23330,N_22628,N_22632);
and U23331 (N_23331,N_22556,N_22500);
nand U23332 (N_23332,N_22816,N_22722);
and U23333 (N_23333,N_22868,N_22740);
xor U23334 (N_23334,N_22501,N_22709);
and U23335 (N_23335,N_22887,N_22510);
and U23336 (N_23336,N_22756,N_22907);
xnor U23337 (N_23337,N_22923,N_22635);
or U23338 (N_23338,N_22962,N_22898);
xnor U23339 (N_23339,N_22930,N_22731);
or U23340 (N_23340,N_22763,N_22847);
nand U23341 (N_23341,N_22545,N_22786);
nand U23342 (N_23342,N_22782,N_22730);
xnor U23343 (N_23343,N_22577,N_22974);
nor U23344 (N_23344,N_22640,N_22969);
or U23345 (N_23345,N_22786,N_22687);
or U23346 (N_23346,N_22734,N_22679);
and U23347 (N_23347,N_22869,N_22685);
nor U23348 (N_23348,N_22898,N_22881);
or U23349 (N_23349,N_22881,N_22518);
or U23350 (N_23350,N_22773,N_22964);
or U23351 (N_23351,N_22781,N_22830);
nand U23352 (N_23352,N_22960,N_22504);
nor U23353 (N_23353,N_22889,N_22501);
and U23354 (N_23354,N_22846,N_22531);
or U23355 (N_23355,N_22693,N_22521);
xor U23356 (N_23356,N_22899,N_22581);
nand U23357 (N_23357,N_22573,N_22858);
nand U23358 (N_23358,N_22664,N_22873);
nor U23359 (N_23359,N_22552,N_22998);
or U23360 (N_23360,N_22573,N_22571);
and U23361 (N_23361,N_22928,N_22965);
or U23362 (N_23362,N_22742,N_22675);
and U23363 (N_23363,N_22990,N_22790);
xnor U23364 (N_23364,N_22920,N_22983);
or U23365 (N_23365,N_22773,N_22952);
or U23366 (N_23366,N_22591,N_22983);
or U23367 (N_23367,N_22653,N_22741);
or U23368 (N_23368,N_22533,N_22633);
and U23369 (N_23369,N_22621,N_22712);
or U23370 (N_23370,N_22801,N_22918);
and U23371 (N_23371,N_22605,N_22911);
and U23372 (N_23372,N_22814,N_22847);
xor U23373 (N_23373,N_22760,N_22654);
xnor U23374 (N_23374,N_22998,N_22599);
or U23375 (N_23375,N_22552,N_22827);
xnor U23376 (N_23376,N_22921,N_22560);
and U23377 (N_23377,N_22529,N_22772);
or U23378 (N_23378,N_22827,N_22777);
and U23379 (N_23379,N_22561,N_22693);
or U23380 (N_23380,N_22728,N_22507);
and U23381 (N_23381,N_22509,N_22949);
or U23382 (N_23382,N_22987,N_22947);
nand U23383 (N_23383,N_22908,N_22643);
xor U23384 (N_23384,N_22775,N_22972);
or U23385 (N_23385,N_22745,N_22948);
xor U23386 (N_23386,N_22552,N_22554);
xor U23387 (N_23387,N_22666,N_22738);
nor U23388 (N_23388,N_22523,N_22970);
nand U23389 (N_23389,N_22764,N_22861);
nor U23390 (N_23390,N_22654,N_22921);
nand U23391 (N_23391,N_22701,N_22558);
or U23392 (N_23392,N_22603,N_22737);
or U23393 (N_23393,N_22559,N_22544);
xnor U23394 (N_23394,N_22754,N_22537);
nand U23395 (N_23395,N_22501,N_22672);
or U23396 (N_23396,N_22545,N_22740);
nor U23397 (N_23397,N_22860,N_22858);
nand U23398 (N_23398,N_22646,N_22587);
xor U23399 (N_23399,N_22938,N_22978);
nor U23400 (N_23400,N_22936,N_22673);
and U23401 (N_23401,N_22659,N_22878);
and U23402 (N_23402,N_22870,N_22759);
xor U23403 (N_23403,N_22597,N_22713);
xor U23404 (N_23404,N_22617,N_22948);
xnor U23405 (N_23405,N_22583,N_22673);
or U23406 (N_23406,N_22689,N_22713);
nor U23407 (N_23407,N_22609,N_22764);
nand U23408 (N_23408,N_22906,N_22946);
xor U23409 (N_23409,N_22953,N_22728);
nand U23410 (N_23410,N_22767,N_22938);
nor U23411 (N_23411,N_22844,N_22546);
nand U23412 (N_23412,N_22797,N_22599);
xor U23413 (N_23413,N_22669,N_22904);
or U23414 (N_23414,N_22525,N_22537);
nand U23415 (N_23415,N_22999,N_22966);
or U23416 (N_23416,N_22515,N_22787);
and U23417 (N_23417,N_22586,N_22847);
and U23418 (N_23418,N_22732,N_22765);
xnor U23419 (N_23419,N_22609,N_22553);
and U23420 (N_23420,N_22585,N_22752);
or U23421 (N_23421,N_22764,N_22535);
nand U23422 (N_23422,N_22926,N_22860);
nor U23423 (N_23423,N_22824,N_22957);
nand U23424 (N_23424,N_22560,N_22789);
nor U23425 (N_23425,N_22958,N_22502);
xnor U23426 (N_23426,N_22951,N_22531);
nand U23427 (N_23427,N_22864,N_22741);
nor U23428 (N_23428,N_22600,N_22864);
nor U23429 (N_23429,N_22844,N_22830);
xnor U23430 (N_23430,N_22824,N_22818);
and U23431 (N_23431,N_22766,N_22591);
and U23432 (N_23432,N_22659,N_22766);
nand U23433 (N_23433,N_22672,N_22666);
and U23434 (N_23434,N_22638,N_22630);
and U23435 (N_23435,N_22771,N_22879);
nand U23436 (N_23436,N_22891,N_22862);
and U23437 (N_23437,N_22818,N_22577);
nor U23438 (N_23438,N_22576,N_22772);
and U23439 (N_23439,N_22797,N_22788);
nor U23440 (N_23440,N_22860,N_22988);
xnor U23441 (N_23441,N_22813,N_22669);
nand U23442 (N_23442,N_22884,N_22795);
nor U23443 (N_23443,N_22699,N_22714);
nor U23444 (N_23444,N_22771,N_22774);
nor U23445 (N_23445,N_22954,N_22610);
xor U23446 (N_23446,N_22910,N_22842);
xnor U23447 (N_23447,N_22844,N_22801);
nand U23448 (N_23448,N_22709,N_22608);
xnor U23449 (N_23449,N_22990,N_22896);
or U23450 (N_23450,N_22726,N_22972);
xor U23451 (N_23451,N_22967,N_22525);
nand U23452 (N_23452,N_22868,N_22974);
nand U23453 (N_23453,N_22799,N_22870);
nor U23454 (N_23454,N_22896,N_22703);
xnor U23455 (N_23455,N_22682,N_22545);
and U23456 (N_23456,N_22890,N_22717);
nor U23457 (N_23457,N_22638,N_22825);
nand U23458 (N_23458,N_22639,N_22867);
and U23459 (N_23459,N_22736,N_22803);
and U23460 (N_23460,N_22811,N_22609);
nor U23461 (N_23461,N_22607,N_22719);
nor U23462 (N_23462,N_22895,N_22753);
and U23463 (N_23463,N_22512,N_22987);
xor U23464 (N_23464,N_22592,N_22526);
or U23465 (N_23465,N_22992,N_22867);
or U23466 (N_23466,N_22924,N_22507);
or U23467 (N_23467,N_22674,N_22700);
and U23468 (N_23468,N_22859,N_22829);
or U23469 (N_23469,N_22661,N_22510);
and U23470 (N_23470,N_22879,N_22920);
xor U23471 (N_23471,N_22745,N_22765);
or U23472 (N_23472,N_22892,N_22770);
and U23473 (N_23473,N_22821,N_22993);
or U23474 (N_23474,N_22512,N_22617);
xor U23475 (N_23475,N_22686,N_22662);
nor U23476 (N_23476,N_22540,N_22749);
nor U23477 (N_23477,N_22664,N_22747);
xor U23478 (N_23478,N_22535,N_22508);
xor U23479 (N_23479,N_22640,N_22685);
nand U23480 (N_23480,N_22548,N_22522);
nor U23481 (N_23481,N_22955,N_22690);
nand U23482 (N_23482,N_22648,N_22832);
nand U23483 (N_23483,N_22543,N_22545);
nor U23484 (N_23484,N_22597,N_22550);
nor U23485 (N_23485,N_22645,N_22991);
nand U23486 (N_23486,N_22868,N_22750);
nand U23487 (N_23487,N_22655,N_22717);
xor U23488 (N_23488,N_22597,N_22694);
nand U23489 (N_23489,N_22677,N_22761);
or U23490 (N_23490,N_22869,N_22637);
or U23491 (N_23491,N_22616,N_22683);
or U23492 (N_23492,N_22724,N_22981);
nand U23493 (N_23493,N_22730,N_22528);
nand U23494 (N_23494,N_22849,N_22535);
nor U23495 (N_23495,N_22530,N_22605);
and U23496 (N_23496,N_22826,N_22563);
or U23497 (N_23497,N_22926,N_22670);
or U23498 (N_23498,N_22759,N_22529);
nor U23499 (N_23499,N_22973,N_22751);
and U23500 (N_23500,N_23003,N_23207);
nor U23501 (N_23501,N_23216,N_23442);
xnor U23502 (N_23502,N_23149,N_23370);
nand U23503 (N_23503,N_23336,N_23381);
nor U23504 (N_23504,N_23300,N_23431);
nor U23505 (N_23505,N_23103,N_23189);
and U23506 (N_23506,N_23126,N_23254);
nor U23507 (N_23507,N_23277,N_23340);
nand U23508 (N_23508,N_23470,N_23422);
nand U23509 (N_23509,N_23112,N_23265);
and U23510 (N_23510,N_23440,N_23402);
nor U23511 (N_23511,N_23233,N_23087);
nand U23512 (N_23512,N_23161,N_23091);
xor U23513 (N_23513,N_23141,N_23117);
xnor U23514 (N_23514,N_23223,N_23373);
or U23515 (N_23515,N_23142,N_23342);
nand U23516 (N_23516,N_23248,N_23485);
xnor U23517 (N_23517,N_23190,N_23101);
or U23518 (N_23518,N_23034,N_23261);
xnor U23519 (N_23519,N_23455,N_23097);
nor U23520 (N_23520,N_23408,N_23247);
nand U23521 (N_23521,N_23317,N_23219);
xnor U23522 (N_23522,N_23390,N_23081);
nand U23523 (N_23523,N_23028,N_23228);
xnor U23524 (N_23524,N_23295,N_23169);
or U23525 (N_23525,N_23392,N_23365);
and U23526 (N_23526,N_23287,N_23058);
and U23527 (N_23527,N_23291,N_23038);
xnor U23528 (N_23528,N_23331,N_23154);
nor U23529 (N_23529,N_23480,N_23472);
nand U23530 (N_23530,N_23089,N_23242);
or U23531 (N_23531,N_23118,N_23129);
and U23532 (N_23532,N_23498,N_23096);
or U23533 (N_23533,N_23424,N_23380);
or U23534 (N_23534,N_23030,N_23301);
xnor U23535 (N_23535,N_23187,N_23397);
and U23536 (N_23536,N_23086,N_23309);
xor U23537 (N_23537,N_23150,N_23155);
xor U23538 (N_23538,N_23235,N_23490);
nor U23539 (N_23539,N_23180,N_23040);
and U23540 (N_23540,N_23178,N_23196);
xnor U23541 (N_23541,N_23256,N_23182);
nor U23542 (N_23542,N_23462,N_23352);
nor U23543 (N_23543,N_23362,N_23115);
nand U23544 (N_23544,N_23446,N_23168);
and U23545 (N_23545,N_23374,N_23227);
or U23546 (N_23546,N_23218,N_23104);
xor U23547 (N_23547,N_23298,N_23044);
and U23548 (N_23548,N_23361,N_23023);
xnor U23549 (N_23549,N_23267,N_23240);
nand U23550 (N_23550,N_23131,N_23499);
or U23551 (N_23551,N_23092,N_23139);
or U23552 (N_23552,N_23318,N_23035);
nand U23553 (N_23553,N_23222,N_23324);
or U23554 (N_23554,N_23181,N_23201);
or U23555 (N_23555,N_23215,N_23013);
nor U23556 (N_23556,N_23193,N_23010);
or U23557 (N_23557,N_23417,N_23311);
or U23558 (N_23558,N_23186,N_23458);
xnor U23559 (N_23559,N_23330,N_23494);
nand U23560 (N_23560,N_23429,N_23226);
xor U23561 (N_23561,N_23310,N_23478);
xor U23562 (N_23562,N_23477,N_23461);
and U23563 (N_23563,N_23171,N_23453);
nor U23564 (N_23564,N_23093,N_23204);
and U23565 (N_23565,N_23275,N_23366);
xor U23566 (N_23566,N_23276,N_23338);
nand U23567 (N_23567,N_23077,N_23341);
or U23568 (N_23568,N_23120,N_23349);
nand U23569 (N_23569,N_23107,N_23283);
xnor U23570 (N_23570,N_23136,N_23414);
or U23571 (N_23571,N_23019,N_23386);
nand U23572 (N_23572,N_23050,N_23083);
nand U23573 (N_23573,N_23128,N_23290);
nand U23574 (N_23574,N_23151,N_23108);
or U23575 (N_23575,N_23060,N_23243);
nor U23576 (N_23576,N_23444,N_23153);
xnor U23577 (N_23577,N_23114,N_23017);
nand U23578 (N_23578,N_23172,N_23075);
and U23579 (N_23579,N_23231,N_23213);
nor U23580 (N_23580,N_23183,N_23328);
nor U23581 (N_23581,N_23005,N_23007);
nor U23582 (N_23582,N_23157,N_23135);
nand U23583 (N_23583,N_23438,N_23111);
nor U23584 (N_23584,N_23071,N_23257);
or U23585 (N_23585,N_23162,N_23140);
nand U23586 (N_23586,N_23170,N_23449);
nand U23587 (N_23587,N_23122,N_23069);
nor U23588 (N_23588,N_23173,N_23369);
or U23589 (N_23589,N_23329,N_23066);
nor U23590 (N_23590,N_23262,N_23379);
or U23591 (N_23591,N_23441,N_23133);
and U23592 (N_23592,N_23082,N_23410);
nand U23593 (N_23593,N_23351,N_23259);
or U23594 (N_23594,N_23008,N_23177);
nor U23595 (N_23595,N_23281,N_23258);
or U23596 (N_23596,N_23127,N_23016);
nor U23597 (N_23597,N_23405,N_23347);
nor U23598 (N_23598,N_23305,N_23252);
and U23599 (N_23599,N_23466,N_23430);
nor U23600 (N_23600,N_23230,N_23326);
and U23601 (N_23601,N_23100,N_23263);
and U23602 (N_23602,N_23481,N_23288);
nor U23603 (N_23603,N_23110,N_23316);
xor U23604 (N_23604,N_23320,N_23345);
nor U23605 (N_23605,N_23260,N_23297);
and U23606 (N_23606,N_23421,N_23018);
nor U23607 (N_23607,N_23033,N_23443);
nand U23608 (N_23608,N_23280,N_23428);
xnor U23609 (N_23609,N_23067,N_23109);
and U23610 (N_23610,N_23073,N_23469);
xnor U23611 (N_23611,N_23147,N_23105);
xnor U23612 (N_23612,N_23409,N_23388);
xor U23613 (N_23613,N_23367,N_23074);
and U23614 (N_23614,N_23085,N_23099);
nand U23615 (N_23615,N_23184,N_23335);
and U23616 (N_23616,N_23296,N_23202);
or U23617 (N_23617,N_23197,N_23179);
nand U23618 (N_23618,N_23354,N_23237);
or U23619 (N_23619,N_23253,N_23394);
or U23620 (N_23620,N_23403,N_23460);
and U23621 (N_23621,N_23239,N_23493);
xor U23622 (N_23622,N_23479,N_23415);
nor U23623 (N_23623,N_23489,N_23425);
xnor U23624 (N_23624,N_23176,N_23212);
nor U23625 (N_23625,N_23175,N_23464);
and U23626 (N_23626,N_23113,N_23163);
and U23627 (N_23627,N_23393,N_23174);
xor U23628 (N_23628,N_23051,N_23241);
and U23629 (N_23629,N_23497,N_23188);
and U23630 (N_23630,N_23418,N_23080);
nor U23631 (N_23631,N_23344,N_23439);
or U23632 (N_23632,N_23383,N_23395);
xnor U23633 (N_23633,N_23057,N_23491);
nor U23634 (N_23634,N_23321,N_23268);
nand U23635 (N_23635,N_23286,N_23377);
nor U23636 (N_23636,N_23376,N_23400);
or U23637 (N_23637,N_23468,N_23307);
nor U23638 (N_23638,N_23411,N_23052);
or U23639 (N_23639,N_23121,N_23124);
and U23640 (N_23640,N_23088,N_23378);
and U23641 (N_23641,N_23015,N_23358);
nor U23642 (N_23642,N_23244,N_23220);
nor U23643 (N_23643,N_23482,N_23137);
or U23644 (N_23644,N_23236,N_23200);
or U23645 (N_23645,N_23055,N_23284);
and U23646 (N_23646,N_23056,N_23021);
xor U23647 (N_23647,N_23156,N_23313);
xor U23648 (N_23648,N_23473,N_23053);
xor U23649 (N_23649,N_23457,N_23245);
and U23650 (N_23650,N_23487,N_23238);
nand U23651 (N_23651,N_23483,N_23266);
and U23652 (N_23652,N_23484,N_23454);
and U23653 (N_23653,N_23094,N_23372);
xnor U23654 (N_23654,N_23492,N_23356);
nor U23655 (N_23655,N_23315,N_23125);
xnor U23656 (N_23656,N_23199,N_23399);
xor U23657 (N_23657,N_23269,N_23339);
nand U23658 (N_23658,N_23046,N_23043);
xnor U23659 (N_23659,N_23130,N_23278);
nor U23660 (N_23660,N_23041,N_23232);
nand U23661 (N_23661,N_23045,N_23203);
or U23662 (N_23662,N_23138,N_23387);
or U23663 (N_23663,N_23412,N_23273);
and U23664 (N_23664,N_23420,N_23319);
or U23665 (N_23665,N_23450,N_23123);
and U23666 (N_23666,N_23433,N_23132);
xnor U23667 (N_23667,N_23078,N_23471);
nand U23668 (N_23668,N_23039,N_23465);
or U23669 (N_23669,N_23432,N_23452);
and U23670 (N_23670,N_23285,N_23012);
xnor U23671 (N_23671,N_23146,N_23049);
and U23672 (N_23672,N_23225,N_23385);
or U23673 (N_23673,N_23002,N_23448);
xnor U23674 (N_23674,N_23363,N_23032);
or U23675 (N_23675,N_23025,N_23072);
xnor U23676 (N_23676,N_23195,N_23334);
xor U23677 (N_23677,N_23217,N_23014);
or U23678 (N_23678,N_23191,N_23264);
nor U23679 (N_23679,N_23333,N_23210);
or U23680 (N_23680,N_23144,N_23348);
and U23681 (N_23681,N_23360,N_23355);
and U23682 (N_23682,N_23293,N_23134);
nand U23683 (N_23683,N_23022,N_23368);
nor U23684 (N_23684,N_23416,N_23160);
nor U23685 (N_23685,N_23451,N_23337);
nor U23686 (N_23686,N_23221,N_23084);
or U23687 (N_23687,N_23389,N_23185);
nor U23688 (N_23688,N_23322,N_23206);
and U23689 (N_23689,N_23048,N_23068);
xor U23690 (N_23690,N_23167,N_23192);
xor U23691 (N_23691,N_23475,N_23274);
and U23692 (N_23692,N_23289,N_23061);
or U23693 (N_23693,N_23398,N_23435);
or U23694 (N_23694,N_23312,N_23353);
or U23695 (N_23695,N_23119,N_23364);
nand U23696 (N_23696,N_23194,N_23371);
xnor U23697 (N_23697,N_23406,N_23343);
xnor U23698 (N_23698,N_23476,N_23255);
nand U23699 (N_23699,N_23325,N_23426);
nor U23700 (N_23700,N_23198,N_23314);
or U23701 (N_23701,N_23357,N_23024);
or U23702 (N_23702,N_23495,N_23098);
and U23703 (N_23703,N_23159,N_23423);
nor U23704 (N_23704,N_23419,N_23294);
nor U23705 (N_23705,N_23165,N_23224);
and U23706 (N_23706,N_23059,N_23346);
nand U23707 (N_23707,N_23279,N_23020);
or U23708 (N_23708,N_23384,N_23407);
nor U23709 (N_23709,N_23359,N_23308);
nor U23710 (N_23710,N_23404,N_23303);
nor U23711 (N_23711,N_23401,N_23076);
nand U23712 (N_23712,N_23064,N_23486);
or U23713 (N_23713,N_23026,N_23001);
xnor U23714 (N_23714,N_23158,N_23332);
nand U23715 (N_23715,N_23447,N_23095);
nor U23716 (N_23716,N_23234,N_23270);
nand U23717 (N_23717,N_23292,N_23164);
and U23718 (N_23718,N_23063,N_23145);
nor U23719 (N_23719,N_23116,N_23211);
nand U23720 (N_23720,N_23306,N_23047);
xnor U23721 (N_23721,N_23434,N_23413);
or U23722 (N_23722,N_23090,N_23036);
or U23723 (N_23723,N_23029,N_23246);
and U23724 (N_23724,N_23323,N_23391);
xnor U23725 (N_23725,N_23102,N_23079);
nand U23726 (N_23726,N_23250,N_23437);
nor U23727 (N_23727,N_23272,N_23037);
nor U23728 (N_23728,N_23299,N_23282);
or U23729 (N_23729,N_23350,N_23463);
nor U23730 (N_23730,N_23427,N_23106);
nand U23731 (N_23731,N_23031,N_23143);
xnor U23732 (N_23732,N_23249,N_23065);
nor U23733 (N_23733,N_23208,N_23152);
xor U23734 (N_23734,N_23327,N_23496);
nand U23735 (N_23735,N_23488,N_23436);
or U23736 (N_23736,N_23467,N_23027);
nor U23737 (N_23737,N_23205,N_23474);
xor U23738 (N_23738,N_23302,N_23148);
nor U23739 (N_23739,N_23445,N_23271);
xor U23740 (N_23740,N_23011,N_23382);
xor U23741 (N_23741,N_23042,N_23009);
or U23742 (N_23742,N_23375,N_23006);
or U23743 (N_23743,N_23004,N_23304);
or U23744 (N_23744,N_23000,N_23166);
nand U23745 (N_23745,N_23456,N_23054);
nor U23746 (N_23746,N_23396,N_23070);
nand U23747 (N_23747,N_23062,N_23214);
and U23748 (N_23748,N_23251,N_23209);
nor U23749 (N_23749,N_23459,N_23229);
or U23750 (N_23750,N_23033,N_23473);
nor U23751 (N_23751,N_23297,N_23411);
and U23752 (N_23752,N_23169,N_23377);
nand U23753 (N_23753,N_23169,N_23387);
or U23754 (N_23754,N_23230,N_23077);
nor U23755 (N_23755,N_23247,N_23335);
xnor U23756 (N_23756,N_23050,N_23041);
or U23757 (N_23757,N_23447,N_23153);
and U23758 (N_23758,N_23457,N_23458);
and U23759 (N_23759,N_23193,N_23123);
nand U23760 (N_23760,N_23243,N_23419);
and U23761 (N_23761,N_23418,N_23185);
and U23762 (N_23762,N_23082,N_23227);
and U23763 (N_23763,N_23264,N_23326);
nor U23764 (N_23764,N_23031,N_23056);
or U23765 (N_23765,N_23168,N_23221);
or U23766 (N_23766,N_23432,N_23441);
nand U23767 (N_23767,N_23024,N_23219);
nand U23768 (N_23768,N_23170,N_23245);
and U23769 (N_23769,N_23028,N_23471);
or U23770 (N_23770,N_23489,N_23149);
nand U23771 (N_23771,N_23481,N_23271);
or U23772 (N_23772,N_23047,N_23416);
or U23773 (N_23773,N_23284,N_23325);
nand U23774 (N_23774,N_23209,N_23077);
or U23775 (N_23775,N_23025,N_23148);
and U23776 (N_23776,N_23437,N_23255);
and U23777 (N_23777,N_23347,N_23098);
or U23778 (N_23778,N_23401,N_23348);
nor U23779 (N_23779,N_23406,N_23232);
xnor U23780 (N_23780,N_23130,N_23061);
xor U23781 (N_23781,N_23076,N_23063);
or U23782 (N_23782,N_23091,N_23189);
and U23783 (N_23783,N_23318,N_23208);
nand U23784 (N_23784,N_23324,N_23097);
nor U23785 (N_23785,N_23273,N_23106);
xnor U23786 (N_23786,N_23478,N_23270);
or U23787 (N_23787,N_23418,N_23078);
xor U23788 (N_23788,N_23176,N_23092);
xnor U23789 (N_23789,N_23316,N_23233);
or U23790 (N_23790,N_23222,N_23359);
nor U23791 (N_23791,N_23149,N_23119);
nand U23792 (N_23792,N_23144,N_23337);
and U23793 (N_23793,N_23258,N_23416);
or U23794 (N_23794,N_23402,N_23170);
xor U23795 (N_23795,N_23330,N_23095);
nor U23796 (N_23796,N_23084,N_23012);
xnor U23797 (N_23797,N_23498,N_23330);
nand U23798 (N_23798,N_23093,N_23450);
or U23799 (N_23799,N_23470,N_23472);
nor U23800 (N_23800,N_23160,N_23316);
nand U23801 (N_23801,N_23102,N_23274);
or U23802 (N_23802,N_23018,N_23416);
nor U23803 (N_23803,N_23226,N_23202);
nand U23804 (N_23804,N_23107,N_23039);
xor U23805 (N_23805,N_23104,N_23231);
nand U23806 (N_23806,N_23143,N_23446);
or U23807 (N_23807,N_23222,N_23184);
nor U23808 (N_23808,N_23459,N_23024);
nand U23809 (N_23809,N_23376,N_23135);
or U23810 (N_23810,N_23375,N_23330);
xnor U23811 (N_23811,N_23472,N_23029);
nand U23812 (N_23812,N_23231,N_23252);
and U23813 (N_23813,N_23190,N_23181);
xor U23814 (N_23814,N_23355,N_23163);
or U23815 (N_23815,N_23254,N_23092);
xor U23816 (N_23816,N_23249,N_23313);
and U23817 (N_23817,N_23196,N_23219);
nor U23818 (N_23818,N_23025,N_23084);
or U23819 (N_23819,N_23356,N_23357);
xor U23820 (N_23820,N_23333,N_23278);
nor U23821 (N_23821,N_23269,N_23412);
xnor U23822 (N_23822,N_23194,N_23168);
and U23823 (N_23823,N_23027,N_23123);
xor U23824 (N_23824,N_23260,N_23186);
xor U23825 (N_23825,N_23416,N_23009);
nor U23826 (N_23826,N_23014,N_23011);
and U23827 (N_23827,N_23389,N_23252);
and U23828 (N_23828,N_23119,N_23495);
nor U23829 (N_23829,N_23219,N_23494);
and U23830 (N_23830,N_23438,N_23128);
or U23831 (N_23831,N_23439,N_23185);
nand U23832 (N_23832,N_23206,N_23187);
xor U23833 (N_23833,N_23308,N_23187);
xor U23834 (N_23834,N_23491,N_23179);
xor U23835 (N_23835,N_23298,N_23341);
or U23836 (N_23836,N_23179,N_23400);
and U23837 (N_23837,N_23194,N_23010);
xnor U23838 (N_23838,N_23161,N_23012);
nand U23839 (N_23839,N_23343,N_23301);
or U23840 (N_23840,N_23290,N_23449);
and U23841 (N_23841,N_23025,N_23284);
and U23842 (N_23842,N_23373,N_23266);
and U23843 (N_23843,N_23454,N_23265);
and U23844 (N_23844,N_23105,N_23011);
and U23845 (N_23845,N_23393,N_23402);
and U23846 (N_23846,N_23480,N_23112);
nand U23847 (N_23847,N_23112,N_23204);
xor U23848 (N_23848,N_23188,N_23189);
xnor U23849 (N_23849,N_23307,N_23480);
and U23850 (N_23850,N_23346,N_23483);
nand U23851 (N_23851,N_23006,N_23352);
nor U23852 (N_23852,N_23286,N_23462);
or U23853 (N_23853,N_23490,N_23342);
xnor U23854 (N_23854,N_23272,N_23059);
xor U23855 (N_23855,N_23470,N_23036);
xnor U23856 (N_23856,N_23138,N_23482);
nand U23857 (N_23857,N_23206,N_23117);
and U23858 (N_23858,N_23285,N_23121);
nor U23859 (N_23859,N_23163,N_23120);
and U23860 (N_23860,N_23488,N_23338);
and U23861 (N_23861,N_23306,N_23484);
or U23862 (N_23862,N_23042,N_23479);
or U23863 (N_23863,N_23008,N_23341);
nand U23864 (N_23864,N_23289,N_23290);
xor U23865 (N_23865,N_23044,N_23295);
nand U23866 (N_23866,N_23124,N_23473);
or U23867 (N_23867,N_23362,N_23329);
or U23868 (N_23868,N_23272,N_23312);
and U23869 (N_23869,N_23208,N_23292);
or U23870 (N_23870,N_23063,N_23155);
nand U23871 (N_23871,N_23395,N_23126);
nor U23872 (N_23872,N_23401,N_23247);
nand U23873 (N_23873,N_23120,N_23148);
and U23874 (N_23874,N_23004,N_23246);
nor U23875 (N_23875,N_23199,N_23000);
and U23876 (N_23876,N_23353,N_23019);
and U23877 (N_23877,N_23268,N_23193);
nor U23878 (N_23878,N_23441,N_23150);
xnor U23879 (N_23879,N_23329,N_23071);
and U23880 (N_23880,N_23112,N_23378);
nor U23881 (N_23881,N_23268,N_23459);
and U23882 (N_23882,N_23259,N_23251);
xnor U23883 (N_23883,N_23050,N_23376);
xor U23884 (N_23884,N_23275,N_23404);
or U23885 (N_23885,N_23025,N_23200);
xor U23886 (N_23886,N_23041,N_23098);
xnor U23887 (N_23887,N_23416,N_23241);
xnor U23888 (N_23888,N_23360,N_23035);
and U23889 (N_23889,N_23272,N_23471);
or U23890 (N_23890,N_23378,N_23093);
or U23891 (N_23891,N_23210,N_23417);
nor U23892 (N_23892,N_23153,N_23409);
nor U23893 (N_23893,N_23199,N_23469);
nor U23894 (N_23894,N_23066,N_23055);
nor U23895 (N_23895,N_23247,N_23071);
nand U23896 (N_23896,N_23168,N_23295);
nor U23897 (N_23897,N_23324,N_23076);
or U23898 (N_23898,N_23163,N_23490);
or U23899 (N_23899,N_23328,N_23376);
and U23900 (N_23900,N_23303,N_23454);
or U23901 (N_23901,N_23494,N_23095);
nor U23902 (N_23902,N_23487,N_23232);
and U23903 (N_23903,N_23268,N_23095);
nor U23904 (N_23904,N_23439,N_23214);
xnor U23905 (N_23905,N_23237,N_23072);
or U23906 (N_23906,N_23393,N_23449);
xor U23907 (N_23907,N_23026,N_23420);
or U23908 (N_23908,N_23488,N_23403);
xor U23909 (N_23909,N_23436,N_23264);
nor U23910 (N_23910,N_23187,N_23470);
nand U23911 (N_23911,N_23494,N_23360);
nand U23912 (N_23912,N_23493,N_23245);
nor U23913 (N_23913,N_23181,N_23046);
and U23914 (N_23914,N_23045,N_23225);
xor U23915 (N_23915,N_23073,N_23309);
nor U23916 (N_23916,N_23340,N_23289);
or U23917 (N_23917,N_23457,N_23135);
nor U23918 (N_23918,N_23262,N_23389);
xor U23919 (N_23919,N_23154,N_23252);
and U23920 (N_23920,N_23246,N_23024);
or U23921 (N_23921,N_23410,N_23499);
or U23922 (N_23922,N_23011,N_23261);
xor U23923 (N_23923,N_23278,N_23038);
xor U23924 (N_23924,N_23131,N_23208);
or U23925 (N_23925,N_23394,N_23430);
nor U23926 (N_23926,N_23398,N_23264);
and U23927 (N_23927,N_23372,N_23344);
and U23928 (N_23928,N_23350,N_23230);
and U23929 (N_23929,N_23337,N_23056);
or U23930 (N_23930,N_23319,N_23169);
and U23931 (N_23931,N_23108,N_23252);
or U23932 (N_23932,N_23282,N_23191);
xor U23933 (N_23933,N_23403,N_23060);
or U23934 (N_23934,N_23283,N_23230);
nor U23935 (N_23935,N_23063,N_23373);
nand U23936 (N_23936,N_23415,N_23150);
xor U23937 (N_23937,N_23203,N_23442);
xnor U23938 (N_23938,N_23223,N_23375);
nor U23939 (N_23939,N_23316,N_23388);
or U23940 (N_23940,N_23273,N_23025);
nor U23941 (N_23941,N_23470,N_23369);
xnor U23942 (N_23942,N_23388,N_23405);
xor U23943 (N_23943,N_23040,N_23174);
nand U23944 (N_23944,N_23469,N_23222);
and U23945 (N_23945,N_23042,N_23495);
xnor U23946 (N_23946,N_23265,N_23226);
and U23947 (N_23947,N_23229,N_23016);
nand U23948 (N_23948,N_23499,N_23303);
and U23949 (N_23949,N_23221,N_23474);
nor U23950 (N_23950,N_23197,N_23444);
xor U23951 (N_23951,N_23310,N_23486);
or U23952 (N_23952,N_23030,N_23331);
nand U23953 (N_23953,N_23373,N_23331);
nor U23954 (N_23954,N_23182,N_23025);
or U23955 (N_23955,N_23476,N_23241);
xor U23956 (N_23956,N_23494,N_23166);
nand U23957 (N_23957,N_23229,N_23387);
nand U23958 (N_23958,N_23324,N_23011);
or U23959 (N_23959,N_23173,N_23398);
xnor U23960 (N_23960,N_23367,N_23040);
nor U23961 (N_23961,N_23459,N_23418);
nor U23962 (N_23962,N_23012,N_23198);
nand U23963 (N_23963,N_23159,N_23454);
nand U23964 (N_23964,N_23005,N_23224);
and U23965 (N_23965,N_23175,N_23375);
and U23966 (N_23966,N_23302,N_23443);
and U23967 (N_23967,N_23435,N_23338);
or U23968 (N_23968,N_23260,N_23430);
xor U23969 (N_23969,N_23474,N_23054);
and U23970 (N_23970,N_23322,N_23029);
or U23971 (N_23971,N_23373,N_23297);
or U23972 (N_23972,N_23000,N_23409);
xor U23973 (N_23973,N_23327,N_23025);
nand U23974 (N_23974,N_23400,N_23269);
and U23975 (N_23975,N_23357,N_23078);
xnor U23976 (N_23976,N_23182,N_23297);
xnor U23977 (N_23977,N_23459,N_23405);
or U23978 (N_23978,N_23185,N_23206);
nor U23979 (N_23979,N_23306,N_23491);
nand U23980 (N_23980,N_23240,N_23173);
nand U23981 (N_23981,N_23315,N_23088);
or U23982 (N_23982,N_23447,N_23052);
nor U23983 (N_23983,N_23216,N_23196);
xor U23984 (N_23984,N_23161,N_23074);
or U23985 (N_23985,N_23276,N_23102);
nor U23986 (N_23986,N_23416,N_23434);
nand U23987 (N_23987,N_23160,N_23216);
nand U23988 (N_23988,N_23183,N_23163);
nor U23989 (N_23989,N_23074,N_23033);
nand U23990 (N_23990,N_23339,N_23272);
nand U23991 (N_23991,N_23054,N_23350);
nor U23992 (N_23992,N_23177,N_23345);
and U23993 (N_23993,N_23462,N_23327);
or U23994 (N_23994,N_23131,N_23009);
nand U23995 (N_23995,N_23335,N_23258);
and U23996 (N_23996,N_23086,N_23094);
xor U23997 (N_23997,N_23286,N_23039);
or U23998 (N_23998,N_23030,N_23440);
and U23999 (N_23999,N_23433,N_23362);
nand U24000 (N_24000,N_23526,N_23605);
nand U24001 (N_24001,N_23715,N_23887);
xnor U24002 (N_24002,N_23676,N_23838);
nor U24003 (N_24003,N_23757,N_23942);
nand U24004 (N_24004,N_23567,N_23731);
or U24005 (N_24005,N_23694,N_23827);
xor U24006 (N_24006,N_23535,N_23790);
or U24007 (N_24007,N_23699,N_23750);
and U24008 (N_24008,N_23586,N_23821);
or U24009 (N_24009,N_23621,N_23990);
xnor U24010 (N_24010,N_23620,N_23582);
xnor U24011 (N_24011,N_23890,N_23716);
nor U24012 (N_24012,N_23612,N_23880);
nor U24013 (N_24013,N_23579,N_23834);
and U24014 (N_24014,N_23888,N_23979);
and U24015 (N_24015,N_23957,N_23743);
nor U24016 (N_24016,N_23938,N_23769);
xor U24017 (N_24017,N_23613,N_23517);
xnor U24018 (N_24018,N_23959,N_23958);
or U24019 (N_24019,N_23984,N_23639);
xnor U24020 (N_24020,N_23799,N_23983);
or U24021 (N_24021,N_23927,N_23812);
nor U24022 (N_24022,N_23875,N_23836);
nor U24023 (N_24023,N_23987,N_23897);
nand U24024 (N_24024,N_23903,N_23645);
nand U24025 (N_24025,N_23633,N_23504);
or U24026 (N_24026,N_23801,N_23764);
or U24027 (N_24027,N_23525,N_23720);
and U24028 (N_24028,N_23532,N_23963);
xnor U24029 (N_24029,N_23693,N_23843);
xnor U24030 (N_24030,N_23617,N_23895);
or U24031 (N_24031,N_23929,N_23690);
nor U24032 (N_24032,N_23589,N_23695);
and U24033 (N_24033,N_23865,N_23817);
nand U24034 (N_24034,N_23892,N_23746);
or U24035 (N_24035,N_23629,N_23671);
nor U24036 (N_24036,N_23980,N_23735);
nor U24037 (N_24037,N_23528,N_23505);
and U24038 (N_24038,N_23747,N_23792);
nor U24039 (N_24039,N_23849,N_23719);
or U24040 (N_24040,N_23833,N_23575);
nor U24041 (N_24041,N_23931,N_23919);
nand U24042 (N_24042,N_23922,N_23610);
xor U24043 (N_24043,N_23661,N_23891);
nand U24044 (N_24044,N_23564,N_23996);
and U24045 (N_24045,N_23732,N_23804);
xnor U24046 (N_24046,N_23837,N_23646);
nor U24047 (N_24047,N_23924,N_23728);
or U24048 (N_24048,N_23783,N_23755);
xor U24049 (N_24049,N_23828,N_23596);
or U24050 (N_24050,N_23855,N_23878);
xnor U24051 (N_24051,N_23513,N_23508);
or U24052 (N_24052,N_23889,N_23544);
xor U24053 (N_24053,N_23696,N_23642);
nand U24054 (N_24054,N_23763,N_23982);
xnor U24055 (N_24055,N_23847,N_23651);
xor U24056 (N_24056,N_23541,N_23970);
or U24057 (N_24057,N_23933,N_23944);
xor U24058 (N_24058,N_23717,N_23636);
or U24059 (N_24059,N_23823,N_23785);
or U24060 (N_24060,N_23820,N_23722);
xor U24061 (N_24061,N_23592,N_23687);
nand U24062 (N_24062,N_23818,N_23908);
nand U24063 (N_24063,N_23991,N_23688);
or U24064 (N_24064,N_23653,N_23861);
xnor U24065 (N_24065,N_23604,N_23992);
and U24066 (N_24066,N_23733,N_23576);
or U24067 (N_24067,N_23841,N_23704);
and U24068 (N_24068,N_23913,N_23697);
nor U24069 (N_24069,N_23530,N_23635);
nand U24070 (N_24070,N_23862,N_23973);
and U24071 (N_24071,N_23680,N_23802);
nor U24072 (N_24072,N_23540,N_23725);
nand U24073 (N_24073,N_23910,N_23858);
or U24074 (N_24074,N_23914,N_23854);
nor U24075 (N_24075,N_23916,N_23758);
nand U24076 (N_24076,N_23711,N_23806);
or U24077 (N_24077,N_23864,N_23700);
and U24078 (N_24078,N_23898,N_23684);
and U24079 (N_24079,N_23807,N_23603);
xor U24080 (N_24080,N_23886,N_23516);
nand U24081 (N_24081,N_23707,N_23580);
xor U24082 (N_24082,N_23658,N_23870);
and U24083 (N_24083,N_23968,N_23630);
xnor U24084 (N_24084,N_23826,N_23930);
nor U24085 (N_24085,N_23718,N_23559);
nor U24086 (N_24086,N_23588,N_23730);
nor U24087 (N_24087,N_23714,N_23782);
and U24088 (N_24088,N_23593,N_23830);
nand U24089 (N_24089,N_23527,N_23840);
nand U24090 (N_24090,N_23668,N_23523);
xnor U24091 (N_24091,N_23831,N_23647);
and U24092 (N_24092,N_23558,N_23967);
nand U24093 (N_24093,N_23551,N_23573);
xor U24094 (N_24094,N_23839,N_23578);
or U24095 (N_24095,N_23925,N_23751);
nor U24096 (N_24096,N_23926,N_23951);
xor U24097 (N_24097,N_23917,N_23881);
nor U24098 (N_24098,N_23666,N_23737);
xnor U24099 (N_24099,N_23947,N_23591);
nor U24100 (N_24100,N_23872,N_23797);
nand U24101 (N_24101,N_23809,N_23616);
and U24102 (N_24102,N_23902,N_23899);
nor U24103 (N_24103,N_23997,N_23936);
or U24104 (N_24104,N_23637,N_23557);
nand U24105 (N_24105,N_23618,N_23698);
or U24106 (N_24106,N_23848,N_23901);
nand U24107 (N_24107,N_23904,N_23681);
xnor U24108 (N_24108,N_23813,N_23771);
or U24109 (N_24109,N_23608,N_23953);
or U24110 (N_24110,N_23561,N_23650);
nand U24111 (N_24111,N_23562,N_23853);
nor U24112 (N_24112,N_23954,N_23611);
nand U24113 (N_24113,N_23803,N_23524);
xor U24114 (N_24114,N_23814,N_23772);
nor U24115 (N_24115,N_23590,N_23538);
nand U24116 (N_24116,N_23577,N_23940);
nor U24117 (N_24117,N_23753,N_23631);
or U24118 (N_24118,N_23868,N_23943);
nand U24119 (N_24119,N_23531,N_23533);
nor U24120 (N_24120,N_23978,N_23542);
or U24121 (N_24121,N_23689,N_23655);
nor U24122 (N_24122,N_23547,N_23657);
nor U24123 (N_24123,N_23768,N_23955);
or U24124 (N_24124,N_23816,N_23822);
and U24125 (N_24125,N_23824,N_23789);
xor U24126 (N_24126,N_23765,N_23842);
and U24127 (N_24127,N_23598,N_23602);
xnor U24128 (N_24128,N_23866,N_23556);
nor U24129 (N_24129,N_23994,N_23972);
or U24130 (N_24130,N_23546,N_23705);
and U24131 (N_24131,N_23738,N_23566);
xor U24132 (N_24132,N_23572,N_23545);
nand U24133 (N_24133,N_23503,N_23601);
and U24134 (N_24134,N_23643,N_23739);
nor U24135 (N_24135,N_23784,N_23798);
nor U24136 (N_24136,N_23779,N_23918);
xnor U24137 (N_24137,N_23921,N_23548);
nor U24138 (N_24138,N_23752,N_23829);
and U24139 (N_24139,N_23665,N_23937);
and U24140 (N_24140,N_23932,N_23835);
or U24141 (N_24141,N_23894,N_23993);
nand U24142 (N_24142,N_23787,N_23935);
xor U24143 (N_24143,N_23640,N_23729);
or U24144 (N_24144,N_23948,N_23884);
nor U24145 (N_24145,N_23685,N_23501);
nor U24146 (N_24146,N_23911,N_23985);
or U24147 (N_24147,N_23805,N_23662);
nand U24148 (N_24148,N_23781,N_23879);
nor U24149 (N_24149,N_23565,N_23946);
or U24150 (N_24150,N_23509,N_23975);
nand U24151 (N_24151,N_23702,N_23766);
nor U24152 (N_24152,N_23974,N_23521);
and U24153 (N_24153,N_23624,N_23713);
nor U24154 (N_24154,N_23560,N_23909);
nor U24155 (N_24155,N_23672,N_23554);
and U24156 (N_24156,N_23748,N_23710);
nand U24157 (N_24157,N_23734,N_23669);
and U24158 (N_24158,N_23776,N_23905);
nand U24159 (N_24159,N_23760,N_23543);
or U24160 (N_24160,N_23563,N_23597);
nor U24161 (N_24161,N_23584,N_23851);
and U24162 (N_24162,N_23966,N_23759);
nand U24163 (N_24163,N_23896,N_23950);
nor U24164 (N_24164,N_23534,N_23941);
xnor U24165 (N_24165,N_23721,N_23632);
nand U24166 (N_24166,N_23507,N_23587);
and U24167 (N_24167,N_23912,N_23773);
or U24168 (N_24168,N_23863,N_23876);
nor U24169 (N_24169,N_23529,N_23569);
and U24170 (N_24170,N_23740,N_23988);
xor U24171 (N_24171,N_23619,N_23701);
or U24172 (N_24172,N_23915,N_23885);
or U24173 (N_24173,N_23920,N_23762);
and U24174 (N_24174,N_23519,N_23522);
nor U24175 (N_24175,N_23960,N_23585);
or U24176 (N_24176,N_23500,N_23767);
nand U24177 (N_24177,N_23846,N_23778);
and U24178 (N_24178,N_23989,N_23686);
nand U24179 (N_24179,N_23742,N_23795);
nor U24180 (N_24180,N_23670,N_23770);
xnor U24181 (N_24181,N_23788,N_23574);
xor U24182 (N_24182,N_23663,N_23999);
nand U24183 (N_24183,N_23599,N_23708);
nor U24184 (N_24184,N_23756,N_23825);
and U24185 (N_24185,N_23638,N_23883);
nand U24186 (N_24186,N_23679,N_23706);
or U24187 (N_24187,N_23774,N_23786);
xor U24188 (N_24188,N_23900,N_23850);
or U24189 (N_24189,N_23845,N_23869);
xor U24190 (N_24190,N_23800,N_23873);
nor U24191 (N_24191,N_23832,N_23518);
xor U24192 (N_24192,N_23678,N_23511);
nor U24193 (N_24193,N_23682,N_23754);
nand U24194 (N_24194,N_23907,N_23780);
or U24195 (N_24195,N_23514,N_23606);
and U24196 (N_24196,N_23981,N_23741);
or U24197 (N_24197,N_23520,N_23815);
nor U24198 (N_24198,N_23736,N_23857);
xnor U24199 (N_24199,N_23810,N_23712);
and U24200 (N_24200,N_23675,N_23793);
xnor U24201 (N_24201,N_23581,N_23971);
nor U24202 (N_24202,N_23595,N_23726);
nor U24203 (N_24203,N_23724,N_23844);
and U24204 (N_24204,N_23703,N_23995);
xnor U24205 (N_24205,N_23723,N_23674);
nor U24206 (N_24206,N_23691,N_23976);
or U24207 (N_24207,N_23623,N_23512);
nor U24208 (N_24208,N_23860,N_23928);
nor U24209 (N_24209,N_23761,N_23744);
nor U24210 (N_24210,N_23506,N_23867);
or U24211 (N_24211,N_23819,N_23537);
nand U24212 (N_24212,N_23874,N_23502);
xor U24213 (N_24213,N_23660,N_23893);
nor U24214 (N_24214,N_23571,N_23923);
or U24215 (N_24215,N_23791,N_23656);
nand U24216 (N_24216,N_23856,N_23622);
and U24217 (N_24217,N_23536,N_23553);
nor U24218 (N_24218,N_23652,N_23555);
or U24219 (N_24219,N_23969,N_23515);
and U24220 (N_24220,N_23625,N_23583);
or U24221 (N_24221,N_23607,N_23709);
nor U24222 (N_24222,N_23796,N_23648);
or U24223 (N_24223,N_23964,N_23634);
xor U24224 (N_24224,N_23934,N_23539);
and U24225 (N_24225,N_23626,N_23871);
or U24226 (N_24226,N_23727,N_23673);
nor U24227 (N_24227,N_23949,N_23627);
nor U24228 (N_24228,N_23552,N_23644);
and U24229 (N_24229,N_23745,N_23986);
or U24230 (N_24230,N_23654,N_23962);
nand U24231 (N_24231,N_23641,N_23549);
and U24232 (N_24232,N_23614,N_23906);
nor U24233 (N_24233,N_23882,N_23811);
and U24234 (N_24234,N_23977,N_23794);
xor U24235 (N_24235,N_23952,N_23692);
and U24236 (N_24236,N_23550,N_23600);
and U24237 (N_24237,N_23852,N_23510);
nor U24238 (N_24238,N_23664,N_23808);
xnor U24239 (N_24239,N_23568,N_23998);
xor U24240 (N_24240,N_23775,N_23961);
and U24241 (N_24241,N_23956,N_23609);
nand U24242 (N_24242,N_23667,N_23594);
xor U24243 (N_24243,N_23677,N_23615);
and U24244 (N_24244,N_23945,N_23939);
xor U24245 (N_24245,N_23659,N_23649);
xor U24246 (N_24246,N_23777,N_23628);
nor U24247 (N_24247,N_23859,N_23749);
and U24248 (N_24248,N_23570,N_23683);
xnor U24249 (N_24249,N_23965,N_23877);
and U24250 (N_24250,N_23596,N_23901);
nor U24251 (N_24251,N_23907,N_23648);
and U24252 (N_24252,N_23926,N_23963);
nand U24253 (N_24253,N_23973,N_23545);
or U24254 (N_24254,N_23860,N_23693);
and U24255 (N_24255,N_23878,N_23563);
and U24256 (N_24256,N_23949,N_23823);
and U24257 (N_24257,N_23844,N_23597);
and U24258 (N_24258,N_23616,N_23580);
and U24259 (N_24259,N_23754,N_23695);
or U24260 (N_24260,N_23591,N_23535);
nor U24261 (N_24261,N_23809,N_23870);
nor U24262 (N_24262,N_23927,N_23525);
and U24263 (N_24263,N_23875,N_23605);
nor U24264 (N_24264,N_23649,N_23823);
nand U24265 (N_24265,N_23632,N_23616);
or U24266 (N_24266,N_23957,N_23613);
and U24267 (N_24267,N_23703,N_23743);
xnor U24268 (N_24268,N_23560,N_23636);
and U24269 (N_24269,N_23937,N_23795);
or U24270 (N_24270,N_23868,N_23720);
or U24271 (N_24271,N_23945,N_23953);
xnor U24272 (N_24272,N_23649,N_23859);
and U24273 (N_24273,N_23741,N_23811);
or U24274 (N_24274,N_23699,N_23871);
nand U24275 (N_24275,N_23988,N_23841);
xor U24276 (N_24276,N_23859,N_23514);
nand U24277 (N_24277,N_23641,N_23637);
or U24278 (N_24278,N_23617,N_23792);
nor U24279 (N_24279,N_23836,N_23698);
or U24280 (N_24280,N_23654,N_23971);
nand U24281 (N_24281,N_23941,N_23740);
xnor U24282 (N_24282,N_23710,N_23892);
nand U24283 (N_24283,N_23969,N_23596);
and U24284 (N_24284,N_23602,N_23659);
nor U24285 (N_24285,N_23663,N_23608);
or U24286 (N_24286,N_23644,N_23669);
nand U24287 (N_24287,N_23707,N_23513);
or U24288 (N_24288,N_23918,N_23580);
xnor U24289 (N_24289,N_23506,N_23792);
xor U24290 (N_24290,N_23951,N_23728);
or U24291 (N_24291,N_23741,N_23947);
nand U24292 (N_24292,N_23622,N_23987);
nor U24293 (N_24293,N_23588,N_23953);
or U24294 (N_24294,N_23616,N_23950);
and U24295 (N_24295,N_23976,N_23562);
nor U24296 (N_24296,N_23683,N_23798);
and U24297 (N_24297,N_23749,N_23533);
nand U24298 (N_24298,N_23628,N_23570);
xnor U24299 (N_24299,N_23922,N_23609);
or U24300 (N_24300,N_23565,N_23776);
and U24301 (N_24301,N_23780,N_23937);
and U24302 (N_24302,N_23568,N_23831);
xor U24303 (N_24303,N_23548,N_23784);
nand U24304 (N_24304,N_23551,N_23844);
nand U24305 (N_24305,N_23906,N_23687);
or U24306 (N_24306,N_23837,N_23603);
or U24307 (N_24307,N_23778,N_23987);
and U24308 (N_24308,N_23807,N_23819);
or U24309 (N_24309,N_23898,N_23929);
xor U24310 (N_24310,N_23587,N_23592);
nand U24311 (N_24311,N_23758,N_23643);
xor U24312 (N_24312,N_23736,N_23522);
nor U24313 (N_24313,N_23855,N_23792);
and U24314 (N_24314,N_23782,N_23688);
nand U24315 (N_24315,N_23969,N_23501);
xor U24316 (N_24316,N_23525,N_23832);
and U24317 (N_24317,N_23688,N_23521);
and U24318 (N_24318,N_23539,N_23859);
nor U24319 (N_24319,N_23593,N_23811);
nand U24320 (N_24320,N_23550,N_23899);
or U24321 (N_24321,N_23571,N_23784);
and U24322 (N_24322,N_23992,N_23970);
xnor U24323 (N_24323,N_23909,N_23758);
and U24324 (N_24324,N_23572,N_23845);
and U24325 (N_24325,N_23970,N_23543);
and U24326 (N_24326,N_23673,N_23639);
and U24327 (N_24327,N_23815,N_23860);
or U24328 (N_24328,N_23586,N_23911);
and U24329 (N_24329,N_23908,N_23978);
xnor U24330 (N_24330,N_23928,N_23743);
nor U24331 (N_24331,N_23578,N_23568);
xor U24332 (N_24332,N_23672,N_23757);
nor U24333 (N_24333,N_23540,N_23803);
or U24334 (N_24334,N_23668,N_23699);
or U24335 (N_24335,N_23725,N_23580);
xnor U24336 (N_24336,N_23675,N_23766);
and U24337 (N_24337,N_23906,N_23661);
nand U24338 (N_24338,N_23590,N_23906);
or U24339 (N_24339,N_23843,N_23824);
xnor U24340 (N_24340,N_23720,N_23555);
xor U24341 (N_24341,N_23618,N_23619);
or U24342 (N_24342,N_23592,N_23646);
nand U24343 (N_24343,N_23726,N_23746);
and U24344 (N_24344,N_23640,N_23926);
and U24345 (N_24345,N_23624,N_23684);
xor U24346 (N_24346,N_23820,N_23729);
and U24347 (N_24347,N_23578,N_23536);
and U24348 (N_24348,N_23586,N_23632);
and U24349 (N_24349,N_23727,N_23835);
xor U24350 (N_24350,N_23855,N_23546);
nor U24351 (N_24351,N_23711,N_23848);
and U24352 (N_24352,N_23980,N_23809);
or U24353 (N_24353,N_23935,N_23659);
and U24354 (N_24354,N_23702,N_23877);
nand U24355 (N_24355,N_23605,N_23888);
nor U24356 (N_24356,N_23518,N_23658);
nor U24357 (N_24357,N_23565,N_23799);
nand U24358 (N_24358,N_23979,N_23711);
xnor U24359 (N_24359,N_23908,N_23648);
or U24360 (N_24360,N_23573,N_23602);
nand U24361 (N_24361,N_23509,N_23638);
or U24362 (N_24362,N_23632,N_23857);
and U24363 (N_24363,N_23898,N_23741);
or U24364 (N_24364,N_23785,N_23969);
or U24365 (N_24365,N_23594,N_23976);
xor U24366 (N_24366,N_23711,N_23967);
and U24367 (N_24367,N_23615,N_23624);
nand U24368 (N_24368,N_23827,N_23697);
or U24369 (N_24369,N_23816,N_23527);
xnor U24370 (N_24370,N_23616,N_23943);
and U24371 (N_24371,N_23692,N_23792);
and U24372 (N_24372,N_23540,N_23872);
and U24373 (N_24373,N_23675,N_23960);
and U24374 (N_24374,N_23690,N_23956);
and U24375 (N_24375,N_23773,N_23668);
and U24376 (N_24376,N_23623,N_23689);
and U24377 (N_24377,N_23609,N_23504);
and U24378 (N_24378,N_23934,N_23758);
xor U24379 (N_24379,N_23831,N_23796);
xor U24380 (N_24380,N_23940,N_23774);
or U24381 (N_24381,N_23904,N_23917);
nand U24382 (N_24382,N_23696,N_23651);
or U24383 (N_24383,N_23846,N_23537);
and U24384 (N_24384,N_23687,N_23741);
and U24385 (N_24385,N_23697,N_23680);
and U24386 (N_24386,N_23809,N_23869);
nand U24387 (N_24387,N_23733,N_23781);
xnor U24388 (N_24388,N_23631,N_23898);
and U24389 (N_24389,N_23995,N_23813);
nor U24390 (N_24390,N_23888,N_23856);
xnor U24391 (N_24391,N_23691,N_23953);
nand U24392 (N_24392,N_23602,N_23835);
or U24393 (N_24393,N_23881,N_23912);
or U24394 (N_24394,N_23990,N_23996);
xor U24395 (N_24395,N_23755,N_23840);
xnor U24396 (N_24396,N_23695,N_23744);
and U24397 (N_24397,N_23709,N_23860);
nor U24398 (N_24398,N_23997,N_23609);
xor U24399 (N_24399,N_23523,N_23635);
nand U24400 (N_24400,N_23718,N_23641);
or U24401 (N_24401,N_23650,N_23630);
xnor U24402 (N_24402,N_23755,N_23631);
nand U24403 (N_24403,N_23524,N_23521);
and U24404 (N_24404,N_23660,N_23705);
and U24405 (N_24405,N_23679,N_23506);
and U24406 (N_24406,N_23600,N_23761);
nor U24407 (N_24407,N_23667,N_23748);
xnor U24408 (N_24408,N_23686,N_23864);
xor U24409 (N_24409,N_23746,N_23817);
nor U24410 (N_24410,N_23658,N_23502);
xnor U24411 (N_24411,N_23723,N_23804);
nor U24412 (N_24412,N_23727,N_23593);
nand U24413 (N_24413,N_23814,N_23742);
or U24414 (N_24414,N_23914,N_23740);
xnor U24415 (N_24415,N_23881,N_23908);
nor U24416 (N_24416,N_23714,N_23772);
nor U24417 (N_24417,N_23657,N_23855);
nor U24418 (N_24418,N_23726,N_23897);
xnor U24419 (N_24419,N_23629,N_23644);
or U24420 (N_24420,N_23937,N_23547);
nor U24421 (N_24421,N_23846,N_23856);
nand U24422 (N_24422,N_23689,N_23727);
nor U24423 (N_24423,N_23735,N_23579);
nand U24424 (N_24424,N_23874,N_23536);
or U24425 (N_24425,N_23752,N_23679);
or U24426 (N_24426,N_23611,N_23701);
and U24427 (N_24427,N_23735,N_23662);
or U24428 (N_24428,N_23940,N_23532);
nor U24429 (N_24429,N_23832,N_23593);
nor U24430 (N_24430,N_23826,N_23622);
and U24431 (N_24431,N_23681,N_23876);
nand U24432 (N_24432,N_23862,N_23964);
or U24433 (N_24433,N_23898,N_23671);
nand U24434 (N_24434,N_23975,N_23630);
xnor U24435 (N_24435,N_23511,N_23818);
xor U24436 (N_24436,N_23945,N_23638);
or U24437 (N_24437,N_23661,N_23910);
xor U24438 (N_24438,N_23771,N_23947);
nand U24439 (N_24439,N_23564,N_23599);
nor U24440 (N_24440,N_23698,N_23768);
and U24441 (N_24441,N_23534,N_23993);
xnor U24442 (N_24442,N_23966,N_23583);
nand U24443 (N_24443,N_23776,N_23855);
nand U24444 (N_24444,N_23899,N_23999);
nand U24445 (N_24445,N_23879,N_23906);
xnor U24446 (N_24446,N_23570,N_23836);
or U24447 (N_24447,N_23934,N_23760);
or U24448 (N_24448,N_23501,N_23547);
nand U24449 (N_24449,N_23980,N_23648);
and U24450 (N_24450,N_23726,N_23904);
nand U24451 (N_24451,N_23887,N_23601);
nor U24452 (N_24452,N_23827,N_23869);
and U24453 (N_24453,N_23720,N_23707);
or U24454 (N_24454,N_23658,N_23597);
nor U24455 (N_24455,N_23589,N_23996);
nand U24456 (N_24456,N_23946,N_23535);
xor U24457 (N_24457,N_23991,N_23855);
and U24458 (N_24458,N_23777,N_23929);
or U24459 (N_24459,N_23705,N_23561);
and U24460 (N_24460,N_23541,N_23898);
xnor U24461 (N_24461,N_23721,N_23742);
or U24462 (N_24462,N_23961,N_23634);
xnor U24463 (N_24463,N_23721,N_23627);
or U24464 (N_24464,N_23798,N_23960);
or U24465 (N_24465,N_23961,N_23647);
nor U24466 (N_24466,N_23930,N_23858);
and U24467 (N_24467,N_23824,N_23651);
xnor U24468 (N_24468,N_23577,N_23756);
xor U24469 (N_24469,N_23840,N_23772);
nand U24470 (N_24470,N_23825,N_23974);
nand U24471 (N_24471,N_23869,N_23992);
nor U24472 (N_24472,N_23750,N_23619);
or U24473 (N_24473,N_23577,N_23568);
nor U24474 (N_24474,N_23574,N_23590);
nor U24475 (N_24475,N_23650,N_23786);
nor U24476 (N_24476,N_23968,N_23687);
or U24477 (N_24477,N_23754,N_23926);
and U24478 (N_24478,N_23761,N_23584);
and U24479 (N_24479,N_23887,N_23730);
xnor U24480 (N_24480,N_23888,N_23947);
and U24481 (N_24481,N_23834,N_23742);
nand U24482 (N_24482,N_23536,N_23934);
nand U24483 (N_24483,N_23503,N_23898);
xnor U24484 (N_24484,N_23743,N_23722);
xnor U24485 (N_24485,N_23609,N_23674);
nor U24486 (N_24486,N_23729,N_23839);
nand U24487 (N_24487,N_23519,N_23740);
nand U24488 (N_24488,N_23656,N_23553);
or U24489 (N_24489,N_23985,N_23776);
xnor U24490 (N_24490,N_23994,N_23558);
xor U24491 (N_24491,N_23641,N_23719);
nor U24492 (N_24492,N_23515,N_23569);
and U24493 (N_24493,N_23905,N_23762);
xnor U24494 (N_24494,N_23765,N_23645);
nor U24495 (N_24495,N_23743,N_23584);
and U24496 (N_24496,N_23767,N_23513);
nand U24497 (N_24497,N_23974,N_23776);
nand U24498 (N_24498,N_23610,N_23750);
and U24499 (N_24499,N_23683,N_23611);
nor U24500 (N_24500,N_24328,N_24408);
xor U24501 (N_24501,N_24324,N_24020);
and U24502 (N_24502,N_24225,N_24430);
or U24503 (N_24503,N_24148,N_24068);
xnor U24504 (N_24504,N_24144,N_24235);
xor U24505 (N_24505,N_24478,N_24207);
nand U24506 (N_24506,N_24186,N_24047);
or U24507 (N_24507,N_24042,N_24264);
or U24508 (N_24508,N_24142,N_24476);
xor U24509 (N_24509,N_24256,N_24385);
nor U24510 (N_24510,N_24445,N_24287);
xnor U24511 (N_24511,N_24062,N_24475);
or U24512 (N_24512,N_24325,N_24352);
nor U24513 (N_24513,N_24080,N_24432);
xor U24514 (N_24514,N_24409,N_24064);
and U24515 (N_24515,N_24129,N_24340);
nor U24516 (N_24516,N_24234,N_24279);
xnor U24517 (N_24517,N_24053,N_24184);
xnor U24518 (N_24518,N_24003,N_24447);
or U24519 (N_24519,N_24307,N_24378);
nand U24520 (N_24520,N_24260,N_24030);
and U24521 (N_24521,N_24451,N_24433);
or U24522 (N_24522,N_24078,N_24212);
nor U24523 (N_24523,N_24336,N_24175);
or U24524 (N_24524,N_24092,N_24002);
and U24525 (N_24525,N_24190,N_24061);
nor U24526 (N_24526,N_24481,N_24288);
nand U24527 (N_24527,N_24330,N_24227);
and U24528 (N_24528,N_24077,N_24115);
and U24529 (N_24529,N_24365,N_24166);
and U24530 (N_24530,N_24008,N_24405);
and U24531 (N_24531,N_24333,N_24320);
nand U24532 (N_24532,N_24254,N_24195);
nor U24533 (N_24533,N_24347,N_24209);
or U24534 (N_24534,N_24130,N_24236);
or U24535 (N_24535,N_24420,N_24419);
and U24536 (N_24536,N_24259,N_24073);
or U24537 (N_24537,N_24194,N_24048);
or U24538 (N_24538,N_24238,N_24012);
nor U24539 (N_24539,N_24453,N_24263);
xor U24540 (N_24540,N_24458,N_24007);
and U24541 (N_24541,N_24470,N_24120);
nand U24542 (N_24542,N_24465,N_24389);
xor U24543 (N_24543,N_24494,N_24442);
xnor U24544 (N_24544,N_24444,N_24271);
or U24545 (N_24545,N_24170,N_24362);
and U24546 (N_24546,N_24449,N_24055);
nand U24547 (N_24547,N_24486,N_24049);
nand U24548 (N_24548,N_24329,N_24474);
and U24549 (N_24549,N_24150,N_24122);
nand U24550 (N_24550,N_24317,N_24377);
and U24551 (N_24551,N_24063,N_24398);
or U24552 (N_24552,N_24344,N_24106);
xor U24553 (N_24553,N_24276,N_24498);
or U24554 (N_24554,N_24174,N_24431);
nand U24555 (N_24555,N_24114,N_24381);
xor U24556 (N_24556,N_24233,N_24286);
nor U24557 (N_24557,N_24125,N_24318);
nor U24558 (N_24558,N_24487,N_24483);
and U24559 (N_24559,N_24229,N_24066);
nand U24560 (N_24560,N_24240,N_24350);
xor U24561 (N_24561,N_24023,N_24164);
nor U24562 (N_24562,N_24069,N_24363);
nand U24563 (N_24563,N_24090,N_24121);
nand U24564 (N_24564,N_24479,N_24272);
or U24565 (N_24565,N_24079,N_24436);
xor U24566 (N_24566,N_24414,N_24163);
nor U24567 (N_24567,N_24282,N_24089);
xnor U24568 (N_24568,N_24241,N_24201);
nor U24569 (N_24569,N_24216,N_24117);
nor U24570 (N_24570,N_24057,N_24313);
nor U24571 (N_24571,N_24252,N_24428);
and U24572 (N_24572,N_24327,N_24232);
xnor U24573 (N_24573,N_24133,N_24348);
xnor U24574 (N_24574,N_24422,N_24167);
nand U24575 (N_24575,N_24031,N_24218);
or U24576 (N_24576,N_24192,N_24308);
or U24577 (N_24577,N_24116,N_24492);
nand U24578 (N_24578,N_24197,N_24354);
and U24579 (N_24579,N_24102,N_24024);
and U24580 (N_24580,N_24322,N_24208);
nor U24581 (N_24581,N_24056,N_24305);
or U24582 (N_24582,N_24037,N_24403);
and U24583 (N_24583,N_24257,N_24132);
nand U24584 (N_24584,N_24391,N_24342);
xor U24585 (N_24585,N_24370,N_24438);
or U24586 (N_24586,N_24247,N_24179);
nand U24587 (N_24587,N_24112,N_24338);
nand U24588 (N_24588,N_24085,N_24104);
and U24589 (N_24589,N_24110,N_24400);
nor U24590 (N_24590,N_24154,N_24346);
nand U24591 (N_24591,N_24375,N_24119);
and U24592 (N_24592,N_24022,N_24267);
xor U24593 (N_24593,N_24001,N_24337);
nor U24594 (N_24594,N_24395,N_24332);
nor U24595 (N_24595,N_24415,N_24147);
nor U24596 (N_24596,N_24457,N_24095);
nand U24597 (N_24597,N_24183,N_24484);
nand U24598 (N_24598,N_24326,N_24178);
xnor U24599 (N_24599,N_24343,N_24000);
and U24600 (N_24600,N_24357,N_24032);
or U24601 (N_24601,N_24151,N_24364);
nand U24602 (N_24602,N_24171,N_24412);
nand U24603 (N_24603,N_24226,N_24406);
or U24604 (N_24604,N_24118,N_24416);
xnor U24605 (N_24605,N_24137,N_24250);
and U24606 (N_24606,N_24262,N_24138);
xor U24607 (N_24607,N_24456,N_24189);
nand U24608 (N_24608,N_24244,N_24108);
nand U24609 (N_24609,N_24488,N_24152);
nand U24610 (N_24610,N_24221,N_24161);
and U24611 (N_24611,N_24081,N_24316);
nand U24612 (N_24612,N_24499,N_24071);
nand U24613 (N_24613,N_24345,N_24396);
and U24614 (N_24614,N_24156,N_24141);
nor U24615 (N_24615,N_24295,N_24127);
xnor U24616 (N_24616,N_24176,N_24004);
nor U24617 (N_24617,N_24452,N_24160);
nor U24618 (N_24618,N_24390,N_24467);
and U24619 (N_24619,N_24297,N_24426);
or U24620 (N_24620,N_24304,N_24018);
and U24621 (N_24621,N_24205,N_24468);
or U24622 (N_24622,N_24029,N_24113);
and U24623 (N_24623,N_24311,N_24392);
or U24624 (N_24624,N_24482,N_24014);
nand U24625 (N_24625,N_24334,N_24314);
and U24626 (N_24626,N_24045,N_24265);
or U24627 (N_24627,N_24315,N_24097);
nor U24628 (N_24628,N_24427,N_24477);
and U24629 (N_24629,N_24341,N_24070);
or U24630 (N_24630,N_24067,N_24107);
nand U24631 (N_24631,N_24373,N_24228);
xnor U24632 (N_24632,N_24075,N_24182);
nand U24633 (N_24633,N_24302,N_24083);
and U24634 (N_24634,N_24323,N_24196);
nor U24635 (N_24635,N_24054,N_24177);
and U24636 (N_24636,N_24051,N_24367);
or U24637 (N_24637,N_24006,N_24242);
and U24638 (N_24638,N_24251,N_24417);
xor U24639 (N_24639,N_24215,N_24038);
nand U24640 (N_24640,N_24084,N_24497);
nor U24641 (N_24641,N_24010,N_24404);
nor U24642 (N_24642,N_24036,N_24026);
xnor U24643 (N_24643,N_24394,N_24128);
or U24644 (N_24644,N_24027,N_24383);
nor U24645 (N_24645,N_24371,N_24096);
or U24646 (N_24646,N_24149,N_24423);
xor U24647 (N_24647,N_24335,N_24019);
and U24648 (N_24648,N_24123,N_24319);
nor U24649 (N_24649,N_24039,N_24299);
nand U24650 (N_24650,N_24139,N_24169);
xor U24651 (N_24651,N_24243,N_24380);
or U24652 (N_24652,N_24076,N_24015);
xnor U24653 (N_24653,N_24165,N_24294);
or U24654 (N_24654,N_24065,N_24495);
nand U24655 (N_24655,N_24253,N_24270);
or U24656 (N_24656,N_24283,N_24249);
nand U24657 (N_24657,N_24025,N_24155);
or U24658 (N_24658,N_24134,N_24440);
nor U24659 (N_24659,N_24044,N_24017);
nor U24660 (N_24660,N_24289,N_24368);
and U24661 (N_24661,N_24086,N_24005);
nand U24662 (N_24662,N_24258,N_24493);
or U24663 (N_24663,N_24473,N_24437);
xor U24664 (N_24664,N_24421,N_24074);
nor U24665 (N_24665,N_24459,N_24248);
or U24666 (N_24666,N_24162,N_24461);
and U24667 (N_24667,N_24496,N_24399);
and U24668 (N_24668,N_24094,N_24101);
and U24669 (N_24669,N_24360,N_24187);
xnor U24670 (N_24670,N_24050,N_24463);
nor U24671 (N_24671,N_24376,N_24193);
xor U24672 (N_24672,N_24091,N_24131);
or U24673 (N_24673,N_24281,N_24200);
and U24674 (N_24674,N_24448,N_24093);
nand U24675 (N_24675,N_24231,N_24312);
or U24676 (N_24676,N_24213,N_24266);
xor U24677 (N_24677,N_24016,N_24491);
nand U24678 (N_24678,N_24041,N_24220);
nand U24679 (N_24679,N_24035,N_24136);
nand U24680 (N_24680,N_24278,N_24387);
nand U24681 (N_24681,N_24339,N_24046);
nand U24682 (N_24682,N_24157,N_24361);
xnor U24683 (N_24683,N_24306,N_24273);
nand U24684 (N_24684,N_24489,N_24309);
and U24685 (N_24685,N_24425,N_24393);
and U24686 (N_24686,N_24296,N_24100);
and U24687 (N_24687,N_24087,N_24210);
xnor U24688 (N_24688,N_24105,N_24028);
or U24689 (N_24689,N_24413,N_24202);
and U24690 (N_24690,N_24379,N_24124);
or U24691 (N_24691,N_24203,N_24058);
and U24692 (N_24692,N_24460,N_24172);
xnor U24693 (N_24693,N_24211,N_24464);
xnor U24694 (N_24694,N_24454,N_24462);
or U24695 (N_24695,N_24407,N_24135);
and U24696 (N_24696,N_24145,N_24274);
or U24697 (N_24697,N_24011,N_24198);
or U24698 (N_24698,N_24206,N_24374);
nand U24699 (N_24699,N_24034,N_24386);
or U24700 (N_24700,N_24280,N_24052);
or U24701 (N_24701,N_24181,N_24300);
nor U24702 (N_24702,N_24410,N_24217);
xnor U24703 (N_24703,N_24103,N_24298);
xor U24704 (N_24704,N_24140,N_24111);
xor U24705 (N_24705,N_24446,N_24275);
nand U24706 (N_24706,N_24043,N_24472);
or U24707 (N_24707,N_24237,N_24366);
nand U24708 (N_24708,N_24480,N_24222);
xnor U24709 (N_24709,N_24099,N_24098);
nand U24710 (N_24710,N_24033,N_24388);
nor U24711 (N_24711,N_24369,N_24424);
xor U24712 (N_24712,N_24013,N_24418);
or U24713 (N_24713,N_24469,N_24301);
and U24714 (N_24714,N_24466,N_24261);
nor U24715 (N_24715,N_24402,N_24355);
and U24716 (N_24716,N_24450,N_24292);
nor U24717 (N_24717,N_24159,N_24358);
and U24718 (N_24718,N_24223,N_24321);
xor U24719 (N_24719,N_24291,N_24021);
xor U24720 (N_24720,N_24191,N_24285);
and U24721 (N_24721,N_24382,N_24303);
nand U24722 (N_24722,N_24401,N_24429);
nor U24723 (N_24723,N_24219,N_24353);
xor U24724 (N_24724,N_24310,N_24351);
nor U24725 (N_24725,N_24397,N_24143);
nand U24726 (N_24726,N_24255,N_24441);
nor U24727 (N_24727,N_24146,N_24214);
nand U24728 (N_24728,N_24331,N_24173);
xor U24729 (N_24729,N_24372,N_24435);
nand U24730 (N_24730,N_24434,N_24060);
nand U24731 (N_24731,N_24204,N_24239);
and U24732 (N_24732,N_24040,N_24439);
and U24733 (N_24733,N_24199,N_24471);
nor U24734 (N_24734,N_24293,N_24168);
xnor U24735 (N_24735,N_24185,N_24158);
xnor U24736 (N_24736,N_24109,N_24268);
nor U24737 (N_24737,N_24284,N_24072);
nor U24738 (N_24738,N_24277,N_24126);
nor U24739 (N_24739,N_24443,N_24455);
xor U24740 (N_24740,N_24009,N_24384);
nand U24741 (N_24741,N_24153,N_24290);
xor U24742 (N_24742,N_24180,N_24490);
nand U24743 (N_24743,N_24059,N_24224);
xor U24744 (N_24744,N_24245,N_24088);
or U24745 (N_24745,N_24356,N_24411);
nand U24746 (N_24746,N_24230,N_24188);
nor U24747 (N_24747,N_24349,N_24485);
and U24748 (N_24748,N_24246,N_24359);
nand U24749 (N_24749,N_24269,N_24082);
and U24750 (N_24750,N_24427,N_24066);
or U24751 (N_24751,N_24286,N_24253);
xnor U24752 (N_24752,N_24102,N_24463);
and U24753 (N_24753,N_24136,N_24075);
xnor U24754 (N_24754,N_24094,N_24450);
nor U24755 (N_24755,N_24096,N_24323);
or U24756 (N_24756,N_24011,N_24123);
xor U24757 (N_24757,N_24097,N_24395);
nor U24758 (N_24758,N_24458,N_24093);
nand U24759 (N_24759,N_24121,N_24044);
nand U24760 (N_24760,N_24364,N_24490);
nand U24761 (N_24761,N_24248,N_24422);
and U24762 (N_24762,N_24065,N_24398);
or U24763 (N_24763,N_24229,N_24301);
xnor U24764 (N_24764,N_24200,N_24046);
nor U24765 (N_24765,N_24496,N_24435);
nand U24766 (N_24766,N_24209,N_24334);
nor U24767 (N_24767,N_24096,N_24289);
or U24768 (N_24768,N_24157,N_24420);
nand U24769 (N_24769,N_24136,N_24271);
xor U24770 (N_24770,N_24433,N_24106);
and U24771 (N_24771,N_24370,N_24363);
nand U24772 (N_24772,N_24047,N_24147);
nand U24773 (N_24773,N_24352,N_24356);
and U24774 (N_24774,N_24236,N_24248);
nor U24775 (N_24775,N_24329,N_24223);
or U24776 (N_24776,N_24005,N_24195);
nor U24777 (N_24777,N_24261,N_24142);
nor U24778 (N_24778,N_24111,N_24010);
or U24779 (N_24779,N_24006,N_24463);
nor U24780 (N_24780,N_24399,N_24485);
xnor U24781 (N_24781,N_24269,N_24384);
xnor U24782 (N_24782,N_24145,N_24480);
or U24783 (N_24783,N_24156,N_24329);
nand U24784 (N_24784,N_24061,N_24477);
nor U24785 (N_24785,N_24321,N_24094);
nand U24786 (N_24786,N_24383,N_24231);
nor U24787 (N_24787,N_24428,N_24082);
xnor U24788 (N_24788,N_24253,N_24384);
or U24789 (N_24789,N_24060,N_24183);
and U24790 (N_24790,N_24022,N_24428);
or U24791 (N_24791,N_24113,N_24117);
nor U24792 (N_24792,N_24233,N_24005);
nand U24793 (N_24793,N_24461,N_24414);
nor U24794 (N_24794,N_24230,N_24063);
nor U24795 (N_24795,N_24214,N_24430);
and U24796 (N_24796,N_24226,N_24035);
or U24797 (N_24797,N_24099,N_24411);
and U24798 (N_24798,N_24469,N_24212);
or U24799 (N_24799,N_24358,N_24483);
nand U24800 (N_24800,N_24353,N_24212);
xor U24801 (N_24801,N_24156,N_24359);
or U24802 (N_24802,N_24464,N_24234);
nor U24803 (N_24803,N_24397,N_24200);
nor U24804 (N_24804,N_24129,N_24342);
xnor U24805 (N_24805,N_24212,N_24499);
and U24806 (N_24806,N_24486,N_24479);
xnor U24807 (N_24807,N_24360,N_24007);
nor U24808 (N_24808,N_24461,N_24294);
and U24809 (N_24809,N_24357,N_24170);
nand U24810 (N_24810,N_24302,N_24289);
and U24811 (N_24811,N_24178,N_24093);
nand U24812 (N_24812,N_24108,N_24046);
or U24813 (N_24813,N_24025,N_24295);
nor U24814 (N_24814,N_24456,N_24012);
nor U24815 (N_24815,N_24268,N_24085);
nor U24816 (N_24816,N_24482,N_24390);
nor U24817 (N_24817,N_24192,N_24126);
and U24818 (N_24818,N_24384,N_24211);
nor U24819 (N_24819,N_24424,N_24381);
nand U24820 (N_24820,N_24227,N_24258);
nand U24821 (N_24821,N_24477,N_24273);
nor U24822 (N_24822,N_24326,N_24484);
or U24823 (N_24823,N_24025,N_24159);
xor U24824 (N_24824,N_24499,N_24317);
xnor U24825 (N_24825,N_24298,N_24309);
or U24826 (N_24826,N_24151,N_24485);
and U24827 (N_24827,N_24484,N_24448);
and U24828 (N_24828,N_24020,N_24255);
nand U24829 (N_24829,N_24365,N_24175);
or U24830 (N_24830,N_24251,N_24135);
or U24831 (N_24831,N_24324,N_24224);
nand U24832 (N_24832,N_24281,N_24063);
and U24833 (N_24833,N_24039,N_24192);
xnor U24834 (N_24834,N_24281,N_24093);
or U24835 (N_24835,N_24216,N_24351);
xor U24836 (N_24836,N_24247,N_24200);
xnor U24837 (N_24837,N_24259,N_24394);
and U24838 (N_24838,N_24375,N_24340);
or U24839 (N_24839,N_24443,N_24299);
and U24840 (N_24840,N_24497,N_24106);
nand U24841 (N_24841,N_24422,N_24467);
xnor U24842 (N_24842,N_24242,N_24447);
nor U24843 (N_24843,N_24399,N_24169);
nand U24844 (N_24844,N_24169,N_24292);
or U24845 (N_24845,N_24374,N_24055);
xor U24846 (N_24846,N_24067,N_24126);
and U24847 (N_24847,N_24311,N_24354);
and U24848 (N_24848,N_24302,N_24250);
and U24849 (N_24849,N_24299,N_24095);
and U24850 (N_24850,N_24328,N_24262);
or U24851 (N_24851,N_24234,N_24445);
nor U24852 (N_24852,N_24454,N_24298);
and U24853 (N_24853,N_24252,N_24455);
nand U24854 (N_24854,N_24208,N_24153);
xnor U24855 (N_24855,N_24195,N_24255);
and U24856 (N_24856,N_24482,N_24059);
nor U24857 (N_24857,N_24443,N_24051);
nand U24858 (N_24858,N_24352,N_24372);
or U24859 (N_24859,N_24408,N_24361);
xor U24860 (N_24860,N_24019,N_24295);
and U24861 (N_24861,N_24070,N_24095);
nor U24862 (N_24862,N_24100,N_24347);
and U24863 (N_24863,N_24433,N_24156);
nand U24864 (N_24864,N_24178,N_24366);
nand U24865 (N_24865,N_24059,N_24403);
nand U24866 (N_24866,N_24200,N_24476);
xor U24867 (N_24867,N_24252,N_24438);
or U24868 (N_24868,N_24221,N_24148);
nor U24869 (N_24869,N_24187,N_24349);
and U24870 (N_24870,N_24404,N_24193);
nand U24871 (N_24871,N_24304,N_24136);
xor U24872 (N_24872,N_24342,N_24387);
nand U24873 (N_24873,N_24269,N_24323);
nand U24874 (N_24874,N_24382,N_24165);
nor U24875 (N_24875,N_24098,N_24109);
xnor U24876 (N_24876,N_24187,N_24182);
and U24877 (N_24877,N_24025,N_24338);
and U24878 (N_24878,N_24464,N_24240);
or U24879 (N_24879,N_24270,N_24296);
nand U24880 (N_24880,N_24015,N_24199);
nor U24881 (N_24881,N_24094,N_24245);
xnor U24882 (N_24882,N_24350,N_24471);
nand U24883 (N_24883,N_24170,N_24484);
nand U24884 (N_24884,N_24430,N_24491);
xor U24885 (N_24885,N_24034,N_24242);
nor U24886 (N_24886,N_24202,N_24118);
or U24887 (N_24887,N_24195,N_24093);
or U24888 (N_24888,N_24462,N_24340);
or U24889 (N_24889,N_24178,N_24261);
and U24890 (N_24890,N_24352,N_24208);
nand U24891 (N_24891,N_24264,N_24005);
and U24892 (N_24892,N_24194,N_24142);
xnor U24893 (N_24893,N_24226,N_24246);
nand U24894 (N_24894,N_24084,N_24275);
and U24895 (N_24895,N_24469,N_24109);
and U24896 (N_24896,N_24022,N_24480);
nor U24897 (N_24897,N_24477,N_24010);
nand U24898 (N_24898,N_24331,N_24289);
or U24899 (N_24899,N_24087,N_24409);
or U24900 (N_24900,N_24245,N_24442);
nand U24901 (N_24901,N_24101,N_24216);
and U24902 (N_24902,N_24164,N_24467);
and U24903 (N_24903,N_24175,N_24204);
nand U24904 (N_24904,N_24143,N_24227);
or U24905 (N_24905,N_24304,N_24457);
nor U24906 (N_24906,N_24444,N_24480);
nor U24907 (N_24907,N_24076,N_24498);
nor U24908 (N_24908,N_24288,N_24282);
and U24909 (N_24909,N_24217,N_24237);
nor U24910 (N_24910,N_24047,N_24219);
nand U24911 (N_24911,N_24118,N_24174);
xnor U24912 (N_24912,N_24070,N_24272);
nand U24913 (N_24913,N_24490,N_24173);
xor U24914 (N_24914,N_24043,N_24463);
or U24915 (N_24915,N_24235,N_24478);
nor U24916 (N_24916,N_24477,N_24171);
xnor U24917 (N_24917,N_24370,N_24392);
xnor U24918 (N_24918,N_24079,N_24477);
and U24919 (N_24919,N_24358,N_24182);
nand U24920 (N_24920,N_24469,N_24026);
nand U24921 (N_24921,N_24169,N_24043);
nand U24922 (N_24922,N_24016,N_24050);
nand U24923 (N_24923,N_24074,N_24214);
nor U24924 (N_24924,N_24276,N_24314);
nor U24925 (N_24925,N_24470,N_24427);
xnor U24926 (N_24926,N_24160,N_24408);
xnor U24927 (N_24927,N_24070,N_24132);
nand U24928 (N_24928,N_24302,N_24148);
or U24929 (N_24929,N_24410,N_24022);
nand U24930 (N_24930,N_24407,N_24323);
and U24931 (N_24931,N_24261,N_24250);
or U24932 (N_24932,N_24421,N_24139);
xor U24933 (N_24933,N_24011,N_24401);
and U24934 (N_24934,N_24133,N_24069);
nand U24935 (N_24935,N_24334,N_24385);
xor U24936 (N_24936,N_24408,N_24474);
xnor U24937 (N_24937,N_24308,N_24110);
xnor U24938 (N_24938,N_24143,N_24045);
xnor U24939 (N_24939,N_24197,N_24298);
and U24940 (N_24940,N_24125,N_24244);
xor U24941 (N_24941,N_24186,N_24017);
and U24942 (N_24942,N_24051,N_24361);
nor U24943 (N_24943,N_24426,N_24100);
xor U24944 (N_24944,N_24350,N_24283);
xor U24945 (N_24945,N_24039,N_24328);
nor U24946 (N_24946,N_24353,N_24021);
or U24947 (N_24947,N_24443,N_24342);
nor U24948 (N_24948,N_24239,N_24126);
xnor U24949 (N_24949,N_24304,N_24372);
and U24950 (N_24950,N_24417,N_24200);
nor U24951 (N_24951,N_24326,N_24240);
or U24952 (N_24952,N_24226,N_24159);
xor U24953 (N_24953,N_24047,N_24189);
nand U24954 (N_24954,N_24419,N_24471);
or U24955 (N_24955,N_24341,N_24499);
nand U24956 (N_24956,N_24391,N_24381);
and U24957 (N_24957,N_24452,N_24306);
or U24958 (N_24958,N_24116,N_24081);
and U24959 (N_24959,N_24290,N_24253);
and U24960 (N_24960,N_24201,N_24050);
and U24961 (N_24961,N_24138,N_24030);
nand U24962 (N_24962,N_24260,N_24136);
nand U24963 (N_24963,N_24233,N_24002);
nand U24964 (N_24964,N_24074,N_24369);
and U24965 (N_24965,N_24139,N_24271);
xnor U24966 (N_24966,N_24283,N_24456);
and U24967 (N_24967,N_24157,N_24477);
and U24968 (N_24968,N_24458,N_24307);
or U24969 (N_24969,N_24155,N_24117);
and U24970 (N_24970,N_24140,N_24307);
and U24971 (N_24971,N_24289,N_24257);
or U24972 (N_24972,N_24299,N_24111);
xor U24973 (N_24973,N_24355,N_24427);
xor U24974 (N_24974,N_24351,N_24421);
or U24975 (N_24975,N_24076,N_24171);
nor U24976 (N_24976,N_24085,N_24495);
or U24977 (N_24977,N_24075,N_24086);
nor U24978 (N_24978,N_24196,N_24183);
and U24979 (N_24979,N_24459,N_24375);
or U24980 (N_24980,N_24246,N_24399);
nor U24981 (N_24981,N_24427,N_24021);
or U24982 (N_24982,N_24000,N_24109);
and U24983 (N_24983,N_24391,N_24497);
and U24984 (N_24984,N_24494,N_24370);
nand U24985 (N_24985,N_24272,N_24155);
or U24986 (N_24986,N_24421,N_24036);
nand U24987 (N_24987,N_24191,N_24338);
nor U24988 (N_24988,N_24045,N_24154);
nand U24989 (N_24989,N_24089,N_24117);
nand U24990 (N_24990,N_24050,N_24021);
nand U24991 (N_24991,N_24283,N_24443);
and U24992 (N_24992,N_24056,N_24271);
nor U24993 (N_24993,N_24295,N_24260);
nor U24994 (N_24994,N_24078,N_24382);
and U24995 (N_24995,N_24096,N_24234);
xor U24996 (N_24996,N_24183,N_24194);
nor U24997 (N_24997,N_24236,N_24371);
or U24998 (N_24998,N_24482,N_24483);
nor U24999 (N_24999,N_24069,N_24344);
and UO_0 (O_0,N_24683,N_24669);
nand UO_1 (O_1,N_24995,N_24779);
and UO_2 (O_2,N_24920,N_24513);
nand UO_3 (O_3,N_24719,N_24908);
nor UO_4 (O_4,N_24838,N_24962);
nand UO_5 (O_5,N_24703,N_24604);
and UO_6 (O_6,N_24944,N_24953);
nor UO_7 (O_7,N_24810,N_24957);
xnor UO_8 (O_8,N_24510,N_24980);
xnor UO_9 (O_9,N_24599,N_24538);
xnor UO_10 (O_10,N_24654,N_24742);
nand UO_11 (O_11,N_24998,N_24682);
or UO_12 (O_12,N_24557,N_24675);
nand UO_13 (O_13,N_24800,N_24859);
nor UO_14 (O_14,N_24961,N_24782);
and UO_15 (O_15,N_24815,N_24596);
xnor UO_16 (O_16,N_24569,N_24680);
nand UO_17 (O_17,N_24631,N_24977);
nor UO_18 (O_18,N_24520,N_24646);
nor UO_19 (O_19,N_24605,N_24902);
xor UO_20 (O_20,N_24664,N_24583);
nand UO_21 (O_21,N_24656,N_24602);
and UO_22 (O_22,N_24935,N_24861);
or UO_23 (O_23,N_24907,N_24526);
nor UO_24 (O_24,N_24891,N_24756);
or UO_25 (O_25,N_24571,N_24919);
nand UO_26 (O_26,N_24796,N_24867);
nor UO_27 (O_27,N_24644,N_24738);
xnor UO_28 (O_28,N_24514,N_24823);
nor UO_29 (O_29,N_24831,N_24572);
xor UO_30 (O_30,N_24870,N_24570);
nor UO_31 (O_31,N_24874,N_24608);
nand UO_32 (O_32,N_24521,N_24876);
xor UO_33 (O_33,N_24610,N_24992);
nand UO_34 (O_34,N_24938,N_24543);
nand UO_35 (O_35,N_24840,N_24777);
xnor UO_36 (O_36,N_24670,N_24626);
nor UO_37 (O_37,N_24746,N_24890);
or UO_38 (O_38,N_24733,N_24798);
and UO_39 (O_39,N_24883,N_24619);
nor UO_40 (O_40,N_24906,N_24630);
or UO_41 (O_41,N_24974,N_24780);
nand UO_42 (O_42,N_24587,N_24533);
nand UO_43 (O_43,N_24614,N_24504);
nand UO_44 (O_44,N_24704,N_24707);
or UO_45 (O_45,N_24681,N_24553);
and UO_46 (O_46,N_24794,N_24633);
nor UO_47 (O_47,N_24639,N_24835);
nor UO_48 (O_48,N_24555,N_24793);
nor UO_49 (O_49,N_24851,N_24624);
or UO_50 (O_50,N_24548,N_24581);
xnor UO_51 (O_51,N_24611,N_24997);
or UO_52 (O_52,N_24546,N_24727);
xnor UO_53 (O_53,N_24667,N_24647);
and UO_54 (O_54,N_24672,N_24556);
or UO_55 (O_55,N_24772,N_24922);
nor UO_56 (O_56,N_24658,N_24858);
nand UO_57 (O_57,N_24714,N_24887);
or UO_58 (O_58,N_24984,N_24685);
and UO_59 (O_59,N_24702,N_24747);
nand UO_60 (O_60,N_24886,N_24894);
or UO_61 (O_61,N_24588,N_24989);
and UO_62 (O_62,N_24807,N_24928);
or UO_63 (O_63,N_24659,N_24885);
nor UO_64 (O_64,N_24817,N_24722);
and UO_65 (O_65,N_24732,N_24561);
nand UO_66 (O_66,N_24735,N_24970);
nand UO_67 (O_67,N_24506,N_24750);
or UO_68 (O_68,N_24763,N_24550);
or UO_69 (O_69,N_24591,N_24927);
nand UO_70 (O_70,N_24509,N_24551);
nor UO_71 (O_71,N_24934,N_24966);
or UO_72 (O_72,N_24806,N_24924);
nor UO_73 (O_73,N_24842,N_24862);
or UO_74 (O_74,N_24687,N_24905);
and UO_75 (O_75,N_24567,N_24503);
nand UO_76 (O_76,N_24893,N_24979);
and UO_77 (O_77,N_24988,N_24712);
and UO_78 (O_78,N_24603,N_24651);
and UO_79 (O_79,N_24617,N_24730);
nor UO_80 (O_80,N_24573,N_24741);
nand UO_81 (O_81,N_24769,N_24845);
and UO_82 (O_82,N_24762,N_24788);
or UO_83 (O_83,N_24837,N_24959);
nand UO_84 (O_84,N_24637,N_24575);
nor UO_85 (O_85,N_24695,N_24697);
and UO_86 (O_86,N_24519,N_24811);
nor UO_87 (O_87,N_24801,N_24868);
and UO_88 (O_88,N_24592,N_24558);
or UO_89 (O_89,N_24776,N_24755);
and UO_90 (O_90,N_24698,N_24700);
xnor UO_91 (O_91,N_24554,N_24530);
nor UO_92 (O_92,N_24715,N_24875);
nand UO_93 (O_93,N_24736,N_24559);
or UO_94 (O_94,N_24650,N_24824);
nand UO_95 (O_95,N_24662,N_24663);
nand UO_96 (O_96,N_24724,N_24694);
and UO_97 (O_97,N_24535,N_24879);
nor UO_98 (O_98,N_24758,N_24812);
or UO_99 (O_99,N_24860,N_24643);
nor UO_100 (O_100,N_24562,N_24737);
and UO_101 (O_101,N_24754,N_24525);
and UO_102 (O_102,N_24954,N_24524);
nand UO_103 (O_103,N_24589,N_24760);
or UO_104 (O_104,N_24889,N_24790);
nand UO_105 (O_105,N_24783,N_24648);
and UO_106 (O_106,N_24690,N_24991);
and UO_107 (O_107,N_24785,N_24795);
nand UO_108 (O_108,N_24729,N_24549);
nand UO_109 (O_109,N_24799,N_24895);
nand UO_110 (O_110,N_24821,N_24999);
and UO_111 (O_111,N_24711,N_24689);
or UO_112 (O_112,N_24500,N_24863);
xnor UO_113 (O_113,N_24918,N_24809);
nor UO_114 (O_114,N_24641,N_24576);
nor UO_115 (O_115,N_24621,N_24940);
xnor UO_116 (O_116,N_24691,N_24540);
xor UO_117 (O_117,N_24882,N_24502);
xnor UO_118 (O_118,N_24964,N_24676);
nand UO_119 (O_119,N_24849,N_24749);
and UO_120 (O_120,N_24774,N_24996);
xor UO_121 (O_121,N_24566,N_24726);
nand UO_122 (O_122,N_24814,N_24518);
xnor UO_123 (O_123,N_24965,N_24797);
nand UO_124 (O_124,N_24973,N_24616);
xnor UO_125 (O_125,N_24734,N_24731);
and UO_126 (O_126,N_24925,N_24808);
nor UO_127 (O_127,N_24655,N_24901);
xnor UO_128 (O_128,N_24686,N_24710);
or UO_129 (O_129,N_24640,N_24916);
nor UO_130 (O_130,N_24773,N_24652);
and UO_131 (O_131,N_24911,N_24818);
nand UO_132 (O_132,N_24822,N_24872);
xnor UO_133 (O_133,N_24743,N_24947);
xor UO_134 (O_134,N_24926,N_24828);
or UO_135 (O_135,N_24657,N_24986);
nand UO_136 (O_136,N_24900,N_24665);
and UO_137 (O_137,N_24515,N_24508);
nor UO_138 (O_138,N_24945,N_24767);
nand UO_139 (O_139,N_24841,N_24668);
nor UO_140 (O_140,N_24620,N_24759);
xnor UO_141 (O_141,N_24660,N_24787);
nand UO_142 (O_142,N_24582,N_24545);
nand UO_143 (O_143,N_24942,N_24949);
and UO_144 (O_144,N_24871,N_24560);
and UO_145 (O_145,N_24850,N_24606);
and UO_146 (O_146,N_24932,N_24802);
and UO_147 (O_147,N_24791,N_24720);
and UO_148 (O_148,N_24615,N_24717);
or UO_149 (O_149,N_24751,N_24847);
nor UO_150 (O_150,N_24666,N_24607);
xor UO_151 (O_151,N_24634,N_24623);
nand UO_152 (O_152,N_24976,N_24856);
nor UO_153 (O_153,N_24930,N_24541);
and UO_154 (O_154,N_24909,N_24903);
xor UO_155 (O_155,N_24910,N_24899);
and UO_156 (O_156,N_24915,N_24718);
nand UO_157 (O_157,N_24881,N_24565);
nor UO_158 (O_158,N_24568,N_24878);
or UO_159 (O_159,N_24931,N_24951);
xnor UO_160 (O_160,N_24590,N_24649);
nand UO_161 (O_161,N_24877,N_24843);
xor UO_162 (O_162,N_24642,N_24725);
nor UO_163 (O_163,N_24766,N_24805);
xnor UO_164 (O_164,N_24739,N_24688);
xor UO_165 (O_165,N_24829,N_24771);
nor UO_166 (O_166,N_24511,N_24967);
and UO_167 (O_167,N_24701,N_24638);
xor UO_168 (O_168,N_24748,N_24869);
and UO_169 (O_169,N_24827,N_24578);
nand UO_170 (O_170,N_24752,N_24792);
xnor UO_171 (O_171,N_24969,N_24941);
xnor UO_172 (O_172,N_24677,N_24753);
or UO_173 (O_173,N_24913,N_24834);
xor UO_174 (O_174,N_24598,N_24593);
or UO_175 (O_175,N_24507,N_24804);
and UO_176 (O_176,N_24852,N_24981);
or UO_177 (O_177,N_24904,N_24857);
nand UO_178 (O_178,N_24537,N_24833);
xor UO_179 (O_179,N_24968,N_24552);
or UO_180 (O_180,N_24622,N_24536);
xnor UO_181 (O_181,N_24740,N_24505);
nand UO_182 (O_182,N_24542,N_24819);
xor UO_183 (O_183,N_24693,N_24594);
xnor UO_184 (O_184,N_24601,N_24597);
and UO_185 (O_185,N_24985,N_24896);
nand UO_186 (O_186,N_24723,N_24564);
xnor UO_187 (O_187,N_24531,N_24994);
and UO_188 (O_188,N_24661,N_24609);
and UO_189 (O_189,N_24635,N_24826);
and UO_190 (O_190,N_24937,N_24613);
or UO_191 (O_191,N_24645,N_24708);
nand UO_192 (O_192,N_24990,N_24699);
and UO_193 (O_193,N_24864,N_24830);
or UO_194 (O_194,N_24539,N_24955);
xnor UO_195 (O_195,N_24775,N_24943);
nor UO_196 (O_196,N_24770,N_24705);
nand UO_197 (O_197,N_24855,N_24696);
xor UO_198 (O_198,N_24888,N_24761);
nor UO_199 (O_199,N_24892,N_24716);
xnor UO_200 (O_200,N_24972,N_24618);
nor UO_201 (O_201,N_24745,N_24692);
nor UO_202 (O_202,N_24684,N_24728);
and UO_203 (O_203,N_24936,N_24721);
nor UO_204 (O_204,N_24674,N_24939);
nand UO_205 (O_205,N_24584,N_24854);
and UO_206 (O_206,N_24516,N_24816);
or UO_207 (O_207,N_24595,N_24586);
xnor UO_208 (O_208,N_24982,N_24679);
or UO_209 (O_209,N_24636,N_24706);
and UO_210 (O_210,N_24933,N_24832);
and UO_211 (O_211,N_24678,N_24563);
or UO_212 (O_212,N_24912,N_24574);
nor UO_213 (O_213,N_24534,N_24713);
xnor UO_214 (O_214,N_24848,N_24873);
and UO_215 (O_215,N_24709,N_24786);
nor UO_216 (O_216,N_24501,N_24522);
nand UO_217 (O_217,N_24836,N_24880);
xnor UO_218 (O_218,N_24844,N_24527);
or UO_219 (O_219,N_24921,N_24853);
nor UO_220 (O_220,N_24612,N_24946);
nor UO_221 (O_221,N_24765,N_24585);
and UO_222 (O_222,N_24789,N_24512);
xor UO_223 (O_223,N_24778,N_24529);
xnor UO_224 (O_224,N_24914,N_24839);
or UO_225 (O_225,N_24866,N_24963);
nor UO_226 (O_226,N_24579,N_24784);
or UO_227 (O_227,N_24917,N_24577);
and UO_228 (O_228,N_24625,N_24825);
or UO_229 (O_229,N_24627,N_24757);
or UO_230 (O_230,N_24629,N_24971);
and UO_231 (O_231,N_24632,N_24983);
xor UO_232 (O_232,N_24846,N_24948);
and UO_233 (O_233,N_24952,N_24950);
xnor UO_234 (O_234,N_24884,N_24768);
xnor UO_235 (O_235,N_24673,N_24923);
or UO_236 (O_236,N_24781,N_24958);
or UO_237 (O_237,N_24813,N_24580);
nand UO_238 (O_238,N_24532,N_24993);
nor UO_239 (O_239,N_24956,N_24820);
nand UO_240 (O_240,N_24528,N_24960);
and UO_241 (O_241,N_24744,N_24600);
nor UO_242 (O_242,N_24987,N_24978);
nand UO_243 (O_243,N_24865,N_24523);
and UO_244 (O_244,N_24547,N_24898);
nor UO_245 (O_245,N_24764,N_24803);
xor UO_246 (O_246,N_24628,N_24897);
or UO_247 (O_247,N_24975,N_24653);
or UO_248 (O_248,N_24544,N_24517);
or UO_249 (O_249,N_24671,N_24929);
and UO_250 (O_250,N_24999,N_24848);
nand UO_251 (O_251,N_24944,N_24589);
nand UO_252 (O_252,N_24878,N_24876);
nor UO_253 (O_253,N_24915,N_24743);
and UO_254 (O_254,N_24916,N_24938);
nand UO_255 (O_255,N_24761,N_24606);
and UO_256 (O_256,N_24642,N_24740);
and UO_257 (O_257,N_24649,N_24941);
or UO_258 (O_258,N_24805,N_24961);
nand UO_259 (O_259,N_24935,N_24773);
or UO_260 (O_260,N_24803,N_24734);
nor UO_261 (O_261,N_24973,N_24935);
nand UO_262 (O_262,N_24594,N_24554);
nor UO_263 (O_263,N_24553,N_24859);
xnor UO_264 (O_264,N_24715,N_24847);
nand UO_265 (O_265,N_24576,N_24748);
nor UO_266 (O_266,N_24792,N_24770);
nand UO_267 (O_267,N_24849,N_24824);
nand UO_268 (O_268,N_24725,N_24553);
nand UO_269 (O_269,N_24977,N_24699);
nor UO_270 (O_270,N_24975,N_24691);
nand UO_271 (O_271,N_24855,N_24541);
nand UO_272 (O_272,N_24710,N_24943);
and UO_273 (O_273,N_24719,N_24842);
or UO_274 (O_274,N_24747,N_24766);
or UO_275 (O_275,N_24804,N_24917);
and UO_276 (O_276,N_24578,N_24754);
xnor UO_277 (O_277,N_24600,N_24927);
nor UO_278 (O_278,N_24514,N_24557);
and UO_279 (O_279,N_24814,N_24513);
nor UO_280 (O_280,N_24541,N_24592);
nand UO_281 (O_281,N_24625,N_24999);
or UO_282 (O_282,N_24975,N_24675);
and UO_283 (O_283,N_24672,N_24996);
and UO_284 (O_284,N_24893,N_24905);
and UO_285 (O_285,N_24675,N_24711);
or UO_286 (O_286,N_24740,N_24753);
nor UO_287 (O_287,N_24841,N_24674);
and UO_288 (O_288,N_24701,N_24706);
nand UO_289 (O_289,N_24510,N_24519);
nor UO_290 (O_290,N_24869,N_24534);
xor UO_291 (O_291,N_24532,N_24756);
or UO_292 (O_292,N_24791,N_24927);
nand UO_293 (O_293,N_24594,N_24805);
and UO_294 (O_294,N_24982,N_24935);
nor UO_295 (O_295,N_24723,N_24852);
nand UO_296 (O_296,N_24803,N_24921);
and UO_297 (O_297,N_24665,N_24991);
xor UO_298 (O_298,N_24634,N_24879);
nand UO_299 (O_299,N_24602,N_24960);
or UO_300 (O_300,N_24566,N_24789);
nand UO_301 (O_301,N_24910,N_24651);
and UO_302 (O_302,N_24624,N_24677);
xor UO_303 (O_303,N_24746,N_24868);
xor UO_304 (O_304,N_24705,N_24939);
nor UO_305 (O_305,N_24858,N_24787);
nand UO_306 (O_306,N_24500,N_24537);
or UO_307 (O_307,N_24895,N_24662);
nand UO_308 (O_308,N_24741,N_24666);
xnor UO_309 (O_309,N_24839,N_24528);
and UO_310 (O_310,N_24807,N_24874);
nor UO_311 (O_311,N_24549,N_24579);
or UO_312 (O_312,N_24983,N_24802);
nand UO_313 (O_313,N_24582,N_24845);
xor UO_314 (O_314,N_24674,N_24831);
nor UO_315 (O_315,N_24827,N_24901);
or UO_316 (O_316,N_24652,N_24992);
and UO_317 (O_317,N_24794,N_24525);
and UO_318 (O_318,N_24590,N_24720);
nor UO_319 (O_319,N_24550,N_24594);
xnor UO_320 (O_320,N_24912,N_24828);
and UO_321 (O_321,N_24583,N_24532);
and UO_322 (O_322,N_24969,N_24693);
nor UO_323 (O_323,N_24624,N_24523);
and UO_324 (O_324,N_24693,N_24962);
nor UO_325 (O_325,N_24623,N_24812);
nand UO_326 (O_326,N_24986,N_24873);
and UO_327 (O_327,N_24749,N_24644);
and UO_328 (O_328,N_24902,N_24904);
and UO_329 (O_329,N_24850,N_24848);
and UO_330 (O_330,N_24521,N_24675);
and UO_331 (O_331,N_24810,N_24769);
and UO_332 (O_332,N_24889,N_24782);
nand UO_333 (O_333,N_24939,N_24529);
and UO_334 (O_334,N_24566,N_24925);
nor UO_335 (O_335,N_24636,N_24728);
xnor UO_336 (O_336,N_24864,N_24716);
nand UO_337 (O_337,N_24953,N_24967);
nand UO_338 (O_338,N_24588,N_24549);
nand UO_339 (O_339,N_24779,N_24925);
xor UO_340 (O_340,N_24664,N_24738);
nand UO_341 (O_341,N_24709,N_24759);
xnor UO_342 (O_342,N_24843,N_24749);
and UO_343 (O_343,N_24950,N_24873);
nand UO_344 (O_344,N_24968,N_24926);
xor UO_345 (O_345,N_24731,N_24620);
or UO_346 (O_346,N_24520,N_24710);
nor UO_347 (O_347,N_24745,N_24793);
nor UO_348 (O_348,N_24735,N_24870);
and UO_349 (O_349,N_24627,N_24711);
nor UO_350 (O_350,N_24786,N_24676);
and UO_351 (O_351,N_24955,N_24678);
and UO_352 (O_352,N_24782,N_24648);
nor UO_353 (O_353,N_24539,N_24745);
nor UO_354 (O_354,N_24560,N_24861);
nand UO_355 (O_355,N_24966,N_24882);
xnor UO_356 (O_356,N_24588,N_24643);
nand UO_357 (O_357,N_24786,N_24720);
or UO_358 (O_358,N_24777,N_24628);
and UO_359 (O_359,N_24903,N_24503);
or UO_360 (O_360,N_24506,N_24627);
nand UO_361 (O_361,N_24580,N_24596);
nand UO_362 (O_362,N_24932,N_24714);
or UO_363 (O_363,N_24804,N_24627);
and UO_364 (O_364,N_24711,N_24826);
xnor UO_365 (O_365,N_24539,N_24713);
nand UO_366 (O_366,N_24629,N_24742);
or UO_367 (O_367,N_24679,N_24897);
and UO_368 (O_368,N_24516,N_24753);
or UO_369 (O_369,N_24640,N_24899);
nor UO_370 (O_370,N_24695,N_24981);
nor UO_371 (O_371,N_24771,N_24535);
xor UO_372 (O_372,N_24956,N_24926);
and UO_373 (O_373,N_24919,N_24774);
or UO_374 (O_374,N_24969,N_24505);
nor UO_375 (O_375,N_24746,N_24748);
nor UO_376 (O_376,N_24736,N_24518);
and UO_377 (O_377,N_24645,N_24537);
or UO_378 (O_378,N_24918,N_24731);
or UO_379 (O_379,N_24940,N_24912);
or UO_380 (O_380,N_24521,N_24767);
xnor UO_381 (O_381,N_24939,N_24582);
nor UO_382 (O_382,N_24819,N_24975);
nor UO_383 (O_383,N_24599,N_24848);
nand UO_384 (O_384,N_24649,N_24575);
xor UO_385 (O_385,N_24730,N_24743);
nand UO_386 (O_386,N_24551,N_24624);
nor UO_387 (O_387,N_24945,N_24875);
xor UO_388 (O_388,N_24639,N_24564);
nor UO_389 (O_389,N_24568,N_24854);
and UO_390 (O_390,N_24896,N_24577);
or UO_391 (O_391,N_24910,N_24711);
nor UO_392 (O_392,N_24778,N_24604);
or UO_393 (O_393,N_24684,N_24609);
and UO_394 (O_394,N_24873,N_24524);
xnor UO_395 (O_395,N_24903,N_24926);
nor UO_396 (O_396,N_24546,N_24656);
and UO_397 (O_397,N_24667,N_24723);
nor UO_398 (O_398,N_24681,N_24692);
or UO_399 (O_399,N_24984,N_24802);
or UO_400 (O_400,N_24584,N_24861);
and UO_401 (O_401,N_24957,N_24571);
or UO_402 (O_402,N_24502,N_24734);
and UO_403 (O_403,N_24819,N_24633);
xor UO_404 (O_404,N_24999,N_24595);
nor UO_405 (O_405,N_24847,N_24741);
nor UO_406 (O_406,N_24931,N_24893);
nor UO_407 (O_407,N_24563,N_24553);
and UO_408 (O_408,N_24756,N_24969);
and UO_409 (O_409,N_24507,N_24635);
and UO_410 (O_410,N_24813,N_24582);
xnor UO_411 (O_411,N_24602,N_24585);
nand UO_412 (O_412,N_24514,N_24526);
nor UO_413 (O_413,N_24567,N_24756);
nand UO_414 (O_414,N_24737,N_24721);
nand UO_415 (O_415,N_24591,N_24948);
xor UO_416 (O_416,N_24609,N_24724);
nor UO_417 (O_417,N_24636,N_24775);
nor UO_418 (O_418,N_24882,N_24725);
and UO_419 (O_419,N_24992,N_24657);
or UO_420 (O_420,N_24803,N_24788);
xnor UO_421 (O_421,N_24582,N_24783);
nand UO_422 (O_422,N_24797,N_24556);
or UO_423 (O_423,N_24679,N_24512);
and UO_424 (O_424,N_24862,N_24714);
nor UO_425 (O_425,N_24551,N_24884);
or UO_426 (O_426,N_24526,N_24539);
nor UO_427 (O_427,N_24725,N_24849);
or UO_428 (O_428,N_24740,N_24628);
nor UO_429 (O_429,N_24895,N_24996);
xnor UO_430 (O_430,N_24703,N_24697);
or UO_431 (O_431,N_24579,N_24731);
nand UO_432 (O_432,N_24777,N_24695);
or UO_433 (O_433,N_24779,N_24583);
nand UO_434 (O_434,N_24630,N_24819);
and UO_435 (O_435,N_24960,N_24951);
xor UO_436 (O_436,N_24663,N_24964);
nor UO_437 (O_437,N_24930,N_24860);
and UO_438 (O_438,N_24976,N_24882);
nand UO_439 (O_439,N_24527,N_24633);
and UO_440 (O_440,N_24548,N_24761);
nand UO_441 (O_441,N_24756,N_24816);
or UO_442 (O_442,N_24785,N_24663);
nor UO_443 (O_443,N_24901,N_24920);
and UO_444 (O_444,N_24608,N_24515);
xor UO_445 (O_445,N_24591,N_24998);
nor UO_446 (O_446,N_24811,N_24820);
and UO_447 (O_447,N_24968,N_24871);
nor UO_448 (O_448,N_24970,N_24656);
xnor UO_449 (O_449,N_24932,N_24906);
or UO_450 (O_450,N_24650,N_24939);
xnor UO_451 (O_451,N_24676,N_24779);
nor UO_452 (O_452,N_24546,N_24716);
and UO_453 (O_453,N_24636,N_24568);
nand UO_454 (O_454,N_24911,N_24861);
and UO_455 (O_455,N_24873,N_24937);
nand UO_456 (O_456,N_24907,N_24658);
nand UO_457 (O_457,N_24962,N_24940);
nor UO_458 (O_458,N_24833,N_24722);
nand UO_459 (O_459,N_24770,N_24543);
nor UO_460 (O_460,N_24703,N_24552);
or UO_461 (O_461,N_24831,N_24853);
xnor UO_462 (O_462,N_24524,N_24529);
nor UO_463 (O_463,N_24751,N_24759);
or UO_464 (O_464,N_24839,N_24729);
nand UO_465 (O_465,N_24657,N_24691);
or UO_466 (O_466,N_24810,N_24513);
xor UO_467 (O_467,N_24829,N_24656);
xor UO_468 (O_468,N_24740,N_24596);
or UO_469 (O_469,N_24739,N_24569);
and UO_470 (O_470,N_24887,N_24725);
nand UO_471 (O_471,N_24534,N_24977);
nand UO_472 (O_472,N_24610,N_24884);
xnor UO_473 (O_473,N_24953,N_24870);
nor UO_474 (O_474,N_24682,N_24792);
nor UO_475 (O_475,N_24866,N_24657);
xnor UO_476 (O_476,N_24737,N_24984);
and UO_477 (O_477,N_24568,N_24654);
and UO_478 (O_478,N_24517,N_24841);
nand UO_479 (O_479,N_24669,N_24852);
or UO_480 (O_480,N_24624,N_24520);
and UO_481 (O_481,N_24618,N_24747);
nand UO_482 (O_482,N_24748,N_24597);
nand UO_483 (O_483,N_24652,N_24637);
nand UO_484 (O_484,N_24929,N_24526);
nor UO_485 (O_485,N_24679,N_24585);
or UO_486 (O_486,N_24984,N_24504);
nand UO_487 (O_487,N_24990,N_24657);
xor UO_488 (O_488,N_24763,N_24918);
nor UO_489 (O_489,N_24577,N_24963);
and UO_490 (O_490,N_24902,N_24964);
nor UO_491 (O_491,N_24888,N_24578);
and UO_492 (O_492,N_24746,N_24747);
or UO_493 (O_493,N_24590,N_24897);
or UO_494 (O_494,N_24624,N_24554);
or UO_495 (O_495,N_24618,N_24756);
nand UO_496 (O_496,N_24791,N_24788);
and UO_497 (O_497,N_24821,N_24839);
or UO_498 (O_498,N_24505,N_24811);
nor UO_499 (O_499,N_24536,N_24599);
nor UO_500 (O_500,N_24711,N_24992);
nor UO_501 (O_501,N_24832,N_24640);
or UO_502 (O_502,N_24798,N_24654);
nor UO_503 (O_503,N_24826,N_24771);
xor UO_504 (O_504,N_24520,N_24630);
and UO_505 (O_505,N_24523,N_24872);
nor UO_506 (O_506,N_24997,N_24751);
and UO_507 (O_507,N_24912,N_24889);
nand UO_508 (O_508,N_24509,N_24786);
nand UO_509 (O_509,N_24755,N_24602);
nand UO_510 (O_510,N_24771,N_24503);
or UO_511 (O_511,N_24985,N_24640);
or UO_512 (O_512,N_24707,N_24545);
and UO_513 (O_513,N_24775,N_24528);
or UO_514 (O_514,N_24815,N_24870);
nor UO_515 (O_515,N_24728,N_24726);
xnor UO_516 (O_516,N_24842,N_24638);
xnor UO_517 (O_517,N_24917,N_24823);
nor UO_518 (O_518,N_24798,N_24693);
or UO_519 (O_519,N_24571,N_24936);
or UO_520 (O_520,N_24892,N_24758);
xnor UO_521 (O_521,N_24953,N_24663);
nand UO_522 (O_522,N_24872,N_24637);
and UO_523 (O_523,N_24966,N_24637);
or UO_524 (O_524,N_24614,N_24817);
or UO_525 (O_525,N_24956,N_24602);
nand UO_526 (O_526,N_24975,N_24892);
and UO_527 (O_527,N_24855,N_24763);
and UO_528 (O_528,N_24531,N_24730);
or UO_529 (O_529,N_24726,N_24533);
and UO_530 (O_530,N_24741,N_24912);
or UO_531 (O_531,N_24782,N_24894);
and UO_532 (O_532,N_24961,N_24874);
nor UO_533 (O_533,N_24933,N_24729);
xnor UO_534 (O_534,N_24638,N_24729);
xor UO_535 (O_535,N_24534,N_24991);
nor UO_536 (O_536,N_24692,N_24599);
nand UO_537 (O_537,N_24652,N_24781);
or UO_538 (O_538,N_24502,N_24700);
or UO_539 (O_539,N_24885,N_24732);
and UO_540 (O_540,N_24722,N_24618);
xnor UO_541 (O_541,N_24553,N_24536);
nor UO_542 (O_542,N_24891,N_24796);
nand UO_543 (O_543,N_24912,N_24850);
or UO_544 (O_544,N_24701,N_24745);
nor UO_545 (O_545,N_24900,N_24608);
xnor UO_546 (O_546,N_24616,N_24673);
or UO_547 (O_547,N_24983,N_24873);
and UO_548 (O_548,N_24999,N_24993);
nor UO_549 (O_549,N_24987,N_24730);
or UO_550 (O_550,N_24868,N_24664);
xnor UO_551 (O_551,N_24861,N_24825);
and UO_552 (O_552,N_24969,N_24791);
xnor UO_553 (O_553,N_24627,N_24893);
xor UO_554 (O_554,N_24696,N_24852);
nand UO_555 (O_555,N_24929,N_24993);
nand UO_556 (O_556,N_24823,N_24627);
or UO_557 (O_557,N_24906,N_24940);
and UO_558 (O_558,N_24987,N_24836);
xnor UO_559 (O_559,N_24569,N_24557);
nand UO_560 (O_560,N_24803,N_24905);
and UO_561 (O_561,N_24822,N_24895);
nand UO_562 (O_562,N_24828,N_24507);
nor UO_563 (O_563,N_24714,N_24673);
or UO_564 (O_564,N_24554,N_24715);
xor UO_565 (O_565,N_24831,N_24694);
and UO_566 (O_566,N_24772,N_24871);
nor UO_567 (O_567,N_24829,N_24861);
or UO_568 (O_568,N_24999,N_24816);
and UO_569 (O_569,N_24661,N_24560);
and UO_570 (O_570,N_24903,N_24957);
nand UO_571 (O_571,N_24607,N_24764);
and UO_572 (O_572,N_24569,N_24577);
nand UO_573 (O_573,N_24921,N_24744);
nor UO_574 (O_574,N_24660,N_24899);
nor UO_575 (O_575,N_24681,N_24745);
and UO_576 (O_576,N_24654,N_24853);
and UO_577 (O_577,N_24651,N_24521);
xor UO_578 (O_578,N_24865,N_24870);
nand UO_579 (O_579,N_24894,N_24574);
nand UO_580 (O_580,N_24887,N_24964);
nor UO_581 (O_581,N_24726,N_24580);
and UO_582 (O_582,N_24748,N_24925);
nand UO_583 (O_583,N_24804,N_24803);
or UO_584 (O_584,N_24722,N_24897);
or UO_585 (O_585,N_24678,N_24934);
or UO_586 (O_586,N_24634,N_24508);
nand UO_587 (O_587,N_24564,N_24668);
and UO_588 (O_588,N_24726,N_24780);
and UO_589 (O_589,N_24881,N_24808);
and UO_590 (O_590,N_24942,N_24958);
nor UO_591 (O_591,N_24672,N_24909);
nand UO_592 (O_592,N_24658,N_24985);
xor UO_593 (O_593,N_24657,N_24994);
and UO_594 (O_594,N_24780,N_24681);
and UO_595 (O_595,N_24711,N_24871);
and UO_596 (O_596,N_24907,N_24653);
or UO_597 (O_597,N_24976,N_24794);
and UO_598 (O_598,N_24526,N_24927);
or UO_599 (O_599,N_24528,N_24693);
or UO_600 (O_600,N_24737,N_24862);
nand UO_601 (O_601,N_24508,N_24822);
nor UO_602 (O_602,N_24515,N_24800);
and UO_603 (O_603,N_24558,N_24693);
nand UO_604 (O_604,N_24711,N_24619);
nor UO_605 (O_605,N_24574,N_24880);
or UO_606 (O_606,N_24588,N_24774);
nand UO_607 (O_607,N_24543,N_24596);
xor UO_608 (O_608,N_24628,N_24621);
xnor UO_609 (O_609,N_24712,N_24982);
xor UO_610 (O_610,N_24977,N_24702);
xnor UO_611 (O_611,N_24975,N_24572);
nor UO_612 (O_612,N_24931,N_24899);
xor UO_613 (O_613,N_24814,N_24998);
xnor UO_614 (O_614,N_24681,N_24900);
nand UO_615 (O_615,N_24853,N_24840);
xor UO_616 (O_616,N_24988,N_24832);
nor UO_617 (O_617,N_24688,N_24938);
xor UO_618 (O_618,N_24818,N_24627);
nor UO_619 (O_619,N_24766,N_24981);
nand UO_620 (O_620,N_24756,N_24888);
nand UO_621 (O_621,N_24701,N_24904);
nand UO_622 (O_622,N_24809,N_24610);
nor UO_623 (O_623,N_24643,N_24872);
or UO_624 (O_624,N_24969,N_24625);
nor UO_625 (O_625,N_24774,N_24747);
nand UO_626 (O_626,N_24790,N_24810);
and UO_627 (O_627,N_24532,N_24903);
and UO_628 (O_628,N_24898,N_24600);
nor UO_629 (O_629,N_24976,N_24545);
nor UO_630 (O_630,N_24633,N_24959);
nand UO_631 (O_631,N_24560,N_24500);
or UO_632 (O_632,N_24733,N_24711);
or UO_633 (O_633,N_24905,N_24968);
xnor UO_634 (O_634,N_24979,N_24535);
nor UO_635 (O_635,N_24523,N_24806);
or UO_636 (O_636,N_24813,N_24691);
and UO_637 (O_637,N_24762,N_24579);
xnor UO_638 (O_638,N_24937,N_24962);
and UO_639 (O_639,N_24599,N_24813);
and UO_640 (O_640,N_24643,N_24778);
nor UO_641 (O_641,N_24662,N_24684);
and UO_642 (O_642,N_24608,N_24999);
nand UO_643 (O_643,N_24973,N_24909);
xor UO_644 (O_644,N_24959,N_24746);
or UO_645 (O_645,N_24935,N_24881);
or UO_646 (O_646,N_24879,N_24554);
and UO_647 (O_647,N_24582,N_24519);
nor UO_648 (O_648,N_24688,N_24625);
xor UO_649 (O_649,N_24949,N_24579);
nand UO_650 (O_650,N_24668,N_24855);
and UO_651 (O_651,N_24894,N_24850);
xor UO_652 (O_652,N_24699,N_24832);
and UO_653 (O_653,N_24874,N_24882);
nor UO_654 (O_654,N_24561,N_24906);
nor UO_655 (O_655,N_24994,N_24804);
xor UO_656 (O_656,N_24636,N_24505);
nor UO_657 (O_657,N_24563,N_24518);
or UO_658 (O_658,N_24772,N_24797);
nor UO_659 (O_659,N_24669,N_24924);
nor UO_660 (O_660,N_24650,N_24643);
nor UO_661 (O_661,N_24547,N_24911);
nor UO_662 (O_662,N_24655,N_24862);
nor UO_663 (O_663,N_24504,N_24856);
nand UO_664 (O_664,N_24599,N_24731);
nor UO_665 (O_665,N_24700,N_24922);
and UO_666 (O_666,N_24988,N_24736);
and UO_667 (O_667,N_24832,N_24580);
nand UO_668 (O_668,N_24893,N_24563);
nand UO_669 (O_669,N_24619,N_24631);
nand UO_670 (O_670,N_24995,N_24862);
or UO_671 (O_671,N_24891,N_24774);
xor UO_672 (O_672,N_24578,N_24748);
nor UO_673 (O_673,N_24928,N_24857);
or UO_674 (O_674,N_24801,N_24930);
nor UO_675 (O_675,N_24972,N_24774);
xnor UO_676 (O_676,N_24589,N_24972);
and UO_677 (O_677,N_24610,N_24524);
and UO_678 (O_678,N_24826,N_24751);
nand UO_679 (O_679,N_24753,N_24739);
or UO_680 (O_680,N_24878,N_24914);
xor UO_681 (O_681,N_24555,N_24695);
nand UO_682 (O_682,N_24993,N_24995);
xor UO_683 (O_683,N_24642,N_24509);
nor UO_684 (O_684,N_24528,N_24709);
xnor UO_685 (O_685,N_24950,N_24968);
nand UO_686 (O_686,N_24977,N_24738);
xnor UO_687 (O_687,N_24939,N_24745);
nor UO_688 (O_688,N_24568,N_24970);
nor UO_689 (O_689,N_24894,N_24934);
nor UO_690 (O_690,N_24791,N_24576);
xor UO_691 (O_691,N_24848,N_24613);
and UO_692 (O_692,N_24723,N_24937);
xor UO_693 (O_693,N_24790,N_24780);
xnor UO_694 (O_694,N_24894,N_24940);
and UO_695 (O_695,N_24546,N_24717);
nand UO_696 (O_696,N_24773,N_24808);
xor UO_697 (O_697,N_24799,N_24956);
nand UO_698 (O_698,N_24868,N_24624);
xnor UO_699 (O_699,N_24644,N_24616);
nand UO_700 (O_700,N_24576,N_24770);
and UO_701 (O_701,N_24784,N_24547);
nor UO_702 (O_702,N_24524,N_24864);
or UO_703 (O_703,N_24633,N_24875);
nand UO_704 (O_704,N_24932,N_24820);
xnor UO_705 (O_705,N_24798,N_24877);
and UO_706 (O_706,N_24964,N_24966);
xor UO_707 (O_707,N_24734,N_24862);
nand UO_708 (O_708,N_24611,N_24718);
and UO_709 (O_709,N_24855,N_24960);
or UO_710 (O_710,N_24978,N_24945);
nand UO_711 (O_711,N_24975,N_24866);
or UO_712 (O_712,N_24880,N_24533);
nand UO_713 (O_713,N_24811,N_24641);
nand UO_714 (O_714,N_24976,N_24864);
xor UO_715 (O_715,N_24999,N_24883);
nand UO_716 (O_716,N_24943,N_24963);
nand UO_717 (O_717,N_24631,N_24557);
nand UO_718 (O_718,N_24603,N_24674);
and UO_719 (O_719,N_24818,N_24503);
nor UO_720 (O_720,N_24508,N_24695);
or UO_721 (O_721,N_24904,N_24729);
and UO_722 (O_722,N_24794,N_24972);
xnor UO_723 (O_723,N_24514,N_24869);
or UO_724 (O_724,N_24635,N_24537);
and UO_725 (O_725,N_24770,N_24628);
nand UO_726 (O_726,N_24572,N_24929);
nand UO_727 (O_727,N_24832,N_24519);
or UO_728 (O_728,N_24993,N_24844);
nor UO_729 (O_729,N_24863,N_24559);
nand UO_730 (O_730,N_24842,N_24655);
or UO_731 (O_731,N_24641,N_24519);
xor UO_732 (O_732,N_24829,N_24696);
nand UO_733 (O_733,N_24685,N_24946);
nand UO_734 (O_734,N_24588,N_24616);
nor UO_735 (O_735,N_24637,N_24845);
nand UO_736 (O_736,N_24838,N_24672);
nand UO_737 (O_737,N_24559,N_24609);
xnor UO_738 (O_738,N_24978,N_24778);
nand UO_739 (O_739,N_24578,N_24929);
nand UO_740 (O_740,N_24982,N_24523);
or UO_741 (O_741,N_24898,N_24517);
and UO_742 (O_742,N_24884,N_24595);
nor UO_743 (O_743,N_24686,N_24877);
nand UO_744 (O_744,N_24739,N_24646);
and UO_745 (O_745,N_24629,N_24810);
or UO_746 (O_746,N_24814,N_24978);
nor UO_747 (O_747,N_24814,N_24651);
and UO_748 (O_748,N_24613,N_24555);
or UO_749 (O_749,N_24984,N_24574);
xor UO_750 (O_750,N_24650,N_24745);
nand UO_751 (O_751,N_24965,N_24824);
xor UO_752 (O_752,N_24642,N_24507);
nor UO_753 (O_753,N_24971,N_24952);
and UO_754 (O_754,N_24997,N_24995);
nand UO_755 (O_755,N_24760,N_24846);
nand UO_756 (O_756,N_24703,N_24867);
xor UO_757 (O_757,N_24599,N_24746);
nand UO_758 (O_758,N_24822,N_24661);
nand UO_759 (O_759,N_24823,N_24585);
and UO_760 (O_760,N_24661,N_24964);
nand UO_761 (O_761,N_24681,N_24671);
xnor UO_762 (O_762,N_24683,N_24757);
and UO_763 (O_763,N_24783,N_24747);
nand UO_764 (O_764,N_24726,N_24955);
xnor UO_765 (O_765,N_24884,N_24651);
nor UO_766 (O_766,N_24581,N_24520);
nand UO_767 (O_767,N_24511,N_24723);
and UO_768 (O_768,N_24563,N_24540);
nor UO_769 (O_769,N_24984,N_24657);
xor UO_770 (O_770,N_24916,N_24642);
xnor UO_771 (O_771,N_24582,N_24877);
xor UO_772 (O_772,N_24585,N_24729);
and UO_773 (O_773,N_24636,N_24937);
xor UO_774 (O_774,N_24980,N_24963);
and UO_775 (O_775,N_24833,N_24735);
and UO_776 (O_776,N_24802,N_24663);
nand UO_777 (O_777,N_24518,N_24644);
or UO_778 (O_778,N_24505,N_24520);
or UO_779 (O_779,N_24534,N_24708);
and UO_780 (O_780,N_24869,N_24872);
xor UO_781 (O_781,N_24503,N_24710);
xor UO_782 (O_782,N_24801,N_24662);
or UO_783 (O_783,N_24769,N_24578);
xnor UO_784 (O_784,N_24537,N_24700);
nand UO_785 (O_785,N_24874,N_24520);
or UO_786 (O_786,N_24588,N_24866);
nor UO_787 (O_787,N_24796,N_24765);
nand UO_788 (O_788,N_24591,N_24876);
xnor UO_789 (O_789,N_24856,N_24792);
xnor UO_790 (O_790,N_24762,N_24706);
or UO_791 (O_791,N_24907,N_24814);
or UO_792 (O_792,N_24554,N_24523);
nand UO_793 (O_793,N_24891,N_24600);
nand UO_794 (O_794,N_24841,N_24956);
nand UO_795 (O_795,N_24828,N_24551);
or UO_796 (O_796,N_24941,N_24978);
or UO_797 (O_797,N_24508,N_24594);
or UO_798 (O_798,N_24924,N_24945);
nor UO_799 (O_799,N_24586,N_24994);
nor UO_800 (O_800,N_24881,N_24508);
or UO_801 (O_801,N_24533,N_24811);
nand UO_802 (O_802,N_24540,N_24825);
and UO_803 (O_803,N_24626,N_24657);
xor UO_804 (O_804,N_24846,N_24885);
xnor UO_805 (O_805,N_24947,N_24584);
nor UO_806 (O_806,N_24978,N_24613);
or UO_807 (O_807,N_24935,N_24783);
or UO_808 (O_808,N_24938,N_24652);
or UO_809 (O_809,N_24581,N_24810);
nand UO_810 (O_810,N_24750,N_24613);
xnor UO_811 (O_811,N_24554,N_24686);
and UO_812 (O_812,N_24841,N_24977);
or UO_813 (O_813,N_24889,N_24500);
or UO_814 (O_814,N_24799,N_24728);
and UO_815 (O_815,N_24632,N_24740);
xor UO_816 (O_816,N_24725,N_24740);
xor UO_817 (O_817,N_24926,N_24538);
nor UO_818 (O_818,N_24799,N_24851);
or UO_819 (O_819,N_24916,N_24982);
nor UO_820 (O_820,N_24686,N_24715);
nor UO_821 (O_821,N_24610,N_24737);
or UO_822 (O_822,N_24753,N_24526);
or UO_823 (O_823,N_24589,N_24769);
xor UO_824 (O_824,N_24944,N_24721);
or UO_825 (O_825,N_24891,N_24809);
nand UO_826 (O_826,N_24573,N_24937);
nor UO_827 (O_827,N_24837,N_24657);
and UO_828 (O_828,N_24762,N_24586);
nor UO_829 (O_829,N_24663,N_24869);
nand UO_830 (O_830,N_24929,N_24893);
xor UO_831 (O_831,N_24771,N_24750);
nand UO_832 (O_832,N_24710,N_24988);
or UO_833 (O_833,N_24626,N_24694);
nor UO_834 (O_834,N_24697,N_24519);
nor UO_835 (O_835,N_24552,N_24541);
nor UO_836 (O_836,N_24653,N_24854);
nor UO_837 (O_837,N_24727,N_24734);
xor UO_838 (O_838,N_24680,N_24765);
or UO_839 (O_839,N_24565,N_24900);
nand UO_840 (O_840,N_24635,N_24985);
or UO_841 (O_841,N_24654,N_24851);
nand UO_842 (O_842,N_24943,N_24844);
nor UO_843 (O_843,N_24843,N_24708);
nand UO_844 (O_844,N_24978,N_24615);
xnor UO_845 (O_845,N_24838,N_24976);
nand UO_846 (O_846,N_24891,N_24968);
or UO_847 (O_847,N_24711,N_24899);
or UO_848 (O_848,N_24712,N_24954);
xnor UO_849 (O_849,N_24829,N_24929);
or UO_850 (O_850,N_24907,N_24875);
xor UO_851 (O_851,N_24923,N_24796);
nand UO_852 (O_852,N_24520,N_24689);
xnor UO_853 (O_853,N_24708,N_24511);
nor UO_854 (O_854,N_24592,N_24701);
xor UO_855 (O_855,N_24862,N_24890);
and UO_856 (O_856,N_24818,N_24854);
or UO_857 (O_857,N_24628,N_24739);
and UO_858 (O_858,N_24714,N_24723);
nand UO_859 (O_859,N_24804,N_24626);
nand UO_860 (O_860,N_24683,N_24829);
nand UO_861 (O_861,N_24810,N_24627);
nand UO_862 (O_862,N_24622,N_24890);
nor UO_863 (O_863,N_24666,N_24674);
and UO_864 (O_864,N_24676,N_24539);
and UO_865 (O_865,N_24940,N_24710);
nand UO_866 (O_866,N_24591,N_24991);
nor UO_867 (O_867,N_24791,N_24610);
nand UO_868 (O_868,N_24922,N_24750);
nand UO_869 (O_869,N_24960,N_24879);
or UO_870 (O_870,N_24799,N_24501);
nand UO_871 (O_871,N_24887,N_24549);
or UO_872 (O_872,N_24761,N_24511);
xnor UO_873 (O_873,N_24606,N_24656);
and UO_874 (O_874,N_24785,N_24996);
xor UO_875 (O_875,N_24987,N_24856);
xor UO_876 (O_876,N_24628,N_24543);
xnor UO_877 (O_877,N_24847,N_24864);
xor UO_878 (O_878,N_24741,N_24577);
xnor UO_879 (O_879,N_24675,N_24582);
or UO_880 (O_880,N_24551,N_24587);
or UO_881 (O_881,N_24673,N_24775);
and UO_882 (O_882,N_24848,N_24604);
nand UO_883 (O_883,N_24627,N_24581);
or UO_884 (O_884,N_24781,N_24912);
xnor UO_885 (O_885,N_24781,N_24627);
nand UO_886 (O_886,N_24986,N_24723);
or UO_887 (O_887,N_24895,N_24863);
xnor UO_888 (O_888,N_24989,N_24869);
xor UO_889 (O_889,N_24820,N_24751);
or UO_890 (O_890,N_24723,N_24626);
nand UO_891 (O_891,N_24641,N_24647);
nor UO_892 (O_892,N_24873,N_24567);
nor UO_893 (O_893,N_24881,N_24613);
or UO_894 (O_894,N_24635,N_24696);
or UO_895 (O_895,N_24803,N_24595);
xor UO_896 (O_896,N_24570,N_24592);
nor UO_897 (O_897,N_24950,N_24571);
nor UO_898 (O_898,N_24504,N_24935);
nand UO_899 (O_899,N_24987,N_24607);
xor UO_900 (O_900,N_24533,N_24872);
nand UO_901 (O_901,N_24542,N_24690);
nor UO_902 (O_902,N_24521,N_24586);
nand UO_903 (O_903,N_24616,N_24684);
xnor UO_904 (O_904,N_24513,N_24914);
nor UO_905 (O_905,N_24941,N_24595);
nor UO_906 (O_906,N_24708,N_24990);
nand UO_907 (O_907,N_24881,N_24554);
and UO_908 (O_908,N_24969,N_24606);
nor UO_909 (O_909,N_24570,N_24880);
or UO_910 (O_910,N_24701,N_24917);
and UO_911 (O_911,N_24769,N_24927);
xor UO_912 (O_912,N_24908,N_24827);
and UO_913 (O_913,N_24613,N_24638);
and UO_914 (O_914,N_24933,N_24905);
nor UO_915 (O_915,N_24667,N_24999);
nand UO_916 (O_916,N_24524,N_24683);
xor UO_917 (O_917,N_24729,N_24743);
xnor UO_918 (O_918,N_24904,N_24748);
nand UO_919 (O_919,N_24792,N_24939);
or UO_920 (O_920,N_24597,N_24856);
or UO_921 (O_921,N_24716,N_24615);
nand UO_922 (O_922,N_24694,N_24522);
xnor UO_923 (O_923,N_24705,N_24966);
or UO_924 (O_924,N_24519,N_24592);
xor UO_925 (O_925,N_24618,N_24602);
nor UO_926 (O_926,N_24980,N_24507);
or UO_927 (O_927,N_24651,N_24891);
nor UO_928 (O_928,N_24581,N_24814);
nor UO_929 (O_929,N_24655,N_24687);
or UO_930 (O_930,N_24789,N_24587);
or UO_931 (O_931,N_24760,N_24606);
xor UO_932 (O_932,N_24895,N_24600);
nor UO_933 (O_933,N_24936,N_24603);
and UO_934 (O_934,N_24787,N_24665);
nor UO_935 (O_935,N_24932,N_24848);
nand UO_936 (O_936,N_24762,N_24679);
or UO_937 (O_937,N_24666,N_24939);
nand UO_938 (O_938,N_24932,N_24908);
or UO_939 (O_939,N_24646,N_24834);
nor UO_940 (O_940,N_24949,N_24703);
xnor UO_941 (O_941,N_24679,N_24913);
xnor UO_942 (O_942,N_24676,N_24507);
nor UO_943 (O_943,N_24849,N_24748);
or UO_944 (O_944,N_24533,N_24577);
nand UO_945 (O_945,N_24540,N_24850);
or UO_946 (O_946,N_24728,N_24842);
nand UO_947 (O_947,N_24853,N_24578);
and UO_948 (O_948,N_24519,N_24985);
or UO_949 (O_949,N_24845,N_24664);
nand UO_950 (O_950,N_24538,N_24993);
nand UO_951 (O_951,N_24786,N_24677);
and UO_952 (O_952,N_24750,N_24973);
xnor UO_953 (O_953,N_24948,N_24645);
and UO_954 (O_954,N_24935,N_24646);
or UO_955 (O_955,N_24851,N_24646);
nand UO_956 (O_956,N_24773,N_24627);
and UO_957 (O_957,N_24784,N_24940);
nor UO_958 (O_958,N_24997,N_24714);
or UO_959 (O_959,N_24715,N_24552);
or UO_960 (O_960,N_24606,N_24749);
nor UO_961 (O_961,N_24955,N_24610);
nand UO_962 (O_962,N_24713,N_24601);
nor UO_963 (O_963,N_24799,N_24703);
nand UO_964 (O_964,N_24609,N_24871);
and UO_965 (O_965,N_24805,N_24705);
xnor UO_966 (O_966,N_24673,N_24751);
or UO_967 (O_967,N_24705,N_24624);
nand UO_968 (O_968,N_24869,N_24528);
or UO_969 (O_969,N_24824,N_24894);
and UO_970 (O_970,N_24628,N_24601);
xor UO_971 (O_971,N_24944,N_24875);
nand UO_972 (O_972,N_24577,N_24873);
nand UO_973 (O_973,N_24594,N_24903);
and UO_974 (O_974,N_24508,N_24836);
nor UO_975 (O_975,N_24956,N_24694);
nand UO_976 (O_976,N_24542,N_24858);
nor UO_977 (O_977,N_24830,N_24756);
nor UO_978 (O_978,N_24934,N_24968);
nor UO_979 (O_979,N_24569,N_24809);
or UO_980 (O_980,N_24645,N_24924);
nor UO_981 (O_981,N_24706,N_24734);
nor UO_982 (O_982,N_24801,N_24941);
nand UO_983 (O_983,N_24671,N_24659);
xnor UO_984 (O_984,N_24555,N_24947);
nor UO_985 (O_985,N_24659,N_24606);
or UO_986 (O_986,N_24909,N_24810);
or UO_987 (O_987,N_24835,N_24952);
xor UO_988 (O_988,N_24756,N_24999);
nand UO_989 (O_989,N_24761,N_24937);
or UO_990 (O_990,N_24885,N_24670);
nor UO_991 (O_991,N_24873,N_24977);
and UO_992 (O_992,N_24730,N_24626);
nand UO_993 (O_993,N_24660,N_24955);
or UO_994 (O_994,N_24703,N_24927);
and UO_995 (O_995,N_24798,N_24574);
nand UO_996 (O_996,N_24792,N_24740);
nor UO_997 (O_997,N_24729,N_24641);
nand UO_998 (O_998,N_24509,N_24979);
xnor UO_999 (O_999,N_24600,N_24514);
and UO_1000 (O_1000,N_24755,N_24949);
and UO_1001 (O_1001,N_24585,N_24924);
nor UO_1002 (O_1002,N_24519,N_24861);
or UO_1003 (O_1003,N_24851,N_24987);
nand UO_1004 (O_1004,N_24603,N_24939);
or UO_1005 (O_1005,N_24986,N_24560);
nand UO_1006 (O_1006,N_24652,N_24842);
xnor UO_1007 (O_1007,N_24807,N_24778);
xnor UO_1008 (O_1008,N_24714,N_24553);
xor UO_1009 (O_1009,N_24618,N_24936);
or UO_1010 (O_1010,N_24510,N_24594);
nor UO_1011 (O_1011,N_24766,N_24520);
nor UO_1012 (O_1012,N_24540,N_24725);
xnor UO_1013 (O_1013,N_24811,N_24748);
or UO_1014 (O_1014,N_24697,N_24940);
nand UO_1015 (O_1015,N_24822,N_24600);
xnor UO_1016 (O_1016,N_24980,N_24837);
and UO_1017 (O_1017,N_24943,N_24829);
nor UO_1018 (O_1018,N_24523,N_24934);
nand UO_1019 (O_1019,N_24803,N_24998);
nor UO_1020 (O_1020,N_24679,N_24748);
and UO_1021 (O_1021,N_24538,N_24925);
and UO_1022 (O_1022,N_24631,N_24551);
nand UO_1023 (O_1023,N_24873,N_24802);
nor UO_1024 (O_1024,N_24644,N_24708);
and UO_1025 (O_1025,N_24689,N_24747);
or UO_1026 (O_1026,N_24515,N_24698);
xor UO_1027 (O_1027,N_24877,N_24591);
xor UO_1028 (O_1028,N_24644,N_24958);
xnor UO_1029 (O_1029,N_24922,N_24644);
nor UO_1030 (O_1030,N_24802,N_24720);
xnor UO_1031 (O_1031,N_24885,N_24779);
and UO_1032 (O_1032,N_24863,N_24674);
or UO_1033 (O_1033,N_24570,N_24852);
or UO_1034 (O_1034,N_24990,N_24943);
or UO_1035 (O_1035,N_24971,N_24957);
nor UO_1036 (O_1036,N_24829,N_24523);
or UO_1037 (O_1037,N_24604,N_24719);
nand UO_1038 (O_1038,N_24953,N_24613);
xor UO_1039 (O_1039,N_24993,N_24951);
xnor UO_1040 (O_1040,N_24978,N_24915);
and UO_1041 (O_1041,N_24815,N_24739);
nor UO_1042 (O_1042,N_24881,N_24964);
xor UO_1043 (O_1043,N_24851,N_24867);
nand UO_1044 (O_1044,N_24661,N_24801);
nand UO_1045 (O_1045,N_24562,N_24583);
nor UO_1046 (O_1046,N_24602,N_24600);
xnor UO_1047 (O_1047,N_24996,N_24801);
nor UO_1048 (O_1048,N_24546,N_24700);
or UO_1049 (O_1049,N_24663,N_24832);
nor UO_1050 (O_1050,N_24542,N_24733);
nand UO_1051 (O_1051,N_24569,N_24512);
or UO_1052 (O_1052,N_24867,N_24692);
nand UO_1053 (O_1053,N_24562,N_24690);
xnor UO_1054 (O_1054,N_24829,N_24684);
or UO_1055 (O_1055,N_24990,N_24726);
nor UO_1056 (O_1056,N_24898,N_24621);
nor UO_1057 (O_1057,N_24781,N_24816);
nand UO_1058 (O_1058,N_24932,N_24564);
xnor UO_1059 (O_1059,N_24591,N_24515);
or UO_1060 (O_1060,N_24989,N_24813);
or UO_1061 (O_1061,N_24572,N_24801);
and UO_1062 (O_1062,N_24505,N_24993);
or UO_1063 (O_1063,N_24766,N_24889);
or UO_1064 (O_1064,N_24502,N_24867);
and UO_1065 (O_1065,N_24668,N_24597);
nand UO_1066 (O_1066,N_24561,N_24942);
or UO_1067 (O_1067,N_24626,N_24853);
xor UO_1068 (O_1068,N_24987,N_24640);
nor UO_1069 (O_1069,N_24779,N_24529);
xor UO_1070 (O_1070,N_24549,N_24558);
xor UO_1071 (O_1071,N_24749,N_24984);
and UO_1072 (O_1072,N_24523,N_24543);
nand UO_1073 (O_1073,N_24773,N_24565);
xor UO_1074 (O_1074,N_24908,N_24896);
xnor UO_1075 (O_1075,N_24975,N_24588);
xnor UO_1076 (O_1076,N_24842,N_24710);
nor UO_1077 (O_1077,N_24583,N_24918);
and UO_1078 (O_1078,N_24896,N_24607);
nor UO_1079 (O_1079,N_24737,N_24906);
and UO_1080 (O_1080,N_24713,N_24504);
nand UO_1081 (O_1081,N_24587,N_24876);
xor UO_1082 (O_1082,N_24643,N_24853);
xnor UO_1083 (O_1083,N_24654,N_24926);
nor UO_1084 (O_1084,N_24740,N_24512);
nor UO_1085 (O_1085,N_24984,N_24703);
or UO_1086 (O_1086,N_24660,N_24932);
and UO_1087 (O_1087,N_24614,N_24941);
xnor UO_1088 (O_1088,N_24869,N_24901);
xnor UO_1089 (O_1089,N_24565,N_24747);
nor UO_1090 (O_1090,N_24759,N_24835);
xnor UO_1091 (O_1091,N_24765,N_24904);
nand UO_1092 (O_1092,N_24632,N_24981);
xnor UO_1093 (O_1093,N_24515,N_24502);
nor UO_1094 (O_1094,N_24984,N_24623);
nor UO_1095 (O_1095,N_24673,N_24823);
nand UO_1096 (O_1096,N_24732,N_24775);
and UO_1097 (O_1097,N_24855,N_24898);
nand UO_1098 (O_1098,N_24559,N_24659);
xnor UO_1099 (O_1099,N_24799,N_24938);
nand UO_1100 (O_1100,N_24599,N_24902);
and UO_1101 (O_1101,N_24728,N_24873);
xnor UO_1102 (O_1102,N_24770,N_24500);
nand UO_1103 (O_1103,N_24997,N_24874);
and UO_1104 (O_1104,N_24504,N_24729);
nand UO_1105 (O_1105,N_24994,N_24909);
nor UO_1106 (O_1106,N_24553,N_24541);
or UO_1107 (O_1107,N_24861,N_24654);
nand UO_1108 (O_1108,N_24594,N_24853);
and UO_1109 (O_1109,N_24790,N_24905);
nor UO_1110 (O_1110,N_24526,N_24849);
and UO_1111 (O_1111,N_24608,N_24931);
or UO_1112 (O_1112,N_24677,N_24829);
xor UO_1113 (O_1113,N_24636,N_24796);
or UO_1114 (O_1114,N_24938,N_24693);
or UO_1115 (O_1115,N_24652,N_24880);
nand UO_1116 (O_1116,N_24826,N_24885);
xor UO_1117 (O_1117,N_24724,N_24552);
nand UO_1118 (O_1118,N_24740,N_24503);
nand UO_1119 (O_1119,N_24778,N_24804);
or UO_1120 (O_1120,N_24822,N_24954);
nor UO_1121 (O_1121,N_24698,N_24556);
xnor UO_1122 (O_1122,N_24797,N_24925);
nand UO_1123 (O_1123,N_24524,N_24555);
nand UO_1124 (O_1124,N_24744,N_24532);
or UO_1125 (O_1125,N_24566,N_24718);
xnor UO_1126 (O_1126,N_24845,N_24875);
or UO_1127 (O_1127,N_24534,N_24638);
xnor UO_1128 (O_1128,N_24787,N_24860);
or UO_1129 (O_1129,N_24531,N_24841);
nor UO_1130 (O_1130,N_24553,N_24881);
and UO_1131 (O_1131,N_24725,N_24913);
or UO_1132 (O_1132,N_24976,N_24715);
nand UO_1133 (O_1133,N_24636,N_24591);
or UO_1134 (O_1134,N_24831,N_24624);
nand UO_1135 (O_1135,N_24943,N_24530);
nor UO_1136 (O_1136,N_24792,N_24751);
and UO_1137 (O_1137,N_24577,N_24920);
xor UO_1138 (O_1138,N_24591,N_24776);
nand UO_1139 (O_1139,N_24807,N_24977);
xor UO_1140 (O_1140,N_24856,N_24540);
and UO_1141 (O_1141,N_24629,N_24529);
and UO_1142 (O_1142,N_24987,N_24862);
xnor UO_1143 (O_1143,N_24898,N_24940);
xnor UO_1144 (O_1144,N_24555,N_24637);
and UO_1145 (O_1145,N_24533,N_24585);
nor UO_1146 (O_1146,N_24944,N_24707);
and UO_1147 (O_1147,N_24619,N_24725);
and UO_1148 (O_1148,N_24937,N_24527);
or UO_1149 (O_1149,N_24815,N_24771);
nor UO_1150 (O_1150,N_24578,N_24962);
nand UO_1151 (O_1151,N_24686,N_24945);
and UO_1152 (O_1152,N_24970,N_24690);
and UO_1153 (O_1153,N_24526,N_24633);
and UO_1154 (O_1154,N_24758,N_24945);
nand UO_1155 (O_1155,N_24952,N_24565);
nand UO_1156 (O_1156,N_24918,N_24995);
nand UO_1157 (O_1157,N_24973,N_24631);
nor UO_1158 (O_1158,N_24650,N_24672);
xnor UO_1159 (O_1159,N_24819,N_24744);
and UO_1160 (O_1160,N_24979,N_24710);
xnor UO_1161 (O_1161,N_24692,N_24856);
xnor UO_1162 (O_1162,N_24891,N_24655);
or UO_1163 (O_1163,N_24943,N_24676);
and UO_1164 (O_1164,N_24634,N_24764);
or UO_1165 (O_1165,N_24871,N_24592);
xor UO_1166 (O_1166,N_24898,N_24554);
nor UO_1167 (O_1167,N_24692,N_24866);
or UO_1168 (O_1168,N_24645,N_24515);
or UO_1169 (O_1169,N_24648,N_24513);
nand UO_1170 (O_1170,N_24502,N_24506);
or UO_1171 (O_1171,N_24890,N_24540);
and UO_1172 (O_1172,N_24591,N_24842);
nand UO_1173 (O_1173,N_24716,N_24856);
and UO_1174 (O_1174,N_24941,N_24526);
and UO_1175 (O_1175,N_24791,N_24773);
or UO_1176 (O_1176,N_24879,N_24572);
and UO_1177 (O_1177,N_24588,N_24935);
or UO_1178 (O_1178,N_24509,N_24601);
or UO_1179 (O_1179,N_24823,N_24715);
nor UO_1180 (O_1180,N_24824,N_24581);
nand UO_1181 (O_1181,N_24635,N_24751);
and UO_1182 (O_1182,N_24584,N_24737);
and UO_1183 (O_1183,N_24754,N_24552);
nand UO_1184 (O_1184,N_24970,N_24518);
nor UO_1185 (O_1185,N_24730,N_24843);
nor UO_1186 (O_1186,N_24934,N_24822);
and UO_1187 (O_1187,N_24830,N_24769);
and UO_1188 (O_1188,N_24807,N_24682);
or UO_1189 (O_1189,N_24632,N_24989);
xor UO_1190 (O_1190,N_24540,N_24861);
nor UO_1191 (O_1191,N_24653,N_24890);
nand UO_1192 (O_1192,N_24569,N_24674);
nand UO_1193 (O_1193,N_24517,N_24797);
nor UO_1194 (O_1194,N_24966,N_24726);
nor UO_1195 (O_1195,N_24678,N_24816);
and UO_1196 (O_1196,N_24776,N_24981);
nor UO_1197 (O_1197,N_24970,N_24778);
xnor UO_1198 (O_1198,N_24818,N_24658);
and UO_1199 (O_1199,N_24882,N_24738);
nand UO_1200 (O_1200,N_24792,N_24712);
or UO_1201 (O_1201,N_24989,N_24567);
or UO_1202 (O_1202,N_24590,N_24625);
nand UO_1203 (O_1203,N_24889,N_24705);
nor UO_1204 (O_1204,N_24950,N_24546);
or UO_1205 (O_1205,N_24629,N_24747);
or UO_1206 (O_1206,N_24576,N_24501);
xor UO_1207 (O_1207,N_24522,N_24590);
nor UO_1208 (O_1208,N_24928,N_24568);
nor UO_1209 (O_1209,N_24939,N_24824);
or UO_1210 (O_1210,N_24524,N_24619);
nor UO_1211 (O_1211,N_24887,N_24625);
xnor UO_1212 (O_1212,N_24741,N_24993);
and UO_1213 (O_1213,N_24908,N_24521);
xor UO_1214 (O_1214,N_24920,N_24515);
nand UO_1215 (O_1215,N_24745,N_24601);
nand UO_1216 (O_1216,N_24574,N_24909);
and UO_1217 (O_1217,N_24574,N_24764);
nand UO_1218 (O_1218,N_24866,N_24862);
nor UO_1219 (O_1219,N_24701,N_24810);
and UO_1220 (O_1220,N_24834,N_24998);
or UO_1221 (O_1221,N_24940,N_24855);
nand UO_1222 (O_1222,N_24510,N_24800);
nand UO_1223 (O_1223,N_24765,N_24869);
nand UO_1224 (O_1224,N_24582,N_24837);
or UO_1225 (O_1225,N_24508,N_24943);
nand UO_1226 (O_1226,N_24915,N_24721);
nor UO_1227 (O_1227,N_24518,N_24564);
or UO_1228 (O_1228,N_24935,N_24660);
and UO_1229 (O_1229,N_24519,N_24692);
nor UO_1230 (O_1230,N_24951,N_24778);
nor UO_1231 (O_1231,N_24786,N_24698);
or UO_1232 (O_1232,N_24821,N_24559);
or UO_1233 (O_1233,N_24854,N_24608);
nand UO_1234 (O_1234,N_24779,N_24505);
and UO_1235 (O_1235,N_24543,N_24808);
nor UO_1236 (O_1236,N_24948,N_24587);
and UO_1237 (O_1237,N_24840,N_24575);
nor UO_1238 (O_1238,N_24719,N_24767);
nor UO_1239 (O_1239,N_24837,N_24719);
or UO_1240 (O_1240,N_24647,N_24621);
or UO_1241 (O_1241,N_24812,N_24573);
or UO_1242 (O_1242,N_24905,N_24794);
nor UO_1243 (O_1243,N_24915,N_24793);
nand UO_1244 (O_1244,N_24916,N_24528);
xnor UO_1245 (O_1245,N_24902,N_24802);
and UO_1246 (O_1246,N_24676,N_24907);
and UO_1247 (O_1247,N_24827,N_24949);
nand UO_1248 (O_1248,N_24889,N_24739);
or UO_1249 (O_1249,N_24927,N_24957);
and UO_1250 (O_1250,N_24730,N_24816);
xnor UO_1251 (O_1251,N_24605,N_24893);
and UO_1252 (O_1252,N_24685,N_24913);
xnor UO_1253 (O_1253,N_24770,N_24768);
and UO_1254 (O_1254,N_24887,N_24845);
xor UO_1255 (O_1255,N_24756,N_24981);
xor UO_1256 (O_1256,N_24511,N_24760);
nand UO_1257 (O_1257,N_24846,N_24556);
nor UO_1258 (O_1258,N_24559,N_24546);
nor UO_1259 (O_1259,N_24908,N_24769);
nand UO_1260 (O_1260,N_24952,N_24694);
or UO_1261 (O_1261,N_24954,N_24609);
xnor UO_1262 (O_1262,N_24867,N_24907);
or UO_1263 (O_1263,N_24849,N_24528);
xor UO_1264 (O_1264,N_24981,N_24555);
nor UO_1265 (O_1265,N_24601,N_24894);
or UO_1266 (O_1266,N_24943,N_24723);
nor UO_1267 (O_1267,N_24773,N_24646);
or UO_1268 (O_1268,N_24563,N_24710);
and UO_1269 (O_1269,N_24680,N_24634);
nor UO_1270 (O_1270,N_24703,N_24691);
and UO_1271 (O_1271,N_24788,N_24989);
or UO_1272 (O_1272,N_24908,N_24891);
nand UO_1273 (O_1273,N_24642,N_24803);
nand UO_1274 (O_1274,N_24849,N_24962);
or UO_1275 (O_1275,N_24794,N_24565);
or UO_1276 (O_1276,N_24607,N_24983);
nor UO_1277 (O_1277,N_24872,N_24880);
or UO_1278 (O_1278,N_24922,N_24736);
and UO_1279 (O_1279,N_24832,N_24553);
nand UO_1280 (O_1280,N_24649,N_24595);
nor UO_1281 (O_1281,N_24607,N_24619);
or UO_1282 (O_1282,N_24595,N_24821);
nor UO_1283 (O_1283,N_24510,N_24746);
and UO_1284 (O_1284,N_24733,N_24528);
and UO_1285 (O_1285,N_24738,N_24933);
nor UO_1286 (O_1286,N_24623,N_24608);
or UO_1287 (O_1287,N_24599,N_24704);
or UO_1288 (O_1288,N_24951,N_24767);
or UO_1289 (O_1289,N_24893,N_24626);
nor UO_1290 (O_1290,N_24538,N_24912);
nor UO_1291 (O_1291,N_24829,N_24734);
nor UO_1292 (O_1292,N_24890,N_24626);
and UO_1293 (O_1293,N_24874,N_24827);
nor UO_1294 (O_1294,N_24852,N_24646);
or UO_1295 (O_1295,N_24988,N_24645);
and UO_1296 (O_1296,N_24570,N_24585);
and UO_1297 (O_1297,N_24773,N_24739);
nand UO_1298 (O_1298,N_24800,N_24828);
xor UO_1299 (O_1299,N_24637,N_24572);
or UO_1300 (O_1300,N_24504,N_24900);
and UO_1301 (O_1301,N_24699,N_24691);
and UO_1302 (O_1302,N_24985,N_24711);
nor UO_1303 (O_1303,N_24699,N_24643);
xor UO_1304 (O_1304,N_24832,N_24756);
and UO_1305 (O_1305,N_24704,N_24978);
nor UO_1306 (O_1306,N_24793,N_24529);
xor UO_1307 (O_1307,N_24795,N_24909);
xnor UO_1308 (O_1308,N_24581,N_24935);
nor UO_1309 (O_1309,N_24939,N_24891);
nand UO_1310 (O_1310,N_24706,N_24516);
or UO_1311 (O_1311,N_24626,N_24647);
nor UO_1312 (O_1312,N_24590,N_24807);
or UO_1313 (O_1313,N_24943,N_24589);
nand UO_1314 (O_1314,N_24601,N_24619);
xor UO_1315 (O_1315,N_24514,N_24606);
nand UO_1316 (O_1316,N_24674,N_24580);
nand UO_1317 (O_1317,N_24864,N_24702);
and UO_1318 (O_1318,N_24930,N_24608);
and UO_1319 (O_1319,N_24622,N_24737);
and UO_1320 (O_1320,N_24578,N_24799);
nor UO_1321 (O_1321,N_24818,N_24750);
nand UO_1322 (O_1322,N_24890,N_24973);
nand UO_1323 (O_1323,N_24778,N_24705);
nor UO_1324 (O_1324,N_24945,N_24741);
nor UO_1325 (O_1325,N_24571,N_24574);
or UO_1326 (O_1326,N_24588,N_24880);
nor UO_1327 (O_1327,N_24942,N_24908);
nand UO_1328 (O_1328,N_24539,N_24894);
nor UO_1329 (O_1329,N_24685,N_24875);
nand UO_1330 (O_1330,N_24704,N_24694);
nand UO_1331 (O_1331,N_24646,N_24761);
nand UO_1332 (O_1332,N_24658,N_24526);
nand UO_1333 (O_1333,N_24548,N_24952);
xnor UO_1334 (O_1334,N_24776,N_24949);
or UO_1335 (O_1335,N_24957,N_24889);
or UO_1336 (O_1336,N_24818,N_24929);
nor UO_1337 (O_1337,N_24825,N_24673);
nor UO_1338 (O_1338,N_24624,N_24683);
or UO_1339 (O_1339,N_24662,N_24880);
xor UO_1340 (O_1340,N_24668,N_24857);
or UO_1341 (O_1341,N_24747,N_24953);
nand UO_1342 (O_1342,N_24785,N_24911);
xnor UO_1343 (O_1343,N_24929,N_24656);
nor UO_1344 (O_1344,N_24856,N_24507);
and UO_1345 (O_1345,N_24641,N_24508);
xnor UO_1346 (O_1346,N_24895,N_24872);
nor UO_1347 (O_1347,N_24984,N_24965);
nand UO_1348 (O_1348,N_24668,N_24540);
nor UO_1349 (O_1349,N_24781,N_24756);
xor UO_1350 (O_1350,N_24852,N_24716);
and UO_1351 (O_1351,N_24641,N_24823);
or UO_1352 (O_1352,N_24532,N_24728);
or UO_1353 (O_1353,N_24767,N_24772);
nor UO_1354 (O_1354,N_24919,N_24813);
xor UO_1355 (O_1355,N_24855,N_24535);
nor UO_1356 (O_1356,N_24694,N_24989);
and UO_1357 (O_1357,N_24803,N_24539);
or UO_1358 (O_1358,N_24695,N_24847);
xor UO_1359 (O_1359,N_24622,N_24701);
and UO_1360 (O_1360,N_24822,N_24950);
and UO_1361 (O_1361,N_24989,N_24568);
xnor UO_1362 (O_1362,N_24738,N_24506);
and UO_1363 (O_1363,N_24513,N_24689);
or UO_1364 (O_1364,N_24742,N_24571);
xnor UO_1365 (O_1365,N_24925,N_24916);
nor UO_1366 (O_1366,N_24527,N_24902);
nor UO_1367 (O_1367,N_24610,N_24890);
and UO_1368 (O_1368,N_24721,N_24939);
xnor UO_1369 (O_1369,N_24502,N_24795);
nor UO_1370 (O_1370,N_24951,N_24532);
and UO_1371 (O_1371,N_24582,N_24867);
xnor UO_1372 (O_1372,N_24772,N_24674);
xor UO_1373 (O_1373,N_24657,N_24896);
and UO_1374 (O_1374,N_24557,N_24846);
or UO_1375 (O_1375,N_24597,N_24540);
and UO_1376 (O_1376,N_24956,N_24525);
or UO_1377 (O_1377,N_24642,N_24768);
and UO_1378 (O_1378,N_24721,N_24749);
or UO_1379 (O_1379,N_24637,N_24682);
nor UO_1380 (O_1380,N_24897,N_24581);
nand UO_1381 (O_1381,N_24998,N_24902);
or UO_1382 (O_1382,N_24827,N_24546);
and UO_1383 (O_1383,N_24854,N_24862);
and UO_1384 (O_1384,N_24503,N_24502);
nor UO_1385 (O_1385,N_24793,N_24882);
nand UO_1386 (O_1386,N_24638,N_24504);
xor UO_1387 (O_1387,N_24961,N_24798);
and UO_1388 (O_1388,N_24678,N_24713);
nand UO_1389 (O_1389,N_24536,N_24629);
nor UO_1390 (O_1390,N_24752,N_24700);
nor UO_1391 (O_1391,N_24534,N_24717);
or UO_1392 (O_1392,N_24634,N_24869);
xor UO_1393 (O_1393,N_24532,N_24620);
nand UO_1394 (O_1394,N_24543,N_24842);
and UO_1395 (O_1395,N_24910,N_24634);
and UO_1396 (O_1396,N_24611,N_24970);
and UO_1397 (O_1397,N_24980,N_24677);
and UO_1398 (O_1398,N_24523,N_24756);
and UO_1399 (O_1399,N_24657,N_24652);
or UO_1400 (O_1400,N_24916,N_24926);
nor UO_1401 (O_1401,N_24741,N_24997);
and UO_1402 (O_1402,N_24982,N_24759);
or UO_1403 (O_1403,N_24533,N_24973);
and UO_1404 (O_1404,N_24703,N_24953);
or UO_1405 (O_1405,N_24630,N_24962);
and UO_1406 (O_1406,N_24859,N_24581);
nand UO_1407 (O_1407,N_24935,N_24698);
xnor UO_1408 (O_1408,N_24935,N_24757);
nand UO_1409 (O_1409,N_24570,N_24998);
xor UO_1410 (O_1410,N_24884,N_24839);
xnor UO_1411 (O_1411,N_24799,N_24636);
xor UO_1412 (O_1412,N_24542,N_24997);
and UO_1413 (O_1413,N_24769,N_24882);
or UO_1414 (O_1414,N_24532,N_24573);
or UO_1415 (O_1415,N_24828,N_24652);
or UO_1416 (O_1416,N_24768,N_24973);
or UO_1417 (O_1417,N_24846,N_24511);
nand UO_1418 (O_1418,N_24681,N_24547);
xor UO_1419 (O_1419,N_24678,N_24552);
and UO_1420 (O_1420,N_24809,N_24872);
nor UO_1421 (O_1421,N_24982,N_24995);
or UO_1422 (O_1422,N_24670,N_24554);
nand UO_1423 (O_1423,N_24595,N_24535);
or UO_1424 (O_1424,N_24697,N_24928);
or UO_1425 (O_1425,N_24761,N_24895);
xnor UO_1426 (O_1426,N_24954,N_24831);
or UO_1427 (O_1427,N_24964,N_24803);
nor UO_1428 (O_1428,N_24681,N_24952);
and UO_1429 (O_1429,N_24959,N_24813);
or UO_1430 (O_1430,N_24812,N_24960);
xnor UO_1431 (O_1431,N_24538,N_24833);
nor UO_1432 (O_1432,N_24927,N_24809);
nand UO_1433 (O_1433,N_24520,N_24752);
or UO_1434 (O_1434,N_24597,N_24562);
and UO_1435 (O_1435,N_24619,N_24921);
xor UO_1436 (O_1436,N_24817,N_24521);
or UO_1437 (O_1437,N_24520,N_24983);
nor UO_1438 (O_1438,N_24799,N_24848);
nor UO_1439 (O_1439,N_24995,N_24510);
nand UO_1440 (O_1440,N_24522,N_24647);
xnor UO_1441 (O_1441,N_24895,N_24773);
xor UO_1442 (O_1442,N_24654,N_24588);
nor UO_1443 (O_1443,N_24688,N_24729);
nand UO_1444 (O_1444,N_24896,N_24630);
nand UO_1445 (O_1445,N_24896,N_24521);
xnor UO_1446 (O_1446,N_24938,N_24747);
xor UO_1447 (O_1447,N_24875,N_24757);
and UO_1448 (O_1448,N_24659,N_24681);
and UO_1449 (O_1449,N_24974,N_24503);
and UO_1450 (O_1450,N_24531,N_24844);
nand UO_1451 (O_1451,N_24907,N_24806);
nor UO_1452 (O_1452,N_24882,N_24804);
or UO_1453 (O_1453,N_24834,N_24945);
nor UO_1454 (O_1454,N_24692,N_24735);
xor UO_1455 (O_1455,N_24925,N_24755);
nor UO_1456 (O_1456,N_24745,N_24538);
nand UO_1457 (O_1457,N_24578,N_24550);
and UO_1458 (O_1458,N_24946,N_24601);
or UO_1459 (O_1459,N_24841,N_24899);
nor UO_1460 (O_1460,N_24511,N_24581);
or UO_1461 (O_1461,N_24690,N_24699);
nor UO_1462 (O_1462,N_24814,N_24726);
nor UO_1463 (O_1463,N_24925,N_24660);
xnor UO_1464 (O_1464,N_24902,N_24944);
and UO_1465 (O_1465,N_24535,N_24988);
nand UO_1466 (O_1466,N_24836,N_24861);
nor UO_1467 (O_1467,N_24862,N_24630);
or UO_1468 (O_1468,N_24980,N_24631);
and UO_1469 (O_1469,N_24507,N_24858);
or UO_1470 (O_1470,N_24862,N_24725);
nor UO_1471 (O_1471,N_24840,N_24871);
xnor UO_1472 (O_1472,N_24882,N_24586);
and UO_1473 (O_1473,N_24763,N_24992);
xnor UO_1474 (O_1474,N_24832,N_24631);
nor UO_1475 (O_1475,N_24873,N_24968);
and UO_1476 (O_1476,N_24620,N_24862);
xor UO_1477 (O_1477,N_24631,N_24639);
xnor UO_1478 (O_1478,N_24735,N_24787);
xnor UO_1479 (O_1479,N_24657,N_24653);
and UO_1480 (O_1480,N_24591,N_24655);
nor UO_1481 (O_1481,N_24664,N_24789);
nand UO_1482 (O_1482,N_24518,N_24754);
nor UO_1483 (O_1483,N_24718,N_24907);
nand UO_1484 (O_1484,N_24861,N_24647);
xnor UO_1485 (O_1485,N_24838,N_24899);
and UO_1486 (O_1486,N_24596,N_24769);
nor UO_1487 (O_1487,N_24923,N_24742);
and UO_1488 (O_1488,N_24692,N_24847);
nand UO_1489 (O_1489,N_24770,N_24630);
nand UO_1490 (O_1490,N_24701,N_24647);
nor UO_1491 (O_1491,N_24953,N_24769);
or UO_1492 (O_1492,N_24713,N_24593);
and UO_1493 (O_1493,N_24990,N_24848);
or UO_1494 (O_1494,N_24820,N_24557);
or UO_1495 (O_1495,N_24812,N_24889);
nand UO_1496 (O_1496,N_24559,N_24944);
nor UO_1497 (O_1497,N_24689,N_24791);
and UO_1498 (O_1498,N_24775,N_24808);
nor UO_1499 (O_1499,N_24930,N_24898);
and UO_1500 (O_1500,N_24704,N_24858);
nand UO_1501 (O_1501,N_24855,N_24882);
xor UO_1502 (O_1502,N_24523,N_24888);
nor UO_1503 (O_1503,N_24529,N_24870);
nand UO_1504 (O_1504,N_24529,N_24902);
nor UO_1505 (O_1505,N_24592,N_24770);
nand UO_1506 (O_1506,N_24831,N_24862);
nand UO_1507 (O_1507,N_24817,N_24991);
or UO_1508 (O_1508,N_24840,N_24808);
and UO_1509 (O_1509,N_24568,N_24598);
nand UO_1510 (O_1510,N_24528,N_24794);
nor UO_1511 (O_1511,N_24719,N_24977);
nand UO_1512 (O_1512,N_24911,N_24863);
and UO_1513 (O_1513,N_24993,N_24769);
nand UO_1514 (O_1514,N_24636,N_24867);
xnor UO_1515 (O_1515,N_24859,N_24630);
nor UO_1516 (O_1516,N_24714,N_24666);
and UO_1517 (O_1517,N_24785,N_24704);
and UO_1518 (O_1518,N_24964,N_24683);
nand UO_1519 (O_1519,N_24911,N_24630);
nand UO_1520 (O_1520,N_24918,N_24877);
nand UO_1521 (O_1521,N_24724,N_24972);
or UO_1522 (O_1522,N_24926,N_24714);
and UO_1523 (O_1523,N_24671,N_24996);
nor UO_1524 (O_1524,N_24958,N_24708);
or UO_1525 (O_1525,N_24507,N_24581);
xnor UO_1526 (O_1526,N_24576,N_24927);
xor UO_1527 (O_1527,N_24964,N_24867);
xnor UO_1528 (O_1528,N_24511,N_24805);
nand UO_1529 (O_1529,N_24977,N_24792);
and UO_1530 (O_1530,N_24522,N_24855);
xnor UO_1531 (O_1531,N_24561,N_24722);
nand UO_1532 (O_1532,N_24642,N_24896);
or UO_1533 (O_1533,N_24578,N_24709);
and UO_1534 (O_1534,N_24583,N_24814);
and UO_1535 (O_1535,N_24745,N_24997);
and UO_1536 (O_1536,N_24870,N_24720);
nand UO_1537 (O_1537,N_24578,N_24645);
or UO_1538 (O_1538,N_24967,N_24721);
xor UO_1539 (O_1539,N_24786,N_24718);
nand UO_1540 (O_1540,N_24537,N_24928);
and UO_1541 (O_1541,N_24570,N_24909);
and UO_1542 (O_1542,N_24973,N_24808);
nor UO_1543 (O_1543,N_24779,N_24719);
xnor UO_1544 (O_1544,N_24621,N_24923);
and UO_1545 (O_1545,N_24630,N_24764);
nor UO_1546 (O_1546,N_24805,N_24581);
nor UO_1547 (O_1547,N_24955,N_24619);
nand UO_1548 (O_1548,N_24653,N_24552);
and UO_1549 (O_1549,N_24606,N_24563);
nor UO_1550 (O_1550,N_24672,N_24941);
nand UO_1551 (O_1551,N_24705,N_24750);
and UO_1552 (O_1552,N_24731,N_24864);
nor UO_1553 (O_1553,N_24940,N_24678);
xor UO_1554 (O_1554,N_24814,N_24912);
nand UO_1555 (O_1555,N_24915,N_24529);
nand UO_1556 (O_1556,N_24874,N_24508);
xnor UO_1557 (O_1557,N_24911,N_24646);
nor UO_1558 (O_1558,N_24791,N_24946);
or UO_1559 (O_1559,N_24664,N_24695);
xor UO_1560 (O_1560,N_24793,N_24844);
and UO_1561 (O_1561,N_24927,N_24636);
nor UO_1562 (O_1562,N_24820,N_24684);
nand UO_1563 (O_1563,N_24868,N_24788);
xor UO_1564 (O_1564,N_24581,N_24741);
and UO_1565 (O_1565,N_24640,N_24677);
nor UO_1566 (O_1566,N_24636,N_24508);
nand UO_1567 (O_1567,N_24851,N_24912);
nand UO_1568 (O_1568,N_24739,N_24752);
xor UO_1569 (O_1569,N_24584,N_24704);
or UO_1570 (O_1570,N_24791,N_24843);
xnor UO_1571 (O_1571,N_24877,N_24884);
nor UO_1572 (O_1572,N_24979,N_24897);
or UO_1573 (O_1573,N_24772,N_24808);
and UO_1574 (O_1574,N_24560,N_24686);
nand UO_1575 (O_1575,N_24666,N_24597);
nor UO_1576 (O_1576,N_24661,N_24612);
nor UO_1577 (O_1577,N_24733,N_24522);
nand UO_1578 (O_1578,N_24650,N_24606);
and UO_1579 (O_1579,N_24547,N_24513);
nor UO_1580 (O_1580,N_24989,N_24941);
xnor UO_1581 (O_1581,N_24902,N_24868);
xor UO_1582 (O_1582,N_24970,N_24991);
xor UO_1583 (O_1583,N_24929,N_24659);
and UO_1584 (O_1584,N_24555,N_24727);
and UO_1585 (O_1585,N_24631,N_24814);
nand UO_1586 (O_1586,N_24753,N_24550);
nor UO_1587 (O_1587,N_24568,N_24723);
and UO_1588 (O_1588,N_24609,N_24762);
and UO_1589 (O_1589,N_24521,N_24520);
or UO_1590 (O_1590,N_24763,N_24610);
nor UO_1591 (O_1591,N_24917,N_24716);
and UO_1592 (O_1592,N_24822,N_24834);
nor UO_1593 (O_1593,N_24647,N_24978);
nand UO_1594 (O_1594,N_24592,N_24567);
nand UO_1595 (O_1595,N_24998,N_24926);
nand UO_1596 (O_1596,N_24867,N_24528);
xor UO_1597 (O_1597,N_24975,N_24683);
nand UO_1598 (O_1598,N_24575,N_24915);
xor UO_1599 (O_1599,N_24601,N_24662);
nor UO_1600 (O_1600,N_24647,N_24684);
and UO_1601 (O_1601,N_24605,N_24742);
and UO_1602 (O_1602,N_24897,N_24900);
nand UO_1603 (O_1603,N_24700,N_24562);
nand UO_1604 (O_1604,N_24853,N_24902);
and UO_1605 (O_1605,N_24998,N_24832);
nand UO_1606 (O_1606,N_24946,N_24724);
and UO_1607 (O_1607,N_24759,N_24706);
nor UO_1608 (O_1608,N_24515,N_24791);
or UO_1609 (O_1609,N_24502,N_24903);
nor UO_1610 (O_1610,N_24701,N_24875);
xor UO_1611 (O_1611,N_24569,N_24725);
nand UO_1612 (O_1612,N_24725,N_24810);
and UO_1613 (O_1613,N_24953,N_24662);
xnor UO_1614 (O_1614,N_24570,N_24636);
xnor UO_1615 (O_1615,N_24578,N_24938);
and UO_1616 (O_1616,N_24812,N_24564);
or UO_1617 (O_1617,N_24926,N_24737);
nor UO_1618 (O_1618,N_24913,N_24592);
xor UO_1619 (O_1619,N_24663,N_24807);
or UO_1620 (O_1620,N_24745,N_24628);
and UO_1621 (O_1621,N_24793,N_24872);
nor UO_1622 (O_1622,N_24716,N_24687);
xnor UO_1623 (O_1623,N_24859,N_24638);
or UO_1624 (O_1624,N_24500,N_24933);
and UO_1625 (O_1625,N_24900,N_24902);
xor UO_1626 (O_1626,N_24922,N_24569);
and UO_1627 (O_1627,N_24631,N_24970);
or UO_1628 (O_1628,N_24551,N_24856);
nand UO_1629 (O_1629,N_24667,N_24861);
and UO_1630 (O_1630,N_24634,N_24674);
and UO_1631 (O_1631,N_24717,N_24932);
and UO_1632 (O_1632,N_24585,N_24889);
nand UO_1633 (O_1633,N_24555,N_24777);
nand UO_1634 (O_1634,N_24696,N_24908);
xnor UO_1635 (O_1635,N_24729,N_24605);
or UO_1636 (O_1636,N_24996,N_24642);
or UO_1637 (O_1637,N_24540,N_24651);
or UO_1638 (O_1638,N_24604,N_24510);
and UO_1639 (O_1639,N_24518,N_24833);
xor UO_1640 (O_1640,N_24922,N_24688);
or UO_1641 (O_1641,N_24650,N_24855);
xor UO_1642 (O_1642,N_24951,N_24829);
nand UO_1643 (O_1643,N_24667,N_24929);
and UO_1644 (O_1644,N_24665,N_24878);
and UO_1645 (O_1645,N_24509,N_24953);
nor UO_1646 (O_1646,N_24891,N_24663);
and UO_1647 (O_1647,N_24567,N_24606);
and UO_1648 (O_1648,N_24624,N_24881);
nand UO_1649 (O_1649,N_24961,N_24750);
xor UO_1650 (O_1650,N_24903,N_24550);
xor UO_1651 (O_1651,N_24863,N_24640);
nand UO_1652 (O_1652,N_24809,N_24873);
nand UO_1653 (O_1653,N_24613,N_24770);
nor UO_1654 (O_1654,N_24660,N_24962);
or UO_1655 (O_1655,N_24890,N_24956);
nor UO_1656 (O_1656,N_24855,N_24959);
nand UO_1657 (O_1657,N_24931,N_24838);
nor UO_1658 (O_1658,N_24961,N_24871);
nand UO_1659 (O_1659,N_24989,N_24535);
xor UO_1660 (O_1660,N_24822,N_24594);
nand UO_1661 (O_1661,N_24834,N_24718);
and UO_1662 (O_1662,N_24668,N_24848);
or UO_1663 (O_1663,N_24738,N_24993);
nand UO_1664 (O_1664,N_24965,N_24630);
nand UO_1665 (O_1665,N_24985,N_24885);
or UO_1666 (O_1666,N_24991,N_24999);
or UO_1667 (O_1667,N_24663,N_24700);
nor UO_1668 (O_1668,N_24964,N_24860);
or UO_1669 (O_1669,N_24543,N_24973);
and UO_1670 (O_1670,N_24550,N_24778);
nor UO_1671 (O_1671,N_24553,N_24754);
and UO_1672 (O_1672,N_24566,N_24754);
and UO_1673 (O_1673,N_24540,N_24940);
nor UO_1674 (O_1674,N_24973,N_24784);
and UO_1675 (O_1675,N_24592,N_24722);
nor UO_1676 (O_1676,N_24684,N_24665);
and UO_1677 (O_1677,N_24763,N_24527);
nor UO_1678 (O_1678,N_24974,N_24975);
nor UO_1679 (O_1679,N_24626,N_24965);
nor UO_1680 (O_1680,N_24874,N_24686);
xnor UO_1681 (O_1681,N_24549,N_24716);
xnor UO_1682 (O_1682,N_24748,N_24564);
and UO_1683 (O_1683,N_24967,N_24802);
nand UO_1684 (O_1684,N_24689,N_24532);
and UO_1685 (O_1685,N_24749,N_24617);
or UO_1686 (O_1686,N_24935,N_24964);
nand UO_1687 (O_1687,N_24881,N_24884);
nor UO_1688 (O_1688,N_24652,N_24867);
nor UO_1689 (O_1689,N_24684,N_24747);
nor UO_1690 (O_1690,N_24870,N_24801);
and UO_1691 (O_1691,N_24961,N_24940);
xnor UO_1692 (O_1692,N_24775,N_24796);
and UO_1693 (O_1693,N_24809,N_24756);
nor UO_1694 (O_1694,N_24732,N_24870);
nand UO_1695 (O_1695,N_24547,N_24810);
nand UO_1696 (O_1696,N_24796,N_24669);
and UO_1697 (O_1697,N_24944,N_24653);
nor UO_1698 (O_1698,N_24687,N_24601);
nand UO_1699 (O_1699,N_24510,N_24664);
xor UO_1700 (O_1700,N_24753,N_24705);
or UO_1701 (O_1701,N_24891,N_24788);
xor UO_1702 (O_1702,N_24712,N_24627);
and UO_1703 (O_1703,N_24645,N_24975);
nor UO_1704 (O_1704,N_24943,N_24882);
or UO_1705 (O_1705,N_24995,N_24575);
and UO_1706 (O_1706,N_24575,N_24663);
xnor UO_1707 (O_1707,N_24970,N_24615);
or UO_1708 (O_1708,N_24875,N_24841);
xnor UO_1709 (O_1709,N_24546,N_24771);
xnor UO_1710 (O_1710,N_24906,N_24507);
and UO_1711 (O_1711,N_24567,N_24587);
or UO_1712 (O_1712,N_24775,N_24886);
nand UO_1713 (O_1713,N_24813,N_24567);
nand UO_1714 (O_1714,N_24822,N_24920);
and UO_1715 (O_1715,N_24680,N_24927);
xnor UO_1716 (O_1716,N_24939,N_24566);
nor UO_1717 (O_1717,N_24513,N_24549);
and UO_1718 (O_1718,N_24883,N_24626);
nor UO_1719 (O_1719,N_24884,N_24821);
or UO_1720 (O_1720,N_24942,N_24666);
xor UO_1721 (O_1721,N_24787,N_24718);
or UO_1722 (O_1722,N_24616,N_24810);
nor UO_1723 (O_1723,N_24543,N_24724);
or UO_1724 (O_1724,N_24519,N_24569);
and UO_1725 (O_1725,N_24890,N_24970);
and UO_1726 (O_1726,N_24597,N_24880);
nor UO_1727 (O_1727,N_24852,N_24658);
xnor UO_1728 (O_1728,N_24802,N_24586);
nor UO_1729 (O_1729,N_24529,N_24893);
nor UO_1730 (O_1730,N_24509,N_24835);
xor UO_1731 (O_1731,N_24722,N_24593);
xnor UO_1732 (O_1732,N_24557,N_24571);
or UO_1733 (O_1733,N_24955,N_24644);
and UO_1734 (O_1734,N_24684,N_24597);
and UO_1735 (O_1735,N_24977,N_24693);
and UO_1736 (O_1736,N_24579,N_24685);
xnor UO_1737 (O_1737,N_24810,N_24628);
nor UO_1738 (O_1738,N_24656,N_24503);
and UO_1739 (O_1739,N_24670,N_24524);
nand UO_1740 (O_1740,N_24895,N_24843);
and UO_1741 (O_1741,N_24872,N_24986);
xnor UO_1742 (O_1742,N_24858,N_24941);
nand UO_1743 (O_1743,N_24643,N_24511);
or UO_1744 (O_1744,N_24790,N_24999);
nor UO_1745 (O_1745,N_24709,N_24790);
xor UO_1746 (O_1746,N_24791,N_24553);
nor UO_1747 (O_1747,N_24666,N_24835);
nand UO_1748 (O_1748,N_24971,N_24984);
or UO_1749 (O_1749,N_24626,N_24658);
nand UO_1750 (O_1750,N_24597,N_24720);
nand UO_1751 (O_1751,N_24701,N_24835);
or UO_1752 (O_1752,N_24501,N_24788);
nand UO_1753 (O_1753,N_24630,N_24743);
nand UO_1754 (O_1754,N_24636,N_24868);
nor UO_1755 (O_1755,N_24610,N_24666);
xnor UO_1756 (O_1756,N_24603,N_24805);
nor UO_1757 (O_1757,N_24894,N_24983);
nand UO_1758 (O_1758,N_24900,N_24759);
xnor UO_1759 (O_1759,N_24958,N_24515);
nand UO_1760 (O_1760,N_24535,N_24550);
or UO_1761 (O_1761,N_24535,N_24558);
nor UO_1762 (O_1762,N_24896,N_24780);
or UO_1763 (O_1763,N_24937,N_24970);
nor UO_1764 (O_1764,N_24573,N_24843);
nand UO_1765 (O_1765,N_24956,N_24789);
nand UO_1766 (O_1766,N_24768,N_24517);
xnor UO_1767 (O_1767,N_24510,N_24992);
nand UO_1768 (O_1768,N_24913,N_24664);
xor UO_1769 (O_1769,N_24698,N_24587);
and UO_1770 (O_1770,N_24640,N_24802);
xor UO_1771 (O_1771,N_24516,N_24857);
nor UO_1772 (O_1772,N_24617,N_24711);
nand UO_1773 (O_1773,N_24795,N_24536);
nor UO_1774 (O_1774,N_24739,N_24615);
xor UO_1775 (O_1775,N_24550,N_24836);
and UO_1776 (O_1776,N_24606,N_24929);
and UO_1777 (O_1777,N_24900,N_24809);
nand UO_1778 (O_1778,N_24834,N_24565);
xor UO_1779 (O_1779,N_24990,N_24811);
xor UO_1780 (O_1780,N_24796,N_24767);
nand UO_1781 (O_1781,N_24751,N_24683);
nor UO_1782 (O_1782,N_24835,N_24718);
xor UO_1783 (O_1783,N_24844,N_24557);
and UO_1784 (O_1784,N_24592,N_24786);
and UO_1785 (O_1785,N_24973,N_24737);
nor UO_1786 (O_1786,N_24579,N_24916);
nor UO_1787 (O_1787,N_24694,N_24879);
xnor UO_1788 (O_1788,N_24710,N_24753);
xor UO_1789 (O_1789,N_24842,N_24660);
xor UO_1790 (O_1790,N_24716,N_24656);
or UO_1791 (O_1791,N_24613,N_24882);
and UO_1792 (O_1792,N_24904,N_24763);
nor UO_1793 (O_1793,N_24666,N_24662);
or UO_1794 (O_1794,N_24549,N_24899);
nand UO_1795 (O_1795,N_24799,N_24906);
or UO_1796 (O_1796,N_24508,N_24583);
xnor UO_1797 (O_1797,N_24856,N_24689);
nand UO_1798 (O_1798,N_24816,N_24969);
nor UO_1799 (O_1799,N_24962,N_24718);
nand UO_1800 (O_1800,N_24802,N_24977);
or UO_1801 (O_1801,N_24601,N_24873);
xor UO_1802 (O_1802,N_24512,N_24810);
or UO_1803 (O_1803,N_24635,N_24518);
nand UO_1804 (O_1804,N_24639,N_24736);
and UO_1805 (O_1805,N_24622,N_24649);
nand UO_1806 (O_1806,N_24591,N_24597);
or UO_1807 (O_1807,N_24957,N_24589);
or UO_1808 (O_1808,N_24588,N_24688);
or UO_1809 (O_1809,N_24835,N_24854);
xor UO_1810 (O_1810,N_24761,N_24801);
or UO_1811 (O_1811,N_24889,N_24606);
nor UO_1812 (O_1812,N_24862,N_24798);
or UO_1813 (O_1813,N_24954,N_24660);
nor UO_1814 (O_1814,N_24690,N_24796);
nand UO_1815 (O_1815,N_24744,N_24516);
xnor UO_1816 (O_1816,N_24971,N_24556);
nor UO_1817 (O_1817,N_24598,N_24520);
nand UO_1818 (O_1818,N_24555,N_24607);
nor UO_1819 (O_1819,N_24824,N_24954);
or UO_1820 (O_1820,N_24746,N_24648);
nor UO_1821 (O_1821,N_24971,N_24896);
xnor UO_1822 (O_1822,N_24930,N_24721);
nand UO_1823 (O_1823,N_24595,N_24645);
and UO_1824 (O_1824,N_24814,N_24677);
xnor UO_1825 (O_1825,N_24626,N_24610);
or UO_1826 (O_1826,N_24692,N_24855);
nand UO_1827 (O_1827,N_24945,N_24567);
xor UO_1828 (O_1828,N_24578,N_24956);
nand UO_1829 (O_1829,N_24757,N_24710);
and UO_1830 (O_1830,N_24999,N_24885);
nand UO_1831 (O_1831,N_24702,N_24706);
xor UO_1832 (O_1832,N_24667,N_24578);
nor UO_1833 (O_1833,N_24522,N_24885);
nor UO_1834 (O_1834,N_24536,N_24694);
and UO_1835 (O_1835,N_24961,N_24996);
xnor UO_1836 (O_1836,N_24907,N_24854);
and UO_1837 (O_1837,N_24844,N_24622);
nor UO_1838 (O_1838,N_24755,N_24780);
nand UO_1839 (O_1839,N_24574,N_24512);
nand UO_1840 (O_1840,N_24515,N_24768);
nand UO_1841 (O_1841,N_24749,N_24846);
nand UO_1842 (O_1842,N_24729,N_24653);
nor UO_1843 (O_1843,N_24925,N_24638);
xor UO_1844 (O_1844,N_24720,N_24639);
nor UO_1845 (O_1845,N_24534,N_24989);
xor UO_1846 (O_1846,N_24933,N_24736);
nor UO_1847 (O_1847,N_24535,N_24676);
and UO_1848 (O_1848,N_24980,N_24645);
nor UO_1849 (O_1849,N_24875,N_24500);
xor UO_1850 (O_1850,N_24755,N_24984);
and UO_1851 (O_1851,N_24698,N_24653);
or UO_1852 (O_1852,N_24679,N_24899);
and UO_1853 (O_1853,N_24916,N_24995);
nand UO_1854 (O_1854,N_24751,N_24924);
xor UO_1855 (O_1855,N_24909,N_24771);
or UO_1856 (O_1856,N_24619,N_24507);
or UO_1857 (O_1857,N_24840,N_24600);
or UO_1858 (O_1858,N_24587,N_24504);
nand UO_1859 (O_1859,N_24619,N_24817);
xnor UO_1860 (O_1860,N_24754,N_24997);
nand UO_1861 (O_1861,N_24636,N_24738);
nand UO_1862 (O_1862,N_24790,N_24543);
and UO_1863 (O_1863,N_24661,N_24705);
nand UO_1864 (O_1864,N_24602,N_24718);
nor UO_1865 (O_1865,N_24735,N_24624);
or UO_1866 (O_1866,N_24921,N_24714);
and UO_1867 (O_1867,N_24535,N_24753);
nor UO_1868 (O_1868,N_24997,N_24929);
nor UO_1869 (O_1869,N_24931,N_24847);
nand UO_1870 (O_1870,N_24918,N_24789);
or UO_1871 (O_1871,N_24881,N_24847);
nand UO_1872 (O_1872,N_24814,N_24699);
nor UO_1873 (O_1873,N_24892,N_24907);
xnor UO_1874 (O_1874,N_24726,N_24941);
and UO_1875 (O_1875,N_24865,N_24680);
or UO_1876 (O_1876,N_24856,N_24946);
xnor UO_1877 (O_1877,N_24737,N_24770);
nor UO_1878 (O_1878,N_24663,N_24897);
nor UO_1879 (O_1879,N_24573,N_24588);
nand UO_1880 (O_1880,N_24610,N_24762);
or UO_1881 (O_1881,N_24887,N_24830);
and UO_1882 (O_1882,N_24790,N_24730);
nor UO_1883 (O_1883,N_24728,N_24965);
xnor UO_1884 (O_1884,N_24888,N_24775);
xnor UO_1885 (O_1885,N_24796,N_24935);
xor UO_1886 (O_1886,N_24778,N_24553);
and UO_1887 (O_1887,N_24998,N_24571);
xor UO_1888 (O_1888,N_24875,N_24664);
and UO_1889 (O_1889,N_24812,N_24624);
or UO_1890 (O_1890,N_24521,N_24857);
nand UO_1891 (O_1891,N_24672,N_24792);
nand UO_1892 (O_1892,N_24687,N_24561);
nor UO_1893 (O_1893,N_24761,N_24664);
and UO_1894 (O_1894,N_24901,N_24621);
xor UO_1895 (O_1895,N_24579,N_24856);
nand UO_1896 (O_1896,N_24897,N_24594);
and UO_1897 (O_1897,N_24506,N_24844);
nor UO_1898 (O_1898,N_24996,N_24508);
nand UO_1899 (O_1899,N_24960,N_24629);
and UO_1900 (O_1900,N_24960,N_24950);
and UO_1901 (O_1901,N_24578,N_24525);
xor UO_1902 (O_1902,N_24857,N_24747);
nor UO_1903 (O_1903,N_24683,N_24699);
nor UO_1904 (O_1904,N_24581,N_24596);
nor UO_1905 (O_1905,N_24967,N_24646);
nand UO_1906 (O_1906,N_24935,N_24893);
nand UO_1907 (O_1907,N_24779,N_24748);
nand UO_1908 (O_1908,N_24940,N_24762);
or UO_1909 (O_1909,N_24641,N_24517);
xor UO_1910 (O_1910,N_24741,N_24793);
nor UO_1911 (O_1911,N_24780,N_24918);
xor UO_1912 (O_1912,N_24897,N_24883);
or UO_1913 (O_1913,N_24764,N_24826);
nor UO_1914 (O_1914,N_24946,N_24614);
or UO_1915 (O_1915,N_24815,N_24591);
nor UO_1916 (O_1916,N_24890,N_24587);
or UO_1917 (O_1917,N_24600,N_24823);
and UO_1918 (O_1918,N_24821,N_24758);
xor UO_1919 (O_1919,N_24535,N_24701);
and UO_1920 (O_1920,N_24649,N_24990);
nand UO_1921 (O_1921,N_24630,N_24875);
or UO_1922 (O_1922,N_24641,N_24500);
xnor UO_1923 (O_1923,N_24652,N_24668);
and UO_1924 (O_1924,N_24730,N_24961);
nor UO_1925 (O_1925,N_24869,N_24572);
nor UO_1926 (O_1926,N_24871,N_24562);
and UO_1927 (O_1927,N_24897,N_24969);
nand UO_1928 (O_1928,N_24782,N_24851);
xnor UO_1929 (O_1929,N_24883,N_24639);
xor UO_1930 (O_1930,N_24889,N_24823);
or UO_1931 (O_1931,N_24718,N_24573);
nand UO_1932 (O_1932,N_24958,N_24898);
or UO_1933 (O_1933,N_24644,N_24908);
or UO_1934 (O_1934,N_24896,N_24828);
nand UO_1935 (O_1935,N_24959,N_24509);
xor UO_1936 (O_1936,N_24696,N_24756);
nor UO_1937 (O_1937,N_24562,N_24917);
or UO_1938 (O_1938,N_24859,N_24834);
nor UO_1939 (O_1939,N_24971,N_24830);
xor UO_1940 (O_1940,N_24796,N_24961);
nor UO_1941 (O_1941,N_24541,N_24762);
xor UO_1942 (O_1942,N_24630,N_24979);
nor UO_1943 (O_1943,N_24674,N_24854);
nand UO_1944 (O_1944,N_24777,N_24922);
nor UO_1945 (O_1945,N_24974,N_24532);
nand UO_1946 (O_1946,N_24809,N_24799);
nor UO_1947 (O_1947,N_24544,N_24858);
or UO_1948 (O_1948,N_24551,N_24929);
or UO_1949 (O_1949,N_24596,N_24523);
or UO_1950 (O_1950,N_24819,N_24566);
xnor UO_1951 (O_1951,N_24531,N_24594);
nand UO_1952 (O_1952,N_24853,N_24986);
nand UO_1953 (O_1953,N_24876,N_24974);
or UO_1954 (O_1954,N_24858,N_24693);
xor UO_1955 (O_1955,N_24875,N_24695);
nor UO_1956 (O_1956,N_24636,N_24624);
or UO_1957 (O_1957,N_24825,N_24668);
or UO_1958 (O_1958,N_24643,N_24969);
nand UO_1959 (O_1959,N_24506,N_24557);
or UO_1960 (O_1960,N_24796,N_24673);
nor UO_1961 (O_1961,N_24903,N_24973);
and UO_1962 (O_1962,N_24797,N_24595);
xnor UO_1963 (O_1963,N_24937,N_24786);
and UO_1964 (O_1964,N_24702,N_24858);
xor UO_1965 (O_1965,N_24679,N_24959);
nor UO_1966 (O_1966,N_24831,N_24739);
and UO_1967 (O_1967,N_24828,N_24953);
nor UO_1968 (O_1968,N_24981,N_24649);
xor UO_1969 (O_1969,N_24605,N_24580);
nand UO_1970 (O_1970,N_24561,N_24921);
nor UO_1971 (O_1971,N_24867,N_24963);
or UO_1972 (O_1972,N_24571,N_24625);
and UO_1973 (O_1973,N_24699,N_24539);
nand UO_1974 (O_1974,N_24984,N_24895);
xnor UO_1975 (O_1975,N_24845,N_24893);
nand UO_1976 (O_1976,N_24743,N_24824);
and UO_1977 (O_1977,N_24666,N_24922);
nor UO_1978 (O_1978,N_24941,N_24852);
and UO_1979 (O_1979,N_24674,N_24727);
nor UO_1980 (O_1980,N_24576,N_24633);
nand UO_1981 (O_1981,N_24573,N_24550);
and UO_1982 (O_1982,N_24779,N_24638);
and UO_1983 (O_1983,N_24615,N_24671);
nand UO_1984 (O_1984,N_24823,N_24542);
nor UO_1985 (O_1985,N_24867,N_24943);
nand UO_1986 (O_1986,N_24908,N_24848);
and UO_1987 (O_1987,N_24519,N_24830);
nand UO_1988 (O_1988,N_24662,N_24945);
nand UO_1989 (O_1989,N_24682,N_24711);
nand UO_1990 (O_1990,N_24542,N_24606);
xor UO_1991 (O_1991,N_24512,N_24878);
nor UO_1992 (O_1992,N_24719,N_24551);
nand UO_1993 (O_1993,N_24710,N_24517);
and UO_1994 (O_1994,N_24973,N_24557);
xor UO_1995 (O_1995,N_24999,N_24579);
or UO_1996 (O_1996,N_24987,N_24610);
and UO_1997 (O_1997,N_24621,N_24983);
nor UO_1998 (O_1998,N_24661,N_24635);
nand UO_1999 (O_1999,N_24881,N_24529);
and UO_2000 (O_2000,N_24958,N_24562);
or UO_2001 (O_2001,N_24657,N_24519);
xnor UO_2002 (O_2002,N_24568,N_24520);
xnor UO_2003 (O_2003,N_24883,N_24612);
or UO_2004 (O_2004,N_24547,N_24591);
nor UO_2005 (O_2005,N_24820,N_24830);
nand UO_2006 (O_2006,N_24789,N_24729);
nand UO_2007 (O_2007,N_24650,N_24871);
and UO_2008 (O_2008,N_24578,N_24788);
xor UO_2009 (O_2009,N_24792,N_24976);
nor UO_2010 (O_2010,N_24668,N_24858);
nand UO_2011 (O_2011,N_24751,N_24729);
nor UO_2012 (O_2012,N_24850,N_24856);
xnor UO_2013 (O_2013,N_24793,N_24710);
or UO_2014 (O_2014,N_24593,N_24650);
or UO_2015 (O_2015,N_24867,N_24959);
xor UO_2016 (O_2016,N_24977,N_24630);
nor UO_2017 (O_2017,N_24688,N_24648);
or UO_2018 (O_2018,N_24634,N_24707);
or UO_2019 (O_2019,N_24801,N_24646);
or UO_2020 (O_2020,N_24896,N_24820);
xor UO_2021 (O_2021,N_24673,N_24773);
or UO_2022 (O_2022,N_24915,N_24551);
xor UO_2023 (O_2023,N_24730,N_24972);
and UO_2024 (O_2024,N_24910,N_24884);
or UO_2025 (O_2025,N_24541,N_24632);
xor UO_2026 (O_2026,N_24517,N_24989);
nand UO_2027 (O_2027,N_24733,N_24982);
or UO_2028 (O_2028,N_24985,N_24797);
xnor UO_2029 (O_2029,N_24557,N_24513);
and UO_2030 (O_2030,N_24788,N_24811);
xnor UO_2031 (O_2031,N_24524,N_24512);
nand UO_2032 (O_2032,N_24808,N_24975);
or UO_2033 (O_2033,N_24773,N_24698);
nor UO_2034 (O_2034,N_24945,N_24753);
and UO_2035 (O_2035,N_24537,N_24971);
or UO_2036 (O_2036,N_24813,N_24555);
nand UO_2037 (O_2037,N_24942,N_24895);
nand UO_2038 (O_2038,N_24692,N_24936);
xnor UO_2039 (O_2039,N_24542,N_24947);
nor UO_2040 (O_2040,N_24501,N_24808);
and UO_2041 (O_2041,N_24953,N_24552);
or UO_2042 (O_2042,N_24769,N_24692);
nor UO_2043 (O_2043,N_24648,N_24926);
nand UO_2044 (O_2044,N_24752,N_24742);
and UO_2045 (O_2045,N_24715,N_24702);
nand UO_2046 (O_2046,N_24665,N_24909);
and UO_2047 (O_2047,N_24819,N_24613);
nand UO_2048 (O_2048,N_24867,N_24752);
or UO_2049 (O_2049,N_24655,N_24666);
nand UO_2050 (O_2050,N_24929,N_24515);
xor UO_2051 (O_2051,N_24656,N_24721);
or UO_2052 (O_2052,N_24795,N_24596);
or UO_2053 (O_2053,N_24859,N_24629);
nor UO_2054 (O_2054,N_24911,N_24920);
or UO_2055 (O_2055,N_24677,N_24590);
xor UO_2056 (O_2056,N_24963,N_24528);
nand UO_2057 (O_2057,N_24711,N_24944);
or UO_2058 (O_2058,N_24861,N_24562);
or UO_2059 (O_2059,N_24838,N_24511);
nor UO_2060 (O_2060,N_24645,N_24772);
nand UO_2061 (O_2061,N_24974,N_24970);
and UO_2062 (O_2062,N_24882,N_24515);
or UO_2063 (O_2063,N_24628,N_24903);
and UO_2064 (O_2064,N_24981,N_24572);
xor UO_2065 (O_2065,N_24824,N_24874);
xor UO_2066 (O_2066,N_24808,N_24695);
or UO_2067 (O_2067,N_24838,N_24556);
or UO_2068 (O_2068,N_24706,N_24765);
xnor UO_2069 (O_2069,N_24994,N_24803);
or UO_2070 (O_2070,N_24667,N_24961);
nor UO_2071 (O_2071,N_24716,N_24846);
and UO_2072 (O_2072,N_24749,N_24592);
xnor UO_2073 (O_2073,N_24523,N_24882);
xor UO_2074 (O_2074,N_24828,N_24973);
nor UO_2075 (O_2075,N_24581,N_24816);
and UO_2076 (O_2076,N_24897,N_24517);
or UO_2077 (O_2077,N_24836,N_24524);
nand UO_2078 (O_2078,N_24765,N_24737);
nor UO_2079 (O_2079,N_24655,N_24569);
xnor UO_2080 (O_2080,N_24586,N_24963);
xnor UO_2081 (O_2081,N_24574,N_24992);
and UO_2082 (O_2082,N_24941,N_24925);
nand UO_2083 (O_2083,N_24800,N_24627);
xor UO_2084 (O_2084,N_24999,N_24986);
nand UO_2085 (O_2085,N_24974,N_24684);
nand UO_2086 (O_2086,N_24679,N_24997);
nand UO_2087 (O_2087,N_24701,N_24587);
and UO_2088 (O_2088,N_24947,N_24823);
and UO_2089 (O_2089,N_24527,N_24655);
or UO_2090 (O_2090,N_24513,N_24979);
and UO_2091 (O_2091,N_24694,N_24599);
xnor UO_2092 (O_2092,N_24530,N_24906);
nand UO_2093 (O_2093,N_24695,N_24513);
or UO_2094 (O_2094,N_24752,N_24617);
xor UO_2095 (O_2095,N_24811,N_24660);
nor UO_2096 (O_2096,N_24834,N_24860);
nor UO_2097 (O_2097,N_24881,N_24500);
nand UO_2098 (O_2098,N_24977,N_24507);
xnor UO_2099 (O_2099,N_24820,N_24910);
xnor UO_2100 (O_2100,N_24932,N_24636);
nand UO_2101 (O_2101,N_24897,N_24917);
nand UO_2102 (O_2102,N_24588,N_24835);
nor UO_2103 (O_2103,N_24845,N_24988);
xnor UO_2104 (O_2104,N_24901,N_24752);
or UO_2105 (O_2105,N_24848,N_24740);
nand UO_2106 (O_2106,N_24949,N_24984);
and UO_2107 (O_2107,N_24643,N_24845);
or UO_2108 (O_2108,N_24789,N_24690);
nand UO_2109 (O_2109,N_24946,N_24833);
and UO_2110 (O_2110,N_24932,N_24690);
and UO_2111 (O_2111,N_24512,N_24534);
xor UO_2112 (O_2112,N_24875,N_24707);
nand UO_2113 (O_2113,N_24725,N_24522);
nand UO_2114 (O_2114,N_24520,N_24823);
nand UO_2115 (O_2115,N_24633,N_24729);
nor UO_2116 (O_2116,N_24822,N_24760);
xor UO_2117 (O_2117,N_24806,N_24964);
nor UO_2118 (O_2118,N_24746,N_24664);
nand UO_2119 (O_2119,N_24646,N_24838);
xor UO_2120 (O_2120,N_24827,N_24616);
and UO_2121 (O_2121,N_24552,N_24903);
nand UO_2122 (O_2122,N_24740,N_24645);
and UO_2123 (O_2123,N_24633,N_24975);
nor UO_2124 (O_2124,N_24796,N_24729);
xor UO_2125 (O_2125,N_24575,N_24621);
nor UO_2126 (O_2126,N_24829,N_24804);
nand UO_2127 (O_2127,N_24523,N_24597);
nor UO_2128 (O_2128,N_24866,N_24835);
nand UO_2129 (O_2129,N_24942,N_24675);
nor UO_2130 (O_2130,N_24764,N_24778);
nor UO_2131 (O_2131,N_24793,N_24918);
nand UO_2132 (O_2132,N_24926,N_24888);
and UO_2133 (O_2133,N_24556,N_24710);
or UO_2134 (O_2134,N_24578,N_24898);
nand UO_2135 (O_2135,N_24627,N_24732);
nor UO_2136 (O_2136,N_24976,N_24968);
or UO_2137 (O_2137,N_24920,N_24659);
and UO_2138 (O_2138,N_24921,N_24585);
and UO_2139 (O_2139,N_24786,N_24818);
nor UO_2140 (O_2140,N_24760,N_24999);
nand UO_2141 (O_2141,N_24819,N_24963);
and UO_2142 (O_2142,N_24605,N_24697);
and UO_2143 (O_2143,N_24797,N_24744);
xnor UO_2144 (O_2144,N_24991,N_24615);
nand UO_2145 (O_2145,N_24682,N_24884);
nor UO_2146 (O_2146,N_24999,N_24965);
and UO_2147 (O_2147,N_24535,N_24756);
nor UO_2148 (O_2148,N_24765,N_24625);
or UO_2149 (O_2149,N_24980,N_24947);
xor UO_2150 (O_2150,N_24552,N_24573);
nor UO_2151 (O_2151,N_24833,N_24960);
xor UO_2152 (O_2152,N_24675,N_24938);
nor UO_2153 (O_2153,N_24510,N_24553);
nor UO_2154 (O_2154,N_24588,N_24946);
xnor UO_2155 (O_2155,N_24587,N_24788);
xnor UO_2156 (O_2156,N_24951,N_24869);
or UO_2157 (O_2157,N_24528,N_24716);
or UO_2158 (O_2158,N_24970,N_24572);
and UO_2159 (O_2159,N_24927,N_24602);
nor UO_2160 (O_2160,N_24634,N_24519);
nor UO_2161 (O_2161,N_24819,N_24702);
xnor UO_2162 (O_2162,N_24723,N_24775);
nor UO_2163 (O_2163,N_24971,N_24763);
xor UO_2164 (O_2164,N_24615,N_24826);
nand UO_2165 (O_2165,N_24788,N_24987);
xor UO_2166 (O_2166,N_24501,N_24512);
nor UO_2167 (O_2167,N_24502,N_24835);
and UO_2168 (O_2168,N_24682,N_24714);
nor UO_2169 (O_2169,N_24523,N_24853);
xnor UO_2170 (O_2170,N_24675,N_24792);
and UO_2171 (O_2171,N_24538,N_24888);
or UO_2172 (O_2172,N_24710,N_24885);
or UO_2173 (O_2173,N_24679,N_24975);
or UO_2174 (O_2174,N_24946,N_24837);
and UO_2175 (O_2175,N_24991,N_24945);
nor UO_2176 (O_2176,N_24979,N_24825);
nor UO_2177 (O_2177,N_24670,N_24535);
and UO_2178 (O_2178,N_24795,N_24745);
nor UO_2179 (O_2179,N_24861,N_24653);
nand UO_2180 (O_2180,N_24822,N_24545);
or UO_2181 (O_2181,N_24780,N_24621);
or UO_2182 (O_2182,N_24893,N_24513);
nand UO_2183 (O_2183,N_24567,N_24865);
nor UO_2184 (O_2184,N_24920,N_24877);
nor UO_2185 (O_2185,N_24899,N_24811);
and UO_2186 (O_2186,N_24797,N_24518);
nand UO_2187 (O_2187,N_24775,N_24978);
xor UO_2188 (O_2188,N_24874,N_24610);
and UO_2189 (O_2189,N_24839,N_24567);
nor UO_2190 (O_2190,N_24774,N_24859);
nor UO_2191 (O_2191,N_24665,N_24633);
or UO_2192 (O_2192,N_24668,N_24826);
and UO_2193 (O_2193,N_24690,N_24592);
and UO_2194 (O_2194,N_24987,N_24761);
xnor UO_2195 (O_2195,N_24709,N_24608);
nand UO_2196 (O_2196,N_24937,N_24502);
nor UO_2197 (O_2197,N_24938,N_24983);
and UO_2198 (O_2198,N_24933,N_24792);
nor UO_2199 (O_2199,N_24793,N_24797);
and UO_2200 (O_2200,N_24532,N_24509);
or UO_2201 (O_2201,N_24812,N_24899);
or UO_2202 (O_2202,N_24850,N_24599);
and UO_2203 (O_2203,N_24506,N_24603);
nor UO_2204 (O_2204,N_24920,N_24757);
nor UO_2205 (O_2205,N_24507,N_24834);
and UO_2206 (O_2206,N_24695,N_24886);
nand UO_2207 (O_2207,N_24768,N_24604);
xnor UO_2208 (O_2208,N_24684,N_24926);
nor UO_2209 (O_2209,N_24994,N_24923);
and UO_2210 (O_2210,N_24978,N_24795);
and UO_2211 (O_2211,N_24975,N_24884);
nand UO_2212 (O_2212,N_24556,N_24560);
xor UO_2213 (O_2213,N_24775,N_24719);
nor UO_2214 (O_2214,N_24563,N_24573);
nand UO_2215 (O_2215,N_24948,N_24917);
or UO_2216 (O_2216,N_24837,N_24664);
and UO_2217 (O_2217,N_24834,N_24881);
xnor UO_2218 (O_2218,N_24903,N_24666);
nor UO_2219 (O_2219,N_24641,N_24509);
and UO_2220 (O_2220,N_24736,N_24668);
xnor UO_2221 (O_2221,N_24781,N_24951);
xnor UO_2222 (O_2222,N_24779,N_24827);
and UO_2223 (O_2223,N_24797,N_24865);
nor UO_2224 (O_2224,N_24973,N_24876);
nor UO_2225 (O_2225,N_24606,N_24660);
and UO_2226 (O_2226,N_24750,N_24639);
or UO_2227 (O_2227,N_24930,N_24539);
xor UO_2228 (O_2228,N_24813,N_24881);
and UO_2229 (O_2229,N_24653,N_24934);
or UO_2230 (O_2230,N_24728,N_24679);
nand UO_2231 (O_2231,N_24867,N_24791);
nand UO_2232 (O_2232,N_24549,N_24871);
or UO_2233 (O_2233,N_24878,N_24953);
nand UO_2234 (O_2234,N_24514,N_24685);
nand UO_2235 (O_2235,N_24869,N_24891);
xnor UO_2236 (O_2236,N_24837,N_24558);
nor UO_2237 (O_2237,N_24553,N_24961);
and UO_2238 (O_2238,N_24626,N_24706);
and UO_2239 (O_2239,N_24993,N_24641);
or UO_2240 (O_2240,N_24778,N_24697);
xor UO_2241 (O_2241,N_24833,N_24702);
nor UO_2242 (O_2242,N_24561,N_24931);
nand UO_2243 (O_2243,N_24759,N_24860);
nand UO_2244 (O_2244,N_24847,N_24753);
xnor UO_2245 (O_2245,N_24864,N_24747);
nand UO_2246 (O_2246,N_24914,N_24705);
or UO_2247 (O_2247,N_24965,N_24629);
and UO_2248 (O_2248,N_24559,N_24834);
nor UO_2249 (O_2249,N_24963,N_24557);
xor UO_2250 (O_2250,N_24587,N_24974);
and UO_2251 (O_2251,N_24932,N_24590);
xor UO_2252 (O_2252,N_24606,N_24713);
or UO_2253 (O_2253,N_24855,N_24984);
nand UO_2254 (O_2254,N_24692,N_24923);
xor UO_2255 (O_2255,N_24609,N_24641);
nor UO_2256 (O_2256,N_24563,N_24838);
xnor UO_2257 (O_2257,N_24923,N_24548);
or UO_2258 (O_2258,N_24529,N_24850);
and UO_2259 (O_2259,N_24691,N_24686);
and UO_2260 (O_2260,N_24944,N_24898);
and UO_2261 (O_2261,N_24550,N_24501);
nand UO_2262 (O_2262,N_24633,N_24779);
or UO_2263 (O_2263,N_24650,N_24873);
or UO_2264 (O_2264,N_24805,N_24689);
nand UO_2265 (O_2265,N_24933,N_24996);
nor UO_2266 (O_2266,N_24752,N_24750);
nand UO_2267 (O_2267,N_24573,N_24820);
nor UO_2268 (O_2268,N_24941,N_24949);
or UO_2269 (O_2269,N_24515,N_24701);
or UO_2270 (O_2270,N_24880,N_24953);
and UO_2271 (O_2271,N_24508,N_24717);
nor UO_2272 (O_2272,N_24729,N_24574);
and UO_2273 (O_2273,N_24607,N_24885);
nand UO_2274 (O_2274,N_24655,N_24977);
nand UO_2275 (O_2275,N_24766,N_24971);
nor UO_2276 (O_2276,N_24877,N_24802);
and UO_2277 (O_2277,N_24996,N_24559);
or UO_2278 (O_2278,N_24902,N_24650);
xor UO_2279 (O_2279,N_24568,N_24737);
and UO_2280 (O_2280,N_24808,N_24875);
xor UO_2281 (O_2281,N_24594,N_24912);
and UO_2282 (O_2282,N_24878,N_24815);
nand UO_2283 (O_2283,N_24639,N_24592);
nand UO_2284 (O_2284,N_24844,N_24636);
and UO_2285 (O_2285,N_24696,N_24621);
or UO_2286 (O_2286,N_24842,N_24935);
xor UO_2287 (O_2287,N_24979,N_24554);
and UO_2288 (O_2288,N_24541,N_24680);
xnor UO_2289 (O_2289,N_24842,N_24596);
nand UO_2290 (O_2290,N_24516,N_24974);
xor UO_2291 (O_2291,N_24587,N_24755);
and UO_2292 (O_2292,N_24592,N_24689);
nor UO_2293 (O_2293,N_24584,N_24625);
xor UO_2294 (O_2294,N_24619,N_24807);
or UO_2295 (O_2295,N_24622,N_24789);
and UO_2296 (O_2296,N_24839,N_24675);
and UO_2297 (O_2297,N_24996,N_24758);
and UO_2298 (O_2298,N_24612,N_24809);
or UO_2299 (O_2299,N_24854,N_24987);
and UO_2300 (O_2300,N_24531,N_24850);
xor UO_2301 (O_2301,N_24998,N_24842);
or UO_2302 (O_2302,N_24975,N_24984);
and UO_2303 (O_2303,N_24624,N_24604);
nand UO_2304 (O_2304,N_24797,N_24701);
nor UO_2305 (O_2305,N_24814,N_24694);
xor UO_2306 (O_2306,N_24810,N_24579);
nand UO_2307 (O_2307,N_24924,N_24721);
and UO_2308 (O_2308,N_24630,N_24660);
nand UO_2309 (O_2309,N_24542,N_24687);
or UO_2310 (O_2310,N_24661,N_24510);
or UO_2311 (O_2311,N_24842,N_24647);
nand UO_2312 (O_2312,N_24839,N_24764);
nor UO_2313 (O_2313,N_24952,N_24566);
nor UO_2314 (O_2314,N_24693,N_24923);
nor UO_2315 (O_2315,N_24718,N_24930);
nor UO_2316 (O_2316,N_24911,N_24950);
and UO_2317 (O_2317,N_24865,N_24907);
or UO_2318 (O_2318,N_24673,N_24868);
xor UO_2319 (O_2319,N_24561,N_24892);
nand UO_2320 (O_2320,N_24535,N_24970);
nor UO_2321 (O_2321,N_24991,N_24711);
or UO_2322 (O_2322,N_24626,N_24659);
and UO_2323 (O_2323,N_24662,N_24633);
and UO_2324 (O_2324,N_24824,N_24750);
or UO_2325 (O_2325,N_24520,N_24975);
nor UO_2326 (O_2326,N_24808,N_24860);
and UO_2327 (O_2327,N_24937,N_24552);
nor UO_2328 (O_2328,N_24621,N_24912);
or UO_2329 (O_2329,N_24830,N_24571);
nor UO_2330 (O_2330,N_24821,N_24943);
and UO_2331 (O_2331,N_24541,N_24536);
nor UO_2332 (O_2332,N_24867,N_24694);
or UO_2333 (O_2333,N_24830,N_24856);
nor UO_2334 (O_2334,N_24755,N_24859);
or UO_2335 (O_2335,N_24531,N_24563);
or UO_2336 (O_2336,N_24848,N_24717);
nor UO_2337 (O_2337,N_24766,N_24535);
xor UO_2338 (O_2338,N_24814,N_24798);
or UO_2339 (O_2339,N_24994,N_24821);
and UO_2340 (O_2340,N_24843,N_24935);
nor UO_2341 (O_2341,N_24749,N_24962);
or UO_2342 (O_2342,N_24583,N_24614);
nand UO_2343 (O_2343,N_24884,N_24674);
nand UO_2344 (O_2344,N_24555,N_24955);
xor UO_2345 (O_2345,N_24515,N_24678);
nand UO_2346 (O_2346,N_24708,N_24545);
or UO_2347 (O_2347,N_24584,N_24550);
or UO_2348 (O_2348,N_24692,N_24938);
nand UO_2349 (O_2349,N_24894,N_24690);
nor UO_2350 (O_2350,N_24943,N_24851);
nor UO_2351 (O_2351,N_24695,N_24645);
or UO_2352 (O_2352,N_24660,N_24558);
nand UO_2353 (O_2353,N_24970,N_24665);
xor UO_2354 (O_2354,N_24955,N_24970);
or UO_2355 (O_2355,N_24913,N_24661);
or UO_2356 (O_2356,N_24626,N_24547);
or UO_2357 (O_2357,N_24619,N_24559);
nor UO_2358 (O_2358,N_24773,N_24711);
nor UO_2359 (O_2359,N_24673,N_24824);
xor UO_2360 (O_2360,N_24750,N_24590);
nand UO_2361 (O_2361,N_24816,N_24640);
xor UO_2362 (O_2362,N_24702,N_24628);
and UO_2363 (O_2363,N_24771,N_24741);
nor UO_2364 (O_2364,N_24684,N_24961);
xor UO_2365 (O_2365,N_24851,N_24619);
and UO_2366 (O_2366,N_24720,N_24611);
nor UO_2367 (O_2367,N_24714,N_24809);
nor UO_2368 (O_2368,N_24921,N_24779);
and UO_2369 (O_2369,N_24571,N_24727);
or UO_2370 (O_2370,N_24538,N_24501);
nor UO_2371 (O_2371,N_24785,N_24596);
xnor UO_2372 (O_2372,N_24870,N_24891);
xor UO_2373 (O_2373,N_24983,N_24683);
xor UO_2374 (O_2374,N_24587,N_24730);
or UO_2375 (O_2375,N_24932,N_24797);
or UO_2376 (O_2376,N_24673,N_24618);
xor UO_2377 (O_2377,N_24617,N_24995);
nand UO_2378 (O_2378,N_24870,N_24761);
or UO_2379 (O_2379,N_24781,N_24860);
and UO_2380 (O_2380,N_24881,N_24765);
xnor UO_2381 (O_2381,N_24878,N_24745);
nand UO_2382 (O_2382,N_24671,N_24716);
nand UO_2383 (O_2383,N_24617,N_24865);
nor UO_2384 (O_2384,N_24836,N_24540);
xnor UO_2385 (O_2385,N_24889,N_24720);
nand UO_2386 (O_2386,N_24731,N_24717);
nor UO_2387 (O_2387,N_24891,N_24944);
xnor UO_2388 (O_2388,N_24547,N_24590);
and UO_2389 (O_2389,N_24606,N_24793);
nand UO_2390 (O_2390,N_24886,N_24833);
and UO_2391 (O_2391,N_24701,N_24772);
or UO_2392 (O_2392,N_24555,N_24908);
nor UO_2393 (O_2393,N_24548,N_24508);
and UO_2394 (O_2394,N_24768,N_24772);
nor UO_2395 (O_2395,N_24519,N_24610);
or UO_2396 (O_2396,N_24921,N_24897);
and UO_2397 (O_2397,N_24594,N_24537);
xor UO_2398 (O_2398,N_24990,N_24698);
or UO_2399 (O_2399,N_24774,N_24643);
nand UO_2400 (O_2400,N_24573,N_24633);
xnor UO_2401 (O_2401,N_24696,N_24503);
xnor UO_2402 (O_2402,N_24586,N_24603);
or UO_2403 (O_2403,N_24594,N_24994);
xor UO_2404 (O_2404,N_24801,N_24750);
or UO_2405 (O_2405,N_24863,N_24534);
xnor UO_2406 (O_2406,N_24927,N_24972);
or UO_2407 (O_2407,N_24941,N_24776);
and UO_2408 (O_2408,N_24627,N_24519);
xor UO_2409 (O_2409,N_24745,N_24877);
xnor UO_2410 (O_2410,N_24850,N_24602);
and UO_2411 (O_2411,N_24692,N_24830);
and UO_2412 (O_2412,N_24520,N_24671);
nor UO_2413 (O_2413,N_24910,N_24777);
or UO_2414 (O_2414,N_24974,N_24568);
nor UO_2415 (O_2415,N_24797,N_24694);
and UO_2416 (O_2416,N_24885,N_24980);
nand UO_2417 (O_2417,N_24900,N_24896);
or UO_2418 (O_2418,N_24781,N_24937);
xor UO_2419 (O_2419,N_24671,N_24776);
nand UO_2420 (O_2420,N_24744,N_24535);
nor UO_2421 (O_2421,N_24945,N_24877);
or UO_2422 (O_2422,N_24988,N_24773);
nor UO_2423 (O_2423,N_24931,N_24767);
nor UO_2424 (O_2424,N_24589,N_24653);
nor UO_2425 (O_2425,N_24932,N_24618);
xor UO_2426 (O_2426,N_24838,N_24919);
xnor UO_2427 (O_2427,N_24958,N_24757);
or UO_2428 (O_2428,N_24727,N_24770);
nor UO_2429 (O_2429,N_24595,N_24581);
or UO_2430 (O_2430,N_24860,N_24617);
xor UO_2431 (O_2431,N_24596,N_24964);
or UO_2432 (O_2432,N_24973,N_24611);
nor UO_2433 (O_2433,N_24877,N_24916);
or UO_2434 (O_2434,N_24644,N_24786);
nand UO_2435 (O_2435,N_24727,N_24851);
and UO_2436 (O_2436,N_24650,N_24868);
xor UO_2437 (O_2437,N_24649,N_24536);
xor UO_2438 (O_2438,N_24949,N_24502);
and UO_2439 (O_2439,N_24762,N_24957);
nor UO_2440 (O_2440,N_24635,N_24722);
or UO_2441 (O_2441,N_24702,N_24839);
nand UO_2442 (O_2442,N_24763,N_24823);
nand UO_2443 (O_2443,N_24884,N_24993);
nand UO_2444 (O_2444,N_24623,N_24674);
or UO_2445 (O_2445,N_24995,N_24855);
xnor UO_2446 (O_2446,N_24698,N_24659);
xnor UO_2447 (O_2447,N_24856,N_24868);
or UO_2448 (O_2448,N_24782,N_24946);
nand UO_2449 (O_2449,N_24865,N_24720);
or UO_2450 (O_2450,N_24731,N_24675);
and UO_2451 (O_2451,N_24989,N_24887);
nand UO_2452 (O_2452,N_24797,N_24760);
nor UO_2453 (O_2453,N_24849,N_24914);
xor UO_2454 (O_2454,N_24558,N_24893);
or UO_2455 (O_2455,N_24701,N_24608);
nand UO_2456 (O_2456,N_24632,N_24943);
and UO_2457 (O_2457,N_24831,N_24535);
nand UO_2458 (O_2458,N_24783,N_24771);
nand UO_2459 (O_2459,N_24561,N_24758);
nor UO_2460 (O_2460,N_24543,N_24789);
nand UO_2461 (O_2461,N_24829,N_24790);
nand UO_2462 (O_2462,N_24846,N_24504);
or UO_2463 (O_2463,N_24615,N_24909);
or UO_2464 (O_2464,N_24707,N_24622);
and UO_2465 (O_2465,N_24989,N_24600);
nor UO_2466 (O_2466,N_24762,N_24847);
xnor UO_2467 (O_2467,N_24929,N_24966);
or UO_2468 (O_2468,N_24694,N_24535);
and UO_2469 (O_2469,N_24875,N_24949);
and UO_2470 (O_2470,N_24698,N_24746);
and UO_2471 (O_2471,N_24597,N_24670);
nand UO_2472 (O_2472,N_24899,N_24602);
or UO_2473 (O_2473,N_24764,N_24847);
and UO_2474 (O_2474,N_24837,N_24757);
and UO_2475 (O_2475,N_24975,N_24699);
nor UO_2476 (O_2476,N_24897,N_24701);
and UO_2477 (O_2477,N_24798,N_24790);
or UO_2478 (O_2478,N_24575,N_24588);
nand UO_2479 (O_2479,N_24791,N_24874);
or UO_2480 (O_2480,N_24676,N_24757);
nor UO_2481 (O_2481,N_24517,N_24794);
nor UO_2482 (O_2482,N_24766,N_24839);
nand UO_2483 (O_2483,N_24766,N_24954);
or UO_2484 (O_2484,N_24718,N_24811);
xor UO_2485 (O_2485,N_24627,N_24787);
or UO_2486 (O_2486,N_24773,N_24738);
nor UO_2487 (O_2487,N_24867,N_24553);
nand UO_2488 (O_2488,N_24584,N_24911);
and UO_2489 (O_2489,N_24538,N_24948);
nand UO_2490 (O_2490,N_24905,N_24590);
xor UO_2491 (O_2491,N_24884,N_24879);
nand UO_2492 (O_2492,N_24971,N_24925);
xor UO_2493 (O_2493,N_24997,N_24752);
nand UO_2494 (O_2494,N_24872,N_24605);
xor UO_2495 (O_2495,N_24770,N_24852);
xor UO_2496 (O_2496,N_24981,N_24770);
xor UO_2497 (O_2497,N_24856,N_24807);
nand UO_2498 (O_2498,N_24594,N_24766);
nor UO_2499 (O_2499,N_24559,N_24512);
nand UO_2500 (O_2500,N_24534,N_24834);
xnor UO_2501 (O_2501,N_24995,N_24927);
nor UO_2502 (O_2502,N_24690,N_24544);
and UO_2503 (O_2503,N_24621,N_24974);
and UO_2504 (O_2504,N_24670,N_24813);
or UO_2505 (O_2505,N_24847,N_24918);
and UO_2506 (O_2506,N_24884,N_24524);
nor UO_2507 (O_2507,N_24609,N_24834);
nor UO_2508 (O_2508,N_24819,N_24918);
nor UO_2509 (O_2509,N_24741,N_24537);
nand UO_2510 (O_2510,N_24689,N_24924);
nor UO_2511 (O_2511,N_24645,N_24848);
or UO_2512 (O_2512,N_24888,N_24757);
nand UO_2513 (O_2513,N_24661,N_24897);
xor UO_2514 (O_2514,N_24666,N_24894);
nor UO_2515 (O_2515,N_24843,N_24782);
xnor UO_2516 (O_2516,N_24823,N_24774);
or UO_2517 (O_2517,N_24578,N_24775);
nand UO_2518 (O_2518,N_24756,N_24759);
nand UO_2519 (O_2519,N_24737,N_24713);
or UO_2520 (O_2520,N_24643,N_24727);
or UO_2521 (O_2521,N_24599,N_24512);
or UO_2522 (O_2522,N_24672,N_24519);
nand UO_2523 (O_2523,N_24927,N_24956);
or UO_2524 (O_2524,N_24741,N_24731);
and UO_2525 (O_2525,N_24918,N_24853);
or UO_2526 (O_2526,N_24747,N_24885);
nand UO_2527 (O_2527,N_24931,N_24974);
and UO_2528 (O_2528,N_24823,N_24752);
xnor UO_2529 (O_2529,N_24789,N_24533);
nand UO_2530 (O_2530,N_24622,N_24744);
nor UO_2531 (O_2531,N_24857,N_24658);
nand UO_2532 (O_2532,N_24959,N_24500);
or UO_2533 (O_2533,N_24778,N_24584);
and UO_2534 (O_2534,N_24594,N_24898);
nand UO_2535 (O_2535,N_24594,N_24775);
nand UO_2536 (O_2536,N_24522,N_24538);
xnor UO_2537 (O_2537,N_24579,N_24688);
nand UO_2538 (O_2538,N_24599,N_24818);
or UO_2539 (O_2539,N_24581,N_24588);
nor UO_2540 (O_2540,N_24687,N_24981);
nor UO_2541 (O_2541,N_24953,N_24837);
xor UO_2542 (O_2542,N_24533,N_24764);
nor UO_2543 (O_2543,N_24693,N_24782);
xor UO_2544 (O_2544,N_24659,N_24566);
xnor UO_2545 (O_2545,N_24826,N_24657);
nor UO_2546 (O_2546,N_24688,N_24865);
nor UO_2547 (O_2547,N_24722,N_24771);
or UO_2548 (O_2548,N_24740,N_24854);
nand UO_2549 (O_2549,N_24534,N_24975);
nor UO_2550 (O_2550,N_24705,N_24829);
or UO_2551 (O_2551,N_24641,N_24735);
and UO_2552 (O_2552,N_24590,N_24654);
nand UO_2553 (O_2553,N_24520,N_24704);
nor UO_2554 (O_2554,N_24997,N_24537);
nand UO_2555 (O_2555,N_24792,N_24866);
or UO_2556 (O_2556,N_24669,N_24865);
and UO_2557 (O_2557,N_24967,N_24597);
xnor UO_2558 (O_2558,N_24525,N_24714);
nor UO_2559 (O_2559,N_24649,N_24975);
xnor UO_2560 (O_2560,N_24639,N_24760);
nand UO_2561 (O_2561,N_24936,N_24665);
and UO_2562 (O_2562,N_24880,N_24558);
nand UO_2563 (O_2563,N_24654,N_24932);
or UO_2564 (O_2564,N_24730,N_24953);
and UO_2565 (O_2565,N_24965,N_24739);
nor UO_2566 (O_2566,N_24541,N_24590);
nand UO_2567 (O_2567,N_24973,N_24705);
or UO_2568 (O_2568,N_24572,N_24519);
and UO_2569 (O_2569,N_24695,N_24956);
nor UO_2570 (O_2570,N_24830,N_24501);
xor UO_2571 (O_2571,N_24652,N_24779);
or UO_2572 (O_2572,N_24773,N_24845);
or UO_2573 (O_2573,N_24746,N_24705);
xor UO_2574 (O_2574,N_24697,N_24656);
or UO_2575 (O_2575,N_24936,N_24785);
xor UO_2576 (O_2576,N_24955,N_24798);
and UO_2577 (O_2577,N_24672,N_24958);
and UO_2578 (O_2578,N_24794,N_24515);
nand UO_2579 (O_2579,N_24701,N_24532);
or UO_2580 (O_2580,N_24608,N_24510);
and UO_2581 (O_2581,N_24596,N_24604);
nor UO_2582 (O_2582,N_24642,N_24645);
and UO_2583 (O_2583,N_24976,N_24785);
nor UO_2584 (O_2584,N_24989,N_24637);
nand UO_2585 (O_2585,N_24977,N_24632);
nor UO_2586 (O_2586,N_24702,N_24599);
and UO_2587 (O_2587,N_24524,N_24501);
or UO_2588 (O_2588,N_24837,N_24658);
nor UO_2589 (O_2589,N_24789,N_24964);
or UO_2590 (O_2590,N_24923,N_24871);
and UO_2591 (O_2591,N_24566,N_24543);
or UO_2592 (O_2592,N_24526,N_24837);
xnor UO_2593 (O_2593,N_24512,N_24824);
xor UO_2594 (O_2594,N_24645,N_24680);
and UO_2595 (O_2595,N_24781,N_24832);
nand UO_2596 (O_2596,N_24821,N_24876);
or UO_2597 (O_2597,N_24540,N_24915);
and UO_2598 (O_2598,N_24898,N_24597);
and UO_2599 (O_2599,N_24595,N_24960);
or UO_2600 (O_2600,N_24689,N_24731);
and UO_2601 (O_2601,N_24809,N_24920);
nor UO_2602 (O_2602,N_24901,N_24734);
and UO_2603 (O_2603,N_24556,N_24928);
or UO_2604 (O_2604,N_24834,N_24901);
nand UO_2605 (O_2605,N_24561,N_24529);
xor UO_2606 (O_2606,N_24899,N_24559);
nor UO_2607 (O_2607,N_24594,N_24719);
xnor UO_2608 (O_2608,N_24523,N_24728);
and UO_2609 (O_2609,N_24610,N_24705);
nand UO_2610 (O_2610,N_24848,N_24934);
nor UO_2611 (O_2611,N_24718,N_24537);
xnor UO_2612 (O_2612,N_24995,N_24937);
or UO_2613 (O_2613,N_24898,N_24635);
and UO_2614 (O_2614,N_24975,N_24608);
nand UO_2615 (O_2615,N_24751,N_24725);
or UO_2616 (O_2616,N_24669,N_24580);
nand UO_2617 (O_2617,N_24807,N_24520);
xnor UO_2618 (O_2618,N_24533,N_24581);
and UO_2619 (O_2619,N_24818,N_24808);
nand UO_2620 (O_2620,N_24984,N_24826);
nor UO_2621 (O_2621,N_24668,N_24649);
or UO_2622 (O_2622,N_24665,N_24937);
nor UO_2623 (O_2623,N_24879,N_24912);
xnor UO_2624 (O_2624,N_24802,N_24993);
nor UO_2625 (O_2625,N_24883,N_24904);
xnor UO_2626 (O_2626,N_24547,N_24841);
xnor UO_2627 (O_2627,N_24824,N_24524);
nand UO_2628 (O_2628,N_24852,N_24693);
nor UO_2629 (O_2629,N_24644,N_24906);
nand UO_2630 (O_2630,N_24576,N_24727);
or UO_2631 (O_2631,N_24627,N_24704);
nor UO_2632 (O_2632,N_24830,N_24569);
xor UO_2633 (O_2633,N_24636,N_24612);
nor UO_2634 (O_2634,N_24814,N_24566);
xnor UO_2635 (O_2635,N_24743,N_24832);
and UO_2636 (O_2636,N_24869,N_24829);
nor UO_2637 (O_2637,N_24970,N_24739);
xor UO_2638 (O_2638,N_24520,N_24555);
xnor UO_2639 (O_2639,N_24654,N_24744);
and UO_2640 (O_2640,N_24890,N_24847);
and UO_2641 (O_2641,N_24731,N_24641);
xnor UO_2642 (O_2642,N_24511,N_24730);
nor UO_2643 (O_2643,N_24625,N_24706);
or UO_2644 (O_2644,N_24822,N_24687);
nor UO_2645 (O_2645,N_24814,N_24972);
or UO_2646 (O_2646,N_24825,N_24530);
nor UO_2647 (O_2647,N_24640,N_24653);
nor UO_2648 (O_2648,N_24997,N_24946);
xor UO_2649 (O_2649,N_24622,N_24976);
xnor UO_2650 (O_2650,N_24601,N_24638);
nand UO_2651 (O_2651,N_24581,N_24936);
nor UO_2652 (O_2652,N_24999,N_24913);
and UO_2653 (O_2653,N_24887,N_24800);
nand UO_2654 (O_2654,N_24671,N_24661);
or UO_2655 (O_2655,N_24829,N_24796);
or UO_2656 (O_2656,N_24659,N_24710);
or UO_2657 (O_2657,N_24791,N_24941);
nor UO_2658 (O_2658,N_24908,N_24935);
nor UO_2659 (O_2659,N_24665,N_24570);
xor UO_2660 (O_2660,N_24709,N_24734);
xnor UO_2661 (O_2661,N_24633,N_24912);
xor UO_2662 (O_2662,N_24764,N_24651);
and UO_2663 (O_2663,N_24728,N_24538);
xor UO_2664 (O_2664,N_24588,N_24718);
nand UO_2665 (O_2665,N_24678,N_24742);
or UO_2666 (O_2666,N_24969,N_24546);
nand UO_2667 (O_2667,N_24911,N_24888);
xnor UO_2668 (O_2668,N_24537,N_24569);
and UO_2669 (O_2669,N_24544,N_24677);
nand UO_2670 (O_2670,N_24502,N_24679);
nand UO_2671 (O_2671,N_24911,N_24653);
nor UO_2672 (O_2672,N_24785,N_24768);
nand UO_2673 (O_2673,N_24802,N_24622);
nor UO_2674 (O_2674,N_24812,N_24944);
xor UO_2675 (O_2675,N_24791,N_24533);
nand UO_2676 (O_2676,N_24936,N_24691);
xor UO_2677 (O_2677,N_24849,N_24846);
nor UO_2678 (O_2678,N_24520,N_24690);
nor UO_2679 (O_2679,N_24920,N_24695);
nor UO_2680 (O_2680,N_24716,N_24915);
or UO_2681 (O_2681,N_24691,N_24880);
nand UO_2682 (O_2682,N_24988,N_24862);
and UO_2683 (O_2683,N_24873,N_24692);
nor UO_2684 (O_2684,N_24944,N_24743);
or UO_2685 (O_2685,N_24681,N_24804);
nor UO_2686 (O_2686,N_24988,N_24548);
nand UO_2687 (O_2687,N_24932,N_24688);
xnor UO_2688 (O_2688,N_24757,N_24623);
or UO_2689 (O_2689,N_24791,N_24988);
nor UO_2690 (O_2690,N_24589,N_24735);
or UO_2691 (O_2691,N_24729,N_24863);
nand UO_2692 (O_2692,N_24827,N_24525);
or UO_2693 (O_2693,N_24769,N_24836);
nor UO_2694 (O_2694,N_24905,N_24843);
nor UO_2695 (O_2695,N_24664,N_24933);
and UO_2696 (O_2696,N_24610,N_24677);
and UO_2697 (O_2697,N_24811,N_24626);
and UO_2698 (O_2698,N_24835,N_24958);
xnor UO_2699 (O_2699,N_24770,N_24507);
xor UO_2700 (O_2700,N_24675,N_24628);
and UO_2701 (O_2701,N_24567,N_24667);
and UO_2702 (O_2702,N_24527,N_24791);
nand UO_2703 (O_2703,N_24805,N_24643);
nand UO_2704 (O_2704,N_24859,N_24543);
or UO_2705 (O_2705,N_24527,N_24860);
nor UO_2706 (O_2706,N_24917,N_24784);
and UO_2707 (O_2707,N_24889,N_24732);
nor UO_2708 (O_2708,N_24811,N_24954);
xnor UO_2709 (O_2709,N_24876,N_24516);
or UO_2710 (O_2710,N_24758,N_24863);
or UO_2711 (O_2711,N_24520,N_24587);
nand UO_2712 (O_2712,N_24737,N_24884);
xor UO_2713 (O_2713,N_24760,N_24783);
and UO_2714 (O_2714,N_24990,N_24853);
or UO_2715 (O_2715,N_24591,N_24993);
or UO_2716 (O_2716,N_24547,N_24578);
or UO_2717 (O_2717,N_24899,N_24787);
nor UO_2718 (O_2718,N_24587,N_24964);
xnor UO_2719 (O_2719,N_24789,N_24863);
xor UO_2720 (O_2720,N_24605,N_24880);
nor UO_2721 (O_2721,N_24590,N_24966);
nor UO_2722 (O_2722,N_24984,N_24886);
nand UO_2723 (O_2723,N_24814,N_24678);
and UO_2724 (O_2724,N_24603,N_24856);
nand UO_2725 (O_2725,N_24764,N_24890);
xnor UO_2726 (O_2726,N_24792,N_24795);
nor UO_2727 (O_2727,N_24762,N_24831);
and UO_2728 (O_2728,N_24797,N_24508);
nand UO_2729 (O_2729,N_24710,N_24588);
nand UO_2730 (O_2730,N_24523,N_24975);
or UO_2731 (O_2731,N_24787,N_24898);
nand UO_2732 (O_2732,N_24965,N_24548);
and UO_2733 (O_2733,N_24938,N_24759);
and UO_2734 (O_2734,N_24701,N_24666);
and UO_2735 (O_2735,N_24673,N_24644);
nand UO_2736 (O_2736,N_24608,N_24994);
xnor UO_2737 (O_2737,N_24733,N_24690);
nor UO_2738 (O_2738,N_24682,N_24629);
or UO_2739 (O_2739,N_24629,N_24603);
nor UO_2740 (O_2740,N_24613,N_24902);
nor UO_2741 (O_2741,N_24705,N_24595);
nand UO_2742 (O_2742,N_24873,N_24523);
xor UO_2743 (O_2743,N_24760,N_24708);
nand UO_2744 (O_2744,N_24605,N_24919);
and UO_2745 (O_2745,N_24776,N_24759);
xnor UO_2746 (O_2746,N_24699,N_24679);
nor UO_2747 (O_2747,N_24738,N_24921);
nand UO_2748 (O_2748,N_24658,N_24813);
xnor UO_2749 (O_2749,N_24639,N_24584);
xor UO_2750 (O_2750,N_24746,N_24693);
or UO_2751 (O_2751,N_24847,N_24672);
or UO_2752 (O_2752,N_24789,N_24970);
xnor UO_2753 (O_2753,N_24622,N_24550);
nand UO_2754 (O_2754,N_24599,N_24840);
or UO_2755 (O_2755,N_24549,N_24615);
or UO_2756 (O_2756,N_24535,N_24547);
or UO_2757 (O_2757,N_24683,N_24895);
nor UO_2758 (O_2758,N_24789,N_24523);
nand UO_2759 (O_2759,N_24629,N_24930);
and UO_2760 (O_2760,N_24628,N_24780);
nor UO_2761 (O_2761,N_24730,N_24550);
and UO_2762 (O_2762,N_24934,N_24876);
nand UO_2763 (O_2763,N_24567,N_24967);
and UO_2764 (O_2764,N_24952,N_24582);
nand UO_2765 (O_2765,N_24591,N_24889);
nand UO_2766 (O_2766,N_24507,N_24774);
nand UO_2767 (O_2767,N_24769,N_24957);
or UO_2768 (O_2768,N_24899,N_24694);
xor UO_2769 (O_2769,N_24730,N_24829);
and UO_2770 (O_2770,N_24950,N_24550);
nor UO_2771 (O_2771,N_24962,N_24856);
nor UO_2772 (O_2772,N_24754,N_24905);
nor UO_2773 (O_2773,N_24585,N_24750);
and UO_2774 (O_2774,N_24688,N_24644);
or UO_2775 (O_2775,N_24653,N_24630);
or UO_2776 (O_2776,N_24805,N_24750);
or UO_2777 (O_2777,N_24623,N_24743);
and UO_2778 (O_2778,N_24547,N_24583);
nand UO_2779 (O_2779,N_24843,N_24856);
xor UO_2780 (O_2780,N_24859,N_24898);
or UO_2781 (O_2781,N_24618,N_24764);
nand UO_2782 (O_2782,N_24697,N_24562);
or UO_2783 (O_2783,N_24685,N_24887);
nor UO_2784 (O_2784,N_24619,N_24970);
xnor UO_2785 (O_2785,N_24700,N_24764);
nor UO_2786 (O_2786,N_24679,N_24923);
and UO_2787 (O_2787,N_24699,N_24861);
or UO_2788 (O_2788,N_24905,N_24541);
and UO_2789 (O_2789,N_24666,N_24954);
or UO_2790 (O_2790,N_24819,N_24846);
and UO_2791 (O_2791,N_24841,N_24742);
and UO_2792 (O_2792,N_24890,N_24513);
nand UO_2793 (O_2793,N_24756,N_24683);
and UO_2794 (O_2794,N_24643,N_24538);
and UO_2795 (O_2795,N_24830,N_24661);
nor UO_2796 (O_2796,N_24977,N_24778);
nor UO_2797 (O_2797,N_24682,N_24925);
xor UO_2798 (O_2798,N_24725,N_24917);
xor UO_2799 (O_2799,N_24655,N_24649);
or UO_2800 (O_2800,N_24710,N_24766);
or UO_2801 (O_2801,N_24736,N_24871);
nand UO_2802 (O_2802,N_24877,N_24875);
xor UO_2803 (O_2803,N_24614,N_24551);
nand UO_2804 (O_2804,N_24858,N_24522);
xnor UO_2805 (O_2805,N_24781,N_24866);
xor UO_2806 (O_2806,N_24919,N_24722);
or UO_2807 (O_2807,N_24600,N_24732);
and UO_2808 (O_2808,N_24663,N_24637);
and UO_2809 (O_2809,N_24630,N_24904);
nand UO_2810 (O_2810,N_24573,N_24715);
nand UO_2811 (O_2811,N_24936,N_24938);
and UO_2812 (O_2812,N_24958,N_24827);
nor UO_2813 (O_2813,N_24797,N_24558);
nand UO_2814 (O_2814,N_24811,N_24856);
xnor UO_2815 (O_2815,N_24795,N_24579);
nand UO_2816 (O_2816,N_24752,N_24609);
xor UO_2817 (O_2817,N_24624,N_24598);
xnor UO_2818 (O_2818,N_24767,N_24862);
or UO_2819 (O_2819,N_24752,N_24873);
and UO_2820 (O_2820,N_24810,N_24879);
nor UO_2821 (O_2821,N_24605,N_24599);
and UO_2822 (O_2822,N_24764,N_24568);
nand UO_2823 (O_2823,N_24796,N_24866);
nor UO_2824 (O_2824,N_24995,N_24728);
nand UO_2825 (O_2825,N_24523,N_24696);
nand UO_2826 (O_2826,N_24505,N_24977);
nor UO_2827 (O_2827,N_24858,N_24976);
or UO_2828 (O_2828,N_24816,N_24960);
and UO_2829 (O_2829,N_24706,N_24785);
and UO_2830 (O_2830,N_24678,N_24813);
or UO_2831 (O_2831,N_24596,N_24676);
nand UO_2832 (O_2832,N_24892,N_24584);
or UO_2833 (O_2833,N_24876,N_24534);
nand UO_2834 (O_2834,N_24509,N_24569);
xor UO_2835 (O_2835,N_24835,N_24694);
nand UO_2836 (O_2836,N_24550,N_24618);
nand UO_2837 (O_2837,N_24686,N_24681);
and UO_2838 (O_2838,N_24979,N_24911);
xnor UO_2839 (O_2839,N_24804,N_24911);
nor UO_2840 (O_2840,N_24818,N_24979);
and UO_2841 (O_2841,N_24962,N_24725);
and UO_2842 (O_2842,N_24860,N_24939);
nor UO_2843 (O_2843,N_24904,N_24841);
nand UO_2844 (O_2844,N_24628,N_24694);
nand UO_2845 (O_2845,N_24503,N_24811);
or UO_2846 (O_2846,N_24758,N_24822);
nand UO_2847 (O_2847,N_24728,N_24913);
and UO_2848 (O_2848,N_24591,N_24634);
nor UO_2849 (O_2849,N_24682,N_24781);
xor UO_2850 (O_2850,N_24817,N_24727);
xnor UO_2851 (O_2851,N_24842,N_24984);
nand UO_2852 (O_2852,N_24757,N_24899);
or UO_2853 (O_2853,N_24782,N_24780);
nor UO_2854 (O_2854,N_24717,N_24837);
or UO_2855 (O_2855,N_24672,N_24979);
and UO_2856 (O_2856,N_24853,N_24750);
and UO_2857 (O_2857,N_24601,N_24564);
xor UO_2858 (O_2858,N_24970,N_24945);
nor UO_2859 (O_2859,N_24702,N_24888);
and UO_2860 (O_2860,N_24547,N_24560);
nor UO_2861 (O_2861,N_24708,N_24578);
nand UO_2862 (O_2862,N_24888,N_24803);
xor UO_2863 (O_2863,N_24995,N_24843);
or UO_2864 (O_2864,N_24612,N_24856);
and UO_2865 (O_2865,N_24540,N_24998);
nand UO_2866 (O_2866,N_24557,N_24998);
or UO_2867 (O_2867,N_24935,N_24778);
or UO_2868 (O_2868,N_24992,N_24824);
and UO_2869 (O_2869,N_24862,N_24544);
nor UO_2870 (O_2870,N_24909,N_24758);
nand UO_2871 (O_2871,N_24997,N_24822);
and UO_2872 (O_2872,N_24895,N_24954);
or UO_2873 (O_2873,N_24759,N_24929);
nand UO_2874 (O_2874,N_24780,N_24732);
and UO_2875 (O_2875,N_24791,N_24794);
and UO_2876 (O_2876,N_24989,N_24816);
nand UO_2877 (O_2877,N_24705,N_24890);
and UO_2878 (O_2878,N_24949,N_24629);
or UO_2879 (O_2879,N_24634,N_24640);
nor UO_2880 (O_2880,N_24930,N_24533);
xnor UO_2881 (O_2881,N_24850,N_24816);
nor UO_2882 (O_2882,N_24509,N_24834);
or UO_2883 (O_2883,N_24788,N_24718);
and UO_2884 (O_2884,N_24933,N_24946);
nand UO_2885 (O_2885,N_24562,N_24575);
nor UO_2886 (O_2886,N_24919,N_24765);
nand UO_2887 (O_2887,N_24826,N_24537);
or UO_2888 (O_2888,N_24698,N_24671);
xnor UO_2889 (O_2889,N_24954,N_24775);
xor UO_2890 (O_2890,N_24734,N_24609);
xnor UO_2891 (O_2891,N_24551,N_24851);
xor UO_2892 (O_2892,N_24749,N_24945);
nor UO_2893 (O_2893,N_24517,N_24867);
nor UO_2894 (O_2894,N_24846,N_24848);
and UO_2895 (O_2895,N_24882,N_24861);
and UO_2896 (O_2896,N_24566,N_24695);
and UO_2897 (O_2897,N_24935,N_24594);
nand UO_2898 (O_2898,N_24519,N_24730);
and UO_2899 (O_2899,N_24628,N_24619);
or UO_2900 (O_2900,N_24977,N_24646);
nand UO_2901 (O_2901,N_24740,N_24951);
nand UO_2902 (O_2902,N_24723,N_24742);
or UO_2903 (O_2903,N_24835,N_24703);
or UO_2904 (O_2904,N_24535,N_24602);
or UO_2905 (O_2905,N_24606,N_24999);
nand UO_2906 (O_2906,N_24507,N_24965);
xnor UO_2907 (O_2907,N_24641,N_24892);
nor UO_2908 (O_2908,N_24649,N_24507);
and UO_2909 (O_2909,N_24980,N_24757);
and UO_2910 (O_2910,N_24864,N_24793);
nor UO_2911 (O_2911,N_24562,N_24708);
or UO_2912 (O_2912,N_24705,N_24644);
and UO_2913 (O_2913,N_24812,N_24592);
xor UO_2914 (O_2914,N_24774,N_24727);
xor UO_2915 (O_2915,N_24942,N_24917);
nand UO_2916 (O_2916,N_24965,N_24811);
or UO_2917 (O_2917,N_24901,N_24521);
xnor UO_2918 (O_2918,N_24758,N_24895);
nor UO_2919 (O_2919,N_24646,N_24659);
xnor UO_2920 (O_2920,N_24871,N_24638);
nor UO_2921 (O_2921,N_24598,N_24570);
xor UO_2922 (O_2922,N_24972,N_24735);
xor UO_2923 (O_2923,N_24666,N_24559);
nand UO_2924 (O_2924,N_24661,N_24907);
nand UO_2925 (O_2925,N_24717,N_24531);
nand UO_2926 (O_2926,N_24728,N_24572);
nand UO_2927 (O_2927,N_24881,N_24780);
xnor UO_2928 (O_2928,N_24717,N_24968);
nor UO_2929 (O_2929,N_24706,N_24868);
and UO_2930 (O_2930,N_24571,N_24550);
and UO_2931 (O_2931,N_24619,N_24737);
nand UO_2932 (O_2932,N_24828,N_24651);
nor UO_2933 (O_2933,N_24928,N_24909);
nand UO_2934 (O_2934,N_24752,N_24683);
nor UO_2935 (O_2935,N_24965,N_24962);
nand UO_2936 (O_2936,N_24999,N_24701);
or UO_2937 (O_2937,N_24580,N_24579);
xor UO_2938 (O_2938,N_24956,N_24697);
nor UO_2939 (O_2939,N_24981,N_24902);
nor UO_2940 (O_2940,N_24897,N_24816);
or UO_2941 (O_2941,N_24636,N_24713);
xor UO_2942 (O_2942,N_24795,N_24917);
nor UO_2943 (O_2943,N_24743,N_24970);
and UO_2944 (O_2944,N_24867,N_24760);
nor UO_2945 (O_2945,N_24925,N_24972);
nand UO_2946 (O_2946,N_24669,N_24700);
xnor UO_2947 (O_2947,N_24501,N_24702);
xor UO_2948 (O_2948,N_24827,N_24808);
nor UO_2949 (O_2949,N_24534,N_24882);
xnor UO_2950 (O_2950,N_24908,N_24801);
nand UO_2951 (O_2951,N_24946,N_24623);
nand UO_2952 (O_2952,N_24995,N_24827);
nand UO_2953 (O_2953,N_24536,N_24653);
nor UO_2954 (O_2954,N_24719,N_24566);
nor UO_2955 (O_2955,N_24808,N_24559);
nor UO_2956 (O_2956,N_24589,N_24969);
or UO_2957 (O_2957,N_24801,N_24758);
or UO_2958 (O_2958,N_24896,N_24638);
nor UO_2959 (O_2959,N_24529,N_24720);
nor UO_2960 (O_2960,N_24876,N_24704);
or UO_2961 (O_2961,N_24887,N_24926);
or UO_2962 (O_2962,N_24905,N_24606);
xnor UO_2963 (O_2963,N_24686,N_24807);
nor UO_2964 (O_2964,N_24964,N_24825);
nor UO_2965 (O_2965,N_24662,N_24621);
or UO_2966 (O_2966,N_24935,N_24598);
nand UO_2967 (O_2967,N_24711,N_24978);
nor UO_2968 (O_2968,N_24827,N_24886);
xnor UO_2969 (O_2969,N_24844,N_24578);
nand UO_2970 (O_2970,N_24794,N_24629);
nor UO_2971 (O_2971,N_24589,N_24683);
nor UO_2972 (O_2972,N_24527,N_24839);
and UO_2973 (O_2973,N_24903,N_24859);
and UO_2974 (O_2974,N_24996,N_24520);
nor UO_2975 (O_2975,N_24793,N_24672);
or UO_2976 (O_2976,N_24843,N_24957);
or UO_2977 (O_2977,N_24905,N_24825);
nor UO_2978 (O_2978,N_24726,N_24718);
xor UO_2979 (O_2979,N_24881,N_24585);
nor UO_2980 (O_2980,N_24762,N_24818);
xor UO_2981 (O_2981,N_24666,N_24638);
nor UO_2982 (O_2982,N_24787,N_24573);
and UO_2983 (O_2983,N_24881,N_24771);
xnor UO_2984 (O_2984,N_24524,N_24753);
or UO_2985 (O_2985,N_24656,N_24609);
nand UO_2986 (O_2986,N_24901,N_24591);
or UO_2987 (O_2987,N_24744,N_24675);
nand UO_2988 (O_2988,N_24868,N_24853);
or UO_2989 (O_2989,N_24784,N_24837);
nor UO_2990 (O_2990,N_24871,N_24970);
and UO_2991 (O_2991,N_24787,N_24919);
or UO_2992 (O_2992,N_24799,N_24985);
nand UO_2993 (O_2993,N_24858,N_24953);
and UO_2994 (O_2994,N_24581,N_24943);
and UO_2995 (O_2995,N_24628,N_24944);
nor UO_2996 (O_2996,N_24682,N_24790);
and UO_2997 (O_2997,N_24615,N_24942);
and UO_2998 (O_2998,N_24855,N_24836);
or UO_2999 (O_2999,N_24608,N_24997);
endmodule