module basic_5000_50000_5000_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_708,In_3762);
or U1 (N_1,In_4271,In_244);
nand U2 (N_2,In_950,In_1963);
nand U3 (N_3,In_4461,In_3358);
nand U4 (N_4,In_3694,In_114);
xor U5 (N_5,In_4442,In_3424);
and U6 (N_6,In_835,In_4733);
nand U7 (N_7,In_3451,In_4812);
and U8 (N_8,In_1249,In_1267);
or U9 (N_9,In_3136,In_2389);
or U10 (N_10,In_2390,In_398);
xor U11 (N_11,In_3124,In_4299);
xor U12 (N_12,In_1129,In_4476);
nor U13 (N_13,In_1471,In_4776);
nor U14 (N_14,In_4509,In_1259);
nor U15 (N_15,In_627,In_3395);
or U16 (N_16,In_3420,In_4219);
xnor U17 (N_17,In_2560,In_3838);
and U18 (N_18,In_3939,In_3217);
or U19 (N_19,In_3870,In_1698);
nor U20 (N_20,In_3809,In_2945);
or U21 (N_21,In_2882,In_3678);
and U22 (N_22,In_345,In_3251);
nor U23 (N_23,In_1656,In_3575);
nand U24 (N_24,In_3474,In_870);
and U25 (N_25,In_3057,In_1458);
and U26 (N_26,In_427,In_4223);
xor U27 (N_27,In_984,In_1542);
and U28 (N_28,In_1235,In_66);
and U29 (N_29,In_3790,In_2496);
or U30 (N_30,In_921,In_4804);
xor U31 (N_31,In_2043,In_380);
nor U32 (N_32,In_3236,In_1596);
nand U33 (N_33,In_4667,In_3977);
or U34 (N_34,In_1285,In_130);
and U35 (N_35,In_2008,In_3259);
nand U36 (N_36,In_3618,In_3098);
xnor U37 (N_37,In_316,In_3644);
nor U38 (N_38,In_2565,In_2341);
nand U39 (N_39,In_2920,In_758);
nor U40 (N_40,In_4843,In_1992);
nor U41 (N_41,In_1647,In_1104);
nor U42 (N_42,In_4955,In_2388);
nor U43 (N_43,In_3442,In_4847);
nand U44 (N_44,In_3757,In_559);
nor U45 (N_45,In_1303,In_4685);
nor U46 (N_46,In_4810,In_1484);
or U47 (N_47,In_39,In_4424);
nor U48 (N_48,In_985,In_403);
and U49 (N_49,In_2073,In_4606);
and U50 (N_50,In_1167,In_1543);
nand U51 (N_51,In_4489,In_3325);
and U52 (N_52,In_1035,In_2364);
and U53 (N_53,In_4016,In_2527);
nand U54 (N_54,In_4011,In_2475);
nand U55 (N_55,In_386,In_567);
and U56 (N_56,In_1398,In_3907);
xnor U57 (N_57,In_1498,In_4944);
nand U58 (N_58,In_3399,In_4739);
and U59 (N_59,In_2725,In_4576);
nand U60 (N_60,In_2044,In_2233);
and U61 (N_61,In_4942,In_1881);
xor U62 (N_62,In_2023,In_1293);
and U63 (N_63,In_2643,In_4112);
xor U64 (N_64,In_1945,In_4373);
xor U65 (N_65,In_4529,In_1297);
xnor U66 (N_66,In_3211,In_2606);
nor U67 (N_67,In_317,In_385);
nand U68 (N_68,In_3263,In_3924);
and U69 (N_69,In_957,In_4567);
nand U70 (N_70,In_4873,In_397);
nand U71 (N_71,In_2990,In_2720);
nand U72 (N_72,In_3178,In_107);
or U73 (N_73,In_125,In_222);
or U74 (N_74,In_3514,In_1416);
nor U75 (N_75,In_4032,In_4022);
xor U76 (N_76,In_4784,In_516);
or U77 (N_77,In_4494,In_4840);
nor U78 (N_78,In_4959,In_425);
or U79 (N_79,In_3275,In_2531);
and U80 (N_80,In_2052,In_4409);
or U81 (N_81,In_1313,In_1646);
nor U82 (N_82,In_578,In_4599);
or U83 (N_83,In_584,In_2571);
nand U84 (N_84,In_2183,In_4287);
nor U85 (N_85,In_1765,In_3922);
nor U86 (N_86,In_1162,In_2890);
or U87 (N_87,In_3051,In_1770);
nand U88 (N_88,In_2280,In_3620);
xnor U89 (N_89,In_3602,In_1210);
and U90 (N_90,In_3635,In_4423);
nand U91 (N_91,In_1125,In_3680);
nor U92 (N_92,In_2817,In_2141);
nor U93 (N_93,In_4688,In_3883);
xor U94 (N_94,In_3951,In_3265);
and U95 (N_95,In_1304,In_1787);
and U96 (N_96,In_4607,In_2088);
or U97 (N_97,In_2366,In_954);
nor U98 (N_98,In_895,In_3455);
or U99 (N_99,In_866,In_445);
nor U100 (N_100,In_4293,In_1551);
nor U101 (N_101,In_570,In_4181);
nand U102 (N_102,In_3624,In_2266);
and U103 (N_103,In_4258,In_2419);
or U104 (N_104,In_1160,In_4900);
xor U105 (N_105,In_3535,In_3297);
nand U106 (N_106,In_1588,In_3459);
nor U107 (N_107,In_3498,In_638);
or U108 (N_108,In_3414,In_844);
or U109 (N_109,In_4341,In_3106);
nand U110 (N_110,In_3833,In_3955);
nand U111 (N_111,In_3091,In_1080);
or U112 (N_112,In_2328,In_872);
or U113 (N_113,In_736,In_2542);
xnor U114 (N_114,In_3811,In_4918);
xor U115 (N_115,In_373,In_4019);
nand U116 (N_116,In_3341,In_2440);
or U117 (N_117,In_9,In_1119);
nand U118 (N_118,In_2988,In_95);
xnor U119 (N_119,In_591,In_3795);
nor U120 (N_120,In_3377,In_1846);
or U121 (N_121,In_84,In_3042);
nor U122 (N_122,In_4363,In_4389);
nand U123 (N_123,In_147,In_4822);
and U124 (N_124,In_2710,In_1217);
nand U125 (N_125,In_928,In_4943);
and U126 (N_126,In_1287,In_268);
nand U127 (N_127,In_4305,In_230);
xnor U128 (N_128,In_3666,In_2895);
or U129 (N_129,In_1307,In_4296);
and U130 (N_130,In_3534,In_3376);
xor U131 (N_131,In_3486,In_1668);
xnor U132 (N_132,In_3787,In_2788);
or U133 (N_133,In_1037,In_1790);
and U134 (N_134,In_4037,In_2228);
xnor U135 (N_135,In_3643,In_3664);
xnor U136 (N_136,In_1174,In_2463);
nor U137 (N_137,In_4252,In_1366);
nor U138 (N_138,In_3723,In_4745);
xor U139 (N_139,In_530,In_1764);
and U140 (N_140,In_2842,In_3820);
nand U141 (N_141,In_2167,In_4445);
and U142 (N_142,In_1346,In_4267);
and U143 (N_143,In_2264,In_2768);
xnor U144 (N_144,In_1879,In_3957);
or U145 (N_145,In_1394,In_935);
xnor U146 (N_146,In_117,In_1150);
xnor U147 (N_147,In_1888,In_3345);
xor U148 (N_148,In_3765,In_577);
nand U149 (N_149,In_4491,In_3659);
or U150 (N_150,In_1864,In_4613);
and U151 (N_151,In_3167,In_2570);
nand U152 (N_152,In_4141,In_4909);
nor U153 (N_153,In_2752,In_1839);
xor U154 (N_154,In_2513,In_3815);
nand U155 (N_155,In_632,In_3216);
nand U156 (N_156,In_917,In_4973);
xnor U157 (N_157,In_2005,In_1679);
nand U158 (N_158,In_4628,In_3172);
or U159 (N_159,In_4303,In_269);
nand U160 (N_160,In_353,In_3309);
or U161 (N_161,In_1728,In_3674);
nor U162 (N_162,In_4055,In_1612);
xnor U163 (N_163,In_2201,In_1221);
xor U164 (N_164,In_2398,In_701);
or U165 (N_165,In_2405,In_1723);
nand U166 (N_166,In_3403,In_3841);
and U167 (N_167,In_1384,In_3590);
and U168 (N_168,In_978,In_2179);
or U169 (N_169,In_4492,In_4686);
nand U170 (N_170,In_1011,In_473);
nand U171 (N_171,In_2171,In_2604);
or U172 (N_172,In_3565,In_261);
xnor U173 (N_173,In_4856,In_1169);
or U174 (N_174,In_743,In_2071);
xnor U175 (N_175,In_1324,In_650);
or U176 (N_176,In_2656,In_1933);
and U177 (N_177,In_3195,In_4525);
or U178 (N_178,In_1655,In_4538);
nand U179 (N_179,In_4772,In_4937);
or U180 (N_180,In_3385,In_2355);
or U181 (N_181,In_3166,In_2060);
or U182 (N_182,In_391,In_4493);
and U183 (N_183,In_526,In_140);
or U184 (N_184,In_4753,In_441);
xnor U185 (N_185,In_3492,In_3874);
and U186 (N_186,In_1461,In_1318);
nand U187 (N_187,In_4165,In_1623);
xor U188 (N_188,In_1152,In_3701);
nand U189 (N_189,In_2674,In_3721);
xnor U190 (N_190,In_2931,In_4895);
nor U191 (N_191,In_3884,In_2098);
xnor U192 (N_192,In_2787,In_4335);
xor U193 (N_193,In_4199,In_1493);
nand U194 (N_194,In_4440,In_3095);
and U195 (N_195,In_4820,In_1108);
or U196 (N_196,In_740,In_3857);
and U197 (N_197,In_1355,In_99);
and U198 (N_198,In_539,In_658);
nand U199 (N_199,In_1693,In_2711);
nand U200 (N_200,In_3580,In_2761);
xnor U201 (N_201,In_672,In_1424);
or U202 (N_202,In_1525,In_1031);
and U203 (N_203,In_3234,In_143);
nand U204 (N_204,In_2078,In_3375);
nand U205 (N_205,In_3261,In_155);
and U206 (N_206,In_811,In_4605);
or U207 (N_207,In_2629,In_3460);
or U208 (N_208,In_2899,In_3370);
xnor U209 (N_209,In_686,In_1727);
and U210 (N_210,In_479,In_1392);
and U211 (N_211,In_1752,In_2149);
nand U212 (N_212,In_4161,In_3039);
and U213 (N_213,In_4390,In_1476);
or U214 (N_214,In_3796,In_2411);
or U215 (N_215,In_3270,In_3224);
nor U216 (N_216,In_4831,In_1672);
and U217 (N_217,In_4534,In_3764);
xnor U218 (N_218,In_1595,In_4716);
xnor U219 (N_219,In_2451,In_2337);
xnor U220 (N_220,In_123,In_2982);
nor U221 (N_221,In_4782,In_887);
nor U222 (N_222,In_1280,In_202);
and U223 (N_223,In_2384,In_4428);
xor U224 (N_224,In_1956,In_295);
nand U225 (N_225,In_1910,In_2831);
nand U226 (N_226,In_4926,In_3513);
and U227 (N_227,In_242,In_4517);
or U228 (N_228,In_719,In_4325);
xnor U229 (N_229,In_1480,In_3777);
and U230 (N_230,In_3596,In_438);
and U231 (N_231,In_394,In_3452);
nand U232 (N_232,In_2491,In_829);
nor U233 (N_233,In_1795,In_1935);
nand U234 (N_234,In_1601,In_1204);
nor U235 (N_235,In_2404,In_4602);
xor U236 (N_236,In_2220,In_1252);
or U237 (N_237,In_4073,In_784);
or U238 (N_238,In_2443,In_1919);
nor U239 (N_239,In_1171,In_4408);
or U240 (N_240,In_52,In_1427);
and U241 (N_241,In_3927,In_1381);
nand U242 (N_242,In_2038,In_3406);
or U243 (N_243,In_3758,In_2639);
nor U244 (N_244,In_4150,In_3747);
or U245 (N_245,In_4496,In_1740);
and U246 (N_246,In_2198,In_1460);
xnor U247 (N_247,In_1946,In_617);
or U248 (N_248,In_3079,In_2243);
xor U249 (N_249,In_4687,In_318);
or U250 (N_250,In_2151,In_3024);
and U251 (N_251,In_3702,In_2454);
nor U252 (N_252,In_826,In_4903);
nand U253 (N_253,In_493,In_1456);
and U254 (N_254,In_3687,In_4899);
xor U255 (N_255,In_520,In_602);
or U256 (N_256,In_1486,In_630);
xnor U257 (N_257,In_4339,In_4755);
and U258 (N_258,In_694,In_3750);
xor U259 (N_259,In_2575,In_2122);
nor U260 (N_260,In_2836,In_4528);
or U261 (N_261,In_2278,In_1664);
xnor U262 (N_262,In_2354,In_2392);
nand U263 (N_263,In_849,In_3179);
nand U264 (N_264,In_2648,In_958);
nand U265 (N_265,In_4704,In_640);
nor U266 (N_266,In_4592,In_3527);
xnor U267 (N_267,In_4671,In_2336);
nand U268 (N_268,In_1418,In_943);
xnor U269 (N_269,In_426,In_34);
nand U270 (N_270,In_4561,In_4264);
or U271 (N_271,In_1818,In_1047);
nand U272 (N_272,In_2066,In_433);
nor U273 (N_273,In_1799,In_1468);
nor U274 (N_274,In_3262,In_1199);
nand U275 (N_275,In_4052,In_2964);
and U276 (N_276,In_2777,In_3731);
nor U277 (N_277,In_273,In_1531);
xnor U278 (N_278,In_2323,In_1257);
xor U279 (N_279,In_288,In_4164);
and U280 (N_280,In_1220,In_4169);
nand U281 (N_281,In_976,In_4829);
nand U282 (N_282,In_4725,In_2692);
and U283 (N_283,In_680,In_190);
nand U284 (N_284,In_3361,In_457);
xnor U285 (N_285,In_2174,In_1658);
nor U286 (N_286,In_963,In_1262);
and U287 (N_287,In_2321,In_3491);
or U288 (N_288,In_2838,In_3537);
or U289 (N_289,In_3348,In_4066);
and U290 (N_290,In_2103,In_2079);
or U291 (N_291,In_660,In_4781);
nand U292 (N_292,In_3133,In_1943);
xnor U293 (N_293,In_1407,In_4844);
or U294 (N_294,In_3577,In_1576);
or U295 (N_295,In_2507,In_661);
and U296 (N_296,In_2846,In_1213);
nor U297 (N_297,In_1344,In_2640);
or U298 (N_298,In_470,In_2285);
nand U299 (N_299,In_1620,In_2024);
nor U300 (N_300,In_3672,In_615);
or U301 (N_301,In_1907,In_4570);
and U302 (N_302,In_3240,In_2632);
or U303 (N_303,In_3660,In_3165);
and U304 (N_304,In_885,In_2153);
nand U305 (N_305,In_2793,In_128);
nor U306 (N_306,In_197,In_4783);
xor U307 (N_307,In_1721,In_2891);
nor U308 (N_308,In_874,In_601);
nor U309 (N_309,In_1008,In_4524);
nand U310 (N_310,In_1863,In_194);
nand U311 (N_311,In_1944,In_2090);
nor U312 (N_312,In_2946,In_800);
xnor U313 (N_313,In_3778,In_2327);
or U314 (N_314,In_646,In_4385);
xnor U315 (N_315,In_4996,In_2934);
and U316 (N_316,In_1173,In_819);
nor U317 (N_317,In_522,In_2998);
xor U318 (N_318,In_4119,In_301);
xnor U319 (N_319,In_1296,In_4636);
xnor U320 (N_320,In_1995,In_3825);
nor U321 (N_321,In_48,In_384);
or U322 (N_322,In_2340,In_4029);
or U323 (N_323,In_767,In_1265);
or U324 (N_324,In_692,In_3576);
xor U325 (N_325,In_2330,In_673);
xnor U326 (N_326,In_3049,In_1735);
nor U327 (N_327,In_1306,In_4439);
nor U328 (N_328,In_1014,In_3071);
nor U329 (N_329,In_3302,In_2551);
nor U330 (N_330,In_3004,In_4038);
or U331 (N_331,In_36,In_1488);
and U332 (N_332,In_4482,In_4463);
nor U333 (N_333,In_746,In_1283);
nor U334 (N_334,In_1238,In_2203);
and U335 (N_335,In_284,In_3061);
nand U336 (N_336,In_897,In_4194);
xor U337 (N_337,In_1966,In_98);
or U338 (N_338,In_2143,In_3303);
xor U339 (N_339,In_1718,In_2262);
xor U340 (N_340,In_2470,In_4379);
xnor U341 (N_341,In_4545,In_893);
nand U342 (N_342,In_765,In_4604);
or U343 (N_343,In_3917,In_3502);
or U344 (N_344,In_4751,In_3102);
or U345 (N_345,In_4421,In_1836);
or U346 (N_346,In_3,In_880);
nor U347 (N_347,In_1783,In_2509);
or U348 (N_348,In_4794,In_1018);
nor U349 (N_349,In_1900,In_1807);
nor U350 (N_350,In_4458,In_2095);
or U351 (N_351,In_1072,In_3914);
and U352 (N_352,In_3285,In_4234);
or U353 (N_353,In_4283,In_3636);
and U354 (N_354,In_1625,In_1228);
or U355 (N_355,In_3208,In_4912);
nor U356 (N_356,In_2400,In_3794);
nand U357 (N_357,In_463,In_1111);
nand U358 (N_358,In_81,In_422);
xor U359 (N_359,In_1885,In_4091);
nand U360 (N_360,In_3305,In_1560);
nor U361 (N_361,In_2974,In_171);
xor U362 (N_362,In_282,In_232);
xor U363 (N_363,In_3707,In_1290);
and U364 (N_364,In_2414,In_1203);
and U365 (N_365,In_3490,In_2663);
and U366 (N_366,In_752,In_1106);
xor U367 (N_367,In_2635,In_657);
and U368 (N_368,In_4646,In_3688);
nor U369 (N_369,In_240,In_1877);
or U370 (N_370,In_3669,In_1785);
xnor U371 (N_371,In_4789,In_3868);
and U372 (N_372,In_2652,In_3813);
nand U373 (N_373,In_2295,In_820);
xnor U374 (N_374,In_3965,In_3097);
xor U375 (N_375,In_3233,In_2703);
xnor U376 (N_376,In_3088,In_276);
or U377 (N_377,In_2549,In_1929);
nand U378 (N_378,In_1871,In_3926);
nand U379 (N_379,In_4564,In_4707);
nor U380 (N_380,In_2436,In_448);
and U381 (N_381,In_3230,In_4085);
nand U382 (N_382,In_4139,In_2132);
xor U383 (N_383,In_1058,In_351);
nand U384 (N_384,In_179,In_4625);
or U385 (N_385,In_541,In_2284);
and U386 (N_386,In_2181,In_3495);
nor U387 (N_387,In_2630,In_1685);
xnor U388 (N_388,In_2784,In_4519);
and U389 (N_389,In_2863,In_2775);
nand U390 (N_390,In_2795,In_2929);
or U391 (N_391,In_2601,In_32);
or U392 (N_392,In_2274,In_413);
nor U393 (N_393,In_4611,In_3196);
nand U394 (N_394,In_4365,In_2221);
nor U395 (N_395,In_3480,In_2806);
nand U396 (N_396,In_3276,In_3013);
nor U397 (N_397,In_1939,In_2819);
and U398 (N_398,In_996,In_1826);
and U399 (N_399,In_2594,In_361);
nor U400 (N_400,In_2852,In_4936);
xnor U401 (N_401,In_2033,In_1261);
or U402 (N_402,In_4042,In_2712);
nand U403 (N_403,In_2681,In_2086);
xor U404 (N_404,In_990,In_821);
xnor U405 (N_405,In_279,In_4907);
nor U406 (N_406,In_2456,In_4076);
nand U407 (N_407,In_2238,In_1808);
xnor U408 (N_408,In_515,In_2433);
xor U409 (N_409,In_841,In_118);
or U410 (N_410,In_3078,In_1399);
xnor U411 (N_411,In_387,In_1409);
nor U412 (N_412,In_2651,In_1163);
nand U413 (N_413,In_4025,In_371);
nand U414 (N_414,In_4040,In_3437);
and U415 (N_415,In_573,In_4004);
xnor U416 (N_416,In_4930,In_4653);
nand U417 (N_417,In_210,In_2961);
and U418 (N_418,In_4785,In_4284);
xnor U419 (N_419,In_4118,In_1558);
xor U420 (N_420,In_761,In_599);
nor U421 (N_421,In_388,In_964);
nor U422 (N_422,In_3173,In_1385);
and U423 (N_423,In_1295,In_4833);
or U424 (N_424,In_1547,In_2448);
xor U425 (N_425,In_2845,In_3632);
and U426 (N_426,In_4121,In_4795);
and U427 (N_427,In_4897,In_3083);
xor U428 (N_428,In_3626,In_3510);
nor U429 (N_429,In_2807,In_216);
xor U430 (N_430,In_2857,In_734);
nor U431 (N_431,In_3246,In_1237);
or U432 (N_432,In_3554,In_1048);
nor U433 (N_433,In_595,In_3337);
xnor U434 (N_434,In_3328,In_3068);
and U435 (N_435,In_311,In_431);
nor U436 (N_436,In_3372,In_2449);
or U437 (N_437,In_2661,In_4557);
nor U438 (N_438,In_2854,In_1984);
and U439 (N_439,In_2435,In_484);
xor U440 (N_440,In_2734,In_1040);
nor U441 (N_441,In_2403,In_3973);
nand U442 (N_442,In_3402,In_183);
xor U443 (N_443,In_667,In_1338);
or U444 (N_444,In_2772,In_177);
nand U445 (N_445,In_4885,In_4680);
nand U446 (N_446,In_793,In_2347);
xor U447 (N_447,In_1825,In_676);
xnor U448 (N_448,In_2461,In_967);
nor U449 (N_449,In_3988,In_3283);
nand U450 (N_450,In_3836,In_525);
xnor U451 (N_451,In_3053,In_135);
xnor U452 (N_452,In_225,In_2204);
nor U453 (N_453,In_4453,In_1586);
or U454 (N_454,In_2779,In_1082);
nor U455 (N_455,In_2893,In_30);
or U456 (N_456,In_1365,In_1154);
nand U457 (N_457,In_4971,In_2363);
and U458 (N_458,In_2232,In_589);
nand U459 (N_459,In_2995,In_3871);
or U460 (N_460,In_4270,In_1131);
nor U461 (N_461,In_1896,In_993);
and U462 (N_462,In_3999,In_4244);
and U463 (N_463,In_339,In_4009);
and U464 (N_464,In_1834,In_3819);
or U465 (N_465,In_3709,In_2365);
and U466 (N_466,In_4742,In_2120);
nor U467 (N_467,In_228,In_2986);
or U468 (N_468,In_3176,In_605);
nand U469 (N_469,In_3256,In_4413);
xnor U470 (N_470,In_3799,In_1076);
nand U471 (N_471,In_1005,In_4103);
nor U472 (N_472,In_1532,In_2447);
or U473 (N_473,In_1109,In_280);
nand U474 (N_474,In_499,In_804);
nor U475 (N_475,In_1714,In_294);
or U476 (N_476,In_2760,In_908);
xnor U477 (N_477,In_560,In_332);
nand U478 (N_478,In_2292,In_1245);
nand U479 (N_479,In_3986,In_540);
xnor U480 (N_480,In_1107,In_2291);
or U481 (N_481,In_1886,In_1774);
and U482 (N_482,In_2125,In_961);
nand U483 (N_483,In_3096,In_1800);
nand U484 (N_484,In_980,In_3476);
or U485 (N_485,In_4105,In_4449);
nand U486 (N_486,In_2586,In_313);
xor U487 (N_487,In_3950,In_4759);
xnor U488 (N_488,In_2145,In_3422);
nand U489 (N_489,In_4887,In_1861);
nand U490 (N_490,In_3921,In_3899);
and U491 (N_491,In_780,In_3915);
nand U492 (N_492,In_1694,In_2916);
nand U493 (N_493,In_3613,In_3638);
xnor U494 (N_494,In_2165,In_1433);
xnor U495 (N_495,In_1641,In_2526);
nor U496 (N_496,In_2706,In_1909);
nor U497 (N_497,In_2563,In_2210);
nor U498 (N_498,In_3280,In_2927);
nand U499 (N_499,In_4371,In_529);
and U500 (N_500,In_46,In_843);
and U501 (N_501,In_4929,In_4441);
and U502 (N_502,In_4036,In_1786);
nand U503 (N_503,In_2446,In_2896);
nor U504 (N_504,In_4530,In_3858);
or U505 (N_505,In_1027,In_1211);
and U506 (N_506,In_226,In_2708);
nand U507 (N_507,In_4736,In_417);
nand U508 (N_508,In_2673,In_970);
xor U509 (N_509,In_2160,In_472);
and U510 (N_510,In_1371,In_428);
nand U511 (N_511,In_1556,In_2993);
xor U512 (N_512,In_3209,In_4477);
or U513 (N_513,In_999,In_2762);
and U514 (N_514,In_1396,In_4768);
xor U515 (N_515,In_4853,In_3953);
nand U516 (N_516,In_2680,In_4624);
and U517 (N_517,In_1229,In_1678);
nand U518 (N_518,In_1243,In_2359);
xnor U519 (N_519,In_1233,In_945);
nor U520 (N_520,In_4859,In_2387);
or U521 (N_521,In_914,In_3839);
nand U522 (N_522,In_3076,In_2809);
xor U523 (N_523,In_4582,In_4549);
nor U524 (N_524,In_2466,In_1294);
xnor U525 (N_525,In_4865,In_730);
nand U526 (N_526,In_3356,In_2385);
nor U527 (N_527,In_44,In_149);
or U528 (N_528,In_2195,In_3142);
nand U529 (N_529,In_1999,In_4849);
nor U530 (N_530,In_3144,In_3808);
or U531 (N_531,In_468,In_3279);
nand U532 (N_532,In_1059,In_4823);
or U533 (N_533,In_4532,In_467);
nand U534 (N_534,In_1386,In_2245);
nand U535 (N_535,In_3901,In_4372);
or U536 (N_536,In_633,In_3594);
nand U537 (N_537,In_703,In_1206);
xor U538 (N_538,In_170,In_4863);
nor U539 (N_539,In_1156,In_139);
nor U540 (N_540,In_2967,In_2825);
and U541 (N_541,In_642,In_1815);
and U542 (N_542,In_4975,In_852);
or U543 (N_543,In_3062,In_176);
or U544 (N_544,In_801,In_831);
and U545 (N_545,In_1497,In_1135);
or U546 (N_546,In_4522,In_2082);
nand U547 (N_547,In_4107,In_439);
or U548 (N_548,In_2914,In_3340);
nor U549 (N_549,In_1591,In_542);
xor U550 (N_550,In_2031,In_4803);
xor U551 (N_551,In_4750,In_1375);
xnor U552 (N_552,In_3471,In_3300);
nor U553 (N_553,In_3749,In_3605);
or U554 (N_554,In_2287,In_1747);
nand U555 (N_555,In_3508,In_186);
or U556 (N_556,In_1500,In_4343);
nor U557 (N_557,In_4217,In_4210);
nor U558 (N_558,In_1358,In_1506);
nand U559 (N_559,In_2276,In_1938);
xnor U560 (N_560,In_3431,In_1932);
and U561 (N_561,In_4035,In_3706);
nor U562 (N_562,In_4497,In_93);
nand U563 (N_563,In_3368,In_1853);
and U564 (N_564,In_3824,In_73);
xor U565 (N_565,In_2847,In_3075);
nor U566 (N_566,In_4726,In_1134);
xnor U567 (N_567,In_383,In_3628);
nor U568 (N_568,In_369,In_802);
xnor U569 (N_569,In_15,In_481);
or U570 (N_570,In_60,In_4550);
nor U571 (N_571,In_2345,In_1122);
nor U572 (N_572,In_2441,In_1833);
nand U573 (N_573,In_2100,In_247);
nand U574 (N_574,In_1904,In_1382);
and U575 (N_575,In_20,In_2667);
xnor U576 (N_576,In_1844,In_912);
nand U577 (N_577,In_1289,In_864);
and U578 (N_578,In_552,In_3312);
xor U579 (N_579,In_3383,In_4898);
nor U580 (N_580,In_1652,In_4136);
or U581 (N_581,In_3542,In_4488);
nor U582 (N_582,In_944,In_2792);
and U583 (N_583,In_2745,In_451);
nand U584 (N_584,In_3035,In_4867);
nor U585 (N_585,In_1611,In_2131);
nand U586 (N_586,In_4732,In_4817);
xor U587 (N_587,In_248,In_1996);
xnor U588 (N_588,In_3410,In_1251);
xnor U589 (N_589,In_586,In_4559);
xor U590 (N_590,In_582,In_2397);
or U591 (N_591,In_1811,In_4146);
or U592 (N_592,In_368,In_4574);
or U593 (N_593,In_4357,In_4641);
and U594 (N_594,In_1136,In_1766);
xnor U595 (N_595,In_2976,In_4130);
or U596 (N_596,In_1224,In_3609);
nand U597 (N_597,In_4008,In_3805);
nand U598 (N_598,In_1132,In_4923);
and U599 (N_599,In_3289,In_2128);
nand U600 (N_600,In_3245,In_713);
xor U601 (N_601,In_3132,In_1585);
or U602 (N_602,In_2267,In_2334);
and U603 (N_603,In_779,In_2413);
nand U604 (N_604,In_1016,In_1299);
or U605 (N_605,In_3159,In_3016);
nand U606 (N_606,In_3363,In_3568);
nand U607 (N_607,In_153,In_4718);
and U608 (N_608,In_4527,In_2362);
and U609 (N_609,In_1146,In_3685);
and U610 (N_610,In_4498,In_2492);
nand U611 (N_611,In_4526,In_822);
nand U612 (N_612,In_2063,In_1390);
nor U613 (N_613,In_4500,In_1415);
or U614 (N_614,In_2707,In_1600);
or U615 (N_615,In_3732,In_4190);
nand U616 (N_616,In_2780,In_3123);
or U617 (N_617,In_3155,In_4342);
nor U618 (N_618,In_927,In_937);
nand U619 (N_619,In_4003,In_535);
and U620 (N_620,In_2240,In_3791);
nor U621 (N_621,In_1621,In_3017);
xor U622 (N_622,In_1510,In_2175);
nor U623 (N_623,In_4154,In_1868);
or U624 (N_624,In_3093,In_3238);
xnor U625 (N_625,In_1100,In_700);
xor U626 (N_626,In_2331,In_1515);
and U627 (N_627,In_1548,In_1196);
and U628 (N_628,In_1278,In_2423);
or U629 (N_629,In_4705,In_785);
xnor U630 (N_630,In_1631,In_2172);
or U631 (N_631,In_1086,In_4935);
xnor U632 (N_632,In_828,In_593);
or U633 (N_633,In_2670,In_2984);
nand U634 (N_634,In_4106,In_4855);
nor U635 (N_635,In_1639,In_4432);
nor U636 (N_636,In_2932,In_4215);
xnor U637 (N_637,In_4192,In_2089);
nand U638 (N_638,In_689,In_1389);
and U639 (N_639,In_3320,In_3105);
or U640 (N_640,In_2273,In_968);
xnor U641 (N_641,In_1260,In_4544);
xnor U642 (N_642,In_1197,In_2268);
or U643 (N_643,In_3570,In_4170);
and U644 (N_644,In_3031,In_4610);
or U645 (N_645,In_1580,In_698);
xor U646 (N_646,In_2718,In_4661);
and U647 (N_647,In_4020,In_757);
nor U648 (N_648,In_2498,In_4983);
nor U649 (N_649,In_4213,In_2704);
xor U650 (N_650,In_111,In_342);
and U651 (N_651,In_3984,In_4674);
and U652 (N_652,In_3298,In_2558);
or U653 (N_653,In_4239,In_206);
xnor U654 (N_654,In_3864,In_1773);
nand U655 (N_655,In_3656,In_733);
xor U656 (N_656,In_2641,In_1226);
or U657 (N_657,In_4276,In_2649);
nor U658 (N_658,In_4792,In_3475);
xor U659 (N_659,In_3737,In_7);
xor U660 (N_660,In_4336,In_3336);
or U661 (N_661,In_2083,In_414);
or U662 (N_662,In_2117,In_4033);
and U663 (N_663,In_429,In_1269);
or U664 (N_664,In_4122,In_2783);
or U665 (N_665,In_2190,In_3872);
and U666 (N_666,In_4764,In_3330);
nor U667 (N_667,In_3277,In_4345);
nand U668 (N_668,In_1855,In_1145);
nand U669 (N_669,In_1437,In_580);
or U670 (N_670,In_3009,In_2081);
nand U671 (N_671,In_4395,In_2076);
or U672 (N_672,In_4241,In_4260);
nor U673 (N_673,In_4414,In_227);
nor U674 (N_674,In_4248,In_1737);
and U675 (N_675,In_1487,In_4761);
or U676 (N_676,In_4910,In_3162);
xnor U677 (N_677,In_2684,In_4311);
xnor U678 (N_678,In_4581,In_2960);
or U679 (N_679,In_3912,In_53);
nand U680 (N_680,In_4717,In_2878);
or U681 (N_681,In_3464,In_3432);
or U682 (N_682,In_3493,In_4518);
nor U683 (N_683,In_1449,In_2642);
or U684 (N_684,In_3533,In_3367);
or U685 (N_685,In_3900,In_4584);
or U686 (N_686,In_2064,In_3220);
xnor U687 (N_687,In_3503,In_3046);
xnor U688 (N_688,In_3905,In_1333);
and U689 (N_689,In_3553,In_951);
nand U690 (N_690,In_3916,In_4669);
or U691 (N_691,In_1034,In_2377);
nor U692 (N_692,In_1569,In_4352);
and U693 (N_693,In_2823,In_663);
and U694 (N_694,In_4562,In_4263);
xor U695 (N_695,In_4291,In_3047);
nor U696 (N_696,In_1388,In_1378);
xnor U697 (N_697,In_4832,In_3607);
nand U698 (N_698,In_156,In_3994);
xnor U699 (N_699,In_415,In_2593);
nor U700 (N_700,In_2111,In_4703);
and U701 (N_701,In_3793,In_1824);
nand U702 (N_702,In_4153,In_1875);
nand U703 (N_703,In_3895,In_1521);
xnor U704 (N_704,In_4658,In_3980);
nand U705 (N_705,In_704,In_4858);
and U706 (N_706,In_1562,In_4798);
and U707 (N_707,In_4690,In_4182);
or U708 (N_708,In_4741,In_3719);
nor U709 (N_709,In_753,In_102);
or U710 (N_710,In_4196,In_2314);
xor U711 (N_711,In_1127,In_2900);
nor U712 (N_712,In_608,In_722);
or U713 (N_713,In_168,In_2555);
and U714 (N_714,In_3426,In_4368);
and U715 (N_715,In_2477,In_3110);
nand U716 (N_716,In_4979,In_859);
and U717 (N_717,In_4460,In_1719);
nand U718 (N_718,In_61,In_4344);
xor U719 (N_719,In_4444,In_4787);
xor U720 (N_720,In_3177,In_1993);
nor U721 (N_721,In_1748,In_2009);
and U722 (N_722,In_742,In_953);
xor U723 (N_723,In_4516,In_2026);
and U724 (N_724,In_452,In_4773);
nor U725 (N_725,In_1702,In_622);
or U726 (N_726,In_2415,In_4231);
or U727 (N_727,In_1592,In_1991);
nor U728 (N_728,In_1183,In_2004);
and U729 (N_729,In_2417,In_412);
nand U730 (N_730,In_2826,In_2156);
and U731 (N_731,In_842,In_2207);
xor U732 (N_732,In_4364,In_3911);
and U733 (N_733,In_791,In_3654);
nand U734 (N_734,In_783,In_119);
and U735 (N_735,In_3591,In_1634);
nor U736 (N_736,In_4589,In_3188);
nand U737 (N_737,In_2119,In_1329);
and U738 (N_738,In_2696,In_3954);
nor U739 (N_739,In_4242,In_4402);
or U740 (N_740,In_215,In_4665);
and U741 (N_741,In_697,In_4748);
and U742 (N_742,In_4968,In_1330);
nor U743 (N_743,In_2006,In_4848);
nor U744 (N_744,In_241,In_304);
and U745 (N_745,In_2740,In_1732);
and U746 (N_746,In_3023,In_4024);
and U747 (N_747,In_29,In_2770);
nor U748 (N_748,In_401,In_3018);
nor U749 (N_749,In_523,In_2810);
or U750 (N_750,In_916,In_3210);
nand U751 (N_751,In_1821,In_133);
xnor U752 (N_752,In_4997,In_4208);
and U753 (N_753,In_3308,In_347);
nor U754 (N_754,In_507,In_1974);
xnor U755 (N_755,In_2608,In_2540);
and U756 (N_756,In_4947,In_4513);
and U757 (N_757,In_1143,In_2074);
nand U758 (N_758,In_2296,In_4596);
or U759 (N_759,In_1019,In_3304);
nand U760 (N_760,In_2866,In_696);
and U761 (N_761,In_2937,In_896);
nand U762 (N_762,In_2102,In_3637);
and U763 (N_763,In_1376,In_1615);
xor U764 (N_764,In_2519,In_3323);
xnor U765 (N_765,In_4539,In_2450);
nand U766 (N_766,In_2728,In_1835);
nand U767 (N_767,In_2682,In_4790);
nand U768 (N_768,In_106,In_1198);
xor U769 (N_769,In_3048,In_3851);
nor U770 (N_770,In_4288,In_3511);
and U771 (N_771,In_3940,In_4499);
nor U772 (N_772,In_756,In_1186);
nand U773 (N_773,In_4649,In_4374);
or U774 (N_774,In_666,In_3840);
or U775 (N_775,In_4713,In_538);
nor U776 (N_776,In_1009,In_1325);
xnor U777 (N_777,In_3783,In_3499);
xor U778 (N_778,In_2325,In_4369);
xnor U779 (N_779,In_3512,In_3366);
or U780 (N_780,In_2989,In_2472);
or U781 (N_781,In_706,In_1955);
nor U782 (N_782,In_3065,In_1273);
or U783 (N_783,In_358,In_4827);
nor U784 (N_784,In_1589,In_4695);
nand U785 (N_785,In_3121,In_220);
nand U786 (N_786,In_1571,In_4648);
or U787 (N_787,In_3962,In_4974);
xor U788 (N_788,In_4456,In_1216);
and U789 (N_789,In_293,In_3751);
nand U790 (N_790,In_2909,In_2944);
nand U791 (N_791,In_3331,In_3552);
nor U792 (N_792,In_598,In_2832);
or U793 (N_793,In_4361,In_509);
and U794 (N_794,In_4088,In_4924);
nor U795 (N_795,In_356,In_1876);
nor U796 (N_796,In_4796,In_4386);
nand U797 (N_797,In_2583,In_1326);
nor U798 (N_798,In_4426,In_2374);
xnor U799 (N_799,In_360,In_4155);
and U800 (N_800,In_3784,In_3925);
nand U801 (N_801,In_3430,In_374);
nand U802 (N_802,In_4446,In_132);
nor U803 (N_803,In_2493,In_314);
and U804 (N_804,In_3154,In_4752);
xor U805 (N_805,In_64,In_4884);
and U806 (N_806,In_2749,In_930);
and U807 (N_807,In_3557,In_4028);
and U808 (N_808,In_2313,In_3978);
or U809 (N_809,In_3485,In_2155);
nand U810 (N_810,In_789,In_634);
or U811 (N_811,In_986,In_4230);
nand U812 (N_812,In_474,In_1367);
xnor U813 (N_813,In_1377,In_1742);
and U814 (N_814,In_2402,In_2425);
xnor U815 (N_815,In_4981,In_3436);
nand U816 (N_816,In_2613,In_1181);
nand U817 (N_817,In_1049,In_1518);
xnor U818 (N_818,In_1153,In_1412);
xnor U819 (N_819,In_4578,In_2822);
and U820 (N_820,In_1042,In_442);
or U821 (N_821,In_2304,In_1092);
nand U822 (N_822,In_4058,In_3547);
nand U823 (N_823,In_2512,In_4535);
xnor U824 (N_824,In_4870,In_1882);
or U825 (N_825,In_212,In_3716);
xnor U826 (N_826,In_281,In_3818);
nand U827 (N_827,In_3185,In_4200);
xnor U828 (N_828,In_2587,In_2061);
or U829 (N_829,In_847,In_298);
nor U830 (N_830,In_127,In_4422);
nor U831 (N_831,In_1331,In_4472);
or U832 (N_832,In_3129,In_2951);
nor U833 (N_833,In_4129,In_1889);
nor U834 (N_834,In_3489,In_3600);
or U835 (N_835,In_76,In_4697);
or U836 (N_836,In_2067,In_1253);
or U837 (N_837,In_88,In_2338);
and U838 (N_838,In_3441,In_3243);
xnor U839 (N_839,In_3421,In_581);
and U840 (N_840,In_1587,In_869);
or U841 (N_841,In_405,In_3322);
nand U842 (N_842,In_290,In_2802);
and U843 (N_843,In_3610,In_2590);
or U844 (N_844,In_366,In_809);
and U845 (N_845,In_2230,In_2835);
nor U846 (N_846,In_2372,In_1165);
nand U847 (N_847,In_1934,In_4958);
nand U848 (N_848,In_1653,In_2996);
nor U849 (N_849,In_424,In_3763);
or U850 (N_850,In_4204,In_725);
nand U851 (N_851,In_3135,In_2235);
xor U852 (N_852,In_89,In_3743);
xnor U853 (N_853,In_1662,In_1195);
xor U854 (N_854,In_2889,In_3956);
and U855 (N_855,In_2427,In_1772);
xor U856 (N_856,In_3997,In_2351);
and U857 (N_857,In_4046,In_747);
and U858 (N_858,In_1141,In_4202);
xor U859 (N_859,In_3351,In_3886);
xor U860 (N_860,In_3438,In_494);
and U861 (N_861,In_2529,In_3186);
or U862 (N_862,In_4877,In_1779);
and U863 (N_863,In_2778,In_400);
nor U864 (N_864,In_1947,In_447);
or U865 (N_865,In_1369,In_1520);
and U866 (N_866,In_3373,In_3295);
xor U867 (N_867,In_1172,In_4579);
and U868 (N_868,In_340,In_3045);
nor U869 (N_869,In_337,In_3271);
nand U870 (N_870,In_1431,In_3832);
and U871 (N_871,In_4317,In_174);
or U872 (N_872,In_878,In_115);
or U873 (N_873,In_4411,In_4249);
or U874 (N_874,In_3056,In_1832);
xnor U875 (N_875,In_2983,In_4128);
and U876 (N_876,In_4382,In_1892);
and U877 (N_877,In_2041,In_1263);
nor U878 (N_878,In_2283,In_2252);
xnor U879 (N_879,In_3720,In_229);
nor U880 (N_880,In_38,In_2097);
or U881 (N_881,In_2888,In_4960);
nor U882 (N_882,In_2538,In_4627);
or U883 (N_883,In_3880,In_4948);
and U884 (N_884,In_477,In_4443);
xor U885 (N_885,In_2368,In_2633);
xor U886 (N_886,In_3058,In_3803);
xnor U887 (N_887,In_2367,In_5);
nand U888 (N_888,In_169,In_3453);
or U889 (N_889,In_1060,In_3150);
xor U890 (N_890,In_4067,In_4434);
nor U891 (N_891,In_4466,In_3852);
nand U892 (N_892,In_72,In_3496);
nor U893 (N_893,In_2226,In_2380);
or U894 (N_894,In_204,In_1323);
and U895 (N_895,In_3477,In_85);
nor U896 (N_896,In_4079,In_4328);
xor U897 (N_897,In_4643,In_519);
and U898 (N_898,In_2219,In_1332);
or U899 (N_899,In_408,In_3396);
nor U900 (N_900,In_2504,In_3892);
nor U901 (N_901,In_837,In_4786);
and U902 (N_902,In_4490,In_3929);
nor U903 (N_903,In_3364,In_4915);
xor U904 (N_904,In_3500,In_4945);
and U905 (N_905,In_1013,In_3090);
or U906 (N_906,In_4081,In_1534);
or U907 (N_907,In_2113,In_365);
and U908 (N_908,In_4728,In_3319);
xor U909 (N_909,In_2329,In_727);
xnor U910 (N_910,In_2164,In_1317);
and U911 (N_911,In_2841,In_1894);
nor U912 (N_912,In_3587,In_1477);
xnor U913 (N_913,In_862,In_3705);
xnor U914 (N_914,In_4565,In_2689);
and U915 (N_915,In_2687,In_3022);
xor U916 (N_916,In_1915,In_2254);
nand U917 (N_917,In_1413,In_3352);
nand U918 (N_918,In_4427,In_1242);
and U919 (N_919,In_3903,In_4701);
xnor U920 (N_920,In_1067,In_203);
nor U921 (N_921,In_4044,In_3952);
nand U922 (N_922,In_4684,In_795);
nor U923 (N_923,In_1321,In_2046);
or U924 (N_924,In_2458,In_1980);
nand U925 (N_925,In_1789,In_1754);
nand U926 (N_926,In_1715,In_807);
or U927 (N_927,In_3291,In_1470);
xnor U928 (N_928,In_2615,In_3543);
or U929 (N_929,In_443,In_3404);
xor U930 (N_930,In_3286,In_1436);
and U931 (N_931,In_3936,In_1960);
nand U932 (N_932,In_4295,In_4407);
or U933 (N_933,In_4660,In_80);
or U934 (N_934,In_833,In_2409);
and U935 (N_935,In_262,In_2379);
xnor U936 (N_936,In_1023,In_4127);
and U937 (N_937,In_2892,In_3028);
xor U938 (N_938,In_4874,In_1114);
nand U939 (N_939,In_2533,In_2755);
xnor U940 (N_940,In_270,In_25);
xor U941 (N_941,In_185,In_3860);
xnor U942 (N_942,In_3450,In_250);
and U943 (N_943,In_856,In_4433);
nand U944 (N_944,In_258,In_4259);
nor U945 (N_945,In_2482,In_2196);
or U946 (N_946,In_4419,In_671);
nand U947 (N_947,In_3479,In_1570);
and U948 (N_948,In_4801,In_2525);
nor U949 (N_949,In_1644,In_2189);
xor U950 (N_950,In_4125,In_145);
nand U951 (N_951,In_3002,In_2199);
and U952 (N_952,In_1255,In_218);
or U953 (N_953,In_96,In_4824);
xnor U954 (N_954,In_1439,In_421);
nor U955 (N_955,In_1032,In_1282);
xnor U956 (N_956,In_3223,In_3655);
xor U957 (N_957,In_716,In_2319);
nor U958 (N_958,In_574,In_544);
nand U959 (N_959,In_1190,In_2478);
xnor U960 (N_960,In_923,In_1465);
or U961 (N_961,In_2134,In_2879);
nor U962 (N_962,In_157,In_1138);
and U963 (N_963,In_3386,In_2473);
nand U964 (N_964,In_4507,In_3625);
xnor U965 (N_965,In_3111,In_2412);
or U966 (N_966,In_1391,In_2178);
nor U967 (N_967,In_1985,In_2194);
nand U968 (N_968,In_3200,In_4021);
nor U969 (N_969,In_3786,In_4240);
and U970 (N_970,In_3843,In_3682);
and U971 (N_971,In_309,In_4999);
nand U972 (N_972,In_1284,In_2801);
and U973 (N_973,In_4729,In_1387);
nor U974 (N_974,In_411,In_4465);
or U975 (N_975,In_2115,In_3411);
nor U976 (N_976,In_3055,In_4148);
nand U977 (N_977,In_2428,In_4980);
xor U978 (N_978,In_3579,In_3574);
xor U979 (N_979,In_2971,In_1673);
and U980 (N_980,In_338,In_3258);
xor U981 (N_981,In_4010,In_3647);
and U982 (N_982,In_4619,In_319);
xnor U983 (N_983,In_4151,In_2047);
xnor U984 (N_984,In_4447,In_3898);
nand U985 (N_985,In_3725,In_4448);
nand U986 (N_986,In_2936,In_4637);
and U987 (N_987,In_4857,In_1250);
nor U988 (N_988,In_37,In_1990);
nand U989 (N_989,In_3859,In_1775);
xor U990 (N_990,In_3698,In_1854);
xor U991 (N_991,In_4057,In_879);
or U992 (N_992,In_4595,In_2346);
or U993 (N_993,In_1362,In_571);
nor U994 (N_994,In_909,In_2013);
and U995 (N_995,In_748,In_2);
nor U996 (N_996,In_131,In_1360);
nand U997 (N_997,In_4800,In_770);
and U998 (N_998,In_623,In_4229);
xor U999 (N_999,In_4014,In_4939);
nor U1000 (N_1000,In_2992,In_1055);
xor U1001 (N_1001,In_1193,In_3744);
xor U1002 (N_1002,In_4555,In_2729);
xnor U1003 (N_1003,In_2070,In_1276);
nor U1004 (N_1004,In_3775,In_4754);
or U1005 (N_1005,In_3299,In_1666);
or U1006 (N_1006,In_4321,In_321);
nand U1007 (N_1007,In_1298,In_2940);
xnor U1008 (N_1008,In_4381,In_3445);
nand U1009 (N_1009,In_1767,In_1950);
nor U1010 (N_1010,In_154,In_955);
xor U1011 (N_1011,In_4255,In_4851);
and U1012 (N_1012,In_528,In_3695);
nand U1013 (N_1013,In_2877,In_938);
nand U1014 (N_1014,In_3797,In_3444);
or U1015 (N_1015,In_3700,In_1665);
or U1016 (N_1016,In_3287,In_2626);
xnor U1017 (N_1017,In_2962,In_549);
nand U1018 (N_1018,In_187,In_3968);
nor U1019 (N_1019,In_2213,In_2742);
or U1020 (N_1020,In_636,In_440);
nand U1021 (N_1021,In_2576,In_1530);
nand U1022 (N_1022,In_1079,In_4298);
or U1023 (N_1023,In_2099,In_1796);
nand U1024 (N_1024,In_4620,In_1478);
nand U1025 (N_1025,In_3466,In_2489);
and U1026 (N_1026,In_1707,In_2887);
nand U1027 (N_1027,In_899,In_3983);
or U1028 (N_1028,In_1450,In_4137);
nor U1029 (N_1029,In_4951,In_898);
nor U1030 (N_1030,In_3250,In_3329);
nand U1031 (N_1031,In_1528,In_4904);
or U1032 (N_1032,In_4740,In_3292);
and U1033 (N_1033,In_4712,In_3748);
nand U1034 (N_1034,In_4807,In_478);
xnor U1035 (N_1035,In_1760,In_2373);
or U1036 (N_1036,In_3573,In_1232);
nor U1037 (N_1037,In_3229,In_4949);
or U1038 (N_1038,In_4383,In_3310);
nor U1039 (N_1039,In_3708,In_2735);
xnor U1040 (N_1040,In_3889,In_1578);
nand U1041 (N_1041,In_2926,In_4133);
xnor U1042 (N_1042,In_3559,In_3100);
nor U1043 (N_1043,In_2335,In_2981);
or U1044 (N_1044,In_1339,In_4065);
or U1045 (N_1045,In_575,In_2607);
xor U1046 (N_1046,In_4990,In_4451);
nand U1047 (N_1047,In_4152,In_597);
or U1048 (N_1048,In_4332,In_3033);
nand U1049 (N_1049,In_2361,In_702);
nor U1050 (N_1050,In_2733,In_1803);
xnor U1051 (N_1051,In_1065,In_2855);
or U1052 (N_1052,In_547,In_4505);
and U1053 (N_1053,In_4431,In_2508);
xnor U1054 (N_1054,In_3268,In_1254);
nand U1055 (N_1055,In_136,In_3646);
xor U1056 (N_1056,In_256,In_3365);
nor U1057 (N_1057,In_1563,In_1869);
xnor U1058 (N_1058,In_2048,In_1709);
nand U1059 (N_1059,In_1577,In_40);
and U1060 (N_1060,In_419,In_4749);
xnor U1061 (N_1061,In_714,In_4308);
or U1062 (N_1062,In_3603,In_2833);
nor U1063 (N_1063,In_728,In_4896);
and U1064 (N_1064,In_2624,In_3673);
xnor U1065 (N_1065,In_51,In_911);
nor U1066 (N_1066,In_2691,In_4059);
or U1067 (N_1067,In_4304,In_2910);
xor U1068 (N_1068,In_1081,In_1268);
nor U1069 (N_1069,In_2218,In_1349);
nand U1070 (N_1070,In_3252,In_2269);
nand U1071 (N_1071,In_4060,In_711);
and U1072 (N_1072,In_1316,In_104);
nor U1073 (N_1073,In_652,In_129);
xor U1074 (N_1074,In_3992,In_1113);
and U1075 (N_1075,In_2326,In_4864);
nand U1076 (N_1076,In_1062,In_1849);
nand U1077 (N_1077,In_2769,In_3242);
nand U1078 (N_1078,In_1777,In_1151);
nand U1079 (N_1079,In_1605,In_569);
and U1080 (N_1080,In_3085,In_4738);
and U1081 (N_1081,In_688,In_2580);
and U1082 (N_1082,In_4310,In_2000);
xor U1083 (N_1083,In_3670,In_4455);
xnor U1084 (N_1084,In_4285,In_4116);
or U1085 (N_1085,In_3282,In_1912);
xor U1086 (N_1086,In_1969,In_4608);
xor U1087 (N_1087,In_3170,In_4617);
xnor U1088 (N_1088,In_1123,In_483);
nand U1089 (N_1089,In_271,In_988);
nand U1090 (N_1090,In_2012,In_1697);
nand U1091 (N_1091,In_2025,In_3691);
xnor U1092 (N_1092,In_1979,In_4839);
xor U1093 (N_1093,In_2383,In_4160);
or U1094 (N_1094,In_2611,In_2800);
nor U1095 (N_1095,In_1073,In_260);
or U1096 (N_1096,In_4788,In_4566);
and U1097 (N_1097,In_2080,In_2407);
or U1098 (N_1098,In_4318,In_3582);
nor U1099 (N_1099,In_3667,In_1852);
xnor U1100 (N_1100,In_1983,In_2591);
nand U1101 (N_1101,In_4501,In_4315);
and U1102 (N_1102,In_4911,In_2950);
nand U1103 (N_1103,In_1207,In_4193);
xor U1104 (N_1104,In_3000,In_381);
or U1105 (N_1105,In_1021,In_122);
or U1106 (N_1106,In_1649,In_4553);
nor U1107 (N_1107,In_3288,In_846);
nand U1108 (N_1108,In_1057,In_4113);
nand U1109 (N_1109,In_3782,In_4828);
nand U1110 (N_1110,In_1967,In_2873);
xor U1111 (N_1111,In_306,In_1078);
and U1112 (N_1112,In_1692,In_2834);
or U1113 (N_1113,In_2129,In_2827);
nor U1114 (N_1114,In_2050,In_3087);
nand U1115 (N_1115,In_2306,In_4536);
nor U1116 (N_1116,In_94,In_2483);
and U1117 (N_1117,In_3523,In_2432);
nor U1118 (N_1118,In_4104,In_2406);
nor U1119 (N_1119,In_4966,In_4708);
and U1120 (N_1120,In_624,In_33);
nor U1121 (N_1121,In_1246,In_2911);
or U1122 (N_1122,In_2184,In_890);
or U1123 (N_1123,In_751,In_291);
nor U1124 (N_1124,In_1003,In_492);
or U1125 (N_1125,In_3175,In_4114);
nand U1126 (N_1126,In_1372,In_2056);
or U1127 (N_1127,In_4632,In_3781);
and U1128 (N_1128,In_4437,In_3374);
or U1129 (N_1129,In_3651,In_3313);
nand U1130 (N_1130,In_735,In_2867);
nor U1131 (N_1131,In_3470,In_3584);
xor U1132 (N_1132,In_2602,In_2015);
and U1133 (N_1133,In_4086,In_1696);
nor U1134 (N_1134,In_2904,In_2700);
xnor U1135 (N_1135,In_877,In_4012);
nor U1136 (N_1136,In_2352,In_4586);
nand U1137 (N_1137,In_4206,In_4474);
or U1138 (N_1138,In_4590,In_4976);
and U1139 (N_1139,In_1363,In_4145);
xnor U1140 (N_1140,In_1526,In_2716);
or U1141 (N_1141,In_3273,In_3597);
xor U1142 (N_1142,In_1052,In_2453);
nor U1143 (N_1143,In_4868,In_771);
xor U1144 (N_1144,In_4978,In_1566);
nor U1145 (N_1145,In_3226,In_4850);
and U1146 (N_1146,In_2431,In_4228);
nand U1147 (N_1147,In_1494,In_4830);
nand U1148 (N_1148,In_1139,In_3454);
nor U1149 (N_1149,In_946,In_1383);
nor U1150 (N_1150,In_3893,In_1667);
xnor U1151 (N_1151,In_832,In_4183);
or U1152 (N_1152,In_159,In_2371);
nor U1153 (N_1153,In_3350,In_1336);
nand U1154 (N_1154,In_3931,In_2874);
or U1155 (N_1155,In_2055,In_2679);
xnor U1156 (N_1156,In_922,In_695);
or U1157 (N_1157,In_2471,In_382);
nor U1158 (N_1158,In_4573,In_78);
nand U1159 (N_1159,In_902,In_75);
xnor U1160 (N_1160,In_3774,In_3518);
nand U1161 (N_1161,In_4030,In_3623);
nand U1162 (N_1162,In_31,In_2469);
nand U1163 (N_1163,In_3094,In_362);
and U1164 (N_1164,In_213,In_446);
xnor U1165 (N_1165,In_3755,In_4639);
nand U1166 (N_1166,In_3714,In_1271);
nor U1167 (N_1167,In_330,In_2544);
or U1168 (N_1168,In_2256,In_1700);
xor U1169 (N_1169,In_1744,In_1902);
or U1170 (N_1170,In_1397,In_3563);
xor U1171 (N_1171,In_2124,In_3063);
nand U1172 (N_1172,In_3081,In_1098);
or U1173 (N_1173,In_1001,In_3696);
xnor U1174 (N_1174,In_982,In_4061);
nor U1175 (N_1175,In_1632,In_600);
or U1176 (N_1176,In_2690,In_901);
nor U1177 (N_1177,In_2534,In_3504);
nand U1178 (N_1178,In_3448,In_4711);
xor U1179 (N_1179,In_616,In_1725);
xor U1180 (N_1180,In_2973,In_3379);
and U1181 (N_1181,In_4053,In_1473);
or U1182 (N_1182,In_4541,In_4307);
xnor U1183 (N_1183,In_2087,In_3928);
nand U1184 (N_1184,In_1884,In_3650);
xnor U1185 (N_1185,In_2714,In_4256);
xor U1186 (N_1186,In_4612,In_2091);
xor U1187 (N_1187,In_4131,In_2121);
nor U1188 (N_1188,In_683,In_4623);
nand U1189 (N_1189,In_3541,In_2814);
or U1190 (N_1190,In_3164,In_2339);
nand U1191 (N_1191,In_886,In_349);
nor U1192 (N_1192,In_4436,In_2445);
xor U1193 (N_1193,In_257,In_1482);
and U1194 (N_1194,In_4203,In_193);
or U1195 (N_1195,In_690,In_86);
nor U1196 (N_1196,In_3169,In_3156);
xnor U1197 (N_1197,In_3967,In_1716);
nand U1198 (N_1198,In_3995,In_2943);
xor U1199 (N_1199,In_920,In_1837);
xnor U1200 (N_1200,In_22,In_2214);
xor U1201 (N_1201,In_4438,In_2719);
or U1202 (N_1202,In_4316,In_2035);
xor U1203 (N_1203,In_4245,In_4429);
and U1204 (N_1204,In_3652,In_3769);
and U1205 (N_1205,In_1567,In_918);
and U1206 (N_1206,In_4552,In_1776);
xnor U1207 (N_1207,In_2864,In_4156);
and U1208 (N_1208,In_126,In_3247);
or U1209 (N_1209,In_82,In_4892);
and U1210 (N_1210,In_3856,In_987);
and U1211 (N_1211,In_1309,In_2595);
nand U1212 (N_1212,In_1443,In_2668);
nor U1213 (N_1213,In_3943,In_1972);
nand U1214 (N_1214,In_2535,In_3433);
nor U1215 (N_1215,In_4294,In_3324);
or U1216 (N_1216,In_3235,In_3615);
or U1217 (N_1217,In_4919,In_4391);
or U1218 (N_1218,In_4743,In_2884);
xnor U1219 (N_1219,In_267,In_2618);
nor U1220 (N_1220,In_1794,In_3434);
and U1221 (N_1221,In_962,In_3506);
nor U1222 (N_1222,In_2567,In_2107);
nor U1223 (N_1223,In_2212,In_3128);
xor U1224 (N_1224,In_1051,In_934);
and U1225 (N_1225,In_2662,In_1215);
xor U1226 (N_1226,In_2997,In_1977);
or U1227 (N_1227,In_1859,In_4778);
xor U1228 (N_1228,In_2623,In_3228);
xor U1229 (N_1229,In_3307,In_3497);
and U1230 (N_1230,In_3338,In_4631);
xnor U1231 (N_1231,In_1357,In_3735);
or U1232 (N_1232,In_707,In_3740);
xor U1233 (N_1233,In_1435,In_4664);
and U1234 (N_1234,In_1184,In_4714);
and U1235 (N_1235,In_3902,In_323);
nand U1236 (N_1236,In_363,In_4286);
xor U1237 (N_1237,In_1116,In_1699);
xnor U1238 (N_1238,In_1638,In_1077);
xnor U1239 (N_1239,In_1438,In_209);
or U1240 (N_1240,In_3359,In_3427);
or U1241 (N_1241,In_2727,In_1457);
nor U1242 (N_1242,In_444,In_2391);
nand U1243 (N_1243,In_1805,In_277);
nor U1244 (N_1244,In_2744,In_4197);
xor U1245 (N_1245,In_2348,In_4710);
nand U1246 (N_1246,In_3469,In_2596);
and U1247 (N_1247,In_2307,In_1619);
and U1248 (N_1248,In_2741,In_2322);
xnor U1249 (N_1249,In_1225,In_3347);
xor U1250 (N_1250,In_1501,In_2462);
or U1251 (N_1251,In_3788,In_2468);
nand U1252 (N_1252,In_4502,In_4102);
xor U1253 (N_1253,In_4323,In_4852);
xnor U1254 (N_1254,In_3241,In_2239);
or U1255 (N_1255,In_500,In_4089);
or U1256 (N_1256,In_4626,In_4201);
nand U1257 (N_1257,In_1513,In_1370);
nor U1258 (N_1258,In_3745,In_3517);
xor U1259 (N_1259,In_4366,In_4290);
or U1260 (N_1260,In_4819,In_685);
and U1261 (N_1261,In_798,In_2353);
and U1262 (N_1262,In_2072,In_2868);
xnor U1263 (N_1263,In_3528,In_4142);
or U1264 (N_1264,In_3733,In_1085);
nor U1265 (N_1265,In_1177,In_1997);
or U1266 (N_1266,In_3494,In_4815);
nor U1267 (N_1267,In_1236,In_496);
xor U1268 (N_1268,In_1410,In_2484);
or U1269 (N_1269,In_2028,In_1584);
and U1270 (N_1270,In_1002,In_3718);
and U1271 (N_1271,In_4320,In_2299);
nor U1272 (N_1272,In_1155,In_3137);
nor U1273 (N_1273,In_1043,In_8);
nor U1274 (N_1274,In_4763,In_1568);
and U1275 (N_1275,In_865,In_4233);
nor U1276 (N_1276,In_2569,In_553);
nand U1277 (N_1277,In_195,In_4771);
xnor U1278 (N_1278,In_4218,In_2401);
nor U1279 (N_1279,In_3569,In_2020);
and U1280 (N_1280,In_2619,In_3008);
nand U1281 (N_1281,In_233,In_4927);
or U1282 (N_1282,In_4609,In_2612);
nor U1283 (N_1283,In_4077,In_26);
xnor U1284 (N_1284,In_709,In_3676);
and U1285 (N_1285,In_3964,In_327);
or U1286 (N_1286,In_3407,In_3727);
nor U1287 (N_1287,In_3181,In_626);
xor U1288 (N_1288,In_1681,In_2872);
or U1289 (N_1289,In_3641,In_2349);
xor U1290 (N_1290,In_884,In_3054);
nor U1291 (N_1291,In_259,In_1874);
nor U1292 (N_1292,In_3315,In_1348);
or U1293 (N_1293,In_3070,In_3069);
and U1294 (N_1294,In_3041,In_2279);
and U1295 (N_1295,In_4814,In_2803);
or U1296 (N_1296,In_2994,In_1479);
and U1297 (N_1297,In_4917,In_2919);
or U1298 (N_1298,In_1994,In_50);
nor U1299 (N_1299,In_4762,In_4412);
xor U1300 (N_1300,In_2108,In_2694);
xor U1301 (N_1301,In_3989,In_2675);
nand U1302 (N_1302,In_410,In_2722);
and U1303 (N_1303,In_4946,In_3710);
xnor U1304 (N_1304,In_3349,In_2837);
nand U1305 (N_1305,In_3734,In_3598);
nand U1306 (N_1306,In_1426,In_2094);
and U1307 (N_1307,In_816,In_4777);
or U1308 (N_1308,In_142,In_141);
xnor U1309 (N_1309,In_4925,In_769);
and U1310 (N_1310,In_2799,In_4678);
and U1311 (N_1311,In_949,In_2939);
nor U1312 (N_1312,In_3354,In_848);
nand U1313 (N_1313,In_4396,In_2399);
nand U1314 (N_1314,In_845,In_1095);
or U1315 (N_1315,In_1706,In_4715);
nand U1316 (N_1316,In_4866,In_4514);
xnor U1317 (N_1317,In_2298,In_2420);
or U1318 (N_1318,In_4478,In_1279);
or U1319 (N_1319,In_3394,In_2277);
and U1320 (N_1320,In_588,In_3963);
nor U1321 (N_1321,In_285,In_965);
nand U1322 (N_1322,In_3171,In_3861);
nand U1323 (N_1323,In_1522,In_1804);
and U1324 (N_1324,In_2222,In_4099);
xor U1325 (N_1325,In_1746,In_1374);
nand U1326 (N_1326,In_3586,In_3204);
or U1327 (N_1327,In_3754,In_2147);
and U1328 (N_1328,In_3561,In_1093);
and U1329 (N_1329,In_4668,In_975);
and U1330 (N_1330,In_3604,In_4216);
and U1331 (N_1331,In_2856,In_4);
and U1332 (N_1332,In_3153,In_2528);
nand U1333 (N_1333,In_1495,In_653);
nor U1334 (N_1334,In_1504,In_2429);
or U1335 (N_1335,In_977,In_2969);
xnor U1336 (N_1336,In_2631,In_3032);
xor U1337 (N_1337,In_762,In_4261);
xor U1338 (N_1338,In_1755,In_4644);
and U1339 (N_1339,In_792,In_3798);
nand U1340 (N_1340,In_344,In_3066);
nand U1341 (N_1341,In_4987,In_2747);
nand U1342 (N_1342,In_2659,In_4377);
nor U1343 (N_1343,In_3371,In_3202);
nand U1344 (N_1344,In_4319,In_4262);
nor U1345 (N_1345,In_4265,In_87);
xor U1346 (N_1346,In_2622,In_3601);
nand U1347 (N_1347,In_4224,In_4531);
nor U1348 (N_1348,In_4746,In_1684);
and U1349 (N_1349,In_4652,In_4600);
xor U1350 (N_1350,In_1121,In_1546);
xor U1351 (N_1351,In_2564,In_2502);
nor U1352 (N_1352,In_2001,In_1741);
nand U1353 (N_1353,In_3888,In_4634);
or U1354 (N_1354,In_1925,In_1635);
nor U1355 (N_1355,In_4251,In_4475);
or U1356 (N_1356,In_42,In_812);
xnor U1357 (N_1357,In_1549,In_1083);
xnor U1358 (N_1358,In_4134,In_933);
or U1359 (N_1359,In_146,In_2713);
xor U1360 (N_1360,In_3885,In_4082);
nand U1361 (N_1361,In_3932,In_1870);
or U1362 (N_1362,In_2901,In_1445);
and U1363 (N_1363,In_2110,In_2963);
or U1364 (N_1364,In_678,In_3468);
nor U1365 (N_1365,In_2263,In_1781);
or U1366 (N_1366,In_4185,In_1166);
and U1367 (N_1367,In_2764,In_3960);
nor U1368 (N_1368,In_3531,In_2875);
nand U1369 (N_1369,In_3780,In_1704);
and U1370 (N_1370,In_3157,In_372);
nor U1371 (N_1371,In_3681,In_3003);
nand U1372 (N_1372,In_3686,In_1028);
and U1373 (N_1373,In_3558,In_4398);
xor U1374 (N_1374,In_1496,In_489);
or U1375 (N_1375,In_4597,In_2774);
nor U1376 (N_1376,In_357,In_2582);
nand U1377 (N_1377,In_2894,In_2014);
nor U1378 (N_1378,In_2922,In_1105);
nor U1379 (N_1379,In_3429,In_4001);
nor U1380 (N_1380,In_682,In_2970);
nor U1381 (N_1381,In_1102,In_3753);
nor U1382 (N_1382,In_3739,In_3369);
nand U1383 (N_1383,In_3478,In_4556);
nor U1384 (N_1384,In_4334,In_4793);
nor U1385 (N_1385,In_1617,In_4166);
nand U1386 (N_1386,In_1624,In_2062);
xor U1387 (N_1387,In_2300,In_1147);
nor U1388 (N_1388,In_328,In_3222);
xnor U1389 (N_1389,In_2688,In_148);
xnor U1390 (N_1390,In_2532,In_1953);
xnor U1391 (N_1391,In_4622,In_4167);
nand U1392 (N_1392,In_1491,In_4651);
xnor U1393 (N_1393,In_1512,In_556);
nand U1394 (N_1394,In_3384,In_524);
and U1395 (N_1395,In_3160,In_3168);
and U1396 (N_1396,In_1690,In_1175);
or U1397 (N_1397,In_1096,In_4875);
nor U1398 (N_1398,In_2139,In_3461);
xnor U1399 (N_1399,In_3981,In_669);
nor U1400 (N_1400,In_1626,In_882);
or U1401 (N_1401,In_4313,In_755);
xor U1402 (N_1402,In_3640,In_1091);
or U1403 (N_1403,In_3050,In_1);
and U1404 (N_1404,In_3728,In_491);
nor U1405 (N_1405,In_10,In_3897);
nor U1406 (N_1406,In_2609,In_2261);
nand U1407 (N_1407,In_2158,In_205);
nand U1408 (N_1408,In_2935,In_178);
nor U1409 (N_1409,In_1637,In_1680);
xor U1410 (N_1410,In_59,In_4537);
or U1411 (N_1411,In_813,In_4506);
nor U1412 (N_1412,In_3812,In_941);
and U1413 (N_1413,In_3112,In_2485);
and U1414 (N_1414,In_2885,In_2859);
xor U1415 (N_1415,In_610,In_1957);
nand U1416 (N_1416,In_4149,In_2731);
nand U1417 (N_1417,In_234,In_4467);
nand U1418 (N_1418,In_4418,In_1820);
nor U1419 (N_1419,In_3397,In_1782);
and U1420 (N_1420,In_764,In_3122);
nand U1421 (N_1421,In_292,In_4072);
nor U1422 (N_1422,In_2886,In_712);
nand U1423 (N_1423,In_2205,In_3342);
and U1424 (N_1424,In_4394,In_1924);
nor U1425 (N_1425,In_583,In_2678);
and U1426 (N_1426,In_873,In_609);
xor U1427 (N_1427,In_2424,In_3645);
or U1428 (N_1428,In_3961,In_4246);
nor U1429 (N_1429,In_2781,In_2732);
xor U1430 (N_1430,In_2271,In_152);
nand U1431 (N_1431,In_4049,In_3010);
and U1432 (N_1432,In_1756,In_4969);
and U1433 (N_1433,In_2289,In_2758);
and U1434 (N_1434,In_659,In_3634);
xnor U1435 (N_1435,In_1930,In_788);
and U1436 (N_1436,In_3882,In_3715);
nor U1437 (N_1437,In_781,In_1467);
nor U1438 (N_1438,In_475,In_797);
xnor U1439 (N_1439,In_3198,In_4988);
xnor U1440 (N_1440,In_876,In_4087);
and U1441 (N_1441,In_4464,In_1533);
or U1442 (N_1442,In_4158,In_2434);
nand U1443 (N_1443,In_2208,In_2928);
xor U1444 (N_1444,In_1872,In_565);
nor U1445 (N_1445,In_654,In_919);
nand U1446 (N_1446,In_2881,In_4094);
nand U1447 (N_1447,In_4618,In_482);
nand U1448 (N_1448,In_2975,In_724);
or U1449 (N_1449,In_3658,In_4459);
or U1450 (N_1450,In_1270,In_744);
or U1451 (N_1451,In_449,In_235);
xnor U1452 (N_1452,In_4964,In_1414);
xor U1453 (N_1453,In_4487,In_1406);
nor U1454 (N_1454,In_4018,In_1448);
or U1455 (N_1455,In_1535,In_511);
and U1456 (N_1456,In_2697,In_629);
xor U1457 (N_1457,In_857,In_4069);
xor U1458 (N_1458,In_3080,In_2382);
nand U1459 (N_1459,In_2480,In_1124);
and U1460 (N_1460,In_3683,In_1029);
xnor U1461 (N_1461,In_2539,In_3975);
or U1462 (N_1462,In_392,In_1554);
nand U1463 (N_1463,In_3131,In_2265);
nand U1464 (N_1464,In_121,In_3447);
xor U1465 (N_1465,In_1878,In_994);
xor U1466 (N_1466,In_3770,In_1711);
nor U1467 (N_1467,In_3991,In_3388);
and U1468 (N_1468,In_2236,In_1987);
nor U1469 (N_1469,In_3549,In_4236);
or U1470 (N_1470,In_3306,In_3862);
and U1471 (N_1471,In_4356,In_2650);
xor U1472 (N_1472,In_71,In_4543);
or U1473 (N_1473,In_1149,In_997);
and U1474 (N_1474,In_2621,In_1722);
nor U1475 (N_1475,In_4108,In_476);
or U1476 (N_1476,In_4346,In_754);
nor U1477 (N_1477,In_4673,In_2646);
xnor U1478 (N_1478,In_1988,In_1126);
or U1479 (N_1479,In_2980,In_1962);
and U1480 (N_1480,In_4007,In_2036);
xnor U1481 (N_1481,In_3227,In_1717);
and U1482 (N_1482,In_2653,In_1158);
xor U1483 (N_1483,In_2002,In_3418);
or U1484 (N_1484,In_3771,In_2979);
xnor U1485 (N_1485,In_3274,In_4957);
xnor U1486 (N_1486,In_1936,In_379);
nand U1487 (N_1487,In_4083,In_4614);
or U1488 (N_1488,In_4209,In_1749);
xor U1489 (N_1489,In_4111,In_1514);
nor U1490 (N_1490,In_1616,In_4417);
nand U1491 (N_1491,In_2746,In_1168);
nand U1492 (N_1492,In_3038,In_4006);
or U1493 (N_1493,In_1609,In_3239);
and U1494 (N_1494,In_4162,In_3161);
nand U1495 (N_1495,In_1758,In_2206);
xor U1496 (N_1496,In_2865,In_1192);
or U1497 (N_1497,In_4878,In_3127);
and U1498 (N_1498,In_925,In_2248);
nor U1499 (N_1499,In_3207,In_420);
nor U1500 (N_1500,In_4269,In_3197);
nand U1501 (N_1501,In_3842,In_2977);
xor U1502 (N_1502,In_745,In_1463);
xor U1503 (N_1503,In_1813,In_2215);
and U1504 (N_1504,In_4826,In_2290);
xor U1505 (N_1505,In_998,In_4554);
nor U1506 (N_1506,In_4813,In_249);
or U1507 (N_1507,In_4403,In_1793);
nand U1508 (N_1508,In_4124,In_2375);
xor U1509 (N_1509,In_3976,In_2501);
xor U1510 (N_1510,In_4324,In_2051);
nor U1511 (N_1511,In_892,In_2965);
and U1512 (N_1512,In_536,In_2257);
nor U1513 (N_1513,In_3120,In_1817);
xor U1514 (N_1514,In_4724,In_3942);
nor U1515 (N_1515,In_1903,In_3826);
and U1516 (N_1516,In_4682,In_2344);
or U1517 (N_1517,In_952,In_286);
and U1518 (N_1518,In_2144,In_4551);
nand U1519 (N_1519,In_2849,In_4891);
nor U1520 (N_1520,In_2217,In_4175);
nor U1521 (N_1521,In_3266,In_726);
nand U1522 (N_1522,In_3817,In_490);
nor U1523 (N_1523,In_562,In_1906);
nor U1524 (N_1524,In_2669,In_3192);
xor U1525 (N_1525,In_2861,In_334);
or U1526 (N_1526,In_1462,In_1266);
nor U1527 (N_1527,In_2007,In_2112);
nand U1528 (N_1528,In_2985,In_2898);
nand U1529 (N_1529,In_1838,In_3599);
nor U1530 (N_1530,In_4638,In_3387);
nor U1531 (N_1531,In_2159,In_1536);
nand U1532 (N_1532,In_858,In_3378);
or U1533 (N_1533,In_2202,In_776);
nor U1534 (N_1534,In_4758,In_390);
nand U1535 (N_1535,In_670,In_4834);
and U1536 (N_1536,In_4274,In_4253);
nor U1537 (N_1537,In_4515,In_2166);
nand U1538 (N_1538,In_3712,In_1736);
and U1539 (N_1539,In_1356,In_3281);
nand U1540 (N_1540,In_4062,In_1610);
nand U1541 (N_1541,In_1328,In_1056);
nand U1542 (N_1542,In_1812,In_90);
and U1543 (N_1543,In_1865,In_3987);
nor U1544 (N_1544,In_1856,In_303);
nand U1545 (N_1545,In_3906,In_2135);
xor U1546 (N_1546,In_4694,In_2748);
or U1547 (N_1547,In_1552,In_2588);
nand U1548 (N_1548,In_4078,In_4227);
nand U1549 (N_1549,In_4510,In_1890);
xnor U1550 (N_1550,In_4050,In_4115);
or U1551 (N_1551,In_4950,In_590);
nand U1552 (N_1552,In_74,In_2464);
xnor U1553 (N_1553,In_2465,In_1036);
xor U1554 (N_1554,In_2225,In_4854);
nand U1555 (N_1555,In_2614,In_16);
or U1556 (N_1556,In_2677,In_875);
xor U1557 (N_1557,In_3996,In_4735);
nor U1558 (N_1558,In_4163,In_4198);
or U1559 (N_1559,In_1689,In_3913);
or U1560 (N_1560,In_2439,In_2636);
or U1561 (N_1561,In_1128,In_2027);
or U1562 (N_1562,In_2333,In_1629);
and U1563 (N_1563,In_2032,In_4481);
xnor U1564 (N_1564,In_2676,In_4452);
nor U1565 (N_1565,In_4143,In_3571);
xnor U1566 (N_1566,In_2356,In_3206);
xnor U1567 (N_1567,In_3538,In_1579);
nor U1568 (N_1568,In_1921,In_628);
nor U1569 (N_1569,In_3990,In_1516);
or U1570 (N_1570,In_1222,In_2234);
nor U1571 (N_1571,In_1958,In_3072);
or U1572 (N_1572,In_3143,In_2309);
and U1573 (N_1573,In_3007,In_3193);
nor U1574 (N_1574,In_4886,In_4991);
nand U1575 (N_1575,In_243,In_2282);
nor U1576 (N_1576,In_4278,In_3614);
nand U1577 (N_1577,In_1905,In_3134);
xor U1578 (N_1578,In_4410,In_1068);
nand U1579 (N_1579,In_4176,In_2906);
nand U1580 (N_1580,In_2127,In_1315);
or U1581 (N_1581,In_1857,In_4521);
and U1582 (N_1582,In_854,In_253);
or U1583 (N_1583,In_24,In_4601);
or U1584 (N_1584,In_1015,In_3617);
nand U1585 (N_1585,In_1687,In_1423);
nand U1586 (N_1586,In_2293,In_1669);
xnor U1587 (N_1587,In_2460,In_4090);
and U1588 (N_1588,In_4388,In_1164);
and U1589 (N_1589,In_3052,In_4548);
nor U1590 (N_1590,In_3595,In_13);
xnor U1591 (N_1591,In_4180,In_166);
nor U1592 (N_1592,In_2554,In_3335);
nand U1593 (N_1593,In_4486,In_2343);
and U1594 (N_1594,In_1311,In_4405);
nor U1595 (N_1595,In_2511,In_551);
and U1596 (N_1596,In_1024,In_4698);
nand U1597 (N_1597,In_3854,In_4031);
nand U1598 (N_1598,In_4360,In_1750);
nor U1599 (N_1599,In_4890,In_1140);
nand U1600 (N_1600,In_3746,In_1345);
nand U1601 (N_1601,In_2913,In_4908);
nand U1602 (N_1602,In_1537,In_3879);
nor U1603 (N_1603,In_1353,In_4226);
nor U1604 (N_1604,In_4779,In_214);
and U1605 (N_1605,In_2952,In_2360);
or U1606 (N_1606,In_2753,In_192);
xor U1607 (N_1607,In_3001,In_395);
nand U1608 (N_1608,In_3821,In_1695);
or U1609 (N_1609,In_4770,In_883);
nand U1610 (N_1610,In_181,In_1923);
xor U1611 (N_1611,In_905,In_2686);
xor U1612 (N_1612,In_2136,In_3722);
nor U1613 (N_1613,In_4282,In_506);
xor U1614 (N_1614,In_664,In_4692);
xor U1615 (N_1615,In_4920,In_563);
and U1616 (N_1616,In_1771,In_4769);
and U1617 (N_1617,In_3006,In_2620);
nand U1618 (N_1618,In_1305,In_1097);
and U1619 (N_1619,In_3711,In_1848);
and U1620 (N_1620,In_466,In_4953);
nand U1621 (N_1621,In_3948,In_4047);
nor U1622 (N_1622,In_83,In_4468);
xor U1623 (N_1623,In_3344,In_3405);
or U1624 (N_1624,In_4696,In_396);
or U1625 (N_1625,In_3923,In_1422);
xnor U1626 (N_1626,In_4238,In_4222);
xnor U1627 (N_1627,In_1373,In_4045);
nor U1628 (N_1628,In_3174,In_3501);
nor U1629 (N_1629,In_3237,In_1194);
nand U1630 (N_1630,In_3773,In_2705);
or U1631 (N_1631,In_1583,In_4676);
or U1632 (N_1632,In_3689,In_402);
nor U1633 (N_1633,In_4683,In_3151);
nor U1634 (N_1634,In_3005,In_3742);
nand U1635 (N_1635,In_3248,In_418);
and U1636 (N_1636,In_2844,In_1553);
and U1637 (N_1637,In_4962,In_915);
xor U1638 (N_1638,In_116,In_3668);
nand U1639 (N_1639,In_3566,In_1867);
or U1640 (N_1640,In_4333,In_1798);
or U1641 (N_1641,In_4546,In_2625);
xor U1642 (N_1642,In_3630,In_3296);
nor U1643 (N_1643,In_488,In_199);
nor U1644 (N_1644,In_1828,In_3146);
nor U1645 (N_1645,In_3611,In_1564);
nand U1646 (N_1646,In_1502,In_926);
nor U1647 (N_1647,In_4809,In_2851);
nand U1648 (N_1648,In_1089,In_3616);
nor U1649 (N_1649,In_534,In_2075);
nand U1650 (N_1650,In_4818,In_4938);
nand U1651 (N_1651,In_3834,In_1063);
nor U1652 (N_1652,In_4982,In_1565);
or U1653 (N_1653,In_631,In_238);
nor U1654 (N_1654,In_4662,In_1041);
nand U1655 (N_1655,In_550,In_1120);
xor U1656 (N_1656,In_2294,In_2370);
nand U1657 (N_1657,In_1954,In_2137);
nand U1658 (N_1658,In_910,In_3633);
nand U1659 (N_1659,In_2495,In_3827);
nor U1660 (N_1660,In_3103,In_4585);
nor U1661 (N_1661,In_6,In_68);
and U1662 (N_1662,In_4952,In_1231);
xnor U1663 (N_1663,In_252,In_3465);
or U1664 (N_1664,In_3225,In_2281);
or U1665 (N_1665,In_1452,In_3027);
xor U1666 (N_1666,In_92,In_1743);
nor U1667 (N_1667,In_651,In_823);
nand U1668 (N_1668,In_2418,In_2751);
nand U1669 (N_1669,In_4580,In_1400);
or U1670 (N_1670,In_2270,In_3935);
and U1671 (N_1671,In_4471,In_2791);
or U1672 (N_1672,In_4603,In_825);
or U1673 (N_1673,In_2938,In_450);
xor U1674 (N_1674,In_1751,In_2316);
nor U1675 (N_1675,In_3944,In_3627);
nand U1676 (N_1676,In_2259,In_579);
nand U1677 (N_1677,In_592,In_4970);
nand U1678 (N_1678,In_1046,In_2672);
nand U1679 (N_1679,In_1545,In_3814);
and U1680 (N_1680,In_3653,In_2169);
or U1681 (N_1681,In_1087,In_3550);
and U1682 (N_1682,In_4174,In_749);
and U1683 (N_1683,In_1402,In_836);
or U1684 (N_1684,In_948,In_613);
nor U1685 (N_1685,In_1191,In_777);
nand U1686 (N_1686,In_1208,In_3959);
or U1687 (N_1687,In_3082,In_49);
nand U1688 (N_1688,In_3487,In_4861);
and U1689 (N_1689,In_3802,In_3334);
nand U1690 (N_1690,In_3853,In_1982);
and U1691 (N_1691,In_1188,In_4430);
nand U1692 (N_1692,In_3284,In_2804);
nor U1693 (N_1693,In_1729,In_717);
or U1694 (N_1694,In_498,In_3622);
nor U1695 (N_1695,In_510,In_3835);
nand U1696 (N_1696,In_3918,In_1020);
nand U1697 (N_1697,In_3920,In_4250);
or U1698 (N_1698,In_3904,In_296);
or U1699 (N_1699,In_4727,In_1301);
nand U1700 (N_1700,In_810,In_4023);
xnor U1701 (N_1701,In_1110,In_4093);
and U1702 (N_1702,In_3585,In_4931);
or U1703 (N_1703,In_4503,In_3529);
nor U1704 (N_1704,In_3869,In_2408);
nor U1705 (N_1705,In_1582,In_1223);
and U1706 (N_1706,In_2597,In_3760);
or U1707 (N_1707,In_1308,In_3218);
nand U1708 (N_1708,In_555,In_1247);
nand U1709 (N_1709,In_995,In_1359);
nand U1710 (N_1710,In_3934,In_4894);
and U1711 (N_1711,In_3621,In_4266);
nand U1712 (N_1712,In_3692,In_1310);
or U1713 (N_1713,In_407,In_4587);
xnor U1714 (N_1714,In_3849,In_3012);
or U1715 (N_1715,In_2839,In_3214);
nand U1716 (N_1716,In_462,In_4816);
and U1717 (N_1717,In_3631,In_4883);
nand U1718 (N_1718,In_2589,In_1738);
and U1719 (N_1719,In_239,In_2474);
and U1720 (N_1720,In_283,In_2978);
or U1721 (N_1721,In_647,In_173);
and U1722 (N_1722,In_2499,In_4747);
xnor U1723 (N_1723,In_2191,In_2715);
and U1724 (N_1724,In_2146,In_2084);
xor U1725 (N_1725,In_3488,In_2991);
nor U1726 (N_1726,In_3101,In_3855);
or U1727 (N_1727,In_681,In_3114);
and U1728 (N_1728,In_2105,In_2229);
or U1729 (N_1729,In_4965,In_4871);
or U1730 (N_1730,In_3232,In_2494);
nor U1731 (N_1731,In_1256,In_3608);
or U1732 (N_1732,In_4171,In_2185);
xor U1733 (N_1733,In_2152,In_3945);
and U1734 (N_1734,In_460,In_1973);
and U1735 (N_1735,In_2188,In_2869);
or U1736 (N_1736,In_4179,In_1447);
and U1737 (N_1737,In_110,In_11);
nand U1738 (N_1738,In_679,In_471);
nand U1739 (N_1739,In_1446,In_2479);
nand U1740 (N_1740,In_2568,In_4397);
and U1741 (N_1741,In_4577,In_815);
or U1742 (N_1742,In_4370,In_4723);
or U1743 (N_1743,In_3729,In_4095);
nand U1744 (N_1744,In_4138,In_1039);
and U1745 (N_1745,In_1444,In_3140);
and U1746 (N_1746,In_2903,In_1802);
and U1747 (N_1747,In_3560,In_3891);
nor U1748 (N_1748,In_2310,In_3581);
or U1749 (N_1749,In_2843,In_1660);
xor U1750 (N_1750,In_2286,In_3380);
and U1751 (N_1751,In_2396,In_900);
nand U1752 (N_1752,In_3606,In_2302);
nand U1753 (N_1753,In_2790,In_2187);
nor U1754 (N_1754,In_699,In_3390);
nor U1755 (N_1755,In_352,In_1419);
xor U1756 (N_1756,In_3026,In_4998);
or U1757 (N_1757,In_4630,In_4159);
nor U1758 (N_1758,In_1214,In_2305);
nor U1759 (N_1759,In_1606,In_1341);
and U1760 (N_1760,In_4302,In_4722);
xnor U1761 (N_1761,In_1841,In_3736);
or U1762 (N_1762,In_1731,In_3389);
xor U1763 (N_1763,In_1117,In_3766);
nor U1764 (N_1764,In_4211,In_4084);
or U1765 (N_1765,In_2311,In_2324);
xor U1766 (N_1766,In_4232,In_868);
and U1767 (N_1767,In_774,In_1561);
xor U1768 (N_1768,In_3180,In_2182);
and U1769 (N_1769,In_2584,In_3472);
xnor U1770 (N_1770,In_1066,In_3221);
xor U1771 (N_1771,In_172,In_4881);
nor U1772 (N_1772,In_2016,In_3267);
nand U1773 (N_1773,In_108,In_587);
nand U1774 (N_1774,In_4292,In_1998);
and U1775 (N_1775,In_3937,In_3118);
or U1776 (N_1776,In_3381,In_1429);
nand U1777 (N_1777,In_3362,In_2053);
nand U1778 (N_1778,In_223,In_772);
and U1779 (N_1779,In_1713,In_805);
nor U1780 (N_1780,In_3564,In_4691);
and U1781 (N_1781,In_4195,In_2523);
xor U1782 (N_1782,In_2250,In_4135);
nand U1783 (N_1783,In_4806,In_2541);
nor U1784 (N_1784,In_4098,In_3343);
nand U1785 (N_1785,In_4845,In_4358);
xnor U1786 (N_1786,In_4207,In_3183);
nand U1787 (N_1787,In_2830,In_3439);
xor U1788 (N_1788,In_1827,In_4375);
nand U1789 (N_1789,In_2957,In_1074);
nor U1790 (N_1790,In_4172,In_2848);
nor U1791 (N_1791,In_2664,In_1540);
nor U1792 (N_1792,In_1544,In_4615);
or U1793 (N_1793,In_4629,In_721);
or U1794 (N_1794,In_2040,In_1648);
nand U1795 (N_1795,In_3555,In_124);
xnor U1796 (N_1796,In_3333,In_2930);
or U1797 (N_1797,In_3887,In_300);
nand U1798 (N_1798,In_4070,In_1895);
or U1799 (N_1799,In_889,In_2592);
and U1800 (N_1800,In_1421,In_2058);
xor U1801 (N_1801,In_77,In_1142);
nand U1802 (N_1802,In_3059,In_1006);
nand U1803 (N_1803,In_4940,In_487);
xor U1804 (N_1804,In_2942,In_1675);
xnor U1805 (N_1805,In_2717,In_263);
nor U1806 (N_1806,In_1182,In_1897);
or U1807 (N_1807,In_2510,In_4243);
nor U1808 (N_1808,In_2759,In_2724);
and U1809 (N_1809,In_1823,In_3409);
nor U1810 (N_1810,In_2211,In_3979);
nor U1811 (N_1811,In_1428,In_4425);
or U1812 (N_1812,In_4583,In_4110);
nand U1813 (N_1813,In_2142,In_3449);
nor U1814 (N_1814,In_913,In_3829);
nor U1815 (N_1815,In_3257,In_3036);
xnor U1816 (N_1816,In_70,In_2010);
nor U1817 (N_1817,In_4888,In_2776);
and U1818 (N_1818,In_1286,In_2003);
nand U1819 (N_1819,In_2726,In_501);
and U1820 (N_1820,In_4689,In_2258);
or U1821 (N_1821,In_4547,In_4961);
nor U1822 (N_1822,In_989,In_65);
nor U1823 (N_1823,In_4901,In_2168);
nor U1824 (N_1824,In_113,In_3353);
nor U1825 (N_1825,In_324,In_850);
nor U1826 (N_1826,In_3189,In_1981);
nand U1827 (N_1827,In_3326,In_1613);
and U1828 (N_1828,In_786,In_2521);
nor U1829 (N_1829,In_2312,In_137);
or U1830 (N_1830,In_461,In_723);
nor U1831 (N_1831,In_2163,In_2617);
nand U1832 (N_1832,In_1099,In_3019);
and U1833 (N_1833,In_1538,In_150);
and U1834 (N_1834,In_1989,In_1517);
and U1835 (N_1835,In_503,In_4906);
nor U1836 (N_1836,In_2559,In_4054);
nand U1837 (N_1837,In_272,In_3415);
or U1838 (N_1838,In_853,In_3761);
nand U1839 (N_1839,In_4312,In_4109);
nand U1840 (N_1840,In_2253,In_2522);
nor U1841 (N_1841,In_4041,In_375);
xnor U1842 (N_1842,In_4376,In_2227);
xnor U1843 (N_1843,In_1809,In_1507);
or U1844 (N_1844,In_3752,In_4362);
nand U1845 (N_1845,In_1550,In_4774);
and U1846 (N_1846,In_1118,In_100);
xor U1847 (N_1847,In_867,In_3519);
or U1848 (N_1848,In_184,In_4846);
or U1849 (N_1849,In_603,In_1941);
xor U1850 (N_1850,In_2180,In_1179);
nor U1851 (N_1851,In_308,In_1202);
nor U1852 (N_1852,In_3064,In_3425);
nor U1853 (N_1853,In_4034,In_3806);
or U1854 (N_1854,In_782,In_134);
xor U1855 (N_1855,In_3881,In_2548);
or U1856 (N_1856,In_1012,In_1084);
and U1857 (N_1857,In_1788,In_2958);
xor U1858 (N_1858,In_3125,In_325);
xnor U1859 (N_1859,In_739,In_1432);
and U1860 (N_1860,In_2315,In_2054);
or U1861 (N_1861,In_1594,In_2955);
xor U1862 (N_1862,In_2683,In_2933);
or U1863 (N_1863,In_57,In_4300);
and U1864 (N_1864,In_2658,In_2907);
or U1865 (N_1865,In_2029,In_1004);
nand U1866 (N_1866,In_2766,In_1395);
and U1867 (N_1867,In_4186,In_207);
xnor U1868 (N_1868,In_2536,In_1509);
nor U1869 (N_1869,In_3117,In_840);
nand U1870 (N_1870,In_2438,In_1380);
xnor U1871 (N_1871,In_1469,In_2695);
nand U1872 (N_1872,In_2644,In_2317);
nor U1873 (N_1873,In_4914,In_1451);
or U1874 (N_1874,In_1277,In_1178);
nor U1875 (N_1875,In_3108,In_1274);
and U1876 (N_1876,In_4670,In_643);
and U1877 (N_1877,In_1677,In_237);
and U1878 (N_1878,In_1170,In_1453);
and U1879 (N_1879,In_1762,In_1314);
or U1880 (N_1880,In_3941,In_1949);
and U1881 (N_1881,In_4237,In_517);
and U1882 (N_1882,In_2585,In_3972);
and U1883 (N_1883,In_1148,In_2140);
nand U1884 (N_1884,In_3525,In_992);
xor U1885 (N_1885,In_1159,In_2242);
or U1886 (N_1886,In_1940,In_1368);
nand U1887 (N_1887,In_1663,In_1061);
or U1888 (N_1888,In_4836,In_1524);
or U1889 (N_1889,In_2918,In_4808);
nor U1890 (N_1890,In_43,In_3703);
nand U1891 (N_1891,In_4702,In_3104);
or U1892 (N_1892,In_518,In_2297);
xnor U1893 (N_1893,In_2069,In_3194);
nor U1894 (N_1894,In_1768,In_364);
xnor U1895 (N_1895,In_1712,In_3516);
nand U1896 (N_1896,In_4212,In_4734);
xnor U1897 (N_1897,In_1354,In_4454);
nor U1898 (N_1898,In_3830,In_3639);
xor U1899 (N_1899,In_508,In_1671);
or U1900 (N_1900,In_1485,In_3697);
or U1901 (N_1901,In_1640,In_3800);
xor U1902 (N_1902,In_3642,In_2500);
nand U1903 (N_1903,In_2605,In_1088);
nor U1904 (N_1904,In_533,In_2812);
nand U1905 (N_1905,In_4842,In_4659);
or U1906 (N_1906,In_4633,In_1209);
or U1907 (N_1907,In_537,In_527);
and U1908 (N_1908,In_3938,In_2109);
nand U1909 (N_1909,In_817,In_2949);
nand U1910 (N_1910,In_3540,In_2481);
nor U1911 (N_1911,In_2671,In_1434);
xnor U1912 (N_1912,In_3419,In_3231);
nor U1913 (N_1913,In_1734,In_818);
nor U1914 (N_1914,In_2255,In_4709);
nor U1915 (N_1915,In_4254,In_4994);
or U1916 (N_1916,In_3873,In_4621);
nor U1917 (N_1917,In_656,In_4309);
or U1918 (N_1918,In_2860,In_3446);
nand U1919 (N_1919,In_2303,In_14);
and U1920 (N_1920,In_2956,In_3084);
nor U1921 (N_1921,In_3985,In_2915);
or U1922 (N_1922,In_3199,In_3191);
or U1923 (N_1923,In_2824,In_265);
xor U1924 (N_1924,In_2019,In_1227);
xor U1925 (N_1925,In_4392,In_1248);
and U1926 (N_1926,In_4905,In_3391);
xor U1927 (N_1927,In_3699,In_931);
nand U1928 (N_1928,In_4650,In_4593);
nor U1929 (N_1929,In_2821,In_4380);
and U1930 (N_1930,In_1952,In_329);
or U1931 (N_1931,In_729,In_3693);
and U1932 (N_1932,In_4048,In_2736);
xnor U1933 (N_1933,In_546,In_808);
and U1934 (N_1934,In_4654,In_2829);
or U1935 (N_1935,In_3876,In_4760);
or U1936 (N_1936,In_3278,In_4512);
and U1937 (N_1937,In_3043,In_63);
xor U1938 (N_1938,In_437,In_307);
nand U1939 (N_1939,In_4862,In_2953);
nor U1940 (N_1940,In_1688,In_4663);
xnor U1941 (N_1941,In_1926,In_4178);
and U1942 (N_1942,In_2301,In_2488);
and U1943 (N_1943,In_2177,In_1842);
xnor U1944 (N_1944,In_4147,In_2288);
nand U1945 (N_1945,In_1064,In_2421);
nand U1946 (N_1946,In_120,In_3073);
nor U1947 (N_1947,In_3583,In_834);
nor U1948 (N_1948,In_2021,In_3014);
or U1949 (N_1949,In_1557,In_979);
and U1950 (N_1950,In_2030,In_3675);
nand U1951 (N_1951,In_3089,In_3393);
xnor U1952 (N_1952,In_2426,In_2068);
nand U1953 (N_1953,In_2455,In_648);
nor U1954 (N_1954,In_3772,In_2186);
nand U1955 (N_1955,In_3679,In_4220);
and U1956 (N_1956,In_860,In_521);
or U1957 (N_1957,In_2011,In_354);
xnor U1958 (N_1958,In_3021,In_1519);
or U1959 (N_1959,In_0,In_966);
xnor U1960 (N_1960,In_2627,In_28);
xor U1961 (N_1961,In_2275,In_1320);
and U1962 (N_1962,In_1898,In_607);
nand U1963 (N_1963,In_2660,In_773);
xor U1964 (N_1964,In_4986,In_863);
nand U1965 (N_1965,In_2192,In_1753);
and U1966 (N_1966,In_1319,In_4275);
or U1967 (N_1967,In_3423,In_568);
nand U1968 (N_1968,In_2921,In_246);
and U1969 (N_1969,In_2862,In_2883);
and U1970 (N_1970,In_3741,In_480);
nand U1971 (N_1971,In_1636,In_1975);
or U1972 (N_1972,In_3321,In_1927);
xnor U1973 (N_1973,In_343,In_839);
nor U1974 (N_1974,In_4642,In_2161);
nand U1975 (N_1975,In_27,In_1185);
nor U1976 (N_1976,In_430,In_1860);
xnor U1977 (N_1977,In_4616,In_1288);
nand U1978 (N_1978,In_4015,In_715);
nand U1979 (N_1979,In_1347,In_144);
nand U1980 (N_1980,In_2811,In_4841);
nand U1981 (N_1981,In_939,In_566);
and U1982 (N_1982,In_665,In_188);
xnor U1983 (N_1983,In_3828,In_1604);
and U1984 (N_1984,In_4301,In_641);
xnor U1985 (N_1985,In_3398,In_4097);
xnor U1986 (N_1986,In_1503,In_151);
and U1987 (N_1987,In_4956,In_2476);
nand U1988 (N_1988,In_2452,In_2394);
nor U1989 (N_1989,In_3463,In_3382);
nand U1990 (N_1990,In_3092,In_759);
xor U1991 (N_1991,In_502,In_940);
xnor U1992 (N_1992,In_4051,In_2223);
nand U1993 (N_1993,In_4469,In_543);
nand U1994 (N_1994,In_4995,In_2045);
or U1995 (N_1995,In_2506,In_1873);
xor U1996 (N_1996,In_1937,In_2999);
xor U1997 (N_1997,In_4338,In_1670);
xnor U1998 (N_1998,In_2518,In_4932);
nand U1999 (N_1999,In_3130,In_1420);
xor U2000 (N_2000,In_1044,In_4766);
or U2001 (N_2001,In_2308,In_2721);
nor U2002 (N_2002,In_4572,In_2693);
or U2003 (N_2003,In_3847,In_4928);
nand U2004 (N_2004,In_1523,In_4457);
nor U2005 (N_2005,In_799,In_4560);
and U2006 (N_2006,In_2114,In_1425);
and U2007 (N_2007,In_763,In_3272);
xor U2008 (N_2008,In_2941,In_3416);
xor U2009 (N_2009,In_4484,In_4872);
or U2010 (N_2010,In_2430,In_4406);
xor U2011 (N_2011,In_3546,In_4068);
xor U2012 (N_2012,In_3846,In_3946);
xnor U2013 (N_2013,In_1205,In_649);
nand U2014 (N_2014,In_1430,In_45);
xnor U2015 (N_2015,In_3544,In_3119);
nand U2016 (N_2016,In_4922,In_275);
nand U2017 (N_2017,In_3044,In_208);
xor U2018 (N_2018,In_2039,In_1529);
xor U2019 (N_2019,In_3141,In_1090);
and U2020 (N_2020,In_4026,In_947);
nor U2021 (N_2021,In_2037,In_3457);
xnor U2022 (N_2022,In_514,In_3717);
or U2023 (N_2023,In_1322,In_1959);
nand U2024 (N_2024,In_3919,In_1408);
nor U2025 (N_2025,In_4354,In_79);
nand U2026 (N_2026,In_3663,In_3037);
and U2027 (N_2027,In_4337,In_4268);
nor U2028 (N_2028,In_3910,In_4387);
xor U2029 (N_2029,In_1499,In_3205);
and U2030 (N_2030,In_4416,In_803);
nand U2031 (N_2031,In_4681,In_495);
nor U2032 (N_2032,In_1007,In_1628);
xor U2033 (N_2033,In_4297,In_3458);
xnor U2034 (N_2034,In_3767,In_3190);
nor U2035 (N_2035,In_3551,In_2853);
or U2036 (N_2036,In_2497,In_3894);
and U2037 (N_2037,In_287,In_4420);
nor U2038 (N_2038,In_312,In_3040);
or U2039 (N_2039,In_3158,In_1180);
xor U2040 (N_2040,In_3152,In_4721);
and U2041 (N_2041,In_2912,In_3713);
nor U2042 (N_2042,In_3908,In_200);
nor U2043 (N_2043,In_3545,In_2657);
nor U2044 (N_2044,In_2200,In_3588);
nand U2045 (N_2045,In_2850,In_103);
nor U2046 (N_2046,In_4594,In_1379);
nor U2047 (N_2047,In_4017,In_320);
and U2048 (N_2048,In_1633,In_2503);
nor U2049 (N_2049,In_454,In_3435);
nand U2050 (N_2050,In_1505,In_2645);
xor U2051 (N_2051,In_4916,In_4655);
xnor U2052 (N_2052,In_3993,In_1302);
and U2053 (N_2053,In_4533,In_254);
nand U2054 (N_2054,In_4934,In_1466);
and U2055 (N_2055,In_741,In_1176);
xor U2056 (N_2056,In_435,In_91);
and U2057 (N_2057,In_1508,In_1350);
or U2058 (N_2058,In_3440,In_4205);
or U2059 (N_2059,In_4591,In_3971);
xor U2060 (N_2060,In_691,In_1917);
nor U2061 (N_2061,In_4326,In_2514);
xor U2062 (N_2062,In_1572,In_3467);
nand U2063 (N_2063,In_1455,In_2628);
or U2064 (N_2064,In_3726,In_4340);
or U2065 (N_2065,In_2486,In_1730);
xnor U2066 (N_2066,In_3011,In_1071);
nor U2067 (N_2067,In_1614,In_3756);
nand U2068 (N_2068,In_4825,In_4272);
and U2069 (N_2069,In_1033,In_4092);
xnor U2070 (N_2070,In_175,In_4322);
nand U2071 (N_2071,In_1101,In_637);
or U2072 (N_2072,In_760,In_1281);
and U2073 (N_2073,In_1661,In_4173);
or U2074 (N_2074,In_4756,In_1908);
and U2075 (N_2075,In_1361,In_1880);
or U2076 (N_2076,In_705,In_1810);
or U2077 (N_2077,In_710,In_2562);
or U2078 (N_2078,In_2395,In_1701);
nand U2079 (N_2079,In_3145,In_1733);
nor U2080 (N_2080,In_2358,In_2905);
xnor U2081 (N_2081,In_1627,In_497);
and U2082 (N_2082,In_662,In_3657);
xnor U2083 (N_2083,In_2092,In_1335);
and U2084 (N_2084,In_1440,In_1650);
or U2085 (N_2085,In_4647,In_2808);
or U2086 (N_2086,In_434,In_1976);
xnor U2087 (N_2087,In_1201,In_69);
nor U2088 (N_2088,In_4504,In_3408);
nor U2089 (N_2089,In_1705,In_532);
and U2090 (N_2090,In_4000,In_1212);
nor U2091 (N_2091,In_333,In_2923);
or U2092 (N_2092,In_3138,In_2757);
nor U2093 (N_2093,In_21,In_1597);
nand U2094 (N_2094,In_731,In_2123);
and U2095 (N_2095,In_618,In_2773);
xor U2096 (N_2096,In_655,In_871);
xnor U2097 (N_2097,In_97,In_3759);
or U2098 (N_2098,In_830,In_720);
nand U2099 (N_2099,In_1527,In_4838);
or U2100 (N_2100,In_3187,In_2798);
and U2101 (N_2101,In_3219,In_4329);
or U2102 (N_2102,In_2665,In_453);
or U2103 (N_2103,In_1112,In_4635);
and U2104 (N_2104,In_4835,In_1598);
and U2105 (N_2105,In_3401,In_2738);
and U2106 (N_2106,In_3704,In_4495);
or U2107 (N_2107,In_4327,In_3890);
nand U2108 (N_2108,In_3360,In_3690);
nand U2109 (N_2109,In_2138,In_576);
nand U2110 (N_2110,In_465,In_3792);
nor U2111 (N_2111,In_1674,In_224);
nand U2112 (N_2112,In_2782,In_3253);
xnor U2113 (N_2113,In_4797,In_3515);
and U2114 (N_2114,In_2797,In_2057);
or U2115 (N_2115,In_2698,In_469);
or U2116 (N_2116,In_4791,In_1608);
or U2117 (N_2117,In_180,In_1659);
and U2118 (N_2118,In_4563,In_1264);
xnor U2119 (N_2119,In_2543,In_4473);
or U2120 (N_2120,In_219,In_1862);
nand U2121 (N_2121,In_2924,In_4005);
or U2122 (N_2122,In_4540,In_2599);
and U2123 (N_2123,In_3443,In_370);
and U2124 (N_2124,In_2369,In_138);
xor U2125 (N_2125,In_4157,In_814);
nand U2126 (N_2126,In_1784,In_1103);
nor U2127 (N_2127,In_1573,In_2743);
nor U2128 (N_2128,In_1069,In_4893);
nor U2129 (N_2129,In_619,In_973);
nand U2130 (N_2130,In_2515,In_4699);
nor U2131 (N_2131,In_2332,In_4984);
nand U2132 (N_2132,In_971,In_4889);
xor U2133 (N_2133,In_4450,In_3483);
xnor U2134 (N_2134,In_4144,In_4672);
xor U2135 (N_2135,In_3203,In_1901);
xnor U2136 (N_2136,In_1581,In_2876);
nand U2137 (N_2137,In_1272,In_904);
nor U2138 (N_2138,In_1920,In_4400);
xor U2139 (N_2139,In_936,In_3212);
nor U2140 (N_2140,In_1559,In_3966);
nor U2141 (N_2141,In_4542,In_2756);
nand U2142 (N_2142,In_3536,In_3982);
nor U2143 (N_2143,In_3776,In_4693);
or U2144 (N_2144,In_2104,In_1352);
nor U2145 (N_2145,In_302,In_4837);
nor U2146 (N_2146,In_2342,In_585);
and U2147 (N_2147,In_1840,In_4780);
nor U2148 (N_2148,In_4401,In_3030);
nand U2149 (N_2149,In_668,In_2162);
and U2150 (N_2150,In_3877,In_1219);
and U2151 (N_2151,In_1593,In_2654);
nand U2152 (N_2152,In_4348,In_4775);
and U2153 (N_2153,In_557,In_512);
xnor U2154 (N_2154,In_1891,In_3147);
nand U2155 (N_2155,In_906,In_3290);
nor U2156 (N_2156,In_1916,In_2101);
and U2157 (N_2157,In_274,In_455);
nand U2158 (N_2158,In_4120,In_838);
xnor U2159 (N_2159,In_4575,In_903);
xor U2160 (N_2160,In_4096,In_3578);
xnor U2161 (N_2161,In_684,In_1607);
nor U2162 (N_2162,In_3619,In_1676);
nand U2163 (N_2163,In_4367,In_4640);
and U2164 (N_2164,In_1144,In_1801);
and U2165 (N_2165,In_3109,In_3317);
and U2166 (N_2166,In_4645,In_4279);
xor U2167 (N_2167,In_2637,In_1964);
nor U2168 (N_2168,In_4913,In_2049);
xor U2169 (N_2169,In_4765,In_2093);
xnor U2170 (N_2170,In_981,In_1555);
nor U2171 (N_2171,In_1951,In_969);
and U2172 (N_2172,In_3149,In_3831);
or U2173 (N_2173,In_3807,In_4479);
nor U2174 (N_2174,In_2517,In_974);
xor U2175 (N_2175,In_1157,In_1239);
or U2176 (N_2176,In_2459,In_2381);
and U2177 (N_2177,In_4571,In_1887);
or U2178 (N_2178,In_3428,In_2987);
nor U2179 (N_2179,In_1404,In_266);
xnor U2180 (N_2180,In_2813,In_3958);
xnor U2181 (N_2181,In_2378,In_3865);
and U2182 (N_2182,In_635,In_942);
or U2183 (N_2183,In_612,In_1025);
nand U2184 (N_2184,In_2133,In_972);
nand U2185 (N_2185,In_4520,In_326);
and U2186 (N_2186,In_2320,In_1054);
xor U2187 (N_2187,In_367,In_4415);
nand U2188 (N_2188,In_1022,In_4235);
xor U2189 (N_2189,In_1724,In_3969);
nand U2190 (N_2190,In_217,In_2224);
nand U2191 (N_2191,In_1682,In_3671);
xor U2192 (N_2192,In_2959,In_504);
and U2193 (N_2193,In_2017,In_881);
nand U2194 (N_2194,In_1971,In_459);
or U2195 (N_2195,In_1914,In_3649);
or U2196 (N_2196,In_4666,In_18);
nor U2197 (N_2197,In_2118,In_775);
or U2198 (N_2198,In_1010,In_3930);
xor U2199 (N_2199,In_19,In_3339);
xnor U2200 (N_2200,In_3034,In_1411);
and U2201 (N_2201,In_1618,In_1654);
xor U2202 (N_2202,In_2444,In_1968);
nand U2203 (N_2203,In_2702,In_4967);
and U2204 (N_2204,In_196,In_2437);
or U2205 (N_2205,In_4043,In_1686);
or U2206 (N_2206,In_2739,In_3612);
and U2207 (N_2207,In_1218,In_3107);
xnor U2208 (N_2208,In_158,In_3730);
nor U2209 (N_2209,In_3269,In_3522);
or U2210 (N_2210,In_1026,In_54);
xor U2211 (N_2211,In_4277,In_2820);
nand U2212 (N_2212,In_4993,In_1161);
nand U2213 (N_2213,In_1726,In_1603);
nor U2214 (N_2214,In_1602,In_191);
or U2215 (N_2215,In_1000,In_2616);
xnor U2216 (N_2216,In_2701,In_4902);
nor U2217 (N_2217,In_794,In_3311);
xnor U2218 (N_2218,In_1364,In_3357);
and U2219 (N_2219,In_2709,In_3648);
or U2220 (N_2220,In_3532,In_4588);
and U2221 (N_2221,In_4569,In_1778);
nand U2222 (N_2222,In_2077,In_1745);
nand U2223 (N_2223,In_4869,In_3810);
xor U2224 (N_2224,In_621,In_4384);
nand U2225 (N_2225,In_2754,In_109);
xnor U2226 (N_2226,In_2244,In_3316);
and U2227 (N_2227,In_2241,In_1806);
or U2228 (N_2228,In_4132,In_1187);
and U2229 (N_2229,In_305,In_161);
nand U2230 (N_2230,In_3115,In_3684);
or U2231 (N_2231,In_2173,In_2572);
nand U2232 (N_2232,In_1830,In_1819);
and U2233 (N_2233,In_4064,In_3909);
xnor U2234 (N_2234,In_4485,In_1822);
or U2235 (N_2235,In_1441,In_4101);
or U2236 (N_2236,In_1851,In_4331);
xor U2237 (N_2237,In_513,In_3505);
xnor U2238 (N_2238,In_907,In_2376);
and U2239 (N_2239,In_2577,In_348);
xnor U2240 (N_2240,In_56,In_3294);
xnor U2241 (N_2241,In_436,In_2059);
xnor U2242 (N_2242,In_2925,In_4568);
nor U2243 (N_2243,In_3392,In_1986);
xor U2244 (N_2244,In_2209,In_3255);
nor U2245 (N_2245,In_1651,In_4075);
nand U2246 (N_2246,In_35,In_3804);
nand U2247 (N_2247,In_2116,In_264);
or U2248 (N_2248,In_4679,In_572);
xnor U2249 (N_2249,In_806,In_2193);
nor U2250 (N_2250,In_4027,In_4470);
xor U2251 (N_2251,In_851,In_2126);
xnor U2252 (N_2252,In_2106,In_2796);
xnor U2253 (N_2253,In_2871,In_335);
nor U2254 (N_2254,In_1759,In_4002);
nor U2255 (N_2255,In_404,In_4977);
nand U2256 (N_2256,In_2610,In_4013);
xnor U2257 (N_2257,In_1137,In_1342);
or U2258 (N_2258,In_2815,In_2794);
xnor U2259 (N_2259,In_3878,In_1234);
nor U2260 (N_2260,In_2487,In_378);
xnor U2261 (N_2261,In_1130,In_3417);
nor U2262 (N_2262,In_2442,In_687);
nor U2263 (N_2263,In_4656,In_346);
nand U2264 (N_2264,In_4963,In_2467);
nor U2265 (N_2265,In_2556,In_2880);
or U2266 (N_2266,In_236,In_4359);
xnor U2267 (N_2267,In_4523,In_3768);
nand U2268 (N_2268,In_1244,In_983);
nor U2269 (N_2269,In_4657,In_1405);
or U2270 (N_2270,In_4168,In_1454);
xor U2271 (N_2271,In_2176,In_2247);
and U2272 (N_2272,In_310,In_2231);
nor U2273 (N_2273,In_4347,In_1489);
nand U2274 (N_2274,In_2042,In_677);
nand U2275 (N_2275,In_3896,In_2638);
xor U2276 (N_2276,In_2318,In_3244);
nor U2277 (N_2277,In_768,In_2763);
or U2278 (N_2278,In_2737,In_1622);
xor U2279 (N_2279,In_750,In_4700);
or U2280 (N_2280,In_1978,In_4483);
and U2281 (N_2281,In_2148,In_1075);
nor U2282 (N_2282,In_1739,In_4720);
nor U2283 (N_2283,In_693,In_531);
nand U2284 (N_2284,In_4744,In_201);
nand U2285 (N_2285,In_1883,In_1334);
nand U2286 (N_2286,In_718,In_3724);
or U2287 (N_2287,In_1053,In_3184);
xnor U2288 (N_2288,In_554,In_1942);
nand U2289 (N_2289,In_4989,In_2603);
and U2290 (N_2290,In_55,In_3875);
nor U2291 (N_2291,In_3314,In_62);
xnor U2292 (N_2292,In_3593,In_787);
or U2293 (N_2293,In_1472,In_3998);
and U2294 (N_2294,In_2022,In_2573);
nor U2295 (N_2295,In_3738,In_2249);
or U2296 (N_2296,In_3562,In_2553);
and U2297 (N_2297,In_4191,In_1343);
nand U2298 (N_2298,In_1590,In_3355);
and U2299 (N_2299,In_1045,In_2237);
xnor U2300 (N_2300,In_2216,In_2750);
nand U2301 (N_2301,In_2386,In_4314);
or U2302 (N_2302,In_3970,In_2260);
nor U2303 (N_2303,In_4511,In_2490);
nor U2304 (N_2304,In_3822,In_4273);
nor U2305 (N_2305,In_1574,In_2246);
xor U2306 (N_2306,In_4882,In_4933);
xnor U2307 (N_2307,In_1763,In_3318);
xnor U2308 (N_2308,In_4677,In_1757);
nor U2309 (N_2309,In_2566,In_4126);
nor U2310 (N_2310,In_406,In_4558);
or U2311 (N_2311,In_1918,In_2350);
and U2312 (N_2312,In_211,In_604);
nor U2313 (N_2313,In_4811,In_1913);
or U2314 (N_2314,In_67,In_1791);
or U2315 (N_2315,In_738,In_1133);
xor U2316 (N_2316,In_3530,In_548);
xor U2317 (N_2317,In_4188,In_2547);
nor U2318 (N_2318,In_3592,In_3556);
or U2319 (N_2319,In_1931,In_4378);
or U2320 (N_2320,In_3060,In_2150);
nor U2321 (N_2321,In_3866,In_1683);
nor U2322 (N_2322,In_4757,In_2251);
xor U2323 (N_2323,In_737,In_606);
and U2324 (N_2324,In_2520,In_614);
or U2325 (N_2325,In_2765,In_1769);
or U2326 (N_2326,In_2545,In_4767);
nand U2327 (N_2327,In_1866,In_1961);
nor U2328 (N_2328,In_393,In_12);
or U2329 (N_2329,In_1710,In_558);
or U2330 (N_2330,In_1275,In_1911);
xor U2331 (N_2331,In_991,In_2858);
and U2332 (N_2332,In_645,In_3526);
nand U2333 (N_2333,In_1643,In_2600);
and U2334 (N_2334,In_4802,In_4737);
and U2335 (N_2335,In_359,In_545);
or U2336 (N_2336,In_2272,In_1483);
nor U2337 (N_2337,In_2972,In_3572);
nand U2338 (N_2338,In_41,In_4177);
xnor U2339 (N_2339,In_1843,In_2550);
nor U2340 (N_2340,In_4876,In_3974);
xor U2341 (N_2341,In_4289,In_1511);
and U2342 (N_2342,In_1300,In_932);
and U2343 (N_2343,In_1351,In_3332);
nor U2344 (N_2344,In_2065,In_2818);
nor U2345 (N_2345,In_1393,In_1401);
nor U2346 (N_2346,In_416,In_888);
nor U2347 (N_2347,In_1258,In_1858);
xnor U2348 (N_2348,In_101,In_2948);
xor U2349 (N_2349,In_3524,In_4214);
or U2350 (N_2350,In_4462,In_3182);
nor U2351 (N_2351,In_3863,In_625);
or U2352 (N_2352,In_3844,In_1703);
xor U2353 (N_2353,In_2840,In_1442);
and U2354 (N_2354,In_377,In_3456);
xnor U2355 (N_2355,In_17,In_1417);
nand U2356 (N_2356,In_3249,In_2954);
nor U2357 (N_2357,In_3481,In_1030);
nor U2358 (N_2358,In_2530,In_594);
and U2359 (N_2359,In_456,In_336);
or U2360 (N_2360,In_1657,In_1038);
xor U2361 (N_2361,In_4117,In_1831);
nand U2362 (N_2362,In_2816,In_4080);
nor U2363 (N_2363,In_4675,In_611);
nor U2364 (N_2364,In_4353,In_355);
nand U2365 (N_2365,In_960,In_620);
nor U2366 (N_2366,In_3400,In_4805);
or U2367 (N_2367,In_2018,In_1899);
and U2368 (N_2368,In_2723,In_1780);
xor U2369 (N_2369,In_1928,In_675);
nor U2370 (N_2370,In_2634,In_4247);
nand U2371 (N_2371,In_3665,In_289);
nand U2372 (N_2372,In_4187,In_47);
and U2373 (N_2373,In_399,In_3867);
nand U2374 (N_2374,In_3346,In_2647);
xor U2375 (N_2375,In_2767,In_4355);
or U2376 (N_2376,In_1403,In_1337);
or U2377 (N_2377,In_3816,In_1539);
nor U2378 (N_2378,In_596,In_1797);
and U2379 (N_2379,In_3015,In_4225);
nand U2380 (N_2380,In_297,In_3785);
or U2381 (N_2381,In_4730,In_1541);
nand U2382 (N_2382,In_2130,In_3567);
xor U2383 (N_2383,In_1340,In_2685);
and U2384 (N_2384,In_105,In_827);
nand U2385 (N_2385,In_3677,In_2574);
nor U2386 (N_2386,In_2157,In_1312);
and U2387 (N_2387,In_4706,In_4972);
and U2388 (N_2388,In_3845,In_1492);
nand U2389 (N_2389,In_165,In_4393);
and U2390 (N_2390,In_4306,In_1327);
and U2391 (N_2391,In_1115,In_4123);
xor U2392 (N_2392,In_3020,In_1708);
or U2393 (N_2393,In_4189,In_824);
or U2394 (N_2394,In_1189,In_2357);
nand U2395 (N_2395,In_3629,In_4280);
nand U2396 (N_2396,In_3779,In_2561);
nor U2397 (N_2397,In_644,In_4056);
or U2398 (N_2398,In_3086,In_2789);
nand U2399 (N_2399,In_2505,In_3850);
nor U2400 (N_2400,In_4821,In_2947);
nand U2401 (N_2401,In_3801,In_322);
xnor U2402 (N_2402,In_255,In_3837);
xor U2403 (N_2403,In_2537,In_3126);
or U2404 (N_2404,In_2524,In_4731);
nand U2405 (N_2405,In_3823,In_162);
or U2406 (N_2406,In_2805,In_2393);
xnor U2407 (N_2407,In_1814,In_1230);
or U2408 (N_2408,In_1464,In_409);
nor U2409 (N_2409,In_4719,In_929);
or U2410 (N_2410,In_1720,In_564);
or U2411 (N_2411,In_1017,In_924);
nand U2412 (N_2412,In_458,In_2085);
nand U2413 (N_2413,In_1459,In_2557);
nand U2414 (N_2414,In_231,In_2785);
xnor U2415 (N_2415,In_3589,In_3077);
and U2416 (N_2416,In_4100,In_1965);
or U2417 (N_2417,In_2170,In_2422);
or U2418 (N_2418,In_1850,In_4985);
or U2419 (N_2419,In_3484,In_1893);
nor U2420 (N_2420,In_1291,In_3254);
or U2421 (N_2421,In_163,In_3539);
and U2422 (N_2422,In_3413,In_4435);
nor U2423 (N_2423,In_3163,In_894);
and U2424 (N_2424,In_3509,In_959);
xnor U2425 (N_2425,In_1847,In_1490);
nand U2426 (N_2426,In_1241,In_4941);
xnor U2427 (N_2427,In_315,In_4598);
and U2428 (N_2428,In_2771,In_1761);
nand U2429 (N_2429,In_1829,In_3029);
nand U2430 (N_2430,In_2197,In_3507);
or U2431 (N_2431,In_4071,In_376);
or U2432 (N_2432,In_3116,In_2581);
nand U2433 (N_2433,In_1240,In_674);
or U2434 (N_2434,In_1292,In_4074);
xor U2435 (N_2435,In_2552,In_2598);
nand U2436 (N_2436,In_3662,In_1970);
nor U2437 (N_2437,In_778,In_485);
xor U2438 (N_2438,In_1792,In_1948);
or U2439 (N_2439,In_956,In_221);
nand U2440 (N_2440,In_1575,In_3462);
nand U2441 (N_2441,In_4184,In_1599);
or U2442 (N_2442,In_1845,In_2870);
nor U2443 (N_2443,In_3482,In_3949);
nand U2444 (N_2444,In_251,In_4039);
and U2445 (N_2445,In_4063,In_486);
or U2446 (N_2446,In_3293,In_189);
xnor U2447 (N_2447,In_2416,In_4404);
or U2448 (N_2448,In_1630,In_3074);
or U2449 (N_2449,In_1474,In_2096);
nor U2450 (N_2450,In_164,In_4992);
and U2451 (N_2451,In_2730,In_4880);
nand U2452 (N_2452,In_2410,In_2902);
or U2453 (N_2453,In_4349,In_1094);
xor U2454 (N_2454,In_3099,In_1645);
and U2455 (N_2455,In_331,In_4350);
nor U2456 (N_2456,In_3548,In_2666);
or U2457 (N_2457,In_1642,In_1200);
or U2458 (N_2458,In_2516,In_4351);
or U2459 (N_2459,In_2966,In_3947);
nand U2460 (N_2460,In_389,In_2655);
nand U2461 (N_2461,In_1922,In_4860);
nand U2462 (N_2462,In_2828,In_2154);
xnor U2463 (N_2463,In_639,In_350);
xor U2464 (N_2464,In_3521,In_299);
or U2465 (N_2465,In_3201,In_432);
nand U2466 (N_2466,In_2457,In_23);
or U2467 (N_2467,In_1691,In_182);
xnor U2468 (N_2468,In_1481,In_3789);
xor U2469 (N_2469,In_4879,In_2578);
xnor U2470 (N_2470,In_732,In_2917);
nand U2471 (N_2471,In_1816,In_112);
or U2472 (N_2472,In_464,In_3412);
xnor U2473 (N_2473,In_4480,In_891);
nand U2474 (N_2474,In_3301,In_2546);
or U2475 (N_2475,In_2897,In_3473);
and U2476 (N_2476,In_3113,In_1050);
nor U2477 (N_2477,In_3661,In_3264);
nand U2478 (N_2478,In_3213,In_341);
and U2479 (N_2479,In_3215,In_4508);
xor U2480 (N_2480,In_2699,In_790);
and U2481 (N_2481,In_245,In_3260);
and U2482 (N_2482,In_561,In_160);
and U2483 (N_2483,In_198,In_167);
nor U2484 (N_2484,In_855,In_3520);
xor U2485 (N_2485,In_2968,In_3139);
nand U2486 (N_2486,In_2034,In_3327);
xnor U2487 (N_2487,In_4921,In_4399);
xor U2488 (N_2488,In_3025,In_2786);
and U2489 (N_2489,In_58,In_4221);
or U2490 (N_2490,In_423,In_1475);
or U2491 (N_2491,In_3148,In_4257);
nand U2492 (N_2492,In_3933,In_278);
and U2493 (N_2493,In_796,In_861);
or U2494 (N_2494,In_766,In_4140);
nand U2495 (N_2495,In_4954,In_505);
and U2496 (N_2496,In_1070,In_4330);
nand U2497 (N_2497,In_3067,In_3848);
nor U2498 (N_2498,In_2579,In_4281);
nand U2499 (N_2499,In_2908,In_4799);
or U2500 (N_2500,N_703,N_1932);
or U2501 (N_2501,N_1498,N_2111);
and U2502 (N_2502,N_881,N_1416);
nor U2503 (N_2503,N_51,N_1190);
nor U2504 (N_2504,N_181,N_1160);
and U2505 (N_2505,N_1319,N_2469);
or U2506 (N_2506,N_2259,N_906);
nand U2507 (N_2507,N_44,N_784);
and U2508 (N_2508,N_1560,N_235);
and U2509 (N_2509,N_1989,N_158);
nand U2510 (N_2510,N_736,N_615);
and U2511 (N_2511,N_2310,N_1421);
nand U2512 (N_2512,N_350,N_608);
or U2513 (N_2513,N_2209,N_543);
and U2514 (N_2514,N_53,N_1312);
xor U2515 (N_2515,N_102,N_898);
nor U2516 (N_2516,N_1629,N_456);
and U2517 (N_2517,N_336,N_1727);
nand U2518 (N_2518,N_1286,N_2322);
xnor U2519 (N_2519,N_240,N_281);
xor U2520 (N_2520,N_1834,N_1211);
xnor U2521 (N_2521,N_69,N_1783);
or U2522 (N_2522,N_1870,N_1247);
or U2523 (N_2523,N_136,N_2489);
nand U2524 (N_2524,N_513,N_1168);
or U2525 (N_2525,N_2115,N_1674);
nand U2526 (N_2526,N_399,N_512);
xnor U2527 (N_2527,N_269,N_1452);
nor U2528 (N_2528,N_2343,N_172);
and U2529 (N_2529,N_1206,N_1759);
or U2530 (N_2530,N_1990,N_1371);
nand U2531 (N_2531,N_823,N_372);
nor U2532 (N_2532,N_1760,N_54);
nand U2533 (N_2533,N_1335,N_1465);
nor U2534 (N_2534,N_259,N_893);
and U2535 (N_2535,N_483,N_190);
nand U2536 (N_2536,N_1584,N_352);
nand U2537 (N_2537,N_1254,N_790);
nor U2538 (N_2538,N_2023,N_2092);
nand U2539 (N_2539,N_708,N_1695);
xnor U2540 (N_2540,N_1679,N_1652);
nand U2541 (N_2541,N_1151,N_56);
xnor U2542 (N_2542,N_2269,N_980);
nor U2543 (N_2543,N_1896,N_266);
xnor U2544 (N_2544,N_2426,N_2316);
nor U2545 (N_2545,N_320,N_167);
and U2546 (N_2546,N_95,N_359);
and U2547 (N_2547,N_964,N_1924);
nand U2548 (N_2548,N_792,N_272);
and U2549 (N_2549,N_337,N_1737);
and U2550 (N_2550,N_2192,N_2194);
nand U2551 (N_2551,N_1696,N_2490);
or U2552 (N_2552,N_2450,N_1725);
or U2553 (N_2553,N_2327,N_2299);
xor U2554 (N_2554,N_1118,N_1669);
xor U2555 (N_2555,N_1677,N_2168);
nand U2556 (N_2556,N_1174,N_1493);
nand U2557 (N_2557,N_1950,N_2458);
nand U2558 (N_2558,N_846,N_1);
or U2559 (N_2559,N_1154,N_1340);
nor U2560 (N_2560,N_1293,N_1218);
xor U2561 (N_2561,N_2205,N_566);
nor U2562 (N_2562,N_1387,N_1810);
nor U2563 (N_2563,N_2179,N_2271);
and U2564 (N_2564,N_293,N_1794);
xnor U2565 (N_2565,N_1373,N_1266);
or U2566 (N_2566,N_1489,N_1450);
or U2567 (N_2567,N_371,N_870);
and U2568 (N_2568,N_379,N_1278);
nor U2569 (N_2569,N_1890,N_619);
and U2570 (N_2570,N_2027,N_757);
nand U2571 (N_2571,N_1137,N_1649);
xor U2572 (N_2572,N_1277,N_2370);
and U2573 (N_2573,N_1745,N_1280);
xor U2574 (N_2574,N_354,N_459);
nand U2575 (N_2575,N_1210,N_1173);
nand U2576 (N_2576,N_1288,N_1900);
xnor U2577 (N_2577,N_1958,N_341);
xnor U2578 (N_2578,N_1599,N_2474);
xor U2579 (N_2579,N_2176,N_2104);
or U2580 (N_2580,N_1527,N_90);
xor U2581 (N_2581,N_1818,N_2389);
nand U2582 (N_2582,N_2284,N_2238);
nand U2583 (N_2583,N_82,N_1388);
xor U2584 (N_2584,N_205,N_1065);
nand U2585 (N_2585,N_1214,N_1929);
nand U2586 (N_2586,N_816,N_1536);
nand U2587 (N_2587,N_1681,N_103);
nor U2588 (N_2588,N_531,N_67);
nand U2589 (N_2589,N_2409,N_2332);
and U2590 (N_2590,N_774,N_1953);
and U2591 (N_2591,N_2100,N_1079);
nor U2592 (N_2592,N_2208,N_2126);
and U2593 (N_2593,N_106,N_1558);
nor U2594 (N_2594,N_80,N_2277);
and U2595 (N_2595,N_704,N_2479);
and U2596 (N_2596,N_1399,N_1867);
xnor U2597 (N_2597,N_2180,N_671);
and U2598 (N_2598,N_73,N_1843);
and U2599 (N_2599,N_2448,N_1644);
and U2600 (N_2600,N_467,N_125);
nor U2601 (N_2601,N_722,N_1222);
xor U2602 (N_2602,N_2071,N_1094);
and U2603 (N_2603,N_1034,N_872);
xor U2604 (N_2604,N_2273,N_2199);
xnor U2605 (N_2605,N_415,N_1739);
nor U2606 (N_2606,N_177,N_1899);
xor U2607 (N_2607,N_1395,N_1336);
nand U2608 (N_2608,N_2484,N_2321);
nand U2609 (N_2609,N_1510,N_560);
or U2610 (N_2610,N_2442,N_308);
and U2611 (N_2611,N_362,N_1743);
or U2612 (N_2612,N_2401,N_922);
or U2613 (N_2613,N_409,N_1246);
xor U2614 (N_2614,N_1274,N_1878);
nand U2615 (N_2615,N_2497,N_32);
nor U2616 (N_2616,N_546,N_1345);
nor U2617 (N_2617,N_1091,N_1187);
and U2618 (N_2618,N_360,N_123);
or U2619 (N_2619,N_2043,N_681);
nand U2620 (N_2620,N_2211,N_1477);
or U2621 (N_2621,N_1839,N_1035);
or U2622 (N_2622,N_744,N_1242);
nor U2623 (N_2623,N_2283,N_31);
xnor U2624 (N_2624,N_1587,N_977);
xor U2625 (N_2625,N_2174,N_1817);
and U2626 (N_2626,N_861,N_1732);
and U2627 (N_2627,N_641,N_658);
and U2628 (N_2628,N_2364,N_215);
or U2629 (N_2629,N_2013,N_2153);
nand U2630 (N_2630,N_1949,N_2058);
nor U2631 (N_2631,N_316,N_1303);
or U2632 (N_2632,N_1790,N_28);
nand U2633 (N_2633,N_987,N_1486);
nor U2634 (N_2634,N_2415,N_941);
nor U2635 (N_2635,N_1691,N_369);
and U2636 (N_2636,N_763,N_1552);
xor U2637 (N_2637,N_765,N_50);
nor U2638 (N_2638,N_2062,N_1013);
or U2639 (N_2639,N_470,N_1012);
and U2640 (N_2640,N_1177,N_1138);
xor U2641 (N_2641,N_1447,N_322);
xor U2642 (N_2642,N_633,N_1331);
or U2643 (N_2643,N_2292,N_1961);
xor U2644 (N_2644,N_1224,N_135);
xnor U2645 (N_2645,N_755,N_2435);
nor U2646 (N_2646,N_1873,N_113);
nand U2647 (N_2647,N_304,N_1304);
and U2648 (N_2648,N_1577,N_1182);
and U2649 (N_2649,N_1827,N_789);
or U2650 (N_2650,N_2042,N_1802);
xnor U2651 (N_2651,N_1040,N_2025);
xnor U2652 (N_2652,N_2093,N_1009);
or U2653 (N_2653,N_2262,N_2320);
or U2654 (N_2654,N_1750,N_958);
and U2655 (N_2655,N_2339,N_278);
xnor U2656 (N_2656,N_2354,N_26);
nand U2657 (N_2657,N_2375,N_664);
nor U2658 (N_2658,N_217,N_343);
xnor U2659 (N_2659,N_962,N_969);
xnor U2660 (N_2660,N_2207,N_1807);
and U2661 (N_2661,N_1532,N_1162);
or U2662 (N_2662,N_2344,N_1700);
and U2663 (N_2663,N_1730,N_2463);
and U2664 (N_2664,N_234,N_1755);
nand U2665 (N_2665,N_1575,N_168);
or U2666 (N_2666,N_498,N_875);
nand U2667 (N_2667,N_1579,N_1016);
or U2668 (N_2668,N_2380,N_454);
nand U2669 (N_2669,N_1495,N_2066);
nor U2670 (N_2670,N_1578,N_497);
and U2671 (N_2671,N_524,N_2247);
nand U2672 (N_2672,N_594,N_1813);
nor U2673 (N_2673,N_140,N_769);
nor U2674 (N_2674,N_632,N_2480);
and U2675 (N_2675,N_1561,N_1947);
xnor U2676 (N_2676,N_173,N_2477);
nand U2677 (N_2677,N_2172,N_469);
nand U2678 (N_2678,N_808,N_1778);
nor U2679 (N_2679,N_2485,N_1630);
nand U2680 (N_2680,N_685,N_2053);
or U2681 (N_2681,N_1483,N_1586);
nand U2682 (N_2682,N_2252,N_1917);
or U2683 (N_2683,N_2422,N_1951);
or U2684 (N_2684,N_2297,N_1982);
or U2685 (N_2685,N_687,N_2464);
xor U2686 (N_2686,N_1986,N_2219);
and U2687 (N_2687,N_536,N_1291);
nand U2688 (N_2688,N_1604,N_2431);
nor U2689 (N_2689,N_1888,N_559);
nand U2690 (N_2690,N_1757,N_1525);
or U2691 (N_2691,N_1386,N_1339);
and U2692 (N_2692,N_591,N_299);
nand U2693 (N_2693,N_713,N_1364);
nand U2694 (N_2694,N_126,N_265);
nand U2695 (N_2695,N_1927,N_918);
nor U2696 (N_2696,N_1208,N_2487);
xnor U2697 (N_2697,N_923,N_413);
nand U2698 (N_2698,N_41,N_2196);
xnor U2699 (N_2699,N_2157,N_890);
nor U2700 (N_2700,N_212,N_2369);
nor U2701 (N_2701,N_429,N_397);
nor U2702 (N_2702,N_887,N_1686);
or U2703 (N_2703,N_307,N_2360);
and U2704 (N_2704,N_648,N_746);
and U2705 (N_2705,N_2291,N_1786);
and U2706 (N_2706,N_1670,N_2335);
nand U2707 (N_2707,N_1131,N_1188);
xnor U2708 (N_2708,N_766,N_1590);
and U2709 (N_2709,N_2051,N_2390);
xnor U2710 (N_2710,N_1542,N_768);
nand U2711 (N_2711,N_1425,N_1814);
and U2712 (N_2712,N_1112,N_2365);
and U2713 (N_2713,N_1333,N_1824);
xor U2714 (N_2714,N_1053,N_2045);
or U2715 (N_2715,N_400,N_490);
xnor U2716 (N_2716,N_1367,N_14);
and U2717 (N_2717,N_1499,N_1516);
nor U2718 (N_2718,N_282,N_1104);
nor U2719 (N_2719,N_1271,N_1944);
nand U2720 (N_2720,N_1660,N_1627);
and U2721 (N_2721,N_1444,N_2055);
and U2722 (N_2722,N_2187,N_111);
nor U2723 (N_2723,N_1613,N_824);
or U2724 (N_2724,N_907,N_572);
nor U2725 (N_2725,N_2395,N_2307);
xnor U2726 (N_2726,N_2482,N_1791);
nand U2727 (N_2727,N_771,N_2425);
or U2728 (N_2728,N_40,N_1068);
and U2729 (N_2729,N_39,N_1726);
or U2730 (N_2730,N_486,N_461);
nand U2731 (N_2731,N_2381,N_1570);
xor U2732 (N_2732,N_374,N_1565);
nand U2733 (N_2733,N_522,N_2266);
and U2734 (N_2734,N_643,N_2439);
or U2735 (N_2735,N_1683,N_568);
or U2736 (N_2736,N_1087,N_882);
nand U2737 (N_2737,N_1163,N_1909);
or U2738 (N_2738,N_1092,N_6);
and U2739 (N_2739,N_1136,N_1390);
xnor U2740 (N_2740,N_1047,N_740);
and U2741 (N_2741,N_1310,N_1368);
xnor U2742 (N_2742,N_160,N_1838);
xnor U2743 (N_2743,N_2021,N_1698);
nand U2744 (N_2744,N_787,N_1567);
and U2745 (N_2745,N_1402,N_558);
xor U2746 (N_2746,N_1712,N_2315);
nor U2747 (N_2747,N_609,N_837);
or U2748 (N_2748,N_1687,N_196);
xor U2749 (N_2749,N_208,N_2008);
xor U2750 (N_2750,N_447,N_699);
and U2751 (N_2751,N_1635,N_1752);
or U2752 (N_2752,N_1828,N_481);
nor U2753 (N_2753,N_133,N_1892);
nor U2754 (N_2754,N_1530,N_43);
nand U2755 (N_2755,N_812,N_1380);
nor U2756 (N_2756,N_2272,N_1326);
or U2757 (N_2757,N_1167,N_1435);
and U2758 (N_2758,N_59,N_251);
and U2759 (N_2759,N_1245,N_564);
and U2760 (N_2760,N_2248,N_1073);
and U2761 (N_2761,N_2044,N_263);
and U2762 (N_2762,N_1699,N_1563);
or U2763 (N_2763,N_2223,N_2186);
and U2764 (N_2764,N_1366,N_596);
nor U2765 (N_2765,N_2281,N_732);
nor U2766 (N_2766,N_1109,N_2368);
and U2767 (N_2767,N_404,N_2333);
nor U2768 (N_2768,N_383,N_2460);
nor U2769 (N_2769,N_2123,N_2190);
xor U2770 (N_2770,N_244,N_166);
xnor U2771 (N_2771,N_323,N_667);
nand U2772 (N_2772,N_1535,N_2116);
xor U2773 (N_2773,N_395,N_2138);
and U2774 (N_2774,N_2371,N_1777);
nor U2775 (N_2775,N_2363,N_433);
nor U2776 (N_2776,N_302,N_305);
xor U2777 (N_2777,N_2056,N_189);
or U2778 (N_2778,N_1826,N_1939);
or U2779 (N_2779,N_534,N_753);
nor U2780 (N_2780,N_1194,N_2420);
or U2781 (N_2781,N_1327,N_1346);
or U2782 (N_2782,N_2096,N_327);
nor U2783 (N_2783,N_1122,N_795);
and U2784 (N_2784,N_1243,N_2278);
or U2785 (N_2785,N_1815,N_22);
and U2786 (N_2786,N_2134,N_1394);
nor U2787 (N_2787,N_2083,N_1963);
nor U2788 (N_2788,N_612,N_1145);
or U2789 (N_2789,N_1157,N_661);
xor U2790 (N_2790,N_614,N_1809);
nor U2791 (N_2791,N_241,N_567);
xnor U2792 (N_2792,N_63,N_1641);
xnor U2793 (N_2793,N_605,N_822);
xnor U2794 (N_2794,N_1031,N_16);
nor U2795 (N_2795,N_578,N_1466);
or U2796 (N_2796,N_994,N_35);
nand U2797 (N_2797,N_1562,N_1805);
or U2798 (N_2798,N_2089,N_2003);
and U2799 (N_2799,N_321,N_778);
and U2800 (N_2800,N_662,N_672);
nor U2801 (N_2801,N_1370,N_130);
xnor U2802 (N_2802,N_1044,N_1847);
xor U2803 (N_2803,N_1481,N_1966);
nor U2804 (N_2804,N_2127,N_1938);
xor U2805 (N_2805,N_1764,N_132);
nand U2806 (N_2806,N_7,N_506);
nand U2807 (N_2807,N_188,N_1377);
and U2808 (N_2808,N_820,N_1615);
xnor U2809 (N_2809,N_1438,N_2000);
nand U2810 (N_2810,N_474,N_1219);
or U2811 (N_2811,N_1508,N_2032);
xor U2812 (N_2812,N_1857,N_1746);
nand U2813 (N_2813,N_1209,N_2011);
and U2814 (N_2814,N_347,N_296);
nor U2815 (N_2815,N_210,N_1866);
xor U2816 (N_2816,N_1954,N_1609);
xor U2817 (N_2817,N_720,N_2150);
nand U2818 (N_2818,N_280,N_1891);
nand U2819 (N_2819,N_2210,N_1507);
or U2820 (N_2820,N_1522,N_598);
or U2821 (N_2821,N_613,N_1580);
xnor U2822 (N_2822,N_2106,N_1269);
or U2823 (N_2823,N_1614,N_624);
xor U2824 (N_2824,N_209,N_1036);
or U2825 (N_2825,N_1987,N_0);
or U2826 (N_2826,N_1120,N_1877);
or U2827 (N_2827,N_1884,N_2145);
and U2828 (N_2828,N_892,N_1490);
and U2829 (N_2829,N_2323,N_1133);
and U2830 (N_2830,N_2230,N_2374);
xnor U2831 (N_2831,N_2455,N_1569);
nor U2832 (N_2832,N_1284,N_1063);
or U2833 (N_2833,N_220,N_1262);
xnor U2834 (N_2834,N_919,N_2471);
xnor U2835 (N_2835,N_1060,N_948);
xnor U2836 (N_2836,N_1519,N_607);
nand U2837 (N_2837,N_745,N_475);
or U2838 (N_2838,N_500,N_455);
xnor U2839 (N_2839,N_2312,N_1975);
or U2840 (N_2840,N_1868,N_1948);
xnor U2841 (N_2841,N_351,N_439);
xor U2842 (N_2842,N_864,N_192);
xnor U2843 (N_2843,N_714,N_1543);
and U2844 (N_2844,N_1874,N_584);
and U2845 (N_2845,N_1808,N_719);
nand U2846 (N_2846,N_151,N_1841);
nor U2847 (N_2847,N_2202,N_581);
and U2848 (N_2848,N_1476,N_555);
and U2849 (N_2849,N_1022,N_1716);
xor U2850 (N_2850,N_602,N_1375);
and U2851 (N_2851,N_1968,N_1411);
nand U2852 (N_2852,N_734,N_2002);
and U2853 (N_2853,N_1556,N_1229);
nor U2854 (N_2854,N_47,N_911);
nor U2855 (N_2855,N_523,N_972);
and U2856 (N_2856,N_261,N_1008);
and U2857 (N_2857,N_1583,N_1514);
xor U2858 (N_2858,N_1276,N_950);
and U2859 (N_2859,N_865,N_760);
nor U2860 (N_2860,N_457,N_1894);
or U2861 (N_2861,N_1601,N_975);
nor U2862 (N_2862,N_1741,N_1671);
xnor U2863 (N_2863,N_411,N_1066);
xnor U2864 (N_2864,N_2311,N_8);
nor U2865 (N_2865,N_1960,N_1589);
nand U2866 (N_2866,N_174,N_1473);
xor U2867 (N_2867,N_2372,N_1544);
or U2868 (N_2868,N_960,N_2414);
nand U2869 (N_2869,N_1383,N_1610);
nor U2870 (N_2870,N_1665,N_582);
or U2871 (N_2871,N_1771,N_434);
or U2872 (N_2872,N_1523,N_267);
nand U2873 (N_2873,N_2031,N_34);
or U2874 (N_2874,N_1415,N_2366);
xor U2875 (N_2875,N_2005,N_2214);
or U2876 (N_2876,N_1249,N_274);
or U2877 (N_2877,N_1343,N_491);
or U2878 (N_2878,N_1574,N_1959);
or U2879 (N_2879,N_2175,N_1062);
or U2880 (N_2880,N_107,N_696);
or U2881 (N_2881,N_737,N_819);
or U2882 (N_2882,N_2195,N_1547);
nor U2883 (N_2883,N_845,N_554);
or U2884 (N_2884,N_1401,N_81);
xnor U2885 (N_2885,N_742,N_1619);
and U2886 (N_2886,N_1238,N_1082);
nand U2887 (N_2887,N_2029,N_2398);
nand U2888 (N_2888,N_2308,N_2394);
xnor U2889 (N_2889,N_1125,N_1648);
nand U2890 (N_2890,N_157,N_981);
nand U2891 (N_2891,N_1518,N_2275);
and U2892 (N_2892,N_175,N_695);
nor U2893 (N_2893,N_65,N_2251);
or U2894 (N_2894,N_2224,N_599);
xnor U2895 (N_2895,N_940,N_1645);
nor U2896 (N_2896,N_938,N_2416);
and U2897 (N_2897,N_1069,N_23);
nand U2898 (N_2898,N_1296,N_2107);
nor U2899 (N_2899,N_2001,N_2249);
nor U2900 (N_2900,N_1926,N_840);
and U2901 (N_2901,N_473,N_2267);
nand U2902 (N_2902,N_1230,N_1637);
nor U2903 (N_2903,N_1223,N_724);
nand U2904 (N_2904,N_1734,N_248);
xnor U2905 (N_2905,N_488,N_2094);
nand U2906 (N_2906,N_92,N_60);
and U2907 (N_2907,N_1862,N_426);
and U2908 (N_2908,N_1484,N_435);
and U2909 (N_2909,N_2197,N_1124);
nor U2910 (N_2910,N_674,N_2433);
nor U2911 (N_2911,N_2102,N_1148);
xor U2912 (N_2912,N_1311,N_423);
and U2913 (N_2913,N_673,N_381);
nor U2914 (N_2914,N_651,N_636);
nor U2915 (N_2915,N_294,N_1429);
and U2916 (N_2916,N_1275,N_2276);
and U2917 (N_2917,N_348,N_78);
or U2918 (N_2918,N_1299,N_143);
nor U2919 (N_2919,N_1605,N_12);
or U2920 (N_2920,N_2105,N_339);
nor U2921 (N_2921,N_2258,N_1001);
xnor U2922 (N_2922,N_541,N_2498);
nor U2923 (N_2923,N_509,N_1289);
or U2924 (N_2924,N_2155,N_2265);
or U2925 (N_2925,N_1056,N_751);
and U2926 (N_2926,N_219,N_1844);
nor U2927 (N_2927,N_1566,N_1650);
and U2928 (N_2928,N_1309,N_1226);
nand U2929 (N_2929,N_2,N_639);
nor U2930 (N_2930,N_759,N_1272);
xor U2931 (N_2931,N_1397,N_1029);
nor U2932 (N_2932,N_677,N_630);
or U2933 (N_2933,N_33,N_2350);
and U2934 (N_2934,N_2376,N_1685);
and U2935 (N_2935,N_226,N_1135);
or U2936 (N_2936,N_688,N_528);
nor U2937 (N_2937,N_2074,N_206);
xor U2938 (N_2938,N_529,N_585);
or U2939 (N_2939,N_540,N_225);
and U2940 (N_2940,N_1071,N_2481);
or U2941 (N_2941,N_216,N_1225);
nand U2942 (N_2942,N_507,N_398);
xnor U2943 (N_2943,N_1318,N_468);
nand U2944 (N_2944,N_119,N_638);
nor U2945 (N_2945,N_1903,N_1203);
or U2946 (N_2946,N_1895,N_1512);
nor U2947 (N_2947,N_122,N_204);
nand U2948 (N_2948,N_754,N_1026);
nor U2949 (N_2949,N_1179,N_1883);
or U2950 (N_2950,N_1515,N_179);
xnor U2951 (N_2951,N_460,N_995);
xor U2952 (N_2952,N_711,N_1461);
and U2953 (N_2953,N_831,N_653);
nand U2954 (N_2954,N_373,N_869);
xor U2955 (N_2955,N_752,N_1634);
nand U2956 (N_2956,N_668,N_2411);
and U2957 (N_2957,N_1920,N_463);
xnor U2958 (N_2958,N_905,N_1740);
nor U2959 (N_2959,N_561,N_1680);
nor U2960 (N_2960,N_1253,N_929);
or U2961 (N_2961,N_164,N_1405);
nor U2962 (N_2962,N_2392,N_1200);
nor U2963 (N_2963,N_691,N_1553);
or U2964 (N_2964,N_1462,N_1240);
nand U2965 (N_2965,N_2462,N_178);
nor U2966 (N_2966,N_1820,N_1096);
nand U2967 (N_2967,N_593,N_728);
and U2968 (N_2968,N_1212,N_1172);
nand U2969 (N_2969,N_17,N_1772);
nand U2970 (N_2970,N_569,N_2438);
xor U2971 (N_2971,N_1885,N_1804);
and U2972 (N_2972,N_2038,N_169);
nor U2973 (N_2973,N_389,N_2154);
nor U2974 (N_2974,N_2399,N_2110);
nand U2975 (N_2975,N_1028,N_2143);
or U2976 (N_2976,N_727,N_1362);
or U2977 (N_2977,N_1090,N_1201);
xnor U2978 (N_2978,N_1485,N_1640);
and U2979 (N_2979,N_762,N_1910);
or U2980 (N_2980,N_1761,N_1784);
xnor U2981 (N_2981,N_1612,N_466);
nand U2982 (N_2982,N_334,N_1851);
nor U2983 (N_2983,N_1546,N_254);
nand U2984 (N_2984,N_580,N_973);
nor U2985 (N_2985,N_2324,N_1831);
or U2986 (N_2986,N_2129,N_689);
xor U2987 (N_2987,N_328,N_1250);
nor U2988 (N_2988,N_1502,N_515);
xnor U2989 (N_2989,N_1100,N_2086);
or U2990 (N_2990,N_1598,N_338);
nand U2991 (N_2991,N_2080,N_2421);
and U2992 (N_2992,N_603,N_1500);
nor U2993 (N_2993,N_640,N_252);
nor U2994 (N_2994,N_2383,N_1541);
and U2995 (N_2995,N_68,N_1350);
or U2996 (N_2996,N_967,N_156);
nand U2997 (N_2997,N_2181,N_1018);
nor U2998 (N_2998,N_1014,N_1710);
nor U2999 (N_2999,N_618,N_2470);
and U3000 (N_3000,N_2405,N_1651);
nor U3001 (N_3001,N_2402,N_1393);
nand U3002 (N_3002,N_2212,N_1875);
nor U3003 (N_3003,N_108,N_717);
and U3004 (N_3004,N_1775,N_1093);
nor U3005 (N_3005,N_1113,N_642);
xnor U3006 (N_3006,N_849,N_200);
and U3007 (N_3007,N_1297,N_1381);
and U3008 (N_3008,N_1349,N_2408);
or U3009 (N_3009,N_2136,N_419);
or U3010 (N_3010,N_2028,N_535);
nor U3011 (N_3011,N_64,N_1835);
or U3012 (N_3012,N_325,N_935);
or U3013 (N_3013,N_257,N_2254);
and U3014 (N_3014,N_828,N_1863);
nor U3015 (N_3015,N_1357,N_303);
nand U3016 (N_3016,N_74,N_1192);
or U3017 (N_3017,N_516,N_1731);
or U3018 (N_3018,N_2353,N_2077);
nand U3019 (N_3019,N_2349,N_2280);
nor U3020 (N_3020,N_1689,N_2120);
nand U3021 (N_3021,N_723,N_418);
and U3022 (N_3022,N_1440,N_983);
or U3023 (N_3023,N_1636,N_2237);
nor U3024 (N_3024,N_197,N_1642);
nor U3025 (N_3025,N_2076,N_27);
and U3026 (N_3026,N_853,N_796);
nor U3027 (N_3027,N_444,N_1032);
and U3028 (N_3028,N_2033,N_1769);
nor U3029 (N_3029,N_2290,N_1721);
nand U3030 (N_3030,N_145,N_1736);
xnor U3031 (N_3031,N_1454,N_1302);
xor U3032 (N_3032,N_1528,N_625);
nand U3033 (N_3033,N_57,N_1703);
and U3034 (N_3034,N_465,N_377);
nand U3035 (N_3035,N_914,N_2139);
nand U3036 (N_3036,N_2114,N_1618);
xnor U3037 (N_3037,N_1889,N_1153);
and U3038 (N_3038,N_2457,N_79);
and U3039 (N_3039,N_1017,N_937);
nand U3040 (N_3040,N_521,N_1942);
xnor U3041 (N_3041,N_503,N_2418);
xor U3042 (N_3042,N_1389,N_2377);
xor U3043 (N_3043,N_2164,N_984);
xnor U3044 (N_3044,N_2410,N_21);
or U3045 (N_3045,N_1709,N_436);
or U3046 (N_3046,N_2367,N_184);
xnor U3047 (N_3047,N_2170,N_2300);
or U3048 (N_3048,N_1418,N_291);
nand U3049 (N_3049,N_709,N_161);
nor U3050 (N_3050,N_1251,N_2052);
or U3051 (N_3051,N_1232,N_236);
or U3052 (N_3052,N_1753,N_1596);
or U3053 (N_3053,N_2459,N_165);
nand U3054 (N_3054,N_390,N_1840);
nor U3055 (N_3055,N_187,N_904);
or U3056 (N_3056,N_364,N_227);
nor U3057 (N_3057,N_1735,N_2012);
nand U3058 (N_3058,N_895,N_479);
nor U3059 (N_3059,N_944,N_15);
nand U3060 (N_3060,N_1796,N_83);
xor U3061 (N_3061,N_1799,N_1592);
xnor U3062 (N_3062,N_1756,N_270);
or U3063 (N_3063,N_1983,N_213);
nand U3064 (N_3064,N_729,N_903);
and U3065 (N_3065,N_1907,N_833);
xor U3066 (N_3066,N_1748,N_1161);
xor U3067 (N_3067,N_76,N_1085);
xnor U3068 (N_3068,N_55,N_1105);
xnor U3069 (N_3069,N_75,N_182);
or U3070 (N_3070,N_2447,N_1404);
xor U3071 (N_3071,N_1384,N_588);
nor U3072 (N_3072,N_2040,N_859);
or U3073 (N_3073,N_138,N_611);
or U3074 (N_3074,N_562,N_91);
and U3075 (N_3075,N_1555,N_1554);
xor U3076 (N_3076,N_1880,N_211);
and U3077 (N_3077,N_1228,N_798);
nor U3078 (N_3078,N_579,N_1198);
and U3079 (N_3079,N_1011,N_1655);
and U3080 (N_3080,N_587,N_453);
nor U3081 (N_3081,N_926,N_510);
nor U3082 (N_3082,N_1170,N_425);
xnor U3083 (N_3083,N_2355,N_675);
and U3084 (N_3084,N_834,N_124);
or U3085 (N_3085,N_2213,N_2039);
nor U3086 (N_3086,N_1114,N_2215);
and U3087 (N_3087,N_647,N_1633);
nor U3088 (N_3088,N_367,N_368);
xor U3089 (N_3089,N_1720,N_1607);
nand U3090 (N_3090,N_1491,N_659);
or U3091 (N_3091,N_620,N_1705);
nor U3092 (N_3092,N_1392,N_862);
xnor U3093 (N_3093,N_366,N_2064);
or U3094 (N_3094,N_1916,N_1130);
or U3095 (N_3095,N_1905,N_2075);
or U3096 (N_3096,N_1306,N_452);
and U3097 (N_3097,N_2304,N_255);
or U3098 (N_3098,N_1197,N_1997);
or U3099 (N_3099,N_809,N_2302);
or U3100 (N_3100,N_1882,N_1952);
nand U3101 (N_3101,N_979,N_2148);
nand U3102 (N_3102,N_1268,N_183);
and U3103 (N_3103,N_700,N_1023);
nor U3104 (N_3104,N_799,N_1559);
or U3105 (N_3105,N_644,N_1342);
or U3106 (N_3106,N_2351,N_2020);
or U3107 (N_3107,N_670,N_1064);
and U3108 (N_3108,N_1766,N_378);
nor U3109 (N_3109,N_1825,N_1436);
nand U3110 (N_3110,N_901,N_1973);
and U3111 (N_3111,N_646,N_894);
nand U3112 (N_3112,N_577,N_802);
xor U3113 (N_3113,N_1315,N_2048);
nor U3114 (N_3114,N_764,N_520);
or U3115 (N_3115,N_574,N_1142);
xor U3116 (N_3116,N_295,N_966);
nor U3117 (N_3117,N_810,N_735);
and U3118 (N_3118,N_159,N_1144);
nor U3119 (N_3119,N_2218,N_2274);
nor U3120 (N_3120,N_1363,N_195);
nand U3121 (N_3121,N_249,N_1919);
nand U3122 (N_3122,N_2108,N_1460);
or U3123 (N_3123,N_2030,N_1617);
xor U3124 (N_3124,N_1913,N_121);
xnor U3125 (N_3125,N_715,N_1787);
xor U3126 (N_3126,N_1098,N_772);
nor U3127 (N_3127,N_1141,N_2090);
nand U3128 (N_3128,N_2309,N_982);
nor U3129 (N_3129,N_109,N_3);
or U3130 (N_3130,N_896,N_1765);
or U3131 (N_3131,N_1773,N_185);
nor U3132 (N_3132,N_1722,N_1398);
nand U3133 (N_3133,N_2050,N_1850);
nor U3134 (N_3134,N_1849,N_1445);
nand U3135 (N_3135,N_13,N_2069);
nand U3136 (N_3136,N_1255,N_657);
xnor U3137 (N_3137,N_416,N_889);
nor U3138 (N_3138,N_340,N_120);
or U3139 (N_3139,N_2347,N_1027);
and U3140 (N_3140,N_2159,N_1789);
xor U3141 (N_3141,N_2362,N_841);
nor U3142 (N_3142,N_1196,N_1202);
xnor U3143 (N_3143,N_925,N_98);
nand U3144 (N_3144,N_1075,N_408);
xor U3145 (N_3145,N_1321,N_542);
nor U3146 (N_3146,N_1059,N_2009);
nand U3147 (N_3147,N_85,N_2151);
nor U3148 (N_3148,N_963,N_2486);
or U3149 (N_3149,N_1996,N_868);
and U3150 (N_3150,N_2198,N_87);
nor U3151 (N_3151,N_19,N_573);
nand U3152 (N_3152,N_239,N_45);
and U3153 (N_3153,N_1758,N_2178);
and U3154 (N_3154,N_298,N_2004);
nand U3155 (N_3155,N_1494,N_1836);
and U3156 (N_3156,N_1539,N_1833);
or U3157 (N_3157,N_1993,N_1505);
xnor U3158 (N_3158,N_1051,N_781);
and U3159 (N_3159,N_1412,N_2496);
xnor U3160 (N_3160,N_827,N_1622);
nand U3161 (N_3161,N_2006,N_1659);
nor U3162 (N_3162,N_924,N_897);
xnor U3163 (N_3163,N_2432,N_1822);
and U3164 (N_3164,N_1119,N_1290);
and U3165 (N_3165,N_317,N_1511);
nor U3166 (N_3166,N_701,N_1496);
or U3167 (N_3167,N_1852,N_800);
nor U3168 (N_3168,N_1664,N_551);
xor U3169 (N_3169,N_1358,N_358);
nand U3170 (N_3170,N_2041,N_2289);
or U3171 (N_3171,N_803,N_1608);
nand U3172 (N_3172,N_2356,N_2095);
xnor U3173 (N_3173,N_2059,N_2279);
nor U3174 (N_3174,N_1904,N_176);
and U3175 (N_3175,N_2156,N_1526);
xor U3176 (N_3176,N_2255,N_353);
or U3177 (N_3177,N_565,N_1189);
nor U3178 (N_3178,N_1267,N_1803);
nand U3179 (N_3179,N_2419,N_617);
and U3180 (N_3180,N_20,N_501);
and U3181 (N_3181,N_264,N_750);
nor U3182 (N_3182,N_968,N_1538);
and U3183 (N_3183,N_1072,N_242);
nand U3184 (N_3184,N_306,N_330);
nand U3185 (N_3185,N_1382,N_1602);
nand U3186 (N_3186,N_1155,N_2423);
and U3187 (N_3187,N_1690,N_1420);
and U3188 (N_3188,N_575,N_2449);
nand U3189 (N_3189,N_66,N_2081);
or U3190 (N_3190,N_933,N_877);
nor U3191 (N_3191,N_1931,N_557);
or U3192 (N_3192,N_1647,N_1003);
and U3193 (N_3193,N_2303,N_910);
xnor U3194 (N_3194,N_545,N_1751);
and U3195 (N_3195,N_978,N_526);
and U3196 (N_3196,N_1821,N_1682);
nor U3197 (N_3197,N_88,N_1441);
nor U3198 (N_3198,N_84,N_1205);
or U3199 (N_3199,N_505,N_2429);
nor U3200 (N_3200,N_1451,N_725);
or U3201 (N_3201,N_2221,N_446);
nand U3202 (N_3202,N_2085,N_2428);
and U3203 (N_3203,N_18,N_1854);
nor U3204 (N_3204,N_2494,N_139);
or U3205 (N_3205,N_2229,N_1534);
nand U3206 (N_3206,N_2453,N_669);
and U3207 (N_3207,N_1159,N_626);
and U3208 (N_3208,N_484,N_443);
and U3209 (N_3209,N_1437,N_2413);
and U3210 (N_3210,N_1127,N_250);
xor U3211 (N_3211,N_405,N_544);
xor U3212 (N_3212,N_144,N_856);
and U3213 (N_3213,N_1832,N_2326);
nor U3214 (N_3214,N_1934,N_2446);
and U3215 (N_3215,N_945,N_2162);
or U3216 (N_3216,N_2067,N_221);
or U3217 (N_3217,N_2357,N_989);
or U3218 (N_3218,N_1045,N_814);
xor U3219 (N_3219,N_1684,N_464);
nand U3220 (N_3220,N_2220,N_1467);
and U3221 (N_3221,N_1893,N_1918);
nand U3222 (N_3222,N_1470,N_29);
nand U3223 (N_3223,N_2203,N_335);
and U3224 (N_3224,N_288,N_863);
or U3225 (N_3225,N_142,N_1221);
nand U3226 (N_3226,N_301,N_830);
nand U3227 (N_3227,N_1995,N_635);
and U3228 (N_3228,N_432,N_2184);
and U3229 (N_3229,N_1646,N_857);
or U3230 (N_3230,N_1463,N_2112);
nor U3231 (N_3231,N_705,N_902);
and U3232 (N_3232,N_94,N_1503);
and U3233 (N_3233,N_2424,N_2403);
nand U3234 (N_3234,N_2443,N_2019);
nor U3235 (N_3235,N_1178,N_1865);
and U3236 (N_3236,N_2387,N_2022);
and U3237 (N_3237,N_1455,N_1517);
nor U3238 (N_3238,N_2293,N_1468);
nor U3239 (N_3239,N_48,N_2165);
nor U3240 (N_3240,N_1132,N_417);
or U3241 (N_3241,N_370,N_131);
nor U3242 (N_3242,N_844,N_1049);
xnor U3243 (N_3243,N_1353,N_676);
nor U3244 (N_3244,N_253,N_1005);
and U3245 (N_3245,N_1859,N_1322);
and U3246 (N_3246,N_2160,N_1307);
nand U3247 (N_3247,N_843,N_2206);
nand U3248 (N_3248,N_1688,N_2345);
and U3249 (N_3249,N_915,N_1729);
nor U3250 (N_3250,N_2060,N_2036);
nand U3251 (N_3251,N_1067,N_2386);
and U3252 (N_3252,N_2338,N_1236);
nand U3253 (N_3253,N_2440,N_616);
xnor U3254 (N_3254,N_951,N_1344);
and U3255 (N_3255,N_115,N_2146);
nand U3256 (N_3256,N_1422,N_485);
nand U3257 (N_3257,N_117,N_1330);
or U3258 (N_3258,N_782,N_2167);
or U3259 (N_3259,N_518,N_46);
nor U3260 (N_3260,N_749,N_1706);
xnor U3261 (N_3261,N_1457,N_2234);
nor U3262 (N_3262,N_116,N_1754);
nand U3263 (N_3263,N_748,N_597);
and U3264 (N_3264,N_1749,N_1744);
and U3265 (N_3265,N_363,N_1025);
nor U3266 (N_3266,N_1693,N_1428);
nand U3267 (N_3267,N_2270,N_1128);
xor U3268 (N_3268,N_2467,N_2226);
or U3269 (N_3269,N_1139,N_2121);
or U3270 (N_3270,N_276,N_1978);
xor U3271 (N_3271,N_2306,N_2239);
nand U3272 (N_3272,N_1300,N_1207);
nor U3273 (N_3273,N_1733,N_716);
nor U3274 (N_3274,N_2097,N_586);
nand U3275 (N_3275,N_821,N_794);
nand U3276 (N_3276,N_1434,N_1943);
nor U3277 (N_3277,N_1906,N_1427);
or U3278 (N_3278,N_2244,N_2070);
or U3279 (N_3279,N_2131,N_1252);
or U3280 (N_3280,N_1061,N_780);
or U3281 (N_3281,N_1475,N_1213);
nor U3282 (N_3282,N_788,N_86);
and U3283 (N_3283,N_866,N_739);
or U3284 (N_3284,N_1914,N_49);
nor U3285 (N_3285,N_1724,N_238);
and U3286 (N_3286,N_1600,N_1248);
nor U3287 (N_3287,N_319,N_1738);
xor U3288 (N_3288,N_148,N_62);
or U3289 (N_3289,N_1270,N_2404);
nor U3290 (N_3290,N_1097,N_2245);
nor U3291 (N_3291,N_180,N_1626);
nand U3292 (N_3292,N_2235,N_2049);
and U3293 (N_3293,N_472,N_2430);
nor U3294 (N_3294,N_2122,N_1860);
or U3295 (N_3295,N_1776,N_871);
and U3296 (N_3296,N_1115,N_1728);
or U3297 (N_3297,N_899,N_860);
nor U3298 (N_3298,N_712,N_1359);
nor U3299 (N_3299,N_1911,N_2444);
nand U3300 (N_3300,N_783,N_952);
or U3301 (N_3301,N_2427,N_442);
or U3302 (N_3302,N_943,N_961);
xor U3303 (N_3303,N_1830,N_420);
and U3304 (N_3304,N_271,N_1458);
nand U3305 (N_3305,N_548,N_1287);
nand U3306 (N_3306,N_886,N_504);
nor U3307 (N_3307,N_1423,N_1385);
xor U3308 (N_3308,N_698,N_2499);
and U3309 (N_3309,N_1768,N_198);
and U3310 (N_3310,N_127,N_1365);
nor U3311 (N_3311,N_4,N_527);
nor U3312 (N_3312,N_1298,N_1487);
nand U3313 (N_3313,N_519,N_422);
nor U3314 (N_3314,N_1360,N_1106);
and U3315 (N_3315,N_5,N_1785);
and U3316 (N_3316,N_1439,N_1842);
xnor U3317 (N_3317,N_949,N_1998);
or U3318 (N_3318,N_1661,N_2285);
nand U3319 (N_3319,N_1623,N_2185);
nand U3320 (N_3320,N_920,N_888);
or U3321 (N_3321,N_1676,N_1537);
xor U3322 (N_3322,N_1043,N_825);
or U3323 (N_3323,N_202,N_1233);
xnor U3324 (N_3324,N_201,N_2024);
or U3325 (N_3325,N_959,N_838);
nand U3326 (N_3326,N_229,N_2461);
nor U3327 (N_3327,N_477,N_448);
nor U3328 (N_3328,N_1984,N_9);
nand U3329 (N_3329,N_1372,N_957);
nor U3330 (N_3330,N_530,N_692);
and U3331 (N_3331,N_1994,N_2261);
xnor U3332 (N_3332,N_1957,N_1673);
or U3333 (N_3333,N_224,N_680);
xor U3334 (N_3334,N_2331,N_878);
nand U3335 (N_3335,N_761,N_697);
nor U3336 (N_3336,N_621,N_1175);
nand U3337 (N_3337,N_105,N_2317);
xor U3338 (N_3338,N_1081,N_1872);
or U3339 (N_3339,N_1928,N_1576);
nor U3340 (N_3340,N_1763,N_480);
nor U3341 (N_3341,N_2407,N_932);
nor U3342 (N_3342,N_2476,N_2253);
nor U3343 (N_3343,N_2243,N_1320);
nand U3344 (N_3344,N_333,N_1991);
nor U3345 (N_3345,N_1147,N_1316);
and U3346 (N_3346,N_839,N_883);
or U3347 (N_3347,N_955,N_538);
or U3348 (N_3348,N_885,N_1779);
and U3349 (N_3349,N_71,N_1478);
nor U3350 (N_3350,N_634,N_230);
nand U3351 (N_3351,N_1504,N_1662);
nor U3352 (N_3352,N_70,N_990);
nand U3353 (N_3353,N_1407,N_2305);
xnor U3354 (N_3354,N_2065,N_909);
nor U3355 (N_3355,N_1829,N_1265);
nand U3356 (N_3356,N_1191,N_733);
and U3357 (N_3357,N_346,N_1241);
xnor U3358 (N_3358,N_1697,N_2342);
and U3359 (N_3359,N_1980,N_590);
and U3360 (N_3360,N_2257,N_2472);
nand U3361 (N_3361,N_2296,N_492);
or U3362 (N_3362,N_1301,N_629);
xnor U3363 (N_3363,N_1121,N_260);
or U3364 (N_3364,N_499,N_1702);
nand U3365 (N_3365,N_396,N_137);
xnor U3366 (N_3366,N_832,N_747);
nand U3367 (N_3367,N_1616,N_2478);
nor U3368 (N_3368,N_1446,N_2135);
and U3369 (N_3369,N_1054,N_300);
and U3370 (N_3370,N_867,N_2465);
and U3371 (N_3371,N_985,N_654);
nand U3372 (N_3372,N_1042,N_1158);
or U3373 (N_3373,N_1876,N_1988);
nand U3374 (N_3374,N_2406,N_592);
xor U3375 (N_3375,N_279,N_1631);
xor U3376 (N_3376,N_154,N_2456);
or U3377 (N_3377,N_2140,N_1846);
nor U3378 (N_3378,N_112,N_2014);
nand U3379 (N_3379,N_1713,N_939);
and U3380 (N_3380,N_1143,N_1453);
nand U3381 (N_3381,N_1313,N_232);
nor U3382 (N_3382,N_1374,N_1123);
nand U3383 (N_3383,N_954,N_1898);
or U3384 (N_3384,N_30,N_2396);
and U3385 (N_3385,N_1317,N_1704);
nand U3386 (N_3386,N_1603,N_693);
nor U3387 (N_3387,N_2132,N_1985);
xnor U3388 (N_3388,N_1666,N_2018);
nor U3389 (N_3389,N_1935,N_1974);
or U3390 (N_3390,N_256,N_1006);
nand U3391 (N_3391,N_191,N_2491);
xnor U3392 (N_3392,N_1718,N_682);
nor U3393 (N_3393,N_1855,N_2241);
or U3394 (N_3394,N_2373,N_462);
or U3395 (N_3395,N_1591,N_1979);
or U3396 (N_3396,N_406,N_1432);
and U3397 (N_3397,N_2445,N_1356);
xor U3398 (N_3398,N_1379,N_149);
nor U3399 (N_3399,N_679,N_2341);
xnor U3400 (N_3400,N_2225,N_292);
nand U3401 (N_3401,N_1925,N_2382);
nand U3402 (N_3402,N_1199,N_424);
or U3403 (N_3403,N_817,N_880);
nor U3404 (N_3404,N_1879,N_1823);
and U3405 (N_3405,N_1922,N_2171);
nor U3406 (N_3406,N_1089,N_152);
nor U3407 (N_3407,N_970,N_1263);
nor U3408 (N_3408,N_1482,N_891);
xnor U3409 (N_3409,N_2158,N_836);
nand U3410 (N_3410,N_141,N_1480);
xnor U3411 (N_3411,N_758,N_1396);
nor U3412 (N_3412,N_1095,N_277);
nand U3413 (N_3413,N_283,N_998);
xnor U3414 (N_3414,N_1261,N_1324);
nor U3415 (N_3415,N_1176,N_1711);
nand U3416 (N_3416,N_314,N_2348);
and U3417 (N_3417,N_356,N_1431);
nand U3418 (N_3418,N_2183,N_2358);
nor U3419 (N_3419,N_1150,N_171);
nand U3420 (N_3420,N_2201,N_1520);
nor U3421 (N_3421,N_851,N_900);
xnor U3422 (N_3422,N_37,N_1620);
nand U3423 (N_3423,N_365,N_153);
xnor U3424 (N_3424,N_690,N_2379);
nand U3425 (N_3425,N_2260,N_1654);
nand U3426 (N_3426,N_421,N_2232);
and U3427 (N_3427,N_826,N_600);
nor U3428 (N_3428,N_1747,N_410);
nand U3429 (N_3429,N_1260,N_2010);
nor U3430 (N_3430,N_2352,N_414);
or U3431 (N_3431,N_495,N_502);
xnor U3432 (N_3432,N_1348,N_2325);
and U3433 (N_3433,N_2128,N_2378);
nand U3434 (N_3434,N_134,N_482);
nand U3435 (N_3435,N_1046,N_2054);
nor U3436 (N_3436,N_1052,N_726);
and U3437 (N_3437,N_976,N_2088);
nand U3438 (N_3438,N_532,N_1571);
xor U3439 (N_3439,N_986,N_1456);
and U3440 (N_3440,N_694,N_2130);
nand U3441 (N_3441,N_1338,N_1050);
nor U3442 (N_3442,N_539,N_552);
and U3443 (N_3443,N_1506,N_1244);
or U3444 (N_3444,N_1719,N_450);
nand U3445 (N_3445,N_1156,N_496);
xnor U3446 (N_3446,N_1971,N_927);
and U3447 (N_3447,N_2047,N_549);
xor U3448 (N_3448,N_1010,N_2295);
xor U3449 (N_3449,N_2073,N_627);
xnor U3450 (N_3450,N_649,N_1845);
nor U3451 (N_3451,N_850,N_391);
nand U3452 (N_3452,N_1858,N_1086);
nor U3453 (N_3453,N_2177,N_2034);
nor U3454 (N_3454,N_1004,N_223);
and U3455 (N_3455,N_1816,N_1955);
nand U3456 (N_3456,N_285,N_785);
or U3457 (N_3457,N_2388,N_199);
nand U3458 (N_3458,N_1037,N_1129);
and U3459 (N_3459,N_1708,N_487);
xor U3460 (N_3460,N_1283,N_1715);
and U3461 (N_3461,N_1328,N_1419);
and U3462 (N_3462,N_1165,N_848);
and U3463 (N_3463,N_1116,N_876);
nor U3464 (N_3464,N_25,N_971);
nand U3465 (N_3465,N_1220,N_247);
and U3466 (N_3466,N_1282,N_2492);
xor U3467 (N_3467,N_382,N_2361);
or U3468 (N_3468,N_1533,N_1403);
nand U3469 (N_3469,N_1234,N_1361);
nand U3470 (N_3470,N_207,N_1164);
nand U3471 (N_3471,N_550,N_2313);
or U3472 (N_3472,N_1169,N_1308);
and U3473 (N_3473,N_2098,N_1256);
nor U3474 (N_3474,N_1442,N_2264);
nor U3475 (N_3475,N_2057,N_1762);
and U3476 (N_3476,N_2400,N_2182);
xor U3477 (N_3477,N_2334,N_1279);
xor U3478 (N_3478,N_412,N_1798);
and U3479 (N_3479,N_847,N_1295);
xnor U3480 (N_3480,N_194,N_246);
or U3481 (N_3481,N_2250,N_1354);
and U3482 (N_3482,N_1410,N_858);
nor U3483 (N_3483,N_428,N_222);
nor U3484 (N_3484,N_942,N_2191);
and U3485 (N_3485,N_2473,N_791);
nor U3486 (N_3486,N_290,N_375);
xor U3487 (N_3487,N_1513,N_1897);
nor U3488 (N_3488,N_993,N_770);
nand U3489 (N_3489,N_517,N_1540);
and U3490 (N_3490,N_401,N_786);
and U3491 (N_3491,N_2493,N_854);
and U3492 (N_3492,N_1030,N_686);
xnor U3493 (N_3493,N_493,N_1083);
nand U3494 (N_3494,N_262,N_1325);
xor U3495 (N_3495,N_1788,N_1107);
and U3496 (N_3496,N_2301,N_52);
xnor U3497 (N_3497,N_1881,N_1992);
nor U3498 (N_3498,N_1692,N_683);
or U3499 (N_3499,N_2124,N_228);
nor U3500 (N_3500,N_1853,N_1171);
nand U3501 (N_3501,N_1594,N_2216);
and U3502 (N_3502,N_2314,N_268);
nor U3503 (N_3503,N_2451,N_1448);
and U3504 (N_3504,N_622,N_1101);
nor U3505 (N_3505,N_1632,N_793);
nand U3506 (N_3506,N_874,N_2101);
and U3507 (N_3507,N_1531,N_2330);
and U3508 (N_3508,N_1770,N_1545);
or U3509 (N_3509,N_2231,N_767);
and U3510 (N_3510,N_42,N_427);
and U3511 (N_3511,N_1146,N_2161);
nor U3512 (N_3512,N_811,N_1663);
nand U3513 (N_3513,N_2222,N_946);
xnor U3514 (N_3514,N_589,N_997);
and U3515 (N_3515,N_1294,N_996);
nor U3516 (N_3516,N_1656,N_2287);
xnor U3517 (N_3517,N_2152,N_1237);
nand U3518 (N_3518,N_361,N_1564);
or U3519 (N_3519,N_99,N_162);
and U3520 (N_3520,N_394,N_1084);
and U3521 (N_3521,N_2468,N_1078);
xor U3522 (N_3522,N_928,N_1572);
and U3523 (N_3523,N_1329,N_1070);
nor U3524 (N_3524,N_936,N_245);
nor U3525 (N_3525,N_2217,N_2078);
nor U3526 (N_3526,N_2117,N_163);
nand U3527 (N_3527,N_1915,N_884);
or U3528 (N_3528,N_1800,N_2328);
nand U3529 (N_3529,N_2436,N_1548);
xor U3530 (N_3530,N_128,N_1110);
nor U3531 (N_3531,N_1976,N_1378);
nor U3532 (N_3532,N_999,N_2099);
and U3533 (N_3533,N_2488,N_1341);
xor U3534 (N_3534,N_1923,N_1152);
nand U3535 (N_3535,N_1941,N_1007);
nor U3536 (N_3536,N_988,N_331);
nand U3537 (N_3537,N_10,N_2068);
xnor U3538 (N_3538,N_386,N_150);
and U3539 (N_3539,N_511,N_1074);
nand U3540 (N_3540,N_660,N_114);
and U3541 (N_3541,N_1479,N_2026);
or U3542 (N_3542,N_1638,N_1956);
or U3543 (N_3543,N_2204,N_1117);
and U3544 (N_3544,N_1057,N_275);
and U3545 (N_3545,N_1355,N_934);
and U3546 (N_3546,N_1227,N_1019);
nor U3547 (N_3547,N_1285,N_1811);
nand U3548 (N_3548,N_1921,N_2118);
xnor U3549 (N_3549,N_2087,N_1166);
and U3550 (N_3550,N_2483,N_1305);
xor U3551 (N_3551,N_1781,N_2188);
or U3552 (N_3552,N_1337,N_11);
nand U3553 (N_3553,N_1549,N_1582);
nand U3554 (N_3554,N_533,N_852);
or U3555 (N_3555,N_741,N_1443);
xnor U3556 (N_3556,N_186,N_101);
or U3557 (N_3557,N_576,N_2133);
or U3558 (N_3558,N_563,N_1901);
or U3559 (N_3559,N_1643,N_835);
or U3560 (N_3560,N_1861,N_738);
or U3561 (N_3561,N_97,N_1593);
xnor U3562 (N_3562,N_233,N_345);
nor U3563 (N_3563,N_2441,N_218);
nor U3564 (N_3564,N_1945,N_1819);
or U3565 (N_3565,N_1869,N_1406);
and U3566 (N_3566,N_1793,N_1568);
nand U3567 (N_3567,N_1624,N_628);
xnor U3568 (N_3568,N_129,N_237);
xor U3569 (N_3569,N_96,N_2434);
or U3570 (N_3570,N_1717,N_1391);
and U3571 (N_3571,N_326,N_1801);
and U3572 (N_3572,N_908,N_1088);
nor U3573 (N_3573,N_1058,N_437);
nor U3574 (N_3574,N_2007,N_2046);
nor U3575 (N_3575,N_706,N_1216);
nand U3576 (N_3576,N_2016,N_631);
and U3577 (N_3577,N_1257,N_730);
nor U3578 (N_3578,N_1126,N_842);
nor U3579 (N_3579,N_2082,N_815);
and U3580 (N_3580,N_1181,N_1886);
and U3581 (N_3581,N_476,N_606);
nand U3582 (N_3582,N_2475,N_1551);
and U3583 (N_3583,N_118,N_100);
or U3584 (N_3584,N_1871,N_1887);
xnor U3585 (N_3585,N_329,N_1108);
nor U3586 (N_3586,N_1550,N_1474);
nand U3587 (N_3587,N_1426,N_1471);
xor U3588 (N_3588,N_991,N_721);
or U3589 (N_3589,N_231,N_1204);
or U3590 (N_3590,N_1000,N_813);
or U3591 (N_3591,N_2298,N_1430);
xor U3592 (N_3592,N_376,N_655);
or U3593 (N_3593,N_1332,N_1424);
nor U3594 (N_3594,N_1970,N_1433);
xor U3595 (N_3595,N_2119,N_1449);
xor U3596 (N_3596,N_1723,N_1334);
nand U3597 (N_3597,N_2288,N_1908);
or U3598 (N_3598,N_623,N_2200);
nand U3599 (N_3599,N_1134,N_1657);
nor U3600 (N_3600,N_953,N_388);
xnor U3601 (N_3601,N_2233,N_1041);
and U3602 (N_3602,N_678,N_297);
nand U3603 (N_3603,N_777,N_921);
nor U3604 (N_3604,N_1459,N_2242);
xnor U3605 (N_3605,N_756,N_1239);
and U3606 (N_3606,N_1215,N_2037);
and U3607 (N_3607,N_1413,N_2393);
or U3608 (N_3608,N_2282,N_478);
nor U3609 (N_3609,N_93,N_947);
nand U3610 (N_3610,N_1653,N_829);
xor U3611 (N_3611,N_1668,N_2359);
nand U3612 (N_3612,N_1667,N_1055);
and U3613 (N_3613,N_1902,N_916);
nand U3614 (N_3614,N_310,N_1967);
and U3615 (N_3615,N_1409,N_2319);
or U3616 (N_3616,N_1323,N_775);
and U3617 (N_3617,N_1180,N_1281);
nand U3618 (N_3618,N_1472,N_855);
nor U3619 (N_3619,N_315,N_1195);
or U3620 (N_3620,N_313,N_684);
xnor U3621 (N_3621,N_707,N_1611);
or U3622 (N_3622,N_974,N_2147);
and U3623 (N_3623,N_1347,N_104);
or U3624 (N_3624,N_170,N_1352);
xnor U3625 (N_3625,N_1217,N_77);
xor U3626 (N_3626,N_2318,N_2113);
and U3627 (N_3627,N_289,N_380);
and U3628 (N_3628,N_2079,N_1707);
and U3629 (N_3629,N_1015,N_1658);
or U3630 (N_3630,N_1369,N_494);
or U3631 (N_3631,N_1856,N_652);
or U3632 (N_3632,N_385,N_1774);
nor U3633 (N_3633,N_2246,N_992);
and U3634 (N_3634,N_1021,N_1231);
nor U3635 (N_3635,N_595,N_1972);
or U3636 (N_3636,N_2385,N_1597);
nand U3637 (N_3637,N_344,N_438);
or U3638 (N_3638,N_2149,N_1837);
xor U3639 (N_3639,N_2397,N_1581);
or U3640 (N_3640,N_806,N_1464);
nand U3641 (N_3641,N_1806,N_645);
or U3642 (N_3642,N_2166,N_2103);
and U3643 (N_3643,N_879,N_1639);
nand U3644 (N_3644,N_392,N_1595);
nor U3645 (N_3645,N_1585,N_666);
and U3646 (N_3646,N_1185,N_556);
and U3647 (N_3647,N_1376,N_1408);
nor U3648 (N_3648,N_1792,N_801);
or U3649 (N_3649,N_818,N_2091);
and U3650 (N_3650,N_407,N_1492);
or U3651 (N_3651,N_332,N_1039);
nor U3652 (N_3652,N_1351,N_1675);
and U3653 (N_3653,N_440,N_287);
and U3654 (N_3654,N_553,N_1077);
nand U3655 (N_3655,N_1628,N_1076);
or U3656 (N_3656,N_284,N_36);
nand U3657 (N_3657,N_1184,N_355);
nand U3658 (N_3658,N_445,N_1930);
nor U3659 (N_3659,N_1529,N_2417);
nor U3660 (N_3660,N_805,N_665);
xor U3661 (N_3661,N_797,N_2329);
or U3662 (N_3662,N_912,N_1714);
nor U3663 (N_3663,N_1521,N_2137);
xnor U3664 (N_3664,N_807,N_1193);
nand U3665 (N_3665,N_2193,N_917);
or U3666 (N_3666,N_2437,N_1186);
nor U3667 (N_3667,N_451,N_702);
and U3668 (N_3668,N_1038,N_24);
nand U3669 (N_3669,N_2236,N_203);
xnor U3670 (N_3670,N_146,N_2163);
nand U3671 (N_3671,N_710,N_547);
or U3672 (N_3672,N_1497,N_1103);
nand U3673 (N_3673,N_2286,N_2035);
and U3674 (N_3674,N_1940,N_1111);
and U3675 (N_3675,N_1080,N_604);
and U3676 (N_3676,N_1024,N_525);
xor U3677 (N_3677,N_349,N_1099);
or U3678 (N_3678,N_610,N_1969);
nor U3679 (N_3679,N_804,N_1780);
and U3680 (N_3680,N_956,N_1488);
xnor U3681 (N_3681,N_1259,N_656);
nand U3682 (N_3682,N_2189,N_650);
nor U3683 (N_3683,N_2227,N_2125);
xor U3684 (N_3684,N_2169,N_2141);
nand U3685 (N_3685,N_393,N_913);
or U3686 (N_3686,N_471,N_776);
and U3687 (N_3687,N_1678,N_258);
and U3688 (N_3688,N_357,N_1742);
and U3689 (N_3689,N_243,N_1936);
or U3690 (N_3690,N_273,N_214);
nor U3691 (N_3691,N_1812,N_2268);
or U3692 (N_3692,N_1140,N_387);
nor U3693 (N_3693,N_1795,N_663);
xnor U3694 (N_3694,N_2412,N_1102);
nand U3695 (N_3695,N_731,N_58);
nand U3696 (N_3696,N_1414,N_2340);
nor U3697 (N_3697,N_318,N_1767);
or U3698 (N_3698,N_2391,N_2144);
nand U3699 (N_3699,N_743,N_2240);
xor U3700 (N_3700,N_537,N_601);
xnor U3701 (N_3701,N_2061,N_2084);
or U3702 (N_3702,N_312,N_1694);
or U3703 (N_3703,N_38,N_61);
xnor U3704 (N_3704,N_2454,N_1672);
nor U3705 (N_3705,N_1501,N_1797);
nor U3706 (N_3706,N_2256,N_571);
or U3707 (N_3707,N_1701,N_1264);
and U3708 (N_3708,N_309,N_1946);
and U3709 (N_3709,N_1524,N_2015);
and U3710 (N_3710,N_1273,N_402);
xor U3711 (N_3711,N_2017,N_779);
xnor U3712 (N_3712,N_2336,N_431);
nand U3713 (N_3713,N_147,N_1977);
nor U3714 (N_3714,N_1292,N_2263);
nand U3715 (N_3715,N_286,N_514);
or U3716 (N_3716,N_1848,N_1235);
nand U3717 (N_3717,N_193,N_1033);
or U3718 (N_3718,N_89,N_1509);
and U3719 (N_3719,N_449,N_2109);
nand U3720 (N_3720,N_1965,N_1149);
and U3721 (N_3721,N_1002,N_311);
nor U3722 (N_3722,N_384,N_1933);
nor U3723 (N_3723,N_2346,N_441);
and U3724 (N_3724,N_718,N_2228);
nor U3725 (N_3725,N_1048,N_773);
or U3726 (N_3726,N_1258,N_1588);
nand U3727 (N_3727,N_1314,N_403);
nand U3728 (N_3728,N_1912,N_72);
nand U3729 (N_3729,N_2173,N_342);
nor U3730 (N_3730,N_508,N_2384);
or U3731 (N_3731,N_2466,N_1981);
or U3732 (N_3732,N_1962,N_155);
or U3733 (N_3733,N_1400,N_430);
xnor U3734 (N_3734,N_2452,N_110);
and U3735 (N_3735,N_965,N_2072);
nor U3736 (N_3736,N_2495,N_1937);
nand U3737 (N_3737,N_324,N_1020);
and U3738 (N_3738,N_1183,N_1417);
nor U3739 (N_3739,N_1864,N_1621);
and U3740 (N_3740,N_930,N_1999);
nor U3741 (N_3741,N_1469,N_2294);
xor U3742 (N_3742,N_1557,N_873);
or U3743 (N_3743,N_489,N_458);
xor U3744 (N_3744,N_2142,N_637);
nand U3745 (N_3745,N_1606,N_2337);
and U3746 (N_3746,N_931,N_1625);
xnor U3747 (N_3747,N_2063,N_583);
nor U3748 (N_3748,N_1573,N_1782);
nand U3749 (N_3749,N_1964,N_570);
or U3750 (N_3750,N_1375,N_2226);
xor U3751 (N_3751,N_1534,N_2267);
nor U3752 (N_3752,N_136,N_1928);
xnor U3753 (N_3753,N_1933,N_1033);
or U3754 (N_3754,N_182,N_85);
and U3755 (N_3755,N_1327,N_1128);
or U3756 (N_3756,N_1420,N_79);
xor U3757 (N_3757,N_1021,N_1609);
xnor U3758 (N_3758,N_855,N_1767);
nand U3759 (N_3759,N_757,N_2312);
and U3760 (N_3760,N_1854,N_815);
and U3761 (N_3761,N_1348,N_633);
nand U3762 (N_3762,N_1627,N_2025);
and U3763 (N_3763,N_933,N_1433);
or U3764 (N_3764,N_2067,N_431);
nand U3765 (N_3765,N_1728,N_444);
nand U3766 (N_3766,N_1443,N_516);
nor U3767 (N_3767,N_2131,N_663);
and U3768 (N_3768,N_2314,N_183);
nand U3769 (N_3769,N_1466,N_767);
and U3770 (N_3770,N_1962,N_2305);
and U3771 (N_3771,N_972,N_338);
nand U3772 (N_3772,N_359,N_1486);
and U3773 (N_3773,N_397,N_892);
xnor U3774 (N_3774,N_1299,N_2004);
nand U3775 (N_3775,N_1211,N_1109);
nor U3776 (N_3776,N_1585,N_1462);
and U3777 (N_3777,N_604,N_2196);
nor U3778 (N_3778,N_71,N_1618);
xnor U3779 (N_3779,N_1143,N_1947);
nand U3780 (N_3780,N_75,N_2433);
and U3781 (N_3781,N_2174,N_1206);
xor U3782 (N_3782,N_1787,N_1539);
xor U3783 (N_3783,N_1922,N_1542);
xnor U3784 (N_3784,N_1678,N_897);
and U3785 (N_3785,N_701,N_1889);
nor U3786 (N_3786,N_1882,N_2213);
and U3787 (N_3787,N_263,N_2036);
or U3788 (N_3788,N_1874,N_1706);
nand U3789 (N_3789,N_1594,N_1769);
nand U3790 (N_3790,N_1070,N_291);
xor U3791 (N_3791,N_715,N_1435);
xnor U3792 (N_3792,N_890,N_0);
or U3793 (N_3793,N_2213,N_1740);
or U3794 (N_3794,N_1915,N_1181);
nor U3795 (N_3795,N_2496,N_605);
nor U3796 (N_3796,N_976,N_434);
nand U3797 (N_3797,N_595,N_2317);
and U3798 (N_3798,N_1306,N_859);
or U3799 (N_3799,N_1588,N_1534);
nor U3800 (N_3800,N_2020,N_1453);
and U3801 (N_3801,N_1358,N_1554);
and U3802 (N_3802,N_1492,N_1233);
xnor U3803 (N_3803,N_1746,N_622);
xor U3804 (N_3804,N_950,N_915);
nand U3805 (N_3805,N_1236,N_463);
or U3806 (N_3806,N_2494,N_1161);
nor U3807 (N_3807,N_2457,N_2310);
nand U3808 (N_3808,N_1512,N_82);
and U3809 (N_3809,N_1297,N_1699);
and U3810 (N_3810,N_795,N_528);
or U3811 (N_3811,N_354,N_502);
nand U3812 (N_3812,N_1668,N_52);
nand U3813 (N_3813,N_1078,N_673);
nor U3814 (N_3814,N_756,N_732);
xnor U3815 (N_3815,N_385,N_1299);
and U3816 (N_3816,N_1032,N_579);
nor U3817 (N_3817,N_2439,N_1120);
and U3818 (N_3818,N_949,N_1049);
and U3819 (N_3819,N_2469,N_1177);
or U3820 (N_3820,N_2183,N_421);
or U3821 (N_3821,N_1149,N_1532);
xnor U3822 (N_3822,N_965,N_1407);
xnor U3823 (N_3823,N_1325,N_1495);
and U3824 (N_3824,N_620,N_14);
nand U3825 (N_3825,N_850,N_1224);
nor U3826 (N_3826,N_672,N_779);
nor U3827 (N_3827,N_1778,N_1662);
xnor U3828 (N_3828,N_2045,N_1480);
or U3829 (N_3829,N_2317,N_188);
nand U3830 (N_3830,N_1544,N_289);
and U3831 (N_3831,N_1193,N_1747);
nor U3832 (N_3832,N_2155,N_1056);
or U3833 (N_3833,N_975,N_2082);
and U3834 (N_3834,N_621,N_733);
nand U3835 (N_3835,N_1413,N_793);
nand U3836 (N_3836,N_259,N_665);
nand U3837 (N_3837,N_1456,N_310);
nand U3838 (N_3838,N_1615,N_1058);
nand U3839 (N_3839,N_594,N_1691);
xnor U3840 (N_3840,N_953,N_1991);
or U3841 (N_3841,N_2344,N_2366);
or U3842 (N_3842,N_1623,N_231);
nand U3843 (N_3843,N_17,N_2446);
nor U3844 (N_3844,N_1164,N_1796);
nand U3845 (N_3845,N_119,N_1280);
and U3846 (N_3846,N_144,N_887);
xnor U3847 (N_3847,N_651,N_2118);
nor U3848 (N_3848,N_73,N_1297);
xor U3849 (N_3849,N_2107,N_779);
nor U3850 (N_3850,N_754,N_2161);
and U3851 (N_3851,N_1113,N_689);
nand U3852 (N_3852,N_1525,N_678);
or U3853 (N_3853,N_6,N_428);
or U3854 (N_3854,N_2468,N_1757);
nor U3855 (N_3855,N_1508,N_2108);
nor U3856 (N_3856,N_805,N_948);
nor U3857 (N_3857,N_1690,N_1953);
nor U3858 (N_3858,N_1659,N_1963);
nand U3859 (N_3859,N_1840,N_2064);
nor U3860 (N_3860,N_555,N_1158);
nor U3861 (N_3861,N_1305,N_303);
xnor U3862 (N_3862,N_1757,N_580);
nor U3863 (N_3863,N_1179,N_1596);
nand U3864 (N_3864,N_2214,N_469);
or U3865 (N_3865,N_1830,N_990);
and U3866 (N_3866,N_2287,N_49);
and U3867 (N_3867,N_1933,N_1889);
nand U3868 (N_3868,N_448,N_1402);
nor U3869 (N_3869,N_1464,N_1535);
nor U3870 (N_3870,N_2490,N_1042);
or U3871 (N_3871,N_1963,N_1410);
or U3872 (N_3872,N_2489,N_193);
and U3873 (N_3873,N_2382,N_926);
nor U3874 (N_3874,N_1499,N_2204);
and U3875 (N_3875,N_2414,N_1518);
nand U3876 (N_3876,N_1691,N_1150);
and U3877 (N_3877,N_256,N_84);
nor U3878 (N_3878,N_2097,N_2010);
xor U3879 (N_3879,N_1662,N_1931);
or U3880 (N_3880,N_1879,N_308);
nand U3881 (N_3881,N_84,N_2171);
or U3882 (N_3882,N_2132,N_656);
or U3883 (N_3883,N_2227,N_2374);
nand U3884 (N_3884,N_1679,N_570);
and U3885 (N_3885,N_1605,N_2493);
nand U3886 (N_3886,N_1410,N_2076);
and U3887 (N_3887,N_446,N_610);
nand U3888 (N_3888,N_1149,N_1537);
nor U3889 (N_3889,N_591,N_294);
xor U3890 (N_3890,N_1214,N_2395);
and U3891 (N_3891,N_386,N_2426);
nor U3892 (N_3892,N_1017,N_2466);
or U3893 (N_3893,N_1312,N_2404);
nand U3894 (N_3894,N_1691,N_1738);
nor U3895 (N_3895,N_2183,N_2300);
nor U3896 (N_3896,N_2155,N_2044);
or U3897 (N_3897,N_544,N_524);
nand U3898 (N_3898,N_2459,N_1265);
or U3899 (N_3899,N_511,N_1902);
nand U3900 (N_3900,N_1374,N_931);
nand U3901 (N_3901,N_1747,N_1159);
or U3902 (N_3902,N_145,N_1797);
nand U3903 (N_3903,N_1157,N_2062);
and U3904 (N_3904,N_401,N_1964);
nor U3905 (N_3905,N_826,N_370);
xnor U3906 (N_3906,N_544,N_342);
or U3907 (N_3907,N_2156,N_1003);
or U3908 (N_3908,N_1168,N_347);
nor U3909 (N_3909,N_1388,N_1191);
and U3910 (N_3910,N_577,N_2193);
xor U3911 (N_3911,N_1352,N_59);
nand U3912 (N_3912,N_1396,N_937);
and U3913 (N_3913,N_2026,N_2060);
nor U3914 (N_3914,N_1891,N_1441);
xnor U3915 (N_3915,N_1814,N_2395);
nand U3916 (N_3916,N_1659,N_2475);
nor U3917 (N_3917,N_1590,N_1761);
xnor U3918 (N_3918,N_27,N_1108);
or U3919 (N_3919,N_717,N_1218);
nor U3920 (N_3920,N_1651,N_1365);
nor U3921 (N_3921,N_1232,N_255);
xor U3922 (N_3922,N_1186,N_201);
nand U3923 (N_3923,N_1442,N_2087);
or U3924 (N_3924,N_532,N_1385);
and U3925 (N_3925,N_2012,N_63);
and U3926 (N_3926,N_1757,N_1129);
or U3927 (N_3927,N_1487,N_626);
or U3928 (N_3928,N_391,N_924);
xor U3929 (N_3929,N_2281,N_43);
and U3930 (N_3930,N_1632,N_2444);
nor U3931 (N_3931,N_2058,N_656);
or U3932 (N_3932,N_1412,N_522);
or U3933 (N_3933,N_2387,N_1146);
xnor U3934 (N_3934,N_1097,N_9);
or U3935 (N_3935,N_353,N_2151);
or U3936 (N_3936,N_1961,N_2484);
xor U3937 (N_3937,N_1002,N_1643);
nor U3938 (N_3938,N_319,N_1162);
nand U3939 (N_3939,N_828,N_1229);
or U3940 (N_3940,N_2406,N_2065);
xnor U3941 (N_3941,N_2388,N_585);
nor U3942 (N_3942,N_1081,N_1285);
xor U3943 (N_3943,N_2067,N_1686);
and U3944 (N_3944,N_2189,N_488);
nand U3945 (N_3945,N_321,N_1980);
or U3946 (N_3946,N_555,N_1284);
nand U3947 (N_3947,N_369,N_338);
and U3948 (N_3948,N_568,N_392);
or U3949 (N_3949,N_2280,N_2409);
nor U3950 (N_3950,N_2471,N_533);
or U3951 (N_3951,N_2409,N_407);
and U3952 (N_3952,N_2094,N_1762);
xor U3953 (N_3953,N_758,N_1889);
or U3954 (N_3954,N_343,N_1170);
nand U3955 (N_3955,N_2201,N_1559);
nor U3956 (N_3956,N_1067,N_1560);
nand U3957 (N_3957,N_1839,N_1900);
xor U3958 (N_3958,N_1446,N_1942);
nor U3959 (N_3959,N_706,N_188);
and U3960 (N_3960,N_591,N_1462);
or U3961 (N_3961,N_20,N_166);
nor U3962 (N_3962,N_107,N_206);
and U3963 (N_3963,N_1801,N_1334);
and U3964 (N_3964,N_306,N_1370);
and U3965 (N_3965,N_2139,N_2365);
and U3966 (N_3966,N_1577,N_378);
nor U3967 (N_3967,N_1691,N_1358);
nand U3968 (N_3968,N_629,N_1592);
and U3969 (N_3969,N_1692,N_713);
nor U3970 (N_3970,N_563,N_1076);
nand U3971 (N_3971,N_2490,N_2072);
or U3972 (N_3972,N_2324,N_156);
nor U3973 (N_3973,N_241,N_1204);
xnor U3974 (N_3974,N_616,N_1749);
and U3975 (N_3975,N_441,N_217);
nand U3976 (N_3976,N_343,N_288);
nor U3977 (N_3977,N_2158,N_2359);
nor U3978 (N_3978,N_1498,N_72);
and U3979 (N_3979,N_2440,N_1254);
nor U3980 (N_3980,N_969,N_570);
nand U3981 (N_3981,N_656,N_732);
xor U3982 (N_3982,N_2379,N_1242);
and U3983 (N_3983,N_1016,N_1269);
or U3984 (N_3984,N_1641,N_502);
nand U3985 (N_3985,N_1170,N_421);
and U3986 (N_3986,N_2328,N_1375);
xnor U3987 (N_3987,N_1561,N_2444);
xor U3988 (N_3988,N_2017,N_231);
or U3989 (N_3989,N_1638,N_869);
xor U3990 (N_3990,N_2433,N_1077);
xor U3991 (N_3991,N_244,N_753);
nor U3992 (N_3992,N_2436,N_1362);
nor U3993 (N_3993,N_1204,N_1961);
xnor U3994 (N_3994,N_2454,N_943);
nand U3995 (N_3995,N_1404,N_59);
nand U3996 (N_3996,N_1283,N_564);
nand U3997 (N_3997,N_2453,N_1158);
nor U3998 (N_3998,N_1931,N_60);
xor U3999 (N_3999,N_1753,N_2182);
nand U4000 (N_4000,N_886,N_2188);
nor U4001 (N_4001,N_2361,N_451);
xor U4002 (N_4002,N_287,N_1070);
nor U4003 (N_4003,N_2164,N_1823);
xnor U4004 (N_4004,N_1030,N_822);
or U4005 (N_4005,N_1769,N_28);
or U4006 (N_4006,N_387,N_1883);
nor U4007 (N_4007,N_2115,N_2347);
and U4008 (N_4008,N_593,N_1817);
and U4009 (N_4009,N_203,N_441);
and U4010 (N_4010,N_614,N_2255);
nand U4011 (N_4011,N_1700,N_2053);
or U4012 (N_4012,N_1719,N_1746);
and U4013 (N_4013,N_1873,N_2306);
nand U4014 (N_4014,N_1774,N_1220);
and U4015 (N_4015,N_1514,N_42);
and U4016 (N_4016,N_1585,N_762);
or U4017 (N_4017,N_459,N_1013);
nor U4018 (N_4018,N_1657,N_268);
xor U4019 (N_4019,N_1295,N_852);
nor U4020 (N_4020,N_227,N_1721);
and U4021 (N_4021,N_1013,N_1406);
nor U4022 (N_4022,N_739,N_1877);
nand U4023 (N_4023,N_729,N_2453);
and U4024 (N_4024,N_2378,N_2295);
xnor U4025 (N_4025,N_868,N_125);
nand U4026 (N_4026,N_1765,N_290);
or U4027 (N_4027,N_1858,N_313);
nor U4028 (N_4028,N_203,N_2138);
xnor U4029 (N_4029,N_1300,N_1433);
xor U4030 (N_4030,N_2344,N_2239);
nor U4031 (N_4031,N_2370,N_664);
and U4032 (N_4032,N_821,N_880);
nand U4033 (N_4033,N_2441,N_142);
nand U4034 (N_4034,N_575,N_2446);
xnor U4035 (N_4035,N_1264,N_1029);
and U4036 (N_4036,N_783,N_1825);
nand U4037 (N_4037,N_674,N_1337);
and U4038 (N_4038,N_385,N_1042);
or U4039 (N_4039,N_1761,N_1783);
nand U4040 (N_4040,N_1362,N_2042);
xor U4041 (N_4041,N_480,N_2248);
or U4042 (N_4042,N_2496,N_571);
nor U4043 (N_4043,N_1437,N_1092);
and U4044 (N_4044,N_926,N_535);
and U4045 (N_4045,N_2132,N_2365);
xor U4046 (N_4046,N_56,N_2287);
nand U4047 (N_4047,N_1245,N_1430);
or U4048 (N_4048,N_2146,N_1786);
or U4049 (N_4049,N_1796,N_1515);
nand U4050 (N_4050,N_1341,N_1238);
or U4051 (N_4051,N_2047,N_1871);
or U4052 (N_4052,N_1872,N_2177);
xnor U4053 (N_4053,N_175,N_1016);
xnor U4054 (N_4054,N_1557,N_2351);
xor U4055 (N_4055,N_1035,N_1118);
or U4056 (N_4056,N_2147,N_2249);
nand U4057 (N_4057,N_1076,N_2090);
or U4058 (N_4058,N_1133,N_1207);
nand U4059 (N_4059,N_1797,N_758);
and U4060 (N_4060,N_1493,N_1884);
and U4061 (N_4061,N_1193,N_632);
nand U4062 (N_4062,N_572,N_266);
nor U4063 (N_4063,N_67,N_288);
and U4064 (N_4064,N_2367,N_968);
nand U4065 (N_4065,N_2060,N_923);
nor U4066 (N_4066,N_1497,N_7);
or U4067 (N_4067,N_937,N_922);
nand U4068 (N_4068,N_877,N_1860);
nor U4069 (N_4069,N_1664,N_1116);
and U4070 (N_4070,N_122,N_348);
xor U4071 (N_4071,N_1980,N_661);
nor U4072 (N_4072,N_2304,N_890);
or U4073 (N_4073,N_2117,N_349);
nand U4074 (N_4074,N_1728,N_1558);
and U4075 (N_4075,N_869,N_1304);
and U4076 (N_4076,N_2422,N_2287);
or U4077 (N_4077,N_1299,N_2224);
and U4078 (N_4078,N_738,N_1141);
xnor U4079 (N_4079,N_2405,N_2478);
and U4080 (N_4080,N_785,N_811);
and U4081 (N_4081,N_319,N_1845);
nor U4082 (N_4082,N_1157,N_1577);
and U4083 (N_4083,N_1269,N_1518);
nor U4084 (N_4084,N_574,N_399);
nor U4085 (N_4085,N_1941,N_2061);
xnor U4086 (N_4086,N_1806,N_868);
nand U4087 (N_4087,N_2374,N_866);
xor U4088 (N_4088,N_1338,N_108);
and U4089 (N_4089,N_1901,N_1768);
xor U4090 (N_4090,N_1466,N_15);
nand U4091 (N_4091,N_751,N_1560);
nor U4092 (N_4092,N_442,N_1306);
or U4093 (N_4093,N_2494,N_1675);
nor U4094 (N_4094,N_786,N_622);
xnor U4095 (N_4095,N_2489,N_170);
nand U4096 (N_4096,N_362,N_683);
nand U4097 (N_4097,N_2066,N_806);
nand U4098 (N_4098,N_1639,N_1497);
xnor U4099 (N_4099,N_1135,N_1909);
or U4100 (N_4100,N_874,N_537);
or U4101 (N_4101,N_1651,N_1523);
nor U4102 (N_4102,N_1774,N_1983);
nand U4103 (N_4103,N_2104,N_1904);
xor U4104 (N_4104,N_432,N_785);
xor U4105 (N_4105,N_1308,N_886);
and U4106 (N_4106,N_186,N_1632);
xnor U4107 (N_4107,N_949,N_2380);
nor U4108 (N_4108,N_869,N_519);
or U4109 (N_4109,N_249,N_1820);
or U4110 (N_4110,N_174,N_2212);
nor U4111 (N_4111,N_1238,N_2096);
nand U4112 (N_4112,N_1183,N_580);
and U4113 (N_4113,N_1459,N_1398);
nor U4114 (N_4114,N_2186,N_460);
xor U4115 (N_4115,N_2428,N_1735);
or U4116 (N_4116,N_314,N_638);
nor U4117 (N_4117,N_1826,N_1816);
nand U4118 (N_4118,N_329,N_540);
or U4119 (N_4119,N_45,N_1720);
xnor U4120 (N_4120,N_1199,N_2497);
or U4121 (N_4121,N_1706,N_381);
nor U4122 (N_4122,N_2227,N_1416);
and U4123 (N_4123,N_810,N_1724);
nand U4124 (N_4124,N_2157,N_273);
or U4125 (N_4125,N_1840,N_642);
nand U4126 (N_4126,N_2462,N_153);
and U4127 (N_4127,N_2476,N_95);
and U4128 (N_4128,N_520,N_2108);
nor U4129 (N_4129,N_1520,N_756);
nand U4130 (N_4130,N_694,N_1698);
nor U4131 (N_4131,N_496,N_1358);
nand U4132 (N_4132,N_2176,N_1745);
nor U4133 (N_4133,N_64,N_728);
nand U4134 (N_4134,N_894,N_1883);
xor U4135 (N_4135,N_1965,N_82);
nand U4136 (N_4136,N_628,N_1540);
and U4137 (N_4137,N_1375,N_1644);
nor U4138 (N_4138,N_680,N_110);
nor U4139 (N_4139,N_1219,N_2171);
nand U4140 (N_4140,N_628,N_815);
xor U4141 (N_4141,N_1806,N_175);
and U4142 (N_4142,N_53,N_2463);
nor U4143 (N_4143,N_1125,N_1836);
nand U4144 (N_4144,N_2209,N_2100);
and U4145 (N_4145,N_2103,N_184);
nor U4146 (N_4146,N_2372,N_302);
or U4147 (N_4147,N_350,N_2189);
nand U4148 (N_4148,N_2372,N_680);
or U4149 (N_4149,N_2272,N_2152);
nor U4150 (N_4150,N_1507,N_253);
nor U4151 (N_4151,N_410,N_1641);
nor U4152 (N_4152,N_2426,N_1533);
xor U4153 (N_4153,N_870,N_1650);
xnor U4154 (N_4154,N_1456,N_1342);
and U4155 (N_4155,N_27,N_1455);
xnor U4156 (N_4156,N_104,N_1373);
nand U4157 (N_4157,N_1644,N_2016);
xnor U4158 (N_4158,N_524,N_157);
xor U4159 (N_4159,N_1693,N_856);
xor U4160 (N_4160,N_728,N_990);
and U4161 (N_4161,N_1601,N_390);
xor U4162 (N_4162,N_875,N_142);
and U4163 (N_4163,N_2053,N_2418);
nand U4164 (N_4164,N_159,N_1520);
nor U4165 (N_4165,N_1357,N_504);
and U4166 (N_4166,N_568,N_800);
xnor U4167 (N_4167,N_1646,N_2027);
nor U4168 (N_4168,N_2283,N_1713);
xnor U4169 (N_4169,N_1526,N_1231);
or U4170 (N_4170,N_818,N_981);
xnor U4171 (N_4171,N_2199,N_1742);
nand U4172 (N_4172,N_2003,N_1019);
xnor U4173 (N_4173,N_1370,N_2020);
or U4174 (N_4174,N_1186,N_508);
or U4175 (N_4175,N_1822,N_1283);
nand U4176 (N_4176,N_1547,N_2025);
and U4177 (N_4177,N_1379,N_102);
nand U4178 (N_4178,N_458,N_2334);
nand U4179 (N_4179,N_581,N_1608);
nand U4180 (N_4180,N_2155,N_635);
nor U4181 (N_4181,N_875,N_983);
and U4182 (N_4182,N_1475,N_758);
xor U4183 (N_4183,N_496,N_867);
and U4184 (N_4184,N_1061,N_1575);
xor U4185 (N_4185,N_886,N_678);
xor U4186 (N_4186,N_2072,N_1015);
xnor U4187 (N_4187,N_1926,N_2230);
xor U4188 (N_4188,N_1697,N_2010);
or U4189 (N_4189,N_1013,N_2257);
nand U4190 (N_4190,N_2315,N_2489);
nor U4191 (N_4191,N_1496,N_1419);
and U4192 (N_4192,N_521,N_445);
or U4193 (N_4193,N_2058,N_2099);
or U4194 (N_4194,N_1415,N_1009);
xor U4195 (N_4195,N_22,N_1731);
xnor U4196 (N_4196,N_1065,N_2130);
and U4197 (N_4197,N_2374,N_610);
nor U4198 (N_4198,N_1965,N_1911);
or U4199 (N_4199,N_434,N_586);
nand U4200 (N_4200,N_850,N_1642);
nor U4201 (N_4201,N_2006,N_930);
or U4202 (N_4202,N_759,N_885);
nand U4203 (N_4203,N_1219,N_961);
and U4204 (N_4204,N_1201,N_64);
nor U4205 (N_4205,N_1122,N_1624);
and U4206 (N_4206,N_2137,N_1541);
or U4207 (N_4207,N_361,N_16);
and U4208 (N_4208,N_901,N_1914);
or U4209 (N_4209,N_2343,N_2115);
nor U4210 (N_4210,N_648,N_602);
nand U4211 (N_4211,N_2155,N_1822);
xnor U4212 (N_4212,N_1182,N_654);
and U4213 (N_4213,N_1730,N_535);
nand U4214 (N_4214,N_1916,N_887);
or U4215 (N_4215,N_947,N_2187);
nor U4216 (N_4216,N_36,N_1126);
or U4217 (N_4217,N_421,N_2101);
and U4218 (N_4218,N_1215,N_836);
or U4219 (N_4219,N_250,N_1363);
nor U4220 (N_4220,N_1121,N_2217);
nor U4221 (N_4221,N_124,N_2449);
and U4222 (N_4222,N_1403,N_1025);
and U4223 (N_4223,N_182,N_1969);
nand U4224 (N_4224,N_2285,N_1901);
and U4225 (N_4225,N_30,N_282);
or U4226 (N_4226,N_2236,N_190);
or U4227 (N_4227,N_1898,N_1277);
nand U4228 (N_4228,N_924,N_824);
xnor U4229 (N_4229,N_1653,N_1820);
or U4230 (N_4230,N_408,N_434);
and U4231 (N_4231,N_2064,N_465);
or U4232 (N_4232,N_2232,N_1586);
or U4233 (N_4233,N_2272,N_476);
or U4234 (N_4234,N_526,N_812);
nor U4235 (N_4235,N_775,N_2160);
and U4236 (N_4236,N_1100,N_1448);
and U4237 (N_4237,N_2171,N_2158);
nand U4238 (N_4238,N_1666,N_494);
xor U4239 (N_4239,N_546,N_1295);
xor U4240 (N_4240,N_1560,N_1702);
xor U4241 (N_4241,N_2202,N_1210);
nand U4242 (N_4242,N_1647,N_2449);
and U4243 (N_4243,N_910,N_1999);
or U4244 (N_4244,N_1959,N_1515);
nor U4245 (N_4245,N_384,N_480);
and U4246 (N_4246,N_1789,N_428);
nor U4247 (N_4247,N_1127,N_156);
nor U4248 (N_4248,N_300,N_244);
or U4249 (N_4249,N_1678,N_2226);
and U4250 (N_4250,N_1894,N_1138);
and U4251 (N_4251,N_1717,N_221);
nor U4252 (N_4252,N_1698,N_448);
and U4253 (N_4253,N_2046,N_606);
and U4254 (N_4254,N_1159,N_633);
xor U4255 (N_4255,N_1999,N_1692);
nor U4256 (N_4256,N_2253,N_469);
nand U4257 (N_4257,N_1663,N_817);
and U4258 (N_4258,N_762,N_1201);
or U4259 (N_4259,N_769,N_219);
or U4260 (N_4260,N_1379,N_1133);
nor U4261 (N_4261,N_317,N_1796);
nand U4262 (N_4262,N_14,N_366);
nor U4263 (N_4263,N_349,N_345);
and U4264 (N_4264,N_1145,N_985);
and U4265 (N_4265,N_1946,N_1137);
and U4266 (N_4266,N_141,N_287);
xor U4267 (N_4267,N_127,N_2492);
and U4268 (N_4268,N_937,N_439);
or U4269 (N_4269,N_441,N_2369);
nor U4270 (N_4270,N_564,N_1030);
nor U4271 (N_4271,N_473,N_581);
xnor U4272 (N_4272,N_1348,N_1195);
xnor U4273 (N_4273,N_1114,N_524);
or U4274 (N_4274,N_805,N_2396);
xnor U4275 (N_4275,N_1192,N_1271);
nor U4276 (N_4276,N_2473,N_2117);
nand U4277 (N_4277,N_81,N_488);
or U4278 (N_4278,N_1726,N_1409);
nor U4279 (N_4279,N_803,N_1265);
nor U4280 (N_4280,N_450,N_309);
nor U4281 (N_4281,N_327,N_1830);
and U4282 (N_4282,N_36,N_2476);
nand U4283 (N_4283,N_1686,N_829);
xor U4284 (N_4284,N_190,N_1032);
or U4285 (N_4285,N_1090,N_1408);
nor U4286 (N_4286,N_2491,N_146);
and U4287 (N_4287,N_2420,N_2055);
nor U4288 (N_4288,N_124,N_393);
nor U4289 (N_4289,N_1758,N_742);
and U4290 (N_4290,N_357,N_2460);
nor U4291 (N_4291,N_1327,N_153);
or U4292 (N_4292,N_1394,N_2412);
xnor U4293 (N_4293,N_1559,N_865);
and U4294 (N_4294,N_514,N_431);
and U4295 (N_4295,N_1367,N_142);
or U4296 (N_4296,N_238,N_2010);
and U4297 (N_4297,N_1309,N_653);
nand U4298 (N_4298,N_755,N_2098);
nor U4299 (N_4299,N_1983,N_2375);
xor U4300 (N_4300,N_1409,N_742);
and U4301 (N_4301,N_483,N_1916);
and U4302 (N_4302,N_1062,N_632);
xnor U4303 (N_4303,N_521,N_2343);
xor U4304 (N_4304,N_271,N_1578);
or U4305 (N_4305,N_1572,N_625);
xor U4306 (N_4306,N_1008,N_707);
or U4307 (N_4307,N_298,N_1110);
xor U4308 (N_4308,N_1429,N_609);
nand U4309 (N_4309,N_1882,N_256);
nor U4310 (N_4310,N_1676,N_303);
nor U4311 (N_4311,N_1681,N_891);
nand U4312 (N_4312,N_2473,N_476);
and U4313 (N_4313,N_2282,N_1601);
and U4314 (N_4314,N_1121,N_1404);
nor U4315 (N_4315,N_1225,N_904);
or U4316 (N_4316,N_1870,N_1582);
xnor U4317 (N_4317,N_1692,N_1537);
or U4318 (N_4318,N_424,N_2223);
nand U4319 (N_4319,N_1118,N_2488);
and U4320 (N_4320,N_514,N_9);
nor U4321 (N_4321,N_1442,N_485);
nand U4322 (N_4322,N_1550,N_826);
nor U4323 (N_4323,N_218,N_859);
nand U4324 (N_4324,N_1728,N_373);
nor U4325 (N_4325,N_2222,N_1997);
nand U4326 (N_4326,N_1201,N_569);
xnor U4327 (N_4327,N_488,N_361);
xnor U4328 (N_4328,N_954,N_412);
nor U4329 (N_4329,N_760,N_2328);
or U4330 (N_4330,N_1407,N_1889);
nand U4331 (N_4331,N_2170,N_1797);
nor U4332 (N_4332,N_2060,N_627);
and U4333 (N_4333,N_1221,N_2479);
and U4334 (N_4334,N_2396,N_73);
and U4335 (N_4335,N_1322,N_110);
and U4336 (N_4336,N_743,N_1029);
xor U4337 (N_4337,N_1793,N_2409);
nand U4338 (N_4338,N_1486,N_2044);
nor U4339 (N_4339,N_120,N_1370);
xnor U4340 (N_4340,N_551,N_365);
nor U4341 (N_4341,N_2297,N_941);
nor U4342 (N_4342,N_1546,N_1731);
or U4343 (N_4343,N_1267,N_1875);
nor U4344 (N_4344,N_612,N_239);
and U4345 (N_4345,N_1592,N_1983);
or U4346 (N_4346,N_2466,N_1988);
or U4347 (N_4347,N_1291,N_477);
xor U4348 (N_4348,N_1742,N_1355);
xor U4349 (N_4349,N_1543,N_2119);
and U4350 (N_4350,N_2393,N_769);
nor U4351 (N_4351,N_2138,N_325);
nand U4352 (N_4352,N_267,N_457);
or U4353 (N_4353,N_2121,N_94);
and U4354 (N_4354,N_270,N_809);
and U4355 (N_4355,N_2082,N_2251);
and U4356 (N_4356,N_1845,N_1159);
nor U4357 (N_4357,N_89,N_1876);
xnor U4358 (N_4358,N_588,N_721);
nor U4359 (N_4359,N_336,N_922);
nor U4360 (N_4360,N_2033,N_1486);
xnor U4361 (N_4361,N_263,N_562);
nor U4362 (N_4362,N_101,N_918);
or U4363 (N_4363,N_1658,N_2091);
nand U4364 (N_4364,N_952,N_970);
nor U4365 (N_4365,N_1298,N_2327);
nand U4366 (N_4366,N_2309,N_2469);
and U4367 (N_4367,N_2454,N_287);
or U4368 (N_4368,N_787,N_7);
or U4369 (N_4369,N_1182,N_2287);
and U4370 (N_4370,N_960,N_1401);
nor U4371 (N_4371,N_1331,N_1173);
and U4372 (N_4372,N_47,N_78);
or U4373 (N_4373,N_1515,N_2312);
xnor U4374 (N_4374,N_1176,N_849);
and U4375 (N_4375,N_1313,N_742);
xor U4376 (N_4376,N_492,N_484);
and U4377 (N_4377,N_16,N_1648);
or U4378 (N_4378,N_1816,N_2086);
nor U4379 (N_4379,N_1037,N_1321);
nand U4380 (N_4380,N_136,N_652);
and U4381 (N_4381,N_395,N_294);
nor U4382 (N_4382,N_1690,N_628);
nand U4383 (N_4383,N_1425,N_247);
nor U4384 (N_4384,N_1322,N_2485);
nand U4385 (N_4385,N_2490,N_11);
and U4386 (N_4386,N_1742,N_906);
or U4387 (N_4387,N_2226,N_655);
or U4388 (N_4388,N_1250,N_2105);
and U4389 (N_4389,N_1588,N_2421);
nor U4390 (N_4390,N_495,N_922);
or U4391 (N_4391,N_1613,N_480);
or U4392 (N_4392,N_2376,N_1689);
and U4393 (N_4393,N_2377,N_1422);
and U4394 (N_4394,N_1935,N_346);
or U4395 (N_4395,N_2459,N_561);
nor U4396 (N_4396,N_1299,N_1968);
nor U4397 (N_4397,N_1818,N_1232);
xnor U4398 (N_4398,N_951,N_1168);
nor U4399 (N_4399,N_1503,N_2087);
nor U4400 (N_4400,N_1226,N_2196);
xor U4401 (N_4401,N_1818,N_2310);
or U4402 (N_4402,N_569,N_553);
xnor U4403 (N_4403,N_312,N_758);
and U4404 (N_4404,N_448,N_2211);
nand U4405 (N_4405,N_628,N_876);
nand U4406 (N_4406,N_1375,N_2223);
nand U4407 (N_4407,N_58,N_464);
xnor U4408 (N_4408,N_2356,N_1453);
and U4409 (N_4409,N_118,N_1775);
xnor U4410 (N_4410,N_250,N_1498);
nor U4411 (N_4411,N_828,N_603);
xor U4412 (N_4412,N_787,N_2485);
and U4413 (N_4413,N_28,N_238);
xnor U4414 (N_4414,N_2402,N_2);
and U4415 (N_4415,N_2240,N_854);
and U4416 (N_4416,N_288,N_1292);
nor U4417 (N_4417,N_975,N_2313);
xnor U4418 (N_4418,N_1552,N_1116);
nand U4419 (N_4419,N_1548,N_1425);
nor U4420 (N_4420,N_2120,N_511);
and U4421 (N_4421,N_1217,N_167);
nand U4422 (N_4422,N_892,N_1199);
nand U4423 (N_4423,N_476,N_748);
xnor U4424 (N_4424,N_1575,N_1659);
and U4425 (N_4425,N_1448,N_1883);
nor U4426 (N_4426,N_2418,N_1529);
or U4427 (N_4427,N_2297,N_1448);
nor U4428 (N_4428,N_686,N_1839);
or U4429 (N_4429,N_2482,N_1202);
and U4430 (N_4430,N_1385,N_1644);
and U4431 (N_4431,N_1374,N_987);
and U4432 (N_4432,N_238,N_2233);
and U4433 (N_4433,N_790,N_1480);
or U4434 (N_4434,N_139,N_1494);
nor U4435 (N_4435,N_1382,N_648);
nand U4436 (N_4436,N_848,N_205);
nor U4437 (N_4437,N_230,N_555);
and U4438 (N_4438,N_1759,N_1317);
and U4439 (N_4439,N_1000,N_312);
xnor U4440 (N_4440,N_1299,N_1653);
nor U4441 (N_4441,N_1154,N_970);
xor U4442 (N_4442,N_2080,N_1231);
nand U4443 (N_4443,N_1029,N_1513);
xnor U4444 (N_4444,N_261,N_1344);
and U4445 (N_4445,N_1353,N_528);
nor U4446 (N_4446,N_349,N_1373);
nor U4447 (N_4447,N_2447,N_1256);
nand U4448 (N_4448,N_1428,N_1268);
xnor U4449 (N_4449,N_809,N_1589);
or U4450 (N_4450,N_1662,N_1679);
nand U4451 (N_4451,N_2138,N_1999);
or U4452 (N_4452,N_1835,N_1345);
nand U4453 (N_4453,N_2403,N_226);
and U4454 (N_4454,N_59,N_1483);
nand U4455 (N_4455,N_1881,N_2456);
or U4456 (N_4456,N_1188,N_2400);
nand U4457 (N_4457,N_14,N_452);
nand U4458 (N_4458,N_1952,N_83);
nor U4459 (N_4459,N_207,N_41);
and U4460 (N_4460,N_92,N_519);
xnor U4461 (N_4461,N_497,N_2177);
xor U4462 (N_4462,N_2119,N_2428);
and U4463 (N_4463,N_600,N_1119);
xor U4464 (N_4464,N_1965,N_1359);
xor U4465 (N_4465,N_1085,N_27);
nand U4466 (N_4466,N_66,N_1581);
nand U4467 (N_4467,N_1380,N_1016);
nor U4468 (N_4468,N_87,N_1008);
xor U4469 (N_4469,N_2003,N_661);
and U4470 (N_4470,N_2038,N_801);
nand U4471 (N_4471,N_2100,N_1271);
and U4472 (N_4472,N_219,N_1020);
nor U4473 (N_4473,N_1821,N_1348);
and U4474 (N_4474,N_1812,N_1947);
and U4475 (N_4475,N_1501,N_2262);
nand U4476 (N_4476,N_426,N_536);
nor U4477 (N_4477,N_720,N_646);
or U4478 (N_4478,N_1361,N_2181);
or U4479 (N_4479,N_1858,N_1123);
or U4480 (N_4480,N_2195,N_2481);
or U4481 (N_4481,N_2348,N_54);
nand U4482 (N_4482,N_2213,N_1427);
nor U4483 (N_4483,N_1403,N_218);
and U4484 (N_4484,N_395,N_1102);
or U4485 (N_4485,N_2373,N_1518);
xor U4486 (N_4486,N_1526,N_426);
xor U4487 (N_4487,N_1666,N_2329);
and U4488 (N_4488,N_489,N_49);
nand U4489 (N_4489,N_641,N_1406);
or U4490 (N_4490,N_2089,N_2117);
nor U4491 (N_4491,N_82,N_151);
or U4492 (N_4492,N_257,N_1088);
and U4493 (N_4493,N_2265,N_2260);
nor U4494 (N_4494,N_531,N_65);
and U4495 (N_4495,N_1788,N_1834);
and U4496 (N_4496,N_1172,N_1694);
nand U4497 (N_4497,N_674,N_76);
nor U4498 (N_4498,N_1346,N_1420);
nand U4499 (N_4499,N_2009,N_2120);
nor U4500 (N_4500,N_1643,N_429);
or U4501 (N_4501,N_1646,N_580);
xor U4502 (N_4502,N_57,N_934);
or U4503 (N_4503,N_1413,N_1384);
xor U4504 (N_4504,N_422,N_176);
and U4505 (N_4505,N_1452,N_37);
or U4506 (N_4506,N_318,N_2423);
and U4507 (N_4507,N_1094,N_1236);
or U4508 (N_4508,N_47,N_1499);
xor U4509 (N_4509,N_1554,N_2450);
or U4510 (N_4510,N_871,N_344);
or U4511 (N_4511,N_1216,N_1605);
or U4512 (N_4512,N_1789,N_1181);
nand U4513 (N_4513,N_2149,N_2336);
nor U4514 (N_4514,N_380,N_1092);
nand U4515 (N_4515,N_863,N_553);
nor U4516 (N_4516,N_37,N_996);
and U4517 (N_4517,N_2179,N_454);
nor U4518 (N_4518,N_2232,N_759);
and U4519 (N_4519,N_1721,N_1634);
or U4520 (N_4520,N_561,N_2064);
nor U4521 (N_4521,N_552,N_936);
xnor U4522 (N_4522,N_1642,N_2320);
xnor U4523 (N_4523,N_1382,N_588);
xnor U4524 (N_4524,N_767,N_856);
nor U4525 (N_4525,N_2386,N_2224);
nor U4526 (N_4526,N_732,N_365);
nand U4527 (N_4527,N_1708,N_2223);
or U4528 (N_4528,N_1563,N_1269);
nor U4529 (N_4529,N_1195,N_1853);
and U4530 (N_4530,N_2426,N_409);
or U4531 (N_4531,N_1649,N_738);
and U4532 (N_4532,N_1461,N_2404);
and U4533 (N_4533,N_1272,N_2008);
nor U4534 (N_4534,N_1544,N_2457);
xnor U4535 (N_4535,N_1773,N_1191);
or U4536 (N_4536,N_1067,N_2418);
xnor U4537 (N_4537,N_1255,N_566);
nand U4538 (N_4538,N_636,N_1054);
nand U4539 (N_4539,N_1712,N_766);
and U4540 (N_4540,N_362,N_1092);
or U4541 (N_4541,N_727,N_2084);
nand U4542 (N_4542,N_233,N_993);
or U4543 (N_4543,N_2444,N_1244);
nor U4544 (N_4544,N_2478,N_636);
and U4545 (N_4545,N_2370,N_1718);
nor U4546 (N_4546,N_794,N_48);
and U4547 (N_4547,N_49,N_1207);
xnor U4548 (N_4548,N_1697,N_2346);
xor U4549 (N_4549,N_535,N_1979);
or U4550 (N_4550,N_2089,N_1779);
or U4551 (N_4551,N_1344,N_1066);
nor U4552 (N_4552,N_703,N_1620);
and U4553 (N_4553,N_109,N_1432);
nor U4554 (N_4554,N_1877,N_2367);
and U4555 (N_4555,N_2368,N_1235);
xor U4556 (N_4556,N_1073,N_892);
and U4557 (N_4557,N_10,N_1551);
nor U4558 (N_4558,N_1719,N_1491);
nor U4559 (N_4559,N_2449,N_1404);
nor U4560 (N_4560,N_211,N_624);
nor U4561 (N_4561,N_289,N_1912);
and U4562 (N_4562,N_1346,N_1408);
xor U4563 (N_4563,N_1139,N_2336);
nand U4564 (N_4564,N_1648,N_2290);
xor U4565 (N_4565,N_576,N_2387);
nor U4566 (N_4566,N_2271,N_1446);
nand U4567 (N_4567,N_1061,N_2416);
or U4568 (N_4568,N_384,N_2307);
xor U4569 (N_4569,N_2279,N_717);
nor U4570 (N_4570,N_2214,N_850);
nor U4571 (N_4571,N_2180,N_41);
xnor U4572 (N_4572,N_1311,N_1403);
xnor U4573 (N_4573,N_554,N_1820);
or U4574 (N_4574,N_950,N_190);
xnor U4575 (N_4575,N_933,N_1128);
nand U4576 (N_4576,N_88,N_1622);
and U4577 (N_4577,N_250,N_1866);
nand U4578 (N_4578,N_431,N_452);
nor U4579 (N_4579,N_1138,N_2453);
nand U4580 (N_4580,N_1983,N_82);
xor U4581 (N_4581,N_703,N_1261);
nand U4582 (N_4582,N_2224,N_871);
nor U4583 (N_4583,N_1701,N_1433);
and U4584 (N_4584,N_756,N_331);
nor U4585 (N_4585,N_596,N_805);
nor U4586 (N_4586,N_1261,N_394);
nor U4587 (N_4587,N_1902,N_1128);
and U4588 (N_4588,N_1812,N_2064);
nand U4589 (N_4589,N_1853,N_241);
or U4590 (N_4590,N_692,N_1770);
nand U4591 (N_4591,N_1639,N_2497);
and U4592 (N_4592,N_2205,N_2358);
nor U4593 (N_4593,N_1005,N_2345);
nand U4594 (N_4594,N_509,N_1846);
xor U4595 (N_4595,N_520,N_959);
or U4596 (N_4596,N_896,N_1688);
nor U4597 (N_4597,N_212,N_2237);
nor U4598 (N_4598,N_126,N_1784);
nor U4599 (N_4599,N_414,N_969);
xnor U4600 (N_4600,N_1383,N_1471);
and U4601 (N_4601,N_1452,N_427);
nor U4602 (N_4602,N_1389,N_1244);
nand U4603 (N_4603,N_1349,N_1450);
and U4604 (N_4604,N_108,N_31);
or U4605 (N_4605,N_1665,N_648);
or U4606 (N_4606,N_1649,N_300);
or U4607 (N_4607,N_1770,N_2404);
nor U4608 (N_4608,N_2444,N_441);
xnor U4609 (N_4609,N_1141,N_1470);
xor U4610 (N_4610,N_179,N_2313);
xnor U4611 (N_4611,N_1162,N_1990);
nand U4612 (N_4612,N_1006,N_255);
nor U4613 (N_4613,N_1310,N_947);
nand U4614 (N_4614,N_1579,N_911);
or U4615 (N_4615,N_943,N_1428);
nor U4616 (N_4616,N_951,N_1777);
nand U4617 (N_4617,N_273,N_2123);
nand U4618 (N_4618,N_1461,N_1312);
nor U4619 (N_4619,N_1726,N_517);
xor U4620 (N_4620,N_722,N_2397);
nand U4621 (N_4621,N_772,N_532);
nor U4622 (N_4622,N_1676,N_1833);
and U4623 (N_4623,N_2099,N_583);
xor U4624 (N_4624,N_1882,N_1649);
and U4625 (N_4625,N_178,N_1398);
and U4626 (N_4626,N_2491,N_2318);
or U4627 (N_4627,N_1294,N_2360);
nand U4628 (N_4628,N_1280,N_801);
and U4629 (N_4629,N_2233,N_263);
nand U4630 (N_4630,N_1166,N_849);
and U4631 (N_4631,N_187,N_49);
nand U4632 (N_4632,N_147,N_1188);
and U4633 (N_4633,N_1669,N_2272);
or U4634 (N_4634,N_575,N_2489);
and U4635 (N_4635,N_908,N_293);
nand U4636 (N_4636,N_190,N_1681);
nand U4637 (N_4637,N_1722,N_1047);
and U4638 (N_4638,N_39,N_326);
xor U4639 (N_4639,N_840,N_710);
and U4640 (N_4640,N_997,N_1890);
xor U4641 (N_4641,N_1489,N_1537);
nand U4642 (N_4642,N_2070,N_242);
or U4643 (N_4643,N_1309,N_1994);
nand U4644 (N_4644,N_1546,N_740);
nand U4645 (N_4645,N_1412,N_91);
nand U4646 (N_4646,N_1380,N_112);
nand U4647 (N_4647,N_559,N_820);
nor U4648 (N_4648,N_152,N_1102);
nand U4649 (N_4649,N_121,N_189);
or U4650 (N_4650,N_590,N_2412);
or U4651 (N_4651,N_1882,N_1254);
nor U4652 (N_4652,N_445,N_1793);
and U4653 (N_4653,N_1790,N_724);
or U4654 (N_4654,N_768,N_1705);
and U4655 (N_4655,N_149,N_1812);
and U4656 (N_4656,N_1824,N_351);
or U4657 (N_4657,N_890,N_1364);
xnor U4658 (N_4658,N_1672,N_433);
and U4659 (N_4659,N_1900,N_360);
and U4660 (N_4660,N_788,N_1343);
nor U4661 (N_4661,N_777,N_1837);
nand U4662 (N_4662,N_2219,N_1537);
xnor U4663 (N_4663,N_143,N_597);
and U4664 (N_4664,N_2252,N_299);
nor U4665 (N_4665,N_631,N_1897);
or U4666 (N_4666,N_687,N_702);
nor U4667 (N_4667,N_588,N_1810);
and U4668 (N_4668,N_1713,N_1968);
nand U4669 (N_4669,N_658,N_2068);
nor U4670 (N_4670,N_448,N_2128);
nor U4671 (N_4671,N_2363,N_176);
nand U4672 (N_4672,N_903,N_1511);
or U4673 (N_4673,N_64,N_1473);
xnor U4674 (N_4674,N_1653,N_478);
or U4675 (N_4675,N_1981,N_1502);
xor U4676 (N_4676,N_1945,N_1775);
xor U4677 (N_4677,N_1162,N_1684);
xor U4678 (N_4678,N_167,N_2440);
xnor U4679 (N_4679,N_981,N_1416);
and U4680 (N_4680,N_1665,N_1716);
and U4681 (N_4681,N_871,N_2349);
nor U4682 (N_4682,N_23,N_1755);
xor U4683 (N_4683,N_1932,N_1161);
nand U4684 (N_4684,N_483,N_1611);
and U4685 (N_4685,N_1934,N_2341);
and U4686 (N_4686,N_2125,N_1906);
xnor U4687 (N_4687,N_1863,N_1913);
or U4688 (N_4688,N_452,N_1676);
nor U4689 (N_4689,N_29,N_1870);
or U4690 (N_4690,N_1875,N_52);
or U4691 (N_4691,N_487,N_1412);
or U4692 (N_4692,N_1479,N_2085);
nand U4693 (N_4693,N_1655,N_409);
and U4694 (N_4694,N_291,N_427);
xor U4695 (N_4695,N_966,N_354);
or U4696 (N_4696,N_1450,N_402);
nand U4697 (N_4697,N_921,N_2063);
and U4698 (N_4698,N_1472,N_2315);
or U4699 (N_4699,N_1304,N_481);
nand U4700 (N_4700,N_2238,N_1625);
xor U4701 (N_4701,N_2237,N_1915);
nor U4702 (N_4702,N_2175,N_2227);
nor U4703 (N_4703,N_2468,N_2434);
or U4704 (N_4704,N_2207,N_1795);
nand U4705 (N_4705,N_1134,N_1866);
and U4706 (N_4706,N_1278,N_1153);
nor U4707 (N_4707,N_797,N_2266);
and U4708 (N_4708,N_958,N_388);
and U4709 (N_4709,N_239,N_1632);
xor U4710 (N_4710,N_638,N_742);
and U4711 (N_4711,N_4,N_165);
and U4712 (N_4712,N_1957,N_2340);
nor U4713 (N_4713,N_1217,N_292);
nand U4714 (N_4714,N_2235,N_1996);
or U4715 (N_4715,N_265,N_1246);
nand U4716 (N_4716,N_2275,N_218);
or U4717 (N_4717,N_2251,N_2020);
nor U4718 (N_4718,N_604,N_1860);
and U4719 (N_4719,N_1435,N_914);
and U4720 (N_4720,N_1109,N_1755);
xnor U4721 (N_4721,N_1967,N_959);
xnor U4722 (N_4722,N_2023,N_1815);
xor U4723 (N_4723,N_218,N_1935);
or U4724 (N_4724,N_1530,N_1658);
or U4725 (N_4725,N_841,N_2377);
xor U4726 (N_4726,N_1050,N_792);
nand U4727 (N_4727,N_839,N_1987);
nor U4728 (N_4728,N_1505,N_1085);
xor U4729 (N_4729,N_1304,N_1651);
nor U4730 (N_4730,N_214,N_1549);
nor U4731 (N_4731,N_740,N_1234);
nand U4732 (N_4732,N_2108,N_2406);
and U4733 (N_4733,N_805,N_1655);
xnor U4734 (N_4734,N_408,N_2347);
xnor U4735 (N_4735,N_1598,N_2167);
nor U4736 (N_4736,N_109,N_877);
and U4737 (N_4737,N_1623,N_874);
xor U4738 (N_4738,N_2417,N_1992);
or U4739 (N_4739,N_519,N_2227);
nand U4740 (N_4740,N_348,N_820);
xnor U4741 (N_4741,N_2308,N_1279);
nor U4742 (N_4742,N_2055,N_1531);
nor U4743 (N_4743,N_419,N_1538);
nand U4744 (N_4744,N_2477,N_1613);
xor U4745 (N_4745,N_2016,N_1556);
or U4746 (N_4746,N_2023,N_2413);
nand U4747 (N_4747,N_1597,N_562);
xnor U4748 (N_4748,N_841,N_302);
nor U4749 (N_4749,N_1502,N_1315);
xor U4750 (N_4750,N_378,N_2023);
xor U4751 (N_4751,N_2280,N_1589);
nor U4752 (N_4752,N_493,N_1515);
and U4753 (N_4753,N_86,N_408);
xor U4754 (N_4754,N_54,N_1879);
or U4755 (N_4755,N_649,N_1360);
and U4756 (N_4756,N_1679,N_2260);
and U4757 (N_4757,N_1646,N_2294);
and U4758 (N_4758,N_360,N_2215);
nand U4759 (N_4759,N_2066,N_1895);
nand U4760 (N_4760,N_649,N_2224);
nor U4761 (N_4761,N_163,N_2210);
xor U4762 (N_4762,N_2007,N_584);
xor U4763 (N_4763,N_2154,N_2279);
nor U4764 (N_4764,N_502,N_590);
and U4765 (N_4765,N_2490,N_1156);
nor U4766 (N_4766,N_1305,N_1222);
or U4767 (N_4767,N_762,N_2457);
xnor U4768 (N_4768,N_487,N_1011);
nor U4769 (N_4769,N_1670,N_2135);
and U4770 (N_4770,N_1554,N_571);
xor U4771 (N_4771,N_785,N_2095);
xnor U4772 (N_4772,N_1241,N_1834);
nand U4773 (N_4773,N_1871,N_2136);
and U4774 (N_4774,N_1853,N_1271);
nand U4775 (N_4775,N_479,N_550);
nand U4776 (N_4776,N_1059,N_1642);
nor U4777 (N_4777,N_1323,N_2064);
nand U4778 (N_4778,N_1540,N_2471);
xnor U4779 (N_4779,N_1469,N_893);
or U4780 (N_4780,N_1291,N_1075);
xor U4781 (N_4781,N_1816,N_2038);
or U4782 (N_4782,N_842,N_365);
or U4783 (N_4783,N_241,N_1536);
nor U4784 (N_4784,N_1091,N_1839);
nand U4785 (N_4785,N_582,N_1165);
nor U4786 (N_4786,N_2372,N_771);
nor U4787 (N_4787,N_190,N_1335);
and U4788 (N_4788,N_1502,N_1516);
xor U4789 (N_4789,N_2385,N_1348);
nor U4790 (N_4790,N_260,N_94);
nand U4791 (N_4791,N_650,N_122);
or U4792 (N_4792,N_1978,N_1473);
xor U4793 (N_4793,N_208,N_1047);
xnor U4794 (N_4794,N_1034,N_962);
xor U4795 (N_4795,N_1923,N_2147);
nand U4796 (N_4796,N_1835,N_1390);
nand U4797 (N_4797,N_421,N_1621);
nand U4798 (N_4798,N_584,N_467);
nand U4799 (N_4799,N_1567,N_2260);
xnor U4800 (N_4800,N_267,N_302);
nor U4801 (N_4801,N_1550,N_1549);
nor U4802 (N_4802,N_159,N_2082);
nor U4803 (N_4803,N_704,N_2219);
nand U4804 (N_4804,N_1382,N_2385);
xor U4805 (N_4805,N_1025,N_523);
and U4806 (N_4806,N_1140,N_406);
or U4807 (N_4807,N_1308,N_360);
or U4808 (N_4808,N_2246,N_2043);
and U4809 (N_4809,N_1752,N_497);
and U4810 (N_4810,N_1379,N_1715);
nor U4811 (N_4811,N_1556,N_1701);
xnor U4812 (N_4812,N_910,N_2000);
or U4813 (N_4813,N_1900,N_303);
xor U4814 (N_4814,N_1217,N_2099);
or U4815 (N_4815,N_685,N_141);
nor U4816 (N_4816,N_1152,N_157);
or U4817 (N_4817,N_1831,N_1749);
and U4818 (N_4818,N_1491,N_699);
xnor U4819 (N_4819,N_994,N_499);
nor U4820 (N_4820,N_1487,N_1879);
xor U4821 (N_4821,N_2238,N_2179);
xor U4822 (N_4822,N_2025,N_668);
nor U4823 (N_4823,N_1336,N_1680);
nor U4824 (N_4824,N_2343,N_2200);
xnor U4825 (N_4825,N_2295,N_221);
nand U4826 (N_4826,N_721,N_1995);
nand U4827 (N_4827,N_274,N_1418);
and U4828 (N_4828,N_1804,N_1643);
xor U4829 (N_4829,N_385,N_1626);
nor U4830 (N_4830,N_1606,N_2273);
nor U4831 (N_4831,N_2488,N_883);
nand U4832 (N_4832,N_1021,N_598);
nand U4833 (N_4833,N_774,N_63);
and U4834 (N_4834,N_1268,N_1767);
nor U4835 (N_4835,N_218,N_2212);
or U4836 (N_4836,N_216,N_2253);
and U4837 (N_4837,N_1788,N_60);
or U4838 (N_4838,N_1899,N_1505);
xor U4839 (N_4839,N_709,N_893);
xor U4840 (N_4840,N_1335,N_923);
xor U4841 (N_4841,N_184,N_1998);
nand U4842 (N_4842,N_1345,N_1351);
nor U4843 (N_4843,N_189,N_1857);
and U4844 (N_4844,N_2352,N_2345);
or U4845 (N_4845,N_57,N_1901);
and U4846 (N_4846,N_258,N_2102);
nor U4847 (N_4847,N_1591,N_1018);
and U4848 (N_4848,N_1179,N_257);
xor U4849 (N_4849,N_1395,N_2385);
nor U4850 (N_4850,N_2237,N_1615);
or U4851 (N_4851,N_2289,N_1568);
or U4852 (N_4852,N_1278,N_2264);
nand U4853 (N_4853,N_547,N_1096);
or U4854 (N_4854,N_1886,N_1673);
or U4855 (N_4855,N_2315,N_1228);
or U4856 (N_4856,N_2199,N_904);
xor U4857 (N_4857,N_1708,N_404);
xor U4858 (N_4858,N_2014,N_843);
or U4859 (N_4859,N_2387,N_1499);
nor U4860 (N_4860,N_1683,N_1029);
nor U4861 (N_4861,N_1395,N_1545);
xnor U4862 (N_4862,N_1459,N_248);
and U4863 (N_4863,N_326,N_2263);
or U4864 (N_4864,N_2357,N_2380);
or U4865 (N_4865,N_872,N_906);
xnor U4866 (N_4866,N_29,N_98);
xnor U4867 (N_4867,N_896,N_1970);
or U4868 (N_4868,N_540,N_256);
nor U4869 (N_4869,N_367,N_1074);
xor U4870 (N_4870,N_451,N_2002);
xor U4871 (N_4871,N_2097,N_776);
and U4872 (N_4872,N_533,N_1539);
nor U4873 (N_4873,N_1457,N_487);
or U4874 (N_4874,N_1502,N_2303);
or U4875 (N_4875,N_2016,N_130);
and U4876 (N_4876,N_2149,N_103);
or U4877 (N_4877,N_1987,N_2273);
and U4878 (N_4878,N_915,N_592);
nand U4879 (N_4879,N_1824,N_1715);
or U4880 (N_4880,N_1320,N_640);
and U4881 (N_4881,N_298,N_790);
or U4882 (N_4882,N_1616,N_1543);
nor U4883 (N_4883,N_1979,N_1064);
nor U4884 (N_4884,N_1435,N_1355);
and U4885 (N_4885,N_1252,N_874);
and U4886 (N_4886,N_1162,N_1857);
nor U4887 (N_4887,N_1253,N_184);
or U4888 (N_4888,N_852,N_245);
nor U4889 (N_4889,N_1206,N_1995);
nand U4890 (N_4890,N_1859,N_169);
xnor U4891 (N_4891,N_240,N_882);
nand U4892 (N_4892,N_773,N_2105);
and U4893 (N_4893,N_987,N_2246);
nor U4894 (N_4894,N_299,N_847);
and U4895 (N_4895,N_1687,N_1168);
or U4896 (N_4896,N_2182,N_2058);
and U4897 (N_4897,N_375,N_1830);
nand U4898 (N_4898,N_2408,N_823);
xnor U4899 (N_4899,N_297,N_1256);
nor U4900 (N_4900,N_162,N_1531);
xnor U4901 (N_4901,N_2303,N_1155);
or U4902 (N_4902,N_749,N_1607);
and U4903 (N_4903,N_1889,N_69);
xor U4904 (N_4904,N_1241,N_2433);
and U4905 (N_4905,N_1088,N_285);
nand U4906 (N_4906,N_345,N_1593);
xor U4907 (N_4907,N_1847,N_1959);
nor U4908 (N_4908,N_1981,N_1180);
nor U4909 (N_4909,N_1272,N_111);
or U4910 (N_4910,N_2112,N_482);
or U4911 (N_4911,N_2428,N_861);
and U4912 (N_4912,N_2411,N_1619);
nor U4913 (N_4913,N_1848,N_1715);
or U4914 (N_4914,N_149,N_122);
xnor U4915 (N_4915,N_2380,N_2155);
or U4916 (N_4916,N_582,N_2376);
and U4917 (N_4917,N_1237,N_1418);
and U4918 (N_4918,N_420,N_11);
xor U4919 (N_4919,N_230,N_1045);
and U4920 (N_4920,N_1355,N_647);
nand U4921 (N_4921,N_2149,N_425);
or U4922 (N_4922,N_888,N_461);
nor U4923 (N_4923,N_2401,N_2466);
or U4924 (N_4924,N_804,N_1779);
or U4925 (N_4925,N_2083,N_1116);
nor U4926 (N_4926,N_286,N_2433);
or U4927 (N_4927,N_879,N_63);
xnor U4928 (N_4928,N_185,N_182);
xor U4929 (N_4929,N_292,N_2298);
xor U4930 (N_4930,N_2385,N_771);
xor U4931 (N_4931,N_107,N_342);
nand U4932 (N_4932,N_826,N_1994);
xor U4933 (N_4933,N_1245,N_2392);
nand U4934 (N_4934,N_2497,N_963);
and U4935 (N_4935,N_1885,N_1205);
nor U4936 (N_4936,N_907,N_583);
xor U4937 (N_4937,N_1337,N_805);
nand U4938 (N_4938,N_2300,N_750);
nor U4939 (N_4939,N_1,N_2085);
nand U4940 (N_4940,N_541,N_602);
xnor U4941 (N_4941,N_1065,N_2406);
and U4942 (N_4942,N_2082,N_1461);
xnor U4943 (N_4943,N_2476,N_1955);
and U4944 (N_4944,N_2087,N_444);
nor U4945 (N_4945,N_1389,N_36);
nor U4946 (N_4946,N_1225,N_1470);
and U4947 (N_4947,N_622,N_2086);
nor U4948 (N_4948,N_2460,N_223);
nand U4949 (N_4949,N_683,N_1123);
xor U4950 (N_4950,N_59,N_781);
or U4951 (N_4951,N_869,N_2274);
or U4952 (N_4952,N_2393,N_762);
nor U4953 (N_4953,N_1224,N_114);
and U4954 (N_4954,N_1101,N_42);
nand U4955 (N_4955,N_362,N_1698);
nor U4956 (N_4956,N_2271,N_897);
or U4957 (N_4957,N_144,N_1950);
xor U4958 (N_4958,N_1892,N_1101);
nand U4959 (N_4959,N_2060,N_1897);
nor U4960 (N_4960,N_1771,N_1239);
and U4961 (N_4961,N_473,N_1878);
xor U4962 (N_4962,N_1538,N_2270);
and U4963 (N_4963,N_1903,N_1946);
nor U4964 (N_4964,N_1825,N_172);
xnor U4965 (N_4965,N_2216,N_1477);
or U4966 (N_4966,N_1637,N_0);
and U4967 (N_4967,N_2374,N_2381);
xnor U4968 (N_4968,N_2238,N_890);
or U4969 (N_4969,N_1788,N_2489);
nor U4970 (N_4970,N_435,N_291);
and U4971 (N_4971,N_1393,N_1047);
nor U4972 (N_4972,N_1009,N_2363);
and U4973 (N_4973,N_1694,N_1678);
and U4974 (N_4974,N_1384,N_95);
nand U4975 (N_4975,N_2195,N_1129);
nand U4976 (N_4976,N_942,N_1224);
nand U4977 (N_4977,N_1136,N_1823);
and U4978 (N_4978,N_1420,N_181);
nor U4979 (N_4979,N_1111,N_1893);
and U4980 (N_4980,N_1655,N_2240);
nand U4981 (N_4981,N_480,N_2154);
xnor U4982 (N_4982,N_1129,N_3);
or U4983 (N_4983,N_1752,N_514);
xnor U4984 (N_4984,N_244,N_726);
nor U4985 (N_4985,N_618,N_2488);
nand U4986 (N_4986,N_1655,N_1609);
and U4987 (N_4987,N_1806,N_2429);
and U4988 (N_4988,N_399,N_1555);
xnor U4989 (N_4989,N_2053,N_1336);
and U4990 (N_4990,N_1259,N_2444);
and U4991 (N_4991,N_1163,N_999);
xnor U4992 (N_4992,N_30,N_304);
xor U4993 (N_4993,N_327,N_2263);
and U4994 (N_4994,N_1783,N_553);
nor U4995 (N_4995,N_1173,N_1925);
xnor U4996 (N_4996,N_1283,N_2037);
xor U4997 (N_4997,N_1283,N_659);
and U4998 (N_4998,N_1111,N_874);
or U4999 (N_4999,N_1658,N_1389);
nor U5000 (N_5000,N_4711,N_2631);
nor U5001 (N_5001,N_2868,N_2582);
xor U5002 (N_5002,N_4354,N_4168);
nor U5003 (N_5003,N_3877,N_3208);
xor U5004 (N_5004,N_2802,N_4413);
or U5005 (N_5005,N_4063,N_4167);
nand U5006 (N_5006,N_3021,N_2745);
or U5007 (N_5007,N_4608,N_4991);
and U5008 (N_5008,N_3794,N_3912);
and U5009 (N_5009,N_4118,N_4443);
nand U5010 (N_5010,N_3569,N_3029);
nor U5011 (N_5011,N_3823,N_3496);
and U5012 (N_5012,N_4427,N_3750);
or U5013 (N_5013,N_4982,N_2981);
nor U5014 (N_5014,N_4646,N_3350);
or U5015 (N_5015,N_4075,N_4417);
nor U5016 (N_5016,N_4231,N_2939);
and U5017 (N_5017,N_3653,N_4130);
xor U5018 (N_5018,N_4154,N_3742);
or U5019 (N_5019,N_4432,N_3722);
xor U5020 (N_5020,N_3594,N_4885);
xnor U5021 (N_5021,N_3515,N_3634);
or U5022 (N_5022,N_2852,N_2533);
nand U5023 (N_5023,N_3774,N_2504);
nand U5024 (N_5024,N_3777,N_4724);
and U5025 (N_5025,N_3534,N_3730);
and U5026 (N_5026,N_3733,N_3150);
or U5027 (N_5027,N_4198,N_4401);
nand U5028 (N_5028,N_2508,N_4203);
xor U5029 (N_5029,N_4103,N_3367);
or U5030 (N_5030,N_3511,N_2727);
xnor U5031 (N_5031,N_4833,N_3537);
xnor U5032 (N_5032,N_3163,N_2874);
nor U5033 (N_5033,N_3577,N_4993);
or U5034 (N_5034,N_4683,N_3828);
nor U5035 (N_5035,N_3861,N_2731);
or U5036 (N_5036,N_4852,N_4194);
nor U5037 (N_5037,N_2865,N_3455);
nand U5038 (N_5038,N_4364,N_3476);
nor U5039 (N_5039,N_3636,N_3749);
xnor U5040 (N_5040,N_2553,N_4738);
xor U5041 (N_5041,N_4291,N_3473);
nor U5042 (N_5042,N_2902,N_4987);
and U5043 (N_5043,N_4763,N_4326);
xnor U5044 (N_5044,N_3919,N_3528);
and U5045 (N_5045,N_3045,N_2552);
xor U5046 (N_5046,N_4623,N_2517);
and U5047 (N_5047,N_2624,N_3746);
nor U5048 (N_5048,N_3082,N_4228);
and U5049 (N_5049,N_2707,N_2664);
nand U5050 (N_5050,N_3505,N_4193);
or U5051 (N_5051,N_3372,N_3624);
xnor U5052 (N_5052,N_2503,N_2895);
and U5053 (N_5053,N_4361,N_2539);
nand U5054 (N_5054,N_3761,N_3425);
nand U5055 (N_5055,N_3457,N_4334);
nor U5056 (N_5056,N_4640,N_4458);
xnor U5057 (N_5057,N_4902,N_2914);
nand U5058 (N_5058,N_3259,N_4003);
xor U5059 (N_5059,N_3380,N_3377);
and U5060 (N_5060,N_3701,N_2775);
xnor U5061 (N_5061,N_4406,N_3504);
or U5062 (N_5062,N_4642,N_2773);
nand U5063 (N_5063,N_4282,N_4524);
nor U5064 (N_5064,N_3519,N_3024);
nor U5065 (N_5065,N_3487,N_3293);
xor U5066 (N_5066,N_4855,N_3226);
or U5067 (N_5067,N_4884,N_2521);
nor U5068 (N_5068,N_3558,N_4302);
or U5069 (N_5069,N_4058,N_4355);
xnor U5070 (N_5070,N_3379,N_3681);
nor U5071 (N_5071,N_4025,N_4582);
nor U5072 (N_5072,N_4834,N_3939);
and U5073 (N_5073,N_4077,N_4467);
nor U5074 (N_5074,N_4150,N_4593);
or U5075 (N_5075,N_2938,N_2755);
and U5076 (N_5076,N_3429,N_2659);
or U5077 (N_5077,N_2655,N_4717);
nor U5078 (N_5078,N_2681,N_2764);
xnor U5079 (N_5079,N_3878,N_2821);
and U5080 (N_5080,N_3467,N_2602);
and U5081 (N_5081,N_4470,N_2563);
nor U5082 (N_5082,N_2726,N_3518);
nor U5083 (N_5083,N_2728,N_2722);
xor U5084 (N_5084,N_3093,N_2928);
nand U5085 (N_5085,N_3724,N_3098);
nand U5086 (N_5086,N_4370,N_4612);
and U5087 (N_5087,N_2592,N_4534);
or U5088 (N_5088,N_3755,N_3116);
nor U5089 (N_5089,N_4903,N_3371);
nor U5090 (N_5090,N_3507,N_3885);
nor U5091 (N_5091,N_4638,N_3644);
xnor U5092 (N_5092,N_2875,N_4658);
nand U5093 (N_5093,N_2640,N_3227);
or U5094 (N_5094,N_3531,N_4665);
nor U5095 (N_5095,N_4229,N_4791);
xnor U5096 (N_5096,N_2679,N_3203);
nand U5097 (N_5097,N_3073,N_3276);
nor U5098 (N_5098,N_4125,N_4986);
or U5099 (N_5099,N_3946,N_3005);
nor U5100 (N_5100,N_3252,N_3584);
nand U5101 (N_5101,N_3941,N_4343);
and U5102 (N_5102,N_2639,N_3545);
nor U5103 (N_5103,N_4807,N_2823);
xor U5104 (N_5104,N_4006,N_4924);
nand U5105 (N_5105,N_2693,N_3326);
and U5106 (N_5106,N_2965,N_4021);
and U5107 (N_5107,N_3810,N_4525);
and U5108 (N_5108,N_3028,N_3396);
and U5109 (N_5109,N_4615,N_2729);
nand U5110 (N_5110,N_4328,N_3205);
or U5111 (N_5111,N_3143,N_3931);
nor U5112 (N_5112,N_3542,N_3744);
nand U5113 (N_5113,N_4731,N_2564);
and U5114 (N_5114,N_3954,N_4743);
nor U5115 (N_5115,N_4165,N_2571);
or U5116 (N_5116,N_4286,N_2557);
xnor U5117 (N_5117,N_4671,N_4105);
nand U5118 (N_5118,N_3443,N_2923);
nand U5119 (N_5119,N_4297,N_2919);
and U5120 (N_5120,N_4380,N_2792);
or U5121 (N_5121,N_4464,N_2565);
or U5122 (N_5122,N_3466,N_3780);
nor U5123 (N_5123,N_3402,N_4974);
or U5124 (N_5124,N_3513,N_3277);
or U5125 (N_5125,N_4871,N_4622);
or U5126 (N_5126,N_3019,N_4869);
nand U5127 (N_5127,N_3138,N_3663);
nor U5128 (N_5128,N_4914,N_4283);
nor U5129 (N_5129,N_3732,N_4880);
nand U5130 (N_5130,N_3933,N_3959);
or U5131 (N_5131,N_4350,N_4800);
and U5132 (N_5132,N_3612,N_4489);
nand U5133 (N_5133,N_3178,N_3450);
or U5134 (N_5134,N_3963,N_4416);
or U5135 (N_5135,N_3273,N_3614);
xnor U5136 (N_5136,N_3391,N_3084);
nand U5137 (N_5137,N_2628,N_3540);
or U5138 (N_5138,N_3386,N_2635);
or U5139 (N_5139,N_4318,N_3211);
xnor U5140 (N_5140,N_3876,N_4245);
xnor U5141 (N_5141,N_4476,N_4053);
or U5142 (N_5142,N_2860,N_3307);
or U5143 (N_5143,N_3144,N_3482);
or U5144 (N_5144,N_3123,N_4779);
nor U5145 (N_5145,N_3710,N_3925);
nor U5146 (N_5146,N_4862,N_2912);
xnor U5147 (N_5147,N_3392,N_3888);
or U5148 (N_5148,N_4492,N_2851);
nor U5149 (N_5149,N_3659,N_3587);
or U5150 (N_5150,N_3906,N_4358);
xor U5151 (N_5151,N_3171,N_4342);
nand U5152 (N_5152,N_4842,N_4338);
or U5153 (N_5153,N_4261,N_4044);
xor U5154 (N_5154,N_4230,N_2814);
nor U5155 (N_5155,N_3210,N_4752);
nand U5156 (N_5156,N_2870,N_4528);
xor U5157 (N_5157,N_4189,N_3824);
nor U5158 (N_5158,N_3341,N_4760);
xor U5159 (N_5159,N_3129,N_3279);
nor U5160 (N_5160,N_4221,N_4035);
xor U5161 (N_5161,N_3385,N_2772);
and U5162 (N_5162,N_3983,N_4259);
xor U5163 (N_5163,N_4875,N_4817);
and U5164 (N_5164,N_3025,N_4945);
or U5165 (N_5165,N_4312,N_4687);
nor U5166 (N_5166,N_4661,N_4888);
nand U5167 (N_5167,N_2534,N_3059);
nor U5168 (N_5168,N_3866,N_4072);
nor U5169 (N_5169,N_3217,N_4722);
nor U5170 (N_5170,N_2793,N_2621);
and U5171 (N_5171,N_3982,N_2600);
or U5172 (N_5172,N_4904,N_4576);
and U5173 (N_5173,N_3686,N_3928);
nor U5174 (N_5174,N_4466,N_2518);
xor U5175 (N_5175,N_3109,N_4162);
nor U5176 (N_5176,N_4776,N_2990);
or U5177 (N_5177,N_4839,N_3685);
or U5178 (N_5178,N_3023,N_3146);
nor U5179 (N_5179,N_3621,N_2616);
or U5180 (N_5180,N_4596,N_4728);
and U5181 (N_5181,N_4357,N_4200);
nand U5182 (N_5182,N_3239,N_3674);
and U5183 (N_5183,N_4271,N_4998);
xor U5184 (N_5184,N_4246,N_3311);
nand U5185 (N_5185,N_3676,N_4627);
xor U5186 (N_5186,N_3923,N_3281);
xnor U5187 (N_5187,N_3533,N_3860);
nand U5188 (N_5188,N_3057,N_3892);
or U5189 (N_5189,N_4511,N_4136);
nand U5190 (N_5190,N_3107,N_4621);
nor U5191 (N_5191,N_2893,N_4497);
xor U5192 (N_5192,N_4521,N_4101);
xor U5193 (N_5193,N_4698,N_4586);
nand U5194 (N_5194,N_3297,N_4241);
nor U5195 (N_5195,N_3099,N_3100);
and U5196 (N_5196,N_2915,N_4634);
and U5197 (N_5197,N_3543,N_4854);
and U5198 (N_5198,N_2654,N_2837);
nor U5199 (N_5199,N_4295,N_4404);
nand U5200 (N_5200,N_2846,N_2546);
and U5201 (N_5201,N_4048,N_4649);
or U5202 (N_5202,N_2697,N_4268);
nand U5203 (N_5203,N_3419,N_2716);
xnor U5204 (N_5204,N_4152,N_4647);
and U5205 (N_5205,N_2530,N_3638);
xnor U5206 (N_5206,N_4997,N_3200);
or U5207 (N_5207,N_3909,N_3817);
and U5208 (N_5208,N_3228,N_2765);
and U5209 (N_5209,N_3497,N_2766);
and U5210 (N_5210,N_4990,N_4918);
nor U5211 (N_5211,N_2918,N_4867);
or U5212 (N_5212,N_3535,N_3344);
and U5213 (N_5213,N_3837,N_2979);
or U5214 (N_5214,N_4068,N_4614);
or U5215 (N_5215,N_4996,N_3435);
or U5216 (N_5216,N_3426,N_3743);
nor U5217 (N_5217,N_4789,N_3563);
xor U5218 (N_5218,N_4653,N_3575);
nor U5219 (N_5219,N_4509,N_4478);
xor U5220 (N_5220,N_4104,N_3940);
xor U5221 (N_5221,N_3026,N_4149);
and U5222 (N_5222,N_2827,N_3413);
or U5223 (N_5223,N_3723,N_4694);
nor U5224 (N_5224,N_2647,N_3104);
and U5225 (N_5225,N_3458,N_3369);
nor U5226 (N_5226,N_4824,N_3167);
or U5227 (N_5227,N_4465,N_2669);
nand U5228 (N_5228,N_4151,N_4702);
or U5229 (N_5229,N_3207,N_2858);
nand U5230 (N_5230,N_3499,N_3718);
or U5231 (N_5231,N_4056,N_3949);
nor U5232 (N_5232,N_3921,N_4147);
or U5233 (N_5233,N_3671,N_3110);
nor U5234 (N_5234,N_3838,N_3713);
nand U5235 (N_5235,N_3186,N_2587);
nand U5236 (N_5236,N_4898,N_4292);
nor U5237 (N_5237,N_4022,N_2898);
nor U5238 (N_5238,N_3992,N_4392);
xor U5239 (N_5239,N_4662,N_2833);
or U5240 (N_5240,N_2543,N_3619);
nand U5241 (N_5241,N_4878,N_3596);
xnor U5242 (N_5242,N_2760,N_3296);
nor U5243 (N_5243,N_4611,N_4493);
and U5244 (N_5244,N_4305,N_3647);
nor U5245 (N_5245,N_4303,N_4428);
or U5246 (N_5246,N_3404,N_2883);
and U5247 (N_5247,N_3215,N_2817);
xnor U5248 (N_5248,N_2732,N_4617);
xnor U5249 (N_5249,N_3738,N_4337);
and U5250 (N_5250,N_2540,N_3305);
and U5251 (N_5251,N_3679,N_3154);
or U5252 (N_5252,N_4609,N_4106);
or U5253 (N_5253,N_3915,N_4995);
xor U5254 (N_5254,N_4561,N_4923);
or U5255 (N_5255,N_3822,N_3937);
nand U5256 (N_5256,N_3855,N_4197);
nand U5257 (N_5257,N_4774,N_2615);
or U5258 (N_5258,N_3424,N_3630);
nor U5259 (N_5259,N_4759,N_3074);
and U5260 (N_5260,N_4232,N_3971);
and U5261 (N_5261,N_2597,N_3834);
nand U5262 (N_5262,N_3920,N_3945);
and U5263 (N_5263,N_3908,N_3856);
and U5264 (N_5264,N_2854,N_4157);
and U5265 (N_5265,N_3054,N_4316);
and U5266 (N_5266,N_3248,N_3398);
nand U5267 (N_5267,N_4396,N_4090);
nand U5268 (N_5268,N_4570,N_3632);
nor U5269 (N_5269,N_4515,N_2550);
nor U5270 (N_5270,N_3598,N_3720);
or U5271 (N_5271,N_4459,N_2700);
nand U5272 (N_5272,N_4159,N_3149);
or U5273 (N_5273,N_4043,N_2819);
nand U5274 (N_5274,N_4641,N_4186);
nand U5275 (N_5275,N_3654,N_2670);
and U5276 (N_5276,N_4349,N_4868);
or U5277 (N_5277,N_3020,N_2513);
nand U5278 (N_5278,N_4138,N_4474);
nor U5279 (N_5279,N_4856,N_4933);
and U5280 (N_5280,N_3683,N_4893);
xnor U5281 (N_5281,N_3826,N_3825);
nand U5282 (N_5282,N_3571,N_4607);
xnor U5283 (N_5283,N_3265,N_3807);
xnor U5284 (N_5284,N_4681,N_4659);
xnor U5285 (N_5285,N_3183,N_4543);
nor U5286 (N_5286,N_4429,N_3649);
nand U5287 (N_5287,N_2523,N_4411);
nor U5288 (N_5288,N_2831,N_2801);
xor U5289 (N_5289,N_4439,N_4169);
or U5290 (N_5290,N_3844,N_3223);
or U5291 (N_5291,N_2864,N_2863);
nor U5292 (N_5292,N_3373,N_4005);
xnor U5293 (N_5293,N_2542,N_3105);
xnor U5294 (N_5294,N_4385,N_4772);
or U5295 (N_5295,N_3845,N_3484);
xor U5296 (N_5296,N_3661,N_3974);
and U5297 (N_5297,N_4420,N_3400);
nand U5298 (N_5298,N_2694,N_2838);
nand U5299 (N_5299,N_4244,N_4705);
or U5300 (N_5300,N_3101,N_4500);
or U5301 (N_5301,N_4346,N_2704);
and U5302 (N_5302,N_3264,N_3597);
nor U5303 (N_5303,N_2808,N_2673);
and U5304 (N_5304,N_3585,N_4966);
nand U5305 (N_5305,N_3873,N_3117);
xor U5306 (N_5306,N_4573,N_2871);
xnor U5307 (N_5307,N_4889,N_2934);
and U5308 (N_5308,N_3890,N_3280);
nor U5309 (N_5309,N_3986,N_3330);
and U5310 (N_5310,N_2715,N_4423);
or U5311 (N_5311,N_2607,N_3960);
or U5312 (N_5312,N_3014,N_4600);
nor U5313 (N_5313,N_4676,N_3754);
and U5314 (N_5314,N_3604,N_4947);
nor U5315 (N_5315,N_4656,N_4989);
or U5316 (N_5316,N_3829,N_4587);
xor U5317 (N_5317,N_3078,N_3030);
or U5318 (N_5318,N_2782,N_3670);
and U5319 (N_5319,N_3263,N_4133);
or U5320 (N_5320,N_4045,N_2964);
and U5321 (N_5321,N_3871,N_2737);
nand U5322 (N_5322,N_3793,N_2690);
and U5323 (N_5323,N_2929,N_3075);
nor U5324 (N_5324,N_2859,N_3643);
nand U5325 (N_5325,N_4613,N_3325);
nor U5326 (N_5326,N_2904,N_4529);
or U5327 (N_5327,N_2889,N_4213);
nand U5328 (N_5328,N_2507,N_4844);
xnor U5329 (N_5329,N_4374,N_4007);
xor U5330 (N_5330,N_4667,N_2734);
xnor U5331 (N_5331,N_3290,N_4547);
nor U5332 (N_5332,N_3648,N_3234);
xor U5333 (N_5333,N_4802,N_2840);
nor U5334 (N_5334,N_2830,N_4107);
or U5335 (N_5335,N_3141,N_3040);
nor U5336 (N_5336,N_4287,N_4532);
xor U5337 (N_5337,N_3573,N_3288);
xor U5338 (N_5338,N_4873,N_3089);
or U5339 (N_5339,N_3121,N_3990);
or U5340 (N_5340,N_2596,N_3682);
xor U5341 (N_5341,N_3382,N_3756);
or U5342 (N_5342,N_2701,N_3464);
or U5343 (N_5343,N_3352,N_3463);
xor U5344 (N_5344,N_4601,N_2834);
nor U5345 (N_5345,N_4272,N_2574);
nand U5346 (N_5346,N_2959,N_4356);
or U5347 (N_5347,N_3389,N_3453);
or U5348 (N_5348,N_4757,N_4121);
and U5349 (N_5349,N_3375,N_2933);
nand U5350 (N_5350,N_3486,N_3606);
xor U5351 (N_5351,N_4351,N_3355);
and U5352 (N_5352,N_3492,N_2541);
or U5353 (N_5353,N_3887,N_2535);
nand U5354 (N_5354,N_3401,N_3079);
and U5355 (N_5355,N_4657,N_4102);
nand U5356 (N_5356,N_2985,N_3480);
and U5357 (N_5357,N_3997,N_4333);
xnor U5358 (N_5358,N_4093,N_3405);
and U5359 (N_5359,N_3033,N_4843);
nand U5360 (N_5360,N_4463,N_3697);
nor U5361 (N_5361,N_3578,N_4412);
or U5362 (N_5362,N_4896,N_3656);
nand U5363 (N_5363,N_2551,N_2759);
nand U5364 (N_5364,N_3795,N_4360);
nand U5365 (N_5365,N_2672,N_4375);
xnor U5366 (N_5366,N_4001,N_3969);
nor U5367 (N_5367,N_3706,N_4379);
nand U5368 (N_5368,N_3693,N_2974);
nor U5369 (N_5369,N_4215,N_3741);
xnor U5370 (N_5370,N_3176,N_4536);
xor U5371 (N_5371,N_3962,N_2709);
xor U5372 (N_5372,N_3867,N_4250);
or U5373 (N_5373,N_3745,N_4688);
nand U5374 (N_5374,N_3036,N_4270);
nor U5375 (N_5375,N_4483,N_3814);
nand U5376 (N_5376,N_4899,N_4444);
and U5377 (N_5377,N_4218,N_4739);
nor U5378 (N_5378,N_3368,N_3802);
or U5379 (N_5379,N_4940,N_2586);
nor U5380 (N_5380,N_3917,N_3006);
nor U5381 (N_5381,N_3813,N_4881);
or U5382 (N_5382,N_3771,N_4279);
nor U5383 (N_5383,N_3695,N_3727);
or U5384 (N_5384,N_4796,N_4762);
nand U5385 (N_5385,N_4978,N_4616);
nand U5386 (N_5386,N_4011,N_3633);
or U5387 (N_5387,N_4849,N_2812);
nor U5388 (N_5388,N_4519,N_4745);
nand U5389 (N_5389,N_3348,N_3524);
nor U5390 (N_5390,N_4184,N_4435);
nor U5391 (N_5391,N_4384,N_4115);
or U5392 (N_5392,N_2991,N_3488);
xor U5393 (N_5393,N_4803,N_2950);
or U5394 (N_5394,N_4679,N_3160);
and U5395 (N_5395,N_3610,N_3832);
or U5396 (N_5396,N_3397,N_3880);
and U5397 (N_5397,N_3995,N_2894);
xor U5398 (N_5398,N_3615,N_3553);
or U5399 (N_5399,N_4087,N_2698);
or U5400 (N_5400,N_2751,N_3346);
xnor U5401 (N_5401,N_4517,N_4794);
nor U5402 (N_5402,N_4141,N_3835);
or U5403 (N_5403,N_3471,N_3156);
or U5404 (N_5404,N_3132,N_4178);
nor U5405 (N_5405,N_3274,N_4340);
nand U5406 (N_5406,N_2853,N_4716);
nor U5407 (N_5407,N_3555,N_2572);
or U5408 (N_5408,N_2580,N_3874);
nand U5409 (N_5409,N_3423,N_4243);
nand U5410 (N_5410,N_3283,N_4002);
nand U5411 (N_5411,N_4541,N_3700);
xor U5412 (N_5412,N_2931,N_3491);
xor U5413 (N_5413,N_2869,N_4818);
or U5414 (N_5414,N_4498,N_3652);
nor U5415 (N_5415,N_2780,N_4161);
and U5416 (N_5416,N_4256,N_4949);
and U5417 (N_5417,N_3192,N_3190);
and U5418 (N_5418,N_3953,N_2560);
nor U5419 (N_5419,N_2544,N_2998);
xnor U5420 (N_5420,N_4965,N_4954);
nor U5421 (N_5421,N_4486,N_4835);
or U5422 (N_5422,N_3015,N_3981);
nor U5423 (N_5423,N_4567,N_3094);
xor U5424 (N_5424,N_4512,N_3417);
or U5425 (N_5425,N_3852,N_3329);
nor U5426 (N_5426,N_4266,N_4344);
or U5427 (N_5427,N_2652,N_4037);
nor U5428 (N_5428,N_3310,N_3605);
xor U5429 (N_5429,N_4253,N_4183);
and U5430 (N_5430,N_2921,N_4734);
nor U5431 (N_5431,N_4377,N_2506);
xnor U5432 (N_5432,N_4790,N_4019);
nand U5433 (N_5433,N_3688,N_3879);
and U5434 (N_5434,N_3895,N_4274);
and U5435 (N_5435,N_3820,N_4258);
and U5436 (N_5436,N_3383,N_3193);
or U5437 (N_5437,N_3851,N_2969);
nand U5438 (N_5438,N_4806,N_3529);
xnor U5439 (N_5439,N_4594,N_4678);
xor U5440 (N_5440,N_4624,N_4700);
or U5441 (N_5441,N_4650,N_4129);
and U5442 (N_5442,N_4188,N_4958);
nor U5443 (N_5443,N_3593,N_3198);
nor U5444 (N_5444,N_3646,N_2601);
and U5445 (N_5445,N_3140,N_2649);
or U5446 (N_5446,N_3284,N_3616);
nor U5447 (N_5447,N_2908,N_3699);
or U5448 (N_5448,N_4325,N_4826);
xnor U5449 (N_5449,N_3570,N_3153);
and U5450 (N_5450,N_4092,N_3765);
nor U5451 (N_5451,N_2595,N_4632);
nand U5452 (N_5452,N_3336,N_4919);
nand U5453 (N_5453,N_4581,N_4260);
xnor U5454 (N_5454,N_2899,N_3261);
nor U5455 (N_5455,N_3185,N_3009);
nor U5456 (N_5456,N_3759,N_4648);
nor U5457 (N_5457,N_3351,N_2967);
and U5458 (N_5458,N_3053,N_4487);
nand U5459 (N_5459,N_3347,N_4477);
or U5460 (N_5460,N_2712,N_3189);
nor U5461 (N_5461,N_3113,N_3017);
and U5462 (N_5462,N_4792,N_4199);
nor U5463 (N_5463,N_4363,N_3958);
nand U5464 (N_5464,N_4526,N_2749);
or U5465 (N_5465,N_4315,N_3358);
xnor U5466 (N_5466,N_2547,N_2684);
or U5467 (N_5467,N_2588,N_3043);
nor U5468 (N_5468,N_4057,N_3902);
nand U5469 (N_5469,N_3320,N_3254);
nor U5470 (N_5470,N_3595,N_3857);
xor U5471 (N_5471,N_3119,N_4145);
xor U5472 (N_5472,N_4571,N_3678);
nand U5473 (N_5473,N_3291,N_3112);
or U5474 (N_5474,N_4216,N_3165);
and U5475 (N_5475,N_3905,N_4639);
nand U5476 (N_5476,N_3797,N_2963);
and U5477 (N_5477,N_4780,N_3804);
nor U5478 (N_5478,N_4335,N_4929);
xnor U5479 (N_5479,N_3734,N_2515);
and U5480 (N_5480,N_2613,N_4905);
nor U5481 (N_5481,N_2630,N_3586);
nor U5482 (N_5482,N_3349,N_4516);
and U5483 (N_5483,N_4367,N_2810);
nor U5484 (N_5484,N_2768,N_2536);
xnor U5485 (N_5485,N_4693,N_2785);
nor U5486 (N_5486,N_2767,N_3312);
xor U5487 (N_5487,N_3422,N_3831);
nand U5488 (N_5488,N_3664,N_4016);
xor U5489 (N_5489,N_4079,N_2641);
xor U5490 (N_5490,N_3843,N_3712);
nor U5491 (N_5491,N_2680,N_2932);
nor U5492 (N_5492,N_4372,N_4715);
or U5493 (N_5493,N_3984,N_3539);
nand U5494 (N_5494,N_3442,N_2980);
and U5495 (N_5495,N_4391,N_4501);
xor U5496 (N_5496,N_3818,N_4430);
xor U5497 (N_5497,N_2862,N_3896);
or U5498 (N_5498,N_3083,N_3196);
or U5499 (N_5499,N_2975,N_3475);
nand U5500 (N_5500,N_4701,N_3478);
or U5501 (N_5501,N_4442,N_2994);
or U5502 (N_5502,N_4848,N_2519);
and U5503 (N_5503,N_4504,N_4052);
nor U5504 (N_5504,N_4014,N_3527);
or U5505 (N_5505,N_2825,N_4957);
nand U5506 (N_5506,N_4010,N_4740);
xnor U5507 (N_5507,N_3256,N_3973);
xnor U5508 (N_5508,N_3894,N_4505);
and U5509 (N_5509,N_3222,N_4564);
nor U5510 (N_5510,N_3016,N_4164);
nand U5511 (N_5511,N_3447,N_2591);
or U5512 (N_5512,N_3628,N_4675);
nor U5513 (N_5513,N_3667,N_2777);
and U5514 (N_5514,N_2763,N_2579);
or U5515 (N_5515,N_3108,N_2984);
or U5516 (N_5516,N_4636,N_2516);
nor U5517 (N_5517,N_4955,N_4506);
xnor U5518 (N_5518,N_3035,N_4395);
and U5519 (N_5519,N_2538,N_4083);
or U5520 (N_5520,N_3428,N_4710);
nor U5521 (N_5521,N_2911,N_3481);
xor U5522 (N_5522,N_3942,N_4247);
xor U5523 (N_5523,N_3080,N_2548);
nor U5524 (N_5524,N_3213,N_3270);
xnor U5525 (N_5525,N_3479,N_2815);
or U5526 (N_5526,N_2798,N_2752);
or U5527 (N_5527,N_4767,N_2770);
or U5528 (N_5528,N_4579,N_4225);
nand U5529 (N_5529,N_2527,N_3547);
nor U5530 (N_5530,N_4643,N_4985);
and U5531 (N_5531,N_2997,N_2946);
or U5532 (N_5532,N_4475,N_2855);
nand U5533 (N_5533,N_2968,N_3936);
nor U5534 (N_5534,N_4602,N_2692);
nand U5535 (N_5535,N_4719,N_3427);
xnor U5536 (N_5536,N_2906,N_4744);
nand U5537 (N_5537,N_3651,N_4112);
and U5538 (N_5538,N_4882,N_3631);
or U5539 (N_5539,N_4032,N_4264);
and U5540 (N_5540,N_3245,N_3924);
nor U5541 (N_5541,N_3356,N_4494);
nor U5542 (N_5542,N_4931,N_4301);
and U5543 (N_5543,N_4455,N_3195);
xnor U5544 (N_5544,N_3139,N_3526);
or U5545 (N_5545,N_4387,N_4906);
and U5546 (N_5546,N_3739,N_3785);
xnor U5547 (N_5547,N_4599,N_3763);
and U5548 (N_5548,N_4122,N_3267);
or U5549 (N_5549,N_3206,N_3275);
and U5550 (N_5550,N_3181,N_3412);
or U5551 (N_5551,N_2897,N_2797);
or U5552 (N_5552,N_2593,N_4962);
nand U5553 (N_5553,N_3846,N_4838);
xnor U5554 (N_5554,N_4359,N_2537);
and U5555 (N_5555,N_2942,N_3776);
or U5556 (N_5556,N_3833,N_3063);
nor U5557 (N_5557,N_2747,N_2920);
or U5558 (N_5558,N_3175,N_4309);
nor U5559 (N_5559,N_2976,N_3556);
nor U5560 (N_5560,N_3840,N_3010);
or U5561 (N_5561,N_2957,N_4108);
and U5562 (N_5562,N_3907,N_3572);
or U5563 (N_5563,N_4578,N_4540);
xnor U5564 (N_5564,N_3120,N_3980);
or U5565 (N_5565,N_4827,N_3691);
xor U5566 (N_5566,N_2555,N_2804);
nor U5567 (N_5567,N_3965,N_4362);
nand U5568 (N_5568,N_4422,N_3414);
or U5569 (N_5569,N_4299,N_3506);
nor U5570 (N_5570,N_2944,N_4620);
or U5571 (N_5571,N_2645,N_4670);
or U5572 (N_5572,N_3174,N_3581);
xor U5573 (N_5573,N_4706,N_4858);
nand U5574 (N_5574,N_3926,N_2608);
nand U5575 (N_5575,N_3411,N_4321);
xor U5576 (N_5576,N_3011,N_3042);
and U5577 (N_5577,N_3768,N_3438);
and U5578 (N_5578,N_4015,N_4733);
xor U5579 (N_5579,N_2524,N_4936);
or U5580 (N_5580,N_4319,N_4174);
nor U5581 (N_5581,N_4160,N_3058);
xnor U5582 (N_5582,N_4591,N_2696);
nor U5583 (N_5583,N_3255,N_4371);
nor U5584 (N_5584,N_4574,N_4263);
nor U5585 (N_5585,N_3444,N_4708);
xor U5586 (N_5586,N_2790,N_2717);
and U5587 (N_5587,N_4836,N_2653);
nor U5588 (N_5588,N_4748,N_3362);
nor U5589 (N_5589,N_4897,N_3590);
or U5590 (N_5590,N_3791,N_4088);
or U5591 (N_5591,N_3418,N_4211);
and U5592 (N_5592,N_4039,N_4482);
xor U5593 (N_5593,N_4434,N_4988);
or U5594 (N_5594,N_3673,N_4964);
and U5595 (N_5595,N_3399,N_4631);
or U5596 (N_5596,N_4262,N_4009);
xnor U5597 (N_5597,N_4214,N_3301);
nor U5598 (N_5598,N_4961,N_3177);
nand U5599 (N_5599,N_3434,N_4114);
or U5600 (N_5600,N_2805,N_3219);
xor U5601 (N_5601,N_4131,N_4403);
or U5602 (N_5602,N_4273,N_4255);
or U5603 (N_5603,N_2901,N_4436);
xnor U5604 (N_5604,N_2987,N_3240);
nand U5605 (N_5605,N_2839,N_3258);
nor U5606 (N_5606,N_4669,N_3753);
nand U5607 (N_5607,N_4389,N_4963);
nor U5608 (N_5608,N_4566,N_4139);
nor U5609 (N_5609,N_3853,N_2636);
nand U5610 (N_5610,N_3993,N_3069);
nand U5611 (N_5611,N_3501,N_3135);
and U5612 (N_5612,N_2970,N_3237);
nor U5613 (N_5613,N_4222,N_4144);
nand U5614 (N_5614,N_3007,N_3952);
or U5615 (N_5615,N_4651,N_4341);
nand U5616 (N_5616,N_4453,N_4210);
nand U5617 (N_5617,N_4064,N_2992);
nand U5618 (N_5618,N_4099,N_3787);
nor U5619 (N_5619,N_3182,N_4191);
nand U5620 (N_5620,N_3257,N_4984);
and U5621 (N_5621,N_4097,N_4583);
nor U5622 (N_5622,N_4251,N_4510);
nor U5623 (N_5623,N_3209,N_4126);
xor U5624 (N_5624,N_3557,N_3134);
xor U5625 (N_5625,N_4055,N_2663);
or U5626 (N_5626,N_3989,N_3039);
nand U5627 (N_5627,N_3188,N_2526);
nand U5628 (N_5628,N_4322,N_3436);
nor U5629 (N_5629,N_3180,N_3420);
nor U5630 (N_5630,N_2657,N_2916);
and U5631 (N_5631,N_3477,N_3448);
nor U5632 (N_5632,N_3809,N_3031);
xnor U5633 (N_5633,N_4071,N_2907);
and U5634 (N_5634,N_2581,N_3157);
nor U5635 (N_5635,N_2794,N_3875);
nor U5636 (N_5636,N_4234,N_3898);
xnor U5637 (N_5637,N_3294,N_3292);
nand U5638 (N_5638,N_3748,N_3740);
xor U5639 (N_5639,N_4450,N_2556);
nand U5640 (N_5640,N_2720,N_4267);
and U5641 (N_5641,N_4153,N_4076);
and U5642 (N_5642,N_3914,N_2962);
nor U5643 (N_5643,N_4202,N_2584);
xnor U5644 (N_5644,N_3022,N_4408);
nor U5645 (N_5645,N_2744,N_3088);
or U5646 (N_5646,N_3944,N_3977);
nor U5647 (N_5647,N_4249,N_3081);
nand U5648 (N_5648,N_4329,N_2633);
nand U5649 (N_5649,N_4668,N_4808);
and U5650 (N_5650,N_3202,N_2660);
xnor U5651 (N_5651,N_3361,N_2638);
nand U5652 (N_5652,N_3884,N_2999);
nand U5653 (N_5653,N_3096,N_4397);
nor U5654 (N_5654,N_4294,N_4785);
and U5655 (N_5655,N_2926,N_3886);
and U5656 (N_5656,N_4111,N_4204);
xnor U5657 (N_5657,N_2995,N_3468);
and U5658 (N_5658,N_4753,N_4535);
xor U5659 (N_5659,N_3967,N_4801);
xnor U5660 (N_5660,N_4732,N_4331);
xnor U5661 (N_5661,N_4179,N_3766);
or U5662 (N_5662,N_3836,N_3561);
or U5663 (N_5663,N_4712,N_3354);
or U5664 (N_5664,N_2844,N_3242);
or U5665 (N_5665,N_4876,N_4994);
nor U5666 (N_5666,N_3943,N_3179);
nor U5667 (N_5667,N_4448,N_4883);
or U5668 (N_5668,N_3131,N_2566);
and U5669 (N_5669,N_4913,N_3583);
nor U5670 (N_5670,N_4495,N_2936);
nor U5671 (N_5671,N_3608,N_2958);
and U5672 (N_5672,N_3403,N_3639);
nand U5673 (N_5673,N_2612,N_4447);
xnor U5674 (N_5674,N_4673,N_4750);
or U5675 (N_5675,N_3576,N_3253);
nor U5676 (N_5676,N_4481,N_2813);
or U5677 (N_5677,N_2622,N_3359);
and U5678 (N_5678,N_4059,N_2940);
or U5679 (N_5679,N_4376,N_3864);
nand U5680 (N_5680,N_3801,N_3137);
nand U5681 (N_5681,N_3999,N_4554);
nor U5682 (N_5682,N_2960,N_3847);
xnor U5683 (N_5683,N_4799,N_4499);
or U5684 (N_5684,N_4180,N_3978);
or U5685 (N_5685,N_4777,N_3018);
nand U5686 (N_5686,N_3929,N_4451);
and U5687 (N_5687,N_4588,N_4028);
nor U5688 (N_5688,N_4438,N_4604);
nor U5689 (N_5689,N_4415,N_2849);
xor U5690 (N_5690,N_4804,N_4365);
and U5691 (N_5691,N_4550,N_4518);
or U5692 (N_5692,N_4718,N_3067);
or U5693 (N_5693,N_2986,N_4503);
nand U5694 (N_5694,N_4672,N_2856);
or U5695 (N_5695,N_3806,N_2675);
nor U5696 (N_5696,N_2873,N_3530);
nand U5697 (N_5697,N_4575,N_3650);
nand U5698 (N_5698,N_4684,N_3126);
xor U5699 (N_5699,N_3068,N_4116);
xnor U5700 (N_5700,N_2758,N_4944);
or U5701 (N_5701,N_3439,N_4910);
nand U5702 (N_5702,N_2956,N_3151);
nor U5703 (N_5703,N_3410,N_4426);
or U5704 (N_5704,N_3955,N_4461);
or U5705 (N_5705,N_3287,N_4555);
nor U5706 (N_5706,N_4117,N_2861);
nand U5707 (N_5707,N_3514,N_3538);
nand U5708 (N_5708,N_3841,N_3469);
and U5709 (N_5709,N_3680,N_4786);
nand U5710 (N_5710,N_3269,N_3815);
nand U5711 (N_5711,N_3328,N_4530);
or U5712 (N_5712,N_3574,N_3086);
nand U5713 (N_5713,N_2835,N_2665);
and U5714 (N_5714,N_2617,N_3148);
or U5715 (N_5715,N_3601,N_3900);
or U5716 (N_5716,N_4680,N_4419);
xor U5717 (N_5717,N_2662,N_3360);
or U5718 (N_5718,N_4637,N_4082);
nand U5719 (N_5719,N_3049,N_4081);
nand U5720 (N_5720,N_2748,N_4484);
and U5721 (N_5721,N_2501,N_3158);
xnor U5722 (N_5722,N_4782,N_4078);
xnor U5723 (N_5723,N_3947,N_2611);
nor U5724 (N_5724,N_3767,N_4046);
and U5725 (N_5725,N_3830,N_4825);
xor U5726 (N_5726,N_2948,N_3964);
and U5727 (N_5727,N_3169,N_2756);
or U5728 (N_5728,N_4832,N_4290);
and U5729 (N_5729,N_4870,N_3617);
xor U5730 (N_5730,N_3516,N_2637);
and U5731 (N_5731,N_3607,N_3164);
and U5732 (N_5732,N_4992,N_3339);
nor U5733 (N_5733,N_3304,N_3050);
xor U5734 (N_5734,N_3696,N_3041);
nor U5735 (N_5735,N_4238,N_3390);
nand U5736 (N_5736,N_4853,N_3001);
and U5737 (N_5737,N_2677,N_3125);
nand U5738 (N_5738,N_2880,N_4257);
xor U5739 (N_5739,N_3065,N_4281);
nor U5740 (N_5740,N_3002,N_3246);
xnor U5741 (N_5741,N_3332,N_4239);
or U5742 (N_5742,N_3087,N_4927);
xnor U5743 (N_5743,N_4327,N_4073);
nand U5744 (N_5744,N_2710,N_4192);
xnor U5745 (N_5745,N_3788,N_3554);
nor U5746 (N_5746,N_4831,N_4908);
nor U5747 (N_5747,N_3168,N_3901);
or U5748 (N_5748,N_3620,N_3322);
or U5749 (N_5749,N_4381,N_3805);
nor U5750 (N_5750,N_4606,N_4857);
or U5751 (N_5751,N_3930,N_4548);
and U5752 (N_5752,N_3214,N_4860);
and U5753 (N_5753,N_3549,N_2702);
xnor U5754 (N_5754,N_4968,N_4932);
nor U5755 (N_5755,N_4747,N_2576);
nor U5756 (N_5756,N_4040,N_2558);
xnor U5757 (N_5757,N_3935,N_4840);
nor U5758 (N_5758,N_4556,N_2896);
nand U5759 (N_5759,N_4714,N_2753);
or U5760 (N_5760,N_2522,N_2650);
xnor U5761 (N_5761,N_2809,N_3698);
xor U5762 (N_5762,N_4110,N_3839);
nand U5763 (N_5763,N_3152,N_3579);
or U5764 (N_5764,N_3869,N_3064);
nand U5765 (N_5765,N_4182,N_2993);
and U5766 (N_5766,N_4764,N_3201);
and U5767 (N_5767,N_4382,N_4036);
nor U5768 (N_5768,N_2978,N_3147);
nand U5769 (N_5769,N_4237,N_4018);
xnor U5770 (N_5770,N_3461,N_3523);
and U5771 (N_5771,N_3918,N_3051);
nor U5772 (N_5772,N_4207,N_3792);
or U5773 (N_5773,N_4288,N_4797);
and U5774 (N_5774,N_4689,N_4727);
and U5775 (N_5775,N_3565,N_2514);
or U5776 (N_5776,N_4460,N_4172);
xnor U5777 (N_5777,N_3394,N_4663);
nor U5778 (N_5778,N_3934,N_2623);
xor U5779 (N_5779,N_3449,N_4959);
xnor U5780 (N_5780,N_4851,N_4813);
nand U5781 (N_5781,N_4124,N_4185);
nand U5782 (N_5782,N_3452,N_3522);
nand U5783 (N_5783,N_3692,N_3314);
and U5784 (N_5784,N_3266,N_2724);
or U5785 (N_5785,N_4749,N_3046);
or U5786 (N_5786,N_4398,N_4031);
xnor U5787 (N_5787,N_4020,N_4027);
or U5788 (N_5788,N_2847,N_3395);
nor U5789 (N_5789,N_4348,N_2909);
and U5790 (N_5790,N_4085,N_4148);
nor U5791 (N_5791,N_2609,N_3191);
xor U5792 (N_5792,N_4953,N_2605);
xnor U5793 (N_5793,N_2922,N_3658);
or U5794 (N_5794,N_2528,N_3451);
xnor U5795 (N_5795,N_3772,N_4024);
nand U5796 (N_5796,N_3308,N_4907);
or U5797 (N_5797,N_3799,N_3409);
nor U5798 (N_5798,N_3249,N_3863);
nor U5799 (N_5799,N_3662,N_3872);
xnor U5800 (N_5800,N_3076,N_2682);
nand U5801 (N_5801,N_4823,N_4941);
or U5802 (N_5802,N_3220,N_3927);
xnor U5803 (N_5803,N_2816,N_4584);
and U5804 (N_5804,N_4773,N_2779);
xor U5805 (N_5805,N_2656,N_2982);
nand U5806 (N_5806,N_3784,N_3221);
nor U5807 (N_5807,N_4837,N_4879);
xnor U5808 (N_5808,N_2567,N_4156);
and U5809 (N_5809,N_3988,N_4386);
nand U5810 (N_5810,N_3600,N_4452);
nor U5811 (N_5811,N_4619,N_3541);
nand U5812 (N_5812,N_4553,N_3333);
and U5813 (N_5813,N_4770,N_2930);
xor U5814 (N_5814,N_3085,N_4388);
and U5815 (N_5815,N_2549,N_3235);
and U5816 (N_5816,N_3762,N_4096);
and U5817 (N_5817,N_4177,N_4874);
nor U5818 (N_5818,N_3133,N_3324);
xnor U5819 (N_5819,N_4061,N_3970);
or U5820 (N_5820,N_2800,N_3611);
or U5821 (N_5821,N_4877,N_3603);
xnor U5822 (N_5822,N_2626,N_4580);
nand U5823 (N_5823,N_3056,N_2573);
nand U5824 (N_5824,N_3868,N_4713);
and U5825 (N_5825,N_4960,N_4520);
or U5826 (N_5826,N_4674,N_4937);
nand U5827 (N_5827,N_4563,N_4916);
nor U5828 (N_5828,N_4469,N_4240);
nand U5829 (N_5829,N_3913,N_4000);
xor U5830 (N_5830,N_4545,N_4741);
or U5831 (N_5831,N_3363,N_4502);
nor U5832 (N_5832,N_4926,N_4746);
nor U5833 (N_5833,N_4980,N_3922);
nand U5834 (N_5834,N_3376,N_4822);
nor U5835 (N_5835,N_3038,N_3364);
nor U5836 (N_5836,N_4707,N_3250);
and U5837 (N_5837,N_2510,N_3493);
nor U5838 (N_5838,N_3055,N_3961);
and U5839 (N_5839,N_4793,N_3289);
or U5840 (N_5840,N_4755,N_3779);
nand U5841 (N_5841,N_2741,N_3842);
nor U5842 (N_5842,N_3708,N_3731);
xnor U5843 (N_5843,N_4912,N_3736);
and U5844 (N_5844,N_3091,N_3987);
nor U5845 (N_5845,N_4726,N_4819);
xor U5846 (N_5846,N_4699,N_2787);
nand U5847 (N_5847,N_4399,N_2644);
nor U5848 (N_5848,N_4778,N_4023);
nand U5849 (N_5849,N_3735,N_3821);
nand U5850 (N_5850,N_4017,N_4173);
or U5851 (N_5851,N_2661,N_4280);
nor U5852 (N_5852,N_3588,N_3315);
nand U5853 (N_5853,N_4013,N_4697);
nor U5854 (N_5854,N_2845,N_4507);
nand U5855 (N_5855,N_4560,N_3687);
xor U5856 (N_5856,N_3459,N_2826);
nand U5857 (N_5857,N_2691,N_3582);
and U5858 (N_5858,N_2953,N_3548);
nor U5859 (N_5859,N_4783,N_4051);
xnor U5860 (N_5860,N_3285,N_3672);
or U5861 (N_5861,N_4558,N_4449);
nand U5862 (N_5862,N_3798,N_3462);
or U5863 (N_5863,N_4496,N_3640);
nor U5864 (N_5864,N_3800,N_3170);
and U5865 (N_5865,N_4490,N_4066);
nor U5866 (N_5866,N_3702,N_4485);
xor U5867 (N_5867,N_4265,N_4224);
and U5868 (N_5868,N_4254,N_3637);
or U5869 (N_5869,N_4917,N_3559);
xnor U5870 (N_5870,N_2502,N_4682);
or U5871 (N_5871,N_2807,N_3972);
nand U5872 (N_5872,N_4212,N_4074);
and U5873 (N_5873,N_4049,N_3550);
nor U5874 (N_5874,N_3758,N_4223);
nand U5875 (N_5875,N_2585,N_4170);
nand U5876 (N_5876,N_4635,N_3489);
and U5877 (N_5877,N_4533,N_3345);
xnor U5878 (N_5878,N_3976,N_4472);
and U5879 (N_5879,N_4330,N_3319);
nand U5880 (N_5880,N_2598,N_4033);
xnor U5881 (N_5881,N_2525,N_3128);
xnor U5882 (N_5882,N_3911,N_4393);
nor U5883 (N_5883,N_3951,N_3204);
or U5884 (N_5884,N_2703,N_3525);
nand U5885 (N_5885,N_4323,N_3008);
nor U5886 (N_5886,N_3430,N_3998);
nand U5887 (N_5887,N_3566,N_4527);
xnor U5888 (N_5888,N_2778,N_4431);
and U5889 (N_5889,N_4977,N_3897);
nand U5890 (N_5890,N_3318,N_3904);
or U5891 (N_5891,N_3694,N_4065);
nand U5892 (N_5892,N_3609,N_4508);
or U5893 (N_5893,N_4300,N_2666);
nand U5894 (N_5894,N_3244,N_4187);
nand U5895 (N_5895,N_3613,N_3052);
xor U5896 (N_5896,N_4654,N_2559);
xnor U5897 (N_5897,N_4633,N_4948);
and U5898 (N_5898,N_2648,N_2881);
nor U5899 (N_5899,N_3432,N_2520);
xnor U5900 (N_5900,N_4983,N_3127);
and U5901 (N_5901,N_2575,N_4866);
nand U5902 (N_5902,N_4551,N_4720);
xnor U5903 (N_5903,N_4278,N_2951);
nor U5904 (N_5904,N_4109,N_2725);
or U5905 (N_5905,N_4976,N_4971);
and U5906 (N_5906,N_3381,N_4951);
nor U5907 (N_5907,N_2625,N_3374);
or U5908 (N_5908,N_4135,N_4690);
nor U5909 (N_5909,N_3725,N_3985);
or U5910 (N_5910,N_4236,N_4421);
or U5911 (N_5911,N_4805,N_2818);
nand U5912 (N_5912,N_2836,N_4557);
or U5913 (N_5913,N_2771,N_2651);
xor U5914 (N_5914,N_2676,N_4242);
and U5915 (N_5915,N_4407,N_4441);
and U5916 (N_5916,N_4595,N_3470);
and U5917 (N_5917,N_4771,N_4886);
and U5918 (N_5918,N_3161,N_3306);
or U5919 (N_5919,N_3711,N_3562);
nor U5920 (N_5920,N_4892,N_4433);
nor U5921 (N_5921,N_3812,N_4336);
nor U5922 (N_5922,N_3717,N_4209);
xor U5923 (N_5923,N_3197,N_3854);
or U5924 (N_5924,N_2719,N_4655);
nand U5925 (N_5925,N_4815,N_2872);
xor U5926 (N_5926,N_3827,N_4437);
and U5927 (N_5927,N_3645,N_3979);
nand U5928 (N_5928,N_3689,N_4787);
nor U5929 (N_5929,N_4725,N_4479);
xnor U5930 (N_5930,N_4537,N_4798);
nor U5931 (N_5931,N_2791,N_4378);
nor U5932 (N_5932,N_4950,N_4695);
or U5933 (N_5933,N_3184,N_3483);
nand U5934 (N_5934,N_3665,N_3789);
nand U5935 (N_5935,N_3456,N_3716);
xnor U5936 (N_5936,N_2743,N_2884);
nand U5937 (N_5937,N_4742,N_4175);
xnor U5938 (N_5938,N_4754,N_4414);
and U5939 (N_5939,N_4166,N_3551);
or U5940 (N_5940,N_4220,N_3034);
or U5941 (N_5941,N_3061,N_3415);
nor U5942 (N_5942,N_2952,N_4390);
nand U5943 (N_5943,N_4737,N_4067);
nand U5944 (N_5944,N_4310,N_3342);
xnor U5945 (N_5945,N_4425,N_4546);
nor U5946 (N_5946,N_3421,N_4488);
and U5947 (N_5947,N_4758,N_4872);
xor U5948 (N_5948,N_4195,N_3726);
or U5949 (N_5949,N_4369,N_2811);
and U5950 (N_5950,N_2658,N_3532);
or U5951 (N_5951,N_3635,N_2738);
and U5952 (N_5952,N_4696,N_4730);
or U5953 (N_5953,N_4206,N_4054);
and U5954 (N_5954,N_4308,N_2789);
nand U5955 (N_5955,N_4943,N_3719);
and U5956 (N_5956,N_3916,N_4972);
and U5957 (N_5957,N_2614,N_4590);
nor U5958 (N_5958,N_2730,N_4775);
nor U5959 (N_5959,N_3095,N_4630);
and U5960 (N_5960,N_4373,N_3521);
nand U5961 (N_5961,N_3599,N_4645);
nor U5962 (N_5962,N_4830,N_2688);
nand U5963 (N_5963,N_2509,N_2945);
nor U5964 (N_5964,N_4895,N_4973);
or U5965 (N_5965,N_4863,N_4751);
and U5966 (N_5966,N_3229,N_3278);
nor U5967 (N_5967,N_4967,N_3474);
xnor U5968 (N_5968,N_3552,N_2879);
nor U5969 (N_5969,N_4952,N_3300);
and U5970 (N_5970,N_2634,N_3037);
nand U5971 (N_5971,N_4569,N_3938);
and U5972 (N_5972,N_3286,N_4320);
and U5973 (N_5973,N_3760,N_3337);
or U5974 (N_5974,N_3517,N_3657);
nor U5975 (N_5975,N_4562,N_3387);
and U5976 (N_5976,N_2888,N_4394);
nor U5977 (N_5977,N_2971,N_3406);
nor U5978 (N_5978,N_3236,N_4795);
nand U5979 (N_5979,N_3102,N_2803);
nand U5980 (N_5980,N_4366,N_4277);
nand U5981 (N_5981,N_4756,N_4400);
or U5982 (N_5982,N_3675,N_4119);
and U5983 (N_5983,N_4190,N_4736);
xnor U5984 (N_5984,N_4457,N_3260);
nand U5985 (N_5985,N_4784,N_4142);
and U5986 (N_5986,N_4592,N_2532);
and U5987 (N_5987,N_4456,N_2892);
or U5988 (N_5988,N_3757,N_3950);
xor U5989 (N_5989,N_2706,N_4935);
nor U5990 (N_5990,N_4163,N_4820);
or U5991 (N_5991,N_2562,N_3865);
nor U5992 (N_5992,N_3384,N_4513);
and U5993 (N_5993,N_4454,N_3327);
and U5994 (N_5994,N_4577,N_2890);
nand U5995 (N_5995,N_3331,N_4552);
nor U5996 (N_5996,N_3216,N_4565);
and U5997 (N_5997,N_4900,N_4781);
nor U5998 (N_5998,N_4004,N_2885);
nor U5999 (N_5999,N_4597,N_2762);
nand U6000 (N_6000,N_3684,N_4709);
nor U6001 (N_6001,N_4181,N_3568);
nand U6002 (N_6002,N_4810,N_3299);
and U6003 (N_6003,N_4677,N_4514);
xnor U6004 (N_6004,N_2583,N_2708);
xnor U6005 (N_6005,N_3460,N_3472);
nand U6006 (N_6006,N_3194,N_4629);
xor U6007 (N_6007,N_4491,N_2799);
nand U6008 (N_6008,N_3773,N_3893);
nor U6009 (N_6009,N_2705,N_4311);
xor U6010 (N_6010,N_4766,N_2983);
or U6011 (N_6011,N_4939,N_4070);
xnor U6012 (N_6012,N_4603,N_4686);
nor U6013 (N_6013,N_2687,N_3626);
or U6014 (N_6014,N_3769,N_4468);
or U6015 (N_6015,N_2714,N_2599);
and U6016 (N_6016,N_3668,N_3544);
nand U6017 (N_6017,N_2935,N_3302);
nor U6018 (N_6018,N_4008,N_2989);
nand U6019 (N_6019,N_2713,N_3510);
nor U6020 (N_6020,N_3321,N_2678);
and U6021 (N_6021,N_3494,N_4666);
nor U6022 (N_6022,N_3669,N_3786);
nor U6023 (N_6023,N_3343,N_4901);
and U6024 (N_6024,N_2795,N_3849);
xnor U6025 (N_6025,N_2642,N_3032);
nor U6026 (N_6026,N_4306,N_3077);
nor U6027 (N_6027,N_4134,N_4196);
nor U6028 (N_6028,N_2828,N_4729);
xnor U6029 (N_6029,N_3618,N_4094);
and U6030 (N_6030,N_4252,N_3282);
nand U6031 (N_6031,N_4069,N_3232);
nand U6032 (N_6032,N_3295,N_3932);
or U6033 (N_6033,N_4894,N_4304);
nor U6034 (N_6034,N_3303,N_2900);
nor U6035 (N_6035,N_4841,N_3495);
xnor U6036 (N_6036,N_4946,N_2955);
and U6037 (N_6037,N_3317,N_2554);
nand U6038 (N_6038,N_2842,N_4956);
or U6039 (N_6039,N_3848,N_3975);
xnor U6040 (N_6040,N_2603,N_2806);
xnor U6041 (N_6041,N_4610,N_4307);
xnor U6042 (N_6042,N_4761,N_3013);
xor U6043 (N_6043,N_3991,N_3948);
or U6044 (N_6044,N_2746,N_4703);
nand U6045 (N_6045,N_2820,N_4284);
or U6046 (N_6046,N_3704,N_3366);
or U6047 (N_6047,N_3251,N_3509);
nand U6048 (N_6048,N_4809,N_4539);
xor U6049 (N_6049,N_3338,N_4589);
and U6050 (N_6050,N_4091,N_4930);
xnor U6051 (N_6051,N_3660,N_4970);
xor U6052 (N_6052,N_3728,N_2913);
nand U6053 (N_6053,N_2627,N_2561);
or U6054 (N_6054,N_4981,N_4969);
xor U6055 (N_6055,N_4445,N_4047);
or U6056 (N_6056,N_2689,N_3625);
or U6057 (N_6057,N_3714,N_3770);
xor U6058 (N_6058,N_4999,N_3500);
xnor U6059 (N_6059,N_3407,N_4585);
or U6060 (N_6060,N_4029,N_3512);
and U6061 (N_6061,N_3243,N_3378);
xnor U6062 (N_6062,N_4531,N_2866);
xnor U6063 (N_6063,N_3627,N_4089);
nand U6064 (N_6064,N_3783,N_2786);
and U6065 (N_6065,N_2850,N_4605);
nand U6066 (N_6066,N_3090,N_2857);
xnor U6067 (N_6067,N_3155,N_2832);
nand U6068 (N_6068,N_3166,N_2977);
nor U6069 (N_6069,N_2629,N_3721);
and U6070 (N_6070,N_3889,N_2876);
or U6071 (N_6071,N_4176,N_2761);
nor U6072 (N_6072,N_4692,N_4332);
nand U6073 (N_6073,N_2578,N_2877);
and U6074 (N_6074,N_3503,N_2723);
or U6075 (N_6075,N_3173,N_3233);
nor U6076 (N_6076,N_4446,N_3782);
nor U6077 (N_6077,N_3536,N_4652);
and U6078 (N_6078,N_4925,N_3271);
nor U6079 (N_6079,N_3677,N_2954);
or U6080 (N_6080,N_3816,N_2742);
nor U6081 (N_6081,N_4345,N_3891);
nand U6082 (N_6082,N_3858,N_2733);
xor U6083 (N_6083,N_4821,N_3881);
and U6084 (N_6084,N_2796,N_3641);
nor U6085 (N_6085,N_2594,N_2973);
nor U6086 (N_6086,N_3060,N_3996);
and U6087 (N_6087,N_2618,N_2739);
nand U6088 (N_6088,N_2577,N_3747);
nand U6089 (N_6089,N_4146,N_3622);
nand U6090 (N_6090,N_3062,N_2512);
xor U6091 (N_6091,N_3591,N_2917);
nor U6092 (N_6092,N_3956,N_4691);
or U6093 (N_6093,N_4317,N_2643);
nor U6094 (N_6094,N_3145,N_3365);
or U6095 (N_6095,N_2589,N_3044);
xnor U6096 (N_6096,N_4298,N_4915);
nor U6097 (N_6097,N_4205,N_3238);
or U6098 (N_6098,N_4424,N_3003);
or U6099 (N_6099,N_4060,N_2711);
nand U6100 (N_6100,N_4890,N_3224);
nor U6101 (N_6101,N_2754,N_4975);
nor U6102 (N_6102,N_3370,N_3729);
nor U6103 (N_6103,N_4314,N_4208);
nor U6104 (N_6104,N_4471,N_3560);
nor U6105 (N_6105,N_3004,N_2646);
or U6106 (N_6106,N_4405,N_4891);
and U6107 (N_6107,N_4248,N_2925);
nor U6108 (N_6108,N_4289,N_4409);
nand U6109 (N_6109,N_3247,N_4572);
xor U6110 (N_6110,N_3262,N_4829);
and U6111 (N_6111,N_4352,N_2937);
and U6112 (N_6112,N_3115,N_4313);
nand U6113 (N_6113,N_3508,N_2882);
and U6114 (N_6114,N_4462,N_3623);
xor U6115 (N_6115,N_2878,N_4721);
nor U6116 (N_6116,N_4143,N_3130);
xnor U6117 (N_6117,N_4549,N_2685);
and U6118 (N_6118,N_3218,N_4942);
nand U6119 (N_6119,N_3546,N_2736);
nor U6120 (N_6120,N_3092,N_3431);
nand U6121 (N_6121,N_3567,N_4538);
and U6122 (N_6122,N_2941,N_3124);
nor U6123 (N_6123,N_3071,N_3903);
nor U6124 (N_6124,N_4544,N_2568);
or U6125 (N_6125,N_3416,N_4155);
nand U6126 (N_6126,N_3709,N_4861);
and U6127 (N_6127,N_2905,N_3441);
nand U6128 (N_6128,N_3272,N_3408);
nor U6129 (N_6129,N_4685,N_2619);
xor U6130 (N_6130,N_3564,N_4038);
or U6131 (N_6131,N_4660,N_3968);
xnor U6132 (N_6132,N_4353,N_3111);
nand U6133 (N_6133,N_3136,N_3899);
xor U6134 (N_6134,N_4864,N_4226);
xor U6135 (N_6135,N_4269,N_2943);
and U6136 (N_6136,N_2674,N_3340);
and U6137 (N_6137,N_2683,N_3000);
and U6138 (N_6138,N_3142,N_4140);
and U6139 (N_6139,N_4383,N_3446);
xnor U6140 (N_6140,N_3862,N_3012);
and U6141 (N_6141,N_3883,N_3592);
nor U6142 (N_6142,N_4158,N_3882);
or U6143 (N_6143,N_2686,N_2695);
or U6144 (N_6144,N_3114,N_4275);
xor U6145 (N_6145,N_4276,N_3072);
or U6146 (N_6146,N_2996,N_4846);
xor U6147 (N_6147,N_3819,N_4522);
xnor U6148 (N_6148,N_3316,N_3353);
nand U6149 (N_6149,N_4480,N_2757);
and U6150 (N_6150,N_3485,N_4938);
xnor U6151 (N_6151,N_4127,N_3957);
or U6152 (N_6152,N_2903,N_2947);
or U6153 (N_6153,N_3118,N_4418);
xor U6154 (N_6154,N_3445,N_2781);
xnor U6155 (N_6155,N_3047,N_4233);
or U6156 (N_6156,N_4723,N_3796);
nor U6157 (N_6157,N_3966,N_2718);
xnor U6158 (N_6158,N_4235,N_2604);
or U6159 (N_6159,N_2699,N_2529);
and U6160 (N_6160,N_4123,N_4911);
or U6161 (N_6161,N_4814,N_4568);
and U6162 (N_6162,N_3298,N_4098);
nand U6163 (N_6163,N_4293,N_2569);
and U6164 (N_6164,N_4473,N_2511);
nor U6165 (N_6165,N_2545,N_4227);
nand U6166 (N_6166,N_4410,N_4440);
and U6167 (N_6167,N_2784,N_4219);
and U6168 (N_6168,N_2750,N_2500);
xnor U6169 (N_6169,N_3433,N_4137);
or U6170 (N_6170,N_2721,N_4598);
xnor U6171 (N_6171,N_3910,N_4086);
nand U6172 (N_6172,N_3122,N_3268);
nand U6173 (N_6173,N_3666,N_3066);
nand U6174 (N_6174,N_2966,N_4084);
and U6175 (N_6175,N_3520,N_2570);
nor U6176 (N_6176,N_4128,N_2740);
and U6177 (N_6177,N_4171,N_3859);
nand U6178 (N_6178,N_4768,N_4626);
nand U6179 (N_6179,N_3241,N_4618);
nand U6180 (N_6180,N_2606,N_4217);
xnor U6181 (N_6181,N_4523,N_3715);
or U6182 (N_6182,N_4859,N_2783);
or U6183 (N_6183,N_4095,N_3172);
or U6184 (N_6184,N_3502,N_3655);
nand U6185 (N_6185,N_3602,N_3703);
or U6186 (N_6186,N_4559,N_4812);
or U6187 (N_6187,N_3335,N_4847);
and U6188 (N_6188,N_4324,N_4034);
xor U6189 (N_6189,N_2961,N_3808);
nand U6190 (N_6190,N_3751,N_3231);
and U6191 (N_6191,N_3048,N_3323);
nand U6192 (N_6192,N_3103,N_3870);
or U6193 (N_6193,N_2735,N_3334);
nor U6194 (N_6194,N_3811,N_3737);
xnor U6195 (N_6195,N_4120,N_3106);
nor U6196 (N_6196,N_2891,N_4909);
nor U6197 (N_6197,N_4100,N_4062);
nand U6198 (N_6198,N_4922,N_4296);
and U6199 (N_6199,N_3850,N_4828);
and U6200 (N_6200,N_4542,N_2927);
xnor U6201 (N_6201,N_2667,N_2610);
and U6202 (N_6202,N_2910,N_3790);
nand U6203 (N_6203,N_4845,N_3187);
and U6204 (N_6204,N_4041,N_4979);
nand U6205 (N_6205,N_4050,N_2867);
nand U6206 (N_6206,N_3440,N_4928);
and U6207 (N_6207,N_2887,N_2824);
xor U6208 (N_6208,N_3465,N_3212);
or U6209 (N_6209,N_4788,N_3225);
and U6210 (N_6210,N_4765,N_2769);
or U6211 (N_6211,N_3642,N_4347);
or U6212 (N_6212,N_2668,N_4735);
and U6213 (N_6213,N_3629,N_2776);
nor U6214 (N_6214,N_2848,N_2531);
xor U6215 (N_6215,N_4339,N_3357);
nor U6216 (N_6216,N_3775,N_2843);
or U6217 (N_6217,N_4625,N_3199);
or U6218 (N_6218,N_2886,N_2822);
nand U6219 (N_6219,N_2972,N_2988);
nand U6220 (N_6220,N_3778,N_4030);
xor U6221 (N_6221,N_4042,N_4920);
and U6222 (N_6222,N_3162,N_3705);
or U6223 (N_6223,N_4664,N_4402);
and U6224 (N_6224,N_4201,N_2590);
xnor U6225 (N_6225,N_4368,N_2924);
and U6226 (N_6226,N_3589,N_4285);
and U6227 (N_6227,N_4012,N_3159);
xor U6228 (N_6228,N_2949,N_4811);
and U6229 (N_6229,N_4887,N_2632);
nor U6230 (N_6230,N_2829,N_3454);
xnor U6231 (N_6231,N_3498,N_4865);
nand U6232 (N_6232,N_3070,N_2774);
xor U6233 (N_6233,N_3490,N_3764);
nor U6234 (N_6234,N_2620,N_4921);
or U6235 (N_6235,N_4769,N_3803);
or U6236 (N_6236,N_3707,N_4132);
nor U6237 (N_6237,N_4026,N_3230);
nand U6238 (N_6238,N_4850,N_3781);
nand U6239 (N_6239,N_3309,N_3388);
or U6240 (N_6240,N_3994,N_2671);
xor U6241 (N_6241,N_2841,N_4644);
and U6242 (N_6242,N_4080,N_3027);
or U6243 (N_6243,N_4628,N_4704);
nor U6244 (N_6244,N_4816,N_4113);
and U6245 (N_6245,N_3690,N_3580);
nor U6246 (N_6246,N_3393,N_3752);
xor U6247 (N_6247,N_3437,N_4934);
and U6248 (N_6248,N_2505,N_3313);
nor U6249 (N_6249,N_3097,N_2788);
or U6250 (N_6250,N_4216,N_3868);
or U6251 (N_6251,N_3651,N_4484);
nand U6252 (N_6252,N_3209,N_2772);
or U6253 (N_6253,N_2891,N_4477);
nor U6254 (N_6254,N_2992,N_3930);
nand U6255 (N_6255,N_2583,N_4729);
nand U6256 (N_6256,N_4271,N_4680);
and U6257 (N_6257,N_3579,N_3945);
nand U6258 (N_6258,N_2532,N_3613);
xnor U6259 (N_6259,N_2636,N_3369);
nand U6260 (N_6260,N_2557,N_2578);
nor U6261 (N_6261,N_2725,N_4679);
xnor U6262 (N_6262,N_4218,N_4491);
xor U6263 (N_6263,N_3020,N_4252);
xnor U6264 (N_6264,N_4714,N_3472);
and U6265 (N_6265,N_3931,N_2792);
nand U6266 (N_6266,N_3349,N_3134);
or U6267 (N_6267,N_3705,N_4919);
xor U6268 (N_6268,N_2719,N_4065);
and U6269 (N_6269,N_3183,N_2983);
nor U6270 (N_6270,N_3269,N_3892);
and U6271 (N_6271,N_3273,N_3272);
nand U6272 (N_6272,N_4559,N_4705);
xor U6273 (N_6273,N_3278,N_4428);
or U6274 (N_6274,N_3287,N_2820);
or U6275 (N_6275,N_4029,N_4966);
or U6276 (N_6276,N_3116,N_3066);
or U6277 (N_6277,N_3282,N_2526);
or U6278 (N_6278,N_2926,N_4451);
nand U6279 (N_6279,N_3818,N_2960);
or U6280 (N_6280,N_3579,N_3667);
nor U6281 (N_6281,N_4121,N_4108);
xnor U6282 (N_6282,N_4062,N_4287);
or U6283 (N_6283,N_4205,N_3973);
or U6284 (N_6284,N_4294,N_4124);
or U6285 (N_6285,N_2720,N_3628);
xnor U6286 (N_6286,N_3322,N_4430);
nand U6287 (N_6287,N_4458,N_3163);
xor U6288 (N_6288,N_3474,N_2646);
and U6289 (N_6289,N_2606,N_2940);
and U6290 (N_6290,N_4295,N_4008);
xor U6291 (N_6291,N_4244,N_4589);
xnor U6292 (N_6292,N_3075,N_2896);
nor U6293 (N_6293,N_4256,N_4970);
and U6294 (N_6294,N_4824,N_2643);
xor U6295 (N_6295,N_4910,N_2959);
xor U6296 (N_6296,N_4324,N_4025);
xor U6297 (N_6297,N_3895,N_3814);
and U6298 (N_6298,N_3501,N_3351);
and U6299 (N_6299,N_3919,N_2744);
nand U6300 (N_6300,N_3053,N_4743);
nor U6301 (N_6301,N_2652,N_3454);
xnor U6302 (N_6302,N_4343,N_3890);
nand U6303 (N_6303,N_4612,N_4149);
xor U6304 (N_6304,N_3300,N_4994);
nand U6305 (N_6305,N_3972,N_4157);
or U6306 (N_6306,N_4215,N_2784);
xor U6307 (N_6307,N_4621,N_2894);
or U6308 (N_6308,N_2628,N_4482);
or U6309 (N_6309,N_4187,N_3374);
nand U6310 (N_6310,N_3993,N_3796);
and U6311 (N_6311,N_3137,N_4826);
or U6312 (N_6312,N_2540,N_3948);
xor U6313 (N_6313,N_4034,N_2539);
and U6314 (N_6314,N_4125,N_4882);
and U6315 (N_6315,N_4033,N_2705);
and U6316 (N_6316,N_3235,N_4454);
and U6317 (N_6317,N_4180,N_3670);
xnor U6318 (N_6318,N_4033,N_2584);
and U6319 (N_6319,N_3412,N_4080);
nor U6320 (N_6320,N_3485,N_3704);
nor U6321 (N_6321,N_4865,N_3233);
xnor U6322 (N_6322,N_2902,N_3923);
and U6323 (N_6323,N_4864,N_3689);
nand U6324 (N_6324,N_3981,N_4196);
or U6325 (N_6325,N_3786,N_4336);
nand U6326 (N_6326,N_4545,N_3265);
or U6327 (N_6327,N_4307,N_3580);
xor U6328 (N_6328,N_3181,N_2651);
and U6329 (N_6329,N_4408,N_4413);
nor U6330 (N_6330,N_2755,N_3116);
nand U6331 (N_6331,N_4889,N_4593);
or U6332 (N_6332,N_4609,N_2653);
and U6333 (N_6333,N_4353,N_4817);
xnor U6334 (N_6334,N_4621,N_3712);
nand U6335 (N_6335,N_3501,N_3807);
xnor U6336 (N_6336,N_4237,N_4345);
nor U6337 (N_6337,N_4704,N_4668);
xor U6338 (N_6338,N_3509,N_4225);
nor U6339 (N_6339,N_3785,N_3932);
nor U6340 (N_6340,N_3219,N_4446);
nand U6341 (N_6341,N_3005,N_4368);
nand U6342 (N_6342,N_2931,N_3825);
and U6343 (N_6343,N_2560,N_3872);
xor U6344 (N_6344,N_4634,N_4765);
and U6345 (N_6345,N_4535,N_3094);
nand U6346 (N_6346,N_3016,N_4738);
nor U6347 (N_6347,N_4757,N_4375);
nor U6348 (N_6348,N_4198,N_3641);
xnor U6349 (N_6349,N_3871,N_4903);
nand U6350 (N_6350,N_2967,N_3938);
xor U6351 (N_6351,N_4106,N_4938);
nor U6352 (N_6352,N_4684,N_3323);
and U6353 (N_6353,N_4843,N_3820);
or U6354 (N_6354,N_3359,N_4286);
nor U6355 (N_6355,N_2796,N_4496);
nor U6356 (N_6356,N_3690,N_3914);
and U6357 (N_6357,N_4568,N_4883);
nor U6358 (N_6358,N_4799,N_4182);
or U6359 (N_6359,N_2817,N_3570);
nand U6360 (N_6360,N_2890,N_4754);
and U6361 (N_6361,N_4575,N_3040);
or U6362 (N_6362,N_4408,N_3391);
nand U6363 (N_6363,N_3552,N_3438);
or U6364 (N_6364,N_3908,N_3005);
nor U6365 (N_6365,N_2826,N_3383);
xnor U6366 (N_6366,N_2879,N_3103);
nor U6367 (N_6367,N_4875,N_4792);
xnor U6368 (N_6368,N_4737,N_4189);
and U6369 (N_6369,N_3813,N_4431);
nand U6370 (N_6370,N_3886,N_2883);
nor U6371 (N_6371,N_3392,N_4640);
nor U6372 (N_6372,N_3969,N_2979);
or U6373 (N_6373,N_2681,N_4950);
nor U6374 (N_6374,N_3607,N_3276);
nor U6375 (N_6375,N_3897,N_4031);
nor U6376 (N_6376,N_4786,N_4487);
and U6377 (N_6377,N_3361,N_3140);
xnor U6378 (N_6378,N_4083,N_2934);
or U6379 (N_6379,N_3363,N_3025);
nor U6380 (N_6380,N_3416,N_4308);
nand U6381 (N_6381,N_3478,N_4275);
nor U6382 (N_6382,N_3703,N_4522);
nand U6383 (N_6383,N_3246,N_4907);
nor U6384 (N_6384,N_3458,N_4757);
nor U6385 (N_6385,N_2502,N_4806);
xor U6386 (N_6386,N_4115,N_2527);
or U6387 (N_6387,N_2807,N_4695);
and U6388 (N_6388,N_3640,N_4697);
xnor U6389 (N_6389,N_2763,N_4432);
nor U6390 (N_6390,N_4079,N_3135);
xor U6391 (N_6391,N_4355,N_3085);
nor U6392 (N_6392,N_4855,N_4445);
or U6393 (N_6393,N_4989,N_3804);
nand U6394 (N_6394,N_3724,N_3793);
or U6395 (N_6395,N_3703,N_3010);
xnor U6396 (N_6396,N_3733,N_3096);
nor U6397 (N_6397,N_4498,N_4982);
nor U6398 (N_6398,N_4578,N_4710);
nand U6399 (N_6399,N_2861,N_3140);
xnor U6400 (N_6400,N_2836,N_2506);
xor U6401 (N_6401,N_3018,N_4654);
xnor U6402 (N_6402,N_4572,N_3556);
or U6403 (N_6403,N_4022,N_3405);
nor U6404 (N_6404,N_4677,N_3750);
or U6405 (N_6405,N_2595,N_4680);
and U6406 (N_6406,N_4503,N_2664);
or U6407 (N_6407,N_2879,N_3892);
nor U6408 (N_6408,N_3935,N_4317);
nor U6409 (N_6409,N_4285,N_3717);
and U6410 (N_6410,N_4731,N_3283);
or U6411 (N_6411,N_2551,N_3644);
or U6412 (N_6412,N_4359,N_4733);
or U6413 (N_6413,N_3031,N_4836);
xnor U6414 (N_6414,N_3905,N_4100);
nor U6415 (N_6415,N_3010,N_3486);
or U6416 (N_6416,N_3038,N_3879);
xor U6417 (N_6417,N_3266,N_3457);
or U6418 (N_6418,N_3414,N_2518);
or U6419 (N_6419,N_4294,N_4724);
xor U6420 (N_6420,N_2668,N_3815);
or U6421 (N_6421,N_2517,N_3240);
nor U6422 (N_6422,N_3189,N_4527);
xor U6423 (N_6423,N_3283,N_4844);
and U6424 (N_6424,N_4320,N_3195);
xnor U6425 (N_6425,N_3975,N_4890);
or U6426 (N_6426,N_4652,N_3226);
and U6427 (N_6427,N_2782,N_4797);
xnor U6428 (N_6428,N_3183,N_3948);
nor U6429 (N_6429,N_4796,N_3507);
xnor U6430 (N_6430,N_3556,N_3618);
or U6431 (N_6431,N_4236,N_3948);
nor U6432 (N_6432,N_3476,N_3395);
and U6433 (N_6433,N_3458,N_4408);
xor U6434 (N_6434,N_3759,N_2667);
xor U6435 (N_6435,N_3665,N_3447);
nor U6436 (N_6436,N_3028,N_3647);
and U6437 (N_6437,N_3241,N_2719);
nor U6438 (N_6438,N_3080,N_2797);
nand U6439 (N_6439,N_3909,N_3233);
xnor U6440 (N_6440,N_4443,N_4125);
or U6441 (N_6441,N_4273,N_4937);
nor U6442 (N_6442,N_4276,N_4509);
and U6443 (N_6443,N_4634,N_2916);
nor U6444 (N_6444,N_4828,N_4242);
nor U6445 (N_6445,N_2810,N_3914);
nor U6446 (N_6446,N_4622,N_3710);
xnor U6447 (N_6447,N_4361,N_4228);
xnor U6448 (N_6448,N_3100,N_3878);
and U6449 (N_6449,N_4895,N_4438);
or U6450 (N_6450,N_4971,N_3208);
xnor U6451 (N_6451,N_4876,N_2746);
nor U6452 (N_6452,N_3626,N_4249);
or U6453 (N_6453,N_2542,N_4617);
or U6454 (N_6454,N_4553,N_4323);
or U6455 (N_6455,N_4658,N_3963);
xor U6456 (N_6456,N_3056,N_4515);
and U6457 (N_6457,N_4083,N_3302);
xnor U6458 (N_6458,N_2774,N_3013);
nor U6459 (N_6459,N_2780,N_3510);
nor U6460 (N_6460,N_4115,N_3140);
and U6461 (N_6461,N_4422,N_4972);
or U6462 (N_6462,N_3444,N_4343);
and U6463 (N_6463,N_4790,N_3330);
or U6464 (N_6464,N_3141,N_3655);
nor U6465 (N_6465,N_4886,N_2514);
nor U6466 (N_6466,N_2544,N_2909);
or U6467 (N_6467,N_4497,N_2773);
nand U6468 (N_6468,N_4656,N_2949);
xor U6469 (N_6469,N_2586,N_3709);
or U6470 (N_6470,N_2981,N_4539);
and U6471 (N_6471,N_3840,N_3781);
nor U6472 (N_6472,N_3344,N_4718);
and U6473 (N_6473,N_4975,N_4745);
and U6474 (N_6474,N_2580,N_4849);
xnor U6475 (N_6475,N_3701,N_2875);
xor U6476 (N_6476,N_4478,N_4951);
nand U6477 (N_6477,N_4711,N_3504);
nand U6478 (N_6478,N_2777,N_4777);
nand U6479 (N_6479,N_2827,N_4460);
nand U6480 (N_6480,N_2927,N_2587);
and U6481 (N_6481,N_2745,N_3996);
nand U6482 (N_6482,N_3803,N_4739);
or U6483 (N_6483,N_3278,N_3165);
xnor U6484 (N_6484,N_3355,N_4545);
or U6485 (N_6485,N_4035,N_3240);
nor U6486 (N_6486,N_3383,N_4928);
nor U6487 (N_6487,N_3525,N_3980);
nand U6488 (N_6488,N_4547,N_4040);
nand U6489 (N_6489,N_4831,N_3957);
nand U6490 (N_6490,N_4879,N_2527);
nor U6491 (N_6491,N_2589,N_2686);
or U6492 (N_6492,N_3329,N_3424);
nand U6493 (N_6493,N_3829,N_4199);
xnor U6494 (N_6494,N_4754,N_4835);
nand U6495 (N_6495,N_4905,N_3958);
xnor U6496 (N_6496,N_4214,N_3572);
xor U6497 (N_6497,N_4910,N_4758);
xnor U6498 (N_6498,N_3769,N_4501);
nor U6499 (N_6499,N_3520,N_2808);
nand U6500 (N_6500,N_2599,N_4422);
xor U6501 (N_6501,N_3505,N_3551);
and U6502 (N_6502,N_3721,N_2750);
nand U6503 (N_6503,N_3831,N_3595);
and U6504 (N_6504,N_4820,N_3357);
nand U6505 (N_6505,N_3081,N_3764);
nor U6506 (N_6506,N_3826,N_2883);
nand U6507 (N_6507,N_3389,N_4537);
nand U6508 (N_6508,N_3724,N_3884);
xnor U6509 (N_6509,N_2531,N_3659);
nor U6510 (N_6510,N_2556,N_4053);
xor U6511 (N_6511,N_4856,N_4840);
xnor U6512 (N_6512,N_2940,N_4283);
xor U6513 (N_6513,N_4080,N_4287);
or U6514 (N_6514,N_4594,N_4739);
and U6515 (N_6515,N_3388,N_2512);
xor U6516 (N_6516,N_3935,N_3207);
or U6517 (N_6517,N_3648,N_4835);
xnor U6518 (N_6518,N_2520,N_4959);
nand U6519 (N_6519,N_4133,N_4489);
nor U6520 (N_6520,N_4091,N_4221);
nand U6521 (N_6521,N_3874,N_4462);
and U6522 (N_6522,N_2583,N_4811);
or U6523 (N_6523,N_3924,N_2998);
nor U6524 (N_6524,N_4908,N_4014);
xnor U6525 (N_6525,N_2818,N_4921);
and U6526 (N_6526,N_3814,N_3533);
nand U6527 (N_6527,N_2987,N_4116);
and U6528 (N_6528,N_3062,N_4109);
and U6529 (N_6529,N_3390,N_4683);
nor U6530 (N_6530,N_3815,N_3582);
nand U6531 (N_6531,N_3012,N_2724);
nand U6532 (N_6532,N_4263,N_4054);
nand U6533 (N_6533,N_4806,N_4070);
xnor U6534 (N_6534,N_3135,N_3371);
xor U6535 (N_6535,N_3897,N_3485);
xor U6536 (N_6536,N_3124,N_2628);
xor U6537 (N_6537,N_3434,N_2919);
nand U6538 (N_6538,N_4859,N_4001);
nand U6539 (N_6539,N_3073,N_4630);
xnor U6540 (N_6540,N_4451,N_2811);
nand U6541 (N_6541,N_3235,N_4735);
nor U6542 (N_6542,N_4464,N_4971);
xor U6543 (N_6543,N_3131,N_2764);
or U6544 (N_6544,N_3336,N_3945);
nand U6545 (N_6545,N_4544,N_2562);
and U6546 (N_6546,N_2532,N_4531);
and U6547 (N_6547,N_3104,N_3729);
nor U6548 (N_6548,N_2959,N_4648);
nor U6549 (N_6549,N_3351,N_4890);
and U6550 (N_6550,N_4331,N_4310);
and U6551 (N_6551,N_4518,N_4672);
nand U6552 (N_6552,N_3662,N_2528);
nor U6553 (N_6553,N_3997,N_3727);
nor U6554 (N_6554,N_3454,N_4335);
xnor U6555 (N_6555,N_3646,N_4519);
and U6556 (N_6556,N_4298,N_3054);
or U6557 (N_6557,N_4584,N_3319);
xor U6558 (N_6558,N_4136,N_3189);
nor U6559 (N_6559,N_3610,N_3310);
nand U6560 (N_6560,N_4427,N_3795);
and U6561 (N_6561,N_3410,N_3556);
or U6562 (N_6562,N_4449,N_3321);
nor U6563 (N_6563,N_4306,N_4270);
nand U6564 (N_6564,N_2677,N_4848);
nor U6565 (N_6565,N_2537,N_2678);
nor U6566 (N_6566,N_4321,N_3326);
nor U6567 (N_6567,N_3113,N_4394);
and U6568 (N_6568,N_4041,N_3166);
nand U6569 (N_6569,N_2520,N_3996);
or U6570 (N_6570,N_4734,N_4756);
nor U6571 (N_6571,N_3387,N_4038);
and U6572 (N_6572,N_3571,N_4751);
or U6573 (N_6573,N_3347,N_2765);
nand U6574 (N_6574,N_2590,N_3930);
xor U6575 (N_6575,N_3011,N_4470);
and U6576 (N_6576,N_4034,N_3843);
and U6577 (N_6577,N_4400,N_2751);
nor U6578 (N_6578,N_3774,N_3095);
xnor U6579 (N_6579,N_4436,N_4008);
nor U6580 (N_6580,N_2575,N_3610);
xor U6581 (N_6581,N_3432,N_4618);
or U6582 (N_6582,N_2864,N_3245);
and U6583 (N_6583,N_2665,N_4102);
nand U6584 (N_6584,N_4429,N_3035);
nand U6585 (N_6585,N_2578,N_4477);
nand U6586 (N_6586,N_4784,N_2912);
and U6587 (N_6587,N_2990,N_3246);
nand U6588 (N_6588,N_4853,N_3678);
xnor U6589 (N_6589,N_4444,N_4308);
and U6590 (N_6590,N_2551,N_2895);
nor U6591 (N_6591,N_4907,N_2733);
and U6592 (N_6592,N_4764,N_3944);
xor U6593 (N_6593,N_4004,N_3917);
or U6594 (N_6594,N_4733,N_3174);
xor U6595 (N_6595,N_2866,N_3303);
and U6596 (N_6596,N_2955,N_4170);
xor U6597 (N_6597,N_4644,N_2557);
xor U6598 (N_6598,N_2659,N_2901);
and U6599 (N_6599,N_2857,N_2937);
and U6600 (N_6600,N_3951,N_3061);
nand U6601 (N_6601,N_2709,N_4202);
nand U6602 (N_6602,N_4029,N_3190);
xnor U6603 (N_6603,N_4071,N_4277);
or U6604 (N_6604,N_4413,N_4489);
or U6605 (N_6605,N_3295,N_4388);
and U6606 (N_6606,N_4371,N_2785);
nor U6607 (N_6607,N_4887,N_3663);
and U6608 (N_6608,N_2705,N_4848);
or U6609 (N_6609,N_2541,N_4809);
or U6610 (N_6610,N_4146,N_4997);
or U6611 (N_6611,N_4753,N_2614);
or U6612 (N_6612,N_4046,N_3664);
or U6613 (N_6613,N_2949,N_3725);
and U6614 (N_6614,N_3368,N_4147);
or U6615 (N_6615,N_3918,N_3443);
nor U6616 (N_6616,N_4689,N_4813);
xnor U6617 (N_6617,N_2598,N_3362);
and U6618 (N_6618,N_4433,N_4432);
nor U6619 (N_6619,N_2717,N_3822);
nand U6620 (N_6620,N_3318,N_4209);
xor U6621 (N_6621,N_2874,N_4926);
nor U6622 (N_6622,N_3450,N_3716);
xor U6623 (N_6623,N_4266,N_2637);
nand U6624 (N_6624,N_4109,N_4104);
or U6625 (N_6625,N_2975,N_3172);
or U6626 (N_6626,N_3960,N_3911);
nand U6627 (N_6627,N_3488,N_4335);
xor U6628 (N_6628,N_2962,N_4860);
and U6629 (N_6629,N_3695,N_2511);
nor U6630 (N_6630,N_3617,N_2613);
or U6631 (N_6631,N_4988,N_3468);
nand U6632 (N_6632,N_4891,N_4430);
xnor U6633 (N_6633,N_3505,N_4555);
nor U6634 (N_6634,N_4848,N_4183);
nor U6635 (N_6635,N_3547,N_3021);
and U6636 (N_6636,N_2786,N_3215);
and U6637 (N_6637,N_4803,N_3837);
nor U6638 (N_6638,N_2875,N_4970);
nand U6639 (N_6639,N_2787,N_4161);
nand U6640 (N_6640,N_4058,N_3812);
xnor U6641 (N_6641,N_2911,N_3816);
and U6642 (N_6642,N_2561,N_3732);
nor U6643 (N_6643,N_3669,N_2610);
nor U6644 (N_6644,N_4346,N_3287);
and U6645 (N_6645,N_3318,N_3963);
or U6646 (N_6646,N_4828,N_3572);
xor U6647 (N_6647,N_4820,N_2940);
or U6648 (N_6648,N_2790,N_2752);
and U6649 (N_6649,N_3164,N_4699);
and U6650 (N_6650,N_3169,N_4753);
or U6651 (N_6651,N_4171,N_4760);
xnor U6652 (N_6652,N_4764,N_3269);
nor U6653 (N_6653,N_3789,N_2628);
nor U6654 (N_6654,N_4368,N_3541);
xnor U6655 (N_6655,N_4365,N_3525);
or U6656 (N_6656,N_2954,N_4275);
or U6657 (N_6657,N_2822,N_4079);
and U6658 (N_6658,N_4631,N_3332);
nor U6659 (N_6659,N_2563,N_2907);
and U6660 (N_6660,N_3123,N_3267);
nor U6661 (N_6661,N_4077,N_4553);
and U6662 (N_6662,N_4426,N_2532);
nor U6663 (N_6663,N_4487,N_2508);
or U6664 (N_6664,N_2794,N_3178);
or U6665 (N_6665,N_3925,N_2914);
nor U6666 (N_6666,N_3284,N_4296);
nor U6667 (N_6667,N_3066,N_3528);
or U6668 (N_6668,N_4573,N_3743);
and U6669 (N_6669,N_3974,N_4084);
and U6670 (N_6670,N_4609,N_3563);
nor U6671 (N_6671,N_4240,N_3878);
nor U6672 (N_6672,N_4895,N_4931);
nand U6673 (N_6673,N_2779,N_4574);
nand U6674 (N_6674,N_4975,N_2773);
nand U6675 (N_6675,N_3016,N_4384);
nor U6676 (N_6676,N_4524,N_4344);
and U6677 (N_6677,N_2951,N_4441);
and U6678 (N_6678,N_4239,N_3929);
xor U6679 (N_6679,N_4385,N_4606);
nand U6680 (N_6680,N_3609,N_4389);
xnor U6681 (N_6681,N_4467,N_4854);
or U6682 (N_6682,N_4298,N_3115);
and U6683 (N_6683,N_3575,N_4684);
or U6684 (N_6684,N_3741,N_3915);
nand U6685 (N_6685,N_3062,N_4114);
nand U6686 (N_6686,N_2790,N_2690);
nor U6687 (N_6687,N_3284,N_4521);
nor U6688 (N_6688,N_4387,N_2550);
or U6689 (N_6689,N_3915,N_3746);
xor U6690 (N_6690,N_2642,N_2618);
xnor U6691 (N_6691,N_4007,N_4993);
nor U6692 (N_6692,N_3640,N_2648);
or U6693 (N_6693,N_4688,N_4747);
or U6694 (N_6694,N_4568,N_4244);
or U6695 (N_6695,N_3548,N_2958);
nor U6696 (N_6696,N_2649,N_3490);
nand U6697 (N_6697,N_4754,N_2761);
nor U6698 (N_6698,N_4197,N_3008);
xor U6699 (N_6699,N_3239,N_3371);
nand U6700 (N_6700,N_3890,N_2636);
nand U6701 (N_6701,N_2829,N_3865);
or U6702 (N_6702,N_4565,N_3135);
and U6703 (N_6703,N_4499,N_4031);
or U6704 (N_6704,N_2553,N_3154);
nand U6705 (N_6705,N_3272,N_2555);
or U6706 (N_6706,N_3523,N_4202);
and U6707 (N_6707,N_4956,N_4790);
nand U6708 (N_6708,N_3137,N_4243);
xor U6709 (N_6709,N_2728,N_3639);
and U6710 (N_6710,N_2547,N_4731);
and U6711 (N_6711,N_4106,N_3575);
nand U6712 (N_6712,N_4549,N_2610);
and U6713 (N_6713,N_4861,N_2726);
and U6714 (N_6714,N_4775,N_2798);
xor U6715 (N_6715,N_3269,N_3999);
xnor U6716 (N_6716,N_2912,N_3037);
or U6717 (N_6717,N_3592,N_3368);
nor U6718 (N_6718,N_3109,N_3401);
and U6719 (N_6719,N_2660,N_3267);
nor U6720 (N_6720,N_3645,N_4272);
xor U6721 (N_6721,N_4175,N_3516);
xnor U6722 (N_6722,N_2909,N_2605);
nand U6723 (N_6723,N_2547,N_3223);
or U6724 (N_6724,N_4902,N_3488);
nor U6725 (N_6725,N_3345,N_2829);
and U6726 (N_6726,N_2711,N_3837);
nor U6727 (N_6727,N_4702,N_3391);
or U6728 (N_6728,N_4004,N_3236);
nand U6729 (N_6729,N_2979,N_2737);
and U6730 (N_6730,N_3993,N_4632);
nor U6731 (N_6731,N_4875,N_4422);
nor U6732 (N_6732,N_2576,N_3474);
xor U6733 (N_6733,N_3145,N_2707);
or U6734 (N_6734,N_3445,N_4464);
nor U6735 (N_6735,N_3401,N_3411);
nor U6736 (N_6736,N_2613,N_3730);
and U6737 (N_6737,N_4627,N_3888);
nand U6738 (N_6738,N_4348,N_3992);
or U6739 (N_6739,N_2621,N_4616);
xor U6740 (N_6740,N_4251,N_4602);
nand U6741 (N_6741,N_4177,N_2680);
and U6742 (N_6742,N_2724,N_3938);
and U6743 (N_6743,N_3949,N_3399);
nand U6744 (N_6744,N_2718,N_4564);
and U6745 (N_6745,N_3586,N_3801);
xnor U6746 (N_6746,N_3086,N_3392);
nor U6747 (N_6747,N_4169,N_3159);
and U6748 (N_6748,N_3522,N_2792);
and U6749 (N_6749,N_4944,N_2525);
nor U6750 (N_6750,N_3179,N_3898);
xnor U6751 (N_6751,N_4784,N_2539);
and U6752 (N_6752,N_3886,N_3812);
and U6753 (N_6753,N_2715,N_3272);
xnor U6754 (N_6754,N_2788,N_3688);
or U6755 (N_6755,N_4870,N_3927);
or U6756 (N_6756,N_3196,N_3398);
and U6757 (N_6757,N_2981,N_2552);
nand U6758 (N_6758,N_2604,N_4378);
nand U6759 (N_6759,N_4663,N_2820);
nor U6760 (N_6760,N_3426,N_2507);
xnor U6761 (N_6761,N_4373,N_3795);
nor U6762 (N_6762,N_4270,N_4530);
nand U6763 (N_6763,N_4337,N_4001);
nand U6764 (N_6764,N_3144,N_2859);
and U6765 (N_6765,N_2808,N_3652);
nor U6766 (N_6766,N_4966,N_4205);
and U6767 (N_6767,N_4899,N_3992);
nand U6768 (N_6768,N_3901,N_3380);
or U6769 (N_6769,N_3541,N_4077);
or U6770 (N_6770,N_4546,N_3117);
nor U6771 (N_6771,N_4360,N_4192);
nor U6772 (N_6772,N_2926,N_4258);
or U6773 (N_6773,N_4979,N_2983);
and U6774 (N_6774,N_3772,N_4010);
nor U6775 (N_6775,N_4228,N_3804);
nor U6776 (N_6776,N_4877,N_3316);
and U6777 (N_6777,N_2654,N_3925);
or U6778 (N_6778,N_4076,N_3871);
or U6779 (N_6779,N_4244,N_3807);
xnor U6780 (N_6780,N_2951,N_4295);
or U6781 (N_6781,N_4968,N_4509);
and U6782 (N_6782,N_4761,N_4122);
nand U6783 (N_6783,N_4136,N_2901);
nor U6784 (N_6784,N_3264,N_4343);
and U6785 (N_6785,N_4329,N_4590);
nand U6786 (N_6786,N_4494,N_3991);
nor U6787 (N_6787,N_4901,N_3172);
or U6788 (N_6788,N_4820,N_3359);
xnor U6789 (N_6789,N_3668,N_3305);
and U6790 (N_6790,N_4298,N_2812);
nor U6791 (N_6791,N_3212,N_3555);
and U6792 (N_6792,N_3394,N_3847);
nor U6793 (N_6793,N_4802,N_4607);
nor U6794 (N_6794,N_2992,N_2765);
xor U6795 (N_6795,N_4152,N_3143);
and U6796 (N_6796,N_3271,N_3900);
nor U6797 (N_6797,N_2544,N_2727);
nor U6798 (N_6798,N_3907,N_4715);
nor U6799 (N_6799,N_2921,N_4522);
nand U6800 (N_6800,N_4613,N_3881);
and U6801 (N_6801,N_4315,N_2924);
nand U6802 (N_6802,N_3221,N_4686);
or U6803 (N_6803,N_2906,N_2674);
xor U6804 (N_6804,N_3372,N_2968);
nand U6805 (N_6805,N_4049,N_4437);
nand U6806 (N_6806,N_3682,N_3987);
and U6807 (N_6807,N_2683,N_3646);
and U6808 (N_6808,N_3268,N_4975);
xnor U6809 (N_6809,N_4536,N_2686);
and U6810 (N_6810,N_3027,N_4887);
nand U6811 (N_6811,N_3971,N_3155);
xor U6812 (N_6812,N_4859,N_4164);
and U6813 (N_6813,N_4952,N_2845);
nor U6814 (N_6814,N_3401,N_2517);
nand U6815 (N_6815,N_3311,N_2551);
or U6816 (N_6816,N_3797,N_3437);
nor U6817 (N_6817,N_2879,N_3802);
nor U6818 (N_6818,N_2878,N_3837);
or U6819 (N_6819,N_3653,N_2842);
xor U6820 (N_6820,N_2792,N_2658);
nand U6821 (N_6821,N_3133,N_4389);
and U6822 (N_6822,N_4442,N_4166);
nand U6823 (N_6823,N_2873,N_4821);
nor U6824 (N_6824,N_2847,N_3953);
or U6825 (N_6825,N_3762,N_2604);
or U6826 (N_6826,N_3220,N_4136);
nor U6827 (N_6827,N_3470,N_3380);
nand U6828 (N_6828,N_4872,N_4119);
and U6829 (N_6829,N_3113,N_4402);
or U6830 (N_6830,N_3618,N_3913);
nand U6831 (N_6831,N_3300,N_3083);
and U6832 (N_6832,N_4792,N_2568);
nor U6833 (N_6833,N_3424,N_2612);
nor U6834 (N_6834,N_3623,N_3239);
nand U6835 (N_6835,N_4600,N_3101);
and U6836 (N_6836,N_4115,N_4436);
or U6837 (N_6837,N_4546,N_2593);
nand U6838 (N_6838,N_2706,N_3255);
or U6839 (N_6839,N_3631,N_3373);
and U6840 (N_6840,N_2512,N_4116);
and U6841 (N_6841,N_3205,N_2585);
nor U6842 (N_6842,N_4590,N_4723);
nand U6843 (N_6843,N_2617,N_3242);
or U6844 (N_6844,N_2966,N_3542);
xor U6845 (N_6845,N_4749,N_3607);
or U6846 (N_6846,N_3857,N_4466);
nor U6847 (N_6847,N_3588,N_3162);
or U6848 (N_6848,N_4069,N_3256);
nor U6849 (N_6849,N_2868,N_2979);
nand U6850 (N_6850,N_4653,N_3522);
xor U6851 (N_6851,N_3921,N_2642);
or U6852 (N_6852,N_3879,N_3714);
xnor U6853 (N_6853,N_3777,N_4102);
xor U6854 (N_6854,N_4747,N_4810);
nand U6855 (N_6855,N_3134,N_4848);
nand U6856 (N_6856,N_2874,N_4840);
and U6857 (N_6857,N_4851,N_4573);
xor U6858 (N_6858,N_3213,N_3087);
or U6859 (N_6859,N_3454,N_3568);
nor U6860 (N_6860,N_4973,N_4517);
xnor U6861 (N_6861,N_4698,N_2948);
and U6862 (N_6862,N_3386,N_3224);
nand U6863 (N_6863,N_4087,N_2606);
and U6864 (N_6864,N_3235,N_3687);
and U6865 (N_6865,N_4456,N_4306);
nor U6866 (N_6866,N_4863,N_2581);
or U6867 (N_6867,N_4543,N_3477);
and U6868 (N_6868,N_2610,N_3453);
xnor U6869 (N_6869,N_3628,N_3078);
and U6870 (N_6870,N_2757,N_3891);
xor U6871 (N_6871,N_3355,N_4038);
xnor U6872 (N_6872,N_4802,N_4870);
xor U6873 (N_6873,N_3035,N_3591);
nor U6874 (N_6874,N_3138,N_2622);
xnor U6875 (N_6875,N_3913,N_3724);
and U6876 (N_6876,N_4166,N_3447);
nand U6877 (N_6877,N_4802,N_3779);
nor U6878 (N_6878,N_3009,N_4035);
and U6879 (N_6879,N_4280,N_4687);
xnor U6880 (N_6880,N_2939,N_2768);
or U6881 (N_6881,N_3287,N_3636);
nor U6882 (N_6882,N_4237,N_4496);
or U6883 (N_6883,N_3913,N_3243);
and U6884 (N_6884,N_3752,N_3320);
xnor U6885 (N_6885,N_3932,N_4534);
nor U6886 (N_6886,N_4885,N_3194);
xnor U6887 (N_6887,N_3797,N_4995);
nor U6888 (N_6888,N_2633,N_4412);
or U6889 (N_6889,N_3105,N_3306);
nor U6890 (N_6890,N_4711,N_3733);
xnor U6891 (N_6891,N_3000,N_4947);
nor U6892 (N_6892,N_4519,N_4276);
xor U6893 (N_6893,N_3823,N_3684);
and U6894 (N_6894,N_3141,N_3637);
nor U6895 (N_6895,N_3971,N_3582);
or U6896 (N_6896,N_3008,N_4412);
nand U6897 (N_6897,N_3275,N_3957);
nor U6898 (N_6898,N_3819,N_2966);
nand U6899 (N_6899,N_2530,N_4006);
or U6900 (N_6900,N_3327,N_4155);
nor U6901 (N_6901,N_4181,N_3409);
and U6902 (N_6902,N_2896,N_4964);
xnor U6903 (N_6903,N_3497,N_4234);
nand U6904 (N_6904,N_4931,N_2882);
and U6905 (N_6905,N_3287,N_2613);
or U6906 (N_6906,N_2644,N_3925);
nand U6907 (N_6907,N_2857,N_4057);
and U6908 (N_6908,N_3119,N_4530);
nand U6909 (N_6909,N_4957,N_4733);
and U6910 (N_6910,N_3251,N_4041);
nand U6911 (N_6911,N_3563,N_3176);
xnor U6912 (N_6912,N_4146,N_3280);
nor U6913 (N_6913,N_4756,N_3927);
nor U6914 (N_6914,N_3162,N_3730);
or U6915 (N_6915,N_4126,N_4155);
and U6916 (N_6916,N_4281,N_2861);
nand U6917 (N_6917,N_3161,N_3750);
and U6918 (N_6918,N_3878,N_4825);
xnor U6919 (N_6919,N_2847,N_4731);
nand U6920 (N_6920,N_3024,N_4102);
xor U6921 (N_6921,N_2796,N_3194);
nand U6922 (N_6922,N_4884,N_4590);
xor U6923 (N_6923,N_3671,N_3779);
nor U6924 (N_6924,N_3005,N_2907);
xnor U6925 (N_6925,N_3431,N_2604);
or U6926 (N_6926,N_4693,N_4805);
xnor U6927 (N_6927,N_4359,N_3321);
nand U6928 (N_6928,N_3831,N_3289);
nand U6929 (N_6929,N_4032,N_2636);
nand U6930 (N_6930,N_3572,N_4768);
xor U6931 (N_6931,N_4421,N_4833);
nor U6932 (N_6932,N_2913,N_2595);
and U6933 (N_6933,N_3640,N_4448);
or U6934 (N_6934,N_2993,N_3985);
nand U6935 (N_6935,N_3076,N_4317);
nand U6936 (N_6936,N_3445,N_4836);
nand U6937 (N_6937,N_2714,N_3286);
xnor U6938 (N_6938,N_4474,N_2826);
nor U6939 (N_6939,N_4648,N_3010);
and U6940 (N_6940,N_2788,N_2696);
or U6941 (N_6941,N_4501,N_3300);
xnor U6942 (N_6942,N_3356,N_3426);
and U6943 (N_6943,N_3295,N_2745);
nor U6944 (N_6944,N_3147,N_4915);
xor U6945 (N_6945,N_3525,N_4932);
nor U6946 (N_6946,N_4152,N_4081);
and U6947 (N_6947,N_3113,N_2635);
xnor U6948 (N_6948,N_3491,N_3931);
or U6949 (N_6949,N_2920,N_3872);
nor U6950 (N_6950,N_3493,N_4138);
xnor U6951 (N_6951,N_3470,N_3933);
nor U6952 (N_6952,N_3998,N_4865);
or U6953 (N_6953,N_2603,N_3520);
and U6954 (N_6954,N_2806,N_4146);
nand U6955 (N_6955,N_2947,N_3695);
nor U6956 (N_6956,N_4612,N_3896);
or U6957 (N_6957,N_3099,N_3774);
nor U6958 (N_6958,N_2908,N_4483);
nor U6959 (N_6959,N_4290,N_4863);
nor U6960 (N_6960,N_2950,N_4235);
or U6961 (N_6961,N_3827,N_3752);
or U6962 (N_6962,N_2827,N_4205);
nand U6963 (N_6963,N_4597,N_4133);
nor U6964 (N_6964,N_2729,N_2509);
and U6965 (N_6965,N_2791,N_3107);
or U6966 (N_6966,N_3806,N_2715);
xor U6967 (N_6967,N_3949,N_4450);
and U6968 (N_6968,N_4200,N_4189);
and U6969 (N_6969,N_4046,N_4007);
and U6970 (N_6970,N_4352,N_4133);
xnor U6971 (N_6971,N_4868,N_3827);
and U6972 (N_6972,N_3315,N_3807);
or U6973 (N_6973,N_3632,N_2928);
nand U6974 (N_6974,N_4339,N_3395);
nor U6975 (N_6975,N_4111,N_3715);
nand U6976 (N_6976,N_4293,N_3262);
or U6977 (N_6977,N_4899,N_4549);
xor U6978 (N_6978,N_3859,N_3088);
xnor U6979 (N_6979,N_4273,N_4796);
xor U6980 (N_6980,N_4244,N_3441);
xnor U6981 (N_6981,N_2513,N_3974);
xnor U6982 (N_6982,N_4604,N_2540);
nand U6983 (N_6983,N_2876,N_4004);
nand U6984 (N_6984,N_4779,N_4643);
xor U6985 (N_6985,N_4994,N_4707);
or U6986 (N_6986,N_4945,N_4077);
and U6987 (N_6987,N_4187,N_4201);
or U6988 (N_6988,N_4822,N_3931);
and U6989 (N_6989,N_3786,N_4006);
nor U6990 (N_6990,N_3733,N_4765);
nor U6991 (N_6991,N_3268,N_3040);
nor U6992 (N_6992,N_4534,N_2647);
nand U6993 (N_6993,N_2727,N_4600);
nor U6994 (N_6994,N_3139,N_3125);
nand U6995 (N_6995,N_4543,N_4905);
nor U6996 (N_6996,N_2680,N_3340);
xor U6997 (N_6997,N_4418,N_4499);
and U6998 (N_6998,N_4691,N_3751);
xor U6999 (N_6999,N_3702,N_2826);
nor U7000 (N_7000,N_3349,N_3479);
xor U7001 (N_7001,N_4500,N_4178);
or U7002 (N_7002,N_2500,N_3011);
or U7003 (N_7003,N_4933,N_4169);
or U7004 (N_7004,N_4420,N_4147);
xor U7005 (N_7005,N_4925,N_3000);
xor U7006 (N_7006,N_3825,N_4681);
nor U7007 (N_7007,N_2641,N_4754);
or U7008 (N_7008,N_4290,N_4837);
nor U7009 (N_7009,N_3072,N_4355);
nor U7010 (N_7010,N_3071,N_4472);
xor U7011 (N_7011,N_4827,N_4157);
xnor U7012 (N_7012,N_3040,N_4313);
nor U7013 (N_7013,N_4003,N_3764);
nand U7014 (N_7014,N_3010,N_3146);
nor U7015 (N_7015,N_4255,N_3881);
nand U7016 (N_7016,N_4756,N_3641);
nor U7017 (N_7017,N_2822,N_2500);
xor U7018 (N_7018,N_4521,N_4223);
or U7019 (N_7019,N_3304,N_3068);
xor U7020 (N_7020,N_4512,N_3892);
and U7021 (N_7021,N_4734,N_3146);
or U7022 (N_7022,N_4385,N_2609);
nor U7023 (N_7023,N_3290,N_3547);
and U7024 (N_7024,N_4828,N_3798);
xor U7025 (N_7025,N_2951,N_4297);
nand U7026 (N_7026,N_2674,N_4131);
xnor U7027 (N_7027,N_4309,N_4648);
nor U7028 (N_7028,N_4395,N_3464);
nor U7029 (N_7029,N_4247,N_4925);
xor U7030 (N_7030,N_2809,N_4828);
and U7031 (N_7031,N_4934,N_3856);
or U7032 (N_7032,N_3065,N_3501);
or U7033 (N_7033,N_3419,N_3809);
nor U7034 (N_7034,N_4271,N_3580);
nor U7035 (N_7035,N_3294,N_4380);
and U7036 (N_7036,N_4914,N_4605);
and U7037 (N_7037,N_3219,N_4143);
xor U7038 (N_7038,N_4334,N_4962);
xor U7039 (N_7039,N_3841,N_3996);
or U7040 (N_7040,N_3228,N_4415);
nand U7041 (N_7041,N_4782,N_4802);
nor U7042 (N_7042,N_3739,N_3897);
nand U7043 (N_7043,N_3438,N_3613);
nor U7044 (N_7044,N_4214,N_4991);
or U7045 (N_7045,N_4901,N_2599);
nor U7046 (N_7046,N_3854,N_4499);
and U7047 (N_7047,N_3032,N_3625);
or U7048 (N_7048,N_3873,N_4927);
nand U7049 (N_7049,N_4946,N_4964);
nand U7050 (N_7050,N_2675,N_4539);
nor U7051 (N_7051,N_4161,N_3974);
xnor U7052 (N_7052,N_3980,N_3057);
and U7053 (N_7053,N_2670,N_2776);
and U7054 (N_7054,N_2565,N_3749);
xnor U7055 (N_7055,N_4809,N_2872);
nand U7056 (N_7056,N_3665,N_4959);
or U7057 (N_7057,N_3158,N_3299);
xor U7058 (N_7058,N_4303,N_3692);
and U7059 (N_7059,N_4244,N_3252);
nor U7060 (N_7060,N_4365,N_3850);
nand U7061 (N_7061,N_3434,N_3198);
nand U7062 (N_7062,N_4621,N_3501);
xnor U7063 (N_7063,N_3840,N_3240);
and U7064 (N_7064,N_2636,N_4508);
xor U7065 (N_7065,N_3557,N_2936);
xnor U7066 (N_7066,N_3759,N_3418);
xnor U7067 (N_7067,N_3140,N_4808);
nand U7068 (N_7068,N_3986,N_4147);
xor U7069 (N_7069,N_4323,N_4049);
nor U7070 (N_7070,N_4783,N_4792);
nor U7071 (N_7071,N_3571,N_3370);
or U7072 (N_7072,N_3367,N_3901);
nand U7073 (N_7073,N_3084,N_2775);
and U7074 (N_7074,N_4600,N_4200);
or U7075 (N_7075,N_4587,N_4999);
and U7076 (N_7076,N_4062,N_2652);
nor U7077 (N_7077,N_2553,N_4759);
and U7078 (N_7078,N_2795,N_3683);
or U7079 (N_7079,N_4957,N_4870);
xnor U7080 (N_7080,N_3970,N_4119);
and U7081 (N_7081,N_3956,N_4666);
or U7082 (N_7082,N_4364,N_4878);
nor U7083 (N_7083,N_2837,N_3848);
nand U7084 (N_7084,N_3865,N_3776);
or U7085 (N_7085,N_4251,N_2915);
and U7086 (N_7086,N_4111,N_4356);
xor U7087 (N_7087,N_4815,N_2986);
nand U7088 (N_7088,N_4378,N_3105);
xor U7089 (N_7089,N_3656,N_3371);
or U7090 (N_7090,N_3303,N_2524);
nand U7091 (N_7091,N_4853,N_4534);
nor U7092 (N_7092,N_4931,N_3285);
xor U7093 (N_7093,N_4789,N_2829);
and U7094 (N_7094,N_4125,N_2867);
nor U7095 (N_7095,N_3881,N_3099);
nand U7096 (N_7096,N_4124,N_2558);
nor U7097 (N_7097,N_4960,N_3053);
nand U7098 (N_7098,N_4110,N_3449);
nand U7099 (N_7099,N_2595,N_4965);
nand U7100 (N_7100,N_4093,N_2737);
nand U7101 (N_7101,N_3361,N_3436);
nor U7102 (N_7102,N_2737,N_4315);
or U7103 (N_7103,N_3824,N_4006);
or U7104 (N_7104,N_4027,N_3739);
nor U7105 (N_7105,N_3255,N_4432);
nand U7106 (N_7106,N_3388,N_4457);
and U7107 (N_7107,N_4453,N_3246);
nor U7108 (N_7108,N_4235,N_3370);
or U7109 (N_7109,N_4509,N_2849);
and U7110 (N_7110,N_2964,N_3236);
or U7111 (N_7111,N_3407,N_3421);
and U7112 (N_7112,N_4653,N_2885);
and U7113 (N_7113,N_4386,N_3400);
nand U7114 (N_7114,N_4672,N_3700);
and U7115 (N_7115,N_3654,N_2975);
and U7116 (N_7116,N_3435,N_4821);
or U7117 (N_7117,N_4960,N_4025);
nor U7118 (N_7118,N_3416,N_3594);
nand U7119 (N_7119,N_3175,N_3942);
nor U7120 (N_7120,N_3699,N_3386);
or U7121 (N_7121,N_2583,N_3788);
and U7122 (N_7122,N_4759,N_4289);
or U7123 (N_7123,N_4933,N_3725);
xnor U7124 (N_7124,N_3453,N_2569);
or U7125 (N_7125,N_3147,N_3621);
and U7126 (N_7126,N_3215,N_4718);
nor U7127 (N_7127,N_3238,N_4958);
xnor U7128 (N_7128,N_3632,N_4267);
nand U7129 (N_7129,N_2652,N_3229);
nand U7130 (N_7130,N_4722,N_3895);
nand U7131 (N_7131,N_3233,N_4607);
xnor U7132 (N_7132,N_3206,N_4062);
or U7133 (N_7133,N_4443,N_4498);
and U7134 (N_7134,N_3509,N_2580);
xnor U7135 (N_7135,N_4527,N_4093);
and U7136 (N_7136,N_3267,N_3728);
nor U7137 (N_7137,N_4352,N_3367);
nand U7138 (N_7138,N_3021,N_4633);
nor U7139 (N_7139,N_3199,N_4463);
or U7140 (N_7140,N_3559,N_3342);
xor U7141 (N_7141,N_3264,N_4281);
nor U7142 (N_7142,N_3500,N_4859);
xnor U7143 (N_7143,N_3678,N_2926);
or U7144 (N_7144,N_2932,N_2914);
nand U7145 (N_7145,N_2748,N_3163);
xnor U7146 (N_7146,N_2509,N_3135);
xor U7147 (N_7147,N_2793,N_4490);
xnor U7148 (N_7148,N_3914,N_3809);
xnor U7149 (N_7149,N_4432,N_3560);
nand U7150 (N_7150,N_4504,N_3038);
nor U7151 (N_7151,N_4965,N_4703);
nor U7152 (N_7152,N_3847,N_3238);
nand U7153 (N_7153,N_4385,N_2865);
nor U7154 (N_7154,N_3059,N_4099);
or U7155 (N_7155,N_4584,N_4816);
nand U7156 (N_7156,N_3641,N_2593);
or U7157 (N_7157,N_4914,N_2670);
nand U7158 (N_7158,N_4722,N_4486);
and U7159 (N_7159,N_4969,N_4047);
or U7160 (N_7160,N_3650,N_3114);
or U7161 (N_7161,N_3096,N_4918);
nand U7162 (N_7162,N_4650,N_3226);
xnor U7163 (N_7163,N_4640,N_2970);
nor U7164 (N_7164,N_4267,N_3014);
nand U7165 (N_7165,N_2889,N_4987);
or U7166 (N_7166,N_3997,N_4552);
xor U7167 (N_7167,N_3427,N_3594);
nor U7168 (N_7168,N_2585,N_3918);
xnor U7169 (N_7169,N_3528,N_3463);
or U7170 (N_7170,N_4515,N_3301);
xnor U7171 (N_7171,N_2914,N_2566);
nand U7172 (N_7172,N_2714,N_4989);
nand U7173 (N_7173,N_2570,N_4325);
or U7174 (N_7174,N_3172,N_4706);
and U7175 (N_7175,N_2923,N_3537);
nor U7176 (N_7176,N_4458,N_3059);
xor U7177 (N_7177,N_4872,N_4635);
xnor U7178 (N_7178,N_4087,N_2736);
or U7179 (N_7179,N_3500,N_4604);
and U7180 (N_7180,N_4141,N_3408);
and U7181 (N_7181,N_4757,N_3971);
nor U7182 (N_7182,N_4145,N_4542);
and U7183 (N_7183,N_4209,N_4258);
nand U7184 (N_7184,N_3388,N_2994);
nor U7185 (N_7185,N_3355,N_2989);
or U7186 (N_7186,N_4602,N_4405);
nor U7187 (N_7187,N_3613,N_4595);
xnor U7188 (N_7188,N_3308,N_4702);
and U7189 (N_7189,N_3146,N_4727);
nand U7190 (N_7190,N_4166,N_3224);
nand U7191 (N_7191,N_4408,N_2960);
xor U7192 (N_7192,N_4584,N_3021);
or U7193 (N_7193,N_2913,N_3221);
nand U7194 (N_7194,N_4136,N_4170);
xor U7195 (N_7195,N_3943,N_3201);
and U7196 (N_7196,N_3068,N_2580);
nand U7197 (N_7197,N_4763,N_3709);
and U7198 (N_7198,N_3624,N_3448);
xnor U7199 (N_7199,N_4810,N_4906);
nor U7200 (N_7200,N_3906,N_2977);
and U7201 (N_7201,N_4657,N_3032);
nand U7202 (N_7202,N_3146,N_3136);
and U7203 (N_7203,N_3210,N_4111);
nor U7204 (N_7204,N_4596,N_4983);
nor U7205 (N_7205,N_3529,N_2726);
or U7206 (N_7206,N_3538,N_2924);
nor U7207 (N_7207,N_3696,N_4118);
or U7208 (N_7208,N_3436,N_3883);
xor U7209 (N_7209,N_3386,N_3151);
xnor U7210 (N_7210,N_4369,N_4969);
and U7211 (N_7211,N_4493,N_4868);
xnor U7212 (N_7212,N_3408,N_3293);
xnor U7213 (N_7213,N_2758,N_2836);
nor U7214 (N_7214,N_4057,N_2759);
nor U7215 (N_7215,N_3080,N_4932);
nor U7216 (N_7216,N_3452,N_4989);
nor U7217 (N_7217,N_4280,N_2698);
and U7218 (N_7218,N_4720,N_3658);
nand U7219 (N_7219,N_4058,N_3395);
and U7220 (N_7220,N_3651,N_4552);
xnor U7221 (N_7221,N_3956,N_2638);
xnor U7222 (N_7222,N_3614,N_3453);
nor U7223 (N_7223,N_4889,N_3042);
nor U7224 (N_7224,N_3848,N_4379);
xor U7225 (N_7225,N_4229,N_2607);
or U7226 (N_7226,N_4639,N_4490);
nor U7227 (N_7227,N_4421,N_3924);
or U7228 (N_7228,N_4564,N_3542);
nor U7229 (N_7229,N_3354,N_2685);
or U7230 (N_7230,N_3334,N_4663);
nor U7231 (N_7231,N_3563,N_4293);
nor U7232 (N_7232,N_4019,N_4440);
nor U7233 (N_7233,N_4573,N_3066);
xnor U7234 (N_7234,N_4115,N_3690);
nor U7235 (N_7235,N_4356,N_4738);
or U7236 (N_7236,N_3357,N_3924);
or U7237 (N_7237,N_3090,N_3849);
or U7238 (N_7238,N_2964,N_4051);
and U7239 (N_7239,N_3398,N_2729);
and U7240 (N_7240,N_4627,N_3014);
nand U7241 (N_7241,N_4583,N_4014);
nor U7242 (N_7242,N_4857,N_3550);
xor U7243 (N_7243,N_3622,N_2608);
xor U7244 (N_7244,N_2771,N_4237);
nand U7245 (N_7245,N_3660,N_3501);
and U7246 (N_7246,N_3149,N_4840);
xnor U7247 (N_7247,N_4461,N_2935);
or U7248 (N_7248,N_4297,N_3609);
or U7249 (N_7249,N_3606,N_3029);
nor U7250 (N_7250,N_4356,N_2868);
or U7251 (N_7251,N_4994,N_4660);
or U7252 (N_7252,N_2854,N_3810);
or U7253 (N_7253,N_3998,N_4082);
and U7254 (N_7254,N_2904,N_2968);
or U7255 (N_7255,N_3963,N_4563);
or U7256 (N_7256,N_2622,N_3194);
and U7257 (N_7257,N_4378,N_3476);
and U7258 (N_7258,N_2986,N_2804);
nand U7259 (N_7259,N_4642,N_4177);
nor U7260 (N_7260,N_4547,N_4748);
or U7261 (N_7261,N_2575,N_4965);
nand U7262 (N_7262,N_3843,N_4893);
xnor U7263 (N_7263,N_4918,N_3664);
and U7264 (N_7264,N_2944,N_3834);
and U7265 (N_7265,N_4920,N_4119);
xnor U7266 (N_7266,N_2667,N_4263);
and U7267 (N_7267,N_3527,N_3894);
nand U7268 (N_7268,N_4209,N_2671);
or U7269 (N_7269,N_3119,N_2657);
and U7270 (N_7270,N_3200,N_3848);
nor U7271 (N_7271,N_3331,N_4686);
nand U7272 (N_7272,N_4183,N_3944);
nand U7273 (N_7273,N_3293,N_2529);
nor U7274 (N_7274,N_4874,N_3733);
xor U7275 (N_7275,N_3664,N_3298);
or U7276 (N_7276,N_2940,N_2669);
and U7277 (N_7277,N_3367,N_3403);
nand U7278 (N_7278,N_3876,N_3827);
or U7279 (N_7279,N_4523,N_3850);
xnor U7280 (N_7280,N_2896,N_2736);
xor U7281 (N_7281,N_4681,N_4933);
and U7282 (N_7282,N_4153,N_4117);
xor U7283 (N_7283,N_4911,N_3501);
nor U7284 (N_7284,N_3104,N_3931);
and U7285 (N_7285,N_3197,N_2860);
and U7286 (N_7286,N_4239,N_4715);
nand U7287 (N_7287,N_3698,N_3581);
and U7288 (N_7288,N_3111,N_4924);
or U7289 (N_7289,N_3567,N_2534);
xor U7290 (N_7290,N_3808,N_4967);
xor U7291 (N_7291,N_4555,N_2774);
nand U7292 (N_7292,N_2878,N_4589);
and U7293 (N_7293,N_4176,N_3364);
nand U7294 (N_7294,N_3012,N_3925);
or U7295 (N_7295,N_3714,N_2556);
and U7296 (N_7296,N_3707,N_3007);
nor U7297 (N_7297,N_3853,N_4074);
nand U7298 (N_7298,N_3266,N_3512);
xor U7299 (N_7299,N_4044,N_4710);
xor U7300 (N_7300,N_3109,N_4416);
or U7301 (N_7301,N_2599,N_3647);
and U7302 (N_7302,N_3177,N_3043);
xnor U7303 (N_7303,N_2914,N_4151);
nand U7304 (N_7304,N_3009,N_4767);
and U7305 (N_7305,N_2713,N_3280);
xnor U7306 (N_7306,N_2792,N_3835);
and U7307 (N_7307,N_4059,N_2880);
or U7308 (N_7308,N_3252,N_3242);
nor U7309 (N_7309,N_3598,N_4765);
and U7310 (N_7310,N_4502,N_3179);
nand U7311 (N_7311,N_4839,N_3236);
and U7312 (N_7312,N_3521,N_3057);
xor U7313 (N_7313,N_2954,N_4998);
nor U7314 (N_7314,N_3103,N_3765);
nand U7315 (N_7315,N_2981,N_2816);
and U7316 (N_7316,N_4728,N_4307);
and U7317 (N_7317,N_2860,N_3714);
or U7318 (N_7318,N_4371,N_4480);
or U7319 (N_7319,N_3463,N_2555);
nand U7320 (N_7320,N_3023,N_4216);
and U7321 (N_7321,N_3386,N_2750);
nand U7322 (N_7322,N_4705,N_3463);
and U7323 (N_7323,N_4587,N_2603);
nor U7324 (N_7324,N_2854,N_2874);
nand U7325 (N_7325,N_3423,N_4481);
xor U7326 (N_7326,N_4280,N_4639);
or U7327 (N_7327,N_4095,N_3861);
or U7328 (N_7328,N_2918,N_2848);
or U7329 (N_7329,N_2685,N_4284);
and U7330 (N_7330,N_2647,N_3904);
xor U7331 (N_7331,N_3955,N_4815);
nor U7332 (N_7332,N_3197,N_3168);
nor U7333 (N_7333,N_3219,N_3553);
or U7334 (N_7334,N_2681,N_3152);
xor U7335 (N_7335,N_3995,N_2986);
or U7336 (N_7336,N_3019,N_4576);
xor U7337 (N_7337,N_3141,N_4277);
nand U7338 (N_7338,N_2796,N_4559);
or U7339 (N_7339,N_4126,N_3339);
or U7340 (N_7340,N_4435,N_4081);
or U7341 (N_7341,N_3916,N_2928);
xor U7342 (N_7342,N_4182,N_3140);
nand U7343 (N_7343,N_3294,N_3564);
nor U7344 (N_7344,N_3788,N_2621);
xor U7345 (N_7345,N_2900,N_4589);
xor U7346 (N_7346,N_2962,N_4128);
or U7347 (N_7347,N_4929,N_4138);
nand U7348 (N_7348,N_3044,N_2835);
nand U7349 (N_7349,N_4062,N_2853);
nor U7350 (N_7350,N_3856,N_2837);
xnor U7351 (N_7351,N_4554,N_4403);
xnor U7352 (N_7352,N_4835,N_2969);
and U7353 (N_7353,N_4723,N_3547);
nand U7354 (N_7354,N_2703,N_4897);
nand U7355 (N_7355,N_2754,N_2710);
xor U7356 (N_7356,N_3515,N_3169);
xor U7357 (N_7357,N_3502,N_3855);
or U7358 (N_7358,N_3895,N_4192);
and U7359 (N_7359,N_4016,N_2639);
nor U7360 (N_7360,N_4222,N_4301);
nor U7361 (N_7361,N_4348,N_2640);
nor U7362 (N_7362,N_3852,N_4851);
and U7363 (N_7363,N_4690,N_4170);
nor U7364 (N_7364,N_3336,N_2554);
and U7365 (N_7365,N_4782,N_4715);
nor U7366 (N_7366,N_4512,N_4312);
nand U7367 (N_7367,N_4225,N_3918);
nor U7368 (N_7368,N_3879,N_2529);
or U7369 (N_7369,N_2786,N_3109);
nand U7370 (N_7370,N_3657,N_2589);
or U7371 (N_7371,N_4515,N_3359);
nor U7372 (N_7372,N_3420,N_3215);
nor U7373 (N_7373,N_3912,N_3204);
nor U7374 (N_7374,N_4859,N_3260);
nor U7375 (N_7375,N_4002,N_3049);
or U7376 (N_7376,N_4844,N_4150);
nand U7377 (N_7377,N_2850,N_3925);
nand U7378 (N_7378,N_3286,N_2856);
or U7379 (N_7379,N_4867,N_3752);
xor U7380 (N_7380,N_3423,N_4304);
nand U7381 (N_7381,N_4933,N_2955);
nor U7382 (N_7382,N_3388,N_4841);
nor U7383 (N_7383,N_4790,N_3466);
nand U7384 (N_7384,N_3583,N_3138);
nor U7385 (N_7385,N_2553,N_4402);
and U7386 (N_7386,N_3779,N_3347);
xnor U7387 (N_7387,N_4122,N_4169);
xor U7388 (N_7388,N_4121,N_2736);
nand U7389 (N_7389,N_4183,N_3501);
nor U7390 (N_7390,N_4438,N_2742);
nand U7391 (N_7391,N_2893,N_3700);
and U7392 (N_7392,N_4458,N_2798);
and U7393 (N_7393,N_3269,N_2703);
xnor U7394 (N_7394,N_3265,N_4780);
and U7395 (N_7395,N_3913,N_4846);
and U7396 (N_7396,N_4176,N_2880);
xor U7397 (N_7397,N_4421,N_3083);
xor U7398 (N_7398,N_3277,N_2903);
nor U7399 (N_7399,N_2922,N_4586);
or U7400 (N_7400,N_4373,N_4437);
and U7401 (N_7401,N_4312,N_3195);
and U7402 (N_7402,N_3573,N_4625);
nor U7403 (N_7403,N_3376,N_2671);
nor U7404 (N_7404,N_4696,N_4494);
or U7405 (N_7405,N_3999,N_4601);
nor U7406 (N_7406,N_4305,N_4740);
or U7407 (N_7407,N_3079,N_4380);
nor U7408 (N_7408,N_3535,N_3407);
or U7409 (N_7409,N_3819,N_3933);
nor U7410 (N_7410,N_3436,N_4506);
and U7411 (N_7411,N_4898,N_3193);
nor U7412 (N_7412,N_4555,N_4608);
xor U7413 (N_7413,N_4538,N_4332);
nor U7414 (N_7414,N_4571,N_4811);
and U7415 (N_7415,N_3135,N_3917);
nor U7416 (N_7416,N_3468,N_3151);
nand U7417 (N_7417,N_3211,N_3543);
nand U7418 (N_7418,N_2844,N_4293);
or U7419 (N_7419,N_3289,N_4174);
and U7420 (N_7420,N_3942,N_3730);
and U7421 (N_7421,N_4803,N_4341);
nor U7422 (N_7422,N_2909,N_4016);
nand U7423 (N_7423,N_4621,N_4244);
nand U7424 (N_7424,N_4012,N_4191);
xnor U7425 (N_7425,N_3856,N_2561);
and U7426 (N_7426,N_3197,N_4594);
xnor U7427 (N_7427,N_4522,N_4875);
or U7428 (N_7428,N_3155,N_4863);
nor U7429 (N_7429,N_4647,N_3015);
and U7430 (N_7430,N_4355,N_4025);
or U7431 (N_7431,N_4418,N_4425);
and U7432 (N_7432,N_3270,N_2829);
and U7433 (N_7433,N_4762,N_4301);
xor U7434 (N_7434,N_3306,N_4173);
nor U7435 (N_7435,N_2954,N_3053);
or U7436 (N_7436,N_3137,N_2850);
xnor U7437 (N_7437,N_4142,N_3381);
nor U7438 (N_7438,N_4152,N_4657);
nor U7439 (N_7439,N_2612,N_4488);
or U7440 (N_7440,N_2906,N_3412);
and U7441 (N_7441,N_4544,N_3447);
nand U7442 (N_7442,N_2605,N_3611);
and U7443 (N_7443,N_4961,N_4685);
xor U7444 (N_7444,N_2898,N_4636);
nor U7445 (N_7445,N_4653,N_3494);
and U7446 (N_7446,N_4346,N_4136);
nand U7447 (N_7447,N_3511,N_4078);
or U7448 (N_7448,N_4175,N_4400);
xnor U7449 (N_7449,N_2818,N_4174);
nor U7450 (N_7450,N_4048,N_4844);
or U7451 (N_7451,N_2983,N_2680);
or U7452 (N_7452,N_4903,N_4570);
nand U7453 (N_7453,N_3585,N_2661);
or U7454 (N_7454,N_4417,N_3181);
or U7455 (N_7455,N_4897,N_3099);
nand U7456 (N_7456,N_4795,N_2749);
or U7457 (N_7457,N_4477,N_4556);
or U7458 (N_7458,N_3141,N_3922);
xor U7459 (N_7459,N_3046,N_4811);
or U7460 (N_7460,N_4370,N_3484);
or U7461 (N_7461,N_4520,N_2604);
and U7462 (N_7462,N_3193,N_3629);
and U7463 (N_7463,N_3100,N_4139);
xor U7464 (N_7464,N_2735,N_4648);
nor U7465 (N_7465,N_3024,N_4335);
nand U7466 (N_7466,N_4005,N_3454);
nor U7467 (N_7467,N_4940,N_4173);
xnor U7468 (N_7468,N_4880,N_3922);
nor U7469 (N_7469,N_4074,N_4313);
xnor U7470 (N_7470,N_4460,N_3431);
or U7471 (N_7471,N_4244,N_4535);
xor U7472 (N_7472,N_3125,N_4679);
nand U7473 (N_7473,N_3804,N_2995);
and U7474 (N_7474,N_3695,N_4157);
xnor U7475 (N_7475,N_3716,N_3524);
and U7476 (N_7476,N_2969,N_4781);
nand U7477 (N_7477,N_3461,N_3544);
nand U7478 (N_7478,N_4539,N_3875);
xnor U7479 (N_7479,N_4772,N_4090);
xor U7480 (N_7480,N_3746,N_4655);
nor U7481 (N_7481,N_3409,N_2840);
or U7482 (N_7482,N_3169,N_4358);
and U7483 (N_7483,N_3484,N_2615);
and U7484 (N_7484,N_4841,N_3526);
xnor U7485 (N_7485,N_4431,N_3917);
nand U7486 (N_7486,N_4264,N_2575);
or U7487 (N_7487,N_2518,N_3990);
xnor U7488 (N_7488,N_4996,N_2640);
or U7489 (N_7489,N_3313,N_4764);
nor U7490 (N_7490,N_4486,N_2505);
or U7491 (N_7491,N_2676,N_4493);
xnor U7492 (N_7492,N_4705,N_3676);
nor U7493 (N_7493,N_4674,N_4448);
and U7494 (N_7494,N_2974,N_3736);
nor U7495 (N_7495,N_3291,N_3932);
nand U7496 (N_7496,N_3520,N_3694);
and U7497 (N_7497,N_4970,N_2981);
xnor U7498 (N_7498,N_3808,N_3813);
nand U7499 (N_7499,N_4253,N_3492);
and U7500 (N_7500,N_5908,N_6748);
or U7501 (N_7501,N_7199,N_6092);
nand U7502 (N_7502,N_6007,N_6674);
and U7503 (N_7503,N_5442,N_5099);
xor U7504 (N_7504,N_5862,N_6433);
nor U7505 (N_7505,N_5218,N_6199);
nor U7506 (N_7506,N_6905,N_7310);
or U7507 (N_7507,N_5669,N_5162);
nor U7508 (N_7508,N_5065,N_5976);
or U7509 (N_7509,N_5420,N_7362);
xor U7510 (N_7510,N_6628,N_6936);
or U7511 (N_7511,N_6062,N_6590);
xor U7512 (N_7512,N_7309,N_6190);
or U7513 (N_7513,N_6696,N_6086);
xor U7514 (N_7514,N_6323,N_6453);
or U7515 (N_7515,N_5175,N_5901);
nand U7516 (N_7516,N_6601,N_7358);
xor U7517 (N_7517,N_5907,N_5252);
and U7518 (N_7518,N_7042,N_5878);
or U7519 (N_7519,N_5048,N_6795);
nor U7520 (N_7520,N_6621,N_7256);
nor U7521 (N_7521,N_5847,N_5251);
and U7522 (N_7522,N_5438,N_7235);
nor U7523 (N_7523,N_6799,N_5685);
and U7524 (N_7524,N_6931,N_5414);
nand U7525 (N_7525,N_6700,N_6355);
and U7526 (N_7526,N_6247,N_6720);
nor U7527 (N_7527,N_6450,N_5645);
or U7528 (N_7528,N_7018,N_6763);
and U7529 (N_7529,N_5947,N_5702);
nor U7530 (N_7530,N_6192,N_6363);
or U7531 (N_7531,N_5422,N_6903);
or U7532 (N_7532,N_6438,N_7385);
nand U7533 (N_7533,N_5443,N_6978);
nand U7534 (N_7534,N_6717,N_5143);
nand U7535 (N_7535,N_6786,N_6727);
nand U7536 (N_7536,N_5830,N_6980);
and U7537 (N_7537,N_5350,N_5011);
or U7538 (N_7538,N_6530,N_6558);
or U7539 (N_7539,N_5558,N_7110);
nand U7540 (N_7540,N_6859,N_6298);
xnor U7541 (N_7541,N_5581,N_7477);
or U7542 (N_7542,N_5625,N_5803);
or U7543 (N_7543,N_6507,N_6402);
nand U7544 (N_7544,N_6326,N_6569);
nor U7545 (N_7545,N_7194,N_5063);
nor U7546 (N_7546,N_6752,N_7205);
xnor U7547 (N_7547,N_7340,N_6833);
nor U7548 (N_7548,N_5681,N_6739);
and U7549 (N_7549,N_5486,N_6877);
or U7550 (N_7550,N_6102,N_7287);
or U7551 (N_7551,N_6059,N_7471);
and U7552 (N_7552,N_6879,N_5144);
or U7553 (N_7553,N_6504,N_7293);
nand U7554 (N_7554,N_6571,N_7258);
and U7555 (N_7555,N_6112,N_6626);
xor U7556 (N_7556,N_7103,N_6774);
nand U7557 (N_7557,N_5870,N_7388);
nand U7558 (N_7558,N_7043,N_6406);
or U7559 (N_7559,N_6452,N_5651);
nand U7560 (N_7560,N_6224,N_5551);
nor U7561 (N_7561,N_5899,N_6339);
nor U7562 (N_7562,N_5305,N_6275);
or U7563 (N_7563,N_5409,N_5723);
xor U7564 (N_7564,N_6580,N_6635);
nor U7565 (N_7565,N_5891,N_5731);
or U7566 (N_7566,N_5391,N_6297);
xnor U7567 (N_7567,N_7026,N_5761);
and U7568 (N_7568,N_5642,N_5213);
and U7569 (N_7569,N_5936,N_6058);
and U7570 (N_7570,N_6501,N_5410);
and U7571 (N_7571,N_6460,N_6971);
xnor U7572 (N_7572,N_5676,N_6565);
xnor U7573 (N_7573,N_5521,N_7137);
nand U7574 (N_7574,N_5666,N_5147);
or U7575 (N_7575,N_5224,N_5017);
xor U7576 (N_7576,N_5186,N_6087);
or U7577 (N_7577,N_5079,N_7443);
nor U7578 (N_7578,N_6898,N_7476);
and U7579 (N_7579,N_5054,N_6074);
xnor U7580 (N_7580,N_6459,N_5771);
nand U7581 (N_7581,N_5270,N_6437);
or U7582 (N_7582,N_7459,N_5788);
nor U7583 (N_7583,N_7207,N_5254);
or U7584 (N_7584,N_5539,N_6187);
nand U7585 (N_7585,N_7263,N_7010);
xor U7586 (N_7586,N_5248,N_5961);
or U7587 (N_7587,N_5717,N_7058);
and U7588 (N_7588,N_5366,N_5025);
or U7589 (N_7589,N_5868,N_6928);
or U7590 (N_7590,N_6364,N_6334);
or U7591 (N_7591,N_6630,N_5603);
and U7592 (N_7592,N_5670,N_5720);
xor U7593 (N_7593,N_7143,N_6746);
xor U7594 (N_7594,N_6867,N_6647);
nand U7595 (N_7595,N_7463,N_5596);
nand U7596 (N_7596,N_5841,N_5534);
xor U7597 (N_7597,N_6979,N_6408);
nand U7598 (N_7598,N_7253,N_7360);
and U7599 (N_7599,N_6473,N_5902);
or U7600 (N_7600,N_5972,N_6890);
nand U7601 (N_7601,N_6889,N_5996);
or U7602 (N_7602,N_6117,N_6732);
nand U7603 (N_7603,N_7370,N_5335);
or U7604 (N_7604,N_5879,N_5544);
nor U7605 (N_7605,N_7461,N_6616);
xnor U7606 (N_7606,N_6693,N_6308);
nor U7607 (N_7607,N_5797,N_6857);
nand U7608 (N_7608,N_5986,N_6232);
and U7609 (N_7609,N_6900,N_6722);
nor U7610 (N_7610,N_6332,N_5705);
or U7611 (N_7611,N_5455,N_5880);
or U7612 (N_7612,N_6950,N_6745);
or U7613 (N_7613,N_5524,N_5106);
nor U7614 (N_7614,N_6728,N_6330);
nor U7615 (N_7615,N_5641,N_6123);
nor U7616 (N_7616,N_6065,N_6870);
nand U7617 (N_7617,N_6049,N_5363);
and U7618 (N_7618,N_5062,N_7341);
nor U7619 (N_7619,N_6083,N_6424);
nor U7620 (N_7620,N_5174,N_6855);
or U7621 (N_7621,N_7254,N_5703);
xnor U7622 (N_7622,N_7333,N_5662);
or U7623 (N_7623,N_5495,N_5450);
and U7624 (N_7624,N_7474,N_6362);
and U7625 (N_7625,N_6317,N_5574);
or U7626 (N_7626,N_6506,N_5719);
and U7627 (N_7627,N_6482,N_5914);
nand U7628 (N_7628,N_5272,N_6038);
xnor U7629 (N_7629,N_6425,N_7037);
or U7630 (N_7630,N_7180,N_6243);
nand U7631 (N_7631,N_7086,N_6932);
xnor U7632 (N_7632,N_6798,N_6961);
nor U7633 (N_7633,N_6707,N_5142);
xnor U7634 (N_7634,N_5597,N_5009);
xor U7635 (N_7635,N_6860,N_6228);
nor U7636 (N_7636,N_5289,N_6288);
nor U7637 (N_7637,N_5056,N_6962);
nand U7638 (N_7638,N_6073,N_5741);
nor U7639 (N_7639,N_5206,N_5917);
and U7640 (N_7640,N_5141,N_7068);
or U7641 (N_7641,N_6815,N_5814);
and U7642 (N_7642,N_5547,N_5449);
xor U7643 (N_7643,N_6060,N_6706);
nand U7644 (N_7644,N_6909,N_7150);
and U7645 (N_7645,N_6515,N_6529);
nand U7646 (N_7646,N_5707,N_5822);
nand U7647 (N_7647,N_6120,N_5842);
and U7648 (N_7648,N_6607,N_6213);
and U7649 (N_7649,N_5619,N_5858);
or U7650 (N_7650,N_5714,N_5145);
or U7651 (N_7651,N_6524,N_6201);
nor U7652 (N_7652,N_7378,N_7190);
xor U7653 (N_7653,N_6742,N_5713);
and U7654 (N_7654,N_5831,N_5284);
nor U7655 (N_7655,N_5857,N_6015);
and U7656 (N_7656,N_5237,N_5390);
and U7657 (N_7657,N_6109,N_6066);
and U7658 (N_7658,N_6446,N_6785);
xor U7659 (N_7659,N_5983,N_6651);
nand U7660 (N_7660,N_5088,N_5828);
xnor U7661 (N_7661,N_7383,N_5211);
or U7662 (N_7662,N_5989,N_6119);
or U7663 (N_7663,N_5392,N_5834);
nand U7664 (N_7664,N_7130,N_6027);
nand U7665 (N_7665,N_6531,N_5968);
nand U7666 (N_7666,N_5884,N_5140);
nand U7667 (N_7667,N_7300,N_6411);
xnor U7668 (N_7668,N_6555,N_6078);
or U7669 (N_7669,N_6612,N_6067);
or U7670 (N_7670,N_5281,N_6891);
or U7671 (N_7671,N_6988,N_7078);
nand U7672 (N_7672,N_6142,N_6668);
nand U7673 (N_7673,N_7319,N_6287);
and U7674 (N_7674,N_6395,N_6248);
nor U7675 (N_7675,N_6577,N_7415);
and U7676 (N_7676,N_5733,N_5630);
nand U7677 (N_7677,N_5308,N_6002);
or U7678 (N_7678,N_5837,N_5718);
nor U7679 (N_7679,N_6274,N_5529);
and U7680 (N_7680,N_7246,N_7083);
nand U7681 (N_7681,N_6465,N_6495);
xor U7682 (N_7682,N_5214,N_6904);
or U7683 (N_7683,N_5624,N_6672);
and U7684 (N_7684,N_7040,N_5698);
nand U7685 (N_7685,N_6510,N_7065);
nand U7686 (N_7686,N_7070,N_6851);
or U7687 (N_7687,N_6829,N_6773);
or U7688 (N_7688,N_6464,N_5192);
xor U7689 (N_7689,N_5941,N_6794);
nand U7690 (N_7690,N_6563,N_7213);
nand U7691 (N_7691,N_6939,N_6412);
xnor U7692 (N_7692,N_6675,N_6549);
and U7693 (N_7693,N_5098,N_5607);
or U7694 (N_7694,N_5960,N_6309);
nor U7695 (N_7695,N_5052,N_6350);
or U7696 (N_7696,N_5935,N_6695);
xnor U7697 (N_7697,N_6296,N_6995);
xnor U7698 (N_7698,N_6152,N_7116);
xnor U7699 (N_7699,N_7326,N_6692);
nor U7700 (N_7700,N_6862,N_5474);
xnor U7701 (N_7701,N_5523,N_7311);
and U7702 (N_7702,N_5944,N_5688);
nand U7703 (N_7703,N_7303,N_7033);
and U7704 (N_7704,N_5038,N_6155);
nand U7705 (N_7705,N_6907,N_6172);
nand U7706 (N_7706,N_6743,N_5673);
xnor U7707 (N_7707,N_6861,N_7422);
nor U7708 (N_7708,N_6500,N_6440);
xor U7709 (N_7709,N_7075,N_6705);
nand U7710 (N_7710,N_6113,N_6699);
nor U7711 (N_7711,N_7000,N_5776);
nand U7712 (N_7712,N_5752,N_6656);
and U7713 (N_7713,N_5490,N_5484);
nand U7714 (N_7714,N_6384,N_7283);
nor U7715 (N_7715,N_6535,N_6345);
nand U7716 (N_7716,N_5362,N_7494);
or U7717 (N_7717,N_6589,N_7134);
xor U7718 (N_7718,N_5924,N_5854);
and U7719 (N_7719,N_6873,N_5105);
nand U7720 (N_7720,N_6373,N_6250);
and U7721 (N_7721,N_7330,N_6998);
xor U7722 (N_7722,N_6044,N_5006);
or U7723 (N_7723,N_5792,N_5058);
or U7724 (N_7724,N_6088,N_7483);
xnor U7725 (N_7725,N_7406,N_5877);
nor U7726 (N_7726,N_5791,N_7302);
and U7727 (N_7727,N_5087,N_7423);
xor U7728 (N_7728,N_5093,N_6263);
or U7729 (N_7729,N_5037,N_6755);
xnor U7730 (N_7730,N_5253,N_5709);
nor U7731 (N_7731,N_5588,N_6477);
nand U7732 (N_7732,N_5617,N_6340);
and U7733 (N_7733,N_5153,N_7465);
nand U7734 (N_7734,N_5601,N_6753);
xnor U7735 (N_7735,N_6645,N_6806);
nand U7736 (N_7736,N_6356,N_5781);
or U7737 (N_7737,N_5602,N_6603);
nand U7738 (N_7738,N_6377,N_5311);
or U7739 (N_7739,N_5202,N_7499);
or U7740 (N_7740,N_5234,N_5347);
xor U7741 (N_7741,N_6709,N_6761);
or U7742 (N_7742,N_7480,N_5198);
or U7743 (N_7743,N_5659,N_5282);
nor U7744 (N_7744,N_7136,N_6121);
or U7745 (N_7745,N_6631,N_6085);
nor U7746 (N_7746,N_5897,N_5262);
xor U7747 (N_7747,N_6012,N_7401);
and U7748 (N_7748,N_6959,N_6032);
and U7749 (N_7749,N_7280,N_7184);
nor U7750 (N_7750,N_6104,N_5783);
nand U7751 (N_7751,N_5326,N_5321);
nand U7752 (N_7752,N_6294,N_5775);
and U7753 (N_7753,N_5667,N_6467);
and U7754 (N_7754,N_6511,N_7023);
xnor U7755 (N_7755,N_5405,N_7251);
and U7756 (N_7756,N_6319,N_5616);
xnor U7757 (N_7757,N_6726,N_6649);
and U7758 (N_7758,N_7455,N_7453);
nor U7759 (N_7759,N_6416,N_6574);
or U7760 (N_7760,N_6608,N_6866);
and U7761 (N_7761,N_5955,N_6286);
xnor U7762 (N_7762,N_7234,N_5869);
nor U7763 (N_7763,N_5779,N_5991);
or U7764 (N_7764,N_7097,N_6548);
nand U7765 (N_7765,N_5090,N_5905);
and U7766 (N_7766,N_6846,N_5297);
nand U7767 (N_7767,N_5351,N_6354);
nor U7768 (N_7768,N_5375,N_6167);
nand U7769 (N_7769,N_7284,N_7131);
xnor U7770 (N_7770,N_5389,N_6272);
xnor U7771 (N_7771,N_6533,N_5816);
and U7772 (N_7772,N_7346,N_6754);
or U7773 (N_7773,N_6780,N_7305);
and U7774 (N_7774,N_7266,N_5122);
nor U7775 (N_7775,N_6600,N_6069);
and U7776 (N_7776,N_7357,N_5100);
or U7777 (N_7777,N_5456,N_5463);
nand U7778 (N_7778,N_5760,N_6783);
nor U7779 (N_7779,N_6756,N_5344);
xor U7780 (N_7780,N_7336,N_6893);
xor U7781 (N_7781,N_7030,N_5593);
or U7782 (N_7782,N_6037,N_6215);
xor U7783 (N_7783,N_5313,N_6987);
xnor U7784 (N_7784,N_6981,N_7306);
xnor U7785 (N_7785,N_5137,N_5113);
and U7786 (N_7786,N_7090,N_6994);
or U7787 (N_7787,N_6999,N_5554);
and U7788 (N_7788,N_6912,N_5888);
or U7789 (N_7789,N_5235,N_7087);
xnor U7790 (N_7790,N_6305,N_7249);
or U7791 (N_7791,N_6071,N_5999);
xor U7792 (N_7792,N_6797,N_6982);
or U7793 (N_7793,N_5967,N_5277);
and U7794 (N_7794,N_5700,N_6264);
and U7795 (N_7795,N_5077,N_6702);
nand U7796 (N_7796,N_6441,N_5686);
and U7797 (N_7797,N_6772,N_6749);
nor U7798 (N_7798,N_6986,N_7329);
and U7799 (N_7799,N_5710,N_6919);
xnor U7800 (N_7800,N_6771,N_5876);
nor U7801 (N_7801,N_5892,N_6249);
nor U7802 (N_7802,N_5171,N_5610);
nand U7803 (N_7803,N_6644,N_7486);
and U7804 (N_7804,N_7104,N_7387);
nor U7805 (N_7805,N_7301,N_5419);
or U7806 (N_7806,N_5992,N_7117);
nand U7807 (N_7807,N_7394,N_6239);
and U7808 (N_7808,N_5061,N_5606);
nand U7809 (N_7809,N_6947,N_7482);
nand U7810 (N_7810,N_5833,N_6646);
or U7811 (N_7811,N_6141,N_5158);
xnor U7812 (N_7812,N_5342,N_6874);
and U7813 (N_7813,N_7107,N_6256);
and U7814 (N_7814,N_7105,N_6137);
nand U7815 (N_7815,N_6942,N_7392);
nor U7816 (N_7816,N_6267,N_7487);
nor U7817 (N_7817,N_5071,N_5930);
nor U7818 (N_7818,N_6016,N_7007);
nor U7819 (N_7819,N_7160,N_5346);
and U7820 (N_7820,N_7414,N_6856);
nor U7821 (N_7821,N_6337,N_5356);
nand U7822 (N_7822,N_6127,N_6481);
xnor U7823 (N_7823,N_5107,N_6953);
xor U7824 (N_7824,N_6985,N_6399);
nand U7825 (N_7825,N_6366,N_5818);
and U7826 (N_7826,N_6144,N_5029);
xor U7827 (N_7827,N_7331,N_5369);
xor U7828 (N_7828,N_5839,N_6901);
nand U7829 (N_7829,N_7462,N_6368);
and U7830 (N_7830,N_5314,N_7203);
xnor U7831 (N_7831,N_5469,N_6906);
xnor U7832 (N_7832,N_5291,N_5926);
and U7833 (N_7833,N_5033,N_5993);
xnor U7834 (N_7834,N_6487,N_5806);
xnor U7835 (N_7835,N_5287,N_6642);
xor U7836 (N_7836,N_6552,N_7032);
nor U7837 (N_7837,N_5959,N_6423);
nor U7838 (N_7838,N_5382,N_6610);
nand U7839 (N_7839,N_7091,N_6878);
xnor U7840 (N_7840,N_6760,N_7402);
nand U7841 (N_7841,N_6976,N_6301);
or U7842 (N_7842,N_5373,N_7475);
xor U7843 (N_7843,N_5019,N_7397);
nand U7844 (N_7844,N_7100,N_5078);
nor U7845 (N_7845,N_7322,N_5358);
nand U7846 (N_7846,N_5750,N_5937);
or U7847 (N_7847,N_5751,N_6945);
xor U7848 (N_7848,N_7257,N_7400);
and U7849 (N_7849,N_5125,N_7288);
and U7850 (N_7850,N_6544,N_7156);
nand U7851 (N_7851,N_6394,N_6389);
and U7852 (N_7852,N_5525,N_6385);
and U7853 (N_7853,N_5827,N_5678);
or U7854 (N_7854,N_6843,N_7048);
and U7855 (N_7855,N_7237,N_5694);
nor U7856 (N_7856,N_5478,N_5181);
nor U7857 (N_7857,N_6129,N_6240);
nand U7858 (N_7858,N_6028,N_7489);
or U7859 (N_7859,N_7404,N_5051);
nand U7860 (N_7860,N_6850,N_6973);
nor U7861 (N_7861,N_5004,N_6039);
xor U7862 (N_7862,N_5221,N_5126);
and U7863 (N_7863,N_5467,N_5608);
or U7864 (N_7864,N_5501,N_6790);
xor U7865 (N_7865,N_5454,N_5911);
nand U7866 (N_7866,N_6946,N_6639);
and U7867 (N_7867,N_5819,N_6949);
xor U7868 (N_7868,N_5365,N_5368);
or U7869 (N_7869,N_6824,N_6072);
xor U7870 (N_7870,N_6220,N_6318);
and U7871 (N_7871,N_7095,N_6892);
or U7872 (N_7872,N_5757,N_7147);
or U7873 (N_7873,N_6367,N_6966);
xnor U7874 (N_7874,N_6740,N_6871);
or U7875 (N_7875,N_5782,N_6951);
xnor U7876 (N_7876,N_6253,N_5337);
nand U7877 (N_7877,N_5777,N_7270);
or U7878 (N_7878,N_6744,N_5549);
nor U7879 (N_7879,N_6210,N_6415);
nand U7880 (N_7880,N_5426,N_5430);
nand U7881 (N_7881,N_7098,N_6703);
nor U7882 (N_7882,N_7313,N_5998);
nand U7883 (N_7883,N_6004,N_6047);
nand U7884 (N_7884,N_6403,N_5039);
nand U7885 (N_7885,N_7102,N_6943);
nor U7886 (N_7886,N_6324,N_5505);
xor U7887 (N_7887,N_5894,N_5226);
and U7888 (N_7888,N_5191,N_6204);
or U7889 (N_7889,N_5860,N_5049);
and U7890 (N_7890,N_7279,N_5560);
or U7891 (N_7891,N_5200,N_5903);
and U7892 (N_7892,N_6392,N_6054);
nand U7893 (N_7893,N_5498,N_6081);
or U7894 (N_7894,N_6184,N_6025);
nor U7895 (N_7895,N_5349,N_5159);
or U7896 (N_7896,N_5031,N_7248);
or U7897 (N_7897,N_6788,N_6005);
nand U7898 (N_7898,N_6875,N_5249);
xnor U7899 (N_7899,N_7044,N_7114);
nor U7900 (N_7900,N_5292,N_6684);
nand U7901 (N_7901,N_5925,N_5487);
nor U7902 (N_7902,N_7332,N_5725);
or U7903 (N_7903,N_6321,N_5339);
and U7904 (N_7904,N_5728,N_5084);
and U7905 (N_7905,N_6920,N_5399);
nand U7906 (N_7906,N_5408,N_5121);
xor U7907 (N_7907,N_6822,N_5429);
nor U7908 (N_7908,N_6338,N_6478);
or U7909 (N_7909,N_7294,N_6536);
xor U7910 (N_7910,N_6082,N_6447);
and U7911 (N_7911,N_6398,N_7316);
or U7912 (N_7912,N_6808,N_7082);
nand U7913 (N_7913,N_5310,N_6602);
or U7914 (N_7914,N_7013,N_5473);
or U7915 (N_7915,N_6553,N_5280);
nor U7916 (N_7916,N_6230,N_5010);
or U7917 (N_7917,N_7093,N_6923);
and U7918 (N_7918,N_5974,N_5599);
nand U7919 (N_7919,N_6386,N_6370);
xor U7920 (N_7920,N_6114,N_6801);
nor U7921 (N_7921,N_5739,N_6200);
nand U7922 (N_7922,N_6781,N_5178);
nand U7923 (N_7923,N_6479,N_6770);
or U7924 (N_7924,N_7276,N_5464);
or U7925 (N_7925,N_6681,N_7118);
nand U7926 (N_7926,N_6992,N_5811);
or U7927 (N_7927,N_6925,N_5510);
xnor U7928 (N_7928,N_5848,N_7315);
and U7929 (N_7929,N_6758,N_6993);
nor U7930 (N_7930,N_6352,N_6880);
xor U7931 (N_7931,N_7009,N_5359);
or U7932 (N_7932,N_6970,N_5805);
and U7933 (N_7933,N_5433,N_5264);
or U7934 (N_7934,N_6276,N_6365);
and U7935 (N_7935,N_5747,N_5795);
and U7936 (N_7936,N_6048,N_6838);
and U7937 (N_7937,N_5067,N_5222);
xnor U7938 (N_7938,N_5655,N_7012);
nor U7939 (N_7939,N_5290,N_6343);
or U7940 (N_7940,N_7430,N_6108);
nand U7941 (N_7941,N_7014,N_6849);
xnor U7942 (N_7942,N_6390,N_5118);
xor U7943 (N_7943,N_7011,N_7324);
nand U7944 (N_7944,N_6793,N_5954);
xor U7945 (N_7945,N_5123,N_6528);
nor U7946 (N_7946,N_7005,N_5453);
and U7947 (N_7947,N_5384,N_5555);
nor U7948 (N_7948,N_5568,N_7435);
nand U7949 (N_7949,N_6842,N_5030);
nand U7950 (N_7950,N_7432,N_6492);
nand U7951 (N_7951,N_5519,N_5613);
nand U7952 (N_7952,N_6115,N_5522);
and U7953 (N_7953,N_6217,N_7488);
and U7954 (N_7954,N_5851,N_5329);
and U7955 (N_7955,N_6181,N_6764);
nand U7956 (N_7956,N_5266,N_6568);
and U7957 (N_7957,N_5016,N_5117);
nand U7958 (N_7958,N_7186,N_5537);
and U7959 (N_7959,N_6844,N_6462);
nand U7960 (N_7960,N_6671,N_5288);
xor U7961 (N_7961,N_6295,N_5950);
xnor U7962 (N_7962,N_5278,N_7212);
and U7963 (N_7963,N_6592,N_7157);
or U7964 (N_7964,N_5507,N_5397);
nor U7965 (N_7965,N_5825,N_7445);
xnor U7966 (N_7966,N_6111,N_7250);
nand U7967 (N_7967,N_7245,N_5503);
nand U7968 (N_7968,N_5623,N_5789);
xnor U7969 (N_7969,N_5977,N_6451);
nor U7970 (N_7970,N_5912,N_7493);
and U7971 (N_7971,N_7144,N_5546);
and U7972 (N_7972,N_5824,N_5132);
xor U7973 (N_7973,N_6599,N_5843);
or U7974 (N_7974,N_5708,N_6261);
and U7975 (N_7975,N_7289,N_7099);
xor U7976 (N_7976,N_5661,N_5732);
xnor U7977 (N_7977,N_6101,N_6730);
or U7978 (N_7978,N_6554,N_6227);
nand U7979 (N_7979,N_5590,N_5157);
or U7980 (N_7980,N_7365,N_5518);
and U7981 (N_7981,N_5784,N_6211);
or U7982 (N_7982,N_5866,N_6526);
or U7983 (N_7983,N_5459,N_5418);
or U7984 (N_7984,N_5324,N_7449);
or U7985 (N_7985,N_5561,N_6502);
nor U7986 (N_7986,N_6997,N_6143);
and U7987 (N_7987,N_6733,N_5167);
and U7988 (N_7988,N_6245,N_6461);
nand U7989 (N_7989,N_5953,N_6140);
nor U7990 (N_7990,N_5730,N_5479);
and U7991 (N_7991,N_6654,N_7307);
or U7992 (N_7992,N_7101,N_7175);
nor U7993 (N_7993,N_5753,N_7063);
nor U7994 (N_7994,N_7154,N_6594);
nand U7995 (N_7995,N_6050,N_6591);
and U7996 (N_7996,N_6666,N_6596);
nor U7997 (N_7997,N_6328,N_7218);
nor U7998 (N_7998,N_5548,N_5923);
or U7999 (N_7999,N_6562,N_6151);
and U8000 (N_8000,N_7338,N_6960);
xor U8001 (N_8001,N_7084,N_6010);
xnor U8002 (N_8002,N_6159,N_5677);
nor U8003 (N_8003,N_6434,N_6523);
or U8004 (N_8004,N_6279,N_6831);
xnor U8005 (N_8005,N_5279,N_5327);
nand U8006 (N_8006,N_5244,N_5425);
and U8007 (N_8007,N_7233,N_6494);
or U8008 (N_8008,N_7354,N_6063);
or U8009 (N_8009,N_7368,N_6517);
and U8010 (N_8010,N_6872,N_6229);
or U8011 (N_8011,N_7490,N_7495);
xor U8012 (N_8012,N_5471,N_5040);
or U8013 (N_8013,N_6314,N_7062);
nor U8014 (N_8014,N_5563,N_7373);
nor U8015 (N_8015,N_5691,N_6405);
or U8016 (N_8016,N_6916,N_5909);
or U8017 (N_8017,N_5207,N_5074);
nand U8018 (N_8018,N_6107,N_5746);
nor U8019 (N_8019,N_5300,N_6029);
nand U8020 (N_8020,N_6952,N_7413);
and U8021 (N_8021,N_5570,N_7122);
and U8022 (N_8022,N_5982,N_6439);
xor U8023 (N_8023,N_5436,N_5097);
nor U8024 (N_8024,N_6463,N_5002);
nor U8025 (N_8025,N_6964,N_5813);
xor U8026 (N_8026,N_6735,N_6431);
and U8027 (N_8027,N_5451,N_5780);
nand U8028 (N_8028,N_7051,N_6096);
xor U8029 (N_8029,N_7252,N_5682);
nand U8030 (N_8030,N_7229,N_6218);
nor U8031 (N_8031,N_7106,N_5726);
or U8032 (N_8032,N_6629,N_6698);
nand U8033 (N_8033,N_7049,N_5829);
nor U8034 (N_8034,N_6404,N_5383);
and U8035 (N_8035,N_7056,N_6381);
and U8036 (N_8036,N_7451,N_5190);
xnor U8037 (N_8037,N_7159,N_7200);
nor U8038 (N_8038,N_7420,N_6673);
nor U8039 (N_8039,N_6154,N_6382);
nor U8040 (N_8040,N_5388,N_7496);
nand U8041 (N_8041,N_7377,N_6475);
xnor U8042 (N_8042,N_5721,N_6257);
nand U8043 (N_8043,N_6921,N_6924);
nand U8044 (N_8044,N_5578,N_6000);
nand U8045 (N_8045,N_6282,N_7345);
nand U8046 (N_8046,N_5742,N_7225);
xnor U8047 (N_8047,N_6711,N_6346);
or U8048 (N_8048,N_6813,N_7464);
xor U8049 (N_8049,N_5800,N_6704);
or U8050 (N_8050,N_5904,N_5353);
and U8051 (N_8051,N_5874,N_6055);
and U8052 (N_8052,N_5745,N_7418);
xor U8053 (N_8053,N_5406,N_5396);
nand U8054 (N_8054,N_6469,N_7066);
nand U8055 (N_8055,N_7391,N_5990);
and U8056 (N_8056,N_5526,N_5809);
nor U8057 (N_8057,N_5626,N_5023);
nor U8058 (N_8058,N_7439,N_5265);
nor U8059 (N_8059,N_7328,N_6271);
or U8060 (N_8060,N_6858,N_6930);
and U8061 (N_8061,N_7046,N_5650);
xnor U8062 (N_8062,N_7408,N_7369);
or U8063 (N_8063,N_7281,N_5786);
xnor U8064 (N_8064,N_7168,N_6202);
xor U8065 (N_8065,N_5500,N_7450);
or U8066 (N_8066,N_6255,N_5758);
nor U8067 (N_8067,N_6676,N_6372);
nor U8068 (N_8068,N_5423,N_5958);
nand U8069 (N_8069,N_7210,N_6490);
or U8070 (N_8070,N_5330,N_7409);
xnor U8071 (N_8071,N_5116,N_5021);
nor U8072 (N_8072,N_6214,N_5386);
and U8073 (N_8073,N_7024,N_6614);
xnor U8074 (N_8074,N_5115,N_6197);
nor U8075 (N_8075,N_5274,N_6226);
xnor U8076 (N_8076,N_6811,N_6225);
nand U8077 (N_8077,N_5629,N_6812);
and U8078 (N_8078,N_6887,N_5364);
xor U8079 (N_8079,N_6254,N_6216);
nand U8080 (N_8080,N_5693,N_5695);
nand U8081 (N_8081,N_6077,N_7457);
or U8082 (N_8082,N_6358,N_5835);
and U8083 (N_8083,N_7427,N_6299);
or U8084 (N_8084,N_5542,N_6804);
or U8085 (N_8085,N_5172,N_6166);
or U8086 (N_8086,N_6410,N_7327);
nand U8087 (N_8087,N_5690,N_5577);
xnor U8088 (N_8088,N_7299,N_5873);
nor U8089 (N_8089,N_6194,N_5127);
xor U8090 (N_8090,N_6882,N_5296);
nor U8091 (N_8091,N_5494,N_7416);
or U8092 (N_8092,N_5150,N_5807);
nand U8093 (N_8093,N_7440,N_7272);
xnor U8094 (N_8094,N_5769,N_5319);
xor U8095 (N_8095,N_7460,N_7298);
nand U8096 (N_8096,N_7113,N_6331);
xor U8097 (N_8097,N_5711,N_6863);
and U8098 (N_8098,N_7077,N_7374);
or U8099 (N_8099,N_5832,N_5258);
nor U8100 (N_8100,N_5504,N_5671);
xnor U8101 (N_8101,N_6598,N_7167);
xnor U8102 (N_8102,N_5081,N_6899);
nor U8103 (N_8103,N_6348,N_5493);
or U8104 (N_8104,N_5286,N_6219);
nor U8105 (N_8105,N_6653,N_6277);
xor U8106 (N_8106,N_5462,N_6570);
nor U8107 (N_8107,N_7479,N_5155);
xor U8108 (N_8108,N_6725,N_6868);
nand U8109 (N_8109,N_6185,N_6958);
or U8110 (N_8110,N_6546,N_5799);
or U8111 (N_8111,N_5579,N_7208);
nand U8112 (N_8112,N_7164,N_7189);
nand U8113 (N_8113,N_5759,N_6662);
and U8114 (N_8114,N_7073,N_7431);
and U8115 (N_8115,N_5885,N_5437);
xor U8116 (N_8116,N_6241,N_6158);
and U8117 (N_8117,N_6915,N_7031);
and U8118 (N_8118,N_6430,N_5212);
or U8119 (N_8119,N_6513,N_6508);
nand U8120 (N_8120,N_5483,N_5727);
nor U8121 (N_8121,N_5315,N_5036);
and U8122 (N_8122,N_5910,N_5299);
and U8123 (N_8123,N_5082,N_6168);
or U8124 (N_8124,N_6902,N_5083);
or U8125 (N_8125,N_5592,N_5639);
nor U8126 (N_8126,N_5005,N_6948);
and U8127 (N_8127,N_6283,N_6131);
xnor U8128 (N_8128,N_7004,N_5496);
and U8129 (N_8129,N_5774,N_5257);
nor U8130 (N_8130,N_6619,N_6413);
xor U8131 (N_8131,N_6051,N_6658);
or U8132 (N_8132,N_5715,N_6556);
and U8133 (N_8133,N_7220,N_5943);
xnor U8134 (N_8134,N_6024,N_5595);
xor U8135 (N_8135,N_7193,N_7219);
or U8136 (N_8136,N_6669,N_6729);
xor U8137 (N_8137,N_7129,N_6036);
and U8138 (N_8138,N_7149,N_6180);
or U8139 (N_8139,N_6203,N_6816);
xnor U8140 (N_8140,N_6509,N_5565);
nand U8141 (N_8141,N_6940,N_5699);
or U8142 (N_8142,N_5638,N_5663);
nand U8143 (N_8143,N_5367,N_7216);
or U8144 (N_8144,N_6587,N_6586);
nor U8145 (N_8145,N_7055,N_6606);
or U8146 (N_8146,N_5101,N_6678);
nand U8147 (N_8147,N_5867,N_6963);
or U8148 (N_8148,N_6106,N_6496);
xnor U8149 (N_8149,N_6179,N_7076);
and U8150 (N_8150,N_6984,N_5053);
and U8151 (N_8151,N_5801,N_7291);
and U8152 (N_8152,N_5772,N_5114);
and U8153 (N_8153,N_5325,N_6933);
nand U8154 (N_8154,N_6826,N_6972);
or U8155 (N_8155,N_6712,N_6110);
xor U8156 (N_8156,N_7278,N_6623);
or U8157 (N_8157,N_6830,N_5530);
nand U8158 (N_8158,N_6270,N_5243);
or U8159 (N_8159,N_6655,N_5648);
nand U8160 (N_8160,N_5401,N_6777);
xnor U8161 (N_8161,N_6342,N_5863);
nor U8162 (N_8162,N_7396,N_7458);
xnor U8163 (N_8163,N_5239,N_7215);
xor U8164 (N_8164,N_5355,N_5204);
or U8165 (N_8165,N_6116,N_6022);
and U8166 (N_8166,N_5587,N_7241);
or U8167 (N_8167,N_6146,N_5952);
or U8168 (N_8168,N_7041,N_6819);
or U8169 (N_8169,N_7297,N_5089);
or U8170 (N_8170,N_5164,N_6768);
and U8171 (N_8171,N_6125,N_5154);
or U8172 (N_8172,N_5020,N_6575);
or U8173 (N_8173,N_6307,N_5108);
xnor U8174 (N_8174,N_7242,N_7067);
nor U8175 (N_8175,N_6126,N_6557);
nor U8176 (N_8176,N_5431,N_6710);
or U8177 (N_8177,N_6076,N_5883);
xnor U8178 (N_8178,N_5970,N_7191);
nor U8179 (N_8179,N_5184,N_7262);
nor U8180 (N_8180,N_6944,N_6518);
xor U8181 (N_8181,N_6075,N_5763);
and U8182 (N_8182,N_5918,N_5247);
and U8183 (N_8183,N_6436,N_6327);
or U8184 (N_8184,N_5506,N_5582);
nand U8185 (N_8185,N_5815,N_5612);
nor U8186 (N_8186,N_6968,N_6757);
xor U8187 (N_8187,N_7403,N_7197);
nand U8188 (N_8188,N_7438,N_7059);
or U8189 (N_8189,N_5767,N_5584);
nand U8190 (N_8190,N_7174,N_6260);
and U8191 (N_8191,N_5550,N_5804);
xnor U8192 (N_8192,N_6622,N_5156);
and U8193 (N_8193,N_5656,N_6374);
xor U8194 (N_8194,N_7389,N_5267);
and U8195 (N_8195,N_7339,N_5447);
nor U8196 (N_8196,N_5104,N_6708);
and U8197 (N_8197,N_6336,N_6604);
xor U8198 (N_8198,N_6262,N_6911);
xor U8199 (N_8199,N_6841,N_5263);
nor U8200 (N_8200,N_6787,N_7172);
and U8201 (N_8201,N_5209,N_5152);
nor U8202 (N_8202,N_5231,N_5657);
and U8203 (N_8203,N_6448,N_6927);
nor U8204 (N_8204,N_7071,N_6769);
nand U8205 (N_8205,N_6231,N_5424);
and U8206 (N_8206,N_6694,N_6387);
xnor U8207 (N_8207,N_6664,N_5945);
nor U8208 (N_8208,N_5460,N_6539);
nor U8209 (N_8209,N_6817,N_5415);
or U8210 (N_8210,N_6564,N_6827);
or U8211 (N_8211,N_5176,N_7481);
or U8212 (N_8212,N_5810,N_5345);
nand U8213 (N_8213,N_6663,N_5472);
nand U8214 (N_8214,N_6414,N_5649);
or U8215 (N_8215,N_6052,N_5994);
nand U8216 (N_8216,N_7029,N_7468);
nand U8217 (N_8217,N_5180,N_7039);
nor U8218 (N_8218,N_5762,N_5875);
or U8219 (N_8219,N_6791,N_6148);
nand U8220 (N_8220,N_7074,N_5881);
nor U8221 (N_8221,N_5273,N_5664);
or U8222 (N_8222,N_7125,N_7467);
xnor U8223 (N_8223,N_7295,N_5855);
xnor U8224 (N_8224,N_6042,N_6776);
nor U8225 (N_8225,N_5594,N_7211);
xor U8226 (N_8226,N_6170,N_5027);
nand U8227 (N_8227,N_7448,N_5749);
nand U8228 (N_8228,N_6864,N_6723);
nor U8229 (N_8229,N_6883,N_6810);
nand U8230 (N_8230,N_6701,N_5307);
nor U8231 (N_8231,N_7411,N_5441);
xnor U8232 (N_8232,N_6079,N_5631);
nand U8233 (N_8233,N_5949,N_5896);
and U8234 (N_8234,N_5482,N_5571);
or U8235 (N_8235,N_7472,N_5380);
or U8236 (N_8236,N_5882,N_6135);
xor U8237 (N_8237,N_5988,N_6320);
xnor U8238 (N_8238,N_6335,N_6097);
nand U8239 (N_8239,N_5163,N_7375);
nand U8240 (N_8240,N_5605,N_5015);
or U8241 (N_8241,N_6908,N_6937);
or U8242 (N_8242,N_5354,N_5285);
and U8243 (N_8243,N_5812,N_6310);
nand U8244 (N_8244,N_5057,N_5785);
and U8245 (N_8245,N_5316,N_6056);
nor U8246 (N_8246,N_5922,N_5528);
and U8247 (N_8247,N_6209,N_6545);
nand U8248 (N_8248,N_5138,N_5407);
or U8249 (N_8249,N_7271,N_5322);
nand U8250 (N_8250,N_5796,N_5124);
xor U8251 (N_8251,N_7003,N_7171);
or U8252 (N_8252,N_6169,N_6174);
and U8253 (N_8253,N_6132,N_5957);
or U8254 (N_8254,N_6035,N_6731);
nor U8255 (N_8255,N_5740,N_6196);
xnor U8256 (N_8256,N_7318,N_6303);
nor U8257 (N_8257,N_6198,N_6443);
and U8258 (N_8258,N_5160,N_5398);
or U8259 (N_8259,N_6238,N_6659);
xnor U8260 (N_8260,N_5336,N_5512);
and U8261 (N_8261,N_7177,N_7223);
and U8262 (N_8262,N_6006,N_6003);
nand U8263 (N_8263,N_6427,N_5440);
and U8264 (N_8264,N_6300,N_5586);
nor U8265 (N_8265,N_6466,N_6388);
or U8266 (N_8266,N_6175,N_6848);
and U8267 (N_8267,N_7379,N_6064);
nand U8268 (N_8268,N_6736,N_6965);
xor U8269 (N_8269,N_6516,N_6359);
nand U8270 (N_8270,N_7108,N_7437);
or U8271 (N_8271,N_6807,N_5573);
xnor U8272 (N_8272,N_6983,N_5689);
and U8273 (N_8273,N_5432,N_6938);
xor U8274 (N_8274,N_7035,N_5497);
and U8275 (N_8275,N_6559,N_6585);
xor U8276 (N_8276,N_5457,N_7016);
or U8277 (N_8277,N_6011,N_5927);
and U8278 (N_8278,N_5674,N_5320);
or U8279 (N_8279,N_5520,N_7492);
nor U8280 (N_8280,N_7202,N_5196);
or U8281 (N_8281,N_6491,N_6660);
xnor U8282 (N_8282,N_5683,N_6178);
nor U8283 (N_8283,N_5716,N_6975);
or U8284 (N_8284,N_6093,N_6967);
and U8285 (N_8285,N_6941,N_6128);
and U8286 (N_8286,N_7181,N_5376);
and U8287 (N_8287,N_7195,N_7355);
and U8288 (N_8288,N_7187,N_5611);
nor U8289 (N_8289,N_6265,N_6521);
and U8290 (N_8290,N_6977,N_7347);
and U8291 (N_8291,N_6313,N_6068);
nand U8292 (N_8292,N_5309,N_5044);
nor U8293 (N_8293,N_6543,N_6480);
and U8294 (N_8294,N_5604,N_7267);
nor U8295 (N_8295,N_5517,N_5470);
and U8296 (N_8296,N_5452,N_6281);
and U8297 (N_8297,N_7222,N_5269);
nand U8298 (N_8298,N_5931,N_6593);
nand U8299 (N_8299,N_7006,N_5210);
or U8300 (N_8300,N_5411,N_6290);
xor U8301 (N_8301,N_5948,N_5738);
nor U8302 (N_8302,N_5333,N_7407);
or U8303 (N_8303,N_7452,N_7268);
and U8304 (N_8304,N_7227,N_5940);
and U8305 (N_8305,N_5640,N_6053);
or U8306 (N_8306,N_6488,N_6422);
and U8307 (N_8307,N_5598,N_5748);
xor U8308 (N_8308,N_5821,N_5338);
or U8309 (N_8309,N_5444,N_6304);
and U8310 (N_8310,N_6173,N_6665);
or U8311 (N_8311,N_6134,N_6040);
xnor U8312 (N_8312,N_6020,N_6657);
and U8313 (N_8313,N_6489,N_7028);
and U8314 (N_8314,N_5734,N_6691);
nand U8315 (N_8315,N_7259,N_5658);
nand U8316 (N_8316,N_6376,N_7206);
and U8317 (N_8317,N_6375,N_6306);
nand U8318 (N_8318,N_5744,N_7151);
and U8319 (N_8319,N_6782,N_7454);
or U8320 (N_8320,N_5059,N_6428);
or U8321 (N_8321,N_6091,N_6778);
nand U8322 (N_8322,N_5514,N_6041);
xnor U8323 (N_8323,N_5572,N_6605);
or U8324 (N_8324,N_5898,N_6233);
or U8325 (N_8325,N_5043,N_7398);
nand U8326 (N_8326,N_7349,N_6547);
xnor U8327 (N_8327,N_6421,N_7317);
or U8328 (N_8328,N_6246,N_7380);
xor U8329 (N_8329,N_5562,N_5533);
xor U8330 (N_8330,N_6130,N_6234);
xnor U8331 (N_8331,N_5971,N_6837);
nor U8332 (N_8332,N_5635,N_7061);
nor U8333 (N_8333,N_5303,N_7050);
nor U8334 (N_8334,N_7085,N_6379);
nand U8335 (N_8335,N_5585,N_6183);
or U8336 (N_8336,N_5531,N_7019);
xor U8337 (N_8337,N_5242,N_5646);
and U8338 (N_8338,N_6640,N_5283);
and U8339 (N_8339,N_6633,N_6688);
nor U8340 (N_8340,N_5600,N_5672);
xor U8341 (N_8341,N_6537,N_7001);
or U8342 (N_8342,N_5553,N_7436);
or U8343 (N_8343,N_6393,N_6186);
nor U8344 (N_8344,N_5012,N_7072);
and U8345 (N_8345,N_5014,N_7045);
nor U8346 (N_8346,N_5480,N_5679);
nand U8347 (N_8347,N_5614,N_7176);
nand U8348 (N_8348,N_6351,N_6268);
or U8349 (N_8349,N_6724,N_7178);
and U8350 (N_8350,N_5778,N_6252);
nor U8351 (N_8351,N_5417,N_6483);
xor U8352 (N_8352,N_7161,N_5893);
xor U8353 (N_8353,N_5465,N_7334);
and U8354 (N_8354,N_6715,N_5932);
nor U8355 (N_8355,N_7163,N_7015);
or U8356 (N_8356,N_5706,N_5232);
nor U8357 (N_8357,N_5633,N_5485);
and U8358 (N_8358,N_6918,N_6624);
and U8359 (N_8359,N_7224,N_6687);
and U8360 (N_8360,N_6136,N_5208);
or U8361 (N_8361,N_5637,N_5393);
or U8362 (N_8362,N_7312,N_6990);
nand U8363 (N_8363,N_6522,N_6207);
nand U8364 (N_8364,N_5238,N_5985);
or U8365 (N_8365,N_7112,N_6818);
or U8366 (N_8366,N_5973,N_6719);
xor U8367 (N_8367,N_6648,N_6697);
and U8368 (N_8368,N_6969,N_5527);
and U8369 (N_8369,N_7456,N_7236);
nand U8370 (N_8370,N_6670,N_6325);
and U8371 (N_8371,N_5766,N_6222);
or U8372 (N_8372,N_6420,N_6609);
or U8373 (N_8373,N_5569,N_5853);
xnor U8374 (N_8374,N_5802,N_6322);
xor U8375 (N_8375,N_5890,N_6514);
or U8376 (N_8376,N_6008,N_6498);
nand U8377 (N_8377,N_6885,N_6718);
nand U8378 (N_8378,N_6145,N_5000);
nand U8379 (N_8379,N_5852,N_5035);
nor U8380 (N_8380,N_5421,N_6845);
or U8381 (N_8381,N_6821,N_5357);
or U8382 (N_8382,N_6836,N_6293);
nand U8383 (N_8383,N_7092,N_5921);
nor U8384 (N_8384,N_6094,N_5887);
xnor U8385 (N_8385,N_5859,N_5580);
nand U8386 (N_8386,N_5439,N_5228);
nor U8387 (N_8387,N_6378,N_7052);
and U8388 (N_8388,N_5628,N_7025);
or U8389 (N_8389,N_6832,N_7274);
or U8390 (N_8390,N_7261,N_6825);
xnor U8391 (N_8391,N_6009,N_5302);
nor U8392 (N_8392,N_6955,N_7285);
or U8393 (N_8393,N_5477,N_5654);
nor U8394 (N_8394,N_5632,N_5294);
or U8395 (N_8395,N_5817,N_5216);
xnor U8396 (N_8396,N_7428,N_5250);
xnor U8397 (N_8397,N_6884,N_6839);
and U8398 (N_8398,N_7140,N_5916);
xor U8399 (N_8399,N_6540,N_5636);
or U8400 (N_8400,N_5865,N_6432);
xnor U8401 (N_8401,N_6682,N_6449);
nand U8402 (N_8402,N_5276,N_7260);
or U8403 (N_8403,N_5736,N_5942);
nor U8404 (N_8404,N_7386,N_6017);
and U8405 (N_8405,N_5729,N_6400);
nor U8406 (N_8406,N_6401,N_5134);
nor U8407 (N_8407,N_5328,N_5445);
or U8408 (N_8408,N_5956,N_6957);
or U8409 (N_8409,N_7162,N_5223);
and U8410 (N_8410,N_7021,N_7204);
xor U8411 (N_8411,N_5446,N_6803);
and U8412 (N_8412,N_6292,N_6341);
nand U8413 (N_8413,N_6156,N_5169);
or U8414 (N_8414,N_5130,N_5435);
nor U8415 (N_8415,N_6472,N_7363);
or U8416 (N_8416,N_5403,N_6429);
and U8417 (N_8417,N_5361,N_6023);
nand U8418 (N_8418,N_6153,N_7352);
or U8419 (N_8419,N_7155,N_7265);
nand U8420 (N_8420,N_6189,N_5575);
and U8421 (N_8421,N_5119,N_5476);
nor U8422 (N_8422,N_6714,N_6470);
nor U8423 (N_8423,N_5755,N_7390);
nand U8424 (N_8424,N_5003,N_6468);
or U8425 (N_8425,N_7096,N_6935);
nand U8426 (N_8426,N_5129,N_5697);
or U8427 (N_8427,N_5050,N_7080);
xnor U8428 (N_8428,N_7244,N_7126);
nor U8429 (N_8429,N_5798,N_5148);
nand U8430 (N_8430,N_6456,N_5980);
or U8431 (N_8431,N_7469,N_5182);
xnor U8432 (N_8432,N_5583,N_5886);
nor U8433 (N_8433,N_5203,N_5913);
nand U8434 (N_8434,N_7342,N_6150);
and U8435 (N_8435,N_5915,N_5215);
and U8436 (N_8436,N_7230,N_7444);
nand U8437 (N_8437,N_5567,N_5647);
xor U8438 (N_8438,N_6349,N_6418);
or U8439 (N_8439,N_6333,N_7290);
xnor U8440 (N_8440,N_7286,N_5306);
nor U8441 (N_8441,N_7491,N_6503);
xor U8442 (N_8442,N_5259,N_5978);
or U8443 (N_8443,N_6716,N_5120);
xor U8444 (N_8444,N_5984,N_6291);
xor U8445 (N_8445,N_5400,N_5665);
and U8446 (N_8446,N_5230,N_5756);
nand U8447 (N_8447,N_6251,N_6235);
or U8448 (N_8448,N_6560,N_6160);
and U8449 (N_8449,N_6486,N_7124);
and U8450 (N_8450,N_5735,N_5293);
nand U8451 (N_8451,N_5965,N_7123);
nand U8452 (N_8452,N_5205,N_5849);
xnor U8453 (N_8453,N_6632,N_5966);
or U8454 (N_8454,N_6854,N_6751);
nand U8455 (N_8455,N_5794,N_6683);
nand U8456 (N_8456,N_5187,N_6652);
and U8457 (N_8457,N_6840,N_5085);
nor U8458 (N_8458,N_5975,N_7121);
xor U8459 (N_8459,N_6765,N_7273);
and U8460 (N_8460,N_7115,N_5969);
nand U8461 (N_8461,N_5787,N_6834);
and U8462 (N_8462,N_6894,N_7376);
nand U8463 (N_8463,N_6505,N_7364);
xor U8464 (N_8464,N_7441,N_5499);
nor U8465 (N_8465,N_5938,N_5871);
nor U8466 (N_8466,N_5271,N_6956);
and U8467 (N_8467,N_7498,N_5395);
or U8468 (N_8468,N_7169,N_5508);
xnor U8469 (N_8469,N_6043,N_5856);
xor U8470 (N_8470,N_5045,N_5173);
xnor U8471 (N_8471,N_5323,N_5591);
nor U8472 (N_8472,N_6061,N_7381);
xor U8473 (N_8473,N_5091,N_6922);
or U8474 (N_8474,N_5404,N_6124);
xor U8475 (N_8475,N_6996,N_6444);
and U8476 (N_8476,N_6627,N_5139);
and U8477 (N_8477,N_5428,N_5199);
nor U8478 (N_8478,N_5644,N_5872);
and U8479 (N_8479,N_7497,N_5229);
xor U8480 (N_8480,N_6278,N_7232);
xnor U8481 (N_8481,N_6493,N_6147);
xor U8482 (N_8482,N_6100,N_5341);
xnor U8483 (N_8483,N_5492,N_7146);
xnor U8484 (N_8484,N_5475,N_5951);
nor U8485 (N_8485,N_7442,N_7170);
nor U8486 (N_8486,N_6057,N_5981);
nor U8487 (N_8487,N_7228,N_7111);
xor U8488 (N_8488,N_5378,N_5042);
nor U8489 (N_8489,N_6579,N_7239);
and U8490 (N_8490,N_5564,N_5183);
and U8491 (N_8491,N_6690,N_6828);
and U8492 (N_8492,N_5028,N_6934);
xor U8493 (N_8493,N_5434,N_7321);
nor U8494 (N_8494,N_6617,N_6357);
or U8495 (N_8495,N_5820,N_5076);
nor U8496 (N_8496,N_6895,N_6926);
nand U8497 (N_8497,N_5068,N_6471);
and U8498 (N_8498,N_5808,N_6280);
nor U8499 (N_8499,N_6741,N_5939);
and U8500 (N_8500,N_7470,N_5371);
nand U8501 (N_8501,N_7002,N_7020);
and U8502 (N_8502,N_7238,N_5458);
xor U8503 (N_8503,N_7393,N_7132);
xnor U8504 (N_8504,N_5185,N_7089);
xnor U8505 (N_8505,N_5620,N_7198);
nand U8506 (N_8506,N_5385,N_5793);
and U8507 (N_8507,N_6519,N_5387);
nor U8508 (N_8508,N_5225,N_6734);
nand U8509 (N_8509,N_7192,N_7269);
nand U8510 (N_8510,N_6852,N_5427);
xor U8511 (N_8511,N_6269,N_5536);
nor U8512 (N_8512,N_6613,N_6775);
or U8513 (N_8513,N_7183,N_6284);
nor U8514 (N_8514,N_6315,N_6566);
xor U8515 (N_8515,N_5509,N_7446);
nor U8516 (N_8516,N_5055,N_7022);
xor U8517 (N_8517,N_5557,N_5236);
and U8518 (N_8518,N_7064,N_7173);
and U8519 (N_8519,N_6713,N_6620);
or U8520 (N_8520,N_5838,N_7335);
or U8521 (N_8521,N_7417,N_6550);
and U8522 (N_8522,N_5468,N_5964);
nand U8523 (N_8523,N_5111,N_7447);
xor U8524 (N_8524,N_5712,N_6361);
and U8525 (N_8525,N_7217,N_5836);
or U8526 (N_8526,N_7188,N_6876);
or U8527 (N_8527,N_7158,N_5652);
xor U8528 (N_8528,N_5275,N_5168);
nor U8529 (N_8529,N_6223,N_5092);
nor U8530 (N_8530,N_5069,N_7424);
nor U8531 (N_8531,N_6031,N_6805);
and U8532 (N_8532,N_6538,N_5060);
and U8533 (N_8533,N_5131,N_7247);
nand U8534 (N_8534,N_5194,N_5095);
and U8535 (N_8535,N_5696,N_6407);
xor U8536 (N_8536,N_6193,N_6679);
xor U8537 (N_8537,N_5701,N_5133);
nor U8538 (N_8538,N_5680,N_7196);
nor U8539 (N_8539,N_6650,N_5007);
nor U8540 (N_8540,N_5704,N_6802);
and U8541 (N_8541,N_5770,N_6019);
or U8542 (N_8542,N_6512,N_5621);
nor U8543 (N_8543,N_7053,N_7348);
or U8544 (N_8544,N_6820,N_7231);
and U8545 (N_8545,N_6767,N_5374);
or U8546 (N_8546,N_7119,N_7399);
xor U8547 (N_8547,N_5962,N_5128);
and U8548 (N_8548,N_5919,N_5268);
and U8549 (N_8549,N_6474,N_5146);
nand U8550 (N_8550,N_6383,N_7323);
nand U8551 (N_8551,N_5540,N_7133);
and U8552 (N_8552,N_6686,N_5094);
xnor U8553 (N_8553,N_6163,N_7325);
and U8554 (N_8554,N_6636,N_6583);
nand U8555 (N_8555,N_5240,N_5013);
and U8556 (N_8556,N_7473,N_5352);
and U8557 (N_8557,N_6792,N_5737);
nand U8558 (N_8558,N_5370,N_5515);
nor U8559 (N_8559,N_6800,N_5255);
or U8560 (N_8560,N_6784,N_7221);
or U8561 (N_8561,N_7384,N_6888);
or U8562 (N_8562,N_5298,N_6581);
xor U8563 (N_8563,N_6347,N_7128);
xnor U8564 (N_8564,N_5394,N_7343);
nor U8565 (N_8565,N_6485,N_6289);
xor U8566 (N_8566,N_7412,N_6221);
or U8567 (N_8567,N_6989,N_5535);
xnor U8568 (N_8568,N_7337,N_7410);
nor U8569 (N_8569,N_5149,N_7017);
or U8570 (N_8570,N_6426,N_6618);
nor U8571 (N_8571,N_6236,N_5773);
xor U8572 (N_8572,N_5109,N_5343);
or U8573 (N_8573,N_6542,N_6014);
xor U8574 (N_8574,N_5193,N_6625);
nand U8575 (N_8575,N_5246,N_5195);
xor U8576 (N_8576,N_7165,N_6638);
and U8577 (N_8577,N_7372,N_7359);
xor U8578 (N_8578,N_5227,N_5692);
nand U8579 (N_8579,N_5179,N_7185);
xnor U8580 (N_8580,N_5687,N_5217);
nand U8581 (N_8581,N_6098,N_6615);
or U8582 (N_8582,N_5627,N_5075);
xnor U8583 (N_8583,N_5041,N_5381);
and U8584 (N_8584,N_6311,N_5764);
nand U8585 (N_8585,N_5850,N_6737);
nor U8586 (N_8586,N_6089,N_5413);
nor U8587 (N_8587,N_6789,N_6244);
nand U8588 (N_8588,N_6177,N_7350);
nand U8589 (N_8589,N_5609,N_6897);
nand U8590 (N_8590,N_7275,N_6182);
and U8591 (N_8591,N_7145,N_6572);
nor U8592 (N_8592,N_5135,N_6195);
nor U8593 (N_8593,N_6157,N_5722);
and U8594 (N_8594,N_6033,N_6853);
nand U8595 (N_8595,N_7292,N_7054);
nand U8596 (N_8596,N_6212,N_5864);
xnor U8597 (N_8597,N_6103,N_7243);
nor U8598 (N_8598,N_5136,N_6457);
nor U8599 (N_8599,N_6080,N_6738);
nand U8600 (N_8600,N_7148,N_6881);
xor U8601 (N_8601,N_5372,N_6034);
or U8602 (N_8602,N_6026,N_5018);
xor U8603 (N_8603,N_5634,N_6532);
xnor U8604 (N_8604,N_6455,N_6105);
nand U8605 (N_8605,N_6021,N_7478);
or U8606 (N_8606,N_5070,N_6090);
nor U8607 (N_8607,N_7485,N_7141);
nor U8608 (N_8608,N_5823,N_6380);
and U8609 (N_8609,N_5889,N_6525);
or U8610 (N_8610,N_7361,N_6139);
xor U8611 (N_8611,N_5340,N_6910);
nand U8612 (N_8612,N_6122,N_6030);
xor U8613 (N_8613,N_6409,N_6353);
xnor U8614 (N_8614,N_6138,N_7419);
or U8615 (N_8615,N_5532,N_5110);
xor U8616 (N_8616,N_5556,N_6582);
nand U8617 (N_8617,N_7142,N_6458);
or U8618 (N_8618,N_5304,N_6913);
or U8619 (N_8619,N_6595,N_7484);
and U8620 (N_8620,N_6520,N_7382);
xnor U8621 (N_8621,N_7081,N_5189);
nand U8622 (N_8622,N_5241,N_6476);
or U8623 (N_8623,N_6896,N_5844);
or U8624 (N_8624,N_5064,N_6417);
or U8625 (N_8625,N_7034,N_5072);
xor U8626 (N_8626,N_7277,N_5348);
or U8627 (N_8627,N_6759,N_7405);
nand U8628 (N_8628,N_5295,N_5301);
nand U8629 (N_8629,N_7038,N_6133);
or U8630 (N_8630,N_5219,N_7209);
and U8631 (N_8631,N_5489,N_5840);
or U8632 (N_8632,N_6242,N_6149);
nand U8633 (N_8633,N_6637,N_5331);
nor U8634 (N_8634,N_6561,N_5491);
nand U8635 (N_8635,N_7240,N_6597);
nor U8636 (N_8636,N_7179,N_5261);
or U8637 (N_8637,N_7421,N_5096);
or U8638 (N_8638,N_6750,N_5928);
nor U8639 (N_8639,N_7314,N_5845);
xor U8640 (N_8640,N_5334,N_6641);
nand U8641 (N_8641,N_6499,N_5112);
nor U8642 (N_8642,N_6045,N_6397);
nand U8643 (N_8643,N_6766,N_5552);
nor U8644 (N_8644,N_7182,N_5080);
xnor U8645 (N_8645,N_7214,N_6541);
and U8646 (N_8646,N_5615,N_5724);
nand U8647 (N_8647,N_6634,N_6176);
nor U8648 (N_8648,N_5743,N_5379);
nor U8649 (N_8649,N_7139,N_6484);
nor U8650 (N_8650,N_5197,N_6188);
xnor U8651 (N_8651,N_7201,N_6070);
xnor U8652 (N_8652,N_6206,N_7255);
nand U8653 (N_8653,N_6809,N_5312);
nand U8654 (N_8654,N_6237,N_6689);
and U8655 (N_8655,N_6584,N_5559);
nor U8656 (N_8656,N_6344,N_6573);
nand U8657 (N_8657,N_5188,N_5416);
nor U8658 (N_8658,N_7094,N_6302);
and U8659 (N_8659,N_5511,N_5765);
or U8660 (N_8660,N_5987,N_7366);
and U8661 (N_8661,N_6046,N_5545);
and U8662 (N_8662,N_6588,N_6435);
xnor U8663 (N_8663,N_5086,N_5412);
xnor U8664 (N_8664,N_5934,N_7109);
xor U8665 (N_8665,N_5513,N_5920);
xor U8666 (N_8666,N_7060,N_5768);
or U8667 (N_8667,N_5317,N_5001);
nor U8668 (N_8668,N_5754,N_6680);
nor U8669 (N_8669,N_6205,N_6208);
xor U8670 (N_8670,N_7429,N_7127);
xnor U8671 (N_8671,N_7282,N_5161);
and U8672 (N_8672,N_5466,N_5502);
nand U8673 (N_8673,N_6567,N_6954);
and U8674 (N_8674,N_5997,N_5979);
or U8675 (N_8675,N_6576,N_5008);
or U8676 (N_8676,N_5576,N_7138);
nand U8677 (N_8677,N_5653,N_6551);
xor U8678 (N_8678,N_5946,N_6266);
xnor U8679 (N_8679,N_5618,N_5151);
or U8680 (N_8680,N_7153,N_6445);
nand U8681 (N_8681,N_6685,N_5103);
nand U8682 (N_8682,N_5066,N_7356);
and U8683 (N_8683,N_7434,N_7057);
nand U8684 (N_8684,N_7308,N_6667);
nor U8685 (N_8685,N_5846,N_5668);
or U8686 (N_8686,N_6835,N_5166);
and U8687 (N_8687,N_6162,N_5995);
xnor U8688 (N_8688,N_5022,N_5201);
nand U8689 (N_8689,N_5622,N_7433);
and U8690 (N_8690,N_5220,N_5377);
nand U8691 (N_8691,N_6762,N_6527);
or U8692 (N_8692,N_5046,N_5538);
nand U8693 (N_8693,N_7344,N_5929);
xnor U8694 (N_8694,N_6171,N_6258);
and U8695 (N_8695,N_6497,N_5260);
nor U8696 (N_8696,N_6454,N_5589);
and U8697 (N_8697,N_6869,N_7395);
or U8698 (N_8698,N_5643,N_6747);
and U8699 (N_8699,N_5488,N_5790);
xor U8700 (N_8700,N_5233,N_5170);
and U8701 (N_8701,N_5318,N_6643);
nor U8702 (N_8702,N_5684,N_6360);
or U8703 (N_8703,N_6316,N_6371);
nand U8704 (N_8704,N_6013,N_6886);
nor U8705 (N_8705,N_7135,N_5245);
nand U8706 (N_8706,N_6929,N_5256);
nand U8707 (N_8707,N_5332,N_6312);
or U8708 (N_8708,N_5177,N_6018);
nand U8709 (N_8709,N_5541,N_6164);
or U8710 (N_8710,N_5895,N_7027);
and U8711 (N_8711,N_6578,N_5675);
nor U8712 (N_8712,N_7047,N_6914);
or U8713 (N_8713,N_5963,N_6191);
nor U8714 (N_8714,N_5906,N_5165);
and U8715 (N_8715,N_7425,N_7088);
or U8716 (N_8716,N_5073,N_6095);
or U8717 (N_8717,N_6847,N_6001);
xnor U8718 (N_8718,N_6329,N_7353);
or U8719 (N_8719,N_5900,N_5660);
nor U8720 (N_8720,N_6611,N_5034);
and U8721 (N_8721,N_6369,N_6442);
or U8722 (N_8722,N_5024,N_6161);
nor U8723 (N_8723,N_6273,N_6165);
and U8724 (N_8724,N_5402,N_7426);
nand U8725 (N_8725,N_7226,N_5543);
and U8726 (N_8726,N_5448,N_5032);
and U8727 (N_8727,N_7296,N_7367);
nor U8728 (N_8728,N_5481,N_6721);
nand U8729 (N_8729,N_5461,N_6865);
and U8730 (N_8730,N_6661,N_7008);
nor U8731 (N_8731,N_5102,N_6419);
nor U8732 (N_8732,N_5826,N_7351);
and U8733 (N_8733,N_7036,N_6099);
and U8734 (N_8734,N_5360,N_6796);
xor U8735 (N_8735,N_7069,N_6285);
nor U8736 (N_8736,N_6814,N_5047);
or U8737 (N_8737,N_5861,N_5026);
and U8738 (N_8738,N_6991,N_6779);
nand U8739 (N_8739,N_7079,N_5516);
xnor U8740 (N_8740,N_6534,N_6823);
nor U8741 (N_8741,N_5933,N_7264);
and U8742 (N_8742,N_6974,N_6677);
nor U8743 (N_8743,N_6118,N_7304);
and U8744 (N_8744,N_6917,N_7166);
or U8745 (N_8745,N_5566,N_7152);
nor U8746 (N_8746,N_7371,N_7120);
nor U8747 (N_8747,N_6259,N_7320);
nand U8748 (N_8748,N_6084,N_6391);
xnor U8749 (N_8749,N_7466,N_6396);
and U8750 (N_8750,N_6469,N_5689);
xor U8751 (N_8751,N_5315,N_5978);
xor U8752 (N_8752,N_6657,N_6748);
xnor U8753 (N_8753,N_6247,N_6244);
nor U8754 (N_8754,N_5003,N_6185);
or U8755 (N_8755,N_7120,N_6015);
nor U8756 (N_8756,N_5433,N_5767);
nand U8757 (N_8757,N_6969,N_7163);
or U8758 (N_8758,N_5427,N_5428);
nand U8759 (N_8759,N_6940,N_6966);
nand U8760 (N_8760,N_6642,N_5767);
nor U8761 (N_8761,N_6022,N_5668);
nand U8762 (N_8762,N_5485,N_5840);
nand U8763 (N_8763,N_7043,N_5749);
or U8764 (N_8764,N_5027,N_6971);
or U8765 (N_8765,N_7049,N_7347);
nor U8766 (N_8766,N_5224,N_6089);
nand U8767 (N_8767,N_5341,N_6800);
and U8768 (N_8768,N_6019,N_7404);
nor U8769 (N_8769,N_6191,N_5864);
nor U8770 (N_8770,N_7460,N_5664);
nor U8771 (N_8771,N_7406,N_5425);
nor U8772 (N_8772,N_6925,N_7301);
nand U8773 (N_8773,N_5162,N_6839);
nand U8774 (N_8774,N_6755,N_5862);
and U8775 (N_8775,N_5228,N_7414);
nand U8776 (N_8776,N_5919,N_5057);
and U8777 (N_8777,N_6944,N_7101);
or U8778 (N_8778,N_6497,N_5023);
and U8779 (N_8779,N_6239,N_7120);
or U8780 (N_8780,N_6047,N_5321);
nor U8781 (N_8781,N_5958,N_6742);
and U8782 (N_8782,N_7332,N_6423);
and U8783 (N_8783,N_5846,N_5000);
or U8784 (N_8784,N_6196,N_6484);
and U8785 (N_8785,N_5766,N_5147);
xor U8786 (N_8786,N_5138,N_6051);
nand U8787 (N_8787,N_6768,N_7024);
and U8788 (N_8788,N_5892,N_5351);
and U8789 (N_8789,N_5989,N_7173);
xnor U8790 (N_8790,N_6417,N_7439);
or U8791 (N_8791,N_5666,N_6513);
and U8792 (N_8792,N_5744,N_7314);
nand U8793 (N_8793,N_5357,N_7474);
xor U8794 (N_8794,N_7444,N_6941);
nor U8795 (N_8795,N_5695,N_6200);
or U8796 (N_8796,N_6647,N_6755);
nor U8797 (N_8797,N_6764,N_5344);
xnor U8798 (N_8798,N_6637,N_6149);
nand U8799 (N_8799,N_7048,N_5845);
nor U8800 (N_8800,N_6687,N_5096);
or U8801 (N_8801,N_6040,N_5821);
nor U8802 (N_8802,N_5130,N_6560);
xor U8803 (N_8803,N_5875,N_6233);
xnor U8804 (N_8804,N_7116,N_6372);
nand U8805 (N_8805,N_7229,N_6298);
nor U8806 (N_8806,N_6469,N_7492);
and U8807 (N_8807,N_6388,N_7000);
or U8808 (N_8808,N_5816,N_6704);
nor U8809 (N_8809,N_5198,N_6217);
nand U8810 (N_8810,N_7200,N_6372);
xor U8811 (N_8811,N_6605,N_7379);
nand U8812 (N_8812,N_7484,N_5516);
nand U8813 (N_8813,N_6964,N_6430);
nor U8814 (N_8814,N_5444,N_7471);
and U8815 (N_8815,N_6832,N_5972);
nand U8816 (N_8816,N_6646,N_6817);
nand U8817 (N_8817,N_6002,N_7465);
nor U8818 (N_8818,N_6624,N_6751);
nand U8819 (N_8819,N_6534,N_6512);
and U8820 (N_8820,N_7276,N_7293);
or U8821 (N_8821,N_6810,N_5091);
or U8822 (N_8822,N_7347,N_6780);
xnor U8823 (N_8823,N_5645,N_5587);
or U8824 (N_8824,N_6437,N_6951);
xor U8825 (N_8825,N_5327,N_5703);
or U8826 (N_8826,N_6479,N_5988);
nor U8827 (N_8827,N_5047,N_6177);
and U8828 (N_8828,N_5856,N_5807);
xor U8829 (N_8829,N_5971,N_7110);
and U8830 (N_8830,N_6880,N_6739);
and U8831 (N_8831,N_6738,N_7283);
or U8832 (N_8832,N_6688,N_7186);
xor U8833 (N_8833,N_5452,N_7279);
and U8834 (N_8834,N_5159,N_5126);
xnor U8835 (N_8835,N_5332,N_7407);
or U8836 (N_8836,N_6609,N_6422);
nor U8837 (N_8837,N_7457,N_6789);
or U8838 (N_8838,N_5966,N_6532);
nand U8839 (N_8839,N_5042,N_6684);
or U8840 (N_8840,N_5762,N_6593);
xor U8841 (N_8841,N_5702,N_7446);
nand U8842 (N_8842,N_6674,N_6471);
and U8843 (N_8843,N_6056,N_7276);
and U8844 (N_8844,N_5847,N_6013);
or U8845 (N_8845,N_6791,N_6707);
nand U8846 (N_8846,N_6094,N_7236);
xnor U8847 (N_8847,N_5303,N_7022);
and U8848 (N_8848,N_5119,N_6725);
and U8849 (N_8849,N_5445,N_5049);
or U8850 (N_8850,N_5138,N_6751);
xnor U8851 (N_8851,N_7082,N_6091);
or U8852 (N_8852,N_6102,N_6536);
or U8853 (N_8853,N_6453,N_5459);
nand U8854 (N_8854,N_6021,N_6020);
and U8855 (N_8855,N_5751,N_5684);
and U8856 (N_8856,N_6323,N_6541);
and U8857 (N_8857,N_5285,N_5149);
nor U8858 (N_8858,N_5701,N_7126);
and U8859 (N_8859,N_5370,N_6180);
or U8860 (N_8860,N_5939,N_6584);
xor U8861 (N_8861,N_7366,N_6470);
nor U8862 (N_8862,N_6725,N_6165);
or U8863 (N_8863,N_5683,N_5737);
and U8864 (N_8864,N_6363,N_5028);
xnor U8865 (N_8865,N_5154,N_7482);
or U8866 (N_8866,N_6179,N_6013);
nor U8867 (N_8867,N_5016,N_6459);
or U8868 (N_8868,N_5467,N_5160);
xnor U8869 (N_8869,N_6437,N_5095);
nor U8870 (N_8870,N_6197,N_6961);
or U8871 (N_8871,N_5806,N_6880);
xnor U8872 (N_8872,N_7175,N_5258);
xor U8873 (N_8873,N_6058,N_6206);
xnor U8874 (N_8874,N_6966,N_5762);
and U8875 (N_8875,N_6494,N_5837);
nor U8876 (N_8876,N_5515,N_5308);
nor U8877 (N_8877,N_6297,N_5134);
or U8878 (N_8878,N_5189,N_5724);
and U8879 (N_8879,N_6014,N_6294);
nor U8880 (N_8880,N_5853,N_5069);
nand U8881 (N_8881,N_6935,N_6437);
and U8882 (N_8882,N_7037,N_6389);
nor U8883 (N_8883,N_5574,N_6336);
nor U8884 (N_8884,N_7261,N_5717);
nor U8885 (N_8885,N_5635,N_7462);
nand U8886 (N_8886,N_5201,N_6943);
and U8887 (N_8887,N_5570,N_5723);
and U8888 (N_8888,N_5662,N_5841);
nor U8889 (N_8889,N_6686,N_5267);
or U8890 (N_8890,N_7010,N_5855);
xnor U8891 (N_8891,N_6267,N_5590);
xor U8892 (N_8892,N_5335,N_6733);
and U8893 (N_8893,N_6864,N_7128);
nand U8894 (N_8894,N_6767,N_5566);
xor U8895 (N_8895,N_6477,N_7061);
nand U8896 (N_8896,N_7315,N_5153);
and U8897 (N_8897,N_7455,N_7323);
xnor U8898 (N_8898,N_5494,N_6105);
or U8899 (N_8899,N_7008,N_5832);
or U8900 (N_8900,N_6291,N_6369);
xor U8901 (N_8901,N_6235,N_6228);
xor U8902 (N_8902,N_5137,N_5452);
or U8903 (N_8903,N_5603,N_6209);
xor U8904 (N_8904,N_5290,N_6338);
nor U8905 (N_8905,N_6510,N_5878);
xnor U8906 (N_8906,N_6460,N_6007);
or U8907 (N_8907,N_7106,N_5785);
and U8908 (N_8908,N_7178,N_5382);
or U8909 (N_8909,N_7291,N_6228);
and U8910 (N_8910,N_6937,N_5645);
and U8911 (N_8911,N_7377,N_5281);
xnor U8912 (N_8912,N_5180,N_6708);
nand U8913 (N_8913,N_6227,N_7341);
and U8914 (N_8914,N_6603,N_6537);
or U8915 (N_8915,N_6457,N_7323);
xor U8916 (N_8916,N_6155,N_5638);
and U8917 (N_8917,N_6373,N_7207);
xor U8918 (N_8918,N_6842,N_6673);
and U8919 (N_8919,N_6970,N_6042);
and U8920 (N_8920,N_5811,N_6846);
nor U8921 (N_8921,N_5063,N_5396);
nand U8922 (N_8922,N_6131,N_5394);
nor U8923 (N_8923,N_7292,N_7463);
nand U8924 (N_8924,N_6601,N_5193);
and U8925 (N_8925,N_7096,N_7100);
nand U8926 (N_8926,N_6248,N_5013);
nand U8927 (N_8927,N_7298,N_5056);
xnor U8928 (N_8928,N_5071,N_5120);
xor U8929 (N_8929,N_7393,N_5977);
nand U8930 (N_8930,N_7129,N_5085);
and U8931 (N_8931,N_6929,N_7279);
nand U8932 (N_8932,N_5285,N_5513);
nand U8933 (N_8933,N_5920,N_7025);
nand U8934 (N_8934,N_7490,N_6552);
xor U8935 (N_8935,N_7154,N_6170);
nor U8936 (N_8936,N_5936,N_6352);
xor U8937 (N_8937,N_5880,N_6878);
and U8938 (N_8938,N_5396,N_5536);
and U8939 (N_8939,N_5714,N_6376);
xnor U8940 (N_8940,N_6408,N_5424);
xnor U8941 (N_8941,N_6082,N_5349);
and U8942 (N_8942,N_5239,N_6107);
nand U8943 (N_8943,N_5177,N_6105);
or U8944 (N_8944,N_7370,N_6259);
or U8945 (N_8945,N_6106,N_5142);
nor U8946 (N_8946,N_7088,N_6104);
xnor U8947 (N_8947,N_6752,N_5722);
and U8948 (N_8948,N_5753,N_7150);
nor U8949 (N_8949,N_6068,N_5229);
nor U8950 (N_8950,N_5448,N_6221);
or U8951 (N_8951,N_6329,N_7027);
and U8952 (N_8952,N_5627,N_6335);
nor U8953 (N_8953,N_6483,N_7338);
nand U8954 (N_8954,N_6717,N_6059);
or U8955 (N_8955,N_7405,N_7425);
or U8956 (N_8956,N_7461,N_5982);
or U8957 (N_8957,N_5630,N_6927);
nor U8958 (N_8958,N_6088,N_6262);
xnor U8959 (N_8959,N_7235,N_7343);
or U8960 (N_8960,N_6851,N_5500);
and U8961 (N_8961,N_7257,N_5945);
nand U8962 (N_8962,N_6980,N_7424);
xor U8963 (N_8963,N_6926,N_5709);
nor U8964 (N_8964,N_6285,N_5728);
nor U8965 (N_8965,N_7293,N_5720);
and U8966 (N_8966,N_5281,N_6558);
or U8967 (N_8967,N_5554,N_6466);
nand U8968 (N_8968,N_6894,N_5473);
and U8969 (N_8969,N_6906,N_5317);
nand U8970 (N_8970,N_6875,N_6111);
or U8971 (N_8971,N_6034,N_6599);
or U8972 (N_8972,N_7037,N_5014);
xor U8973 (N_8973,N_6487,N_5005);
nand U8974 (N_8974,N_5731,N_7231);
or U8975 (N_8975,N_5433,N_5067);
and U8976 (N_8976,N_5850,N_5911);
or U8977 (N_8977,N_6265,N_7187);
xor U8978 (N_8978,N_5216,N_5053);
xor U8979 (N_8979,N_5663,N_7114);
xor U8980 (N_8980,N_6728,N_6570);
or U8981 (N_8981,N_6059,N_6445);
nor U8982 (N_8982,N_5418,N_5070);
nand U8983 (N_8983,N_5221,N_7469);
xnor U8984 (N_8984,N_7467,N_6542);
and U8985 (N_8985,N_5167,N_5691);
nor U8986 (N_8986,N_6260,N_5907);
nand U8987 (N_8987,N_5560,N_6884);
nor U8988 (N_8988,N_5103,N_6120);
nor U8989 (N_8989,N_5410,N_6563);
or U8990 (N_8990,N_7290,N_5101);
and U8991 (N_8991,N_7214,N_5581);
xnor U8992 (N_8992,N_6936,N_5293);
xor U8993 (N_8993,N_7393,N_5198);
or U8994 (N_8994,N_5792,N_6595);
nand U8995 (N_8995,N_5508,N_7209);
and U8996 (N_8996,N_7386,N_6182);
and U8997 (N_8997,N_5372,N_5787);
nor U8998 (N_8998,N_5429,N_7078);
or U8999 (N_8999,N_6931,N_7389);
or U9000 (N_9000,N_6143,N_7405);
and U9001 (N_9001,N_6229,N_6791);
nor U9002 (N_9002,N_7127,N_5814);
or U9003 (N_9003,N_6164,N_6775);
nand U9004 (N_9004,N_5902,N_6562);
and U9005 (N_9005,N_7147,N_6279);
nor U9006 (N_9006,N_6469,N_5172);
xor U9007 (N_9007,N_6169,N_5502);
and U9008 (N_9008,N_5936,N_5933);
nand U9009 (N_9009,N_5078,N_5745);
nor U9010 (N_9010,N_6299,N_5730);
and U9011 (N_9011,N_7411,N_5491);
nor U9012 (N_9012,N_5300,N_5924);
nand U9013 (N_9013,N_6696,N_5180);
nand U9014 (N_9014,N_5772,N_6328);
nor U9015 (N_9015,N_5946,N_5107);
xor U9016 (N_9016,N_7115,N_5297);
and U9017 (N_9017,N_5645,N_5618);
and U9018 (N_9018,N_5597,N_7454);
nand U9019 (N_9019,N_6743,N_6083);
nand U9020 (N_9020,N_6594,N_5134);
xnor U9021 (N_9021,N_5735,N_5932);
and U9022 (N_9022,N_7467,N_5528);
nand U9023 (N_9023,N_6806,N_5313);
nand U9024 (N_9024,N_6276,N_6046);
nor U9025 (N_9025,N_5801,N_5037);
or U9026 (N_9026,N_5521,N_6767);
xnor U9027 (N_9027,N_7288,N_5348);
xnor U9028 (N_9028,N_5324,N_7170);
and U9029 (N_9029,N_7322,N_7166);
xnor U9030 (N_9030,N_5128,N_7272);
xor U9031 (N_9031,N_6157,N_6173);
or U9032 (N_9032,N_5388,N_5268);
and U9033 (N_9033,N_5683,N_6281);
and U9034 (N_9034,N_5873,N_6133);
nor U9035 (N_9035,N_6423,N_6252);
or U9036 (N_9036,N_5896,N_7025);
nand U9037 (N_9037,N_5890,N_6631);
nor U9038 (N_9038,N_5454,N_7310);
or U9039 (N_9039,N_5179,N_5310);
nor U9040 (N_9040,N_7069,N_5565);
and U9041 (N_9041,N_7087,N_6868);
and U9042 (N_9042,N_6837,N_6234);
xnor U9043 (N_9043,N_5633,N_5009);
or U9044 (N_9044,N_6814,N_5298);
nand U9045 (N_9045,N_6238,N_7245);
xor U9046 (N_9046,N_7403,N_6873);
and U9047 (N_9047,N_5676,N_6399);
or U9048 (N_9048,N_5799,N_5713);
or U9049 (N_9049,N_5405,N_5794);
or U9050 (N_9050,N_6882,N_5465);
and U9051 (N_9051,N_5995,N_6940);
nand U9052 (N_9052,N_6300,N_7154);
nor U9053 (N_9053,N_5759,N_5536);
or U9054 (N_9054,N_6021,N_6356);
and U9055 (N_9055,N_6631,N_5153);
and U9056 (N_9056,N_5366,N_6183);
xor U9057 (N_9057,N_5407,N_6870);
nand U9058 (N_9058,N_6331,N_5213);
nand U9059 (N_9059,N_7260,N_7310);
xor U9060 (N_9060,N_7050,N_7375);
nor U9061 (N_9061,N_5640,N_5996);
nor U9062 (N_9062,N_5722,N_7075);
nand U9063 (N_9063,N_6321,N_6436);
and U9064 (N_9064,N_5669,N_5324);
and U9065 (N_9065,N_5872,N_6670);
nand U9066 (N_9066,N_6449,N_5043);
and U9067 (N_9067,N_5691,N_5015);
nand U9068 (N_9068,N_6335,N_6501);
nor U9069 (N_9069,N_7499,N_6615);
xor U9070 (N_9070,N_7397,N_6081);
nor U9071 (N_9071,N_5006,N_6142);
xor U9072 (N_9072,N_6890,N_5001);
xnor U9073 (N_9073,N_5313,N_5960);
or U9074 (N_9074,N_6994,N_6208);
and U9075 (N_9075,N_6283,N_6261);
xnor U9076 (N_9076,N_6784,N_7125);
or U9077 (N_9077,N_6030,N_5829);
nor U9078 (N_9078,N_5818,N_5383);
nor U9079 (N_9079,N_7141,N_5438);
xor U9080 (N_9080,N_5374,N_5253);
xnor U9081 (N_9081,N_5655,N_5133);
or U9082 (N_9082,N_5582,N_5354);
nor U9083 (N_9083,N_6018,N_6751);
nand U9084 (N_9084,N_6474,N_6922);
nor U9085 (N_9085,N_6587,N_6674);
and U9086 (N_9086,N_6827,N_6748);
and U9087 (N_9087,N_7063,N_5488);
nor U9088 (N_9088,N_7188,N_7097);
xnor U9089 (N_9089,N_6714,N_7423);
and U9090 (N_9090,N_6519,N_5873);
or U9091 (N_9091,N_7472,N_6057);
xnor U9092 (N_9092,N_5266,N_6049);
xnor U9093 (N_9093,N_5691,N_6962);
and U9094 (N_9094,N_5471,N_5919);
and U9095 (N_9095,N_7220,N_7050);
or U9096 (N_9096,N_6126,N_6325);
nand U9097 (N_9097,N_5009,N_5222);
nor U9098 (N_9098,N_7381,N_6551);
nor U9099 (N_9099,N_5312,N_7017);
nor U9100 (N_9100,N_6967,N_6470);
and U9101 (N_9101,N_6001,N_6300);
nand U9102 (N_9102,N_7452,N_6264);
or U9103 (N_9103,N_5460,N_5885);
xnor U9104 (N_9104,N_5108,N_6413);
nor U9105 (N_9105,N_5364,N_5967);
xnor U9106 (N_9106,N_5325,N_6069);
or U9107 (N_9107,N_6725,N_5045);
xnor U9108 (N_9108,N_6900,N_5868);
nor U9109 (N_9109,N_7296,N_5736);
nand U9110 (N_9110,N_5026,N_5903);
nor U9111 (N_9111,N_6819,N_6269);
and U9112 (N_9112,N_7403,N_5353);
xnor U9113 (N_9113,N_5834,N_5126);
nand U9114 (N_9114,N_5941,N_5783);
and U9115 (N_9115,N_7368,N_6590);
nand U9116 (N_9116,N_6204,N_7308);
nor U9117 (N_9117,N_5468,N_6640);
or U9118 (N_9118,N_5620,N_6036);
nor U9119 (N_9119,N_7113,N_5714);
and U9120 (N_9120,N_5703,N_5658);
nor U9121 (N_9121,N_6085,N_6856);
xor U9122 (N_9122,N_7415,N_6823);
nor U9123 (N_9123,N_6026,N_7253);
nor U9124 (N_9124,N_7267,N_5212);
nor U9125 (N_9125,N_7393,N_6381);
nor U9126 (N_9126,N_6301,N_7420);
and U9127 (N_9127,N_5466,N_5832);
nand U9128 (N_9128,N_6048,N_6864);
nand U9129 (N_9129,N_5530,N_5896);
and U9130 (N_9130,N_6484,N_5634);
nand U9131 (N_9131,N_6755,N_7346);
nor U9132 (N_9132,N_5623,N_5751);
and U9133 (N_9133,N_5078,N_5682);
or U9134 (N_9134,N_5497,N_5153);
and U9135 (N_9135,N_5164,N_5847);
xnor U9136 (N_9136,N_5774,N_6928);
and U9137 (N_9137,N_5971,N_6171);
and U9138 (N_9138,N_6962,N_6734);
and U9139 (N_9139,N_6630,N_6881);
xor U9140 (N_9140,N_5769,N_6647);
nand U9141 (N_9141,N_6989,N_6417);
and U9142 (N_9142,N_7132,N_7414);
and U9143 (N_9143,N_7196,N_5268);
nand U9144 (N_9144,N_7175,N_5735);
nand U9145 (N_9145,N_6131,N_7302);
nand U9146 (N_9146,N_5967,N_5174);
or U9147 (N_9147,N_6905,N_7357);
nor U9148 (N_9148,N_7295,N_5581);
or U9149 (N_9149,N_5334,N_7475);
xor U9150 (N_9150,N_7376,N_6174);
or U9151 (N_9151,N_6596,N_7107);
nand U9152 (N_9152,N_6523,N_5526);
and U9153 (N_9153,N_7376,N_5392);
xnor U9154 (N_9154,N_6145,N_6179);
and U9155 (N_9155,N_7203,N_5067);
nand U9156 (N_9156,N_7498,N_5243);
xor U9157 (N_9157,N_6132,N_6612);
and U9158 (N_9158,N_7438,N_7068);
or U9159 (N_9159,N_6954,N_5621);
nand U9160 (N_9160,N_5133,N_6267);
xnor U9161 (N_9161,N_7189,N_5440);
nor U9162 (N_9162,N_6760,N_6249);
and U9163 (N_9163,N_6453,N_6558);
nor U9164 (N_9164,N_7110,N_7335);
or U9165 (N_9165,N_5077,N_7107);
nor U9166 (N_9166,N_6727,N_6817);
nand U9167 (N_9167,N_7341,N_6029);
nand U9168 (N_9168,N_5347,N_7155);
nor U9169 (N_9169,N_5237,N_5847);
or U9170 (N_9170,N_6825,N_6625);
or U9171 (N_9171,N_5673,N_7065);
nor U9172 (N_9172,N_6805,N_7262);
xnor U9173 (N_9173,N_6296,N_5416);
and U9174 (N_9174,N_7239,N_6262);
or U9175 (N_9175,N_6228,N_5023);
xor U9176 (N_9176,N_7222,N_5964);
nor U9177 (N_9177,N_6599,N_6768);
or U9178 (N_9178,N_7006,N_5215);
and U9179 (N_9179,N_5623,N_5220);
nand U9180 (N_9180,N_5963,N_6310);
xnor U9181 (N_9181,N_5336,N_6985);
nand U9182 (N_9182,N_7415,N_7306);
xnor U9183 (N_9183,N_7185,N_5353);
nor U9184 (N_9184,N_6705,N_5244);
and U9185 (N_9185,N_6467,N_5089);
nand U9186 (N_9186,N_5419,N_5609);
xnor U9187 (N_9187,N_7003,N_6028);
nand U9188 (N_9188,N_7302,N_5677);
xnor U9189 (N_9189,N_6296,N_5840);
or U9190 (N_9190,N_5042,N_7452);
or U9191 (N_9191,N_6103,N_7443);
nor U9192 (N_9192,N_5754,N_5715);
nand U9193 (N_9193,N_5662,N_6267);
xnor U9194 (N_9194,N_6661,N_7167);
nand U9195 (N_9195,N_5660,N_5997);
or U9196 (N_9196,N_6935,N_6704);
and U9197 (N_9197,N_6505,N_5500);
and U9198 (N_9198,N_7160,N_6227);
nor U9199 (N_9199,N_7283,N_5217);
or U9200 (N_9200,N_5680,N_5102);
or U9201 (N_9201,N_5348,N_5466);
nand U9202 (N_9202,N_6407,N_7110);
nand U9203 (N_9203,N_7289,N_6818);
and U9204 (N_9204,N_6489,N_5020);
xor U9205 (N_9205,N_6780,N_5353);
xor U9206 (N_9206,N_6677,N_6766);
nand U9207 (N_9207,N_5632,N_6785);
nand U9208 (N_9208,N_5635,N_6097);
xnor U9209 (N_9209,N_5535,N_5995);
or U9210 (N_9210,N_6732,N_5027);
or U9211 (N_9211,N_5467,N_7275);
or U9212 (N_9212,N_5658,N_5223);
nor U9213 (N_9213,N_6218,N_5649);
and U9214 (N_9214,N_6647,N_6587);
nand U9215 (N_9215,N_7360,N_6325);
xor U9216 (N_9216,N_5502,N_6575);
or U9217 (N_9217,N_5502,N_5384);
or U9218 (N_9218,N_5025,N_5896);
nor U9219 (N_9219,N_5551,N_5490);
and U9220 (N_9220,N_6061,N_6154);
and U9221 (N_9221,N_5367,N_5541);
or U9222 (N_9222,N_6379,N_5318);
nor U9223 (N_9223,N_6922,N_6462);
nand U9224 (N_9224,N_5076,N_6977);
and U9225 (N_9225,N_7037,N_7103);
and U9226 (N_9226,N_6501,N_6820);
xnor U9227 (N_9227,N_7345,N_6021);
xnor U9228 (N_9228,N_6126,N_6436);
or U9229 (N_9229,N_5901,N_5402);
nor U9230 (N_9230,N_6356,N_6093);
nor U9231 (N_9231,N_7199,N_6409);
or U9232 (N_9232,N_5170,N_5342);
nand U9233 (N_9233,N_5367,N_7070);
and U9234 (N_9234,N_5286,N_6621);
xnor U9235 (N_9235,N_7343,N_5634);
nor U9236 (N_9236,N_5030,N_5578);
and U9237 (N_9237,N_6539,N_6620);
nor U9238 (N_9238,N_6033,N_5700);
nor U9239 (N_9239,N_7249,N_6454);
nand U9240 (N_9240,N_6099,N_5132);
and U9241 (N_9241,N_7356,N_6141);
nand U9242 (N_9242,N_6277,N_6893);
or U9243 (N_9243,N_6478,N_7208);
xnor U9244 (N_9244,N_7225,N_5081);
or U9245 (N_9245,N_6280,N_6254);
xnor U9246 (N_9246,N_6849,N_6790);
or U9247 (N_9247,N_7176,N_6244);
nor U9248 (N_9248,N_7037,N_6948);
xor U9249 (N_9249,N_5352,N_6322);
xnor U9250 (N_9250,N_6052,N_5040);
nor U9251 (N_9251,N_5967,N_5492);
nor U9252 (N_9252,N_6996,N_5582);
or U9253 (N_9253,N_5058,N_7180);
nand U9254 (N_9254,N_7180,N_5951);
xor U9255 (N_9255,N_5782,N_7370);
nor U9256 (N_9256,N_6264,N_5545);
xor U9257 (N_9257,N_6547,N_6649);
or U9258 (N_9258,N_5859,N_6410);
nand U9259 (N_9259,N_5850,N_5874);
nand U9260 (N_9260,N_6515,N_5441);
and U9261 (N_9261,N_7418,N_6206);
and U9262 (N_9262,N_7231,N_6302);
xnor U9263 (N_9263,N_6019,N_7010);
nand U9264 (N_9264,N_7170,N_6482);
xor U9265 (N_9265,N_6885,N_7289);
xnor U9266 (N_9266,N_6271,N_7272);
or U9267 (N_9267,N_5269,N_6420);
nor U9268 (N_9268,N_6570,N_7361);
and U9269 (N_9269,N_6419,N_6193);
and U9270 (N_9270,N_7417,N_5315);
and U9271 (N_9271,N_5608,N_5967);
nand U9272 (N_9272,N_6442,N_6870);
or U9273 (N_9273,N_6570,N_6346);
nor U9274 (N_9274,N_5029,N_6820);
nor U9275 (N_9275,N_6416,N_6318);
nor U9276 (N_9276,N_6486,N_6653);
and U9277 (N_9277,N_5008,N_5664);
xor U9278 (N_9278,N_6632,N_5217);
and U9279 (N_9279,N_5613,N_6782);
nand U9280 (N_9280,N_6879,N_6820);
xor U9281 (N_9281,N_7088,N_5546);
nor U9282 (N_9282,N_7426,N_5588);
or U9283 (N_9283,N_5667,N_5028);
and U9284 (N_9284,N_5029,N_5402);
nand U9285 (N_9285,N_5795,N_5679);
nand U9286 (N_9286,N_6949,N_6865);
and U9287 (N_9287,N_5018,N_7065);
or U9288 (N_9288,N_7310,N_5198);
and U9289 (N_9289,N_6443,N_6678);
or U9290 (N_9290,N_6619,N_6957);
and U9291 (N_9291,N_6687,N_6773);
nand U9292 (N_9292,N_6033,N_7027);
nand U9293 (N_9293,N_6186,N_7062);
nand U9294 (N_9294,N_5193,N_5189);
nor U9295 (N_9295,N_6732,N_6434);
or U9296 (N_9296,N_6794,N_5835);
xor U9297 (N_9297,N_5961,N_6435);
and U9298 (N_9298,N_5169,N_6354);
nor U9299 (N_9299,N_5803,N_6638);
and U9300 (N_9300,N_7037,N_5162);
nor U9301 (N_9301,N_5477,N_6484);
xor U9302 (N_9302,N_6689,N_5428);
or U9303 (N_9303,N_6408,N_6301);
nand U9304 (N_9304,N_5384,N_5752);
xor U9305 (N_9305,N_6350,N_6121);
xor U9306 (N_9306,N_7282,N_7128);
or U9307 (N_9307,N_7272,N_7131);
nor U9308 (N_9308,N_5190,N_6540);
nand U9309 (N_9309,N_7323,N_6801);
nand U9310 (N_9310,N_7229,N_5353);
and U9311 (N_9311,N_7307,N_7191);
and U9312 (N_9312,N_6402,N_6494);
or U9313 (N_9313,N_5444,N_7332);
or U9314 (N_9314,N_7278,N_5962);
xnor U9315 (N_9315,N_7387,N_5714);
and U9316 (N_9316,N_5144,N_6898);
nor U9317 (N_9317,N_6968,N_5393);
nor U9318 (N_9318,N_5069,N_6056);
nand U9319 (N_9319,N_6024,N_6230);
and U9320 (N_9320,N_5675,N_5929);
and U9321 (N_9321,N_6801,N_6857);
and U9322 (N_9322,N_6201,N_7485);
nand U9323 (N_9323,N_6184,N_6398);
nand U9324 (N_9324,N_5047,N_7463);
and U9325 (N_9325,N_5172,N_5798);
and U9326 (N_9326,N_5678,N_5060);
xnor U9327 (N_9327,N_5001,N_5633);
nand U9328 (N_9328,N_6843,N_6449);
nand U9329 (N_9329,N_7045,N_6159);
nor U9330 (N_9330,N_5387,N_5205);
or U9331 (N_9331,N_7235,N_5972);
and U9332 (N_9332,N_6490,N_7241);
or U9333 (N_9333,N_6844,N_7429);
and U9334 (N_9334,N_6000,N_6484);
and U9335 (N_9335,N_7002,N_6594);
xor U9336 (N_9336,N_7486,N_6020);
and U9337 (N_9337,N_7423,N_6687);
xor U9338 (N_9338,N_6012,N_7159);
xnor U9339 (N_9339,N_5487,N_6349);
and U9340 (N_9340,N_6876,N_6840);
nor U9341 (N_9341,N_6357,N_6683);
and U9342 (N_9342,N_5475,N_6402);
or U9343 (N_9343,N_5514,N_6360);
or U9344 (N_9344,N_7223,N_6042);
and U9345 (N_9345,N_5789,N_6892);
xor U9346 (N_9346,N_5263,N_6954);
and U9347 (N_9347,N_5198,N_5274);
nand U9348 (N_9348,N_7150,N_6002);
nand U9349 (N_9349,N_5922,N_5012);
nor U9350 (N_9350,N_5648,N_7020);
xor U9351 (N_9351,N_5193,N_5603);
nor U9352 (N_9352,N_6412,N_7356);
and U9353 (N_9353,N_5139,N_6089);
and U9354 (N_9354,N_6699,N_5952);
or U9355 (N_9355,N_6017,N_5269);
xor U9356 (N_9356,N_6093,N_7257);
and U9357 (N_9357,N_7102,N_5000);
nor U9358 (N_9358,N_7147,N_6679);
xnor U9359 (N_9359,N_6288,N_6895);
xnor U9360 (N_9360,N_5583,N_5240);
and U9361 (N_9361,N_6813,N_6111);
nand U9362 (N_9362,N_7118,N_6988);
nand U9363 (N_9363,N_6955,N_5184);
or U9364 (N_9364,N_7473,N_6816);
nand U9365 (N_9365,N_6236,N_6726);
and U9366 (N_9366,N_5679,N_7289);
nand U9367 (N_9367,N_7066,N_6974);
and U9368 (N_9368,N_6021,N_7237);
nor U9369 (N_9369,N_5328,N_6417);
xor U9370 (N_9370,N_6826,N_6825);
and U9371 (N_9371,N_5743,N_5068);
or U9372 (N_9372,N_7488,N_5938);
nand U9373 (N_9373,N_6260,N_6443);
xor U9374 (N_9374,N_6353,N_5021);
xnor U9375 (N_9375,N_7110,N_7387);
or U9376 (N_9376,N_7331,N_5464);
and U9377 (N_9377,N_7124,N_5378);
xnor U9378 (N_9378,N_5077,N_6658);
or U9379 (N_9379,N_6384,N_7292);
nor U9380 (N_9380,N_5096,N_7327);
xnor U9381 (N_9381,N_5960,N_6369);
xor U9382 (N_9382,N_6052,N_5592);
and U9383 (N_9383,N_6855,N_7221);
xor U9384 (N_9384,N_7312,N_6451);
xor U9385 (N_9385,N_7240,N_6947);
xnor U9386 (N_9386,N_6979,N_5907);
nor U9387 (N_9387,N_6809,N_6077);
xnor U9388 (N_9388,N_5346,N_7251);
nand U9389 (N_9389,N_7498,N_7346);
or U9390 (N_9390,N_7244,N_7324);
and U9391 (N_9391,N_7135,N_6482);
nand U9392 (N_9392,N_5784,N_6560);
nand U9393 (N_9393,N_6132,N_5719);
nor U9394 (N_9394,N_6631,N_6311);
nor U9395 (N_9395,N_7229,N_7184);
or U9396 (N_9396,N_5845,N_7401);
nand U9397 (N_9397,N_7031,N_5357);
and U9398 (N_9398,N_7172,N_6658);
nand U9399 (N_9399,N_7120,N_5748);
nor U9400 (N_9400,N_6211,N_5248);
nor U9401 (N_9401,N_5330,N_7280);
nor U9402 (N_9402,N_5946,N_6416);
or U9403 (N_9403,N_5633,N_6021);
and U9404 (N_9404,N_5561,N_5133);
nor U9405 (N_9405,N_7002,N_5318);
nor U9406 (N_9406,N_5245,N_6921);
and U9407 (N_9407,N_5739,N_7407);
nor U9408 (N_9408,N_7398,N_6331);
and U9409 (N_9409,N_6409,N_5417);
xnor U9410 (N_9410,N_6047,N_5924);
xor U9411 (N_9411,N_7392,N_5072);
and U9412 (N_9412,N_6691,N_6433);
xnor U9413 (N_9413,N_7102,N_5182);
nand U9414 (N_9414,N_6230,N_7123);
nand U9415 (N_9415,N_5209,N_6268);
or U9416 (N_9416,N_6121,N_5986);
nand U9417 (N_9417,N_5367,N_7172);
nand U9418 (N_9418,N_5677,N_5621);
or U9419 (N_9419,N_5696,N_6805);
and U9420 (N_9420,N_6576,N_6652);
and U9421 (N_9421,N_6143,N_7452);
nand U9422 (N_9422,N_6444,N_6431);
xnor U9423 (N_9423,N_5304,N_7093);
or U9424 (N_9424,N_6663,N_7042);
and U9425 (N_9425,N_7056,N_6877);
nor U9426 (N_9426,N_5725,N_5177);
xor U9427 (N_9427,N_6044,N_6772);
nor U9428 (N_9428,N_7263,N_6221);
xor U9429 (N_9429,N_7285,N_6867);
nor U9430 (N_9430,N_7000,N_6052);
and U9431 (N_9431,N_5677,N_6144);
xnor U9432 (N_9432,N_5781,N_5997);
nor U9433 (N_9433,N_5576,N_6167);
nand U9434 (N_9434,N_7404,N_6486);
nor U9435 (N_9435,N_6929,N_6183);
xor U9436 (N_9436,N_6510,N_6831);
or U9437 (N_9437,N_6807,N_7237);
or U9438 (N_9438,N_6114,N_6756);
or U9439 (N_9439,N_6910,N_6485);
nor U9440 (N_9440,N_5845,N_7448);
and U9441 (N_9441,N_6596,N_6323);
and U9442 (N_9442,N_6195,N_7167);
nand U9443 (N_9443,N_6325,N_6299);
xor U9444 (N_9444,N_5103,N_6362);
or U9445 (N_9445,N_6127,N_5889);
nand U9446 (N_9446,N_5720,N_5033);
xnor U9447 (N_9447,N_7111,N_6897);
or U9448 (N_9448,N_6709,N_6908);
xor U9449 (N_9449,N_5953,N_6089);
xnor U9450 (N_9450,N_6582,N_6075);
or U9451 (N_9451,N_5361,N_6728);
nand U9452 (N_9452,N_6193,N_5192);
nand U9453 (N_9453,N_5285,N_6945);
nor U9454 (N_9454,N_5822,N_5100);
nor U9455 (N_9455,N_7273,N_7254);
or U9456 (N_9456,N_6219,N_5958);
nand U9457 (N_9457,N_7436,N_5310);
nor U9458 (N_9458,N_7183,N_6751);
nand U9459 (N_9459,N_6672,N_6766);
and U9460 (N_9460,N_6633,N_7305);
xor U9461 (N_9461,N_6881,N_5613);
nand U9462 (N_9462,N_5390,N_6923);
nand U9463 (N_9463,N_5938,N_6129);
xor U9464 (N_9464,N_7361,N_7032);
and U9465 (N_9465,N_6394,N_6017);
and U9466 (N_9466,N_5265,N_5737);
nand U9467 (N_9467,N_5899,N_6587);
nor U9468 (N_9468,N_6486,N_6580);
nand U9469 (N_9469,N_6460,N_5593);
or U9470 (N_9470,N_6048,N_6229);
nor U9471 (N_9471,N_5502,N_7043);
xor U9472 (N_9472,N_7304,N_6523);
and U9473 (N_9473,N_7441,N_7226);
nand U9474 (N_9474,N_7146,N_6484);
nor U9475 (N_9475,N_7455,N_7288);
xor U9476 (N_9476,N_5550,N_7248);
nand U9477 (N_9477,N_6703,N_6176);
or U9478 (N_9478,N_5330,N_6757);
xor U9479 (N_9479,N_6027,N_7486);
or U9480 (N_9480,N_6508,N_5466);
xor U9481 (N_9481,N_6904,N_5520);
xor U9482 (N_9482,N_6720,N_6039);
nor U9483 (N_9483,N_5453,N_5241);
and U9484 (N_9484,N_7362,N_6986);
nor U9485 (N_9485,N_7283,N_6302);
or U9486 (N_9486,N_6692,N_7261);
xnor U9487 (N_9487,N_7037,N_5853);
nand U9488 (N_9488,N_5573,N_5422);
nor U9489 (N_9489,N_5710,N_5321);
or U9490 (N_9490,N_7064,N_7002);
or U9491 (N_9491,N_5907,N_6195);
nor U9492 (N_9492,N_6355,N_6129);
nor U9493 (N_9493,N_5880,N_7071);
nor U9494 (N_9494,N_5133,N_7429);
nor U9495 (N_9495,N_7022,N_7430);
and U9496 (N_9496,N_6320,N_7341);
or U9497 (N_9497,N_7007,N_6921);
nand U9498 (N_9498,N_6006,N_6768);
nor U9499 (N_9499,N_5329,N_5210);
nand U9500 (N_9500,N_6303,N_6926);
nand U9501 (N_9501,N_5963,N_5335);
or U9502 (N_9502,N_5411,N_6144);
nor U9503 (N_9503,N_5817,N_6607);
nand U9504 (N_9504,N_7397,N_5802);
nor U9505 (N_9505,N_6791,N_5516);
nor U9506 (N_9506,N_7347,N_6657);
xor U9507 (N_9507,N_5270,N_5550);
and U9508 (N_9508,N_6815,N_6782);
nand U9509 (N_9509,N_6896,N_5179);
nand U9510 (N_9510,N_5097,N_5493);
and U9511 (N_9511,N_5191,N_5009);
nand U9512 (N_9512,N_5956,N_7129);
xor U9513 (N_9513,N_7005,N_5388);
nand U9514 (N_9514,N_5836,N_5286);
xnor U9515 (N_9515,N_7000,N_6329);
nand U9516 (N_9516,N_6712,N_6627);
and U9517 (N_9517,N_5500,N_6792);
or U9518 (N_9518,N_7053,N_7430);
xor U9519 (N_9519,N_5393,N_7436);
nor U9520 (N_9520,N_7172,N_7282);
nor U9521 (N_9521,N_6300,N_5085);
xor U9522 (N_9522,N_6213,N_5743);
and U9523 (N_9523,N_7146,N_7235);
xor U9524 (N_9524,N_6711,N_5665);
or U9525 (N_9525,N_5166,N_6621);
xor U9526 (N_9526,N_5529,N_7468);
xnor U9527 (N_9527,N_5882,N_5332);
nor U9528 (N_9528,N_6907,N_6002);
nor U9529 (N_9529,N_5746,N_5688);
xnor U9530 (N_9530,N_5765,N_5634);
and U9531 (N_9531,N_6871,N_5138);
nand U9532 (N_9532,N_7349,N_7111);
nor U9533 (N_9533,N_7005,N_6168);
nor U9534 (N_9534,N_5033,N_7181);
and U9535 (N_9535,N_5093,N_7040);
nor U9536 (N_9536,N_7171,N_5059);
or U9537 (N_9537,N_5819,N_5366);
and U9538 (N_9538,N_6660,N_5746);
or U9539 (N_9539,N_5903,N_7481);
nor U9540 (N_9540,N_7171,N_5856);
xor U9541 (N_9541,N_5691,N_6661);
xnor U9542 (N_9542,N_6763,N_5573);
nor U9543 (N_9543,N_6455,N_5646);
nor U9544 (N_9544,N_7200,N_6225);
nand U9545 (N_9545,N_7449,N_6339);
nor U9546 (N_9546,N_7289,N_6173);
or U9547 (N_9547,N_6174,N_5411);
xnor U9548 (N_9548,N_5392,N_6642);
or U9549 (N_9549,N_6781,N_6415);
nand U9550 (N_9550,N_5379,N_5668);
nor U9551 (N_9551,N_6960,N_6963);
xnor U9552 (N_9552,N_7408,N_5746);
nand U9553 (N_9553,N_6576,N_7200);
xor U9554 (N_9554,N_7485,N_7134);
xnor U9555 (N_9555,N_6215,N_6676);
nor U9556 (N_9556,N_6322,N_5287);
nor U9557 (N_9557,N_6689,N_5072);
nor U9558 (N_9558,N_6339,N_5495);
or U9559 (N_9559,N_5815,N_5535);
or U9560 (N_9560,N_7421,N_5665);
xor U9561 (N_9561,N_5367,N_5177);
xnor U9562 (N_9562,N_7172,N_5820);
or U9563 (N_9563,N_5269,N_5324);
or U9564 (N_9564,N_6721,N_7132);
or U9565 (N_9565,N_6205,N_6800);
nand U9566 (N_9566,N_7080,N_6528);
nor U9567 (N_9567,N_7390,N_5690);
xnor U9568 (N_9568,N_5645,N_6057);
nor U9569 (N_9569,N_5672,N_5034);
nor U9570 (N_9570,N_5603,N_5305);
nand U9571 (N_9571,N_5249,N_6243);
and U9572 (N_9572,N_5433,N_6940);
and U9573 (N_9573,N_6042,N_7386);
or U9574 (N_9574,N_6786,N_6299);
and U9575 (N_9575,N_7154,N_6463);
or U9576 (N_9576,N_6815,N_5867);
nand U9577 (N_9577,N_7082,N_5875);
or U9578 (N_9578,N_6813,N_6569);
and U9579 (N_9579,N_6986,N_6086);
and U9580 (N_9580,N_5861,N_6046);
nor U9581 (N_9581,N_5292,N_6559);
or U9582 (N_9582,N_6593,N_7365);
or U9583 (N_9583,N_5056,N_6789);
or U9584 (N_9584,N_5583,N_5721);
or U9585 (N_9585,N_5889,N_6112);
nor U9586 (N_9586,N_7147,N_6868);
or U9587 (N_9587,N_7167,N_6905);
nor U9588 (N_9588,N_6491,N_6792);
or U9589 (N_9589,N_5078,N_6704);
nand U9590 (N_9590,N_6881,N_5495);
nor U9591 (N_9591,N_6697,N_6800);
and U9592 (N_9592,N_7269,N_6825);
and U9593 (N_9593,N_6892,N_6056);
and U9594 (N_9594,N_5694,N_7487);
or U9595 (N_9595,N_6134,N_5595);
xnor U9596 (N_9596,N_6617,N_7182);
or U9597 (N_9597,N_5747,N_7261);
xnor U9598 (N_9598,N_6549,N_7155);
nor U9599 (N_9599,N_5120,N_6110);
or U9600 (N_9600,N_6260,N_7398);
nor U9601 (N_9601,N_5846,N_6670);
or U9602 (N_9602,N_7104,N_6988);
nand U9603 (N_9603,N_6844,N_5190);
xor U9604 (N_9604,N_5521,N_7177);
and U9605 (N_9605,N_6171,N_6335);
or U9606 (N_9606,N_6319,N_5025);
or U9607 (N_9607,N_7452,N_6176);
nand U9608 (N_9608,N_6870,N_6641);
or U9609 (N_9609,N_6712,N_5448);
nor U9610 (N_9610,N_6892,N_5947);
xor U9611 (N_9611,N_6554,N_6735);
nand U9612 (N_9612,N_7289,N_7144);
or U9613 (N_9613,N_6703,N_6062);
nor U9614 (N_9614,N_7253,N_7343);
nor U9615 (N_9615,N_5798,N_5329);
xnor U9616 (N_9616,N_6309,N_5745);
and U9617 (N_9617,N_6023,N_7020);
nor U9618 (N_9618,N_5837,N_6328);
and U9619 (N_9619,N_7418,N_5204);
and U9620 (N_9620,N_5497,N_6265);
xor U9621 (N_9621,N_5974,N_5665);
nor U9622 (N_9622,N_5186,N_5728);
xor U9623 (N_9623,N_6613,N_6744);
and U9624 (N_9624,N_6092,N_6760);
and U9625 (N_9625,N_5915,N_7080);
nor U9626 (N_9626,N_6433,N_5290);
or U9627 (N_9627,N_5137,N_5585);
and U9628 (N_9628,N_7139,N_6300);
nor U9629 (N_9629,N_5607,N_5957);
nand U9630 (N_9630,N_6450,N_5891);
nand U9631 (N_9631,N_7313,N_5318);
xnor U9632 (N_9632,N_5028,N_5985);
and U9633 (N_9633,N_5121,N_6461);
xnor U9634 (N_9634,N_5161,N_6826);
and U9635 (N_9635,N_5919,N_6095);
and U9636 (N_9636,N_5659,N_7021);
nor U9637 (N_9637,N_5441,N_6965);
nor U9638 (N_9638,N_5581,N_6109);
nand U9639 (N_9639,N_6862,N_6905);
nor U9640 (N_9640,N_7111,N_5781);
or U9641 (N_9641,N_5551,N_6338);
xor U9642 (N_9642,N_6669,N_5935);
or U9643 (N_9643,N_7203,N_5221);
or U9644 (N_9644,N_6071,N_5602);
nor U9645 (N_9645,N_7494,N_6661);
and U9646 (N_9646,N_7251,N_6416);
and U9647 (N_9647,N_5404,N_6371);
nor U9648 (N_9648,N_6835,N_6338);
and U9649 (N_9649,N_5814,N_5332);
xnor U9650 (N_9650,N_7490,N_5434);
or U9651 (N_9651,N_6497,N_5118);
and U9652 (N_9652,N_5572,N_7251);
or U9653 (N_9653,N_5104,N_5054);
or U9654 (N_9654,N_7094,N_5553);
xnor U9655 (N_9655,N_5606,N_6207);
or U9656 (N_9656,N_7052,N_6139);
nor U9657 (N_9657,N_6757,N_6964);
nand U9658 (N_9658,N_7237,N_5014);
nand U9659 (N_9659,N_6744,N_7165);
or U9660 (N_9660,N_6024,N_6445);
or U9661 (N_9661,N_6780,N_6697);
and U9662 (N_9662,N_7184,N_6032);
or U9663 (N_9663,N_6223,N_5953);
nand U9664 (N_9664,N_5855,N_7023);
nand U9665 (N_9665,N_6098,N_6083);
or U9666 (N_9666,N_5337,N_5720);
nand U9667 (N_9667,N_5756,N_6162);
or U9668 (N_9668,N_6721,N_7419);
nand U9669 (N_9669,N_5751,N_6421);
xor U9670 (N_9670,N_5000,N_7047);
nand U9671 (N_9671,N_5643,N_5460);
nand U9672 (N_9672,N_6111,N_6794);
nand U9673 (N_9673,N_5181,N_5227);
nor U9674 (N_9674,N_6461,N_5050);
nor U9675 (N_9675,N_6045,N_5610);
nor U9676 (N_9676,N_5684,N_6536);
xnor U9677 (N_9677,N_6919,N_6923);
and U9678 (N_9678,N_5989,N_5143);
xnor U9679 (N_9679,N_5568,N_5098);
and U9680 (N_9680,N_5917,N_5496);
nor U9681 (N_9681,N_5478,N_6621);
or U9682 (N_9682,N_5705,N_6370);
xor U9683 (N_9683,N_6242,N_7138);
and U9684 (N_9684,N_5918,N_6729);
nand U9685 (N_9685,N_6614,N_7193);
nor U9686 (N_9686,N_6945,N_5142);
and U9687 (N_9687,N_7391,N_5019);
nor U9688 (N_9688,N_7012,N_5295);
nand U9689 (N_9689,N_5401,N_7372);
nor U9690 (N_9690,N_7301,N_7180);
or U9691 (N_9691,N_6342,N_5397);
and U9692 (N_9692,N_6963,N_5363);
xor U9693 (N_9693,N_6099,N_5531);
and U9694 (N_9694,N_6510,N_7473);
and U9695 (N_9695,N_6453,N_5854);
nand U9696 (N_9696,N_6485,N_7022);
and U9697 (N_9697,N_5046,N_6324);
nand U9698 (N_9698,N_7169,N_6590);
and U9699 (N_9699,N_6187,N_6684);
and U9700 (N_9700,N_5196,N_6758);
nor U9701 (N_9701,N_6924,N_5186);
xnor U9702 (N_9702,N_6937,N_7144);
nor U9703 (N_9703,N_6031,N_7138);
or U9704 (N_9704,N_5989,N_5829);
nor U9705 (N_9705,N_5345,N_6870);
nand U9706 (N_9706,N_7307,N_5248);
or U9707 (N_9707,N_7296,N_5975);
nand U9708 (N_9708,N_6490,N_5679);
or U9709 (N_9709,N_5537,N_5174);
xor U9710 (N_9710,N_5617,N_5244);
xor U9711 (N_9711,N_5932,N_5159);
nand U9712 (N_9712,N_6062,N_5648);
or U9713 (N_9713,N_5214,N_7334);
and U9714 (N_9714,N_5458,N_7239);
and U9715 (N_9715,N_5813,N_5698);
nand U9716 (N_9716,N_6011,N_6782);
or U9717 (N_9717,N_5751,N_6088);
and U9718 (N_9718,N_6160,N_6783);
and U9719 (N_9719,N_5904,N_5638);
xnor U9720 (N_9720,N_6037,N_5902);
nand U9721 (N_9721,N_7361,N_6001);
xor U9722 (N_9722,N_6290,N_6342);
nand U9723 (N_9723,N_6419,N_7341);
nand U9724 (N_9724,N_6508,N_6161);
nand U9725 (N_9725,N_5113,N_5707);
or U9726 (N_9726,N_5986,N_5734);
and U9727 (N_9727,N_7442,N_5023);
nand U9728 (N_9728,N_5079,N_7285);
and U9729 (N_9729,N_6468,N_5788);
nor U9730 (N_9730,N_6209,N_6590);
and U9731 (N_9731,N_6117,N_7327);
or U9732 (N_9732,N_6090,N_6140);
xor U9733 (N_9733,N_7380,N_5236);
and U9734 (N_9734,N_7326,N_6473);
nand U9735 (N_9735,N_5414,N_5766);
or U9736 (N_9736,N_6740,N_6818);
or U9737 (N_9737,N_6088,N_5648);
nand U9738 (N_9738,N_5075,N_5811);
nand U9739 (N_9739,N_6584,N_5986);
nand U9740 (N_9740,N_6941,N_5082);
or U9741 (N_9741,N_5450,N_5868);
nor U9742 (N_9742,N_5623,N_7084);
nor U9743 (N_9743,N_7078,N_6641);
or U9744 (N_9744,N_6564,N_6411);
xor U9745 (N_9745,N_5570,N_6925);
nand U9746 (N_9746,N_6183,N_6712);
and U9747 (N_9747,N_6202,N_5319);
nand U9748 (N_9748,N_6643,N_5826);
and U9749 (N_9749,N_5874,N_5044);
nand U9750 (N_9750,N_6964,N_6503);
and U9751 (N_9751,N_6271,N_5426);
or U9752 (N_9752,N_7498,N_6362);
xnor U9753 (N_9753,N_6422,N_7484);
or U9754 (N_9754,N_6678,N_6003);
nand U9755 (N_9755,N_6226,N_6694);
or U9756 (N_9756,N_7020,N_5180);
or U9757 (N_9757,N_7491,N_6176);
or U9758 (N_9758,N_5797,N_7151);
and U9759 (N_9759,N_5969,N_6849);
and U9760 (N_9760,N_5012,N_7076);
and U9761 (N_9761,N_7409,N_6342);
or U9762 (N_9762,N_5691,N_7183);
nand U9763 (N_9763,N_7357,N_5660);
xor U9764 (N_9764,N_5452,N_5007);
and U9765 (N_9765,N_6556,N_7403);
xor U9766 (N_9766,N_5676,N_5668);
and U9767 (N_9767,N_5911,N_5451);
nand U9768 (N_9768,N_5090,N_7388);
xor U9769 (N_9769,N_6541,N_6347);
nand U9770 (N_9770,N_7284,N_6906);
or U9771 (N_9771,N_6716,N_6912);
or U9772 (N_9772,N_6334,N_7488);
nand U9773 (N_9773,N_6029,N_6551);
nor U9774 (N_9774,N_5404,N_5504);
or U9775 (N_9775,N_5578,N_5713);
and U9776 (N_9776,N_5027,N_5324);
nand U9777 (N_9777,N_5141,N_6370);
or U9778 (N_9778,N_5271,N_6056);
xor U9779 (N_9779,N_5364,N_5561);
or U9780 (N_9780,N_5287,N_5021);
nand U9781 (N_9781,N_6712,N_5741);
and U9782 (N_9782,N_6164,N_7217);
or U9783 (N_9783,N_6824,N_5139);
or U9784 (N_9784,N_6731,N_5834);
nor U9785 (N_9785,N_7233,N_6054);
or U9786 (N_9786,N_5605,N_6624);
nand U9787 (N_9787,N_6335,N_5646);
nand U9788 (N_9788,N_5974,N_5550);
and U9789 (N_9789,N_6686,N_7465);
or U9790 (N_9790,N_7446,N_5160);
xor U9791 (N_9791,N_5437,N_5605);
and U9792 (N_9792,N_7077,N_5447);
nand U9793 (N_9793,N_6639,N_5018);
or U9794 (N_9794,N_5260,N_6255);
nor U9795 (N_9795,N_5509,N_7141);
xnor U9796 (N_9796,N_6145,N_5816);
and U9797 (N_9797,N_5763,N_7184);
and U9798 (N_9798,N_6891,N_6354);
nand U9799 (N_9799,N_7145,N_6772);
xnor U9800 (N_9800,N_6795,N_6256);
or U9801 (N_9801,N_7018,N_6914);
or U9802 (N_9802,N_5234,N_5204);
nor U9803 (N_9803,N_6330,N_6687);
or U9804 (N_9804,N_7378,N_5649);
nand U9805 (N_9805,N_7282,N_5576);
nor U9806 (N_9806,N_6136,N_5215);
xnor U9807 (N_9807,N_5747,N_5940);
nand U9808 (N_9808,N_5826,N_5344);
nor U9809 (N_9809,N_5301,N_7423);
nor U9810 (N_9810,N_5192,N_5850);
or U9811 (N_9811,N_5566,N_5875);
or U9812 (N_9812,N_5254,N_5162);
nand U9813 (N_9813,N_5902,N_6633);
nand U9814 (N_9814,N_7168,N_5973);
nor U9815 (N_9815,N_5221,N_5203);
or U9816 (N_9816,N_5513,N_5810);
xnor U9817 (N_9817,N_5931,N_5012);
and U9818 (N_9818,N_6479,N_5388);
nand U9819 (N_9819,N_5673,N_6275);
xor U9820 (N_9820,N_5655,N_7164);
nand U9821 (N_9821,N_5253,N_7223);
nand U9822 (N_9822,N_5345,N_6553);
and U9823 (N_9823,N_6219,N_7229);
xor U9824 (N_9824,N_7455,N_5461);
nor U9825 (N_9825,N_7243,N_5406);
nor U9826 (N_9826,N_5199,N_6750);
nand U9827 (N_9827,N_7122,N_5214);
xnor U9828 (N_9828,N_5341,N_5665);
and U9829 (N_9829,N_6091,N_5194);
or U9830 (N_9830,N_6961,N_7192);
xnor U9831 (N_9831,N_6710,N_7148);
nor U9832 (N_9832,N_7233,N_6975);
or U9833 (N_9833,N_7368,N_6210);
and U9834 (N_9834,N_6530,N_5870);
and U9835 (N_9835,N_5252,N_5511);
xor U9836 (N_9836,N_6718,N_6828);
nand U9837 (N_9837,N_5093,N_5590);
xor U9838 (N_9838,N_5639,N_5427);
nand U9839 (N_9839,N_6604,N_7358);
and U9840 (N_9840,N_5031,N_5979);
and U9841 (N_9841,N_5270,N_7180);
xnor U9842 (N_9842,N_6878,N_5787);
nand U9843 (N_9843,N_6905,N_6316);
nor U9844 (N_9844,N_6160,N_5358);
xnor U9845 (N_9845,N_5304,N_5290);
nand U9846 (N_9846,N_5500,N_6769);
nor U9847 (N_9847,N_5063,N_5735);
nand U9848 (N_9848,N_5445,N_5472);
xnor U9849 (N_9849,N_5503,N_5994);
xor U9850 (N_9850,N_7067,N_5747);
xor U9851 (N_9851,N_6921,N_6917);
or U9852 (N_9852,N_6429,N_5867);
xnor U9853 (N_9853,N_5326,N_7271);
nor U9854 (N_9854,N_6193,N_6045);
xor U9855 (N_9855,N_6788,N_6088);
and U9856 (N_9856,N_7332,N_5125);
nand U9857 (N_9857,N_5054,N_6485);
and U9858 (N_9858,N_6609,N_6911);
or U9859 (N_9859,N_5608,N_5233);
and U9860 (N_9860,N_5604,N_6647);
or U9861 (N_9861,N_5111,N_6842);
nand U9862 (N_9862,N_6655,N_7097);
nand U9863 (N_9863,N_6338,N_5369);
nor U9864 (N_9864,N_6174,N_6824);
nor U9865 (N_9865,N_6888,N_6671);
nand U9866 (N_9866,N_5279,N_7440);
xnor U9867 (N_9867,N_6019,N_6944);
and U9868 (N_9868,N_7143,N_5375);
nand U9869 (N_9869,N_6424,N_7155);
and U9870 (N_9870,N_5098,N_6067);
and U9871 (N_9871,N_5226,N_5677);
and U9872 (N_9872,N_7081,N_5139);
or U9873 (N_9873,N_6670,N_7128);
or U9874 (N_9874,N_5386,N_6022);
and U9875 (N_9875,N_6619,N_5721);
and U9876 (N_9876,N_6153,N_5068);
xor U9877 (N_9877,N_5192,N_5375);
and U9878 (N_9878,N_6977,N_6096);
nand U9879 (N_9879,N_6872,N_5962);
nand U9880 (N_9880,N_5728,N_5996);
and U9881 (N_9881,N_7007,N_7392);
and U9882 (N_9882,N_5010,N_6223);
nand U9883 (N_9883,N_5333,N_6134);
nor U9884 (N_9884,N_5913,N_5214);
and U9885 (N_9885,N_6867,N_7331);
nand U9886 (N_9886,N_6966,N_6851);
or U9887 (N_9887,N_7280,N_5092);
nand U9888 (N_9888,N_5681,N_5972);
or U9889 (N_9889,N_5567,N_5662);
nand U9890 (N_9890,N_6276,N_7286);
xnor U9891 (N_9891,N_6347,N_7107);
nor U9892 (N_9892,N_6843,N_5226);
and U9893 (N_9893,N_5830,N_7440);
nand U9894 (N_9894,N_5712,N_5500);
or U9895 (N_9895,N_5155,N_5747);
xor U9896 (N_9896,N_5739,N_6779);
or U9897 (N_9897,N_6164,N_5000);
and U9898 (N_9898,N_6810,N_5980);
or U9899 (N_9899,N_6986,N_7107);
or U9900 (N_9900,N_7221,N_5005);
nand U9901 (N_9901,N_6212,N_6104);
or U9902 (N_9902,N_5037,N_5432);
or U9903 (N_9903,N_6047,N_6548);
and U9904 (N_9904,N_6953,N_5768);
or U9905 (N_9905,N_6679,N_5840);
or U9906 (N_9906,N_5907,N_6903);
or U9907 (N_9907,N_5262,N_6282);
nand U9908 (N_9908,N_6819,N_6542);
xor U9909 (N_9909,N_6502,N_7483);
nand U9910 (N_9910,N_5595,N_5863);
nand U9911 (N_9911,N_7412,N_5895);
xnor U9912 (N_9912,N_7205,N_6633);
nand U9913 (N_9913,N_5509,N_5171);
nand U9914 (N_9914,N_6528,N_5715);
nor U9915 (N_9915,N_6245,N_5733);
or U9916 (N_9916,N_5281,N_7071);
nand U9917 (N_9917,N_5468,N_5802);
nand U9918 (N_9918,N_6946,N_6816);
and U9919 (N_9919,N_6609,N_7338);
or U9920 (N_9920,N_6553,N_5955);
xor U9921 (N_9921,N_5574,N_6408);
or U9922 (N_9922,N_6679,N_6233);
nand U9923 (N_9923,N_6466,N_6950);
nand U9924 (N_9924,N_5572,N_6496);
and U9925 (N_9925,N_5125,N_6161);
xnor U9926 (N_9926,N_7163,N_5026);
and U9927 (N_9927,N_6395,N_5516);
nor U9928 (N_9928,N_5101,N_6458);
or U9929 (N_9929,N_5857,N_5659);
nor U9930 (N_9930,N_5518,N_5439);
or U9931 (N_9931,N_6073,N_6132);
or U9932 (N_9932,N_7326,N_5192);
nor U9933 (N_9933,N_7337,N_5660);
or U9934 (N_9934,N_6749,N_5218);
or U9935 (N_9935,N_6865,N_7055);
and U9936 (N_9936,N_6109,N_7365);
and U9937 (N_9937,N_5355,N_5787);
xor U9938 (N_9938,N_6313,N_5571);
nand U9939 (N_9939,N_5337,N_5373);
nor U9940 (N_9940,N_5089,N_5663);
nand U9941 (N_9941,N_7167,N_7469);
xnor U9942 (N_9942,N_7347,N_7227);
nand U9943 (N_9943,N_6845,N_7035);
nand U9944 (N_9944,N_5971,N_7135);
or U9945 (N_9945,N_6881,N_7188);
xnor U9946 (N_9946,N_6205,N_6170);
xnor U9947 (N_9947,N_5665,N_7420);
or U9948 (N_9948,N_6281,N_7060);
nand U9949 (N_9949,N_5027,N_5999);
nor U9950 (N_9950,N_7039,N_7069);
nand U9951 (N_9951,N_5537,N_5009);
and U9952 (N_9952,N_5565,N_6967);
nor U9953 (N_9953,N_7258,N_5895);
and U9954 (N_9954,N_5565,N_5711);
and U9955 (N_9955,N_5449,N_7017);
and U9956 (N_9956,N_5701,N_6138);
and U9957 (N_9957,N_6942,N_5215);
nand U9958 (N_9958,N_5729,N_6379);
nand U9959 (N_9959,N_7168,N_5900);
nor U9960 (N_9960,N_5979,N_6638);
and U9961 (N_9961,N_7110,N_7149);
and U9962 (N_9962,N_5639,N_5554);
or U9963 (N_9963,N_7494,N_5095);
or U9964 (N_9964,N_5151,N_5591);
nand U9965 (N_9965,N_7240,N_6042);
and U9966 (N_9966,N_5722,N_7013);
or U9967 (N_9967,N_5776,N_7424);
xor U9968 (N_9968,N_6472,N_5193);
and U9969 (N_9969,N_6943,N_6575);
or U9970 (N_9970,N_5365,N_6362);
xnor U9971 (N_9971,N_6191,N_6057);
nor U9972 (N_9972,N_5904,N_6598);
and U9973 (N_9973,N_6695,N_6928);
xor U9974 (N_9974,N_6951,N_5403);
and U9975 (N_9975,N_6334,N_6899);
and U9976 (N_9976,N_6014,N_7435);
nand U9977 (N_9977,N_6037,N_7267);
and U9978 (N_9978,N_5948,N_6870);
or U9979 (N_9979,N_6058,N_7334);
xnor U9980 (N_9980,N_5912,N_5736);
xor U9981 (N_9981,N_6276,N_6553);
and U9982 (N_9982,N_5475,N_7419);
nor U9983 (N_9983,N_7346,N_6269);
xnor U9984 (N_9984,N_7223,N_7321);
nor U9985 (N_9985,N_7491,N_5464);
nor U9986 (N_9986,N_5085,N_6172);
or U9987 (N_9987,N_6394,N_7309);
or U9988 (N_9988,N_5433,N_6867);
xor U9989 (N_9989,N_6229,N_5085);
nand U9990 (N_9990,N_5230,N_5143);
nor U9991 (N_9991,N_7424,N_6998);
nand U9992 (N_9992,N_7021,N_6921);
and U9993 (N_9993,N_6861,N_5335);
and U9994 (N_9994,N_5406,N_6351);
nand U9995 (N_9995,N_7127,N_7194);
and U9996 (N_9996,N_6596,N_6449);
xor U9997 (N_9997,N_5742,N_5584);
nor U9998 (N_9998,N_5690,N_6638);
or U9999 (N_9999,N_5628,N_7252);
and U10000 (N_10000,N_8948,N_8205);
or U10001 (N_10001,N_9278,N_8080);
or U10002 (N_10002,N_9944,N_9609);
xnor U10003 (N_10003,N_9246,N_9764);
and U10004 (N_10004,N_9589,N_8994);
or U10005 (N_10005,N_8924,N_9530);
xor U10006 (N_10006,N_9146,N_9353);
nor U10007 (N_10007,N_7603,N_8235);
or U10008 (N_10008,N_8331,N_9389);
nor U10009 (N_10009,N_9844,N_7517);
and U10010 (N_10010,N_9721,N_9100);
nor U10011 (N_10011,N_7729,N_8553);
and U10012 (N_10012,N_9688,N_9471);
xnor U10013 (N_10013,N_8022,N_8668);
nor U10014 (N_10014,N_8090,N_9393);
or U10015 (N_10015,N_7730,N_8814);
nand U10016 (N_10016,N_8071,N_9914);
or U10017 (N_10017,N_8393,N_9260);
nor U10018 (N_10018,N_7571,N_8843);
nand U10019 (N_10019,N_8034,N_8474);
and U10020 (N_10020,N_8222,N_8544);
nand U10021 (N_10021,N_9727,N_8023);
nand U10022 (N_10022,N_8761,N_7906);
or U10023 (N_10023,N_8126,N_7907);
nand U10024 (N_10024,N_8236,N_9438);
and U10025 (N_10025,N_8536,N_9758);
xnor U10026 (N_10026,N_8621,N_9494);
or U10027 (N_10027,N_8086,N_9485);
xnor U10028 (N_10028,N_8823,N_9251);
xor U10029 (N_10029,N_7525,N_9015);
nand U10030 (N_10030,N_9941,N_8170);
or U10031 (N_10031,N_9887,N_9524);
and U10032 (N_10032,N_8674,N_9335);
xor U10033 (N_10033,N_8686,N_8442);
xor U10034 (N_10034,N_8152,N_9770);
xnor U10035 (N_10035,N_9558,N_9158);
or U10036 (N_10036,N_8917,N_9405);
xnor U10037 (N_10037,N_8586,N_9479);
and U10038 (N_10038,N_8477,N_8786);
nor U10039 (N_10039,N_8038,N_8996);
and U10040 (N_10040,N_8729,N_8505);
nor U10041 (N_10041,N_8273,N_9352);
or U10042 (N_10042,N_7608,N_9074);
xor U10043 (N_10043,N_8543,N_9965);
or U10044 (N_10044,N_8649,N_9928);
or U10045 (N_10045,N_7966,N_9790);
nor U10046 (N_10046,N_7564,N_7780);
and U10047 (N_10047,N_8787,N_9024);
and U10048 (N_10048,N_8701,N_7577);
xor U10049 (N_10049,N_9414,N_9049);
and U10050 (N_10050,N_9977,N_7929);
nand U10051 (N_10051,N_9952,N_8865);
and U10052 (N_10052,N_9326,N_9384);
xor U10053 (N_10053,N_8945,N_8276);
nor U10054 (N_10054,N_9535,N_9108);
xnor U10055 (N_10055,N_7865,N_8500);
nand U10056 (N_10056,N_8560,N_9749);
nor U10057 (N_10057,N_7764,N_7677);
or U10058 (N_10058,N_9180,N_8971);
nand U10059 (N_10059,N_8319,N_9498);
nor U10060 (N_10060,N_9464,N_9643);
nand U10061 (N_10061,N_7659,N_8252);
nand U10062 (N_10062,N_8730,N_8137);
nand U10063 (N_10063,N_7829,N_8770);
nand U10064 (N_10064,N_8635,N_8282);
nor U10065 (N_10065,N_7628,N_9674);
or U10066 (N_10066,N_9800,N_8470);
nand U10067 (N_10067,N_7832,N_8144);
nand U10068 (N_10068,N_9953,N_8092);
nand U10069 (N_10069,N_7768,N_7546);
and U10070 (N_10070,N_9431,N_8749);
and U10071 (N_10071,N_7711,N_8731);
nand U10072 (N_10072,N_9646,N_9083);
nand U10073 (N_10073,N_7982,N_9968);
nand U10074 (N_10074,N_8661,N_8979);
or U10075 (N_10075,N_7957,N_8293);
xor U10076 (N_10076,N_9415,N_8651);
or U10077 (N_10077,N_8483,N_8875);
nand U10078 (N_10078,N_8400,N_8970);
and U10079 (N_10079,N_9657,N_8502);
xnor U10080 (N_10080,N_8708,N_8617);
and U10081 (N_10081,N_8690,N_9433);
and U10082 (N_10082,N_8744,N_9480);
nor U10083 (N_10083,N_9368,N_7878);
xor U10084 (N_10084,N_8292,N_8112);
nor U10085 (N_10085,N_8892,N_8440);
and U10086 (N_10086,N_8081,N_8489);
xor U10087 (N_10087,N_7720,N_9231);
xor U10088 (N_10088,N_7936,N_7520);
xnor U10089 (N_10089,N_9877,N_7568);
and U10090 (N_10090,N_8135,N_7699);
or U10091 (N_10091,N_8327,N_8532);
xor U10092 (N_10092,N_8431,N_8695);
and U10093 (N_10093,N_8463,N_9762);
and U10094 (N_10094,N_8334,N_9677);
nor U10095 (N_10095,N_8065,N_8703);
and U10096 (N_10096,N_9942,N_7856);
and U10097 (N_10097,N_7594,N_8527);
xor U10098 (N_10098,N_7626,N_8568);
nor U10099 (N_10099,N_7841,N_8029);
and U10100 (N_10100,N_8433,N_8889);
or U10101 (N_10101,N_7978,N_9228);
xnor U10102 (N_10102,N_8115,N_7912);
xnor U10103 (N_10103,N_8202,N_9280);
xor U10104 (N_10104,N_9726,N_9717);
and U10105 (N_10105,N_7821,N_8177);
and U10106 (N_10106,N_8461,N_7536);
or U10107 (N_10107,N_7728,N_9362);
nor U10108 (N_10108,N_8420,N_7977);
and U10109 (N_10109,N_9686,N_8099);
nor U10110 (N_10110,N_7523,N_7782);
and U10111 (N_10111,N_8827,N_8138);
or U10112 (N_10112,N_8852,N_9711);
or U10113 (N_10113,N_8526,N_8165);
xnor U10114 (N_10114,N_7937,N_7923);
xnor U10115 (N_10115,N_9363,N_9864);
or U10116 (N_10116,N_9318,N_9680);
or U10117 (N_10117,N_7621,N_8339);
nor U10118 (N_10118,N_8764,N_9071);
nand U10119 (N_10119,N_8569,N_7875);
and U10120 (N_10120,N_8938,N_8345);
nand U10121 (N_10121,N_8687,N_8610);
or U10122 (N_10122,N_8278,N_8328);
xnor U10123 (N_10123,N_9969,N_9302);
or U10124 (N_10124,N_9059,N_8123);
and U10125 (N_10125,N_8002,N_9736);
nor U10126 (N_10126,N_7514,N_9150);
nor U10127 (N_10127,N_8662,N_8231);
and U10128 (N_10128,N_7548,N_9279);
or U10129 (N_10129,N_8998,N_7814);
and U10130 (N_10130,N_8528,N_8401);
and U10131 (N_10131,N_8897,N_8000);
nand U10132 (N_10132,N_8910,N_9684);
nor U10133 (N_10133,N_9513,N_8270);
or U10134 (N_10134,N_8632,N_7647);
xnor U10135 (N_10135,N_8828,N_7712);
nor U10136 (N_10136,N_7547,N_7749);
nor U10137 (N_10137,N_8845,N_9351);
nor U10138 (N_10138,N_8743,N_8702);
xnor U10139 (N_10139,N_9011,N_7954);
nand U10140 (N_10140,N_8604,N_9295);
nor U10141 (N_10141,N_8941,N_9579);
nand U10142 (N_10142,N_7706,N_9852);
nand U10143 (N_10143,N_9564,N_7917);
or U10144 (N_10144,N_8061,N_8168);
xor U10145 (N_10145,N_9000,N_9078);
nor U10146 (N_10146,N_9585,N_8098);
and U10147 (N_10147,N_7855,N_8836);
or U10148 (N_10148,N_9984,N_9805);
and U10149 (N_10149,N_9731,N_9903);
xnor U10150 (N_10150,N_9744,N_8896);
or U10151 (N_10151,N_9293,N_7962);
xor U10152 (N_10152,N_7817,N_8959);
or U10153 (N_10153,N_9491,N_8009);
or U10154 (N_10154,N_9202,N_8798);
xor U10155 (N_10155,N_9938,N_7785);
xnor U10156 (N_10156,N_8773,N_8486);
xnor U10157 (N_10157,N_8010,N_8296);
or U10158 (N_10158,N_7839,N_8001);
nor U10159 (N_10159,N_7807,N_8371);
xor U10160 (N_10160,N_8559,N_7838);
and U10161 (N_10161,N_7922,N_9216);
or U10162 (N_10162,N_9300,N_9858);
or U10163 (N_10163,N_9014,N_8975);
nor U10164 (N_10164,N_9148,N_9305);
and U10165 (N_10165,N_7913,N_8193);
nand U10166 (N_10166,N_9840,N_8448);
and U10167 (N_10167,N_9937,N_8429);
or U10168 (N_10168,N_9662,N_8057);
nand U10169 (N_10169,N_8771,N_9945);
or U10170 (N_10170,N_9257,N_9547);
nor U10171 (N_10171,N_8343,N_9332);
nor U10172 (N_10172,N_8699,N_7702);
xor U10173 (N_10173,N_9409,N_9529);
nand U10174 (N_10174,N_9194,N_8395);
and U10175 (N_10175,N_7911,N_7823);
nand U10176 (N_10176,N_9271,N_9741);
xnor U10177 (N_10177,N_7794,N_7971);
nand U10178 (N_10178,N_9036,N_8886);
nand U10179 (N_10179,N_8653,N_9930);
nand U10180 (N_10180,N_7770,N_9815);
xnor U10181 (N_10181,N_8375,N_7803);
nand U10182 (N_10182,N_7819,N_9436);
and U10183 (N_10183,N_9678,N_8487);
or U10184 (N_10184,N_8735,N_9812);
or U10185 (N_10185,N_8931,N_8390);
or U10186 (N_10186,N_9706,N_9843);
nand U10187 (N_10187,N_9665,N_9365);
xnor U10188 (N_10188,N_7662,N_8871);
nand U10189 (N_10189,N_8266,N_9313);
xnor U10190 (N_10190,N_9113,N_8605);
nor U10191 (N_10191,N_8321,N_9974);
and U10192 (N_10192,N_8341,N_9110);
or U10193 (N_10193,N_8417,N_9331);
and U10194 (N_10194,N_8885,N_9661);
xor U10195 (N_10195,N_7612,N_9361);
xor U10196 (N_10196,N_9488,N_8707);
nand U10197 (N_10197,N_7715,N_7869);
or U10198 (N_10198,N_8513,N_9077);
or U10199 (N_10199,N_9356,N_7793);
nand U10200 (N_10200,N_9510,N_9693);
and U10201 (N_10201,N_7554,N_8881);
nor U10202 (N_10202,N_8418,N_9329);
and U10203 (N_10203,N_9209,N_7560);
or U10204 (N_10204,N_8226,N_8696);
or U10205 (N_10205,N_8724,N_8893);
nor U10206 (N_10206,N_8146,N_9334);
xnor U10207 (N_10207,N_8655,N_8493);
xor U10208 (N_10208,N_9294,N_8337);
or U10209 (N_10209,N_8563,N_8154);
nor U10210 (N_10210,N_8589,N_9196);
or U10211 (N_10211,N_7501,N_8746);
nor U10212 (N_10212,N_9070,N_7524);
or U10213 (N_10213,N_9712,N_9648);
or U10214 (N_10214,N_8063,N_9574);
nand U10215 (N_10215,N_8973,N_7505);
and U10216 (N_10216,N_9020,N_8025);
xnor U10217 (N_10217,N_9575,N_8925);
nor U10218 (N_10218,N_8723,N_9446);
nor U10219 (N_10219,N_8866,N_8013);
nand U10220 (N_10220,N_7944,N_8113);
and U10221 (N_10221,N_8873,N_9526);
nand U10222 (N_10222,N_7624,N_9270);
and U10223 (N_10223,N_7646,N_9669);
or U10224 (N_10224,N_8272,N_8834);
or U10225 (N_10225,N_9618,N_8336);
nor U10226 (N_10226,N_8241,N_7802);
and U10227 (N_10227,N_9065,N_9986);
nand U10228 (N_10228,N_8076,N_7800);
nand U10229 (N_10229,N_8534,N_9062);
or U10230 (N_10230,N_7736,N_7748);
and U10231 (N_10231,N_8955,N_9003);
nor U10232 (N_10232,N_8715,N_8406);
and U10233 (N_10233,N_9109,N_8101);
xnor U10234 (N_10234,N_8134,N_8084);
and U10235 (N_10235,N_9336,N_8303);
or U10236 (N_10236,N_9555,N_8085);
xnor U10237 (N_10237,N_9568,N_9154);
nor U10238 (N_10238,N_8880,N_9076);
and U10239 (N_10239,N_9732,N_8988);
xnor U10240 (N_10240,N_9068,N_9738);
or U10241 (N_10241,N_9502,N_9814);
nor U10242 (N_10242,N_9989,N_9675);
xor U10243 (N_10243,N_8891,N_9307);
nor U10244 (N_10244,N_9848,N_9652);
nand U10245 (N_10245,N_9052,N_9705);
nand U10246 (N_10246,N_8516,N_9651);
nand U10247 (N_10247,N_9879,N_9614);
nand U10248 (N_10248,N_7527,N_8452);
and U10249 (N_10249,N_9090,N_9911);
xor U10250 (N_10250,N_8570,N_9483);
xnor U10251 (N_10251,N_7602,N_8215);
or U10252 (N_10252,N_8999,N_7726);
nand U10253 (N_10253,N_9772,N_8802);
nor U10254 (N_10254,N_7503,N_7587);
or U10255 (N_10255,N_8186,N_8658);
or U10256 (N_10256,N_9452,N_8369);
nand U10257 (N_10257,N_9343,N_8848);
nand U10258 (N_10258,N_8275,N_7894);
or U10259 (N_10259,N_8567,N_9632);
and U10260 (N_10260,N_8811,N_7790);
nand U10261 (N_10261,N_9262,N_8953);
xnor U10262 (N_10262,N_9364,N_7660);
nor U10263 (N_10263,N_9878,N_9459);
nand U10264 (N_10264,N_9566,N_9897);
and U10265 (N_10265,N_9601,N_8054);
xnor U10266 (N_10266,N_7857,N_8330);
nand U10267 (N_10267,N_8481,N_9640);
nor U10268 (N_10268,N_8779,N_9139);
xnor U10269 (N_10269,N_9865,N_8810);
or U10270 (N_10270,N_9901,N_9277);
and U10271 (N_10271,N_7617,N_8911);
nand U10272 (N_10272,N_9037,N_9048);
nor U10273 (N_10273,N_9315,N_7678);
and U10274 (N_10274,N_9201,N_9173);
or U10275 (N_10275,N_7949,N_9046);
xor U10276 (N_10276,N_9704,N_8874);
xnor U10277 (N_10277,N_7630,N_8310);
and U10278 (N_10278,N_8130,N_9411);
and U10279 (N_10279,N_9912,N_9458);
nand U10280 (N_10280,N_7590,N_8797);
nor U10281 (N_10281,N_9298,N_8815);
or U10282 (N_10282,N_7529,N_8585);
xnor U10283 (N_10283,N_8370,N_9245);
and U10284 (N_10284,N_7787,N_8741);
and U10285 (N_10285,N_7778,N_7583);
nor U10286 (N_10286,N_8851,N_9230);
nand U10287 (N_10287,N_9427,N_8736);
nand U10288 (N_10288,N_7902,N_8195);
nand U10289 (N_10289,N_8041,N_7579);
nand U10290 (N_10290,N_8638,N_8171);
nor U10291 (N_10291,N_8323,N_9666);
and U10292 (N_10292,N_9016,N_9366);
and U10293 (N_10293,N_8571,N_9539);
or U10294 (N_10294,N_7994,N_9103);
and U10295 (N_10295,N_9545,N_9715);
xor U10296 (N_10296,N_8795,N_9337);
and U10297 (N_10297,N_9631,N_8082);
nand U10298 (N_10298,N_9837,N_8407);
xnor U10299 (N_10299,N_8857,N_8684);
and U10300 (N_10300,N_9592,N_8471);
nand U10301 (N_10301,N_9017,N_9779);
xnor U10302 (N_10302,N_7920,N_8385);
nor U10303 (N_10303,N_9166,N_7507);
or U10304 (N_10304,N_8713,N_9185);
nand U10305 (N_10305,N_7989,N_9916);
and U10306 (N_10306,N_9634,N_9587);
xor U10307 (N_10307,N_8618,N_9450);
nand U10308 (N_10308,N_9101,N_8158);
nand U10309 (N_10309,N_8650,N_9080);
xor U10310 (N_10310,N_7940,N_8204);
and U10311 (N_10311,N_7837,N_8225);
xnor U10312 (N_10312,N_8541,N_9475);
and U10313 (N_10313,N_9689,N_9890);
nor U10314 (N_10314,N_9296,N_8249);
or U10315 (N_10315,N_9988,N_8383);
nor U10316 (N_10316,N_9636,N_7588);
or U10317 (N_10317,N_7613,N_8382);
xnor U10318 (N_10318,N_8556,N_9243);
nand U10319 (N_10319,N_9321,N_9456);
or U10320 (N_10320,N_9473,N_7506);
and U10321 (N_10321,N_8676,N_9598);
nand U10322 (N_10322,N_7988,N_9042);
or U10323 (N_10323,N_9633,N_9025);
or U10324 (N_10324,N_7811,N_9033);
nor U10325 (N_10325,N_7885,N_9700);
and U10326 (N_10326,N_8344,N_7597);
nor U10327 (N_10327,N_9818,N_8169);
nor U10328 (N_10328,N_8199,N_9591);
nor U10329 (N_10329,N_9383,N_8265);
and U10330 (N_10330,N_9121,N_7804);
or U10331 (N_10331,N_7903,N_8129);
nor U10332 (N_10332,N_7767,N_9792);
nand U10333 (N_10333,N_9047,N_9492);
xnor U10334 (N_10334,N_7708,N_8167);
or U10335 (N_10335,N_7866,N_7570);
nand U10336 (N_10336,N_8213,N_9917);
or U10337 (N_10337,N_8394,N_7721);
and U10338 (N_10338,N_7609,N_9191);
nor U10339 (N_10339,N_8698,N_7710);
nand U10340 (N_10340,N_9947,N_9908);
nand U10341 (N_10341,N_7655,N_9940);
or U10342 (N_10342,N_9511,N_9958);
nor U10343 (N_10343,N_8105,N_9949);
or U10344 (N_10344,N_8884,N_7561);
nor U10345 (N_10345,N_9217,N_9733);
nor U10346 (N_10346,N_8627,N_7806);
or U10347 (N_10347,N_8190,N_8763);
nor U10348 (N_10348,N_9451,N_9860);
or U10349 (N_10349,N_7834,N_8781);
or U10350 (N_10350,N_8117,N_7663);
or U10351 (N_10351,N_8709,N_8623);
nand U10352 (N_10352,N_8238,N_8829);
nor U10353 (N_10353,N_8333,N_9576);
xnor U10354 (N_10354,N_8943,N_9345);
xnor U10355 (N_10355,N_8007,N_9543);
and U10356 (N_10356,N_8841,N_9416);
nand U10357 (N_10357,N_9716,N_8789);
nor U10358 (N_10358,N_8596,N_8194);
nor U10359 (N_10359,N_9743,N_8965);
or U10360 (N_10360,N_9328,N_7636);
xnor U10361 (N_10361,N_7997,N_8597);
nand U10362 (N_10362,N_7705,N_9820);
and U10363 (N_10363,N_9553,N_8940);
and U10364 (N_10364,N_8475,N_9975);
xnor U10365 (N_10365,N_8855,N_7718);
or U10366 (N_10366,N_9478,N_8267);
nor U10367 (N_10367,N_8986,N_9647);
nor U10368 (N_10368,N_8446,N_9596);
and U10369 (N_10369,N_9541,N_7851);
nand U10370 (N_10370,N_9454,N_8643);
nand U10371 (N_10371,N_8868,N_7614);
nor U10372 (N_10372,N_9867,N_7759);
or U10373 (N_10373,N_8870,N_9099);
and U10374 (N_10374,N_8928,N_9115);
xor U10375 (N_10375,N_9259,N_9323);
xor U10376 (N_10376,N_8290,N_8445);
xnor U10377 (N_10377,N_8862,N_9723);
nor U10378 (N_10378,N_8381,N_8473);
or U10379 (N_10379,N_7969,N_8291);
nor U10380 (N_10380,N_8012,N_8972);
and U10381 (N_10381,N_8737,N_8289);
or U10382 (N_10382,N_8148,N_8042);
and U10383 (N_10383,N_7606,N_8324);
or U10384 (N_10384,N_9578,N_7955);
and U10385 (N_10385,N_9709,N_9525);
nand U10386 (N_10386,N_9420,N_9249);
or U10387 (N_10387,N_8530,N_9274);
and U10388 (N_10388,N_9029,N_9835);
xnor U10389 (N_10389,N_9831,N_8478);
or U10390 (N_10390,N_8982,N_7953);
nand U10391 (N_10391,N_9909,N_7665);
nor U10392 (N_10392,N_9748,N_7863);
and U10393 (N_10393,N_9187,N_9287);
nand U10394 (N_10394,N_9006,N_8537);
nor U10395 (N_10395,N_7552,N_7716);
and U10396 (N_10396,N_9970,N_9240);
nand U10397 (N_10397,N_8738,N_7550);
or U10398 (N_10398,N_9221,N_8325);
nor U10399 (N_10399,N_7941,N_9497);
xnor U10400 (N_10400,N_8279,N_9058);
nand U10401 (N_10401,N_9425,N_9111);
nand U10402 (N_10402,N_9250,N_7596);
and U10403 (N_10403,N_8642,N_8540);
xor U10404 (N_10404,N_7826,N_8326);
or U10405 (N_10405,N_8125,N_9886);
or U10406 (N_10406,N_9181,N_9387);
or U10407 (N_10407,N_7629,N_9208);
nand U10408 (N_10408,N_7927,N_9489);
xor U10409 (N_10409,N_8479,N_8246);
nor U10410 (N_10410,N_8318,N_7796);
and U10411 (N_10411,N_9728,N_8660);
or U10412 (N_10412,N_8392,N_9819);
and U10413 (N_10413,N_7774,N_9962);
xor U10414 (N_10414,N_8286,N_8645);
and U10415 (N_10415,N_8335,N_8634);
xnor U10416 (N_10416,N_8987,N_9169);
or U10417 (N_10417,N_8163,N_9496);
nand U10418 (N_10418,N_9019,N_9195);
or U10419 (N_10419,N_8077,N_7801);
nand U10420 (N_10420,N_9872,N_7859);
nand U10421 (N_10421,N_9045,N_8912);
nand U10422 (N_10422,N_9135,N_8021);
or U10423 (N_10423,N_9399,N_8058);
nand U10424 (N_10424,N_8221,N_8357);
or U10425 (N_10425,N_7893,N_9851);
nand U10426 (N_10426,N_8185,N_8459);
nor U10427 (N_10427,N_8800,N_8759);
nand U10428 (N_10428,N_8320,N_8372);
or U10429 (N_10429,N_8268,N_9849);
nand U10430 (N_10430,N_8842,N_9784);
and U10431 (N_10431,N_7610,N_9934);
xor U10432 (N_10432,N_9972,N_8903);
nand U10433 (N_10433,N_7639,N_9931);
nor U10434 (N_10434,N_7576,N_9403);
or U10435 (N_10435,N_9992,N_9691);
xor U10436 (N_10436,N_8430,N_8712);
nor U10437 (N_10437,N_7792,N_9960);
nor U10438 (N_10438,N_9876,N_7669);
xor U10439 (N_10439,N_7752,N_8719);
nand U10440 (N_10440,N_9220,N_9341);
and U10441 (N_10441,N_9429,N_9737);
nand U10442 (N_10442,N_8514,N_7535);
or U10443 (N_10443,N_9263,N_9299);
nand U10444 (N_10444,N_9594,N_7641);
and U10445 (N_10445,N_9692,N_8710);
and U10446 (N_10446,N_9548,N_9767);
xnor U10447 (N_10447,N_7586,N_8142);
or U10448 (N_10448,N_7582,N_8095);
xnor U10449 (N_10449,N_8316,N_8366);
and U10450 (N_10450,N_9314,N_7513);
nor U10451 (N_10451,N_9789,N_9798);
xor U10452 (N_10452,N_9994,N_8412);
xnor U10453 (N_10453,N_7788,N_7771);
xnor U10454 (N_10454,N_9707,N_8485);
and U10455 (N_10455,N_9829,N_8102);
xor U10456 (N_10456,N_8051,N_8898);
or U10457 (N_10457,N_9040,N_8969);
and U10458 (N_10458,N_8991,N_8673);
nor U10459 (N_10459,N_7541,N_9455);
and U10460 (N_10460,N_9979,N_9740);
nand U10461 (N_10461,N_8467,N_8380);
xnor U10462 (N_10462,N_8636,N_8469);
or U10463 (N_10463,N_8352,N_9826);
xor U10464 (N_10464,N_9856,N_7958);
nor U10465 (N_10465,N_9859,N_8878);
nor U10466 (N_10466,N_9222,N_8260);
and U10467 (N_10467,N_9339,N_8353);
nand U10468 (N_10468,N_9556,N_9204);
or U10469 (N_10469,N_8219,N_7942);
xnor U10470 (N_10470,N_9239,N_8128);
or U10471 (N_10471,N_7762,N_9127);
or U10472 (N_10472,N_7575,N_8601);
xor U10473 (N_10473,N_8824,N_8229);
nor U10474 (N_10474,N_9681,N_9788);
nor U10475 (N_10475,N_9520,N_7965);
nand U10476 (N_10476,N_8685,N_8804);
or U10477 (N_10477,N_8515,N_9285);
and U10478 (N_10478,N_8411,N_7661);
or U10479 (N_10479,N_9563,N_8234);
or U10480 (N_10480,N_8754,N_9390);
nor U10481 (N_10481,N_8872,N_9701);
nor U10482 (N_10482,N_8579,N_9760);
or U10483 (N_10483,N_9129,N_9774);
nor U10484 (N_10484,N_8512,N_9896);
nor U10485 (N_10485,N_8564,N_7504);
nor U10486 (N_10486,N_8960,N_9995);
nand U10487 (N_10487,N_7963,N_9237);
nor U10488 (N_10488,N_9276,N_9883);
nor U10489 (N_10489,N_8173,N_9752);
xnor U10490 (N_10490,N_8631,N_8933);
xor U10491 (N_10491,N_7673,N_9234);
nand U10492 (N_10492,N_8174,N_8611);
and U10493 (N_10493,N_8410,N_8131);
and U10494 (N_10494,N_7670,N_7551);
and U10495 (N_10495,N_8616,N_8523);
or U10496 (N_10496,N_9847,N_8727);
and U10497 (N_10497,N_7599,N_9854);
and U10498 (N_10498,N_7836,N_7620);
nor U10499 (N_10499,N_9540,N_8792);
or U10500 (N_10500,N_9206,N_8518);
nand U10501 (N_10501,N_9742,N_9342);
or U10502 (N_10502,N_9874,N_9667);
or U10503 (N_10503,N_7891,N_8950);
nand U10504 (N_10504,N_8049,N_8967);
xnor U10505 (N_10505,N_9075,N_9283);
xnor U10506 (N_10506,N_7512,N_9768);
nand U10507 (N_10507,N_9963,N_7627);
nand U10508 (N_10508,N_8091,N_9394);
nor U10509 (N_10509,N_8808,N_7760);
or U10510 (N_10510,N_9765,N_9913);
nor U10511 (N_10511,N_8706,N_9573);
nand U10512 (N_10512,N_9385,N_7725);
xor U10513 (N_10513,N_8398,N_9515);
and U10514 (N_10514,N_9224,N_8208);
nand U10515 (N_10515,N_7980,N_8191);
nor U10516 (N_10516,N_8269,N_8005);
xnor U10517 (N_10517,N_9032,N_9229);
nand U10518 (N_10518,N_9645,N_9521);
nor U10519 (N_10519,N_7697,N_9503);
xnor U10520 (N_10520,N_8581,N_8908);
nand U10521 (N_10521,N_9660,N_8338);
or U10522 (N_10522,N_8498,N_9162);
xnor U10523 (N_10523,N_9730,N_9939);
nor U10524 (N_10524,N_9920,N_9924);
and U10525 (N_10525,N_9655,N_8716);
nand U10526 (N_10526,N_7723,N_9442);
or U10527 (N_10527,N_9170,N_9401);
nor U10528 (N_10528,N_9735,N_9120);
xnor U10529 (N_10529,N_8424,N_8722);
nand U10530 (N_10530,N_7680,N_7815);
xnor U10531 (N_10531,N_7905,N_7968);
or U10532 (N_10532,N_9561,N_7964);
and U10533 (N_10533,N_7543,N_9990);
and U10534 (N_10534,N_7611,N_7926);
or U10535 (N_10535,N_8239,N_9532);
xnor U10536 (N_10536,N_8583,N_8035);
nor U10537 (N_10537,N_8801,N_9757);
nor U10538 (N_10538,N_9584,N_9468);
nand U10539 (N_10539,N_9833,N_9621);
or U10540 (N_10540,N_9641,N_9799);
xor U10541 (N_10541,N_9428,N_8700);
nand U10542 (N_10542,N_9720,N_8166);
xnor U10543 (N_10543,N_7717,N_9215);
nor U10544 (N_10544,N_8263,N_8853);
nand U10545 (N_10545,N_8952,N_7648);
xor U10546 (N_10546,N_9569,N_8900);
and U10547 (N_10547,N_7516,N_9906);
and U10548 (N_10548,N_9842,N_8096);
nor U10549 (N_10549,N_8060,N_8745);
or U10550 (N_10550,N_7742,N_7895);
nand U10551 (N_10551,N_8214,N_7945);
xor U10552 (N_10552,N_7578,N_8155);
or U10553 (N_10553,N_9355,N_9499);
or U10554 (N_10554,N_9183,N_9060);
or U10555 (N_10555,N_7990,N_8805);
or U10556 (N_10556,N_9378,N_7709);
and U10557 (N_10557,N_7886,N_8927);
xor U10558 (N_10558,N_8351,N_8046);
nand U10559 (N_10559,N_8663,N_8378);
nor U10560 (N_10560,N_8584,N_9806);
nand U10561 (N_10561,N_9813,N_8577);
xor U10562 (N_10562,N_8230,N_7518);
nand U10563 (N_10563,N_8149,N_8426);
nor U10564 (N_10564,N_8162,N_8666);
nand U10565 (N_10565,N_9694,N_8124);
nor U10566 (N_10566,N_7645,N_9775);
or U10567 (N_10567,N_9698,N_9374);
nand U10568 (N_10568,N_9501,N_8044);
nor U10569 (N_10569,N_8451,N_9344);
nand U10570 (N_10570,N_7996,N_9238);
and U10571 (N_10571,N_8434,N_7592);
or U10572 (N_10572,N_8739,N_9863);
nand U10573 (N_10573,N_8108,N_8078);
or U10574 (N_10574,N_8587,N_9102);
and U10575 (N_10575,N_8818,N_9649);
nor U10576 (N_10576,N_9447,N_9616);
xnor U10577 (N_10577,N_9082,N_8386);
or U10578 (N_10578,N_7510,N_8854);
nand U10579 (N_10579,N_7864,N_9093);
and U10580 (N_10580,N_9626,N_7656);
nand U10581 (N_10581,N_9236,N_8100);
nand U10582 (N_10582,N_8694,N_9957);
xor U10583 (N_10583,N_7756,N_9097);
xor U10584 (N_10584,N_9670,N_8681);
and U10585 (N_10585,N_7714,N_8966);
nand U10586 (N_10586,N_9210,N_9190);
nand U10587 (N_10587,N_9004,N_8796);
nor U10588 (N_10588,N_9954,N_9461);
or U10589 (N_10589,N_9839,N_9892);
and U10590 (N_10590,N_8550,N_8914);
nor U10591 (N_10591,N_9255,N_8311);
and U10592 (N_10592,N_7999,N_8990);
xnor U10593 (N_10593,N_9918,N_7534);
and U10594 (N_10594,N_8097,N_9248);
xor U10595 (N_10595,N_9266,N_9193);
or U10596 (N_10596,N_9611,N_7738);
nand U10597 (N_10597,N_9088,N_8551);
nand U10598 (N_10598,N_9932,N_9889);
and U10599 (N_10599,N_8281,N_9756);
xnor U10600 (N_10600,N_8329,N_9550);
xnor U10601 (N_10601,N_8180,N_9282);
xnor U10602 (N_10602,N_7727,N_8895);
and U10603 (N_10603,N_7668,N_8626);
and U10604 (N_10604,N_8422,N_8522);
nand U10605 (N_10605,N_7675,N_7634);
nand U10606 (N_10606,N_8074,N_9659);
nor U10607 (N_10607,N_9888,N_8340);
and U10608 (N_10608,N_8062,N_8482);
nand U10609 (N_10609,N_7930,N_7544);
or U10610 (N_10610,N_9725,N_7998);
and U10611 (N_10611,N_9448,N_8641);
or U10612 (N_10612,N_8262,N_7810);
nand U10613 (N_10613,N_8508,N_9227);
nand U10614 (N_10614,N_8939,N_7625);
nand U10615 (N_10615,N_9105,N_7844);
or U10616 (N_10616,N_8346,N_8159);
xor U10617 (N_10617,N_9933,N_7731);
and U10618 (N_10618,N_7858,N_9096);
and U10619 (N_10619,N_8612,N_7690);
nor U10620 (N_10620,N_8887,N_9367);
and U10621 (N_10621,N_7862,N_8409);
nor U10622 (N_10622,N_9570,N_9581);
nand U10623 (N_10623,N_9582,N_8143);
xnor U10624 (N_10624,N_7827,N_9147);
nor U10625 (N_10625,N_9226,N_7753);
or U10626 (N_10626,N_9466,N_7537);
xnor U10627 (N_10627,N_8529,N_9797);
nand U10628 (N_10628,N_8421,N_8283);
xnor U10629 (N_10629,N_7696,N_9376);
xor U10630 (N_10630,N_8785,N_8361);
and U10631 (N_10631,N_9369,N_9136);
nor U10632 (N_10632,N_9832,N_8639);
and U10633 (N_10633,N_8628,N_8954);
or U10634 (N_10634,N_7981,N_9755);
xnor U10635 (N_10635,N_8360,N_8902);
nor U10636 (N_10636,N_7882,N_8457);
and U10637 (N_10637,N_9623,N_7861);
and U10638 (N_10638,N_8192,N_8243);
or U10639 (N_10639,N_9590,N_7595);
xor U10640 (N_10640,N_8506,N_9043);
or U10641 (N_10641,N_9031,N_8602);
or U10642 (N_10642,N_9177,N_8748);
or U10643 (N_10643,N_9165,N_9845);
nand U10644 (N_10644,N_8858,N_8995);
nand U10645 (N_10645,N_7654,N_9057);
nor U10646 (N_10646,N_8510,N_7688);
nor U10647 (N_10647,N_9683,N_7924);
nor U10648 (N_10648,N_7781,N_8833);
or U10649 (N_10649,N_8024,N_8750);
and U10650 (N_10650,N_7769,N_8677);
and U10651 (N_10651,N_8688,N_8348);
nand U10652 (N_10652,N_9846,N_9349);
nand U10653 (N_10653,N_8545,N_9622);
nor U10654 (N_10654,N_9021,N_7870);
nand U10655 (N_10655,N_7899,N_8408);
nor U10656 (N_10656,N_8837,N_8145);
or U10657 (N_10657,N_8210,N_8607);
or U10658 (N_10658,N_8139,N_9320);
or U10659 (N_10659,N_9605,N_9654);
or U10660 (N_10660,N_8415,N_9137);
nor U10661 (N_10661,N_9002,N_9493);
nand U10662 (N_10662,N_8877,N_8504);
xnor U10663 (N_10663,N_8026,N_9133);
nor U10664 (N_10664,N_7657,N_9184);
and U10665 (N_10665,N_8413,N_9482);
and U10666 (N_10666,N_8449,N_8274);
nand U10667 (N_10667,N_9303,N_8242);
nor U10668 (N_10668,N_9759,N_8387);
nand U10669 (N_10669,N_8758,N_8447);
nor U10670 (N_10670,N_9413,N_7901);
xor U10671 (N_10671,N_7676,N_9822);
nand U10672 (N_10672,N_9857,N_9073);
nor U10673 (N_10673,N_9027,N_7995);
nand U10674 (N_10674,N_9012,N_9685);
and U10675 (N_10675,N_8312,N_9619);
and U10676 (N_10676,N_7540,N_8388);
and U10677 (N_10677,N_9106,N_8014);
xnor U10678 (N_10678,N_9123,N_7549);
nor U10679 (N_10679,N_8068,N_9050);
nor U10680 (N_10680,N_8578,N_9324);
nand U10681 (N_10681,N_8557,N_9549);
xor U10682 (N_10682,N_8444,N_8576);
xnor U10683 (N_10683,N_8923,N_9516);
xnor U10684 (N_10684,N_9559,N_9978);
or U10685 (N_10685,N_9253,N_9153);
nand U10686 (N_10686,N_8285,N_9971);
and U10687 (N_10687,N_7644,N_8864);
or U10688 (N_10688,N_9747,N_8679);
nor U10689 (N_10689,N_8861,N_7557);
or U10690 (N_10690,N_9777,N_7972);
nand U10691 (N_10691,N_7976,N_9018);
xnor U10692 (N_10692,N_7775,N_9417);
nand U10693 (N_10693,N_9474,N_8240);
and U10694 (N_10694,N_8732,N_7652);
nor U10695 (N_10695,N_8665,N_8968);
and U10696 (N_10696,N_7784,N_9961);
nor U10697 (N_10697,N_8133,N_7569);
xor U10698 (N_10698,N_9424,N_8414);
or U10699 (N_10699,N_9746,N_9713);
or U10700 (N_10700,N_9235,N_9964);
and U10701 (N_10701,N_9481,N_8187);
nand U10702 (N_10702,N_8480,N_8614);
or U10703 (N_10703,N_8625,N_9607);
xnor U10704 (N_10704,N_8572,N_9507);
and U10705 (N_10705,N_8717,N_8630);
nor U10706 (N_10706,N_7640,N_9653);
and U10707 (N_10707,N_9898,N_8300);
nand U10708 (N_10708,N_9695,N_8003);
nand U10709 (N_10709,N_8905,N_8016);
or U10710 (N_10710,N_8692,N_8176);
or U10711 (N_10711,N_8934,N_7777);
nand U10712 (N_10712,N_9407,N_8667);
or U10713 (N_10713,N_9551,N_7746);
or U10714 (N_10714,N_7539,N_9107);
nand U10715 (N_10715,N_8916,N_7685);
or U10716 (N_10716,N_9186,N_8179);
xnor U10717 (N_10717,N_8591,N_9268);
nand U10718 (N_10718,N_9925,N_8791);
and U10719 (N_10719,N_9188,N_8909);
nor U10720 (N_10720,N_8232,N_8742);
nor U10721 (N_10721,N_8981,N_9922);
xnor U10722 (N_10722,N_9610,N_8879);
nand U10723 (N_10723,N_7860,N_8377);
and U10724 (N_10724,N_8066,N_8606);
or U10725 (N_10725,N_8350,N_8992);
or U10726 (N_10726,N_9087,N_8359);
nand U10727 (N_10727,N_7572,N_7671);
xnor U10728 (N_10728,N_8354,N_9642);
or U10729 (N_10729,N_8277,N_7846);
nor U10730 (N_10730,N_7795,N_7741);
nand U10731 (N_10731,N_8284,N_9786);
or U10732 (N_10732,N_9719,N_8691);
and U10733 (N_10733,N_7763,N_7873);
xnor U10734 (N_10734,N_9825,N_7892);
nor U10735 (N_10735,N_8237,N_9039);
or U10736 (N_10736,N_9484,N_9132);
nor U10737 (N_10737,N_8184,N_9308);
nand U10738 (N_10738,N_8188,N_8844);
and U10739 (N_10739,N_9470,N_9690);
and U10740 (N_10740,N_9457,N_8980);
or U10741 (N_10741,N_9714,N_8189);
nand U10742 (N_10742,N_8654,N_9554);
xor U10743 (N_10743,N_9092,N_8151);
nand U10744 (N_10744,N_7848,N_8217);
nand U10745 (N_10745,N_8088,N_9350);
and U10746 (N_10746,N_9834,N_8964);
nor U10747 (N_10747,N_7562,N_9445);
nand U10748 (N_10748,N_8083,N_8069);
or U10749 (N_10749,N_8355,N_8379);
or U10750 (N_10750,N_9375,N_9882);
or U10751 (N_10751,N_8807,N_9325);
and U10752 (N_10752,N_7874,N_8793);
and U10753 (N_10753,N_7933,N_8983);
and U10754 (N_10754,N_9923,N_8490);
and U10755 (N_10755,N_9089,N_8160);
xor U10756 (N_10756,N_7845,N_8883);
nand U10757 (N_10757,N_8157,N_7521);
or U10758 (N_10758,N_8629,N_8768);
nor U10759 (N_10759,N_7952,N_7915);
and U10760 (N_10760,N_8549,N_7538);
and U10761 (N_10761,N_9673,N_7653);
and U10762 (N_10762,N_7872,N_9583);
xnor U10763 (N_10763,N_7908,N_9168);
xor U10764 (N_10764,N_7931,N_7750);
and U10765 (N_10765,N_7532,N_8220);
xor U10766 (N_10766,N_7747,N_8794);
or U10767 (N_10767,N_7692,N_9254);
xnor U10768 (N_10768,N_8890,N_8728);
and U10769 (N_10769,N_8037,N_7773);
nand U10770 (N_10770,N_8777,N_7877);
and U10771 (N_10771,N_9580,N_7943);
nand U10772 (N_10772,N_8863,N_9371);
and U10773 (N_10773,N_7650,N_8720);
nor U10774 (N_10774,N_8547,N_9348);
nor U10775 (N_10775,N_8659,N_8315);
nor U10776 (N_10776,N_8531,N_9951);
nor U10777 (N_10777,N_8767,N_7833);
nand U10778 (N_10778,N_9664,N_8790);
nor U10779 (N_10779,N_8458,N_9412);
nor U10780 (N_10780,N_8297,N_9066);
nand U10781 (N_10781,N_8104,N_8984);
nor U10782 (N_10782,N_9469,N_9312);
nand U10783 (N_10783,N_8944,N_7684);
nand U10784 (N_10784,N_9396,N_8780);
nor U10785 (N_10785,N_9753,N_8314);
or U10786 (N_10786,N_7946,N_8856);
nor U10787 (N_10787,N_9477,N_8740);
and U10788 (N_10788,N_8358,N_8224);
nand U10789 (N_10789,N_8008,N_8111);
nand U10790 (N_10790,N_9506,N_8705);
or U10791 (N_10791,N_9359,N_8182);
or U10792 (N_10792,N_9881,N_8031);
xor U10793 (N_10793,N_7666,N_7830);
and U10794 (N_10794,N_8820,N_9780);
and U10795 (N_10795,N_9317,N_7847);
nor U10796 (N_10796,N_9081,N_8301);
or U10797 (N_10797,N_9130,N_7947);
nand U10798 (N_10798,N_8595,N_9044);
and U10799 (N_10799,N_9761,N_8788);
and U10800 (N_10800,N_8976,N_9868);
xor U10801 (N_10801,N_8309,N_8258);
or U10802 (N_10802,N_8517,N_8664);
and U10803 (N_10803,N_7555,N_9827);
nand U10804 (N_10804,N_7637,N_8064);
xnor U10805 (N_10805,N_7910,N_9739);
or U10806 (N_10806,N_7511,N_9862);
xor U10807 (N_10807,N_8860,N_9948);
xor U10808 (N_10808,N_9437,N_9252);
or U10809 (N_10809,N_9214,N_8609);
and U10810 (N_10810,N_9198,N_7842);
or U10811 (N_10811,N_9604,N_8846);
xor U10812 (N_10812,N_9134,N_9304);
xor U10813 (N_10813,N_9223,N_8127);
xnor U10814 (N_10814,N_8956,N_8637);
xor U10815 (N_10815,N_8460,N_9885);
xnor U10816 (N_10816,N_9866,N_9125);
and U10817 (N_10817,N_9144,N_7651);
nor U10818 (N_10818,N_9247,N_9131);
xor U10819 (N_10819,N_8894,N_8373);
or U10820 (N_10820,N_8760,N_7986);
or U10821 (N_10821,N_9836,N_8977);
and U10822 (N_10822,N_8600,N_8207);
or U10823 (N_10823,N_9943,N_7674);
nand U10824 (N_10824,N_8295,N_8367);
nor U10825 (N_10825,N_7698,N_7679);
nor U10826 (N_10826,N_8562,N_8671);
nor U10827 (N_10827,N_8755,N_7500);
nor U10828 (N_10828,N_8342,N_9009);
nand U10829 (N_10829,N_7918,N_9112);
nor U10830 (N_10830,N_9776,N_7909);
nand U10831 (N_10831,N_9571,N_8622);
and U10832 (N_10832,N_8181,N_7743);
or U10833 (N_10833,N_9023,N_8648);
or U10834 (N_10834,N_8509,N_9891);
nand U10835 (N_10835,N_8298,N_9182);
and U10836 (N_10836,N_8678,N_9386);
nor U10837 (N_10837,N_8588,N_9151);
nor U10838 (N_10838,N_8017,N_8817);
nand U10839 (N_10839,N_8850,N_9104);
or U10840 (N_10840,N_9552,N_9175);
nor U10841 (N_10841,N_9463,N_8669);
xnor U10842 (N_10842,N_9258,N_8580);
or U10843 (N_10843,N_7828,N_9595);
or U10844 (N_10844,N_8554,N_8682);
nor U10845 (N_10845,N_9155,N_8525);
nand U10846 (N_10846,N_9899,N_9627);
or U10847 (N_10847,N_7843,N_9124);
nor U10848 (N_10848,N_9769,N_8918);
nor U10849 (N_10849,N_8961,N_9261);
nor U10850 (N_10850,N_8997,N_8647);
xnor U10851 (N_10851,N_8365,N_8006);
or U10852 (N_10852,N_9311,N_9802);
nor U10853 (N_10853,N_8762,N_9910);
or U10854 (N_10854,N_8052,N_8019);
nand U10855 (N_10855,N_8906,N_7984);
nand U10856 (N_10856,N_7694,N_9007);
xor U10857 (N_10857,N_8443,N_9955);
and U10858 (N_10858,N_8253,N_8436);
nand U10859 (N_10859,N_8399,N_9005);
xnor U10860 (N_10860,N_9272,N_8079);
nand U10861 (N_10861,N_8644,N_9794);
and U10862 (N_10862,N_7631,N_7642);
nor U10863 (N_10863,N_8349,N_7619);
nand U10864 (N_10864,N_9241,N_9275);
and U10865 (N_10865,N_9956,N_7818);
xor U10866 (N_10866,N_9562,N_9486);
or U10867 (N_10867,N_8594,N_7956);
xnor U10868 (N_10868,N_8812,N_7876);
and U10869 (N_10869,N_8094,N_9382);
and U10870 (N_10870,N_9828,N_8455);
nor U10871 (N_10871,N_7565,N_8251);
nor U10872 (N_10872,N_7973,N_7791);
or U10873 (N_10873,N_7761,N_8507);
or U10874 (N_10874,N_8533,N_7887);
nand U10875 (N_10875,N_8175,N_8402);
nor U10876 (N_10876,N_7635,N_7519);
xor U10877 (N_10877,N_7585,N_8620);
xnor U10878 (N_10878,N_9586,N_9803);
nor U10879 (N_10879,N_9460,N_8332);
and U10880 (N_10880,N_7812,N_7938);
or U10881 (N_10881,N_7879,N_8826);
and U10882 (N_10882,N_8294,N_8670);
nand U10883 (N_10883,N_8020,N_9823);
or U10884 (N_10884,N_8305,N_9639);
nand U10885 (N_10885,N_8936,N_8775);
and U10886 (N_10886,N_9810,N_9841);
and U10887 (N_10887,N_7686,N_9542);
or U10888 (N_10888,N_7914,N_9286);
nand U10889 (N_10889,N_9443,N_9161);
and U10890 (N_10890,N_9773,N_8899);
nor U10891 (N_10891,N_9696,N_9319);
xnor U10892 (N_10892,N_9189,N_7664);
nand U10893 (N_10893,N_7605,N_9869);
or U10894 (N_10894,N_8073,N_9038);
nor U10895 (N_10895,N_8876,N_8087);
and U10896 (N_10896,N_9267,N_8472);
nor U10897 (N_10897,N_7542,N_7545);
or U10898 (N_10898,N_8110,N_9771);
and U10899 (N_10899,N_9617,N_8978);
nor U10900 (N_10900,N_9138,N_8751);
xor U10901 (N_10901,N_8806,N_9064);
and U10902 (N_10902,N_9211,N_9306);
nand U10903 (N_10903,N_8391,N_9292);
xor U10904 (N_10904,N_8799,N_9310);
nand U10905 (N_10905,N_8491,N_9531);
xor U10906 (N_10906,N_8776,N_9638);
and U10907 (N_10907,N_8693,N_8070);
nor U10908 (N_10908,N_9998,N_9072);
xor U10909 (N_10909,N_9167,N_9624);
xor U10910 (N_10910,N_7691,N_7573);
or U10911 (N_10911,N_9787,N_7559);
nand U10912 (N_10912,N_7502,N_9218);
nand U10913 (N_10913,N_8494,N_8200);
xnor U10914 (N_10914,N_8985,N_8838);
nor U10915 (N_10915,N_9145,N_9449);
xnor U10916 (N_10916,N_7695,N_9894);
xor U10917 (N_10917,N_7751,N_9870);
nand U10918 (N_10918,N_9534,N_9398);
and U10919 (N_10919,N_9079,N_9392);
nand U10920 (N_10920,N_7740,N_7779);
or U10921 (N_10921,N_9179,N_7799);
or U10922 (N_10922,N_9264,N_8935);
or U10923 (N_10923,N_8178,N_9612);
xnor U10924 (N_10924,N_8869,N_9946);
nor U10925 (N_10925,N_8520,N_9265);
nor U10926 (N_10926,N_9884,N_9781);
xor U10927 (N_10927,N_8264,N_9608);
xor U10928 (N_10928,N_9676,N_8747);
nand U10929 (N_10929,N_9754,N_8437);
nand U10930 (N_10930,N_7745,N_9533);
or U10931 (N_10931,N_9650,N_9603);
and U10932 (N_10932,N_8257,N_9069);
and U10933 (N_10933,N_9976,N_9807);
and U10934 (N_10934,N_8244,N_8697);
xor U10935 (N_10935,N_9861,N_9900);
nor U10936 (N_10936,N_9094,N_8376);
xor U10937 (N_10937,N_8306,N_7522);
or U10938 (N_10938,N_9030,N_8103);
and U10939 (N_10939,N_9297,N_9599);
nor U10940 (N_10940,N_8915,N_9936);
and U10941 (N_10941,N_9927,N_9801);
or U10942 (N_10942,N_9410,N_8419);
xnor U10943 (N_10943,N_9745,N_9061);
xor U10944 (N_10944,N_7724,N_8405);
or U10945 (N_10945,N_7707,N_8476);
nor U10946 (N_10946,N_9528,N_7897);
nor U10947 (N_10947,N_8462,N_9372);
and U10948 (N_10948,N_9128,N_9926);
nand U10949 (N_10949,N_7888,N_7581);
xor U10950 (N_10950,N_9871,N_8714);
xnor U10951 (N_10951,N_8432,N_8821);
or U10952 (N_10952,N_8055,N_7618);
xor U10953 (N_10953,N_8963,N_7992);
and U10954 (N_10954,N_9055,N_7643);
nand U10955 (N_10955,N_9880,N_9232);
and U10956 (N_10956,N_7951,N_7831);
xnor U10957 (N_10957,N_8047,N_9508);
nand U10958 (N_10958,N_8118,N_8711);
nor U10959 (N_10959,N_8164,N_9290);
nand U10960 (N_10960,N_9567,N_8374);
nand U10961 (N_10961,N_9811,N_7703);
nor U10962 (N_10962,N_8734,N_8147);
or U10963 (N_10963,N_8028,N_9291);
nand U10964 (N_10964,N_8920,N_9453);
nor U10965 (N_10965,N_8592,N_7850);
nand U10966 (N_10966,N_9710,N_8535);
or U10967 (N_10967,N_9418,N_9873);
and U10968 (N_10968,N_7667,N_8039);
nor U10969 (N_10969,N_9086,N_8261);
xor U10970 (N_10970,N_9309,N_9523);
and U10971 (N_10971,N_9346,N_8228);
and U10972 (N_10972,N_8859,N_8227);
or U10973 (N_10973,N_7574,N_8045);
or U10974 (N_10974,N_7853,N_9126);
xnor U10975 (N_10975,N_9379,N_8153);
nor U10976 (N_10976,N_7622,N_9380);
and U10977 (N_10977,N_8423,N_8598);
nand U10978 (N_10978,N_9527,N_8004);
or U10979 (N_10979,N_7985,N_8962);
and U10980 (N_10980,N_7970,N_9432);
or U10981 (N_10981,N_8772,N_8196);
nor U10982 (N_10982,N_8652,N_8603);
nand U10983 (N_10983,N_8050,N_7533);
and U10984 (N_10984,N_9656,N_8197);
or U10985 (N_10985,N_8121,N_8203);
and U10986 (N_10986,N_8942,N_8640);
xnor U10987 (N_10987,N_9119,N_8059);
and U10988 (N_10988,N_9495,N_7950);
xor U10989 (N_10989,N_9782,N_9600);
xor U10990 (N_10990,N_9722,N_9791);
nand U10991 (N_10991,N_7925,N_9517);
and U10992 (N_10992,N_9322,N_9991);
nor U10993 (N_10993,N_8599,N_8488);
and U10994 (N_10994,N_9327,N_7822);
and U10995 (N_10995,N_9354,N_8565);
or U10996 (N_10996,N_9316,N_9330);
xnor U10997 (N_10997,N_8271,N_7825);
xor U10998 (N_10998,N_9141,N_9288);
nand U10999 (N_10999,N_9546,N_8036);
or U11000 (N_11000,N_9171,N_8322);
nand U11001 (N_11001,N_9199,N_9518);
nor U11002 (N_11002,N_9163,N_7898);
xor U11003 (N_11003,N_9340,N_8882);
or U11004 (N_11004,N_8922,N_8425);
nand U11005 (N_11005,N_7704,N_9472);
and U11006 (N_11006,N_9143,N_8752);
nand U11007 (N_11007,N_8427,N_8456);
and U11008 (N_11008,N_8646,N_8989);
nor U11009 (N_11009,N_9904,N_9915);
and U11010 (N_11010,N_7852,N_8574);
or U11011 (N_11011,N_9142,N_9644);
and U11012 (N_11012,N_7531,N_7939);
and U11013 (N_11013,N_9625,N_9597);
nand U11014 (N_11014,N_9419,N_9987);
xnor U11015 (N_11015,N_8313,N_9560);
nor U11016 (N_11016,N_9213,N_9347);
and U11017 (N_11017,N_9159,N_9821);
and U11018 (N_11018,N_9514,N_8250);
and U11019 (N_11019,N_9117,N_9441);
nand U11020 (N_11020,N_7974,N_9022);
nor U11021 (N_11021,N_9377,N_8907);
xnor U11022 (N_11022,N_8657,N_9895);
nor U11023 (N_11023,N_9544,N_8396);
xor U11024 (N_11024,N_9783,N_8183);
or U11025 (N_11025,N_7979,N_8813);
xnor U11026 (N_11026,N_7700,N_9207);
or U11027 (N_11027,N_8043,N_9509);
nand U11028 (N_11028,N_8454,N_8256);
or U11029 (N_11029,N_7921,N_9192);
xnor U11030 (N_11030,N_9537,N_7623);
nor U11031 (N_11031,N_7589,N_8901);
nor U11032 (N_11032,N_7840,N_9606);
nand U11033 (N_11033,N_8725,N_7959);
nor U11034 (N_11034,N_7600,N_8633);
nor U11035 (N_11035,N_8439,N_9406);
and U11036 (N_11036,N_8561,N_9853);
and U11037 (N_11037,N_9672,N_9095);
or U11038 (N_11038,N_7772,N_7935);
nor U11039 (N_11039,N_8958,N_8364);
nor U11040 (N_11040,N_8803,N_8255);
nor U11041 (N_11041,N_9628,N_9750);
nor U11042 (N_11042,N_8248,N_7632);
nand U11043 (N_11043,N_8033,N_9176);
and U11044 (N_11044,N_9635,N_9114);
nor U11045 (N_11045,N_8867,N_8492);
nor U11046 (N_11046,N_8756,N_9440);
nor U11047 (N_11047,N_7530,N_9875);
or U11048 (N_11048,N_7816,N_8552);
and U11049 (N_11049,N_8840,N_7733);
xor U11050 (N_11050,N_9373,N_8825);
and U11051 (N_11051,N_8765,N_9699);
nor U11052 (N_11052,N_9830,N_9172);
or U11053 (N_11053,N_8783,N_9702);
or U11054 (N_11054,N_9902,N_8368);
nand U11055 (N_11055,N_9281,N_7649);
nor U11056 (N_11056,N_9679,N_8048);
xnor U11057 (N_11057,N_8929,N_7813);
xor U11058 (N_11058,N_8680,N_7615);
and U11059 (N_11059,N_8849,N_8307);
and U11060 (N_11060,N_8040,N_9205);
xnor U11061 (N_11061,N_9630,N_9421);
and U11062 (N_11062,N_8347,N_8122);
nor U11063 (N_11063,N_7961,N_9504);
nand U11064 (N_11064,N_7604,N_9200);
or U11065 (N_11065,N_7607,N_7693);
or U11066 (N_11066,N_9658,N_8782);
nor U11067 (N_11067,N_8757,N_9122);
xor U11068 (N_11068,N_8317,N_7526);
nand U11069 (N_11069,N_8056,N_9997);
and U11070 (N_11070,N_9565,N_8211);
nand U11071 (N_11071,N_7890,N_9013);
and U11072 (N_11072,N_7754,N_8403);
or U11073 (N_11073,N_9358,N_8212);
or U11074 (N_11074,N_7658,N_9593);
or U11075 (N_11075,N_7868,N_7786);
nand U11076 (N_11076,N_8435,N_7556);
nand U11077 (N_11077,N_9333,N_9500);
xor U11078 (N_11078,N_9010,N_9467);
nand U11079 (N_11079,N_8816,N_8198);
and U11080 (N_11080,N_8356,N_7737);
or U11081 (N_11081,N_8015,N_9850);
xor U11082 (N_11082,N_7683,N_9233);
xor U11083 (N_11083,N_8548,N_7932);
and U11084 (N_11084,N_8888,N_9284);
xor U11085 (N_11085,N_8161,N_8555);
nor U11086 (N_11086,N_8304,N_9817);
or U11087 (N_11087,N_7722,N_8957);
xor U11088 (N_11088,N_8539,N_8774);
xnor U11089 (N_11089,N_8497,N_8389);
or U11090 (N_11090,N_9435,N_8172);
nand U11091 (N_11091,N_9035,N_9557);
and U11092 (N_11092,N_8937,N_7797);
xor U11093 (N_11093,N_9512,N_9360);
nand U11094 (N_11094,N_9620,N_9729);
nor U11095 (N_11095,N_7689,N_9967);
nor U11096 (N_11096,N_7593,N_9668);
nor U11097 (N_11097,N_9269,N_9985);
or U11098 (N_11098,N_9572,N_8216);
nor U11099 (N_11099,N_9613,N_9444);
nand U11100 (N_11100,N_9462,N_7991);
xor U11101 (N_11101,N_7983,N_9423);
nor U11102 (N_11102,N_7776,N_9085);
and U11103 (N_11103,N_8721,N_9703);
nand U11104 (N_11104,N_7871,N_7598);
nand U11105 (N_11105,N_8847,N_9919);
xnor U11106 (N_11106,N_9157,N_9244);
nand U11107 (N_11107,N_9966,N_7616);
nand U11108 (N_11108,N_8438,N_9174);
nor U11109 (N_11109,N_7967,N_9793);
nand U11110 (N_11110,N_8018,N_8946);
and U11111 (N_11111,N_9778,N_8136);
or U11112 (N_11112,N_8932,N_9718);
and U11113 (N_11113,N_7580,N_7820);
xnor U11114 (N_11114,N_9629,N_7508);
xnor U11115 (N_11115,N_7809,N_8362);
and U11116 (N_11116,N_9838,N_7883);
or U11117 (N_11117,N_7735,N_9996);
nand U11118 (N_11118,N_7849,N_9687);
or U11119 (N_11119,N_8919,N_7734);
and U11120 (N_11120,N_7601,N_9051);
nand U11121 (N_11121,N_9273,N_9054);
or U11122 (N_11122,N_9400,N_7755);
xor U11123 (N_11123,N_7884,N_8511);
xor U11124 (N_11124,N_7701,N_7591);
xnor U11125 (N_11125,N_8384,N_9982);
nor U11126 (N_11126,N_7805,N_8223);
and U11127 (N_11127,N_8558,N_9766);
nand U11128 (N_11128,N_8809,N_8521);
or U11129 (N_11129,N_7960,N_8120);
or U11130 (N_11130,N_7732,N_8974);
xnor U11131 (N_11131,N_9301,N_8830);
xor U11132 (N_11132,N_9983,N_8416);
and U11133 (N_11133,N_9536,N_9381);
xnor U11134 (N_11134,N_7975,N_9225);
nor U11135 (N_11135,N_7881,N_9697);
xnor U11136 (N_11136,N_8683,N_9028);
nand U11137 (N_11137,N_7993,N_9395);
nand U11138 (N_11138,N_7880,N_8784);
nor U11139 (N_11139,N_9203,N_7515);
nand U11140 (N_11140,N_8132,N_9197);
and U11141 (N_11141,N_8067,N_9637);
and U11142 (N_11142,N_7948,N_8926);
and U11143 (N_11143,N_9795,N_7987);
xor U11144 (N_11144,N_9402,N_9370);
nor U11145 (N_11145,N_9465,N_9490);
or U11146 (N_11146,N_7889,N_9980);
nor U11147 (N_11147,N_8575,N_7739);
or U11148 (N_11148,N_8141,N_7744);
nor U11149 (N_11149,N_8150,N_7916);
xnor U11150 (N_11150,N_9804,N_8053);
xor U11151 (N_11151,N_8542,N_9588);
or U11152 (N_11152,N_9160,N_9796);
xnor U11153 (N_11153,N_8608,N_8503);
and U11154 (N_11154,N_9116,N_8769);
xor U11155 (N_11155,N_9538,N_9219);
xnor U11156 (N_11156,N_9999,N_9056);
nor U11157 (N_11157,N_8839,N_8245);
nand U11158 (N_11158,N_8116,N_9809);
nand U11159 (N_11159,N_8280,N_9476);
nand U11160 (N_11160,N_9067,N_8904);
or U11161 (N_11161,N_8835,N_7934);
nand U11162 (N_11162,N_8465,N_7757);
nor U11163 (N_11163,N_9708,N_8201);
nand U11164 (N_11164,N_8733,N_8538);
xor U11165 (N_11165,N_9098,N_9084);
xor U11166 (N_11166,N_9242,N_7566);
or U11167 (N_11167,N_8778,N_8299);
xnor U11168 (N_11168,N_8615,N_8450);
xnor U11169 (N_11169,N_7567,N_8593);
or U11170 (N_11170,N_9981,N_7719);
nand U11171 (N_11171,N_8573,N_8464);
and U11172 (N_11172,N_7765,N_9505);
and U11173 (N_11173,N_8254,N_8704);
nand U11174 (N_11174,N_8075,N_8156);
and U11175 (N_11175,N_8993,N_8011);
or U11176 (N_11176,N_7687,N_9152);
xor U11177 (N_11177,N_9091,N_9663);
or U11178 (N_11178,N_7766,N_8428);
nand U11179 (N_11179,N_8726,N_8247);
and U11180 (N_11180,N_9950,N_9893);
xor U11181 (N_11181,N_9816,N_8672);
or U11182 (N_11182,N_7758,N_8822);
nand U11183 (N_11183,N_8524,N_9671);
or U11184 (N_11184,N_8921,N_8233);
or U11185 (N_11185,N_7824,N_8093);
nor U11186 (N_11186,N_9164,N_9041);
and U11187 (N_11187,N_7528,N_7798);
nor U11188 (N_11188,N_8209,N_9439);
nor U11189 (N_11189,N_9430,N_9149);
or U11190 (N_11190,N_9993,N_8287);
xnor U11191 (N_11191,N_7553,N_9397);
or U11192 (N_11192,N_9256,N_8072);
nor U11193 (N_11193,N_7682,N_8119);
nor U11194 (N_11194,N_8089,N_9289);
or U11195 (N_11195,N_9734,N_7919);
nand U11196 (N_11196,N_8308,N_9615);
xor U11197 (N_11197,N_9388,N_8619);
nor U11198 (N_11198,N_8140,N_8566);
and U11199 (N_11199,N_9212,N_9118);
and U11200 (N_11200,N_9404,N_9522);
nand U11201 (N_11201,N_7638,N_7904);
nand U11202 (N_11202,N_9034,N_7867);
nand U11203 (N_11203,N_8499,N_8519);
xor U11204 (N_11204,N_9785,N_9959);
or U11205 (N_11205,N_9434,N_8032);
or U11206 (N_11206,N_9053,N_7835);
and U11207 (N_11207,N_7509,N_9001);
or U11208 (N_11208,N_7681,N_9763);
nor U11209 (N_11209,N_9391,N_9063);
xnor U11210 (N_11210,N_8501,N_8114);
nor U11211 (N_11211,N_8675,N_8689);
nand U11212 (N_11212,N_8441,N_9178);
or U11213 (N_11213,N_9824,N_9426);
and U11214 (N_11214,N_8259,N_7896);
or U11215 (N_11215,N_8613,N_7808);
nand U11216 (N_11216,N_7789,N_8363);
nor U11217 (N_11217,N_8027,N_8656);
or U11218 (N_11218,N_8206,N_7633);
and U11219 (N_11219,N_8951,N_8484);
xor U11220 (N_11220,N_9140,N_9724);
nand U11221 (N_11221,N_7558,N_8109);
and U11222 (N_11222,N_9682,N_9602);
nor U11223 (N_11223,N_9156,N_8949);
nor U11224 (N_11224,N_8832,N_8453);
nand U11225 (N_11225,N_8496,N_9935);
or U11226 (N_11226,N_9855,N_8397);
xnor U11227 (N_11227,N_8468,N_9973);
and U11228 (N_11228,N_8913,N_9751);
nand U11229 (N_11229,N_8930,N_8753);
and U11230 (N_11230,N_8624,N_9008);
and U11231 (N_11231,N_7563,N_7672);
nor U11232 (N_11232,N_8546,N_9929);
nand U11233 (N_11233,N_9338,N_7900);
and U11234 (N_11234,N_8030,N_9907);
nor U11235 (N_11235,N_8218,N_8718);
xor U11236 (N_11236,N_9422,N_8582);
xor U11237 (N_11237,N_8302,N_9905);
nor U11238 (N_11238,N_7713,N_8288);
and U11239 (N_11239,N_8106,N_7783);
and U11240 (N_11240,N_9487,N_8404);
xnor U11241 (N_11241,N_9026,N_8107);
and U11242 (N_11242,N_8466,N_8831);
nor U11243 (N_11243,N_8819,N_8947);
xnor U11244 (N_11244,N_8590,N_9357);
nand U11245 (N_11245,N_8766,N_7584);
nand U11246 (N_11246,N_7928,N_9921);
nand U11247 (N_11247,N_9519,N_7854);
nor U11248 (N_11248,N_9408,N_8495);
nor U11249 (N_11249,N_9808,N_9577);
xnor U11250 (N_11250,N_8873,N_8805);
or U11251 (N_11251,N_8102,N_9027);
xnor U11252 (N_11252,N_8612,N_8460);
xor U11253 (N_11253,N_8582,N_8783);
nand U11254 (N_11254,N_9123,N_9427);
nor U11255 (N_11255,N_9726,N_9728);
xnor U11256 (N_11256,N_8625,N_9624);
nand U11257 (N_11257,N_8302,N_9189);
nand U11258 (N_11258,N_8796,N_9450);
or U11259 (N_11259,N_8265,N_9469);
nor U11260 (N_11260,N_8269,N_7576);
or U11261 (N_11261,N_8411,N_9253);
nor U11262 (N_11262,N_7799,N_7511);
xor U11263 (N_11263,N_8400,N_9646);
nand U11264 (N_11264,N_9445,N_8971);
or U11265 (N_11265,N_8042,N_8969);
nor U11266 (N_11266,N_8760,N_9276);
xnor U11267 (N_11267,N_8653,N_9410);
or U11268 (N_11268,N_9547,N_8625);
and U11269 (N_11269,N_8356,N_8293);
xor U11270 (N_11270,N_8957,N_8457);
or U11271 (N_11271,N_8383,N_9138);
nor U11272 (N_11272,N_9733,N_9041);
and U11273 (N_11273,N_8541,N_9214);
nand U11274 (N_11274,N_9826,N_8126);
xnor U11275 (N_11275,N_7715,N_9006);
or U11276 (N_11276,N_9471,N_8541);
and U11277 (N_11277,N_8413,N_7548);
nand U11278 (N_11278,N_9408,N_9400);
nor U11279 (N_11279,N_8498,N_7566);
xnor U11280 (N_11280,N_7826,N_8865);
nor U11281 (N_11281,N_9803,N_9937);
or U11282 (N_11282,N_9722,N_9762);
nand U11283 (N_11283,N_9184,N_7962);
xor U11284 (N_11284,N_8361,N_7739);
or U11285 (N_11285,N_8434,N_9949);
nor U11286 (N_11286,N_8728,N_9588);
nor U11287 (N_11287,N_8465,N_8174);
and U11288 (N_11288,N_9181,N_9310);
nor U11289 (N_11289,N_8025,N_8887);
nor U11290 (N_11290,N_9500,N_8398);
nor U11291 (N_11291,N_8547,N_8190);
or U11292 (N_11292,N_8108,N_9412);
or U11293 (N_11293,N_9667,N_8770);
nand U11294 (N_11294,N_8698,N_8813);
nand U11295 (N_11295,N_8655,N_7580);
nor U11296 (N_11296,N_9961,N_8862);
xnor U11297 (N_11297,N_8814,N_8421);
or U11298 (N_11298,N_9646,N_8415);
or U11299 (N_11299,N_7711,N_9981);
nor U11300 (N_11300,N_9815,N_7732);
and U11301 (N_11301,N_8751,N_8919);
or U11302 (N_11302,N_8952,N_8954);
nor U11303 (N_11303,N_9122,N_9530);
xor U11304 (N_11304,N_9485,N_8321);
or U11305 (N_11305,N_8112,N_7784);
xnor U11306 (N_11306,N_7678,N_7557);
nand U11307 (N_11307,N_9571,N_9695);
and U11308 (N_11308,N_7879,N_8700);
and U11309 (N_11309,N_8707,N_9933);
or U11310 (N_11310,N_7600,N_9267);
or U11311 (N_11311,N_8072,N_9380);
nor U11312 (N_11312,N_8446,N_9279);
nor U11313 (N_11313,N_8926,N_8236);
or U11314 (N_11314,N_7907,N_9635);
nor U11315 (N_11315,N_9564,N_7610);
and U11316 (N_11316,N_8445,N_9044);
and U11317 (N_11317,N_9680,N_8622);
xor U11318 (N_11318,N_9053,N_8025);
nand U11319 (N_11319,N_9749,N_7572);
nor U11320 (N_11320,N_8764,N_9333);
and U11321 (N_11321,N_7946,N_8260);
or U11322 (N_11322,N_8681,N_9565);
nand U11323 (N_11323,N_9435,N_9240);
xnor U11324 (N_11324,N_7889,N_7845);
nand U11325 (N_11325,N_8769,N_8171);
and U11326 (N_11326,N_9483,N_9921);
nand U11327 (N_11327,N_8055,N_9116);
xnor U11328 (N_11328,N_8709,N_8602);
nand U11329 (N_11329,N_7931,N_9277);
nand U11330 (N_11330,N_8308,N_8549);
nand U11331 (N_11331,N_7933,N_7664);
xor U11332 (N_11332,N_9048,N_8174);
or U11333 (N_11333,N_7951,N_8373);
and U11334 (N_11334,N_9140,N_9618);
xnor U11335 (N_11335,N_8828,N_8409);
nor U11336 (N_11336,N_9907,N_7535);
xnor U11337 (N_11337,N_8346,N_9042);
nor U11338 (N_11338,N_8241,N_7549);
and U11339 (N_11339,N_9683,N_9841);
and U11340 (N_11340,N_8371,N_9797);
nand U11341 (N_11341,N_7964,N_9446);
nor U11342 (N_11342,N_9206,N_8251);
and U11343 (N_11343,N_8405,N_7885);
nand U11344 (N_11344,N_8002,N_8592);
nand U11345 (N_11345,N_9719,N_7521);
xor U11346 (N_11346,N_7861,N_7586);
or U11347 (N_11347,N_7808,N_9022);
xor U11348 (N_11348,N_9737,N_9096);
xor U11349 (N_11349,N_9743,N_8565);
and U11350 (N_11350,N_8423,N_8519);
nor U11351 (N_11351,N_9847,N_9622);
or U11352 (N_11352,N_9656,N_7918);
and U11353 (N_11353,N_8147,N_8188);
or U11354 (N_11354,N_8206,N_7806);
nor U11355 (N_11355,N_9758,N_7750);
nor U11356 (N_11356,N_9018,N_9028);
nor U11357 (N_11357,N_8582,N_8578);
nor U11358 (N_11358,N_8913,N_8627);
or U11359 (N_11359,N_9862,N_9672);
nor U11360 (N_11360,N_8967,N_8513);
and U11361 (N_11361,N_9441,N_8874);
nor U11362 (N_11362,N_8257,N_8857);
nand U11363 (N_11363,N_8586,N_7993);
or U11364 (N_11364,N_8790,N_7506);
nand U11365 (N_11365,N_8152,N_9779);
or U11366 (N_11366,N_8456,N_8430);
nor U11367 (N_11367,N_8768,N_8274);
xnor U11368 (N_11368,N_8983,N_9029);
nand U11369 (N_11369,N_9174,N_7979);
nor U11370 (N_11370,N_8030,N_9754);
nand U11371 (N_11371,N_9121,N_7760);
nand U11372 (N_11372,N_9145,N_9900);
and U11373 (N_11373,N_9772,N_9395);
nand U11374 (N_11374,N_7598,N_8080);
and U11375 (N_11375,N_8645,N_9127);
and U11376 (N_11376,N_8686,N_8702);
xnor U11377 (N_11377,N_7925,N_8703);
nand U11378 (N_11378,N_8492,N_7838);
xnor U11379 (N_11379,N_9822,N_7600);
nand U11380 (N_11380,N_9623,N_7714);
or U11381 (N_11381,N_9756,N_9102);
and U11382 (N_11382,N_9582,N_8020);
nor U11383 (N_11383,N_9595,N_9473);
nand U11384 (N_11384,N_8450,N_8894);
xor U11385 (N_11385,N_9027,N_8734);
nor U11386 (N_11386,N_8556,N_8097);
or U11387 (N_11387,N_8970,N_9760);
or U11388 (N_11388,N_9244,N_8334);
nand U11389 (N_11389,N_9355,N_9376);
and U11390 (N_11390,N_8634,N_9828);
or U11391 (N_11391,N_9387,N_9316);
nor U11392 (N_11392,N_7830,N_7736);
xor U11393 (N_11393,N_9467,N_9049);
or U11394 (N_11394,N_7537,N_8688);
or U11395 (N_11395,N_8947,N_8087);
xnor U11396 (N_11396,N_8744,N_9528);
or U11397 (N_11397,N_9728,N_9844);
nand U11398 (N_11398,N_9343,N_9950);
nand U11399 (N_11399,N_9715,N_8010);
xor U11400 (N_11400,N_7822,N_8318);
xor U11401 (N_11401,N_9429,N_9135);
or U11402 (N_11402,N_8261,N_7500);
xor U11403 (N_11403,N_8457,N_7656);
or U11404 (N_11404,N_9250,N_8769);
or U11405 (N_11405,N_8412,N_8956);
nand U11406 (N_11406,N_7841,N_8824);
nor U11407 (N_11407,N_7920,N_9032);
nor U11408 (N_11408,N_7957,N_9231);
xnor U11409 (N_11409,N_9280,N_8011);
nor U11410 (N_11410,N_9206,N_9392);
or U11411 (N_11411,N_7850,N_9495);
or U11412 (N_11412,N_9453,N_9468);
or U11413 (N_11413,N_9376,N_7940);
nand U11414 (N_11414,N_8196,N_9641);
or U11415 (N_11415,N_8607,N_8691);
nor U11416 (N_11416,N_9134,N_9222);
xor U11417 (N_11417,N_8890,N_8068);
xnor U11418 (N_11418,N_8222,N_9831);
and U11419 (N_11419,N_8022,N_7972);
and U11420 (N_11420,N_8313,N_8231);
nor U11421 (N_11421,N_9967,N_9448);
nor U11422 (N_11422,N_8681,N_8986);
and U11423 (N_11423,N_9028,N_7528);
nand U11424 (N_11424,N_8948,N_8218);
or U11425 (N_11425,N_9086,N_7866);
xor U11426 (N_11426,N_9524,N_9031);
and U11427 (N_11427,N_7800,N_8941);
nand U11428 (N_11428,N_8267,N_9685);
or U11429 (N_11429,N_9120,N_9634);
or U11430 (N_11430,N_7509,N_8636);
and U11431 (N_11431,N_9997,N_8171);
xnor U11432 (N_11432,N_8600,N_7764);
and U11433 (N_11433,N_8935,N_7934);
or U11434 (N_11434,N_7587,N_9274);
nor U11435 (N_11435,N_7676,N_8574);
nor U11436 (N_11436,N_8119,N_9613);
nor U11437 (N_11437,N_9834,N_8801);
and U11438 (N_11438,N_8993,N_9977);
nand U11439 (N_11439,N_9281,N_8739);
xnor U11440 (N_11440,N_8305,N_8577);
xnor U11441 (N_11441,N_9464,N_9094);
or U11442 (N_11442,N_9338,N_8966);
xnor U11443 (N_11443,N_8638,N_9592);
nand U11444 (N_11444,N_8393,N_9699);
xnor U11445 (N_11445,N_9315,N_8632);
xor U11446 (N_11446,N_9056,N_9046);
xor U11447 (N_11447,N_7652,N_8507);
nand U11448 (N_11448,N_9259,N_8870);
nand U11449 (N_11449,N_7817,N_8648);
nand U11450 (N_11450,N_8251,N_7760);
or U11451 (N_11451,N_9822,N_9241);
nor U11452 (N_11452,N_8374,N_8426);
nand U11453 (N_11453,N_8808,N_8910);
and U11454 (N_11454,N_9848,N_8168);
and U11455 (N_11455,N_8187,N_9036);
nor U11456 (N_11456,N_8692,N_7583);
or U11457 (N_11457,N_9885,N_9822);
or U11458 (N_11458,N_8846,N_9000);
nor U11459 (N_11459,N_8222,N_8886);
xor U11460 (N_11460,N_7634,N_7945);
or U11461 (N_11461,N_9466,N_7661);
nand U11462 (N_11462,N_7542,N_7517);
xor U11463 (N_11463,N_9347,N_8034);
nand U11464 (N_11464,N_9947,N_8078);
nor U11465 (N_11465,N_8823,N_8805);
nand U11466 (N_11466,N_8673,N_9949);
or U11467 (N_11467,N_7856,N_9808);
or U11468 (N_11468,N_8255,N_8718);
xnor U11469 (N_11469,N_9510,N_7924);
nand U11470 (N_11470,N_8023,N_7999);
xnor U11471 (N_11471,N_9835,N_8380);
xor U11472 (N_11472,N_9255,N_9228);
nor U11473 (N_11473,N_8892,N_9875);
nand U11474 (N_11474,N_9619,N_9647);
xor U11475 (N_11475,N_8001,N_9365);
nor U11476 (N_11476,N_7565,N_8751);
or U11477 (N_11477,N_9382,N_7573);
or U11478 (N_11478,N_8022,N_8382);
nand U11479 (N_11479,N_7806,N_8112);
nand U11480 (N_11480,N_8017,N_9421);
xnor U11481 (N_11481,N_8196,N_8160);
nand U11482 (N_11482,N_9377,N_8309);
xor U11483 (N_11483,N_9647,N_8091);
or U11484 (N_11484,N_8823,N_8749);
nor U11485 (N_11485,N_9068,N_8390);
or U11486 (N_11486,N_9362,N_7776);
nand U11487 (N_11487,N_8233,N_9208);
nand U11488 (N_11488,N_8429,N_9910);
nor U11489 (N_11489,N_9372,N_9312);
xor U11490 (N_11490,N_8858,N_8483);
nand U11491 (N_11491,N_9059,N_8561);
and U11492 (N_11492,N_7832,N_7735);
and U11493 (N_11493,N_8725,N_7933);
xnor U11494 (N_11494,N_8828,N_8629);
or U11495 (N_11495,N_9124,N_8458);
nand U11496 (N_11496,N_9438,N_8482);
and U11497 (N_11497,N_9177,N_8781);
nand U11498 (N_11498,N_7860,N_8437);
and U11499 (N_11499,N_8726,N_7948);
and U11500 (N_11500,N_9778,N_8767);
nor U11501 (N_11501,N_9251,N_8915);
xor U11502 (N_11502,N_9556,N_9685);
nor U11503 (N_11503,N_9335,N_9193);
xnor U11504 (N_11504,N_7758,N_7752);
nand U11505 (N_11505,N_8422,N_7958);
nand U11506 (N_11506,N_8783,N_7680);
and U11507 (N_11507,N_8797,N_7691);
or U11508 (N_11508,N_9339,N_8426);
nand U11509 (N_11509,N_8794,N_9393);
nor U11510 (N_11510,N_8440,N_8399);
or U11511 (N_11511,N_7730,N_8509);
or U11512 (N_11512,N_9290,N_8026);
or U11513 (N_11513,N_8178,N_8029);
xor U11514 (N_11514,N_9633,N_9060);
nor U11515 (N_11515,N_9861,N_8693);
and U11516 (N_11516,N_8742,N_9973);
and U11517 (N_11517,N_9518,N_9281);
xor U11518 (N_11518,N_9068,N_8213);
nand U11519 (N_11519,N_9846,N_7500);
xor U11520 (N_11520,N_9869,N_9913);
or U11521 (N_11521,N_7697,N_9561);
xnor U11522 (N_11522,N_7859,N_9729);
xor U11523 (N_11523,N_8435,N_7653);
or U11524 (N_11524,N_8898,N_8315);
and U11525 (N_11525,N_9239,N_9216);
nor U11526 (N_11526,N_8940,N_8249);
or U11527 (N_11527,N_8567,N_9777);
nand U11528 (N_11528,N_9576,N_9957);
or U11529 (N_11529,N_7868,N_8759);
nor U11530 (N_11530,N_8623,N_9776);
nor U11531 (N_11531,N_9378,N_9571);
and U11532 (N_11532,N_9606,N_8406);
and U11533 (N_11533,N_7919,N_8025);
xnor U11534 (N_11534,N_9412,N_9690);
and U11535 (N_11535,N_8677,N_8200);
and U11536 (N_11536,N_7538,N_8795);
nand U11537 (N_11537,N_7873,N_9645);
nor U11538 (N_11538,N_8105,N_8462);
xnor U11539 (N_11539,N_9611,N_9907);
or U11540 (N_11540,N_8763,N_8517);
nand U11541 (N_11541,N_9203,N_9977);
or U11542 (N_11542,N_8394,N_9790);
or U11543 (N_11543,N_7731,N_9878);
nor U11544 (N_11544,N_9205,N_9934);
nor U11545 (N_11545,N_9278,N_8178);
nand U11546 (N_11546,N_8489,N_7692);
nor U11547 (N_11547,N_9749,N_7862);
nand U11548 (N_11548,N_8292,N_8052);
nor U11549 (N_11549,N_9974,N_9868);
nand U11550 (N_11550,N_9191,N_9757);
or U11551 (N_11551,N_8039,N_8464);
and U11552 (N_11552,N_9732,N_8599);
nor U11553 (N_11553,N_8486,N_8277);
and U11554 (N_11554,N_8828,N_9044);
xnor U11555 (N_11555,N_8270,N_8237);
nor U11556 (N_11556,N_9365,N_8764);
nand U11557 (N_11557,N_8500,N_8499);
nand U11558 (N_11558,N_9238,N_7682);
or U11559 (N_11559,N_7999,N_8033);
nand U11560 (N_11560,N_7630,N_9580);
and U11561 (N_11561,N_9860,N_7658);
and U11562 (N_11562,N_9346,N_9492);
nor U11563 (N_11563,N_8305,N_9888);
nand U11564 (N_11564,N_8434,N_8659);
and U11565 (N_11565,N_7984,N_9382);
xnor U11566 (N_11566,N_7921,N_9115);
nand U11567 (N_11567,N_9066,N_8128);
xnor U11568 (N_11568,N_8920,N_8946);
or U11569 (N_11569,N_9167,N_9672);
and U11570 (N_11570,N_8211,N_9009);
or U11571 (N_11571,N_8501,N_7859);
or U11572 (N_11572,N_8501,N_9118);
xor U11573 (N_11573,N_7653,N_8244);
xor U11574 (N_11574,N_8962,N_9926);
nor U11575 (N_11575,N_7526,N_7538);
or U11576 (N_11576,N_8073,N_8685);
or U11577 (N_11577,N_7589,N_9598);
xor U11578 (N_11578,N_7890,N_7886);
nor U11579 (N_11579,N_7845,N_9938);
nor U11580 (N_11580,N_8071,N_9056);
or U11581 (N_11581,N_8953,N_8290);
nand U11582 (N_11582,N_8897,N_9419);
nor U11583 (N_11583,N_9501,N_8608);
nand U11584 (N_11584,N_8784,N_7888);
nor U11585 (N_11585,N_9575,N_8012);
or U11586 (N_11586,N_9247,N_8100);
xor U11587 (N_11587,N_8583,N_8102);
xnor U11588 (N_11588,N_9524,N_9081);
or U11589 (N_11589,N_8575,N_8883);
xnor U11590 (N_11590,N_8705,N_9100);
xor U11591 (N_11591,N_9945,N_7546);
and U11592 (N_11592,N_8051,N_7659);
xnor U11593 (N_11593,N_8866,N_8250);
and U11594 (N_11594,N_8382,N_7919);
and U11595 (N_11595,N_9836,N_8542);
and U11596 (N_11596,N_8247,N_9536);
xnor U11597 (N_11597,N_8799,N_9319);
and U11598 (N_11598,N_9231,N_9915);
and U11599 (N_11599,N_9993,N_8966);
or U11600 (N_11600,N_9301,N_9984);
nor U11601 (N_11601,N_9312,N_9949);
or U11602 (N_11602,N_8816,N_8884);
xnor U11603 (N_11603,N_9388,N_7628);
nand U11604 (N_11604,N_8297,N_8841);
and U11605 (N_11605,N_9709,N_9182);
or U11606 (N_11606,N_8986,N_9345);
or U11607 (N_11607,N_9967,N_9389);
or U11608 (N_11608,N_8735,N_8245);
xnor U11609 (N_11609,N_8980,N_9405);
and U11610 (N_11610,N_8166,N_8451);
nand U11611 (N_11611,N_9944,N_8053);
nand U11612 (N_11612,N_9880,N_8176);
nor U11613 (N_11613,N_8690,N_7913);
xor U11614 (N_11614,N_8661,N_9163);
or U11615 (N_11615,N_8710,N_7713);
xnor U11616 (N_11616,N_9400,N_9148);
xnor U11617 (N_11617,N_7864,N_7804);
nor U11618 (N_11618,N_7800,N_8267);
nand U11619 (N_11619,N_8352,N_8724);
xnor U11620 (N_11620,N_7510,N_8273);
nor U11621 (N_11621,N_7711,N_9740);
or U11622 (N_11622,N_8001,N_9289);
nand U11623 (N_11623,N_8335,N_9589);
xnor U11624 (N_11624,N_8573,N_8807);
xnor U11625 (N_11625,N_7961,N_7512);
and U11626 (N_11626,N_7910,N_9852);
xnor U11627 (N_11627,N_8019,N_9173);
or U11628 (N_11628,N_7648,N_8541);
nand U11629 (N_11629,N_8608,N_7919);
nand U11630 (N_11630,N_7886,N_9242);
xor U11631 (N_11631,N_7785,N_9805);
or U11632 (N_11632,N_8674,N_8595);
or U11633 (N_11633,N_8648,N_8911);
or U11634 (N_11634,N_7830,N_7652);
nor U11635 (N_11635,N_7655,N_8281);
nand U11636 (N_11636,N_7906,N_8915);
nor U11637 (N_11637,N_8436,N_7602);
xor U11638 (N_11638,N_8503,N_8027);
nand U11639 (N_11639,N_7813,N_7852);
and U11640 (N_11640,N_9862,N_9888);
nor U11641 (N_11641,N_8351,N_9546);
or U11642 (N_11642,N_9443,N_7712);
nor U11643 (N_11643,N_8835,N_9639);
nand U11644 (N_11644,N_8749,N_9267);
nand U11645 (N_11645,N_7580,N_8868);
nand U11646 (N_11646,N_9137,N_8125);
xnor U11647 (N_11647,N_9302,N_7806);
nand U11648 (N_11648,N_9638,N_8116);
nand U11649 (N_11649,N_9229,N_8539);
or U11650 (N_11650,N_9470,N_8810);
or U11651 (N_11651,N_8758,N_8142);
xnor U11652 (N_11652,N_8074,N_9319);
nand U11653 (N_11653,N_8716,N_8635);
nand U11654 (N_11654,N_9049,N_9522);
xnor U11655 (N_11655,N_9619,N_8311);
xnor U11656 (N_11656,N_8796,N_8079);
and U11657 (N_11657,N_8441,N_9008);
nand U11658 (N_11658,N_7666,N_9883);
nor U11659 (N_11659,N_7834,N_9690);
nand U11660 (N_11660,N_9517,N_8890);
and U11661 (N_11661,N_9355,N_7749);
nand U11662 (N_11662,N_9220,N_8083);
nor U11663 (N_11663,N_7598,N_9507);
nand U11664 (N_11664,N_9138,N_8528);
or U11665 (N_11665,N_8365,N_8460);
or U11666 (N_11666,N_8435,N_7692);
nand U11667 (N_11667,N_7972,N_9234);
nor U11668 (N_11668,N_7665,N_9217);
and U11669 (N_11669,N_8139,N_9946);
nor U11670 (N_11670,N_9019,N_7876);
nand U11671 (N_11671,N_9526,N_7650);
nor U11672 (N_11672,N_9647,N_9552);
nor U11673 (N_11673,N_9847,N_8237);
nor U11674 (N_11674,N_9531,N_9248);
xor U11675 (N_11675,N_9740,N_9280);
or U11676 (N_11676,N_8852,N_8931);
nor U11677 (N_11677,N_9015,N_7692);
and U11678 (N_11678,N_8118,N_8246);
nand U11679 (N_11679,N_9922,N_9044);
and U11680 (N_11680,N_8909,N_7571);
or U11681 (N_11681,N_9043,N_9340);
nand U11682 (N_11682,N_9792,N_8587);
and U11683 (N_11683,N_7588,N_9186);
nand U11684 (N_11684,N_9737,N_7842);
nand U11685 (N_11685,N_7609,N_7794);
xor U11686 (N_11686,N_7529,N_7951);
xnor U11687 (N_11687,N_9980,N_7861);
nor U11688 (N_11688,N_9148,N_7896);
or U11689 (N_11689,N_9074,N_9864);
and U11690 (N_11690,N_8745,N_7602);
nor U11691 (N_11691,N_9257,N_8763);
xnor U11692 (N_11692,N_8266,N_9432);
and U11693 (N_11693,N_8615,N_9821);
xnor U11694 (N_11694,N_7832,N_8874);
xor U11695 (N_11695,N_9446,N_8869);
or U11696 (N_11696,N_9539,N_9845);
or U11697 (N_11697,N_7713,N_7852);
nor U11698 (N_11698,N_7685,N_7887);
nor U11699 (N_11699,N_7689,N_9295);
or U11700 (N_11700,N_8121,N_9655);
and U11701 (N_11701,N_9345,N_8078);
nor U11702 (N_11702,N_9022,N_9881);
and U11703 (N_11703,N_9028,N_8769);
and U11704 (N_11704,N_9732,N_8993);
xor U11705 (N_11705,N_7775,N_8244);
nand U11706 (N_11706,N_9110,N_8078);
xor U11707 (N_11707,N_9995,N_7537);
nor U11708 (N_11708,N_9958,N_7864);
nand U11709 (N_11709,N_8247,N_7553);
nor U11710 (N_11710,N_9247,N_8080);
nand U11711 (N_11711,N_8005,N_7789);
xor U11712 (N_11712,N_9508,N_9341);
xor U11713 (N_11713,N_9639,N_8485);
nor U11714 (N_11714,N_8611,N_8977);
and U11715 (N_11715,N_8438,N_9292);
nor U11716 (N_11716,N_8176,N_8094);
nand U11717 (N_11717,N_7869,N_9344);
xor U11718 (N_11718,N_9809,N_9849);
or U11719 (N_11719,N_8816,N_9149);
nor U11720 (N_11720,N_9587,N_9674);
and U11721 (N_11721,N_9367,N_8280);
nand U11722 (N_11722,N_8959,N_8086);
or U11723 (N_11723,N_9710,N_7642);
or U11724 (N_11724,N_7676,N_8995);
xnor U11725 (N_11725,N_8138,N_7971);
or U11726 (N_11726,N_8229,N_7600);
nand U11727 (N_11727,N_9579,N_9080);
or U11728 (N_11728,N_9608,N_9921);
nor U11729 (N_11729,N_8423,N_7893);
and U11730 (N_11730,N_8232,N_7534);
xor U11731 (N_11731,N_9110,N_8071);
nand U11732 (N_11732,N_9168,N_9594);
xnor U11733 (N_11733,N_8513,N_9276);
xnor U11734 (N_11734,N_9745,N_9995);
nor U11735 (N_11735,N_8500,N_7620);
xor U11736 (N_11736,N_8487,N_9980);
nand U11737 (N_11737,N_7636,N_7601);
nand U11738 (N_11738,N_8186,N_7786);
nor U11739 (N_11739,N_8569,N_9769);
and U11740 (N_11740,N_9382,N_8003);
xnor U11741 (N_11741,N_8205,N_8086);
and U11742 (N_11742,N_9628,N_9309);
and U11743 (N_11743,N_9507,N_8158);
nor U11744 (N_11744,N_8969,N_7886);
or U11745 (N_11745,N_8752,N_9915);
nor U11746 (N_11746,N_7945,N_8639);
xnor U11747 (N_11747,N_7778,N_7998);
xor U11748 (N_11748,N_9348,N_9926);
xor U11749 (N_11749,N_8069,N_8124);
xor U11750 (N_11750,N_8725,N_9171);
and U11751 (N_11751,N_9126,N_8468);
nand U11752 (N_11752,N_8209,N_7777);
or U11753 (N_11753,N_9446,N_7893);
xor U11754 (N_11754,N_8691,N_9616);
nor U11755 (N_11755,N_9635,N_9228);
nand U11756 (N_11756,N_8349,N_9196);
xnor U11757 (N_11757,N_9874,N_8108);
nor U11758 (N_11758,N_8554,N_9810);
nand U11759 (N_11759,N_8590,N_8947);
and U11760 (N_11760,N_7818,N_7648);
or U11761 (N_11761,N_9680,N_8322);
nor U11762 (N_11762,N_8440,N_9940);
nand U11763 (N_11763,N_8151,N_8602);
or U11764 (N_11764,N_9603,N_8865);
or U11765 (N_11765,N_8752,N_7798);
or U11766 (N_11766,N_9902,N_9250);
and U11767 (N_11767,N_8471,N_8563);
nor U11768 (N_11768,N_8969,N_8036);
nor U11769 (N_11769,N_9231,N_9820);
and U11770 (N_11770,N_7702,N_8210);
xnor U11771 (N_11771,N_8442,N_7831);
xnor U11772 (N_11772,N_9065,N_8817);
and U11773 (N_11773,N_8749,N_9094);
and U11774 (N_11774,N_8558,N_9325);
nor U11775 (N_11775,N_9794,N_9644);
nor U11776 (N_11776,N_9018,N_8804);
xnor U11777 (N_11777,N_7990,N_9750);
xnor U11778 (N_11778,N_8293,N_7798);
nand U11779 (N_11779,N_8992,N_8861);
nand U11780 (N_11780,N_9049,N_8664);
nand U11781 (N_11781,N_7658,N_8167);
nor U11782 (N_11782,N_8298,N_9120);
or U11783 (N_11783,N_8105,N_8859);
nand U11784 (N_11784,N_9562,N_8309);
or U11785 (N_11785,N_8149,N_8424);
xnor U11786 (N_11786,N_9435,N_8796);
nor U11787 (N_11787,N_9639,N_8694);
nor U11788 (N_11788,N_9195,N_7729);
nor U11789 (N_11789,N_9610,N_9633);
and U11790 (N_11790,N_7725,N_9730);
xor U11791 (N_11791,N_7596,N_8334);
or U11792 (N_11792,N_7650,N_8818);
xnor U11793 (N_11793,N_9766,N_8188);
nor U11794 (N_11794,N_8030,N_8417);
or U11795 (N_11795,N_7773,N_9118);
or U11796 (N_11796,N_9256,N_7621);
or U11797 (N_11797,N_8528,N_8386);
xor U11798 (N_11798,N_8512,N_8053);
nor U11799 (N_11799,N_9986,N_8588);
nor U11800 (N_11800,N_9273,N_9408);
xor U11801 (N_11801,N_8928,N_9515);
nand U11802 (N_11802,N_8064,N_9241);
xor U11803 (N_11803,N_8157,N_7875);
or U11804 (N_11804,N_8865,N_9175);
and U11805 (N_11805,N_8916,N_7861);
and U11806 (N_11806,N_8216,N_7706);
and U11807 (N_11807,N_8684,N_8757);
nand U11808 (N_11808,N_9874,N_8552);
and U11809 (N_11809,N_8931,N_9389);
and U11810 (N_11810,N_8623,N_7858);
nor U11811 (N_11811,N_9626,N_9741);
nor U11812 (N_11812,N_7929,N_9792);
xnor U11813 (N_11813,N_9376,N_8042);
or U11814 (N_11814,N_9274,N_8634);
xnor U11815 (N_11815,N_9772,N_9420);
nor U11816 (N_11816,N_9639,N_9308);
nor U11817 (N_11817,N_9262,N_9775);
nand U11818 (N_11818,N_8195,N_9486);
or U11819 (N_11819,N_8123,N_8348);
or U11820 (N_11820,N_8869,N_9445);
and U11821 (N_11821,N_9189,N_9632);
nor U11822 (N_11822,N_7673,N_9348);
or U11823 (N_11823,N_9491,N_7873);
or U11824 (N_11824,N_8828,N_9752);
nor U11825 (N_11825,N_7537,N_8844);
and U11826 (N_11826,N_8384,N_9672);
or U11827 (N_11827,N_8567,N_9422);
xnor U11828 (N_11828,N_7680,N_9157);
xnor U11829 (N_11829,N_9179,N_9168);
or U11830 (N_11830,N_9825,N_7502);
or U11831 (N_11831,N_9164,N_7817);
or U11832 (N_11832,N_8167,N_8320);
nor U11833 (N_11833,N_9703,N_8832);
or U11834 (N_11834,N_9238,N_9764);
xnor U11835 (N_11835,N_9254,N_8826);
xnor U11836 (N_11836,N_9235,N_9564);
or U11837 (N_11837,N_7722,N_8526);
or U11838 (N_11838,N_8185,N_9360);
nand U11839 (N_11839,N_8537,N_7999);
xor U11840 (N_11840,N_9789,N_7945);
nand U11841 (N_11841,N_8865,N_9616);
or U11842 (N_11842,N_8516,N_8685);
and U11843 (N_11843,N_7765,N_7744);
xor U11844 (N_11844,N_8755,N_9126);
xor U11845 (N_11845,N_9911,N_7788);
nand U11846 (N_11846,N_7594,N_8014);
or U11847 (N_11847,N_8935,N_8751);
nor U11848 (N_11848,N_9595,N_8495);
nor U11849 (N_11849,N_8529,N_8103);
or U11850 (N_11850,N_7981,N_9156);
and U11851 (N_11851,N_9839,N_8181);
xor U11852 (N_11852,N_9755,N_8839);
or U11853 (N_11853,N_7797,N_9618);
nand U11854 (N_11854,N_9191,N_8326);
nand U11855 (N_11855,N_8500,N_9602);
nor U11856 (N_11856,N_9719,N_8496);
or U11857 (N_11857,N_7828,N_9772);
xnor U11858 (N_11858,N_8371,N_7770);
and U11859 (N_11859,N_8438,N_9325);
nor U11860 (N_11860,N_9507,N_8550);
or U11861 (N_11861,N_7992,N_8804);
nor U11862 (N_11862,N_9558,N_8760);
or U11863 (N_11863,N_8824,N_7650);
xor U11864 (N_11864,N_7522,N_7845);
nor U11865 (N_11865,N_9223,N_7750);
and U11866 (N_11866,N_8039,N_9616);
nand U11867 (N_11867,N_9721,N_8148);
nor U11868 (N_11868,N_8031,N_7864);
or U11869 (N_11869,N_8088,N_9455);
or U11870 (N_11870,N_9643,N_9294);
and U11871 (N_11871,N_8963,N_9588);
and U11872 (N_11872,N_8657,N_9421);
or U11873 (N_11873,N_8287,N_9986);
nand U11874 (N_11874,N_9985,N_8217);
xnor U11875 (N_11875,N_8532,N_8334);
and U11876 (N_11876,N_9382,N_8444);
nor U11877 (N_11877,N_8543,N_9301);
or U11878 (N_11878,N_8269,N_8702);
and U11879 (N_11879,N_7825,N_8331);
nor U11880 (N_11880,N_9362,N_9554);
nand U11881 (N_11881,N_8352,N_8049);
xnor U11882 (N_11882,N_7906,N_9255);
xor U11883 (N_11883,N_7644,N_9078);
or U11884 (N_11884,N_7598,N_7640);
and U11885 (N_11885,N_7989,N_8235);
nor U11886 (N_11886,N_9738,N_7832);
xor U11887 (N_11887,N_7560,N_8506);
or U11888 (N_11888,N_9903,N_8545);
nor U11889 (N_11889,N_9477,N_9999);
or U11890 (N_11890,N_8496,N_7791);
nor U11891 (N_11891,N_7995,N_9242);
or U11892 (N_11892,N_9325,N_8924);
nor U11893 (N_11893,N_9545,N_9320);
nand U11894 (N_11894,N_9916,N_9265);
nand U11895 (N_11895,N_9709,N_8190);
or U11896 (N_11896,N_9508,N_8413);
or U11897 (N_11897,N_8381,N_9017);
xor U11898 (N_11898,N_8522,N_8380);
nand U11899 (N_11899,N_8589,N_9896);
and U11900 (N_11900,N_7610,N_8209);
xor U11901 (N_11901,N_7953,N_8397);
and U11902 (N_11902,N_9860,N_9650);
and U11903 (N_11903,N_8375,N_8792);
xnor U11904 (N_11904,N_8561,N_9093);
xnor U11905 (N_11905,N_7603,N_8854);
nor U11906 (N_11906,N_8720,N_8551);
nand U11907 (N_11907,N_8131,N_7735);
nand U11908 (N_11908,N_9282,N_9614);
xnor U11909 (N_11909,N_9995,N_9382);
xnor U11910 (N_11910,N_7886,N_9577);
and U11911 (N_11911,N_8243,N_7764);
or U11912 (N_11912,N_9121,N_8348);
and U11913 (N_11913,N_9814,N_9694);
and U11914 (N_11914,N_8798,N_7947);
nor U11915 (N_11915,N_7898,N_7917);
nand U11916 (N_11916,N_9077,N_9655);
nand U11917 (N_11917,N_9988,N_8392);
and U11918 (N_11918,N_9696,N_9988);
and U11919 (N_11919,N_9564,N_9321);
or U11920 (N_11920,N_9983,N_9621);
or U11921 (N_11921,N_9317,N_7750);
nor U11922 (N_11922,N_9014,N_8868);
nand U11923 (N_11923,N_9949,N_8469);
or U11924 (N_11924,N_9682,N_9417);
xnor U11925 (N_11925,N_8261,N_8029);
and U11926 (N_11926,N_8938,N_9914);
nand U11927 (N_11927,N_9991,N_7864);
nand U11928 (N_11928,N_8867,N_8096);
and U11929 (N_11929,N_7842,N_9779);
or U11930 (N_11930,N_7881,N_9784);
nand U11931 (N_11931,N_7728,N_9828);
and U11932 (N_11932,N_8663,N_9185);
and U11933 (N_11933,N_8399,N_9466);
or U11934 (N_11934,N_8297,N_8200);
and U11935 (N_11935,N_7915,N_9136);
xnor U11936 (N_11936,N_7949,N_8094);
xor U11937 (N_11937,N_8333,N_9231);
nor U11938 (N_11938,N_8625,N_9849);
or U11939 (N_11939,N_9411,N_9028);
xor U11940 (N_11940,N_9850,N_9853);
and U11941 (N_11941,N_9756,N_8208);
nor U11942 (N_11942,N_8049,N_8384);
or U11943 (N_11943,N_8741,N_9307);
xnor U11944 (N_11944,N_9726,N_7889);
or U11945 (N_11945,N_8800,N_7883);
or U11946 (N_11946,N_8071,N_9931);
nand U11947 (N_11947,N_8908,N_9958);
nand U11948 (N_11948,N_8425,N_9360);
nor U11949 (N_11949,N_9792,N_9644);
nand U11950 (N_11950,N_9801,N_9303);
or U11951 (N_11951,N_8333,N_8611);
xor U11952 (N_11952,N_8985,N_9720);
and U11953 (N_11953,N_9444,N_7976);
xnor U11954 (N_11954,N_7681,N_8624);
nor U11955 (N_11955,N_9542,N_8662);
and U11956 (N_11956,N_8870,N_8113);
nand U11957 (N_11957,N_7559,N_9091);
xnor U11958 (N_11958,N_9966,N_8510);
and U11959 (N_11959,N_7510,N_8316);
xor U11960 (N_11960,N_8242,N_8230);
and U11961 (N_11961,N_9208,N_7637);
and U11962 (N_11962,N_8067,N_9143);
xor U11963 (N_11963,N_9767,N_9041);
nand U11964 (N_11964,N_9630,N_9391);
and U11965 (N_11965,N_8962,N_9654);
xor U11966 (N_11966,N_9485,N_8289);
or U11967 (N_11967,N_9583,N_8504);
xnor U11968 (N_11968,N_8349,N_8981);
nand U11969 (N_11969,N_8840,N_9284);
or U11970 (N_11970,N_8815,N_7793);
xnor U11971 (N_11971,N_9608,N_8853);
nor U11972 (N_11972,N_9172,N_8808);
xor U11973 (N_11973,N_9731,N_8705);
xor U11974 (N_11974,N_8496,N_9042);
and U11975 (N_11975,N_9051,N_9562);
xor U11976 (N_11976,N_9851,N_8114);
and U11977 (N_11977,N_7710,N_7753);
and U11978 (N_11978,N_9064,N_8387);
xor U11979 (N_11979,N_8774,N_8268);
xor U11980 (N_11980,N_9424,N_8914);
and U11981 (N_11981,N_8091,N_9324);
nand U11982 (N_11982,N_8943,N_8874);
nor U11983 (N_11983,N_9197,N_9237);
and U11984 (N_11984,N_9437,N_8663);
and U11985 (N_11985,N_8048,N_9145);
and U11986 (N_11986,N_8473,N_7736);
xnor U11987 (N_11987,N_7907,N_9622);
and U11988 (N_11988,N_8712,N_9915);
nand U11989 (N_11989,N_8243,N_8452);
or U11990 (N_11990,N_8612,N_8965);
and U11991 (N_11991,N_7628,N_9615);
nand U11992 (N_11992,N_8219,N_9108);
or U11993 (N_11993,N_8607,N_7974);
nand U11994 (N_11994,N_9405,N_9919);
and U11995 (N_11995,N_9748,N_9979);
and U11996 (N_11996,N_9260,N_8145);
nand U11997 (N_11997,N_8559,N_7625);
nand U11998 (N_11998,N_9107,N_7634);
or U11999 (N_11999,N_8741,N_9295);
and U12000 (N_12000,N_9775,N_8048);
nor U12001 (N_12001,N_8350,N_8948);
nor U12002 (N_12002,N_9037,N_9859);
nand U12003 (N_12003,N_8608,N_8839);
xor U12004 (N_12004,N_7977,N_8597);
and U12005 (N_12005,N_8327,N_7922);
or U12006 (N_12006,N_9397,N_8599);
or U12007 (N_12007,N_8311,N_9167);
xnor U12008 (N_12008,N_7739,N_8273);
nand U12009 (N_12009,N_9448,N_7620);
and U12010 (N_12010,N_9913,N_7963);
nand U12011 (N_12011,N_8425,N_8186);
or U12012 (N_12012,N_8606,N_7556);
nor U12013 (N_12013,N_9943,N_8305);
xor U12014 (N_12014,N_8982,N_8384);
or U12015 (N_12015,N_7937,N_7655);
and U12016 (N_12016,N_9808,N_9997);
xnor U12017 (N_12017,N_8651,N_9593);
nor U12018 (N_12018,N_8174,N_8541);
nand U12019 (N_12019,N_9048,N_8019);
and U12020 (N_12020,N_9866,N_9426);
xor U12021 (N_12021,N_7717,N_7778);
nor U12022 (N_12022,N_9259,N_8505);
and U12023 (N_12023,N_8457,N_9437);
nor U12024 (N_12024,N_7555,N_9253);
and U12025 (N_12025,N_9704,N_9045);
and U12026 (N_12026,N_7843,N_8178);
nand U12027 (N_12027,N_8187,N_8149);
and U12028 (N_12028,N_7611,N_8506);
or U12029 (N_12029,N_8526,N_8886);
xor U12030 (N_12030,N_8366,N_8469);
xnor U12031 (N_12031,N_8472,N_8312);
and U12032 (N_12032,N_8934,N_9437);
and U12033 (N_12033,N_9680,N_8262);
and U12034 (N_12034,N_9954,N_9152);
nand U12035 (N_12035,N_7758,N_9988);
and U12036 (N_12036,N_7593,N_8626);
and U12037 (N_12037,N_9598,N_9097);
and U12038 (N_12038,N_9108,N_9826);
nor U12039 (N_12039,N_7723,N_7599);
or U12040 (N_12040,N_8481,N_9146);
and U12041 (N_12041,N_8263,N_9463);
xnor U12042 (N_12042,N_7973,N_8504);
nand U12043 (N_12043,N_8505,N_7995);
nand U12044 (N_12044,N_7589,N_8784);
nand U12045 (N_12045,N_8508,N_9300);
or U12046 (N_12046,N_8015,N_8380);
nand U12047 (N_12047,N_8872,N_9410);
or U12048 (N_12048,N_8465,N_8443);
xnor U12049 (N_12049,N_9207,N_7961);
nand U12050 (N_12050,N_9326,N_9987);
xor U12051 (N_12051,N_8850,N_8891);
nor U12052 (N_12052,N_8310,N_9011);
xnor U12053 (N_12053,N_8968,N_9754);
nor U12054 (N_12054,N_7824,N_8202);
nand U12055 (N_12055,N_8096,N_9377);
or U12056 (N_12056,N_8914,N_7688);
and U12057 (N_12057,N_9448,N_8681);
and U12058 (N_12058,N_8116,N_9973);
and U12059 (N_12059,N_9657,N_7674);
xnor U12060 (N_12060,N_9742,N_7684);
nand U12061 (N_12061,N_8121,N_8757);
xnor U12062 (N_12062,N_9848,N_8499);
or U12063 (N_12063,N_7799,N_8512);
or U12064 (N_12064,N_8893,N_8102);
nand U12065 (N_12065,N_8988,N_9003);
nor U12066 (N_12066,N_7772,N_8394);
and U12067 (N_12067,N_9497,N_9071);
nor U12068 (N_12068,N_8669,N_8295);
nor U12069 (N_12069,N_7954,N_8969);
or U12070 (N_12070,N_8606,N_8201);
and U12071 (N_12071,N_8332,N_9739);
nor U12072 (N_12072,N_7652,N_8106);
and U12073 (N_12073,N_8322,N_7652);
nand U12074 (N_12074,N_8503,N_8449);
and U12075 (N_12075,N_9986,N_8010);
or U12076 (N_12076,N_9566,N_9169);
nor U12077 (N_12077,N_9777,N_9812);
or U12078 (N_12078,N_8935,N_9526);
or U12079 (N_12079,N_8712,N_9356);
nor U12080 (N_12080,N_9937,N_9088);
nand U12081 (N_12081,N_8847,N_8864);
nor U12082 (N_12082,N_9158,N_9734);
nor U12083 (N_12083,N_9598,N_8785);
xor U12084 (N_12084,N_9256,N_7797);
or U12085 (N_12085,N_8587,N_9058);
xor U12086 (N_12086,N_7568,N_8030);
and U12087 (N_12087,N_9445,N_9366);
or U12088 (N_12088,N_7731,N_7831);
or U12089 (N_12089,N_7869,N_8084);
and U12090 (N_12090,N_9791,N_9032);
nand U12091 (N_12091,N_8232,N_9287);
and U12092 (N_12092,N_7682,N_9560);
xor U12093 (N_12093,N_9592,N_9248);
nand U12094 (N_12094,N_8623,N_8557);
nand U12095 (N_12095,N_7967,N_9069);
xnor U12096 (N_12096,N_8131,N_9138);
nor U12097 (N_12097,N_8781,N_9540);
and U12098 (N_12098,N_8208,N_9361);
nand U12099 (N_12099,N_9064,N_7807);
and U12100 (N_12100,N_7855,N_7629);
nand U12101 (N_12101,N_9774,N_9909);
and U12102 (N_12102,N_9982,N_7798);
and U12103 (N_12103,N_8225,N_8847);
nand U12104 (N_12104,N_8663,N_8761);
nand U12105 (N_12105,N_8807,N_9012);
nand U12106 (N_12106,N_8748,N_9655);
and U12107 (N_12107,N_9137,N_9341);
nor U12108 (N_12108,N_7893,N_8861);
or U12109 (N_12109,N_9446,N_7578);
xnor U12110 (N_12110,N_8797,N_9000);
nand U12111 (N_12111,N_8000,N_9709);
xor U12112 (N_12112,N_7564,N_8563);
xnor U12113 (N_12113,N_8266,N_9048);
nand U12114 (N_12114,N_7787,N_7799);
or U12115 (N_12115,N_7505,N_8054);
or U12116 (N_12116,N_9774,N_8310);
xnor U12117 (N_12117,N_9464,N_8930);
and U12118 (N_12118,N_9209,N_8380);
or U12119 (N_12119,N_8230,N_9195);
and U12120 (N_12120,N_8806,N_8010);
and U12121 (N_12121,N_8117,N_7677);
or U12122 (N_12122,N_9007,N_7544);
nand U12123 (N_12123,N_8399,N_9163);
nor U12124 (N_12124,N_9700,N_8127);
or U12125 (N_12125,N_8187,N_9629);
and U12126 (N_12126,N_9571,N_8248);
nor U12127 (N_12127,N_9064,N_8976);
xnor U12128 (N_12128,N_8065,N_7881);
nand U12129 (N_12129,N_9776,N_9849);
nor U12130 (N_12130,N_7645,N_8182);
xnor U12131 (N_12131,N_8602,N_7700);
and U12132 (N_12132,N_7770,N_8489);
nor U12133 (N_12133,N_9977,N_8779);
or U12134 (N_12134,N_9731,N_7553);
and U12135 (N_12135,N_8167,N_7838);
xnor U12136 (N_12136,N_9935,N_9319);
and U12137 (N_12137,N_9753,N_8344);
nand U12138 (N_12138,N_8924,N_9186);
and U12139 (N_12139,N_9078,N_9299);
and U12140 (N_12140,N_8537,N_9417);
nor U12141 (N_12141,N_9645,N_7531);
nor U12142 (N_12142,N_7951,N_8693);
nor U12143 (N_12143,N_8178,N_8890);
and U12144 (N_12144,N_8281,N_9909);
nand U12145 (N_12145,N_8485,N_9851);
and U12146 (N_12146,N_8739,N_9785);
nor U12147 (N_12147,N_8784,N_8217);
nand U12148 (N_12148,N_9957,N_9444);
nand U12149 (N_12149,N_7843,N_9195);
nor U12150 (N_12150,N_9649,N_9543);
or U12151 (N_12151,N_7963,N_8604);
or U12152 (N_12152,N_8089,N_8764);
or U12153 (N_12153,N_8239,N_8607);
nand U12154 (N_12154,N_9815,N_9601);
nand U12155 (N_12155,N_9161,N_8570);
xnor U12156 (N_12156,N_9324,N_7800);
nand U12157 (N_12157,N_8168,N_9499);
nand U12158 (N_12158,N_8407,N_8594);
or U12159 (N_12159,N_7692,N_8989);
nor U12160 (N_12160,N_9569,N_8250);
and U12161 (N_12161,N_8994,N_7627);
nor U12162 (N_12162,N_8671,N_9646);
nor U12163 (N_12163,N_8036,N_8776);
and U12164 (N_12164,N_8695,N_8775);
or U12165 (N_12165,N_8725,N_8475);
nand U12166 (N_12166,N_7549,N_8562);
xor U12167 (N_12167,N_7936,N_9321);
and U12168 (N_12168,N_9262,N_7590);
xnor U12169 (N_12169,N_9374,N_9143);
xor U12170 (N_12170,N_9069,N_7510);
nand U12171 (N_12171,N_9052,N_8444);
and U12172 (N_12172,N_9217,N_8957);
or U12173 (N_12173,N_7588,N_7886);
or U12174 (N_12174,N_8853,N_9831);
nand U12175 (N_12175,N_9104,N_9982);
xnor U12176 (N_12176,N_8055,N_8683);
or U12177 (N_12177,N_7877,N_8834);
nor U12178 (N_12178,N_7800,N_8683);
nand U12179 (N_12179,N_9792,N_9516);
nand U12180 (N_12180,N_9889,N_8270);
xnor U12181 (N_12181,N_9840,N_8329);
and U12182 (N_12182,N_8888,N_7646);
nand U12183 (N_12183,N_8750,N_8972);
or U12184 (N_12184,N_8354,N_9037);
nand U12185 (N_12185,N_9421,N_9468);
xor U12186 (N_12186,N_9300,N_8392);
or U12187 (N_12187,N_9626,N_9945);
and U12188 (N_12188,N_9697,N_8188);
and U12189 (N_12189,N_8097,N_9416);
or U12190 (N_12190,N_8443,N_8697);
or U12191 (N_12191,N_9075,N_9424);
nand U12192 (N_12192,N_9238,N_8027);
or U12193 (N_12193,N_8581,N_8977);
or U12194 (N_12194,N_8768,N_8237);
nand U12195 (N_12195,N_8816,N_8567);
nor U12196 (N_12196,N_7616,N_9519);
nor U12197 (N_12197,N_9474,N_7777);
and U12198 (N_12198,N_8814,N_8567);
or U12199 (N_12199,N_8065,N_8361);
or U12200 (N_12200,N_9214,N_8623);
nand U12201 (N_12201,N_7645,N_9468);
or U12202 (N_12202,N_8488,N_9802);
or U12203 (N_12203,N_9500,N_7815);
nor U12204 (N_12204,N_9436,N_8818);
xor U12205 (N_12205,N_8702,N_8986);
and U12206 (N_12206,N_8837,N_8715);
and U12207 (N_12207,N_8341,N_9298);
nor U12208 (N_12208,N_8219,N_7930);
or U12209 (N_12209,N_9299,N_8076);
xor U12210 (N_12210,N_8879,N_9697);
nor U12211 (N_12211,N_7760,N_7862);
or U12212 (N_12212,N_8142,N_8088);
nand U12213 (N_12213,N_7934,N_9711);
xor U12214 (N_12214,N_8057,N_8137);
or U12215 (N_12215,N_7570,N_8021);
xor U12216 (N_12216,N_9452,N_7886);
nand U12217 (N_12217,N_9251,N_9932);
nor U12218 (N_12218,N_8783,N_7803);
nor U12219 (N_12219,N_7969,N_8994);
nand U12220 (N_12220,N_9100,N_7927);
nand U12221 (N_12221,N_7774,N_9903);
xnor U12222 (N_12222,N_7634,N_8833);
and U12223 (N_12223,N_9715,N_8381);
and U12224 (N_12224,N_8870,N_7552);
nor U12225 (N_12225,N_8432,N_9795);
and U12226 (N_12226,N_9759,N_7568);
nand U12227 (N_12227,N_9036,N_7692);
nand U12228 (N_12228,N_8253,N_7628);
nand U12229 (N_12229,N_9795,N_9579);
nor U12230 (N_12230,N_8024,N_8722);
nor U12231 (N_12231,N_8449,N_8871);
and U12232 (N_12232,N_7753,N_8818);
and U12233 (N_12233,N_9025,N_9607);
nor U12234 (N_12234,N_8316,N_8078);
nand U12235 (N_12235,N_9464,N_8018);
or U12236 (N_12236,N_8844,N_9308);
and U12237 (N_12237,N_8917,N_9133);
or U12238 (N_12238,N_8050,N_9100);
nand U12239 (N_12239,N_9885,N_7639);
xnor U12240 (N_12240,N_7882,N_9279);
and U12241 (N_12241,N_8646,N_8029);
nor U12242 (N_12242,N_8665,N_8904);
nor U12243 (N_12243,N_8509,N_8529);
xor U12244 (N_12244,N_7549,N_8239);
nand U12245 (N_12245,N_7723,N_7692);
xor U12246 (N_12246,N_7583,N_8413);
nand U12247 (N_12247,N_7838,N_9356);
and U12248 (N_12248,N_9185,N_9118);
and U12249 (N_12249,N_8788,N_9095);
or U12250 (N_12250,N_7653,N_8927);
nand U12251 (N_12251,N_7529,N_7912);
or U12252 (N_12252,N_9094,N_9441);
nand U12253 (N_12253,N_9759,N_9871);
xor U12254 (N_12254,N_7505,N_9054);
or U12255 (N_12255,N_7965,N_9625);
xnor U12256 (N_12256,N_8079,N_9271);
or U12257 (N_12257,N_9572,N_8212);
nand U12258 (N_12258,N_9085,N_7682);
or U12259 (N_12259,N_8549,N_9049);
or U12260 (N_12260,N_9328,N_8150);
xor U12261 (N_12261,N_9837,N_8153);
nand U12262 (N_12262,N_9329,N_9672);
xnor U12263 (N_12263,N_9832,N_9786);
or U12264 (N_12264,N_7646,N_8738);
and U12265 (N_12265,N_9515,N_9811);
nand U12266 (N_12266,N_8164,N_9277);
xnor U12267 (N_12267,N_9111,N_7562);
or U12268 (N_12268,N_8011,N_9881);
xnor U12269 (N_12269,N_8617,N_8847);
nand U12270 (N_12270,N_9914,N_9304);
and U12271 (N_12271,N_7526,N_8516);
xor U12272 (N_12272,N_7723,N_8938);
xor U12273 (N_12273,N_7571,N_9626);
nor U12274 (N_12274,N_9338,N_8856);
nor U12275 (N_12275,N_9679,N_9235);
xor U12276 (N_12276,N_8585,N_8254);
nor U12277 (N_12277,N_9981,N_8737);
nor U12278 (N_12278,N_9480,N_8912);
nor U12279 (N_12279,N_8159,N_8608);
nor U12280 (N_12280,N_8085,N_7654);
and U12281 (N_12281,N_8556,N_9958);
nor U12282 (N_12282,N_8672,N_9822);
xnor U12283 (N_12283,N_8519,N_8257);
nand U12284 (N_12284,N_8181,N_8638);
and U12285 (N_12285,N_8840,N_9632);
and U12286 (N_12286,N_8793,N_8157);
and U12287 (N_12287,N_7557,N_7967);
and U12288 (N_12288,N_9683,N_9123);
or U12289 (N_12289,N_7675,N_7671);
nor U12290 (N_12290,N_8503,N_9584);
nand U12291 (N_12291,N_9433,N_9428);
nand U12292 (N_12292,N_9588,N_9364);
or U12293 (N_12293,N_9908,N_8179);
xnor U12294 (N_12294,N_9928,N_8418);
or U12295 (N_12295,N_9999,N_7548);
nand U12296 (N_12296,N_8555,N_8459);
nand U12297 (N_12297,N_8709,N_8956);
nand U12298 (N_12298,N_9092,N_9423);
and U12299 (N_12299,N_9226,N_9356);
and U12300 (N_12300,N_9353,N_8583);
nand U12301 (N_12301,N_9754,N_7828);
and U12302 (N_12302,N_8866,N_8255);
nor U12303 (N_12303,N_7945,N_9261);
or U12304 (N_12304,N_8257,N_9665);
xnor U12305 (N_12305,N_7677,N_9505);
nor U12306 (N_12306,N_8950,N_8677);
xnor U12307 (N_12307,N_8684,N_7817);
xor U12308 (N_12308,N_9413,N_9546);
and U12309 (N_12309,N_8916,N_7693);
nor U12310 (N_12310,N_9921,N_9190);
nor U12311 (N_12311,N_8615,N_7521);
nor U12312 (N_12312,N_7541,N_9919);
or U12313 (N_12313,N_8521,N_8905);
nand U12314 (N_12314,N_9390,N_9304);
and U12315 (N_12315,N_8195,N_9037);
xor U12316 (N_12316,N_9379,N_8538);
and U12317 (N_12317,N_9472,N_9998);
xor U12318 (N_12318,N_9387,N_8089);
nor U12319 (N_12319,N_9619,N_8705);
nor U12320 (N_12320,N_8337,N_7570);
nor U12321 (N_12321,N_7546,N_9555);
and U12322 (N_12322,N_9177,N_9726);
xnor U12323 (N_12323,N_8216,N_9505);
xor U12324 (N_12324,N_9841,N_8231);
or U12325 (N_12325,N_8397,N_9223);
xor U12326 (N_12326,N_7553,N_7791);
and U12327 (N_12327,N_9828,N_9866);
and U12328 (N_12328,N_9626,N_8771);
nor U12329 (N_12329,N_9979,N_9309);
nor U12330 (N_12330,N_9513,N_9303);
nor U12331 (N_12331,N_8870,N_8927);
or U12332 (N_12332,N_7748,N_9552);
nor U12333 (N_12333,N_9157,N_9972);
or U12334 (N_12334,N_9512,N_9086);
or U12335 (N_12335,N_7646,N_8617);
nand U12336 (N_12336,N_9348,N_9319);
nor U12337 (N_12337,N_8130,N_8213);
xnor U12338 (N_12338,N_7851,N_9966);
nand U12339 (N_12339,N_9740,N_9990);
xor U12340 (N_12340,N_7870,N_9874);
xor U12341 (N_12341,N_9214,N_7956);
or U12342 (N_12342,N_8259,N_9288);
xor U12343 (N_12343,N_9626,N_9174);
xnor U12344 (N_12344,N_7998,N_8412);
and U12345 (N_12345,N_9785,N_9826);
xnor U12346 (N_12346,N_8031,N_9849);
or U12347 (N_12347,N_8178,N_7623);
and U12348 (N_12348,N_9178,N_8328);
nand U12349 (N_12349,N_7819,N_8167);
nand U12350 (N_12350,N_9870,N_9499);
nand U12351 (N_12351,N_8276,N_8062);
and U12352 (N_12352,N_8081,N_8732);
nor U12353 (N_12353,N_9375,N_8801);
or U12354 (N_12354,N_8438,N_8923);
and U12355 (N_12355,N_7794,N_9790);
or U12356 (N_12356,N_8682,N_9127);
nor U12357 (N_12357,N_7981,N_9226);
nand U12358 (N_12358,N_9045,N_9878);
or U12359 (N_12359,N_9109,N_9786);
and U12360 (N_12360,N_8099,N_8393);
xnor U12361 (N_12361,N_7760,N_7764);
nor U12362 (N_12362,N_8051,N_9986);
xnor U12363 (N_12363,N_9648,N_8710);
and U12364 (N_12364,N_8898,N_8468);
xor U12365 (N_12365,N_9123,N_9380);
or U12366 (N_12366,N_8851,N_7936);
or U12367 (N_12367,N_9844,N_7901);
nor U12368 (N_12368,N_9464,N_9935);
and U12369 (N_12369,N_9811,N_9485);
xnor U12370 (N_12370,N_8369,N_7755);
and U12371 (N_12371,N_9440,N_9497);
xor U12372 (N_12372,N_8021,N_8702);
and U12373 (N_12373,N_8717,N_8435);
nand U12374 (N_12374,N_8902,N_8893);
and U12375 (N_12375,N_7551,N_8428);
nand U12376 (N_12376,N_9985,N_9577);
nor U12377 (N_12377,N_8900,N_9034);
or U12378 (N_12378,N_7586,N_9620);
xnor U12379 (N_12379,N_7959,N_9842);
or U12380 (N_12380,N_8200,N_8449);
xor U12381 (N_12381,N_9335,N_9364);
nand U12382 (N_12382,N_9386,N_9633);
xor U12383 (N_12383,N_8541,N_8027);
or U12384 (N_12384,N_9543,N_8148);
and U12385 (N_12385,N_9857,N_8280);
nand U12386 (N_12386,N_7640,N_8899);
and U12387 (N_12387,N_8868,N_7680);
nor U12388 (N_12388,N_7726,N_8966);
and U12389 (N_12389,N_8848,N_7561);
xor U12390 (N_12390,N_9373,N_9956);
or U12391 (N_12391,N_8753,N_9168);
and U12392 (N_12392,N_9028,N_8277);
nand U12393 (N_12393,N_8875,N_8309);
or U12394 (N_12394,N_7986,N_8495);
xor U12395 (N_12395,N_9569,N_8301);
nor U12396 (N_12396,N_9371,N_9528);
and U12397 (N_12397,N_8729,N_7962);
nand U12398 (N_12398,N_9107,N_8396);
xor U12399 (N_12399,N_7937,N_9222);
xor U12400 (N_12400,N_7828,N_8682);
xor U12401 (N_12401,N_8123,N_8030);
or U12402 (N_12402,N_9885,N_8759);
and U12403 (N_12403,N_8215,N_9492);
xnor U12404 (N_12404,N_8154,N_8363);
and U12405 (N_12405,N_8413,N_9041);
nand U12406 (N_12406,N_7919,N_8215);
and U12407 (N_12407,N_8852,N_7507);
xor U12408 (N_12408,N_8004,N_8813);
or U12409 (N_12409,N_8934,N_8438);
and U12410 (N_12410,N_8813,N_8166);
and U12411 (N_12411,N_9561,N_8081);
and U12412 (N_12412,N_9324,N_7774);
nor U12413 (N_12413,N_9108,N_7958);
and U12414 (N_12414,N_7626,N_8185);
xnor U12415 (N_12415,N_7539,N_9507);
nor U12416 (N_12416,N_8450,N_8400);
nor U12417 (N_12417,N_8157,N_9650);
nand U12418 (N_12418,N_8955,N_7535);
xnor U12419 (N_12419,N_8728,N_8007);
and U12420 (N_12420,N_8329,N_8658);
nand U12421 (N_12421,N_8557,N_9195);
or U12422 (N_12422,N_9584,N_8195);
xnor U12423 (N_12423,N_8088,N_9083);
or U12424 (N_12424,N_8349,N_7706);
or U12425 (N_12425,N_9535,N_8586);
or U12426 (N_12426,N_9167,N_9704);
xnor U12427 (N_12427,N_9365,N_9709);
xor U12428 (N_12428,N_8510,N_9679);
or U12429 (N_12429,N_9495,N_9923);
and U12430 (N_12430,N_9197,N_7941);
nor U12431 (N_12431,N_9327,N_8258);
and U12432 (N_12432,N_8365,N_8852);
nand U12433 (N_12433,N_9284,N_8691);
nand U12434 (N_12434,N_8561,N_8121);
nand U12435 (N_12435,N_9778,N_7720);
xnor U12436 (N_12436,N_8627,N_8966);
xnor U12437 (N_12437,N_8577,N_8560);
nor U12438 (N_12438,N_7847,N_9636);
or U12439 (N_12439,N_8766,N_9340);
nor U12440 (N_12440,N_9331,N_9474);
nand U12441 (N_12441,N_9598,N_8858);
or U12442 (N_12442,N_8443,N_7525);
nor U12443 (N_12443,N_8439,N_9533);
nand U12444 (N_12444,N_9277,N_9000);
nor U12445 (N_12445,N_8683,N_8285);
nand U12446 (N_12446,N_8969,N_9421);
nand U12447 (N_12447,N_8475,N_9824);
and U12448 (N_12448,N_9030,N_8176);
nand U12449 (N_12449,N_7707,N_9325);
nor U12450 (N_12450,N_9078,N_9192);
nor U12451 (N_12451,N_9892,N_9063);
and U12452 (N_12452,N_8779,N_9096);
and U12453 (N_12453,N_7740,N_8324);
nor U12454 (N_12454,N_7939,N_9953);
nand U12455 (N_12455,N_8560,N_9198);
nand U12456 (N_12456,N_8582,N_7557);
xor U12457 (N_12457,N_7803,N_8712);
or U12458 (N_12458,N_8408,N_8146);
nor U12459 (N_12459,N_7794,N_8017);
xnor U12460 (N_12460,N_7833,N_9936);
xnor U12461 (N_12461,N_7910,N_9623);
xnor U12462 (N_12462,N_8036,N_9727);
and U12463 (N_12463,N_8966,N_9500);
and U12464 (N_12464,N_8261,N_9743);
nor U12465 (N_12465,N_9794,N_9903);
nor U12466 (N_12466,N_7592,N_8207);
nor U12467 (N_12467,N_8814,N_9685);
nor U12468 (N_12468,N_7657,N_8744);
or U12469 (N_12469,N_7538,N_9881);
xor U12470 (N_12470,N_8774,N_8502);
or U12471 (N_12471,N_8576,N_9014);
nor U12472 (N_12472,N_7718,N_8641);
and U12473 (N_12473,N_8458,N_9955);
or U12474 (N_12474,N_8317,N_7528);
or U12475 (N_12475,N_8643,N_9528);
or U12476 (N_12476,N_9704,N_9925);
and U12477 (N_12477,N_7797,N_9372);
and U12478 (N_12478,N_7820,N_8874);
nand U12479 (N_12479,N_8593,N_9365);
nand U12480 (N_12480,N_9541,N_9851);
nand U12481 (N_12481,N_7664,N_9630);
nor U12482 (N_12482,N_8910,N_8823);
or U12483 (N_12483,N_7992,N_9473);
nor U12484 (N_12484,N_8601,N_9532);
or U12485 (N_12485,N_9714,N_9553);
nand U12486 (N_12486,N_9598,N_8501);
or U12487 (N_12487,N_8951,N_7755);
xor U12488 (N_12488,N_7552,N_9540);
or U12489 (N_12489,N_9820,N_7681);
and U12490 (N_12490,N_9015,N_7768);
or U12491 (N_12491,N_9441,N_9204);
and U12492 (N_12492,N_8855,N_9924);
nand U12493 (N_12493,N_9057,N_8566);
nand U12494 (N_12494,N_8603,N_8339);
nor U12495 (N_12495,N_7696,N_8939);
or U12496 (N_12496,N_7798,N_8993);
or U12497 (N_12497,N_7566,N_9726);
nand U12498 (N_12498,N_7964,N_8144);
nor U12499 (N_12499,N_8745,N_9847);
nand U12500 (N_12500,N_10875,N_11020);
and U12501 (N_12501,N_10809,N_10766);
nand U12502 (N_12502,N_12427,N_11326);
nor U12503 (N_12503,N_12200,N_11157);
and U12504 (N_12504,N_11409,N_12020);
or U12505 (N_12505,N_11072,N_12231);
or U12506 (N_12506,N_10366,N_11953);
nand U12507 (N_12507,N_11947,N_10682);
nor U12508 (N_12508,N_11758,N_10144);
and U12509 (N_12509,N_12292,N_11145);
or U12510 (N_12510,N_11795,N_11809);
nor U12511 (N_12511,N_11645,N_11931);
or U12512 (N_12512,N_11220,N_11411);
xnor U12513 (N_12513,N_11071,N_10876);
and U12514 (N_12514,N_10793,N_12018);
nand U12515 (N_12515,N_10727,N_11493);
xnor U12516 (N_12516,N_10327,N_10497);
nand U12517 (N_12517,N_12277,N_11537);
nor U12518 (N_12518,N_11100,N_10064);
nor U12519 (N_12519,N_10381,N_11987);
nor U12520 (N_12520,N_10192,N_10012);
nand U12521 (N_12521,N_10191,N_10000);
xnor U12522 (N_12522,N_10966,N_12269);
nand U12523 (N_12523,N_11381,N_11236);
xor U12524 (N_12524,N_11884,N_11569);
or U12525 (N_12525,N_10700,N_10758);
xnor U12526 (N_12526,N_11010,N_10959);
or U12527 (N_12527,N_11615,N_10313);
or U12528 (N_12528,N_11498,N_10276);
nand U12529 (N_12529,N_11548,N_11058);
nor U12530 (N_12530,N_11929,N_10351);
nand U12531 (N_12531,N_10475,N_10707);
and U12532 (N_12532,N_11367,N_11841);
nand U12533 (N_12533,N_11968,N_12023);
nor U12534 (N_12534,N_12214,N_11270);
and U12535 (N_12535,N_10223,N_10342);
nand U12536 (N_12536,N_11310,N_11408);
nand U12537 (N_12537,N_11515,N_11799);
nor U12538 (N_12538,N_10214,N_11040);
xnor U12539 (N_12539,N_12382,N_10234);
nor U12540 (N_12540,N_11756,N_10061);
and U12541 (N_12541,N_10914,N_12286);
nand U12542 (N_12542,N_11422,N_11227);
and U12543 (N_12543,N_12113,N_12156);
nor U12544 (N_12544,N_10826,N_10148);
or U12545 (N_12545,N_11583,N_12021);
xnor U12546 (N_12546,N_11845,N_11494);
or U12547 (N_12547,N_12332,N_11431);
or U12548 (N_12548,N_11142,N_12017);
xor U12549 (N_12549,N_10241,N_10404);
nor U12550 (N_12550,N_10640,N_11673);
nor U12551 (N_12551,N_11005,N_10883);
nor U12552 (N_12552,N_11840,N_10060);
nor U12553 (N_12553,N_11457,N_10090);
nor U12554 (N_12554,N_11394,N_10118);
nor U12555 (N_12555,N_10140,N_12187);
or U12556 (N_12556,N_11032,N_12417);
or U12557 (N_12557,N_10205,N_11539);
nand U12558 (N_12558,N_10812,N_11545);
nand U12559 (N_12559,N_10369,N_10474);
nand U12560 (N_12560,N_11991,N_12103);
nor U12561 (N_12561,N_11577,N_11327);
nand U12562 (N_12562,N_11347,N_10237);
or U12563 (N_12563,N_12080,N_10846);
nor U12564 (N_12564,N_10954,N_12275);
nand U12565 (N_12565,N_10498,N_11544);
nand U12566 (N_12566,N_10218,N_11380);
or U12567 (N_12567,N_10272,N_10273);
and U12568 (N_12568,N_11824,N_10601);
nand U12569 (N_12569,N_10481,N_12250);
nor U12570 (N_12570,N_12479,N_10508);
or U12571 (N_12571,N_12494,N_10319);
nand U12572 (N_12572,N_10861,N_10917);
and U12573 (N_12573,N_10282,N_11039);
nor U12574 (N_12574,N_10910,N_11303);
nand U12575 (N_12575,N_10949,N_10915);
nor U12576 (N_12576,N_11135,N_11774);
nor U12577 (N_12577,N_10219,N_11855);
and U12578 (N_12578,N_12499,N_11762);
nand U12579 (N_12579,N_10538,N_12480);
nor U12580 (N_12580,N_10080,N_11483);
and U12581 (N_12581,N_11649,N_11871);
nand U12582 (N_12582,N_11287,N_10533);
xor U12583 (N_12583,N_12320,N_11143);
and U12584 (N_12584,N_11585,N_11517);
xor U12585 (N_12585,N_10859,N_11410);
nand U12586 (N_12586,N_10057,N_10017);
and U12587 (N_12587,N_10027,N_12439);
nor U12588 (N_12588,N_11998,N_10583);
xor U12589 (N_12589,N_11301,N_10582);
xor U12590 (N_12590,N_11334,N_12450);
or U12591 (N_12591,N_12290,N_11125);
nor U12592 (N_12592,N_11885,N_10246);
nand U12593 (N_12593,N_11925,N_11509);
xor U12594 (N_12594,N_12291,N_10301);
xor U12595 (N_12595,N_10612,N_11862);
and U12596 (N_12596,N_10247,N_10195);
xnor U12597 (N_12597,N_10346,N_11580);
or U12598 (N_12598,N_12133,N_12318);
nor U12599 (N_12599,N_10131,N_10872);
or U12600 (N_12600,N_11798,N_11277);
and U12601 (N_12601,N_12339,N_12203);
nor U12602 (N_12602,N_12165,N_12322);
nor U12603 (N_12603,N_11056,N_11849);
nand U12604 (N_12604,N_12288,N_11065);
and U12605 (N_12605,N_10824,N_10604);
nor U12606 (N_12606,N_12466,N_11802);
or U12607 (N_12607,N_11672,N_10355);
nor U12608 (N_12608,N_11708,N_10922);
and U12609 (N_12609,N_11185,N_11190);
and U12610 (N_12610,N_12425,N_10098);
nor U12611 (N_12611,N_11678,N_11740);
or U12612 (N_12612,N_11863,N_10423);
nand U12613 (N_12613,N_12151,N_10592);
xor U12614 (N_12614,N_10322,N_10734);
nand U12615 (N_12615,N_11526,N_11838);
nor U12616 (N_12616,N_11946,N_10816);
nand U12617 (N_12617,N_10201,N_12493);
and U12618 (N_12618,N_12109,N_10843);
xor U12619 (N_12619,N_10735,N_12063);
or U12620 (N_12620,N_11400,N_10728);
xor U12621 (N_12621,N_10283,N_12378);
nor U12622 (N_12622,N_11727,N_10510);
nand U12623 (N_12623,N_10579,N_10285);
and U12624 (N_12624,N_12350,N_11842);
nand U12625 (N_12625,N_12002,N_11718);
nand U12626 (N_12626,N_11200,N_11426);
nor U12627 (N_12627,N_12311,N_11749);
xnor U12628 (N_12628,N_12010,N_10545);
or U12629 (N_12629,N_11386,N_10504);
nor U12630 (N_12630,N_11133,N_10725);
xor U12631 (N_12631,N_10746,N_10266);
or U12632 (N_12632,N_10400,N_11018);
xnor U12633 (N_12633,N_11805,N_10711);
nor U12634 (N_12634,N_10796,N_11612);
and U12635 (N_12635,N_11746,N_12126);
and U12636 (N_12636,N_10203,N_11048);
nand U12637 (N_12637,N_10033,N_11184);
or U12638 (N_12638,N_10432,N_12475);
or U12639 (N_12639,N_11358,N_11264);
nor U12640 (N_12640,N_11144,N_11835);
or U12641 (N_12641,N_10652,N_11331);
and U12642 (N_12642,N_11549,N_11123);
nor U12643 (N_12643,N_12428,N_10703);
and U12644 (N_12644,N_10335,N_12369);
xnor U12645 (N_12645,N_12478,N_11834);
or U12646 (N_12646,N_11922,N_10597);
and U12647 (N_12647,N_11487,N_11618);
or U12648 (N_12648,N_12278,N_10286);
and U12649 (N_12649,N_10975,N_10985);
xor U12650 (N_12650,N_11722,N_11937);
or U12651 (N_12651,N_12317,N_10124);
and U12652 (N_12652,N_10265,N_10523);
nor U12653 (N_12653,N_10401,N_12367);
nand U12654 (N_12654,N_11042,N_12408);
nand U12655 (N_12655,N_10557,N_11573);
and U12656 (N_12656,N_11883,N_11913);
nand U12657 (N_12657,N_11900,N_11706);
nand U12658 (N_12658,N_10558,N_10349);
or U12659 (N_12659,N_10116,N_11599);
nand U12660 (N_12660,N_11477,N_10486);
or U12661 (N_12661,N_10513,N_10564);
nor U12662 (N_12662,N_12089,N_11342);
nor U12663 (N_12663,N_12364,N_12303);
xnor U12664 (N_12664,N_11240,N_11423);
nor U12665 (N_12665,N_10713,N_11231);
and U12666 (N_12666,N_10186,N_10501);
nor U12667 (N_12667,N_10345,N_10316);
xor U12668 (N_12668,N_11479,N_11070);
nand U12669 (N_12669,N_10665,N_10536);
xnor U12670 (N_12670,N_11711,N_10795);
or U12671 (N_12671,N_12052,N_10947);
nand U12672 (N_12672,N_10177,N_10038);
or U12673 (N_12673,N_11503,N_12132);
or U12674 (N_12674,N_12391,N_11496);
and U12675 (N_12675,N_10965,N_10686);
or U12676 (N_12676,N_10183,N_12129);
nand U12677 (N_12677,N_10441,N_12462);
nor U12678 (N_12678,N_11779,N_10729);
xor U12679 (N_12679,N_12148,N_10855);
xor U12680 (N_12680,N_11606,N_10037);
nor U12681 (N_12681,N_10792,N_12430);
xor U12682 (N_12682,N_12333,N_12101);
and U12683 (N_12683,N_12449,N_10726);
nor U12684 (N_12684,N_11889,N_10906);
xor U12685 (N_12685,N_12219,N_11392);
or U12686 (N_12686,N_12009,N_12003);
and U12687 (N_12687,N_10047,N_10822);
nand U12688 (N_12688,N_11897,N_11516);
nor U12689 (N_12689,N_11547,N_11528);
or U12690 (N_12690,N_10547,N_10695);
nand U12691 (N_12691,N_10304,N_12223);
nor U12692 (N_12692,N_10373,N_11025);
xor U12693 (N_12693,N_10350,N_10014);
xnor U12694 (N_12694,N_11445,N_12040);
nor U12695 (N_12695,N_10937,N_11605);
nand U12696 (N_12696,N_12373,N_11519);
and U12697 (N_12697,N_10264,N_10073);
xnor U12698 (N_12698,N_10680,N_10270);
and U12699 (N_12699,N_11416,N_11560);
and U12700 (N_12700,N_11744,N_10377);
xor U12701 (N_12701,N_10065,N_10537);
or U12702 (N_12702,N_10907,N_12429);
and U12703 (N_12703,N_11846,N_10009);
nor U12704 (N_12704,N_10328,N_10337);
xor U12705 (N_12705,N_12065,N_12432);
or U12706 (N_12706,N_10111,N_10165);
xor U12707 (N_12707,N_12121,N_10622);
and U12708 (N_12708,N_10578,N_10823);
or U12709 (N_12709,N_12074,N_11215);
nand U12710 (N_12710,N_11245,N_10772);
or U12711 (N_12711,N_10455,N_12238);
nor U12712 (N_12712,N_11816,N_11211);
nand U12713 (N_12713,N_11266,N_11576);
nor U12714 (N_12714,N_10275,N_10397);
or U12715 (N_12715,N_10467,N_10150);
and U12716 (N_12716,N_10877,N_12446);
or U12717 (N_12717,N_10331,N_10129);
and U12718 (N_12718,N_11932,N_11844);
and U12719 (N_12719,N_12130,N_11401);
xor U12720 (N_12720,N_11113,N_10412);
nor U12721 (N_12721,N_11742,N_11149);
xor U12722 (N_12722,N_11260,N_11559);
nor U12723 (N_12723,N_12182,N_11873);
or U12724 (N_12724,N_10600,N_10834);
xor U12725 (N_12725,N_12049,N_11435);
and U12726 (N_12726,N_10175,N_10023);
xor U12727 (N_12727,N_11006,N_11434);
or U12728 (N_12728,N_12171,N_10243);
xor U12729 (N_12729,N_11867,N_11781);
xor U12730 (N_12730,N_11500,N_10114);
xnor U12731 (N_12731,N_12304,N_10565);
xor U12732 (N_12732,N_10574,N_10670);
nand U12733 (N_12733,N_10108,N_11087);
xor U12734 (N_12734,N_10886,N_12081);
nand U12735 (N_12735,N_11090,N_10022);
nand U12736 (N_12736,N_11963,N_11419);
xor U12737 (N_12737,N_12345,N_10245);
nor U12738 (N_12738,N_12416,N_12481);
or U12739 (N_12739,N_11354,N_10088);
or U12740 (N_12740,N_11948,N_10093);
and U12741 (N_12741,N_12376,N_10330);
nor U12742 (N_12742,N_10655,N_10015);
nand U12743 (N_12743,N_10961,N_11183);
and U12744 (N_12744,N_10338,N_11420);
nand U12745 (N_12745,N_12349,N_12053);
and U12746 (N_12746,N_10904,N_10030);
nand U12747 (N_12747,N_10839,N_11399);
nor U12748 (N_12748,N_10888,N_11692);
nor U12749 (N_12749,N_12325,N_12404);
nor U12750 (N_12750,N_10576,N_12107);
nor U12751 (N_12751,N_11768,N_10426);
nand U12752 (N_12752,N_10461,N_10387);
or U12753 (N_12753,N_12205,N_10661);
nand U12754 (N_12754,N_12346,N_10664);
nand U12755 (N_12755,N_10198,N_11022);
nor U12756 (N_12756,N_12385,N_10941);
or U12757 (N_12757,N_10468,N_10509);
or U12758 (N_12758,N_11255,N_11764);
or U12759 (N_12759,N_12088,N_10919);
or U12760 (N_12760,N_11314,N_11940);
nor U12761 (N_12761,N_11297,N_12239);
nor U12762 (N_12762,N_11712,N_10650);
or U12763 (N_12763,N_11012,N_11376);
or U12764 (N_12764,N_10935,N_10398);
or U12765 (N_12765,N_11872,N_12414);
nor U12766 (N_12766,N_12236,N_10732);
xnor U12767 (N_12767,N_12242,N_11892);
xnor U12768 (N_12768,N_11134,N_10499);
xnor U12769 (N_12769,N_10981,N_11075);
or U12770 (N_12770,N_10252,N_10067);
nand U12771 (N_12771,N_10750,N_12392);
xnor U12772 (N_12772,N_11624,N_11938);
and U12773 (N_12773,N_10411,N_11276);
xnor U12774 (N_12774,N_10303,N_12190);
or U12775 (N_12775,N_11592,N_11186);
and U12776 (N_12776,N_10176,N_11495);
or U12777 (N_12777,N_12183,N_10543);
or U12778 (N_12778,N_12123,N_10492);
nor U12779 (N_12779,N_11154,N_12038);
nand U12780 (N_12780,N_12441,N_11330);
nand U12781 (N_12781,N_12355,N_10759);
xnor U12782 (N_12782,N_11014,N_10999);
nand U12783 (N_12783,N_11904,N_10208);
and U12784 (N_12784,N_10464,N_10181);
or U12785 (N_12785,N_11957,N_10476);
nand U12786 (N_12786,N_12296,N_11620);
or U12787 (N_12787,N_11653,N_10858);
nor U12788 (N_12788,N_10893,N_11016);
or U12789 (N_12789,N_10251,N_10050);
and U12790 (N_12790,N_11783,N_11888);
nand U12791 (N_12791,N_11902,N_10326);
xnor U12792 (N_12792,N_11473,N_10287);
or U12793 (N_12793,N_11972,N_11374);
nor U12794 (N_12794,N_11403,N_11370);
nor U12795 (N_12795,N_10797,N_10605);
or U12796 (N_12796,N_11172,N_11981);
or U12797 (N_12797,N_10487,N_10048);
and U12798 (N_12798,N_11153,N_10573);
xnor U12799 (N_12799,N_11909,N_10016);
xor U12800 (N_12800,N_11136,N_11436);
nand U12801 (N_12801,N_12323,N_11046);
and U12802 (N_12802,N_10757,N_11782);
and U12803 (N_12803,N_11561,N_12356);
nor U12804 (N_12804,N_10415,N_12381);
nand U12805 (N_12805,N_11086,N_10780);
nand U12806 (N_12806,N_10347,N_11222);
xnor U12807 (N_12807,N_10257,N_11596);
xnor U12808 (N_12808,N_11833,N_11800);
nor U12809 (N_12809,N_12447,N_10168);
nand U12810 (N_12810,N_10685,N_11697);
or U12811 (N_12811,N_12188,N_12173);
nor U12812 (N_12812,N_11489,N_10736);
nor U12813 (N_12813,N_12402,N_12418);
or U12814 (N_12814,N_12154,N_10818);
nand U12815 (N_12815,N_11875,N_11466);
or U12816 (N_12816,N_10344,N_11613);
nand U12817 (N_12817,N_11621,N_11428);
xnor U12818 (N_12818,N_10639,N_11924);
and U12819 (N_12819,N_11208,N_12176);
or U12820 (N_12820,N_10672,N_10676);
xor U12821 (N_12821,N_11508,N_11979);
nand U12822 (N_12822,N_12093,N_11715);
nand U12823 (N_12823,N_12308,N_11066);
or U12824 (N_12824,N_11250,N_10298);
nor U12825 (N_12825,N_12166,N_10375);
and U12826 (N_12826,N_10233,N_12357);
and U12827 (N_12827,N_11322,N_11532);
nand U12828 (N_12828,N_11829,N_10830);
xor U12829 (N_12829,N_10866,N_10649);
or U12830 (N_12830,N_11175,N_10239);
nand U12831 (N_12831,N_10500,N_11108);
or U12832 (N_12832,N_10025,N_11572);
and U12833 (N_12833,N_10609,N_10182);
or U12834 (N_12834,N_12366,N_12315);
and U12835 (N_12835,N_11203,N_11146);
and U12836 (N_12836,N_10852,N_10913);
nand U12837 (N_12837,N_12281,N_11407);
nand U12838 (N_12838,N_11379,N_10180);
xnor U12839 (N_12839,N_10193,N_11660);
nand U12840 (N_12840,N_11602,N_11656);
or U12841 (N_12841,N_10840,N_11761);
xnor U12842 (N_12842,N_11017,N_11284);
nor U12843 (N_12843,N_11769,N_10516);
nor U12844 (N_12844,N_12117,N_11318);
and U12845 (N_12845,N_11556,N_11352);
nor U12846 (N_12846,N_12410,N_10028);
nand U12847 (N_12847,N_12160,N_11189);
nand U12848 (N_12848,N_11732,N_10952);
nor U12849 (N_12849,N_10076,N_10268);
nand U12850 (N_12850,N_11854,N_11249);
or U12851 (N_12851,N_10469,N_12082);
nor U12852 (N_12852,N_11982,N_11955);
or U12853 (N_12853,N_11766,N_11338);
and U12854 (N_12854,N_11648,N_10778);
xnor U12855 (N_12855,N_10152,N_10396);
or U12856 (N_12856,N_10248,N_11207);
nand U12857 (N_12857,N_10932,N_10737);
nand U12858 (N_12858,N_11634,N_10531);
and U12859 (N_12859,N_11346,N_10962);
nor U12860 (N_12860,N_11633,N_10043);
or U12861 (N_12861,N_10957,N_11751);
xor U12862 (N_12862,N_12263,N_10293);
nand U12863 (N_12863,N_10178,N_10606);
and U12864 (N_12864,N_11351,N_10608);
nand U12865 (N_12865,N_10951,N_12328);
nor U12866 (N_12866,N_10767,N_12487);
nor U12867 (N_12867,N_12058,N_11905);
or U12868 (N_12868,N_10221,N_11366);
or U12869 (N_12869,N_10160,N_10967);
or U12870 (N_12870,N_12229,N_10996);
xor U12871 (N_12871,N_11502,N_10333);
and U12872 (N_12872,N_10189,N_10353);
xor U12873 (N_12873,N_10081,N_12180);
or U12874 (N_12874,N_10306,N_10891);
nand U12875 (N_12875,N_10850,N_10388);
or U12876 (N_12876,N_10478,N_12247);
nand U12877 (N_12877,N_10137,N_10071);
and U12878 (N_12878,N_10315,N_10110);
xnor U12879 (N_12879,N_10164,N_12072);
nor U12880 (N_12880,N_12086,N_11879);
nor U12881 (N_12881,N_10117,N_12008);
nor U12882 (N_12882,N_11702,N_10153);
and U12883 (N_12883,N_11076,N_11213);
xor U12884 (N_12884,N_10414,N_10897);
nand U12885 (N_12885,N_10756,N_11669);
nor U12886 (N_12886,N_10638,N_11523);
nand U12887 (N_12887,N_11355,N_11527);
and U12888 (N_12888,N_11480,N_11522);
nand U12889 (N_12889,N_10515,N_11657);
nand U12890 (N_12890,N_10614,N_11206);
and U12891 (N_12891,N_11723,N_10420);
nor U12892 (N_12892,N_12039,N_11514);
or U12893 (N_12893,N_12098,N_10560);
nand U12894 (N_12894,N_11731,N_11343);
nand U12895 (N_12895,N_11155,N_10249);
or U12896 (N_12896,N_10278,N_12299);
and U12897 (N_12897,N_10462,N_10158);
nor U12898 (N_12898,N_10019,N_11292);
and U12899 (N_12899,N_12271,N_11725);
nor U12900 (N_12900,N_11964,N_10918);
xnor U12901 (N_12901,N_10628,N_12228);
nand U12902 (N_12902,N_10699,N_11666);
nand U12903 (N_12903,N_12193,N_10997);
and U12904 (N_12904,N_10280,N_11054);
or U12905 (N_12905,N_10648,N_12094);
and U12906 (N_12906,N_11173,N_11195);
nor U12907 (N_12907,N_10083,N_12297);
or U12908 (N_12908,N_10063,N_12025);
or U12909 (N_12909,N_10145,N_11546);
nor U12910 (N_12910,N_12454,N_11843);
nor U12911 (N_12911,N_11777,N_12336);
nand U12912 (N_12912,N_11893,N_11587);
and U12913 (N_12913,N_11233,N_10740);
xor U12914 (N_12914,N_11551,N_10066);
nor U12915 (N_12915,N_10289,N_11335);
nor U12916 (N_12916,N_10712,N_11707);
xor U12917 (N_12917,N_10225,N_11704);
nand U12918 (N_12918,N_11792,N_11741);
and U12919 (N_12919,N_10663,N_10806);
nor U12920 (N_12920,N_11939,N_10786);
and U12921 (N_12921,N_10151,N_10446);
nand U12922 (N_12922,N_11770,N_10385);
xnor U12923 (N_12923,N_12211,N_11404);
nand U12924 (N_12924,N_11755,N_10585);
xor U12925 (N_12925,N_11131,N_10115);
nand U12926 (N_12926,N_12007,N_11686);
nand U12927 (N_12927,N_10624,N_11282);
or U12928 (N_12928,N_11174,N_11047);
nor U12929 (N_12929,N_10697,N_12226);
nand U12930 (N_12930,N_10970,N_12386);
xnor U12931 (N_12931,N_11162,N_12334);
xor U12932 (N_12932,N_11699,N_11646);
nand U12933 (N_12933,N_10779,N_10004);
nand U12934 (N_12934,N_10358,N_11912);
xor U12935 (N_12935,N_11289,N_11041);
xor U12936 (N_12936,N_10617,N_10754);
or U12937 (N_12937,N_11438,N_11821);
and U12938 (N_12938,N_12326,N_10783);
or U12939 (N_12939,N_10323,N_10568);
nor U12940 (N_12940,N_10845,N_11541);
nand U12941 (N_12941,N_10184,N_11830);
xnor U12942 (N_12942,N_10236,N_10810);
xnor U12943 (N_12943,N_11138,N_12162);
nor U12944 (N_12944,N_12348,N_10172);
and U12945 (N_12945,N_10425,N_11970);
or U12946 (N_12946,N_10626,N_10125);
and U12947 (N_12947,N_10107,N_11994);
nor U12948 (N_12948,N_10804,N_11876);
xnor U12949 (N_12949,N_11349,N_12419);
or U12950 (N_12950,N_12144,N_10041);
and U12951 (N_12951,N_10130,N_10173);
or U12952 (N_12952,N_10698,N_10119);
and U12953 (N_12953,N_10905,N_11652);
xor U12954 (N_12954,N_10668,N_11474);
and U12955 (N_12955,N_11302,N_10874);
or U12956 (N_12956,N_11117,N_10132);
xnor U12957 (N_12957,N_11864,N_12174);
xor U12958 (N_12958,N_10794,N_10517);
nor U12959 (N_12959,N_12091,N_11446);
and U12960 (N_12960,N_10819,N_12116);
nor U12961 (N_12961,N_10798,N_12393);
or U12962 (N_12962,N_11116,N_10157);
and U12963 (N_12963,N_11898,N_12106);
and U12964 (N_12964,N_11826,N_10994);
or U12965 (N_12965,N_12302,N_10895);
or U12966 (N_12966,N_11499,N_10473);
nand U12967 (N_12967,N_11760,N_10109);
nor U12968 (N_12968,N_12233,N_10992);
nand U12969 (N_12969,N_12396,N_10973);
xor U12970 (N_12970,N_10419,N_12047);
nand U12971 (N_12971,N_11819,N_11927);
nand U12972 (N_12972,N_12014,N_10702);
and U12973 (N_12973,N_11817,N_11837);
nor U12974 (N_12974,N_10062,N_10052);
or U12975 (N_12975,N_10853,N_12057);
or U12976 (N_12976,N_12273,N_10405);
xor U12977 (N_12977,N_11969,N_10141);
nor U12978 (N_12978,N_10360,N_11388);
and U12979 (N_12979,N_11714,N_12309);
xnor U12980 (N_12980,N_10296,N_10427);
and U12981 (N_12981,N_11315,N_10921);
nor U12982 (N_12982,N_12136,N_11941);
and U12983 (N_12983,N_10869,N_11470);
or U12984 (N_12984,N_11166,N_10693);
nor U12985 (N_12985,N_11443,N_11321);
and U12986 (N_12986,N_12212,N_12464);
nand U12987 (N_12987,N_11150,N_10135);
and U12988 (N_12988,N_11415,N_10690);
nand U12989 (N_12989,N_10911,N_11990);
and U12990 (N_12990,N_12360,N_10596);
xnor U12991 (N_12991,N_11936,N_11579);
nand U12992 (N_12992,N_12383,N_11642);
and U12993 (N_12993,N_12352,N_10710);
and U12994 (N_12994,N_11716,N_11050);
nor U12995 (N_12995,N_12342,N_11414);
and U12996 (N_12996,N_10969,N_10363);
xor U12997 (N_12997,N_11540,N_11110);
nor U12998 (N_12998,N_11348,N_11647);
nor U12999 (N_12999,N_10607,N_11801);
nor U13000 (N_13000,N_10374,N_11793);
xnor U13001 (N_13001,N_11632,N_11308);
nor U13002 (N_13002,N_12240,N_10217);
or U13003 (N_13003,N_11198,N_11061);
nand U13004 (N_13004,N_11429,N_11051);
and U13005 (N_13005,N_11784,N_10613);
or U13006 (N_13006,N_10658,N_12120);
nor U13007 (N_13007,N_10674,N_11610);
or U13008 (N_13008,N_10989,N_11160);
nand U13009 (N_13009,N_10955,N_10202);
or U13010 (N_13010,N_10139,N_11341);
nand U13011 (N_13011,N_12471,N_11794);
xnor U13012 (N_13012,N_10307,N_11325);
nand U13013 (N_13013,N_11424,N_12215);
xor U13014 (N_13014,N_11966,N_10378);
xor U13015 (N_13015,N_11199,N_11091);
nor U13016 (N_13016,N_11575,N_11031);
or U13017 (N_13017,N_12145,N_11235);
and U13018 (N_13018,N_12175,N_10087);
nor U13019 (N_13019,N_12260,N_11853);
or U13020 (N_13020,N_10944,N_12122);
and U13021 (N_13021,N_11717,N_12407);
nand U13022 (N_13022,N_11158,N_10762);
nor U13023 (N_13023,N_11440,N_11775);
nand U13024 (N_13024,N_10292,N_12184);
xor U13025 (N_13025,N_10552,N_11996);
nand U13026 (N_13026,N_11385,N_10773);
and U13027 (N_13027,N_10867,N_11976);
xnor U13028 (N_13028,N_11590,N_11695);
or U13029 (N_13029,N_12244,N_10774);
or U13030 (N_13030,N_11719,N_10256);
and U13031 (N_13031,N_10817,N_10005);
xnor U13032 (N_13032,N_12489,N_10422);
nand U13033 (N_13033,N_10657,N_10320);
or U13034 (N_13034,N_10185,N_10739);
nand U13035 (N_13035,N_10259,N_11002);
nand U13036 (N_13036,N_10044,N_10653);
nand U13037 (N_13037,N_10733,N_12488);
xor U13038 (N_13038,N_10436,N_11747);
nand U13039 (N_13039,N_10782,N_10741);
nand U13040 (N_13040,N_12405,N_10644);
xor U13041 (N_13041,N_11192,N_10084);
nand U13042 (N_13042,N_10654,N_11670);
nand U13043 (N_13043,N_12201,N_11391);
nor U13044 (N_13044,N_11811,N_12451);
and U13045 (N_13045,N_12256,N_11813);
xor U13046 (N_13046,N_12327,N_10829);
nor U13047 (N_13047,N_10242,N_10988);
or U13048 (N_13048,N_10370,N_10069);
or U13049 (N_13049,N_12210,N_10007);
and U13050 (N_13050,N_12064,N_12196);
nand U13051 (N_13051,N_11677,N_11743);
nand U13052 (N_13052,N_12437,N_10925);
nor U13053 (N_13053,N_10563,N_11271);
or U13054 (N_13054,N_10408,N_11977);
nand U13055 (N_13055,N_12426,N_12310);
and U13056 (N_13056,N_10983,N_12090);
xnor U13057 (N_13057,N_11180,N_10121);
nand U13058 (N_13058,N_12143,N_12150);
nand U13059 (N_13059,N_11458,N_10162);
nor U13060 (N_13060,N_12141,N_10334);
and U13061 (N_13061,N_10254,N_12261);
or U13062 (N_13062,N_10570,N_11974);
xnor U13063 (N_13063,N_11038,N_11194);
nor U13064 (N_13064,N_12246,N_11242);
nand U13065 (N_13065,N_11759,N_10161);
or U13066 (N_13066,N_10465,N_10010);
nor U13067 (N_13067,N_11787,N_12139);
or U13068 (N_13068,N_11983,N_11468);
xor U13069 (N_13069,N_10228,N_10482);
nand U13070 (N_13070,N_10407,N_12252);
and U13071 (N_13071,N_10321,N_10493);
xor U13072 (N_13072,N_10399,N_11027);
or U13073 (N_13073,N_10356,N_10719);
xor U13074 (N_13074,N_10085,N_12204);
xor U13075 (N_13075,N_10212,N_10046);
nand U13076 (N_13076,N_10837,N_11689);
nor U13077 (N_13077,N_10445,N_10953);
nor U13078 (N_13078,N_10011,N_11878);
or U13079 (N_13079,N_11643,N_12397);
nand U13080 (N_13080,N_11665,N_11965);
nand U13081 (N_13081,N_10878,N_11788);
xor U13082 (N_13082,N_11170,N_11141);
nand U13083 (N_13083,N_10382,N_10379);
xor U13084 (N_13084,N_11895,N_10987);
nand U13085 (N_13085,N_12061,N_12026);
and U13086 (N_13086,N_12216,N_12467);
nor U13087 (N_13087,N_11600,N_10194);
and U13088 (N_13088,N_10442,N_10112);
nand U13089 (N_13089,N_10452,N_11030);
nand U13090 (N_13090,N_10684,N_10752);
xnor U13091 (N_13091,N_10260,N_10662);
or U13092 (N_13092,N_11390,N_10744);
nand U13093 (N_13093,N_10021,N_11928);
nor U13094 (N_13094,N_11096,N_10179);
or U13095 (N_13095,N_12012,N_10155);
or U13096 (N_13096,N_11914,N_12055);
nor U13097 (N_13097,N_11193,N_10295);
or U13098 (N_13098,N_11683,N_10637);
nand U13099 (N_13099,N_11626,N_10660);
xor U13100 (N_13100,N_10364,N_10495);
or U13101 (N_13101,N_10091,N_11832);
nand U13102 (N_13102,N_11852,N_11839);
nor U13103 (N_13103,N_11300,N_10651);
and U13104 (N_13104,N_12490,N_12465);
xnor U13105 (N_13105,N_11106,N_10784);
or U13106 (N_13106,N_12368,N_11115);
xor U13107 (N_13107,N_10924,N_10569);
and U13108 (N_13108,N_11533,N_12243);
nor U13109 (N_13109,N_11283,N_12084);
nand U13110 (N_13110,N_10235,N_12387);
nor U13111 (N_13111,N_12284,N_10631);
and U13112 (N_13112,N_11316,N_11412);
and U13113 (N_13113,N_11671,N_10209);
and U13114 (N_13114,N_10594,N_11951);
or U13115 (N_13115,N_12198,N_12206);
or U13116 (N_13116,N_12147,N_12491);
xor U13117 (N_13117,N_10636,N_10300);
xor U13118 (N_13118,N_11272,N_11786);
and U13119 (N_13119,N_12045,N_10122);
nand U13120 (N_13120,N_10956,N_11890);
xnor U13121 (N_13121,N_10716,N_12324);
xnor U13122 (N_13122,N_12372,N_12423);
or U13123 (N_13123,N_10018,N_10760);
or U13124 (N_13124,N_12329,N_10365);
nand U13125 (N_13125,N_10521,N_10930);
and U13126 (N_13126,N_11304,N_10444);
and U13127 (N_13127,N_11950,N_11542);
xnor U13128 (N_13128,N_11285,N_12431);
xnor U13129 (N_13129,N_11393,N_10789);
nor U13130 (N_13130,N_10311,N_12000);
or U13131 (N_13131,N_10329,N_12067);
xnor U13132 (N_13132,N_10715,N_10200);
nor U13133 (N_13133,N_11525,N_10416);
nand U13134 (N_13134,N_11628,N_12313);
or U13135 (N_13135,N_11406,N_11015);
and U13136 (N_13136,N_11934,N_11586);
and U13137 (N_13137,N_10409,N_11033);
xnor U13138 (N_13138,N_10484,N_12168);
or U13139 (N_13139,N_12118,N_11244);
or U13140 (N_13140,N_11497,N_10820);
nand U13141 (N_13141,N_10936,N_11161);
nand U13142 (N_13142,N_10646,N_11942);
or U13143 (N_13143,N_12066,N_10768);
and U13144 (N_13144,N_11880,N_12316);
and U13145 (N_13145,N_11168,N_12413);
xor U13146 (N_13146,N_12270,N_12172);
nor U13147 (N_13147,N_10494,N_10808);
or U13148 (N_13148,N_10838,N_11202);
and U13149 (N_13149,N_12495,N_11044);
nor U13150 (N_13150,N_10053,N_10566);
nor U13151 (N_13151,N_12400,N_11209);
nand U13152 (N_13152,N_12295,N_11815);
nand U13153 (N_13153,N_12482,N_10553);
or U13154 (N_13154,N_10979,N_10525);
nand U13155 (N_13155,N_10472,N_12114);
xnor U13156 (N_13156,N_12477,N_10731);
nand U13157 (N_13157,N_12249,N_11881);
nor U13158 (N_13158,N_11109,N_10174);
and U13159 (N_13159,N_11814,N_11013);
and U13160 (N_13160,N_11631,N_12254);
and U13161 (N_13161,N_11954,N_12164);
or U13162 (N_13162,N_11187,N_10391);
or U13163 (N_13163,N_11651,N_10687);
or U13164 (N_13164,N_12266,N_10673);
nand U13165 (N_13165,N_12004,N_11372);
nand U13166 (N_13166,N_12330,N_12044);
and U13167 (N_13167,N_11114,N_10706);
nand U13168 (N_13168,N_11906,N_11789);
nor U13169 (N_13169,N_11074,N_12051);
and U13170 (N_13170,N_11822,N_11089);
or U13171 (N_13171,N_10916,N_11685);
xnor U13172 (N_13172,N_12022,N_10502);
nand U13173 (N_13173,N_12068,N_12030);
or U13174 (N_13174,N_10410,N_11810);
and U13175 (N_13175,N_10434,N_10453);
and U13176 (N_13176,N_10395,N_10045);
or U13177 (N_13177,N_11856,N_12124);
nand U13178 (N_13178,N_10724,N_12158);
or U13179 (N_13179,N_10632,N_10036);
xor U13180 (N_13180,N_10960,N_11147);
and U13181 (N_13181,N_10099,N_11679);
nor U13182 (N_13182,N_12054,N_10584);
xnor U13183 (N_13183,N_12128,N_10072);
or U13184 (N_13184,N_10933,N_10633);
and U13185 (N_13185,N_11510,N_11578);
nand U13186 (N_13186,N_11619,N_10032);
nand U13187 (N_13187,N_11223,N_10642);
and U13188 (N_13188,N_10908,N_10227);
or U13189 (N_13189,N_10357,N_11636);
and U13190 (N_13190,N_10421,N_12420);
nor U13191 (N_13191,N_11910,N_11165);
nand U13192 (N_13192,N_11312,N_10244);
or U13193 (N_13193,N_12048,N_10535);
nor U13194 (N_13194,N_12340,N_11505);
and U13195 (N_13195,N_11562,N_12347);
nand U13196 (N_13196,N_10394,N_11230);
and U13197 (N_13197,N_10892,N_10898);
xor U13198 (N_13198,N_11735,N_10920);
or U13199 (N_13199,N_11060,N_12031);
xor U13200 (N_13200,N_10743,N_11377);
nand U13201 (N_13201,N_10075,N_11437);
nand U13202 (N_13202,N_12337,N_11239);
nand U13203 (N_13203,N_12379,N_11069);
and U13204 (N_13204,N_10599,N_11566);
or U13205 (N_13205,N_10871,N_12056);
nor U13206 (N_13206,N_10447,N_11265);
or U13207 (N_13207,N_12422,N_11857);
nand U13208 (N_13208,N_10042,N_11305);
nor U13209 (N_13209,N_10591,N_10993);
nand U13210 (N_13210,N_10156,N_11923);
and U13211 (N_13211,N_11122,N_10341);
and U13212 (N_13212,N_11080,N_11248);
or U13213 (N_13213,N_12388,N_10332);
and U13214 (N_13214,N_11796,N_10645);
and U13215 (N_13215,N_10831,N_11703);
xor U13216 (N_13216,N_11320,N_11674);
xor U13217 (N_13217,N_10294,N_12403);
or U13218 (N_13218,N_11188,N_11099);
and U13219 (N_13219,N_10368,N_11571);
nand U13220 (N_13220,N_12276,N_10903);
and U13221 (N_13221,N_10466,N_10863);
or U13222 (N_13222,N_12354,N_11105);
xnor U13223 (N_13223,N_10980,N_10581);
and U13224 (N_13224,N_11698,N_11294);
xor U13225 (N_13225,N_11684,N_10149);
nand U13226 (N_13226,N_10429,N_11280);
nand U13227 (N_13227,N_10790,N_11772);
or U13228 (N_13228,N_10143,N_10745);
xnor U13229 (N_13229,N_10216,N_10889);
nor U13230 (N_13230,N_12208,N_10939);
nor U13231 (N_13231,N_10196,N_11163);
or U13232 (N_13232,N_10616,N_11943);
or U13233 (N_13233,N_11861,N_11073);
and U13234 (N_13234,N_10480,N_11917);
and U13235 (N_13235,N_10559,N_10958);
xnor U13236 (N_13236,N_11364,N_10586);
nand U13237 (N_13237,N_10103,N_10821);
nor U13238 (N_13238,N_11252,N_11550);
nand U13239 (N_13239,N_10231,N_10708);
and U13240 (N_13240,N_10546,N_10479);
and U13241 (N_13241,N_10675,N_11622);
nand U13242 (N_13242,N_10755,N_11095);
or U13243 (N_13243,N_10721,N_10984);
xor U13244 (N_13244,N_12338,N_10856);
and U13245 (N_13245,N_11687,N_12301);
nand U13246 (N_13246,N_10857,N_11353);
xor U13247 (N_13247,N_10738,N_12095);
nand U13248 (N_13248,N_12362,N_10833);
nand U13249 (N_13249,N_11034,N_10006);
xor U13250 (N_13250,N_11247,N_11675);
xnor U13251 (N_13251,N_11396,N_11476);
and U13252 (N_13252,N_12234,N_11780);
xor U13253 (N_13253,N_11710,N_11063);
xnor U13254 (N_13254,N_11345,N_12016);
nand U13255 (N_13255,N_12496,N_10380);
or U13256 (N_13256,N_11971,N_11298);
nand U13257 (N_13257,N_12059,N_10456);
nand U13258 (N_13258,N_12374,N_11081);
nor U13259 (N_13259,N_11908,N_10376);
nand U13260 (N_13260,N_12006,N_10602);
xnor U13261 (N_13261,N_11274,N_10625);
nor U13262 (N_13262,N_12140,N_10880);
nand U13263 (N_13263,N_11915,N_11229);
or U13264 (N_13264,N_10439,N_11529);
nor U13265 (N_13265,N_10146,N_11765);
nand U13266 (N_13266,N_11439,N_11616);
nand U13267 (N_13267,N_10056,N_11009);
or U13268 (N_13268,N_10873,N_12282);
nor U13269 (N_13269,N_12458,N_12389);
or U13270 (N_13270,N_10828,N_12060);
or U13271 (N_13271,N_11043,N_11068);
xor U13272 (N_13272,N_10555,N_10528);
nand U13273 (N_13273,N_11644,N_12321);
xor U13274 (N_13274,N_11471,N_11721);
or U13275 (N_13275,N_11989,N_11427);
xor U13276 (N_13276,N_11945,N_11269);
and U13277 (N_13277,N_12375,N_11557);
nand U13278 (N_13278,N_12033,N_11241);
and U13279 (N_13279,N_11232,N_12001);
nor U13280 (N_13280,N_10159,N_12440);
and U13281 (N_13281,N_11375,N_10490);
nor U13282 (N_13282,N_12245,N_11603);
and U13283 (N_13283,N_10197,N_10931);
or U13284 (N_13284,N_11421,N_12137);
nor U13285 (N_13285,N_12062,N_11639);
xnor U13286 (N_13286,N_11911,N_10912);
and U13287 (N_13287,N_11340,N_11752);
and U13288 (N_13288,N_10595,N_12102);
nand U13289 (N_13289,N_10058,N_12335);
and U13290 (N_13290,N_10643,N_10832);
nor U13291 (N_13291,N_11465,N_10865);
or U13292 (N_13292,N_11739,N_10730);
or U13293 (N_13293,N_10704,N_11894);
or U13294 (N_13294,N_12161,N_12073);
or U13295 (N_13295,N_10694,N_10503);
nand U13296 (N_13296,N_10440,N_10222);
xnor U13297 (N_13297,N_10210,N_10974);
nor U13298 (N_13298,N_12486,N_10305);
or U13299 (N_13299,N_10105,N_10238);
nand U13300 (N_13300,N_11064,N_11901);
or U13301 (N_13301,N_11097,N_10879);
and U13302 (N_13302,N_11467,N_11273);
or U13303 (N_13303,N_11003,N_12306);
nor U13304 (N_13304,N_11754,N_11638);
or U13305 (N_13305,N_10054,N_10938);
nand U13306 (N_13306,N_12476,N_11368);
xor U13307 (N_13307,N_10133,N_10457);
and U13308 (N_13308,N_12222,N_10598);
nor U13309 (N_13309,N_12268,N_10909);
nor U13310 (N_13310,N_12153,N_11167);
or U13311 (N_13311,N_12119,N_11588);
and U13312 (N_13312,N_11103,N_10520);
and U13313 (N_13313,N_12461,N_12037);
or U13314 (N_13314,N_12181,N_10534);
xor U13315 (N_13315,N_11311,N_10449);
nor U13316 (N_13316,N_11625,N_11151);
and U13317 (N_13317,N_10352,N_11129);
xnor U13318 (N_13318,N_11828,N_10881);
nand U13319 (N_13319,N_12015,N_11313);
nand U13320 (N_13320,N_12406,N_11214);
and U13321 (N_13321,N_10113,N_10868);
xnor U13322 (N_13322,N_10611,N_11738);
and U13323 (N_13323,N_10163,N_12146);
nor U13324 (N_13324,N_10518,N_11567);
nor U13325 (N_13325,N_10963,N_10929);
nand U13326 (N_13326,N_11112,N_10890);
nor U13327 (N_13327,N_12359,N_10785);
nor U13328 (N_13328,N_10031,N_10188);
and U13329 (N_13329,N_10001,N_10751);
or U13330 (N_13330,N_11728,N_11958);
xor U13331 (N_13331,N_12170,N_12071);
or U13332 (N_13332,N_11797,N_10170);
or U13333 (N_13333,N_11682,N_10864);
or U13334 (N_13334,N_12399,N_11425);
or U13335 (N_13335,N_11447,N_12395);
and U13336 (N_13336,N_11848,N_10102);
and U13337 (N_13337,N_11691,N_11664);
nor U13338 (N_13338,N_12157,N_11130);
nand U13339 (N_13339,N_11611,N_10026);
or U13340 (N_13340,N_11369,N_11485);
nor U13341 (N_13341,N_12138,N_11806);
nor U13342 (N_13342,N_11137,N_12258);
or U13343 (N_13343,N_10532,N_11444);
or U13344 (N_13344,N_11451,N_10106);
or U13345 (N_13345,N_11920,N_10847);
nand U13346 (N_13346,N_12438,N_11448);
or U13347 (N_13347,N_11899,N_11328);
or U13348 (N_13348,N_10927,N_10742);
or U13349 (N_13349,N_10336,N_11776);
and U13350 (N_13350,N_12011,N_11052);
xor U13351 (N_13351,N_10078,N_12076);
nand U13352 (N_13352,N_10709,N_12075);
or U13353 (N_13353,N_12456,N_10095);
nand U13354 (N_13354,N_11916,N_10527);
xor U13355 (N_13355,N_10870,N_11973);
nor U13356 (N_13356,N_12024,N_10049);
xor U13357 (N_13357,N_12092,N_11417);
nand U13358 (N_13358,N_11251,N_11296);
or U13359 (N_13359,N_11094,N_11608);
nand U13360 (N_13360,N_11169,N_11111);
and U13361 (N_13361,N_11062,N_12300);
nor U13362 (N_13362,N_10827,N_12085);
nor U13363 (N_13363,N_10383,N_11737);
nand U13364 (N_13364,N_10902,N_10986);
nand U13365 (N_13365,N_10389,N_10593);
or U13366 (N_13366,N_11700,N_10807);
and U13367 (N_13367,N_10978,N_10138);
nand U13368 (N_13368,N_10630,N_11734);
xor U13369 (N_13369,N_11986,N_12319);
nor U13370 (N_13370,N_10039,N_10765);
xnor U13371 (N_13371,N_10290,N_12280);
nand U13372 (N_13372,N_10450,N_11000);
and U13373 (N_13373,N_10215,N_11637);
xor U13374 (N_13374,N_11565,N_12424);
nand U13375 (N_13375,N_10274,N_11650);
nand U13376 (N_13376,N_10390,N_12207);
and U13377 (N_13377,N_11221,N_12070);
nand U13378 (N_13378,N_11382,N_11454);
and U13379 (N_13379,N_11745,N_10485);
or U13380 (N_13380,N_12363,N_12457);
and U13381 (N_13381,N_10526,N_10362);
xor U13382 (N_13382,N_10431,N_12248);
xor U13383 (N_13383,N_11093,N_11344);
nor U13384 (N_13384,N_11257,N_10123);
nand U13385 (N_13385,N_10317,N_12343);
and U13386 (N_13386,N_10723,N_11823);
nand U13387 (N_13387,N_10550,N_11663);
and U13388 (N_13388,N_12259,N_11361);
and U13389 (N_13389,N_11205,N_11726);
xor U13390 (N_13390,N_12100,N_10271);
xnor U13391 (N_13391,N_10055,N_11307);
nand U13392 (N_13392,N_11021,N_10483);
nor U13393 (N_13393,N_11999,N_10667);
nor U13394 (N_13394,N_12194,N_12042);
xnor U13395 (N_13395,N_10580,N_10437);
or U13396 (N_13396,N_12028,N_12452);
nor U13397 (N_13397,N_11398,N_10418);
or U13398 (N_13398,N_11668,N_10003);
nand U13399 (N_13399,N_11045,N_11790);
or U13400 (N_13400,N_11323,N_10435);
or U13401 (N_13401,N_10842,N_12445);
nor U13402 (N_13402,N_11132,N_11978);
xnor U13403 (N_13403,N_10549,N_10603);
xor U13404 (N_13404,N_12149,N_10621);
nand U13405 (N_13405,N_10529,N_11827);
and U13406 (N_13406,N_11967,N_10567);
and U13407 (N_13407,N_10051,N_10885);
and U13408 (N_13408,N_12483,N_10656);
xnor U13409 (N_13409,N_10841,N_11753);
and U13410 (N_13410,N_11589,N_10571);
nand U13411 (N_13411,N_12213,N_11825);
nor U13412 (N_13412,N_11290,N_11261);
xnor U13413 (N_13413,N_11373,N_11299);
nand U13414 (N_13414,N_12163,N_11171);
nand U13415 (N_13415,N_10224,N_10589);
nor U13416 (N_13416,N_12436,N_10835);
nor U13417 (N_13417,N_11930,N_10623);
nor U13418 (N_13418,N_11803,N_12365);
nor U13419 (N_13419,N_11119,N_11614);
and U13420 (N_13420,N_10940,N_11088);
nand U13421 (N_13421,N_11641,N_10477);
xor U13422 (N_13422,N_11098,N_11773);
and U13423 (N_13423,N_12361,N_11337);
nor U13424 (N_13424,N_11658,N_11092);
nand U13425 (N_13425,N_11688,N_12351);
or U13426 (N_13426,N_11085,N_11729);
or U13427 (N_13427,N_10284,N_11804);
xor U13428 (N_13428,N_10096,N_10470);
nor U13429 (N_13429,N_11488,N_10458);
nand U13430 (N_13430,N_12134,N_11956);
or U13431 (N_13431,N_11336,N_11278);
nand U13432 (N_13432,N_11363,N_12099);
or U13433 (N_13433,N_11680,N_11191);
or U13434 (N_13434,N_11868,N_10761);
and U13435 (N_13435,N_11812,N_11461);
and U13436 (N_13436,N_11228,N_10454);
or U13437 (N_13437,N_12274,N_10505);
nand U13438 (N_13438,N_10561,N_10154);
nand U13439 (N_13439,N_10291,N_11371);
xnor U13440 (N_13440,N_11791,N_11506);
nor U13441 (N_13441,N_11164,N_11944);
or U13442 (N_13442,N_12307,N_11490);
or U13443 (N_13443,N_11055,N_11659);
or U13444 (N_13444,N_10562,N_11101);
nor U13445 (N_13445,N_11484,N_12265);
nand U13446 (N_13446,N_11176,N_11460);
xnor U13447 (N_13447,N_10688,N_12235);
nor U13448 (N_13448,N_11847,N_11433);
or U13449 (N_13449,N_10572,N_10540);
nand U13450 (N_13450,N_11148,N_11082);
or U13451 (N_13451,N_10354,N_10691);
nor U13452 (N_13452,N_12013,N_10166);
and U13453 (N_13453,N_11217,N_11886);
and U13454 (N_13454,N_10548,N_11104);
and U13455 (N_13455,N_10491,N_10013);
or U13456 (N_13456,N_10126,N_10258);
or U13457 (N_13457,N_11263,N_12224);
and U13458 (N_13458,N_12298,N_10995);
xor U13459 (N_13459,N_10213,N_10438);
xnor U13460 (N_13460,N_11332,N_11317);
nand U13461 (N_13461,N_10588,N_10471);
or U13462 (N_13462,N_10659,N_10430);
and U13463 (N_13463,N_11350,N_11482);
or U13464 (N_13464,N_12257,N_11961);
and U13465 (N_13465,N_11007,N_10424);
nor U13466 (N_13466,N_12197,N_11866);
or U13467 (N_13467,N_10776,N_11339);
or U13468 (N_13468,N_12411,N_11690);
and U13469 (N_13469,N_11521,N_11570);
nor U13470 (N_13470,N_10896,N_12285);
nand U13471 (N_13471,N_11078,N_11785);
nand U13472 (N_13472,N_11219,N_12358);
or U13473 (N_13473,N_11553,N_12443);
xnor U13474 (N_13474,N_11736,N_10506);
nor U13475 (N_13475,N_11179,N_11201);
or U13476 (N_13476,N_10232,N_10769);
and U13477 (N_13477,N_11995,N_10136);
nand U13478 (N_13478,N_11397,N_11975);
and U13479 (N_13479,N_10542,N_10134);
nand U13480 (N_13480,N_10530,N_11256);
xor U13481 (N_13481,N_11558,N_11306);
xnor U13482 (N_13482,N_10190,N_10230);
xor U13483 (N_13483,N_10678,N_10945);
nor U13484 (N_13484,N_10267,N_10692);
or U13485 (N_13485,N_10851,N_11701);
nor U13486 (N_13486,N_10647,N_11402);
or U13487 (N_13487,N_12079,N_12377);
xnor U13488 (N_13488,N_11907,N_10229);
or U13489 (N_13489,N_11462,N_10459);
and U13490 (N_13490,N_11598,N_11696);
or U13491 (N_13491,N_11655,N_10764);
or U13492 (N_13492,N_11869,N_12220);
nor U13493 (N_13493,N_10849,N_12253);
and U13494 (N_13494,N_11024,N_10590);
and U13495 (N_13495,N_10671,N_11204);
xnor U13496 (N_13496,N_11530,N_11019);
and U13497 (N_13497,N_10800,N_11360);
and U13498 (N_13498,N_11709,N_10669);
or U13499 (N_13499,N_11568,N_12185);
xor U13500 (N_13500,N_10689,N_12043);
or U13501 (N_13501,N_10934,N_12032);
nand U13502 (N_13502,N_10035,N_12293);
or U13503 (N_13503,N_10998,N_11574);
and U13504 (N_13504,N_11531,N_10507);
nor U13505 (N_13505,N_10059,N_10288);
or U13506 (N_13506,N_11026,N_12470);
and U13507 (N_13507,N_11238,N_11243);
and U13508 (N_13508,N_11226,N_11654);
or U13509 (N_13509,N_12434,N_12485);
and U13510 (N_13510,N_11455,N_10199);
and U13511 (N_13511,N_11933,N_10433);
nor U13512 (N_13512,N_10443,N_10314);
or U13513 (N_13513,N_11036,N_12186);
and U13514 (N_13514,N_10948,N_10070);
and U13515 (N_13515,N_12468,N_11463);
and U13516 (N_13516,N_10127,N_11362);
or U13517 (N_13517,N_11952,N_12227);
nand U13518 (N_13518,N_10240,N_12108);
xor U13519 (N_13519,N_10226,N_11921);
or U13520 (N_13520,N_11984,N_10950);
or U13521 (N_13521,N_10348,N_11918);
nor U13522 (N_13522,N_11750,N_12097);
xor U13523 (N_13523,N_11555,N_11216);
and U13524 (N_13524,N_10615,N_11281);
and U13525 (N_13525,N_10269,N_12152);
nand U13526 (N_13526,N_10705,N_12178);
xor U13527 (N_13527,N_12255,N_11591);
nor U13528 (N_13528,N_10539,N_10976);
nand U13529 (N_13529,N_11836,N_10770);
and U13530 (N_13530,N_11997,N_11850);
nand U13531 (N_13531,N_12435,N_10901);
nand U13532 (N_13532,N_11383,N_11387);
nand U13533 (N_13533,N_10220,N_10094);
nand U13534 (N_13534,N_11581,N_12191);
or U13535 (N_13535,N_12448,N_10308);
and U13536 (N_13536,N_12179,N_11128);
or U13537 (N_13537,N_11469,N_11384);
xnor U13538 (N_13538,N_12104,N_12127);
nand U13539 (N_13539,N_10923,N_10384);
nor U13540 (N_13540,N_11985,N_12312);
nand U13541 (N_13541,N_10627,N_10544);
nor U13542 (N_13542,N_12344,N_10802);
or U13543 (N_13543,N_12394,N_11218);
nand U13544 (N_13544,N_10575,N_11365);
nand U13545 (N_13545,N_10899,N_10641);
or U13546 (N_13546,N_11442,N_11877);
nand U13547 (N_13547,N_10262,N_10763);
nand U13548 (N_13548,N_10635,N_10894);
or U13549 (N_13549,N_12442,N_11667);
xnor U13550 (N_13550,N_10024,N_11181);
xnor U13551 (N_13551,N_11635,N_11324);
nand U13552 (N_13552,N_11903,N_10551);
nor U13553 (N_13553,N_11988,N_11234);
nor U13554 (N_13554,N_12125,N_12287);
nand U13555 (N_13555,N_12390,N_10309);
or U13556 (N_13556,N_11865,N_10068);
or U13557 (N_13557,N_11107,N_11926);
xnor U13558 (N_13558,N_11472,N_12473);
xor U13559 (N_13559,N_10748,N_11949);
xor U13560 (N_13560,N_10101,N_10803);
xnor U13561 (N_13561,N_10848,N_12497);
nor U13562 (N_13562,N_12341,N_10942);
or U13563 (N_13563,N_11077,N_11156);
xnor U13564 (N_13564,N_11035,N_12472);
or U13565 (N_13565,N_10990,N_12135);
xnor U13566 (N_13566,N_10836,N_11478);
and U13567 (N_13567,N_10717,N_12264);
nand U13568 (N_13568,N_11378,N_12484);
xnor U13569 (N_13569,N_12115,N_10991);
and U13570 (N_13570,N_11001,N_10100);
xnor U13571 (N_13571,N_10860,N_11513);
nand U13572 (N_13572,N_12034,N_12087);
nand U13573 (N_13573,N_10541,N_12096);
nor U13574 (N_13574,N_10771,N_10496);
nand U13575 (N_13575,N_10749,N_11253);
nand U13576 (N_13576,N_11267,N_12289);
xnor U13577 (N_13577,N_12459,N_11767);
nor U13578 (N_13578,N_12195,N_10946);
nor U13579 (N_13579,N_11309,N_10359);
or U13580 (N_13580,N_10799,N_10451);
and U13581 (N_13581,N_11057,N_11748);
nor U13582 (N_13582,N_11980,N_12371);
or U13583 (N_13583,N_10211,N_10402);
and U13584 (N_13584,N_11196,N_10448);
nor U13585 (N_13585,N_11733,N_11919);
nor U13586 (N_13586,N_10324,N_11028);
or U13587 (N_13587,N_11224,N_10900);
and U13588 (N_13588,N_11627,N_12384);
nand U13589 (N_13589,N_11291,N_11501);
nor U13590 (N_13590,N_11520,N_12077);
or U13591 (N_13591,N_11279,N_11771);
nor U13592 (N_13592,N_11359,N_12036);
or U13593 (N_13593,N_10512,N_10020);
and U13594 (N_13594,N_12050,N_11450);
xor U13595 (N_13595,N_10040,N_11441);
xor U13596 (N_13596,N_11534,N_11563);
and U13597 (N_13597,N_12035,N_11512);
xor U13598 (N_13598,N_10299,N_11102);
or U13599 (N_13599,N_11210,N_10318);
xor U13600 (N_13600,N_11860,N_11763);
or U13601 (N_13601,N_10618,N_11449);
nand U13602 (N_13602,N_10092,N_11676);
nor U13603 (N_13603,N_10204,N_11023);
or U13604 (N_13604,N_12230,N_11481);
nand U13605 (N_13605,N_11882,N_11452);
or U13606 (N_13606,N_12110,N_10263);
nand U13607 (N_13607,N_10696,N_11693);
nor U13608 (N_13608,N_10463,N_11262);
or U13609 (N_13609,N_11891,N_11159);
nand U13610 (N_13610,N_10556,N_10844);
xnor U13611 (N_13611,N_10367,N_11831);
nor U13612 (N_13612,N_11456,N_11413);
xnor U13613 (N_13613,N_10577,N_11504);
nor U13614 (N_13614,N_10747,N_10371);
and U13615 (N_13615,N_10428,N_11887);
or U13616 (N_13616,N_12159,N_10255);
nand U13617 (N_13617,N_10825,N_12492);
nand U13618 (N_13618,N_11818,N_11993);
and U13619 (N_13619,N_11604,N_10720);
xor U13620 (N_13620,N_11609,N_11225);
nor U13621 (N_13621,N_11543,N_12209);
nor U13622 (N_13622,N_11126,N_11661);
and U13623 (N_13623,N_11389,N_11935);
nand U13624 (N_13624,N_11554,N_10701);
xnor U13625 (N_13625,N_10634,N_10297);
xor U13626 (N_13626,N_10971,N_11617);
and U13627 (N_13627,N_11593,N_10977);
nor U13628 (N_13628,N_11459,N_10679);
xnor U13629 (N_13629,N_12169,N_12241);
nand U13630 (N_13630,N_10928,N_11705);
or U13631 (N_13631,N_12279,N_11808);
and U13632 (N_13632,N_11268,N_11275);
nor U13633 (N_13633,N_11177,N_10610);
xnor U13634 (N_13634,N_10777,N_11896);
nor U13635 (N_13635,N_11564,N_11757);
or U13636 (N_13636,N_11662,N_10814);
or U13637 (N_13637,N_10488,N_10524);
nand U13638 (N_13638,N_11535,N_10683);
nand U13639 (N_13639,N_12262,N_10406);
and U13640 (N_13640,N_10403,N_10514);
and U13641 (N_13641,N_11713,N_10086);
nor U13642 (N_13642,N_10619,N_12029);
and U13643 (N_13643,N_11720,N_10169);
nor U13644 (N_13644,N_12105,N_11286);
or U13645 (N_13645,N_11237,N_10128);
or U13646 (N_13646,N_11629,N_11333);
xnor U13647 (N_13647,N_12469,N_12167);
nor U13648 (N_13648,N_10167,N_12380);
xnor U13649 (N_13649,N_12314,N_11053);
nor U13650 (N_13650,N_10522,N_11430);
and U13651 (N_13651,N_10805,N_11118);
xor U13652 (N_13652,N_11259,N_12370);
nand U13653 (N_13653,N_10964,N_11630);
nor U13654 (N_13654,N_10077,N_11084);
or U13655 (N_13655,N_11293,N_11037);
or U13656 (N_13656,N_10801,N_10882);
and U13657 (N_13657,N_12283,N_11607);
nand U13658 (N_13658,N_11858,N_12199);
or U13659 (N_13659,N_11601,N_11507);
nor U13660 (N_13660,N_10554,N_12294);
xnor U13661 (N_13661,N_12398,N_11178);
xor U13662 (N_13662,N_10813,N_10187);
and U13663 (N_13663,N_11518,N_10781);
nand U13664 (N_13664,N_10775,N_10250);
or U13665 (N_13665,N_10887,N_12453);
and U13666 (N_13666,N_11594,N_11254);
and U13667 (N_13667,N_11820,N_12237);
or U13668 (N_13668,N_10714,N_10862);
or U13669 (N_13669,N_10171,N_11004);
xor U13670 (N_13670,N_10417,N_10325);
and U13671 (N_13671,N_11182,N_12455);
nand U13672 (N_13672,N_10029,N_10361);
nor U13673 (N_13673,N_11246,N_11859);
nand U13674 (N_13674,N_11724,N_12083);
nand U13675 (N_13675,N_10279,N_10034);
or U13676 (N_13676,N_11008,N_10722);
nand U13677 (N_13677,N_12217,N_11067);
nor U13678 (N_13678,N_12267,N_10811);
and U13679 (N_13679,N_11694,N_10281);
nor U13680 (N_13680,N_10511,N_11395);
nand U13681 (N_13681,N_11524,N_12401);
or U13682 (N_13682,N_11418,N_11120);
nand U13683 (N_13683,N_12177,N_12463);
nor U13684 (N_13684,N_11870,N_11538);
and U13685 (N_13685,N_12409,N_12474);
nand U13686 (N_13686,N_11959,N_11059);
or U13687 (N_13687,N_11584,N_10339);
and U13688 (N_13688,N_11807,N_12221);
and U13689 (N_13689,N_11552,N_10074);
xor U13690 (N_13690,N_12111,N_11623);
or U13691 (N_13691,N_11197,N_10519);
and U13692 (N_13692,N_12046,N_12412);
nand U13693 (N_13693,N_10392,N_11475);
xor U13694 (N_13694,N_10982,N_12415);
or U13695 (N_13695,N_11492,N_10386);
nand U13696 (N_13696,N_11491,N_11152);
xnor U13697 (N_13697,N_10677,N_10261);
xnor U13698 (N_13698,N_12421,N_12112);
or U13699 (N_13699,N_10277,N_12225);
nor U13700 (N_13700,N_11319,N_11139);
nand U13701 (N_13701,N_10413,N_11874);
nand U13702 (N_13702,N_11079,N_11730);
nand U13703 (N_13703,N_12460,N_11681);
xnor U13704 (N_13704,N_11432,N_11357);
nand U13705 (N_13705,N_11486,N_10253);
and U13706 (N_13706,N_12433,N_11212);
and U13707 (N_13707,N_10343,N_10943);
nor U13708 (N_13708,N_10082,N_11140);
nand U13709 (N_13709,N_10147,N_11121);
or U13710 (N_13710,N_11356,N_12331);
xor U13711 (N_13711,N_12131,N_10097);
xor U13712 (N_13712,N_10815,N_12069);
nand U13713 (N_13713,N_11288,N_11329);
or U13714 (N_13714,N_11962,N_11258);
and U13715 (N_13715,N_12078,N_11127);
and U13716 (N_13716,N_10489,N_12192);
or U13717 (N_13717,N_10089,N_10968);
nor U13718 (N_13718,N_11851,N_11453);
or U13719 (N_13719,N_10718,N_10854);
and U13720 (N_13720,N_10788,N_10008);
nor U13721 (N_13721,N_11640,N_11582);
nand U13722 (N_13722,N_10587,N_10460);
nor U13723 (N_13723,N_10620,N_10393);
nor U13724 (N_13724,N_10302,N_12019);
nor U13725 (N_13725,N_10884,N_11049);
xnor U13726 (N_13726,N_12005,N_11597);
nor U13727 (N_13727,N_11124,N_11536);
nand U13728 (N_13728,N_10104,N_10972);
or U13729 (N_13729,N_10312,N_11083);
or U13730 (N_13730,N_10681,N_11029);
nand U13731 (N_13731,N_12232,N_11778);
or U13732 (N_13732,N_10207,N_10142);
or U13733 (N_13733,N_11295,N_12353);
and U13734 (N_13734,N_10629,N_10120);
nand U13735 (N_13735,N_12498,N_10310);
xor U13736 (N_13736,N_10791,N_12218);
nand U13737 (N_13737,N_10787,N_12305);
or U13738 (N_13738,N_11405,N_11011);
or U13739 (N_13739,N_10002,N_10079);
and U13740 (N_13740,N_10372,N_11464);
or U13741 (N_13741,N_10926,N_12251);
and U13742 (N_13742,N_12041,N_10340);
nor U13743 (N_13743,N_11992,N_12444);
nand U13744 (N_13744,N_12189,N_12202);
or U13745 (N_13745,N_11511,N_11595);
xnor U13746 (N_13746,N_12155,N_12027);
and U13747 (N_13747,N_12142,N_11960);
or U13748 (N_13748,N_12272,N_10666);
xnor U13749 (N_13749,N_10753,N_10206);
and U13750 (N_13750,N_11984,N_12423);
and U13751 (N_13751,N_12464,N_10788);
or U13752 (N_13752,N_12296,N_10713);
xor U13753 (N_13753,N_12420,N_11685);
xor U13754 (N_13754,N_11922,N_12283);
nand U13755 (N_13755,N_10920,N_10804);
or U13756 (N_13756,N_10725,N_10326);
or U13757 (N_13757,N_12436,N_10631);
nand U13758 (N_13758,N_10691,N_10995);
nor U13759 (N_13759,N_11419,N_12064);
and U13760 (N_13760,N_10035,N_12058);
nor U13761 (N_13761,N_11924,N_10835);
and U13762 (N_13762,N_10876,N_11701);
nand U13763 (N_13763,N_10270,N_12226);
nand U13764 (N_13764,N_11382,N_10656);
nor U13765 (N_13765,N_11267,N_10448);
nand U13766 (N_13766,N_11056,N_11439);
and U13767 (N_13767,N_11662,N_12265);
and U13768 (N_13768,N_11072,N_12242);
and U13769 (N_13769,N_10653,N_12096);
or U13770 (N_13770,N_10843,N_11533);
xor U13771 (N_13771,N_11969,N_11447);
and U13772 (N_13772,N_10020,N_11631);
nor U13773 (N_13773,N_10714,N_12408);
and U13774 (N_13774,N_10202,N_11786);
and U13775 (N_13775,N_11898,N_12292);
and U13776 (N_13776,N_12422,N_10491);
and U13777 (N_13777,N_11170,N_10943);
or U13778 (N_13778,N_10087,N_11016);
nand U13779 (N_13779,N_10581,N_12499);
nor U13780 (N_13780,N_11743,N_10903);
and U13781 (N_13781,N_11276,N_11939);
nand U13782 (N_13782,N_11664,N_11271);
nand U13783 (N_13783,N_11951,N_12413);
nand U13784 (N_13784,N_11898,N_10385);
xnor U13785 (N_13785,N_11125,N_10543);
nand U13786 (N_13786,N_11930,N_11802);
xnor U13787 (N_13787,N_10793,N_11835);
and U13788 (N_13788,N_12098,N_12303);
and U13789 (N_13789,N_11647,N_10818);
nand U13790 (N_13790,N_11637,N_12488);
and U13791 (N_13791,N_11987,N_11087);
and U13792 (N_13792,N_10987,N_10862);
or U13793 (N_13793,N_11775,N_10721);
xnor U13794 (N_13794,N_11324,N_11660);
and U13795 (N_13795,N_11307,N_10370);
nor U13796 (N_13796,N_10385,N_11263);
or U13797 (N_13797,N_11957,N_11570);
nand U13798 (N_13798,N_12121,N_11826);
xnor U13799 (N_13799,N_11405,N_10829);
nor U13800 (N_13800,N_11183,N_10762);
nor U13801 (N_13801,N_11467,N_12495);
or U13802 (N_13802,N_11406,N_12133);
and U13803 (N_13803,N_10980,N_11637);
nand U13804 (N_13804,N_11639,N_12338);
xor U13805 (N_13805,N_10717,N_12073);
nor U13806 (N_13806,N_11858,N_12469);
nor U13807 (N_13807,N_11484,N_11381);
and U13808 (N_13808,N_11596,N_12329);
or U13809 (N_13809,N_10284,N_10901);
and U13810 (N_13810,N_11525,N_11874);
and U13811 (N_13811,N_11573,N_10239);
xnor U13812 (N_13812,N_12238,N_10360);
nor U13813 (N_13813,N_12232,N_11243);
and U13814 (N_13814,N_10553,N_10956);
or U13815 (N_13815,N_11980,N_10208);
or U13816 (N_13816,N_10072,N_10879);
nand U13817 (N_13817,N_12267,N_11302);
and U13818 (N_13818,N_12189,N_10945);
or U13819 (N_13819,N_10855,N_10829);
nor U13820 (N_13820,N_10658,N_10864);
or U13821 (N_13821,N_12465,N_11866);
xor U13822 (N_13822,N_10523,N_11612);
nor U13823 (N_13823,N_11035,N_10708);
or U13824 (N_13824,N_10257,N_12428);
xnor U13825 (N_13825,N_10276,N_11344);
xnor U13826 (N_13826,N_12432,N_10684);
nand U13827 (N_13827,N_10334,N_10810);
and U13828 (N_13828,N_10597,N_10978);
nor U13829 (N_13829,N_11392,N_12352);
and U13830 (N_13830,N_12129,N_11422);
nand U13831 (N_13831,N_11545,N_11636);
nor U13832 (N_13832,N_10553,N_11979);
or U13833 (N_13833,N_10602,N_11659);
xnor U13834 (N_13834,N_10760,N_10280);
xor U13835 (N_13835,N_10006,N_10463);
xor U13836 (N_13836,N_11874,N_11324);
and U13837 (N_13837,N_11868,N_10947);
and U13838 (N_13838,N_12137,N_12135);
xnor U13839 (N_13839,N_12496,N_11091);
nor U13840 (N_13840,N_11484,N_11520);
and U13841 (N_13841,N_12447,N_11712);
and U13842 (N_13842,N_11952,N_10011);
xnor U13843 (N_13843,N_12128,N_12164);
xnor U13844 (N_13844,N_10592,N_12179);
nand U13845 (N_13845,N_10397,N_11233);
xor U13846 (N_13846,N_12425,N_12080);
and U13847 (N_13847,N_11576,N_10756);
xor U13848 (N_13848,N_10809,N_11846);
or U13849 (N_13849,N_12339,N_10437);
and U13850 (N_13850,N_11748,N_12087);
xnor U13851 (N_13851,N_11343,N_10069);
and U13852 (N_13852,N_12251,N_10925);
or U13853 (N_13853,N_11011,N_11623);
xnor U13854 (N_13854,N_10446,N_10819);
xnor U13855 (N_13855,N_12194,N_11550);
or U13856 (N_13856,N_12465,N_10244);
nand U13857 (N_13857,N_11003,N_11458);
or U13858 (N_13858,N_12441,N_11861);
nor U13859 (N_13859,N_11584,N_10729);
nand U13860 (N_13860,N_10767,N_12213);
or U13861 (N_13861,N_10922,N_11022);
or U13862 (N_13862,N_10088,N_10950);
nor U13863 (N_13863,N_12384,N_11525);
or U13864 (N_13864,N_10059,N_11983);
or U13865 (N_13865,N_10954,N_12360);
nand U13866 (N_13866,N_10243,N_10123);
and U13867 (N_13867,N_11362,N_12464);
nor U13868 (N_13868,N_11368,N_12227);
or U13869 (N_13869,N_12417,N_12147);
and U13870 (N_13870,N_11801,N_10258);
and U13871 (N_13871,N_10903,N_10540);
and U13872 (N_13872,N_11559,N_11677);
and U13873 (N_13873,N_11921,N_10262);
xor U13874 (N_13874,N_12319,N_12377);
or U13875 (N_13875,N_11688,N_10065);
nand U13876 (N_13876,N_12428,N_11399);
and U13877 (N_13877,N_11559,N_11447);
nor U13878 (N_13878,N_12489,N_12087);
nand U13879 (N_13879,N_11372,N_11418);
nor U13880 (N_13880,N_12131,N_11526);
and U13881 (N_13881,N_11927,N_11419);
nor U13882 (N_13882,N_10006,N_11127);
xor U13883 (N_13883,N_10662,N_10689);
or U13884 (N_13884,N_12387,N_10577);
and U13885 (N_13885,N_10924,N_10352);
or U13886 (N_13886,N_10456,N_11905);
nand U13887 (N_13887,N_12361,N_10315);
nor U13888 (N_13888,N_11844,N_10820);
xor U13889 (N_13889,N_10817,N_12027);
xor U13890 (N_13890,N_10077,N_11352);
and U13891 (N_13891,N_11243,N_10498);
xnor U13892 (N_13892,N_12389,N_12223);
nand U13893 (N_13893,N_12112,N_10952);
nor U13894 (N_13894,N_10547,N_10024);
xnor U13895 (N_13895,N_10210,N_11518);
xnor U13896 (N_13896,N_11916,N_10656);
xor U13897 (N_13897,N_12112,N_12320);
xor U13898 (N_13898,N_12386,N_12277);
and U13899 (N_13899,N_10586,N_11275);
and U13900 (N_13900,N_11260,N_10398);
nor U13901 (N_13901,N_12293,N_10283);
or U13902 (N_13902,N_12488,N_10355);
xor U13903 (N_13903,N_10589,N_11363);
nand U13904 (N_13904,N_11912,N_11619);
or U13905 (N_13905,N_10093,N_11774);
nand U13906 (N_13906,N_12119,N_10207);
nand U13907 (N_13907,N_11474,N_10714);
nor U13908 (N_13908,N_11667,N_11016);
nor U13909 (N_13909,N_10814,N_11528);
and U13910 (N_13910,N_11503,N_12039);
nor U13911 (N_13911,N_12276,N_10331);
nor U13912 (N_13912,N_12337,N_12485);
nand U13913 (N_13913,N_11406,N_11384);
and U13914 (N_13914,N_10390,N_12354);
and U13915 (N_13915,N_11109,N_10957);
or U13916 (N_13916,N_11433,N_10551);
and U13917 (N_13917,N_12468,N_11151);
or U13918 (N_13918,N_10391,N_12088);
xnor U13919 (N_13919,N_10490,N_11035);
and U13920 (N_13920,N_11684,N_10897);
xor U13921 (N_13921,N_12261,N_11369);
nor U13922 (N_13922,N_10920,N_11861);
and U13923 (N_13923,N_11052,N_11541);
nand U13924 (N_13924,N_12406,N_10612);
xor U13925 (N_13925,N_11652,N_10257);
nand U13926 (N_13926,N_12416,N_10990);
xor U13927 (N_13927,N_12338,N_10885);
xnor U13928 (N_13928,N_11561,N_11826);
xor U13929 (N_13929,N_11166,N_11310);
nand U13930 (N_13930,N_12222,N_11952);
xnor U13931 (N_13931,N_12174,N_10571);
or U13932 (N_13932,N_10111,N_12023);
and U13933 (N_13933,N_11768,N_12429);
and U13934 (N_13934,N_10003,N_10006);
or U13935 (N_13935,N_10329,N_10662);
or U13936 (N_13936,N_11877,N_10386);
and U13937 (N_13937,N_10347,N_10568);
nand U13938 (N_13938,N_11105,N_10888);
nand U13939 (N_13939,N_11730,N_10148);
nor U13940 (N_13940,N_12191,N_10211);
and U13941 (N_13941,N_12092,N_11415);
or U13942 (N_13942,N_10972,N_12031);
or U13943 (N_13943,N_12123,N_10946);
nand U13944 (N_13944,N_10345,N_10811);
or U13945 (N_13945,N_10522,N_10479);
nor U13946 (N_13946,N_11537,N_12052);
and U13947 (N_13947,N_10951,N_12347);
nor U13948 (N_13948,N_10377,N_11614);
or U13949 (N_13949,N_12241,N_11508);
nand U13950 (N_13950,N_12355,N_12034);
nor U13951 (N_13951,N_12099,N_12133);
nand U13952 (N_13952,N_10110,N_11131);
nand U13953 (N_13953,N_10872,N_11436);
nand U13954 (N_13954,N_11824,N_11652);
nor U13955 (N_13955,N_10379,N_11044);
and U13956 (N_13956,N_10497,N_10989);
or U13957 (N_13957,N_11620,N_10986);
and U13958 (N_13958,N_12285,N_10203);
nand U13959 (N_13959,N_10885,N_10494);
xnor U13960 (N_13960,N_10753,N_10642);
xnor U13961 (N_13961,N_11086,N_10351);
or U13962 (N_13962,N_10976,N_11004);
nor U13963 (N_13963,N_10977,N_10236);
nand U13964 (N_13964,N_11693,N_12084);
nor U13965 (N_13965,N_11638,N_11379);
and U13966 (N_13966,N_10182,N_12144);
nand U13967 (N_13967,N_12146,N_11019);
nand U13968 (N_13968,N_10859,N_11122);
and U13969 (N_13969,N_11629,N_11855);
xor U13970 (N_13970,N_10023,N_10588);
or U13971 (N_13971,N_11058,N_11230);
and U13972 (N_13972,N_12315,N_10224);
xor U13973 (N_13973,N_10002,N_11626);
nand U13974 (N_13974,N_11199,N_10654);
and U13975 (N_13975,N_10720,N_12082);
and U13976 (N_13976,N_10487,N_10119);
and U13977 (N_13977,N_11150,N_11062);
nand U13978 (N_13978,N_11627,N_10801);
nand U13979 (N_13979,N_10483,N_12130);
nor U13980 (N_13980,N_11180,N_10287);
nand U13981 (N_13981,N_11424,N_10737);
or U13982 (N_13982,N_10763,N_10413);
nor U13983 (N_13983,N_12026,N_11931);
nand U13984 (N_13984,N_11582,N_10990);
nand U13985 (N_13985,N_10495,N_12074);
and U13986 (N_13986,N_11419,N_11519);
and U13987 (N_13987,N_10368,N_10659);
nand U13988 (N_13988,N_12293,N_11680);
nand U13989 (N_13989,N_10744,N_11717);
xor U13990 (N_13990,N_10533,N_12277);
xnor U13991 (N_13991,N_10151,N_10082);
and U13992 (N_13992,N_10723,N_12392);
nand U13993 (N_13993,N_10670,N_11553);
nand U13994 (N_13994,N_10445,N_11864);
nor U13995 (N_13995,N_12250,N_10736);
and U13996 (N_13996,N_12468,N_11844);
xor U13997 (N_13997,N_12375,N_11759);
nor U13998 (N_13998,N_10809,N_12389);
and U13999 (N_13999,N_10876,N_11953);
nand U14000 (N_14000,N_11249,N_10431);
nand U14001 (N_14001,N_10328,N_10348);
nand U14002 (N_14002,N_10391,N_10628);
nor U14003 (N_14003,N_11941,N_10846);
nor U14004 (N_14004,N_10829,N_10111);
and U14005 (N_14005,N_11768,N_12106);
xnor U14006 (N_14006,N_11739,N_12322);
xor U14007 (N_14007,N_10766,N_10388);
nor U14008 (N_14008,N_11070,N_11537);
nor U14009 (N_14009,N_10653,N_10993);
and U14010 (N_14010,N_11941,N_10497);
nor U14011 (N_14011,N_11603,N_10343);
nand U14012 (N_14012,N_11939,N_10970);
and U14013 (N_14013,N_10435,N_11393);
nand U14014 (N_14014,N_11503,N_10478);
nand U14015 (N_14015,N_10196,N_11517);
nand U14016 (N_14016,N_10937,N_11054);
nand U14017 (N_14017,N_10963,N_11587);
nand U14018 (N_14018,N_11454,N_10295);
xnor U14019 (N_14019,N_11616,N_10974);
and U14020 (N_14020,N_10030,N_12033);
nand U14021 (N_14021,N_10456,N_12369);
and U14022 (N_14022,N_11798,N_10344);
nor U14023 (N_14023,N_11901,N_10494);
or U14024 (N_14024,N_11086,N_10940);
nor U14025 (N_14025,N_12351,N_12147);
or U14026 (N_14026,N_11005,N_10460);
and U14027 (N_14027,N_10673,N_11458);
or U14028 (N_14028,N_11817,N_11026);
or U14029 (N_14029,N_10000,N_10830);
xor U14030 (N_14030,N_11277,N_10328);
nor U14031 (N_14031,N_10952,N_12359);
nor U14032 (N_14032,N_11604,N_10815);
nand U14033 (N_14033,N_10491,N_10572);
xnor U14034 (N_14034,N_10130,N_10794);
xnor U14035 (N_14035,N_10474,N_11278);
and U14036 (N_14036,N_10384,N_10768);
and U14037 (N_14037,N_11237,N_12299);
nand U14038 (N_14038,N_11068,N_10626);
nand U14039 (N_14039,N_11893,N_11546);
nor U14040 (N_14040,N_11082,N_11170);
xnor U14041 (N_14041,N_11166,N_11241);
nand U14042 (N_14042,N_10879,N_11002);
nor U14043 (N_14043,N_11028,N_11404);
nand U14044 (N_14044,N_11541,N_12158);
nand U14045 (N_14045,N_10503,N_11640);
nand U14046 (N_14046,N_10342,N_10025);
nand U14047 (N_14047,N_12411,N_11499);
nand U14048 (N_14048,N_11483,N_12176);
xor U14049 (N_14049,N_10453,N_12380);
xnor U14050 (N_14050,N_11228,N_10090);
xnor U14051 (N_14051,N_11486,N_11030);
or U14052 (N_14052,N_10813,N_10808);
nor U14053 (N_14053,N_11110,N_12088);
nand U14054 (N_14054,N_11513,N_11423);
or U14055 (N_14055,N_10285,N_10857);
or U14056 (N_14056,N_10453,N_12227);
and U14057 (N_14057,N_10822,N_12363);
nor U14058 (N_14058,N_11152,N_10641);
nor U14059 (N_14059,N_11376,N_10778);
xnor U14060 (N_14060,N_10760,N_12337);
or U14061 (N_14061,N_10209,N_12153);
and U14062 (N_14062,N_10047,N_10200);
and U14063 (N_14063,N_10818,N_10159);
nand U14064 (N_14064,N_12199,N_11769);
and U14065 (N_14065,N_10522,N_11612);
and U14066 (N_14066,N_11264,N_12232);
or U14067 (N_14067,N_10252,N_10411);
nor U14068 (N_14068,N_12465,N_11736);
nand U14069 (N_14069,N_10778,N_10007);
nor U14070 (N_14070,N_10044,N_11148);
or U14071 (N_14071,N_12178,N_10657);
or U14072 (N_14072,N_12399,N_11484);
nand U14073 (N_14073,N_10942,N_11030);
nor U14074 (N_14074,N_12218,N_11005);
nor U14075 (N_14075,N_11643,N_11970);
xnor U14076 (N_14076,N_10997,N_10021);
and U14077 (N_14077,N_10958,N_10017);
nand U14078 (N_14078,N_11079,N_10203);
and U14079 (N_14079,N_11772,N_11715);
xor U14080 (N_14080,N_11632,N_12293);
xor U14081 (N_14081,N_10481,N_12021);
and U14082 (N_14082,N_10636,N_10382);
nand U14083 (N_14083,N_11402,N_12308);
xnor U14084 (N_14084,N_11405,N_10134);
nand U14085 (N_14085,N_10499,N_11316);
nand U14086 (N_14086,N_10013,N_12388);
and U14087 (N_14087,N_11478,N_10372);
and U14088 (N_14088,N_11948,N_11389);
nand U14089 (N_14089,N_11315,N_10538);
or U14090 (N_14090,N_12383,N_11530);
nand U14091 (N_14091,N_12321,N_10412);
and U14092 (N_14092,N_10865,N_11396);
and U14093 (N_14093,N_12089,N_11937);
and U14094 (N_14094,N_11688,N_12312);
and U14095 (N_14095,N_10154,N_10901);
xor U14096 (N_14096,N_11785,N_11616);
nor U14097 (N_14097,N_10105,N_12486);
and U14098 (N_14098,N_11409,N_10771);
and U14099 (N_14099,N_10543,N_11385);
xor U14100 (N_14100,N_11403,N_10001);
xnor U14101 (N_14101,N_11299,N_11933);
xor U14102 (N_14102,N_12371,N_12272);
nor U14103 (N_14103,N_10010,N_12339);
or U14104 (N_14104,N_11978,N_10519);
xnor U14105 (N_14105,N_10683,N_12274);
xor U14106 (N_14106,N_11716,N_12202);
nor U14107 (N_14107,N_11955,N_11895);
or U14108 (N_14108,N_10258,N_11252);
nor U14109 (N_14109,N_10733,N_10656);
xor U14110 (N_14110,N_10418,N_11682);
or U14111 (N_14111,N_10418,N_12457);
xor U14112 (N_14112,N_11685,N_10338);
nand U14113 (N_14113,N_11680,N_11910);
and U14114 (N_14114,N_12237,N_11066);
and U14115 (N_14115,N_11952,N_12349);
or U14116 (N_14116,N_11571,N_12420);
nand U14117 (N_14117,N_11556,N_10697);
nand U14118 (N_14118,N_11506,N_10433);
and U14119 (N_14119,N_11411,N_11778);
nor U14120 (N_14120,N_11630,N_12207);
nand U14121 (N_14121,N_10819,N_11219);
nor U14122 (N_14122,N_11955,N_11925);
nand U14123 (N_14123,N_12090,N_12313);
or U14124 (N_14124,N_10512,N_12397);
nand U14125 (N_14125,N_10950,N_11394);
nor U14126 (N_14126,N_12063,N_12434);
or U14127 (N_14127,N_10556,N_11925);
or U14128 (N_14128,N_10705,N_11395);
or U14129 (N_14129,N_10603,N_11258);
or U14130 (N_14130,N_10411,N_12272);
or U14131 (N_14131,N_10189,N_11064);
or U14132 (N_14132,N_10417,N_12077);
or U14133 (N_14133,N_10436,N_11414);
xor U14134 (N_14134,N_10315,N_11136);
xor U14135 (N_14135,N_11622,N_11919);
nand U14136 (N_14136,N_10873,N_10333);
nor U14137 (N_14137,N_12284,N_11221);
nor U14138 (N_14138,N_10376,N_10262);
and U14139 (N_14139,N_10853,N_10808);
nor U14140 (N_14140,N_11907,N_12195);
nor U14141 (N_14141,N_12372,N_10695);
or U14142 (N_14142,N_11016,N_12001);
or U14143 (N_14143,N_11240,N_12307);
or U14144 (N_14144,N_10780,N_11045);
nand U14145 (N_14145,N_10998,N_10857);
nor U14146 (N_14146,N_10197,N_10221);
nand U14147 (N_14147,N_10698,N_11616);
or U14148 (N_14148,N_10413,N_12465);
and U14149 (N_14149,N_11971,N_11180);
and U14150 (N_14150,N_11525,N_11751);
nand U14151 (N_14151,N_11883,N_10656);
and U14152 (N_14152,N_10906,N_10027);
nor U14153 (N_14153,N_10670,N_10996);
and U14154 (N_14154,N_10194,N_11337);
and U14155 (N_14155,N_10091,N_11723);
xor U14156 (N_14156,N_11558,N_11597);
nand U14157 (N_14157,N_12376,N_12157);
nand U14158 (N_14158,N_10184,N_10463);
nand U14159 (N_14159,N_11012,N_10526);
and U14160 (N_14160,N_12348,N_11610);
xnor U14161 (N_14161,N_12073,N_11163);
xor U14162 (N_14162,N_12007,N_11241);
and U14163 (N_14163,N_11786,N_10727);
nor U14164 (N_14164,N_11351,N_10783);
xor U14165 (N_14165,N_10697,N_11774);
or U14166 (N_14166,N_11682,N_10978);
or U14167 (N_14167,N_10069,N_10218);
and U14168 (N_14168,N_10570,N_11457);
nor U14169 (N_14169,N_11127,N_12267);
or U14170 (N_14170,N_11916,N_10731);
nand U14171 (N_14171,N_11908,N_10656);
nand U14172 (N_14172,N_12058,N_12414);
or U14173 (N_14173,N_11190,N_11772);
nor U14174 (N_14174,N_12011,N_10009);
xnor U14175 (N_14175,N_11947,N_11489);
and U14176 (N_14176,N_11519,N_11489);
and U14177 (N_14177,N_11668,N_10639);
and U14178 (N_14178,N_10992,N_10348);
xnor U14179 (N_14179,N_10288,N_11299);
or U14180 (N_14180,N_10009,N_10655);
nor U14181 (N_14181,N_10357,N_10044);
and U14182 (N_14182,N_11928,N_11745);
nor U14183 (N_14183,N_10659,N_11434);
or U14184 (N_14184,N_11358,N_11732);
and U14185 (N_14185,N_11412,N_10769);
or U14186 (N_14186,N_11915,N_11122);
nor U14187 (N_14187,N_11322,N_10340);
xor U14188 (N_14188,N_11861,N_10894);
xor U14189 (N_14189,N_12424,N_10548);
and U14190 (N_14190,N_12331,N_11883);
nor U14191 (N_14191,N_10081,N_10938);
and U14192 (N_14192,N_11812,N_11454);
or U14193 (N_14193,N_10070,N_11533);
and U14194 (N_14194,N_10759,N_12052);
xnor U14195 (N_14195,N_10924,N_10945);
xor U14196 (N_14196,N_11766,N_10247);
xor U14197 (N_14197,N_11672,N_10445);
xnor U14198 (N_14198,N_11286,N_11223);
nand U14199 (N_14199,N_10841,N_11202);
xor U14200 (N_14200,N_10879,N_12136);
nand U14201 (N_14201,N_11444,N_10429);
nand U14202 (N_14202,N_12125,N_11939);
xnor U14203 (N_14203,N_11195,N_11630);
nor U14204 (N_14204,N_11286,N_12250);
xor U14205 (N_14205,N_10268,N_10997);
nor U14206 (N_14206,N_11163,N_10546);
nand U14207 (N_14207,N_11071,N_10902);
or U14208 (N_14208,N_12432,N_12099);
and U14209 (N_14209,N_11020,N_11333);
and U14210 (N_14210,N_12180,N_10102);
nand U14211 (N_14211,N_11238,N_10736);
nand U14212 (N_14212,N_10851,N_12217);
nand U14213 (N_14213,N_11019,N_11692);
or U14214 (N_14214,N_10770,N_10832);
xnor U14215 (N_14215,N_12175,N_11142);
nand U14216 (N_14216,N_10770,N_10533);
xor U14217 (N_14217,N_12410,N_10422);
and U14218 (N_14218,N_12429,N_10894);
or U14219 (N_14219,N_11754,N_10326);
xnor U14220 (N_14220,N_10069,N_12419);
nor U14221 (N_14221,N_11602,N_10403);
xnor U14222 (N_14222,N_12333,N_11881);
and U14223 (N_14223,N_10931,N_12290);
xor U14224 (N_14224,N_12277,N_12051);
xnor U14225 (N_14225,N_11055,N_10808);
nand U14226 (N_14226,N_11124,N_12415);
and U14227 (N_14227,N_11277,N_12090);
or U14228 (N_14228,N_12441,N_11337);
nor U14229 (N_14229,N_11955,N_11950);
xor U14230 (N_14230,N_11053,N_12105);
or U14231 (N_14231,N_10448,N_10536);
nor U14232 (N_14232,N_11034,N_10299);
and U14233 (N_14233,N_12134,N_11740);
nor U14234 (N_14234,N_11205,N_10759);
or U14235 (N_14235,N_12381,N_10015);
or U14236 (N_14236,N_10627,N_12224);
xnor U14237 (N_14237,N_11339,N_12059);
xor U14238 (N_14238,N_10018,N_11789);
nand U14239 (N_14239,N_10226,N_12407);
nand U14240 (N_14240,N_10529,N_10601);
or U14241 (N_14241,N_11658,N_11917);
xnor U14242 (N_14242,N_10394,N_10493);
or U14243 (N_14243,N_10893,N_10354);
and U14244 (N_14244,N_10056,N_10717);
xnor U14245 (N_14245,N_10839,N_12025);
nand U14246 (N_14246,N_10597,N_11706);
or U14247 (N_14247,N_12317,N_11059);
or U14248 (N_14248,N_11772,N_12146);
nand U14249 (N_14249,N_11210,N_11350);
nand U14250 (N_14250,N_11633,N_11392);
and U14251 (N_14251,N_12062,N_11520);
xnor U14252 (N_14252,N_10922,N_11020);
nor U14253 (N_14253,N_10713,N_10407);
and U14254 (N_14254,N_12349,N_10058);
and U14255 (N_14255,N_10562,N_10700);
nand U14256 (N_14256,N_10920,N_10292);
xnor U14257 (N_14257,N_10661,N_12009);
nand U14258 (N_14258,N_12243,N_10107);
and U14259 (N_14259,N_10143,N_10332);
nor U14260 (N_14260,N_12092,N_10012);
and U14261 (N_14261,N_11785,N_12128);
or U14262 (N_14262,N_10731,N_10177);
or U14263 (N_14263,N_12466,N_11638);
and U14264 (N_14264,N_11498,N_11522);
and U14265 (N_14265,N_12099,N_11480);
or U14266 (N_14266,N_11467,N_12474);
nor U14267 (N_14267,N_10220,N_12326);
and U14268 (N_14268,N_11961,N_10949);
or U14269 (N_14269,N_12406,N_12210);
nand U14270 (N_14270,N_11177,N_12317);
and U14271 (N_14271,N_11924,N_11489);
and U14272 (N_14272,N_12097,N_10777);
and U14273 (N_14273,N_11424,N_11701);
xnor U14274 (N_14274,N_12399,N_11662);
nor U14275 (N_14275,N_11910,N_10121);
xnor U14276 (N_14276,N_10994,N_12314);
nand U14277 (N_14277,N_11316,N_10411);
and U14278 (N_14278,N_10758,N_12112);
and U14279 (N_14279,N_11843,N_12372);
nor U14280 (N_14280,N_11900,N_11686);
or U14281 (N_14281,N_11763,N_11711);
and U14282 (N_14282,N_10782,N_12460);
nor U14283 (N_14283,N_11709,N_10485);
nand U14284 (N_14284,N_11373,N_10461);
and U14285 (N_14285,N_10810,N_12314);
or U14286 (N_14286,N_10262,N_11400);
nand U14287 (N_14287,N_12014,N_11555);
or U14288 (N_14288,N_10530,N_11833);
or U14289 (N_14289,N_11421,N_10879);
and U14290 (N_14290,N_10253,N_12266);
nand U14291 (N_14291,N_10438,N_12247);
or U14292 (N_14292,N_11258,N_11196);
or U14293 (N_14293,N_11935,N_11023);
and U14294 (N_14294,N_12143,N_11977);
and U14295 (N_14295,N_12110,N_10081);
xnor U14296 (N_14296,N_10185,N_10198);
nand U14297 (N_14297,N_10307,N_10473);
nand U14298 (N_14298,N_10452,N_10463);
nand U14299 (N_14299,N_10615,N_11097);
nand U14300 (N_14300,N_10679,N_10740);
nor U14301 (N_14301,N_10727,N_12177);
or U14302 (N_14302,N_10253,N_10770);
nand U14303 (N_14303,N_10417,N_10569);
xnor U14304 (N_14304,N_11050,N_11804);
nand U14305 (N_14305,N_10136,N_12032);
and U14306 (N_14306,N_12249,N_11157);
and U14307 (N_14307,N_11612,N_11511);
xnor U14308 (N_14308,N_12046,N_10746);
nand U14309 (N_14309,N_11225,N_11029);
and U14310 (N_14310,N_11327,N_10389);
xor U14311 (N_14311,N_10506,N_10353);
and U14312 (N_14312,N_10573,N_11018);
nand U14313 (N_14313,N_11802,N_11583);
or U14314 (N_14314,N_10242,N_10334);
and U14315 (N_14315,N_12176,N_12263);
xor U14316 (N_14316,N_12469,N_12431);
and U14317 (N_14317,N_10074,N_11448);
or U14318 (N_14318,N_11275,N_10037);
nand U14319 (N_14319,N_11419,N_12116);
xor U14320 (N_14320,N_10801,N_11049);
nand U14321 (N_14321,N_10838,N_10212);
xnor U14322 (N_14322,N_11460,N_11647);
nor U14323 (N_14323,N_11319,N_12311);
xor U14324 (N_14324,N_12254,N_11867);
or U14325 (N_14325,N_12439,N_12428);
xor U14326 (N_14326,N_10551,N_12459);
or U14327 (N_14327,N_10312,N_12054);
and U14328 (N_14328,N_12491,N_10552);
or U14329 (N_14329,N_12029,N_10544);
xor U14330 (N_14330,N_11321,N_10879);
nand U14331 (N_14331,N_10908,N_10213);
nand U14332 (N_14332,N_10131,N_10316);
nand U14333 (N_14333,N_11595,N_12255);
and U14334 (N_14334,N_12401,N_12268);
or U14335 (N_14335,N_12070,N_10136);
nor U14336 (N_14336,N_12168,N_11802);
xnor U14337 (N_14337,N_12259,N_11213);
or U14338 (N_14338,N_11526,N_11645);
nor U14339 (N_14339,N_10642,N_11894);
nand U14340 (N_14340,N_10381,N_11343);
or U14341 (N_14341,N_11725,N_12024);
xnor U14342 (N_14342,N_11420,N_10511);
xor U14343 (N_14343,N_10636,N_12395);
nand U14344 (N_14344,N_10435,N_11050);
xor U14345 (N_14345,N_10639,N_11273);
nand U14346 (N_14346,N_10988,N_11443);
or U14347 (N_14347,N_11689,N_11757);
nor U14348 (N_14348,N_10257,N_11819);
nor U14349 (N_14349,N_11802,N_10255);
nor U14350 (N_14350,N_10662,N_11671);
and U14351 (N_14351,N_10797,N_10267);
xnor U14352 (N_14352,N_11769,N_10731);
and U14353 (N_14353,N_11596,N_11411);
or U14354 (N_14354,N_10844,N_12498);
nor U14355 (N_14355,N_11177,N_11448);
nor U14356 (N_14356,N_11094,N_10558);
xnor U14357 (N_14357,N_10002,N_11455);
nor U14358 (N_14358,N_11550,N_12032);
xor U14359 (N_14359,N_10342,N_10343);
or U14360 (N_14360,N_11462,N_11300);
xor U14361 (N_14361,N_11852,N_11010);
and U14362 (N_14362,N_12165,N_12327);
nand U14363 (N_14363,N_10337,N_11408);
nor U14364 (N_14364,N_11383,N_10954);
and U14365 (N_14365,N_10650,N_11239);
and U14366 (N_14366,N_10231,N_10286);
nor U14367 (N_14367,N_11571,N_10234);
and U14368 (N_14368,N_11205,N_10246);
and U14369 (N_14369,N_12223,N_11942);
nor U14370 (N_14370,N_10261,N_11175);
or U14371 (N_14371,N_11517,N_11787);
or U14372 (N_14372,N_10213,N_11938);
nand U14373 (N_14373,N_11445,N_12108);
xor U14374 (N_14374,N_11565,N_12044);
and U14375 (N_14375,N_12385,N_11227);
and U14376 (N_14376,N_10930,N_11464);
xor U14377 (N_14377,N_10586,N_10625);
and U14378 (N_14378,N_12165,N_12151);
nand U14379 (N_14379,N_12137,N_12351);
nor U14380 (N_14380,N_10530,N_10082);
and U14381 (N_14381,N_10251,N_11001);
nor U14382 (N_14382,N_12244,N_10868);
nand U14383 (N_14383,N_10535,N_11715);
nand U14384 (N_14384,N_12195,N_11045);
nand U14385 (N_14385,N_12255,N_11657);
xor U14386 (N_14386,N_12247,N_10233);
and U14387 (N_14387,N_11296,N_11050);
or U14388 (N_14388,N_10265,N_12405);
or U14389 (N_14389,N_11802,N_11499);
xnor U14390 (N_14390,N_11852,N_10616);
nand U14391 (N_14391,N_11416,N_11188);
or U14392 (N_14392,N_11833,N_10453);
and U14393 (N_14393,N_10801,N_11894);
nor U14394 (N_14394,N_12059,N_12441);
nor U14395 (N_14395,N_11307,N_12328);
nor U14396 (N_14396,N_10132,N_10676);
xor U14397 (N_14397,N_11449,N_10374);
or U14398 (N_14398,N_11198,N_11530);
or U14399 (N_14399,N_11130,N_11929);
nand U14400 (N_14400,N_11390,N_11991);
nand U14401 (N_14401,N_11308,N_11935);
nand U14402 (N_14402,N_11745,N_10863);
nand U14403 (N_14403,N_12190,N_10869);
nor U14404 (N_14404,N_11212,N_10937);
xnor U14405 (N_14405,N_10281,N_11726);
and U14406 (N_14406,N_10362,N_10654);
nand U14407 (N_14407,N_10414,N_11006);
xnor U14408 (N_14408,N_10786,N_11430);
or U14409 (N_14409,N_10250,N_10555);
nor U14410 (N_14410,N_11266,N_10129);
nor U14411 (N_14411,N_11998,N_10821);
nor U14412 (N_14412,N_12231,N_12168);
nor U14413 (N_14413,N_10980,N_10934);
or U14414 (N_14414,N_10318,N_10027);
or U14415 (N_14415,N_11197,N_10679);
nand U14416 (N_14416,N_12277,N_11686);
nor U14417 (N_14417,N_10938,N_10568);
xnor U14418 (N_14418,N_11451,N_11075);
xnor U14419 (N_14419,N_10207,N_11189);
nand U14420 (N_14420,N_10074,N_11644);
xnor U14421 (N_14421,N_10326,N_11123);
nand U14422 (N_14422,N_11656,N_12314);
nand U14423 (N_14423,N_11789,N_11052);
nand U14424 (N_14424,N_10670,N_10307);
and U14425 (N_14425,N_11826,N_11577);
xnor U14426 (N_14426,N_11847,N_10397);
and U14427 (N_14427,N_11868,N_12439);
and U14428 (N_14428,N_11500,N_11420);
nor U14429 (N_14429,N_12124,N_11783);
nand U14430 (N_14430,N_10939,N_12472);
or U14431 (N_14431,N_10400,N_11497);
or U14432 (N_14432,N_10165,N_10271);
nor U14433 (N_14433,N_11550,N_11973);
nand U14434 (N_14434,N_10625,N_10957);
nand U14435 (N_14435,N_11907,N_10138);
xnor U14436 (N_14436,N_10388,N_10377);
xnor U14437 (N_14437,N_10751,N_10744);
and U14438 (N_14438,N_10082,N_10038);
nor U14439 (N_14439,N_10976,N_12387);
xor U14440 (N_14440,N_11285,N_12181);
nor U14441 (N_14441,N_11572,N_10723);
and U14442 (N_14442,N_12217,N_12109);
or U14443 (N_14443,N_11443,N_11818);
or U14444 (N_14444,N_10687,N_11141);
nor U14445 (N_14445,N_10934,N_12448);
or U14446 (N_14446,N_11739,N_12450);
nor U14447 (N_14447,N_10102,N_11656);
or U14448 (N_14448,N_10197,N_12174);
and U14449 (N_14449,N_12191,N_11499);
xnor U14450 (N_14450,N_11999,N_10364);
nand U14451 (N_14451,N_10686,N_11388);
xor U14452 (N_14452,N_12003,N_12327);
nor U14453 (N_14453,N_11072,N_11725);
nand U14454 (N_14454,N_11723,N_12025);
xnor U14455 (N_14455,N_11888,N_10790);
nor U14456 (N_14456,N_10440,N_11553);
nand U14457 (N_14457,N_12296,N_10116);
and U14458 (N_14458,N_11542,N_11299);
and U14459 (N_14459,N_10671,N_11515);
nor U14460 (N_14460,N_10309,N_11212);
and U14461 (N_14461,N_10661,N_10287);
nor U14462 (N_14462,N_12006,N_11957);
and U14463 (N_14463,N_10931,N_10366);
xor U14464 (N_14464,N_10441,N_11933);
or U14465 (N_14465,N_11069,N_12173);
nor U14466 (N_14466,N_11574,N_10423);
nand U14467 (N_14467,N_10558,N_10364);
nor U14468 (N_14468,N_10642,N_11699);
xor U14469 (N_14469,N_11178,N_10680);
xnor U14470 (N_14470,N_11918,N_10303);
or U14471 (N_14471,N_12332,N_11264);
xor U14472 (N_14472,N_11358,N_10093);
or U14473 (N_14473,N_12408,N_11503);
xor U14474 (N_14474,N_10517,N_10027);
and U14475 (N_14475,N_10489,N_12021);
nor U14476 (N_14476,N_11497,N_11157);
or U14477 (N_14477,N_10721,N_12246);
or U14478 (N_14478,N_11516,N_10692);
nor U14479 (N_14479,N_12340,N_11168);
nor U14480 (N_14480,N_10658,N_12436);
xor U14481 (N_14481,N_10103,N_12038);
nand U14482 (N_14482,N_10054,N_11814);
xnor U14483 (N_14483,N_11246,N_10460);
or U14484 (N_14484,N_10013,N_12426);
nor U14485 (N_14485,N_12133,N_12080);
xor U14486 (N_14486,N_11599,N_12040);
xor U14487 (N_14487,N_10723,N_10675);
xor U14488 (N_14488,N_10105,N_10144);
and U14489 (N_14489,N_11643,N_12133);
xnor U14490 (N_14490,N_10822,N_10597);
xnor U14491 (N_14491,N_11043,N_10807);
xnor U14492 (N_14492,N_12253,N_11792);
and U14493 (N_14493,N_10988,N_10656);
nand U14494 (N_14494,N_10546,N_11226);
and U14495 (N_14495,N_11369,N_11048);
and U14496 (N_14496,N_11693,N_11799);
nor U14497 (N_14497,N_12132,N_10925);
and U14498 (N_14498,N_10273,N_10135);
nand U14499 (N_14499,N_11447,N_12157);
nand U14500 (N_14500,N_11975,N_12399);
nand U14501 (N_14501,N_10158,N_11409);
and U14502 (N_14502,N_11806,N_12134);
nor U14503 (N_14503,N_11361,N_11491);
nand U14504 (N_14504,N_10788,N_12196);
or U14505 (N_14505,N_10602,N_11050);
xor U14506 (N_14506,N_10638,N_10287);
xor U14507 (N_14507,N_11017,N_10447);
nand U14508 (N_14508,N_11505,N_10324);
nand U14509 (N_14509,N_11354,N_11277);
and U14510 (N_14510,N_12337,N_12190);
or U14511 (N_14511,N_10835,N_10207);
or U14512 (N_14512,N_12353,N_12227);
nand U14513 (N_14513,N_10562,N_11263);
nor U14514 (N_14514,N_10252,N_10595);
xnor U14515 (N_14515,N_11533,N_11694);
nand U14516 (N_14516,N_11197,N_10081);
nand U14517 (N_14517,N_11964,N_12276);
xnor U14518 (N_14518,N_11939,N_11954);
nand U14519 (N_14519,N_10260,N_11758);
or U14520 (N_14520,N_11138,N_10222);
nand U14521 (N_14521,N_11831,N_10995);
nor U14522 (N_14522,N_11355,N_10513);
xnor U14523 (N_14523,N_10585,N_11684);
and U14524 (N_14524,N_10861,N_11258);
nand U14525 (N_14525,N_11314,N_12439);
nand U14526 (N_14526,N_11211,N_11533);
xnor U14527 (N_14527,N_11589,N_10834);
nor U14528 (N_14528,N_10871,N_12437);
xor U14529 (N_14529,N_10206,N_10713);
nand U14530 (N_14530,N_12019,N_10039);
or U14531 (N_14531,N_10602,N_10642);
nand U14532 (N_14532,N_11073,N_12026);
nand U14533 (N_14533,N_10369,N_11131);
nand U14534 (N_14534,N_10482,N_11798);
and U14535 (N_14535,N_10093,N_10127);
or U14536 (N_14536,N_12139,N_12403);
or U14537 (N_14537,N_11736,N_11656);
xor U14538 (N_14538,N_10700,N_12384);
nand U14539 (N_14539,N_11645,N_11781);
or U14540 (N_14540,N_11887,N_11008);
nor U14541 (N_14541,N_10956,N_12064);
or U14542 (N_14542,N_10154,N_10057);
or U14543 (N_14543,N_11704,N_11716);
xor U14544 (N_14544,N_12006,N_12270);
xor U14545 (N_14545,N_12497,N_10477);
or U14546 (N_14546,N_10533,N_12320);
xor U14547 (N_14547,N_11582,N_12245);
nand U14548 (N_14548,N_10559,N_10677);
and U14549 (N_14549,N_10394,N_12072);
and U14550 (N_14550,N_11644,N_11564);
and U14551 (N_14551,N_11132,N_10715);
and U14552 (N_14552,N_11364,N_11855);
nor U14553 (N_14553,N_11928,N_10873);
nor U14554 (N_14554,N_12431,N_10578);
or U14555 (N_14555,N_10236,N_10388);
nor U14556 (N_14556,N_11725,N_12167);
xor U14557 (N_14557,N_10813,N_10267);
and U14558 (N_14558,N_10203,N_10940);
nand U14559 (N_14559,N_11878,N_12120);
xnor U14560 (N_14560,N_10866,N_11606);
and U14561 (N_14561,N_10918,N_11099);
nor U14562 (N_14562,N_11287,N_10913);
nand U14563 (N_14563,N_11900,N_11031);
xor U14564 (N_14564,N_10141,N_10507);
nand U14565 (N_14565,N_10720,N_12465);
or U14566 (N_14566,N_10333,N_12395);
and U14567 (N_14567,N_11777,N_10915);
nand U14568 (N_14568,N_11463,N_11234);
or U14569 (N_14569,N_12158,N_10175);
and U14570 (N_14570,N_10085,N_10310);
nand U14571 (N_14571,N_11118,N_11333);
xnor U14572 (N_14572,N_10836,N_11531);
and U14573 (N_14573,N_11544,N_11816);
or U14574 (N_14574,N_11146,N_10029);
nand U14575 (N_14575,N_12486,N_11603);
or U14576 (N_14576,N_12192,N_12077);
nand U14577 (N_14577,N_11423,N_11795);
xnor U14578 (N_14578,N_10315,N_12064);
xor U14579 (N_14579,N_11380,N_10635);
nand U14580 (N_14580,N_11793,N_11623);
and U14581 (N_14581,N_12436,N_10303);
or U14582 (N_14582,N_11855,N_12412);
and U14583 (N_14583,N_11536,N_11380);
nand U14584 (N_14584,N_10564,N_11194);
or U14585 (N_14585,N_11856,N_10142);
or U14586 (N_14586,N_10062,N_11282);
nor U14587 (N_14587,N_11145,N_10069);
xor U14588 (N_14588,N_10812,N_11724);
or U14589 (N_14589,N_10070,N_11398);
and U14590 (N_14590,N_10227,N_11892);
and U14591 (N_14591,N_10942,N_11832);
or U14592 (N_14592,N_11373,N_11170);
or U14593 (N_14593,N_12159,N_12432);
nor U14594 (N_14594,N_11127,N_10187);
xor U14595 (N_14595,N_10992,N_10661);
and U14596 (N_14596,N_10820,N_11625);
xnor U14597 (N_14597,N_10380,N_11069);
and U14598 (N_14598,N_10028,N_11788);
or U14599 (N_14599,N_11603,N_12050);
and U14600 (N_14600,N_10581,N_10227);
and U14601 (N_14601,N_12132,N_12423);
xor U14602 (N_14602,N_10410,N_12063);
or U14603 (N_14603,N_11568,N_12464);
nand U14604 (N_14604,N_11422,N_10674);
nor U14605 (N_14605,N_11698,N_11699);
and U14606 (N_14606,N_10161,N_10383);
nand U14607 (N_14607,N_11161,N_10009);
xor U14608 (N_14608,N_11009,N_11271);
xnor U14609 (N_14609,N_12226,N_11043);
xor U14610 (N_14610,N_11071,N_11579);
xnor U14611 (N_14611,N_11770,N_12261);
and U14612 (N_14612,N_11867,N_11110);
nor U14613 (N_14613,N_10756,N_10342);
and U14614 (N_14614,N_11928,N_11955);
nor U14615 (N_14615,N_11439,N_11662);
and U14616 (N_14616,N_11874,N_11733);
or U14617 (N_14617,N_12086,N_11942);
and U14618 (N_14618,N_11070,N_10981);
or U14619 (N_14619,N_10292,N_11390);
xnor U14620 (N_14620,N_11782,N_11366);
nand U14621 (N_14621,N_10415,N_10802);
xnor U14622 (N_14622,N_10289,N_10535);
and U14623 (N_14623,N_11438,N_11371);
nor U14624 (N_14624,N_11593,N_11665);
nor U14625 (N_14625,N_10510,N_12175);
or U14626 (N_14626,N_11437,N_11689);
or U14627 (N_14627,N_10312,N_10579);
or U14628 (N_14628,N_11882,N_10055);
nor U14629 (N_14629,N_11185,N_10520);
and U14630 (N_14630,N_12359,N_11123);
or U14631 (N_14631,N_11814,N_12142);
nor U14632 (N_14632,N_10953,N_10676);
or U14633 (N_14633,N_10766,N_11733);
nand U14634 (N_14634,N_11230,N_11362);
nand U14635 (N_14635,N_11172,N_11435);
and U14636 (N_14636,N_10816,N_12411);
or U14637 (N_14637,N_12061,N_10406);
or U14638 (N_14638,N_10971,N_10415);
xor U14639 (N_14639,N_11113,N_12308);
nor U14640 (N_14640,N_11105,N_10427);
or U14641 (N_14641,N_11198,N_12327);
xnor U14642 (N_14642,N_11022,N_11388);
or U14643 (N_14643,N_10710,N_10336);
nor U14644 (N_14644,N_12188,N_10918);
nor U14645 (N_14645,N_11137,N_11800);
nor U14646 (N_14646,N_10157,N_11753);
nor U14647 (N_14647,N_11656,N_12454);
and U14648 (N_14648,N_10243,N_12100);
or U14649 (N_14649,N_11298,N_12248);
or U14650 (N_14650,N_10344,N_11252);
nand U14651 (N_14651,N_11162,N_11398);
and U14652 (N_14652,N_10015,N_10061);
xnor U14653 (N_14653,N_11015,N_11366);
and U14654 (N_14654,N_10047,N_12105);
nor U14655 (N_14655,N_10561,N_10209);
nand U14656 (N_14656,N_10744,N_10951);
nand U14657 (N_14657,N_10519,N_11441);
nand U14658 (N_14658,N_12006,N_11192);
or U14659 (N_14659,N_10874,N_11513);
nand U14660 (N_14660,N_10762,N_10153);
or U14661 (N_14661,N_10165,N_12256);
nand U14662 (N_14662,N_11886,N_11449);
nand U14663 (N_14663,N_11799,N_10612);
or U14664 (N_14664,N_10536,N_11974);
nor U14665 (N_14665,N_10151,N_12497);
nand U14666 (N_14666,N_10560,N_11832);
or U14667 (N_14667,N_10597,N_11560);
and U14668 (N_14668,N_11034,N_10796);
nor U14669 (N_14669,N_10308,N_10893);
xnor U14670 (N_14670,N_10611,N_11024);
xor U14671 (N_14671,N_11974,N_11265);
nand U14672 (N_14672,N_11784,N_10871);
or U14673 (N_14673,N_11906,N_10302);
or U14674 (N_14674,N_11435,N_11237);
xnor U14675 (N_14675,N_11712,N_10459);
and U14676 (N_14676,N_11066,N_11792);
nand U14677 (N_14677,N_12334,N_11961);
xnor U14678 (N_14678,N_11090,N_10507);
or U14679 (N_14679,N_11281,N_10005);
nand U14680 (N_14680,N_12225,N_10373);
nor U14681 (N_14681,N_12414,N_10878);
nor U14682 (N_14682,N_10785,N_11541);
or U14683 (N_14683,N_12260,N_10690);
nor U14684 (N_14684,N_10965,N_12358);
or U14685 (N_14685,N_10982,N_11847);
nor U14686 (N_14686,N_10056,N_10012);
or U14687 (N_14687,N_11457,N_12262);
and U14688 (N_14688,N_10226,N_11669);
and U14689 (N_14689,N_10697,N_12287);
or U14690 (N_14690,N_11544,N_12285);
nand U14691 (N_14691,N_10804,N_10495);
or U14692 (N_14692,N_11264,N_10312);
or U14693 (N_14693,N_10401,N_10211);
and U14694 (N_14694,N_11845,N_12340);
nand U14695 (N_14695,N_10839,N_12051);
and U14696 (N_14696,N_12193,N_11549);
and U14697 (N_14697,N_12157,N_10777);
nand U14698 (N_14698,N_11780,N_11118);
and U14699 (N_14699,N_10290,N_11304);
and U14700 (N_14700,N_11209,N_10095);
nand U14701 (N_14701,N_12194,N_10713);
xor U14702 (N_14702,N_12380,N_10576);
or U14703 (N_14703,N_12138,N_10841);
or U14704 (N_14704,N_11664,N_10323);
nand U14705 (N_14705,N_10268,N_12125);
nand U14706 (N_14706,N_10874,N_11466);
nor U14707 (N_14707,N_10958,N_11440);
and U14708 (N_14708,N_10128,N_11850);
nor U14709 (N_14709,N_12056,N_12148);
or U14710 (N_14710,N_10596,N_12422);
xnor U14711 (N_14711,N_11574,N_10586);
xnor U14712 (N_14712,N_10675,N_11792);
or U14713 (N_14713,N_11068,N_11309);
nor U14714 (N_14714,N_12275,N_11663);
xor U14715 (N_14715,N_12257,N_12345);
nand U14716 (N_14716,N_11982,N_11542);
or U14717 (N_14717,N_10794,N_12059);
nand U14718 (N_14718,N_11224,N_12128);
nor U14719 (N_14719,N_11693,N_10960);
nand U14720 (N_14720,N_10920,N_11193);
or U14721 (N_14721,N_10208,N_11524);
nand U14722 (N_14722,N_11810,N_10262);
and U14723 (N_14723,N_10448,N_10525);
or U14724 (N_14724,N_11346,N_12188);
and U14725 (N_14725,N_10798,N_12182);
or U14726 (N_14726,N_10638,N_11908);
xor U14727 (N_14727,N_10276,N_10335);
and U14728 (N_14728,N_11147,N_10380);
xnor U14729 (N_14729,N_10217,N_12104);
or U14730 (N_14730,N_11805,N_12473);
nand U14731 (N_14731,N_10366,N_11700);
xor U14732 (N_14732,N_11474,N_10993);
and U14733 (N_14733,N_10359,N_11667);
or U14734 (N_14734,N_10910,N_11472);
xnor U14735 (N_14735,N_10476,N_10044);
xnor U14736 (N_14736,N_10988,N_10329);
xor U14737 (N_14737,N_10454,N_10356);
nand U14738 (N_14738,N_10745,N_11720);
nand U14739 (N_14739,N_10043,N_11147);
nor U14740 (N_14740,N_10857,N_11396);
and U14741 (N_14741,N_11355,N_12361);
or U14742 (N_14742,N_11965,N_12089);
xnor U14743 (N_14743,N_10003,N_10794);
or U14744 (N_14744,N_11795,N_11350);
xor U14745 (N_14745,N_10417,N_12028);
or U14746 (N_14746,N_10233,N_12383);
xnor U14747 (N_14747,N_10304,N_10776);
or U14748 (N_14748,N_10209,N_10831);
or U14749 (N_14749,N_10412,N_10891);
and U14750 (N_14750,N_12127,N_11863);
nor U14751 (N_14751,N_11115,N_11181);
nor U14752 (N_14752,N_12335,N_10841);
xor U14753 (N_14753,N_10839,N_10711);
or U14754 (N_14754,N_11444,N_11226);
and U14755 (N_14755,N_10992,N_12436);
nor U14756 (N_14756,N_10811,N_11642);
or U14757 (N_14757,N_11855,N_10670);
xnor U14758 (N_14758,N_10461,N_10796);
xnor U14759 (N_14759,N_10959,N_11575);
and U14760 (N_14760,N_10877,N_11999);
nand U14761 (N_14761,N_11747,N_10830);
or U14762 (N_14762,N_11376,N_11584);
or U14763 (N_14763,N_11171,N_10425);
nand U14764 (N_14764,N_11203,N_12153);
and U14765 (N_14765,N_11487,N_12197);
nor U14766 (N_14766,N_10460,N_10811);
or U14767 (N_14767,N_11672,N_11439);
or U14768 (N_14768,N_11172,N_11433);
nand U14769 (N_14769,N_11861,N_12077);
or U14770 (N_14770,N_10090,N_10235);
nand U14771 (N_14771,N_10634,N_12138);
xor U14772 (N_14772,N_11919,N_11523);
xnor U14773 (N_14773,N_10791,N_10035);
or U14774 (N_14774,N_11484,N_10959);
nand U14775 (N_14775,N_11889,N_12431);
nand U14776 (N_14776,N_10564,N_10549);
nor U14777 (N_14777,N_10147,N_11278);
or U14778 (N_14778,N_10817,N_11095);
or U14779 (N_14779,N_10489,N_10496);
nor U14780 (N_14780,N_11348,N_10633);
and U14781 (N_14781,N_11194,N_10736);
and U14782 (N_14782,N_10085,N_10469);
nor U14783 (N_14783,N_10033,N_10891);
nor U14784 (N_14784,N_10269,N_11624);
xor U14785 (N_14785,N_11120,N_11991);
xor U14786 (N_14786,N_12489,N_11300);
nand U14787 (N_14787,N_10298,N_11624);
nor U14788 (N_14788,N_10851,N_10734);
nand U14789 (N_14789,N_10642,N_11207);
xnor U14790 (N_14790,N_10018,N_10471);
xor U14791 (N_14791,N_12229,N_11397);
xor U14792 (N_14792,N_11650,N_10613);
or U14793 (N_14793,N_10588,N_11359);
and U14794 (N_14794,N_12222,N_12424);
nand U14795 (N_14795,N_10025,N_10186);
or U14796 (N_14796,N_12389,N_10994);
or U14797 (N_14797,N_12429,N_10291);
xor U14798 (N_14798,N_12065,N_10966);
xor U14799 (N_14799,N_10513,N_11015);
xor U14800 (N_14800,N_10241,N_11945);
and U14801 (N_14801,N_11675,N_11062);
or U14802 (N_14802,N_10365,N_11796);
and U14803 (N_14803,N_11758,N_11143);
nand U14804 (N_14804,N_11601,N_10971);
nand U14805 (N_14805,N_11359,N_10538);
xnor U14806 (N_14806,N_10973,N_11484);
nand U14807 (N_14807,N_12147,N_10130);
nor U14808 (N_14808,N_10342,N_10196);
or U14809 (N_14809,N_10874,N_11983);
xor U14810 (N_14810,N_11170,N_10456);
or U14811 (N_14811,N_10911,N_11767);
xor U14812 (N_14812,N_10646,N_10507);
or U14813 (N_14813,N_11627,N_10321);
or U14814 (N_14814,N_11357,N_12437);
nor U14815 (N_14815,N_11763,N_11385);
nand U14816 (N_14816,N_12481,N_11294);
or U14817 (N_14817,N_11122,N_11015);
xnor U14818 (N_14818,N_10997,N_12255);
and U14819 (N_14819,N_12400,N_12003);
xnor U14820 (N_14820,N_10174,N_10601);
or U14821 (N_14821,N_10265,N_11710);
nand U14822 (N_14822,N_11997,N_11388);
nor U14823 (N_14823,N_11192,N_11735);
and U14824 (N_14824,N_10196,N_12052);
nand U14825 (N_14825,N_12085,N_11682);
xnor U14826 (N_14826,N_10765,N_10076);
nor U14827 (N_14827,N_11061,N_11810);
nand U14828 (N_14828,N_11601,N_10640);
xnor U14829 (N_14829,N_12261,N_10154);
and U14830 (N_14830,N_11680,N_12373);
xor U14831 (N_14831,N_11939,N_10916);
xor U14832 (N_14832,N_12216,N_11612);
nand U14833 (N_14833,N_11378,N_12061);
nand U14834 (N_14834,N_10642,N_12099);
and U14835 (N_14835,N_11465,N_12136);
nor U14836 (N_14836,N_12250,N_12154);
or U14837 (N_14837,N_10271,N_10259);
xor U14838 (N_14838,N_10413,N_10435);
and U14839 (N_14839,N_10886,N_10782);
xnor U14840 (N_14840,N_12486,N_12017);
xor U14841 (N_14841,N_12311,N_11709);
and U14842 (N_14842,N_11363,N_11611);
and U14843 (N_14843,N_10796,N_11358);
and U14844 (N_14844,N_10052,N_10444);
or U14845 (N_14845,N_10484,N_11711);
xnor U14846 (N_14846,N_10792,N_10901);
nand U14847 (N_14847,N_12029,N_11157);
and U14848 (N_14848,N_12037,N_11968);
nand U14849 (N_14849,N_12252,N_12109);
and U14850 (N_14850,N_11209,N_11045);
and U14851 (N_14851,N_11198,N_10514);
and U14852 (N_14852,N_12341,N_11504);
nor U14853 (N_14853,N_11009,N_11900);
xor U14854 (N_14854,N_11771,N_12465);
xnor U14855 (N_14855,N_10922,N_11419);
nor U14856 (N_14856,N_11096,N_12350);
or U14857 (N_14857,N_12226,N_11333);
nor U14858 (N_14858,N_10643,N_10613);
xnor U14859 (N_14859,N_10486,N_12494);
or U14860 (N_14860,N_10022,N_10463);
nor U14861 (N_14861,N_10697,N_11604);
or U14862 (N_14862,N_12339,N_11352);
and U14863 (N_14863,N_11523,N_11003);
and U14864 (N_14864,N_10436,N_10187);
nor U14865 (N_14865,N_12151,N_11173);
xnor U14866 (N_14866,N_11313,N_11624);
nor U14867 (N_14867,N_12078,N_11642);
or U14868 (N_14868,N_10834,N_11183);
or U14869 (N_14869,N_10871,N_11731);
and U14870 (N_14870,N_10281,N_12456);
xnor U14871 (N_14871,N_12052,N_10242);
nand U14872 (N_14872,N_10100,N_11034);
or U14873 (N_14873,N_12262,N_11049);
xor U14874 (N_14874,N_10960,N_10912);
nor U14875 (N_14875,N_11506,N_10205);
or U14876 (N_14876,N_10548,N_10006);
xor U14877 (N_14877,N_12290,N_10537);
or U14878 (N_14878,N_10319,N_11730);
nand U14879 (N_14879,N_10682,N_11220);
nor U14880 (N_14880,N_11814,N_11601);
nand U14881 (N_14881,N_11670,N_11579);
and U14882 (N_14882,N_10219,N_11203);
or U14883 (N_14883,N_10027,N_11543);
nor U14884 (N_14884,N_11021,N_11168);
or U14885 (N_14885,N_11274,N_10191);
or U14886 (N_14886,N_11948,N_11616);
nand U14887 (N_14887,N_10958,N_11247);
nor U14888 (N_14888,N_11787,N_10072);
xor U14889 (N_14889,N_11545,N_11870);
nand U14890 (N_14890,N_11557,N_10586);
xor U14891 (N_14891,N_11701,N_11482);
xor U14892 (N_14892,N_10449,N_11733);
and U14893 (N_14893,N_10110,N_10261);
xnor U14894 (N_14894,N_11148,N_10625);
nand U14895 (N_14895,N_10179,N_11764);
or U14896 (N_14896,N_12008,N_12155);
nor U14897 (N_14897,N_10186,N_10599);
nand U14898 (N_14898,N_10416,N_10937);
or U14899 (N_14899,N_10461,N_12366);
nor U14900 (N_14900,N_10522,N_10107);
or U14901 (N_14901,N_10479,N_11282);
nand U14902 (N_14902,N_11172,N_10076);
or U14903 (N_14903,N_10239,N_11331);
and U14904 (N_14904,N_12463,N_10091);
and U14905 (N_14905,N_11715,N_12156);
and U14906 (N_14906,N_11268,N_10645);
nand U14907 (N_14907,N_11054,N_11052);
and U14908 (N_14908,N_10064,N_11674);
and U14909 (N_14909,N_11218,N_11478);
and U14910 (N_14910,N_10621,N_10810);
nand U14911 (N_14911,N_10932,N_11809);
and U14912 (N_14912,N_10301,N_12399);
nand U14913 (N_14913,N_12358,N_10349);
xor U14914 (N_14914,N_11674,N_11154);
and U14915 (N_14915,N_12031,N_11141);
nand U14916 (N_14916,N_11483,N_10225);
xor U14917 (N_14917,N_10276,N_12324);
xnor U14918 (N_14918,N_10883,N_11142);
and U14919 (N_14919,N_10865,N_10903);
or U14920 (N_14920,N_11819,N_12252);
nand U14921 (N_14921,N_10090,N_11099);
nor U14922 (N_14922,N_11934,N_10262);
or U14923 (N_14923,N_12272,N_11254);
and U14924 (N_14924,N_10065,N_10241);
and U14925 (N_14925,N_11587,N_11886);
or U14926 (N_14926,N_10817,N_12222);
or U14927 (N_14927,N_12249,N_11956);
or U14928 (N_14928,N_11055,N_12225);
nand U14929 (N_14929,N_11084,N_12313);
nor U14930 (N_14930,N_12413,N_10186);
nand U14931 (N_14931,N_11010,N_12061);
or U14932 (N_14932,N_10084,N_11020);
xnor U14933 (N_14933,N_12484,N_12028);
nand U14934 (N_14934,N_11114,N_11232);
nor U14935 (N_14935,N_10990,N_10880);
nor U14936 (N_14936,N_11834,N_11758);
xor U14937 (N_14937,N_10340,N_11516);
nor U14938 (N_14938,N_10844,N_10766);
nor U14939 (N_14939,N_10177,N_11470);
and U14940 (N_14940,N_10742,N_10624);
and U14941 (N_14941,N_12272,N_11039);
nor U14942 (N_14942,N_10303,N_10893);
nand U14943 (N_14943,N_10527,N_11662);
xor U14944 (N_14944,N_12342,N_12305);
nand U14945 (N_14945,N_10118,N_12144);
xnor U14946 (N_14946,N_12481,N_12164);
nand U14947 (N_14947,N_10794,N_10688);
nand U14948 (N_14948,N_11832,N_11605);
nand U14949 (N_14949,N_11240,N_12439);
or U14950 (N_14950,N_11296,N_12301);
xnor U14951 (N_14951,N_11966,N_11207);
and U14952 (N_14952,N_10886,N_10744);
nand U14953 (N_14953,N_10305,N_10938);
xor U14954 (N_14954,N_10551,N_11041);
and U14955 (N_14955,N_10471,N_10827);
or U14956 (N_14956,N_12338,N_12297);
xor U14957 (N_14957,N_11566,N_10521);
nor U14958 (N_14958,N_12225,N_10841);
xor U14959 (N_14959,N_10051,N_10328);
and U14960 (N_14960,N_11107,N_11580);
xor U14961 (N_14961,N_11795,N_10597);
and U14962 (N_14962,N_11801,N_11211);
nand U14963 (N_14963,N_11777,N_10648);
or U14964 (N_14964,N_10076,N_10323);
or U14965 (N_14965,N_10377,N_10232);
nand U14966 (N_14966,N_11628,N_12272);
xnor U14967 (N_14967,N_11924,N_10583);
and U14968 (N_14968,N_11961,N_11152);
xnor U14969 (N_14969,N_12357,N_11625);
nor U14970 (N_14970,N_11943,N_10468);
or U14971 (N_14971,N_12430,N_12174);
and U14972 (N_14972,N_12329,N_10396);
or U14973 (N_14973,N_11690,N_10811);
nand U14974 (N_14974,N_10540,N_11414);
xor U14975 (N_14975,N_11316,N_11528);
xor U14976 (N_14976,N_11005,N_10408);
nor U14977 (N_14977,N_10025,N_11717);
or U14978 (N_14978,N_12364,N_10930);
nand U14979 (N_14979,N_11567,N_10514);
nor U14980 (N_14980,N_11054,N_12463);
xor U14981 (N_14981,N_10284,N_11760);
or U14982 (N_14982,N_11430,N_11761);
and U14983 (N_14983,N_12446,N_12244);
or U14984 (N_14984,N_11513,N_10455);
xnor U14985 (N_14985,N_11789,N_11166);
nand U14986 (N_14986,N_10956,N_10861);
or U14987 (N_14987,N_12478,N_12195);
and U14988 (N_14988,N_10241,N_12096);
and U14989 (N_14989,N_10119,N_10594);
xnor U14990 (N_14990,N_11213,N_10176);
nor U14991 (N_14991,N_10242,N_11102);
nand U14992 (N_14992,N_12108,N_10803);
nand U14993 (N_14993,N_11137,N_11473);
nor U14994 (N_14994,N_12075,N_12387);
nor U14995 (N_14995,N_11103,N_12239);
xnor U14996 (N_14996,N_12237,N_11659);
xnor U14997 (N_14997,N_11639,N_11719);
and U14998 (N_14998,N_11945,N_10581);
nor U14999 (N_14999,N_10676,N_12348);
nor U15000 (N_15000,N_14817,N_13245);
or U15001 (N_15001,N_12825,N_13725);
nor U15002 (N_15002,N_13110,N_12990);
nor U15003 (N_15003,N_14564,N_14755);
and U15004 (N_15004,N_14391,N_13911);
xor U15005 (N_15005,N_14167,N_14358);
and U15006 (N_15006,N_14542,N_13886);
nand U15007 (N_15007,N_12791,N_14917);
nor U15008 (N_15008,N_13991,N_14856);
nor U15009 (N_15009,N_14614,N_14151);
nor U15010 (N_15010,N_13456,N_13020);
xnor U15011 (N_15011,N_13675,N_14309);
nor U15012 (N_15012,N_13093,N_14387);
nand U15013 (N_15013,N_14348,N_14937);
nor U15014 (N_15014,N_12632,N_13278);
or U15015 (N_15015,N_12555,N_12647);
nor U15016 (N_15016,N_14025,N_14648);
nand U15017 (N_15017,N_13168,N_13510);
nor U15018 (N_15018,N_14770,N_14114);
nand U15019 (N_15019,N_13650,N_14685);
nor U15020 (N_15020,N_14057,N_12787);
nor U15021 (N_15021,N_13274,N_14369);
or U15022 (N_15022,N_13576,N_13430);
nor U15023 (N_15023,N_13363,N_13992);
or U15024 (N_15024,N_14949,N_14950);
or U15025 (N_15025,N_14052,N_13273);
and U15026 (N_15026,N_13705,N_14041);
nand U15027 (N_15027,N_14653,N_14517);
xor U15028 (N_15028,N_12838,N_14735);
xnor U15029 (N_15029,N_13436,N_12640);
or U15030 (N_15030,N_14875,N_13210);
nand U15031 (N_15031,N_13315,N_13328);
xnor U15032 (N_15032,N_12962,N_14142);
or U15033 (N_15033,N_13010,N_12512);
xnor U15034 (N_15034,N_13695,N_14785);
nand U15035 (N_15035,N_13002,N_13798);
nand U15036 (N_15036,N_14488,N_13852);
nor U15037 (N_15037,N_12795,N_13963);
and U15038 (N_15038,N_13643,N_14392);
xnor U15039 (N_15039,N_14959,N_14942);
and U15040 (N_15040,N_14626,N_13302);
nand U15041 (N_15041,N_14760,N_14561);
nand U15042 (N_15042,N_12852,N_14422);
and U15043 (N_15043,N_13387,N_12803);
or U15044 (N_15044,N_12902,N_13803);
nor U15045 (N_15045,N_14809,N_12807);
nor U15046 (N_15046,N_12964,N_12526);
xnor U15047 (N_15047,N_12573,N_14593);
nand U15048 (N_15048,N_13512,N_13945);
and U15049 (N_15049,N_12992,N_14285);
and U15050 (N_15050,N_12592,N_13935);
xnor U15051 (N_15051,N_13007,N_12840);
or U15052 (N_15052,N_14555,N_12725);
nand U15053 (N_15053,N_14427,N_14590);
or U15054 (N_15054,N_12991,N_13413);
nand U15055 (N_15055,N_13636,N_13601);
xor U15056 (N_15056,N_14350,N_14372);
nor U15057 (N_15057,N_12963,N_13897);
xnor U15058 (N_15058,N_14505,N_13174);
nand U15059 (N_15059,N_14191,N_13070);
and U15060 (N_15060,N_13840,N_14676);
or U15061 (N_15061,N_13028,N_12934);
or U15062 (N_15062,N_13600,N_13438);
nand U15063 (N_15063,N_14528,N_14288);
nand U15064 (N_15064,N_13809,N_14076);
xnor U15065 (N_15065,N_13094,N_13022);
or U15066 (N_15066,N_14093,N_13645);
nor U15067 (N_15067,N_12879,N_14107);
or U15068 (N_15068,N_14829,N_14059);
or U15069 (N_15069,N_12843,N_13122);
nand U15070 (N_15070,N_13033,N_14037);
nand U15071 (N_15071,N_13649,N_12811);
nor U15072 (N_15072,N_12846,N_13167);
xnor U15073 (N_15073,N_13810,N_14388);
xnor U15074 (N_15074,N_14174,N_13377);
and U15075 (N_15075,N_14835,N_14644);
nor U15076 (N_15076,N_14603,N_14510);
xnor U15077 (N_15077,N_13147,N_12599);
and U15078 (N_15078,N_14397,N_13773);
nand U15079 (N_15079,N_13637,N_14080);
nand U15080 (N_15080,N_14137,N_13540);
xor U15081 (N_15081,N_14474,N_13763);
or U15082 (N_15082,N_13150,N_14763);
and U15083 (N_15083,N_14814,N_14655);
nor U15084 (N_15084,N_14239,N_13384);
or U15085 (N_15085,N_12862,N_13482);
and U15086 (N_15086,N_14313,N_13907);
nor U15087 (N_15087,N_12643,N_12677);
xor U15088 (N_15088,N_12926,N_14307);
nand U15089 (N_15089,N_13779,N_14342);
and U15090 (N_15090,N_13271,N_14982);
and U15091 (N_15091,N_14922,N_13365);
nor U15092 (N_15092,N_14978,N_12914);
and U15093 (N_15093,N_12808,N_13656);
nand U15094 (N_15094,N_13954,N_12870);
nand U15095 (N_15095,N_14839,N_13348);
nor U15096 (N_15096,N_13241,N_12530);
and U15097 (N_15097,N_12684,N_13104);
xor U15098 (N_15098,N_13874,N_13934);
nor U15099 (N_15099,N_12998,N_13206);
or U15100 (N_15100,N_12804,N_13074);
nor U15101 (N_15101,N_14182,N_14659);
and U15102 (N_15102,N_14617,N_13362);
xnor U15103 (N_15103,N_13865,N_13190);
xnor U15104 (N_15104,N_12777,N_14781);
xnor U15105 (N_15105,N_12924,N_14708);
nand U15106 (N_15106,N_14640,N_14206);
nand U15107 (N_15107,N_14019,N_14627);
nor U15108 (N_15108,N_14103,N_14531);
xor U15109 (N_15109,N_14747,N_14563);
or U15110 (N_15110,N_14975,N_12732);
and U15111 (N_15111,N_13966,N_13528);
nand U15112 (N_15112,N_14165,N_12799);
xnor U15113 (N_15113,N_13744,N_14901);
nand U15114 (N_15114,N_13754,N_13192);
and U15115 (N_15115,N_12848,N_14226);
and U15116 (N_15116,N_12989,N_14569);
nor U15117 (N_15117,N_14273,N_12661);
xor U15118 (N_15118,N_14078,N_12539);
and U15119 (N_15119,N_14988,N_13057);
nor U15120 (N_15120,N_12976,N_12501);
and U15121 (N_15121,N_13898,N_13633);
nand U15122 (N_15122,N_12669,N_13502);
or U15123 (N_15123,N_12778,N_12549);
or U15124 (N_15124,N_13667,N_13938);
nor U15125 (N_15125,N_14144,N_12679);
nor U15126 (N_15126,N_13702,N_12744);
nor U15127 (N_15127,N_13679,N_13193);
xor U15128 (N_15128,N_12750,N_14652);
nor U15129 (N_15129,N_13125,N_13855);
nand U15130 (N_15130,N_12953,N_14623);
xnor U15131 (N_15131,N_14434,N_12961);
xor U15132 (N_15132,N_14301,N_13509);
nor U15133 (N_15133,N_13352,N_14331);
xor U15134 (N_15134,N_14845,N_14351);
xor U15135 (N_15135,N_13771,N_12940);
or U15136 (N_15136,N_14155,N_14981);
nand U15137 (N_15137,N_12701,N_13381);
and U15138 (N_15138,N_14258,N_13928);
and U15139 (N_15139,N_14501,N_13550);
xor U15140 (N_15140,N_12568,N_13851);
nand U15141 (N_15141,N_13914,N_14106);
or U15142 (N_15142,N_14536,N_13979);
and U15143 (N_15143,N_13000,N_12614);
or U15144 (N_15144,N_13857,N_12529);
and U15145 (N_15145,N_13757,N_12663);
nor U15146 (N_15146,N_14046,N_12800);
and U15147 (N_15147,N_14083,N_14240);
xnor U15148 (N_15148,N_13516,N_12812);
or U15149 (N_15149,N_13358,N_13040);
nand U15150 (N_15150,N_14376,N_13390);
xnor U15151 (N_15151,N_12749,N_13506);
nor U15152 (N_15152,N_14218,N_12896);
and U15153 (N_15153,N_13339,N_12875);
and U15154 (N_15154,N_14838,N_14896);
or U15155 (N_15155,N_14112,N_14912);
or U15156 (N_15156,N_12809,N_13998);
nand U15157 (N_15157,N_13681,N_14671);
xnor U15158 (N_15158,N_14525,N_14400);
nor U15159 (N_15159,N_13715,N_14780);
nor U15160 (N_15160,N_13095,N_13969);
and U15161 (N_15161,N_14360,N_13156);
xnor U15162 (N_15162,N_12915,N_13776);
and U15163 (N_15163,N_14330,N_13762);
nand U15164 (N_15164,N_12815,N_12967);
nor U15165 (N_15165,N_13335,N_12721);
or U15166 (N_15166,N_12642,N_13831);
nand U15167 (N_15167,N_13149,N_13234);
nand U15168 (N_15168,N_14911,N_13838);
nor U15169 (N_15169,N_13217,N_12514);
nand U15170 (N_15170,N_13049,N_14418);
nand U15171 (N_15171,N_12925,N_14314);
and U15172 (N_15172,N_13414,N_13289);
or U15173 (N_15173,N_13565,N_13366);
xor U15174 (N_15174,N_13951,N_12861);
xnor U15175 (N_15175,N_14872,N_14003);
and U15176 (N_15176,N_14308,N_14722);
nand U15177 (N_15177,N_12520,N_14195);
xor U15178 (N_15178,N_13918,N_14677);
xor U15179 (N_15179,N_13005,N_13740);
or U15180 (N_15180,N_14599,N_14819);
or U15181 (N_15181,N_14731,N_12880);
nand U15182 (N_15182,N_14322,N_14327);
xor U15183 (N_15183,N_14030,N_14605);
xor U15184 (N_15184,N_14175,N_12891);
nor U15185 (N_15185,N_13747,N_12888);
or U15186 (N_15186,N_12935,N_14633);
and U15187 (N_15187,N_14664,N_14320);
xnor U15188 (N_15188,N_14932,N_14415);
nand U15189 (N_15189,N_13140,N_14183);
xnor U15190 (N_15190,N_14936,N_13367);
and U15191 (N_15191,N_13356,N_14197);
nor U15192 (N_15192,N_12923,N_13662);
xor U15193 (N_15193,N_14656,N_13548);
and U15194 (N_15194,N_13614,N_14717);
and U15195 (N_15195,N_14340,N_14328);
or U15196 (N_15196,N_13325,N_13825);
nand U15197 (N_15197,N_13562,N_13087);
xnor U15198 (N_15198,N_14702,N_14053);
xnor U15199 (N_15199,N_12575,N_12798);
xor U15200 (N_15200,N_13890,N_13625);
and U15201 (N_15201,N_14004,N_12823);
nand U15202 (N_15202,N_13448,N_12546);
and U15203 (N_15203,N_13863,N_13257);
and U15204 (N_15204,N_13287,N_14892);
nor U15205 (N_15205,N_12897,N_13472);
and U15206 (N_15206,N_13872,N_13980);
or U15207 (N_15207,N_12850,N_12841);
nor U15208 (N_15208,N_14798,N_14454);
and U15209 (N_15209,N_13262,N_13652);
xor U15210 (N_15210,N_13485,N_14259);
xor U15211 (N_15211,N_14598,N_14084);
or U15212 (N_15212,N_14668,N_13745);
nor U15213 (N_15213,N_13220,N_14050);
nand U15214 (N_15214,N_13698,N_14442);
nand U15215 (N_15215,N_13144,N_14549);
nand U15216 (N_15216,N_14907,N_14205);
xor U15217 (N_15217,N_13988,N_13768);
nor U15218 (N_15218,N_14486,N_13973);
or U15219 (N_15219,N_12824,N_12782);
nor U15220 (N_15220,N_12541,N_13568);
or U15221 (N_15221,N_14766,N_13431);
or U15222 (N_15222,N_13975,N_14545);
or U15223 (N_15223,N_14271,N_12780);
or U15224 (N_15224,N_14190,N_14077);
xnor U15225 (N_15225,N_13101,N_12927);
or U15226 (N_15226,N_14778,N_13690);
nor U15227 (N_15227,N_13329,N_12607);
and U15228 (N_15228,N_14222,N_14484);
and U15229 (N_15229,N_13183,N_14576);
xnor U15230 (N_15230,N_13739,N_13232);
or U15231 (N_15231,N_13917,N_13288);
nor U15232 (N_15232,N_13466,N_14877);
xnor U15233 (N_15233,N_12973,N_14544);
or U15234 (N_15234,N_13561,N_13617);
nor U15235 (N_15235,N_14746,N_14022);
xor U15236 (N_15236,N_13444,N_13496);
nand U15237 (N_15237,N_14768,N_14807);
or U15238 (N_15238,N_13292,N_14296);
or U15239 (N_15239,N_13296,N_14699);
and U15240 (N_15240,N_14674,N_14177);
nor U15241 (N_15241,N_13378,N_13457);
and U15242 (N_15242,N_14927,N_13107);
nand U15243 (N_15243,N_12689,N_13549);
or U15244 (N_15244,N_14058,N_14697);
or U15245 (N_15245,N_14629,N_13249);
nor U15246 (N_15246,N_14591,N_14141);
or U15247 (N_15247,N_14503,N_13483);
nor U15248 (N_15248,N_12877,N_12613);
and U15249 (N_15249,N_14738,N_14812);
nor U15250 (N_15250,N_14450,N_12887);
and U15251 (N_15251,N_14694,N_14213);
nor U15252 (N_15252,N_12566,N_12601);
and U15253 (N_15253,N_14943,N_14249);
nor U15254 (N_15254,N_13090,N_13470);
and U15255 (N_15255,N_12506,N_12866);
nor U15256 (N_15256,N_13169,N_13712);
and U15257 (N_15257,N_14231,N_13597);
nand U15258 (N_15258,N_13760,N_13950);
or U15259 (N_15259,N_13654,N_14416);
nor U15260 (N_15260,N_14111,N_14235);
xnor U15261 (N_15261,N_14681,N_14577);
nor U15262 (N_15262,N_13326,N_14169);
nand U15263 (N_15263,N_14775,N_13442);
or U15264 (N_15264,N_13808,N_14361);
and U15265 (N_15265,N_14963,N_13513);
nor U15266 (N_15266,N_14009,N_13233);
or U15267 (N_15267,N_13282,N_14651);
nand U15268 (N_15268,N_12633,N_13259);
and U15269 (N_15269,N_13931,N_14396);
nand U15270 (N_15270,N_14601,N_13981);
and U15271 (N_15271,N_14029,N_13011);
xnor U15272 (N_15272,N_13566,N_14749);
nor U15273 (N_15273,N_13788,N_13400);
nand U15274 (N_15274,N_14366,N_13626);
and U15275 (N_15275,N_13563,N_14362);
nor U15276 (N_15276,N_14344,N_13422);
nand U15277 (N_15277,N_14324,N_12708);
nand U15278 (N_15278,N_14667,N_12584);
nand U15279 (N_15279,N_14700,N_14507);
xor U15280 (N_15280,N_13465,N_14953);
nor U15281 (N_15281,N_12569,N_14414);
nand U15282 (N_15282,N_13867,N_13610);
and U15283 (N_15283,N_13923,N_13799);
nand U15284 (N_15284,N_13277,N_14118);
nor U15285 (N_15285,N_12820,N_13364);
xnor U15286 (N_15286,N_14184,N_13284);
xnor U15287 (N_15287,N_14909,N_13678);
nand U15288 (N_15288,N_13404,N_14508);
nand U15289 (N_15289,N_14933,N_12638);
nor U15290 (N_15290,N_13162,N_14830);
xor U15291 (N_15291,N_14200,N_13130);
nand U15292 (N_15292,N_13639,N_12975);
nand U15293 (N_15293,N_12667,N_13211);
xnor U15294 (N_15294,N_13463,N_13571);
and U15295 (N_15295,N_14595,N_14419);
and U15296 (N_15296,N_12564,N_13629);
xnor U15297 (N_15297,N_13572,N_14456);
xnor U15298 (N_15298,N_14773,N_14121);
or U15299 (N_15299,N_13298,N_13632);
nand U15300 (N_15300,N_14161,N_14295);
xnor U15301 (N_15301,N_14672,N_13786);
or U15302 (N_15302,N_14005,N_14990);
or U15303 (N_15303,N_13059,N_14862);
nor U15304 (N_15304,N_12772,N_14039);
nand U15305 (N_15305,N_13882,N_14583);
and U15306 (N_15306,N_14045,N_13878);
and U15307 (N_15307,N_14945,N_13276);
and U15308 (N_15308,N_14269,N_14997);
nor U15309 (N_15309,N_13062,N_13052);
xor U15310 (N_15310,N_13916,N_13620);
nor U15311 (N_15311,N_12785,N_12648);
nand U15312 (N_15312,N_14357,N_12929);
nor U15313 (N_15313,N_13962,N_12695);
or U15314 (N_15314,N_13896,N_14256);
nand U15315 (N_15315,N_14704,N_13114);
or U15316 (N_15316,N_13589,N_13006);
or U15317 (N_15317,N_14712,N_13098);
or U15318 (N_15318,N_14551,N_12646);
nor U15319 (N_15319,N_14958,N_12857);
nor U15320 (N_15320,N_12965,N_13323);
nor U15321 (N_15321,N_13295,N_14759);
nand U15322 (N_15322,N_13957,N_14794);
or U15323 (N_15323,N_13354,N_13802);
nor U15324 (N_15324,N_12682,N_12637);
or U15325 (N_15325,N_14663,N_12715);
or U15326 (N_15326,N_14018,N_14148);
and U15327 (N_15327,N_14102,N_13375);
xnor U15328 (N_15328,N_13688,N_14512);
nor U15329 (N_15329,N_12666,N_14745);
nor U15330 (N_15330,N_14173,N_13453);
xnor U15331 (N_15331,N_14834,N_14268);
xor U15332 (N_15332,N_13504,N_13489);
or U15333 (N_15333,N_14015,N_14618);
nor U15334 (N_15334,N_13887,N_13359);
nor U15335 (N_15335,N_14534,N_14497);
nor U15336 (N_15336,N_13944,N_13791);
and U15337 (N_15337,N_13447,N_14686);
nand U15338 (N_15338,N_14247,N_13205);
xor U15339 (N_15339,N_14385,N_13519);
nor U15340 (N_15340,N_13286,N_14333);
xor U15341 (N_15341,N_12507,N_12656);
or U15342 (N_15342,N_13214,N_14062);
and U15343 (N_15343,N_13397,N_13783);
nand U15344 (N_15344,N_13959,N_13929);
nor U15345 (N_15345,N_13816,N_13642);
nor U15346 (N_15346,N_14260,N_12768);
or U15347 (N_15347,N_12634,N_12955);
and U15348 (N_15348,N_13586,N_14441);
nand U15349 (N_15349,N_12504,N_14675);
or U15350 (N_15350,N_13396,N_12733);
nor U15351 (N_15351,N_12687,N_12776);
nand U15352 (N_15352,N_13733,N_12605);
xnor U15353 (N_15353,N_13829,N_12922);
and U15354 (N_15354,N_12892,N_12793);
nor U15355 (N_15355,N_12884,N_14607);
nand U15356 (N_15356,N_14783,N_13987);
nor U15357 (N_15357,N_13738,N_14225);
and U15358 (N_15358,N_13848,N_12672);
nor U15359 (N_15359,N_14998,N_14924);
nand U15360 (N_15360,N_14880,N_14624);
or U15361 (N_15361,N_13388,N_12931);
nor U15362 (N_15362,N_13879,N_13570);
xnor U15363 (N_15363,N_14034,N_12619);
nand U15364 (N_15364,N_13860,N_14619);
xor U15365 (N_15365,N_14522,N_14606);
nor U15366 (N_15366,N_14223,N_12654);
or U15367 (N_15367,N_12872,N_12783);
nand U15368 (N_15368,N_14787,N_12510);
nand U15369 (N_15369,N_12794,N_13053);
nand U15370 (N_15370,N_14261,N_12760);
nand U15371 (N_15371,N_12538,N_14264);
xnor U15372 (N_15372,N_12860,N_12999);
nand U15373 (N_15373,N_14138,N_14831);
nand U15374 (N_15374,N_13569,N_14451);
nand U15375 (N_15375,N_13534,N_13143);
and U15376 (N_15376,N_14283,N_13047);
and U15377 (N_15377,N_14902,N_14289);
xnor U15378 (N_15378,N_13801,N_12664);
and U15379 (N_15379,N_13452,N_13921);
nor U15380 (N_15380,N_13699,N_13612);
or U15381 (N_15381,N_13955,N_13399);
xnor U15382 (N_15382,N_13846,N_13189);
or U15383 (N_15383,N_13064,N_14002);
nand U15384 (N_15384,N_12545,N_13408);
and U15385 (N_15385,N_14498,N_12580);
nand U15386 (N_15386,N_12690,N_14756);
and U15387 (N_15387,N_13839,N_14297);
xnor U15388 (N_15388,N_13332,N_12868);
and U15389 (N_15389,N_14961,N_12737);
xor U15390 (N_15390,N_14820,N_12764);
and U15391 (N_15391,N_14769,N_13417);
or U15392 (N_15392,N_14262,N_14666);
and U15393 (N_15393,N_13235,N_14394);
nand U15394 (N_15394,N_13297,N_13869);
and U15395 (N_15395,N_13824,N_13222);
and U15396 (N_15396,N_14075,N_13229);
and U15397 (N_15397,N_14305,N_13487);
or U15398 (N_15398,N_13729,N_12842);
nor U15399 (N_15399,N_14691,N_14615);
or U15400 (N_15400,N_14381,N_12641);
nor U15401 (N_15401,N_13596,N_13054);
nor U15402 (N_15402,N_12770,N_14719);
or U15403 (N_15403,N_14854,N_13529);
nand U15404 (N_15404,N_13434,N_13238);
nor U15405 (N_15405,N_12618,N_13443);
and U15406 (N_15406,N_13673,N_14635);
nand U15407 (N_15407,N_14196,N_13781);
xnor U15408 (N_15408,N_13451,N_14424);
and U15409 (N_15409,N_14841,N_14302);
xor U15410 (N_15410,N_14580,N_12711);
and U15411 (N_15411,N_14444,N_13065);
or U15412 (N_15412,N_13027,N_13480);
nor U15413 (N_15413,N_12797,N_14293);
nand U15414 (N_15414,N_14801,N_14791);
nor U15415 (N_15415,N_14962,N_13713);
xor U15416 (N_15416,N_12628,N_12578);
or U15417 (N_15417,N_12600,N_12644);
nand U15418 (N_15418,N_14670,N_13337);
or U15419 (N_15419,N_14405,N_13379);
nor U15420 (N_15420,N_13926,N_14947);
or U15421 (N_15421,N_13710,N_14752);
xnor U15422 (N_15422,N_12984,N_14941);
nor U15423 (N_15423,N_14224,N_12660);
nor U15424 (N_15424,N_12900,N_12767);
or U15425 (N_15425,N_13248,N_14837);
nor U15426 (N_15426,N_13701,N_13728);
nor U15427 (N_15427,N_14478,N_13511);
or U15428 (N_15428,N_13197,N_13903);
or U15429 (N_15429,N_14504,N_13009);
nand U15430 (N_15430,N_13243,N_13063);
nor U15431 (N_15431,N_14439,N_13208);
and U15432 (N_15432,N_14395,N_14960);
and U15433 (N_15433,N_12920,N_13421);
and U15434 (N_15434,N_13254,N_14382);
nand U15435 (N_15435,N_14900,N_14879);
nor U15436 (N_15436,N_14281,N_14566);
and U15437 (N_15437,N_14219,N_13674);
nand U15438 (N_15438,N_14007,N_14951);
nand U15439 (N_15439,N_12942,N_12959);
and U15440 (N_15440,N_13411,N_14412);
nor U15441 (N_15441,N_14379,N_14984);
xnor U15442 (N_15442,N_13163,N_13968);
or U15443 (N_15443,N_14094,N_14110);
xnor U15444 (N_15444,N_12761,N_13567);
xnor U15445 (N_15445,N_13909,N_14915);
and U15446 (N_15446,N_12971,N_14012);
and U15447 (N_15447,N_14091,N_13503);
nor U15448 (N_15448,N_14557,N_14568);
or U15449 (N_15449,N_14952,N_13983);
or U15450 (N_15450,N_13305,N_12859);
or U15451 (N_15451,N_13460,N_14524);
nand U15452 (N_15452,N_12944,N_12528);
or U15453 (N_15453,N_13361,N_14625);
nor U15454 (N_15454,N_12645,N_14466);
nor U15455 (N_15455,N_13306,N_13283);
xnor U15456 (N_15456,N_12518,N_14669);
xnor U15457 (N_15457,N_12784,N_12517);
nand U15458 (N_15458,N_12565,N_14300);
xor U15459 (N_15459,N_12949,N_14447);
and U15460 (N_15460,N_14399,N_12622);
nand U15461 (N_15461,N_13317,N_14554);
and U15462 (N_15462,N_12719,N_13796);
nand U15463 (N_15463,N_14426,N_13355);
nand U15464 (N_15464,N_12542,N_12853);
nor U15465 (N_15465,N_13575,N_13307);
nor U15466 (N_15466,N_12769,N_14526);
nor U15467 (N_15467,N_13251,N_14716);
xor U15468 (N_15468,N_14733,N_12736);
xor U15469 (N_15469,N_14898,N_14847);
xnor U15470 (N_15470,N_14082,N_14265);
and U15471 (N_15471,N_13066,N_13327);
or U15472 (N_15472,N_14567,N_14122);
xnor U15473 (N_15473,N_14168,N_13386);
xnor U15474 (N_15474,N_12593,N_14597);
nor U15475 (N_15475,N_13079,N_12864);
and U15476 (N_15476,N_14253,N_14788);
or U15477 (N_15477,N_14095,N_12839);
nor U15478 (N_15478,N_12835,N_14024);
nand U15479 (N_15479,N_14767,N_13014);
xor U15480 (N_15480,N_13170,N_13398);
xor U15481 (N_15481,N_12818,N_13180);
nor U15482 (N_15482,N_12571,N_14693);
and U15483 (N_15483,N_13461,N_14139);
nor U15484 (N_15484,N_13313,N_13797);
or U15485 (N_15485,N_13994,N_13644);
or U15486 (N_15486,N_13624,N_14529);
nand U15487 (N_15487,N_13209,N_14765);
nor U15488 (N_15488,N_14060,N_13737);
or U15489 (N_15489,N_13578,N_12729);
nor U15490 (N_15490,N_14199,N_14085);
nor U15491 (N_15491,N_13850,N_12854);
or U15492 (N_15492,N_13015,N_13322);
nor U15493 (N_15493,N_14446,N_12983);
or U15494 (N_15494,N_14539,N_14463);
nor U15495 (N_15495,N_12678,N_13160);
or U15496 (N_15496,N_14806,N_12674);
xnor U15497 (N_15497,N_12805,N_14824);
and U15498 (N_15498,N_14968,N_13403);
or U15499 (N_15499,N_14680,N_14616);
and U15500 (N_15500,N_12710,N_13603);
and U15501 (N_15501,N_13227,N_12893);
or U15502 (N_15502,N_14800,N_13727);
xor U15503 (N_15503,N_14345,N_14521);
xor U15504 (N_15504,N_13056,N_13515);
and U15505 (N_15505,N_14572,N_13552);
nand U15506 (N_15506,N_14126,N_14489);
or U15507 (N_15507,N_13201,N_14011);
nand U15508 (N_15508,N_14565,N_14483);
nor U15509 (N_15509,N_14688,N_12617);
nor U15510 (N_15510,N_14695,N_12537);
nand U15511 (N_15511,N_14860,N_14732);
nor U15512 (N_15512,N_14548,N_13591);
and U15513 (N_15513,N_14378,N_12834);
nand U15514 (N_15514,N_14910,N_14753);
or U15515 (N_15515,N_12814,N_12722);
or U15516 (N_15516,N_13123,N_12692);
and U15517 (N_15517,N_13230,N_14202);
xor U15518 (N_15518,N_14355,N_13657);
nand U15519 (N_15519,N_13141,N_13097);
nor U15520 (N_15520,N_14411,N_12620);
nor U15521 (N_15521,N_14125,N_14596);
or U15522 (N_15522,N_13216,N_14401);
and U15523 (N_15523,N_14027,N_12553);
and U15524 (N_15524,N_14304,N_12740);
xor U15525 (N_15525,N_14180,N_12911);
xnor U15526 (N_15526,N_12548,N_13309);
or U15527 (N_15527,N_13684,N_14163);
xnor U15528 (N_15528,N_12958,N_14208);
nand U15529 (N_15529,N_13228,N_13412);
or U15530 (N_15530,N_13105,N_13767);
or U15531 (N_15531,N_14276,N_14147);
nor U15532 (N_15532,N_13545,N_14101);
or U15533 (N_15533,N_12581,N_14889);
and U15534 (N_15534,N_14589,N_13429);
and U15535 (N_15535,N_12594,N_13357);
xor U15536 (N_15536,N_14725,N_13039);
nand U15537 (N_15537,N_14220,N_12806);
nand U15538 (N_15538,N_13401,N_13419);
nor U15539 (N_15539,N_14825,N_14108);
and U15540 (N_15540,N_12844,N_13806);
nor U15541 (N_15541,N_14876,N_14294);
xor U15542 (N_15542,N_13708,N_13560);
nand U15543 (N_15543,N_12603,N_14171);
nor U15544 (N_15544,N_13577,N_13360);
nand U15545 (N_15545,N_14238,N_12788);
and U15546 (N_15546,N_13320,N_14021);
and U15547 (N_15547,N_14146,N_13137);
nor U15548 (N_15548,N_14727,N_13300);
nand U15549 (N_15549,N_13743,N_14852);
nand U15550 (N_15550,N_14865,N_12883);
xor U15551 (N_15551,N_13664,N_13615);
nor U15552 (N_15552,N_13659,N_13118);
xnor U15553 (N_15553,N_14518,N_14443);
nor U15554 (N_15554,N_13524,N_14423);
or U15555 (N_15555,N_12558,N_13099);
or U15556 (N_15556,N_13269,N_13126);
nor U15557 (N_15557,N_12757,N_13016);
nor U15558 (N_15558,N_13961,N_14437);
nand U15559 (N_15559,N_14067,N_13814);
nor U15560 (N_15560,N_14374,N_14178);
or U15561 (N_15561,N_14464,N_12602);
nor U15562 (N_15562,N_13374,N_13580);
nor U15563 (N_15563,N_13541,N_13038);
xnor U15564 (N_15564,N_14858,N_13731);
xor U15565 (N_15565,N_14632,N_14291);
or U15566 (N_15566,N_14864,N_14543);
xor U15567 (N_15567,N_12979,N_12511);
xnor U15568 (N_15568,N_14509,N_13158);
or U15569 (N_15569,N_14185,N_13389);
xnor U15570 (N_15570,N_12681,N_13556);
nor U15571 (N_15571,N_14552,N_12630);
nand U15572 (N_15572,N_14347,N_13693);
xnor U15573 (N_15573,N_12826,N_13507);
and U15574 (N_15574,N_12635,N_13559);
and U15575 (N_15575,N_14332,N_14429);
xnor U15576 (N_15576,N_14919,N_14246);
nor U15577 (N_15577,N_13520,N_14459);
and U15578 (N_15578,N_12574,N_12615);
or U15579 (N_15579,N_13252,N_12588);
or U15580 (N_15580,N_14319,N_13191);
nor U15581 (N_15581,N_13514,N_13653);
xor U15582 (N_15582,N_12702,N_13943);
nand U15583 (N_15583,N_13686,N_12762);
and U15584 (N_15584,N_14194,N_13523);
xor U15585 (N_15585,N_13266,N_13347);
or U15586 (N_15586,N_13427,N_14696);
and U15587 (N_15587,N_14636,N_14530);
nand U15588 (N_15588,N_14315,N_14377);
xnor U15589 (N_15589,N_12981,N_14863);
nor U15590 (N_15590,N_13179,N_14709);
nand U15591 (N_15591,N_13058,N_13888);
xnor U15592 (N_15592,N_12847,N_13018);
or U15593 (N_15593,N_14040,N_12986);
or U15594 (N_15594,N_13815,N_13807);
nand U15595 (N_15595,N_13308,N_14861);
or U15596 (N_15596,N_13665,N_13402);
nand U15597 (N_15597,N_14744,N_13368);
and U15598 (N_15598,N_14871,N_14848);
xor U15599 (N_15599,N_13135,N_14006);
nor U15600 (N_15600,N_13184,N_12727);
nand U15601 (N_15601,N_13486,N_14895);
xnor U15602 (N_15602,N_14365,N_12587);
xor U15603 (N_15603,N_12680,N_13820);
or U15604 (N_15604,N_14255,N_14560);
xor U15605 (N_15605,N_13742,N_13242);
or U15606 (N_15606,N_13493,N_13630);
nand U15607 (N_15607,N_13083,N_14639);
or U15608 (N_15608,N_14939,N_12629);
xnor U15609 (N_15609,N_14683,N_13061);
nand U15610 (N_15610,N_13108,N_13003);
xnor U15611 (N_15611,N_13984,N_13905);
nand U15612 (N_15612,N_14349,N_13155);
and U15613 (N_15613,N_13818,N_14066);
or U15614 (N_15614,N_12724,N_13611);
or U15615 (N_15615,N_13045,N_12707);
and U15616 (N_15616,N_13085,N_12966);
xor U15617 (N_15617,N_14983,N_14609);
nor U15618 (N_15618,N_13758,N_13299);
nor U15619 (N_15619,N_14430,N_14948);
or U15620 (N_15620,N_14380,N_14410);
and U15621 (N_15621,N_13314,N_12505);
and U15622 (N_15622,N_13634,N_13175);
or U15623 (N_15623,N_14516,N_13416);
nand U15624 (N_15624,N_13978,N_14383);
xor U15625 (N_15625,N_13606,N_12941);
or U15626 (N_15626,N_12856,N_13948);
and U15627 (N_15627,N_13112,N_13330);
and U15628 (N_15628,N_14134,N_13500);
and U15629 (N_15629,N_13598,N_14229);
xor U15630 (N_15630,N_14154,N_14730);
and U15631 (N_15631,N_14570,N_14634);
nand U15632 (N_15632,N_13640,N_13718);
or U15633 (N_15633,N_14908,N_14428);
xnor U15634 (N_15634,N_14771,N_14657);
nand U15635 (N_15635,N_13680,N_13247);
nand U15636 (N_15636,N_13004,N_14461);
and U15637 (N_15637,N_14527,N_13393);
nand U15638 (N_15638,N_14808,N_13426);
xor U15639 (N_15639,N_13468,N_13445);
and U15640 (N_15640,N_13720,N_13331);
nor U15641 (N_15641,N_12570,N_14048);
nor U15642 (N_15642,N_14237,N_13789);
nand U15643 (N_15643,N_12899,N_14162);
xor U15644 (N_15644,N_12703,N_13215);
nand U15645 (N_15645,N_12616,N_14757);
nand U15646 (N_15646,N_14017,N_14967);
and U15647 (N_15647,N_12822,N_13953);
or U15648 (N_15648,N_12916,N_13602);
xnor U15649 (N_15649,N_12651,N_13391);
nand U15650 (N_15650,N_12693,N_13925);
xnor U15651 (N_15651,N_14925,N_12543);
xor U15652 (N_15652,N_12921,N_13106);
and U15653 (N_15653,N_13986,N_13076);
xnor U15654 (N_15654,N_13272,N_14187);
xnor U15655 (N_15655,N_13078,N_12882);
nand U15656 (N_15656,N_12746,N_13410);
nor U15657 (N_15657,N_13794,N_14792);
and U15658 (N_15658,N_14353,N_13711);
and U15659 (N_15659,N_14310,N_14203);
or U15660 (N_15660,N_13830,N_14940);
and U15661 (N_15661,N_13035,N_14514);
and U15662 (N_15662,N_13102,N_12755);
nand U15663 (N_15663,N_14119,N_13187);
and U15664 (N_15664,N_14851,N_13342);
and U15665 (N_15665,N_14575,N_14460);
or U15666 (N_15666,N_13912,N_13164);
nor U15667 (N_15667,N_13225,N_12903);
nor U15668 (N_15668,N_13902,N_14602);
nor U15669 (N_15669,N_12625,N_13996);
xnor U15670 (N_15670,N_13660,N_13333);
nor U15671 (N_15671,N_13392,N_13581);
and U15672 (N_15672,N_14097,N_14179);
nand U15673 (N_15673,N_13594,N_12502);
or U15674 (N_15674,N_14957,N_12572);
or U15675 (N_15675,N_14475,N_14023);
xnor U15676 (N_15676,N_13042,N_14881);
nand U15677 (N_15677,N_14592,N_14893);
nand U15678 (N_15678,N_13281,N_13697);
nor U15679 (N_15679,N_14089,N_14087);
xnor U15680 (N_15680,N_14016,N_12996);
xnor U15681 (N_15681,N_13861,N_13748);
and U15682 (N_15682,N_14465,N_13584);
and U15683 (N_15683,N_13780,N_13304);
and U15684 (N_15684,N_13692,N_13942);
nor U15685 (N_15685,N_13476,N_13089);
and U15686 (N_15686,N_12738,N_14390);
or U15687 (N_15687,N_14649,N_14645);
nor U15688 (N_15688,N_14887,N_12943);
xor U15689 (N_15689,N_13756,N_12816);
nor U15690 (N_15690,N_14986,N_13420);
or U15691 (N_15691,N_14329,N_13769);
nand U15692 (N_15692,N_13025,N_13345);
and U15693 (N_15693,N_14499,N_12658);
xnor U15694 (N_15694,N_14726,N_14217);
nor U15695 (N_15695,N_14540,N_14043);
and U15696 (N_15696,N_14425,N_14316);
or U15697 (N_15697,N_13464,N_13293);
or U15698 (N_15698,N_13477,N_12985);
nand U15699 (N_15699,N_13341,N_14128);
nand U15700 (N_15700,N_14888,N_14720);
nor U15701 (N_15701,N_14152,N_14044);
nor U15702 (N_15702,N_14481,N_14317);
nor U15703 (N_15703,N_13256,N_13075);
nand U15704 (N_15704,N_13224,N_13689);
or U15705 (N_15705,N_13877,N_14248);
or U15706 (N_15706,N_12906,N_12751);
nor U15707 (N_15707,N_12889,N_12956);
and U15708 (N_15708,N_14113,N_14176);
nor U15709 (N_15709,N_12714,N_14257);
nor U15710 (N_15710,N_14263,N_12586);
or U15711 (N_15711,N_14153,N_12775);
and U15712 (N_15712,N_12686,N_12904);
and U15713 (N_15713,N_12536,N_13974);
xor U15714 (N_15714,N_13406,N_13812);
nand U15715 (N_15715,N_14761,N_14207);
or U15716 (N_15716,N_13736,N_13670);
or U15717 (N_15717,N_14492,N_14684);
xor U15718 (N_15718,N_14104,N_12609);
or U15719 (N_15719,N_14407,N_12867);
nand U15720 (N_15720,N_14306,N_13995);
or U15721 (N_15721,N_14064,N_13832);
nand U15722 (N_15722,N_13826,N_13709);
and U15723 (N_15723,N_14440,N_13318);
and U15724 (N_15724,N_13795,N_13685);
xor U15725 (N_15725,N_14406,N_13704);
nand U15726 (N_15726,N_14493,N_12726);
xor U15727 (N_15727,N_13219,N_13439);
and U15728 (N_15728,N_13275,N_12972);
xnor U15729 (N_15729,N_13312,N_13765);
or U15730 (N_15730,N_14335,N_13424);
and U15731 (N_15731,N_12781,N_14855);
nor U15732 (N_15732,N_14193,N_13165);
nand U15733 (N_15733,N_14286,N_14679);
nor U15734 (N_15734,N_13121,N_14650);
nand U15735 (N_15735,N_14964,N_12525);
or U15736 (N_15736,N_12773,N_14711);
and U15737 (N_15737,N_13231,N_13949);
nand U15738 (N_15738,N_12865,N_13924);
or U15739 (N_15739,N_12522,N_14124);
and U15740 (N_15740,N_14748,N_13428);
or U15741 (N_15741,N_14170,N_12718);
and U15742 (N_15742,N_12688,N_12551);
nor U15743 (N_15743,N_12562,N_13450);
xor U15744 (N_15744,N_14689,N_12556);
xor U15745 (N_15745,N_12662,N_14928);
or U15746 (N_15746,N_12779,N_12547);
nor U15747 (N_15747,N_13423,N_14063);
or U15748 (N_15748,N_12871,N_14127);
nand U15749 (N_15749,N_12938,N_14799);
nor U15750 (N_15750,N_14638,N_12516);
nor U15751 (N_15751,N_13285,N_13997);
or U15752 (N_15752,N_13590,N_13092);
nor U15753 (N_15753,N_12735,N_13041);
nand U15754 (N_15754,N_13048,N_14776);
xor U15755 (N_15755,N_14364,N_13956);
or U15756 (N_15756,N_13870,N_12917);
and U15757 (N_15757,N_13989,N_12621);
or U15758 (N_15758,N_14622,N_14993);
xor U15759 (N_15759,N_14117,N_14490);
xnor U15760 (N_15760,N_14969,N_13133);
xnor U15761 (N_15761,N_12742,N_12874);
nand U15762 (N_15762,N_14402,N_13533);
xor U15763 (N_15763,N_14403,N_13669);
or U15764 (N_15764,N_12577,N_13250);
and U15765 (N_15765,N_13475,N_14038);
and U15766 (N_15766,N_14797,N_14929);
nand U15767 (N_15767,N_14715,N_14581);
and U15768 (N_15768,N_14994,N_14166);
and U15769 (N_15769,N_12557,N_14532);
and U15770 (N_15770,N_14204,N_13854);
and U15771 (N_15771,N_13967,N_13490);
nor U15772 (N_15772,N_14816,N_14703);
xor U15773 (N_15773,N_14587,N_14946);
nor U15774 (N_15774,N_13539,N_14042);
nor U15775 (N_15775,N_14267,N_13449);
nor U15776 (N_15776,N_13264,N_14010);
and U15777 (N_15777,N_12728,N_14136);
and U15778 (N_15778,N_12765,N_14714);
nor U15779 (N_15779,N_13319,N_13721);
nor U15780 (N_15780,N_13458,N_13790);
nor U15781 (N_15781,N_13415,N_12696);
nor U15782 (N_15782,N_12550,N_13023);
nand U15783 (N_15783,N_12947,N_14956);
and U15784 (N_15784,N_13148,N_14795);
or U15785 (N_15785,N_13766,N_13127);
nand U15786 (N_15786,N_13599,N_14013);
and U15787 (N_15787,N_14035,N_13340);
or U15788 (N_15788,N_13136,N_12717);
xnor U15789 (N_15789,N_14784,N_12855);
nand U15790 (N_15790,N_13723,N_14926);
xor U15791 (N_15791,N_12771,N_12928);
nor U15792 (N_15792,N_13019,N_14899);
xnor U15793 (N_15793,N_14989,N_12561);
nor U15794 (N_15794,N_13706,N_13844);
nand U15795 (N_15795,N_13547,N_14473);
or U15796 (N_15796,N_13154,N_12894);
nor U15797 (N_15797,N_13244,N_13900);
and U15798 (N_15798,N_13467,N_13557);
or U15799 (N_15799,N_12763,N_14367);
or U15800 (N_15800,N_14158,N_14558);
nor U15801 (N_15801,N_14905,N_13495);
nor U15802 (N_15802,N_13491,N_14140);
or U15803 (N_15803,N_14579,N_14869);
nand U15804 (N_15804,N_12716,N_14116);
or U15805 (N_15805,N_14553,N_13972);
nor U15806 (N_15806,N_12954,N_14303);
nand U15807 (N_15807,N_13182,N_14109);
xnor U15808 (N_15808,N_14470,N_13263);
nand U15809 (N_15809,N_14562,N_14736);
nor U15810 (N_15810,N_14803,N_14469);
and U15811 (N_15811,N_14081,N_14790);
nand U15812 (N_15812,N_14188,N_12700);
and U15813 (N_15813,N_13369,N_13069);
or U15814 (N_15814,N_14739,N_14070);
nor U15815 (N_15815,N_13350,N_12950);
nor U15816 (N_15816,N_14904,N_14280);
or U15817 (N_15817,N_14611,N_14115);
nor U15818 (N_15818,N_13344,N_14408);
xnor U15819 (N_15819,N_14815,N_14272);
nand U15820 (N_15820,N_12919,N_12657);
and U15821 (N_15821,N_13138,N_13455);
and U15822 (N_15822,N_13836,N_13750);
or U15823 (N_15823,N_14409,N_14000);
nor U15824 (N_15824,N_13343,N_13585);
or U15825 (N_15825,N_12694,N_12552);
and U15826 (N_15826,N_13819,N_13927);
nand U15827 (N_15827,N_13714,N_14487);
xnor U15828 (N_15828,N_14805,N_13186);
or U15829 (N_15829,N_12591,N_13952);
xnor U15830 (N_15830,N_13346,N_13441);
xor U15831 (N_15831,N_13977,N_14690);
or U15832 (N_15832,N_13109,N_13142);
nor U15833 (N_15833,N_14326,N_14977);
xnor U15834 (N_15834,N_12559,N_14966);
nand U15835 (N_15835,N_14356,N_13349);
and U15836 (N_15836,N_14131,N_13473);
nor U15837 (N_15837,N_13641,N_13380);
nand U15838 (N_15838,N_13761,N_12612);
or U15839 (N_15839,N_13583,N_14859);
xnor U15840 (N_15840,N_13279,N_12789);
nand U15841 (N_15841,N_14071,N_14971);
and U15842 (N_15842,N_14662,N_12881);
or U15843 (N_15843,N_14096,N_14274);
nor U15844 (N_15844,N_13628,N_13582);
and U15845 (N_15845,N_12606,N_13858);
or U15846 (N_15846,N_14891,N_14236);
nor U15847 (N_15847,N_13008,N_13999);
xor U15848 (N_15848,N_12748,N_14088);
or U15849 (N_15849,N_14299,N_13847);
or U15850 (N_15850,N_13471,N_13437);
and U15851 (N_15851,N_13891,N_13532);
nand U15852 (N_15852,N_13303,N_13435);
xnor U15853 (N_15853,N_13051,N_13817);
xnor U15854 (N_15854,N_14192,N_12951);
nand U15855 (N_15855,N_13901,N_13280);
or U15856 (N_15856,N_14973,N_14991);
or U15857 (N_15857,N_14164,N_14890);
and U15858 (N_15858,N_13212,N_12858);
xnor U15859 (N_15859,N_13119,N_14467);
nand U15860 (N_15860,N_12676,N_14346);
nor U15861 (N_15861,N_14072,N_13741);
and U15862 (N_15862,N_12933,N_14215);
nand U15863 (N_15863,N_14074,N_12563);
or U15864 (N_15864,N_14445,N_13941);
and U15865 (N_15865,N_13196,N_14491);
nor U15866 (N_15866,N_13864,N_14724);
nand U15867 (N_15867,N_14547,N_13526);
and U15868 (N_15868,N_13784,N_14032);
or U15869 (N_15869,N_14920,N_12829);
xor U15870 (N_15870,N_14251,N_14150);
xor U15871 (N_15871,N_12523,N_12831);
xnor U15872 (N_15872,N_12712,N_14069);
xnor U15873 (N_15873,N_13828,N_13593);
xnor U15874 (N_15874,N_13200,N_14673);
and U15875 (N_15875,N_12759,N_14600);
xor U15876 (N_15876,N_13395,N_13181);
nor U15877 (N_15877,N_14341,N_14846);
or U15878 (N_15878,N_14417,N_14480);
nand U15879 (N_15879,N_12596,N_12673);
nor U15880 (N_15880,N_13853,N_13117);
or U15881 (N_15881,N_13746,N_12608);
nor U15882 (N_15882,N_12624,N_12997);
or U15883 (N_15883,N_13202,N_14511);
and U15884 (N_15884,N_14646,N_14279);
nor U15885 (N_15885,N_14051,N_12968);
or U15886 (N_15886,N_13383,N_14181);
or U15887 (N_15887,N_14436,N_14086);
or U15888 (N_15888,N_14338,N_14641);
and U15889 (N_15889,N_13535,N_14594);
or U15890 (N_15890,N_12579,N_14212);
nor U15891 (N_15891,N_13100,N_12741);
nor U15892 (N_15892,N_13881,N_13129);
nor U15893 (N_15893,N_14935,N_13055);
or U15894 (N_15894,N_13521,N_13321);
nor U15895 (N_15895,N_13871,N_13876);
and U15896 (N_15896,N_13618,N_13976);
or U15897 (N_15897,N_14758,N_14987);
and U15898 (N_15898,N_14458,N_13338);
nor U15899 (N_15899,N_13694,N_12697);
xnor U15900 (N_15900,N_12988,N_13017);
nand U15901 (N_15901,N_14343,N_13145);
or U15902 (N_15902,N_14129,N_14485);
or U15903 (N_15903,N_13588,N_14786);
xnor U15904 (N_15904,N_12960,N_12827);
or U15905 (N_15905,N_14764,N_12598);
xnor U15906 (N_15906,N_14334,N_14373);
and U15907 (N_15907,N_13001,N_12821);
nor U15908 (N_15908,N_14519,N_12786);
or U15909 (N_15909,N_14630,N_13862);
nand U15910 (N_15910,N_13787,N_13841);
nand U15911 (N_15911,N_12524,N_13082);
and U15912 (N_15912,N_14743,N_14538);
or U15913 (N_15913,N_14384,N_12752);
xnor U15914 (N_15914,N_13542,N_13032);
nand U15915 (N_15915,N_13755,N_13198);
nor U15916 (N_15916,N_13627,N_12898);
xor U15917 (N_15917,N_13753,N_12636);
nand U15918 (N_15918,N_14586,N_14811);
nand U15919 (N_15919,N_13497,N_14621);
or U15920 (N_15920,N_14631,N_14098);
and U15921 (N_15921,N_13544,N_13782);
nand U15922 (N_15922,N_13239,N_14550);
xnor U15923 (N_15923,N_13734,N_13131);
xor U15924 (N_15924,N_14352,N_13868);
nand U15925 (N_15925,N_14955,N_14734);
nor U15926 (N_15926,N_14754,N_13937);
nor U15927 (N_15927,N_13478,N_13631);
xnor U15928 (N_15928,N_12534,N_13111);
and U15929 (N_15929,N_13752,N_14750);
and U15930 (N_15930,N_13261,N_14359);
nand U15931 (N_15931,N_12730,N_13469);
nand U15932 (N_15932,N_14130,N_13376);
and U15933 (N_15933,N_13081,N_12974);
and U15934 (N_15934,N_13554,N_12907);
xor U15935 (N_15935,N_13940,N_14546);
or U15936 (N_15936,N_12792,N_12670);
nand U15937 (N_15937,N_12704,N_14556);
nor U15938 (N_15938,N_14934,N_14156);
or U15939 (N_15939,N_14821,N_13462);
nand U15940 (N_15940,N_14386,N_14897);
or U15941 (N_15941,N_14701,N_13655);
nor U15942 (N_15942,N_14471,N_14737);
nand U15943 (N_15943,N_12756,N_14894);
or U15944 (N_15944,N_12626,N_12595);
or U15945 (N_15945,N_13044,N_14198);
and U15946 (N_15946,N_14438,N_14159);
xor U15947 (N_15947,N_14455,N_13823);
or U15948 (N_15948,N_13246,N_14574);
nand U15949 (N_15949,N_12709,N_14001);
nor U15950 (N_15950,N_14913,N_13834);
or U15951 (N_15951,N_12631,N_12527);
xnor U15952 (N_15952,N_13939,N_14608);
and U15953 (N_15953,N_14995,N_13372);
nor U15954 (N_15954,N_12905,N_12734);
or U15955 (N_15955,N_12977,N_14449);
nand U15956 (N_15956,N_14431,N_14849);
nand U15957 (N_15957,N_13072,N_14515);
xor U15958 (N_15958,N_13592,N_13915);
nand U15959 (N_15959,N_14132,N_12810);
or U15960 (N_15960,N_12623,N_14833);
nand U15961 (N_15961,N_12819,N_14462);
nor U15962 (N_15962,N_13658,N_13433);
nor U15963 (N_15963,N_13604,N_14073);
nand U15964 (N_15964,N_13906,N_13336);
and U15965 (N_15965,N_12754,N_12723);
and U15966 (N_15966,N_13037,N_13034);
and U15967 (N_15967,N_13207,N_14266);
xnor U15968 (N_15968,N_13096,N_12653);
xnor U15969 (N_15969,N_13683,N_12995);
or U15970 (N_15970,N_14277,N_14823);
or U15971 (N_15971,N_13843,N_13351);
nand U15972 (N_15972,N_14741,N_13553);
nor U15973 (N_15973,N_13068,N_14033);
or U15974 (N_15974,N_14201,N_14230);
nor U15975 (N_15975,N_12604,N_14903);
and U15976 (N_15976,N_14844,N_14020);
nand U15977 (N_15977,N_14054,N_12978);
nor U15978 (N_15978,N_13932,N_12817);
nor U15979 (N_15979,N_14729,N_12611);
xnor U15980 (N_15980,N_14339,N_13124);
nand U15981 (N_15981,N_14452,N_12863);
or U15982 (N_15982,N_14448,N_14796);
or U15983 (N_15983,N_12533,N_13894);
and U15984 (N_15984,N_13595,N_13240);
nand U15985 (N_15985,N_14707,N_13668);
or U15986 (N_15986,N_13334,N_14189);
and U15987 (N_15987,N_12828,N_14873);
nand U15988 (N_15988,N_14186,N_13835);
xor U15989 (N_15989,N_14980,N_12836);
nand U15990 (N_15990,N_13370,N_12945);
xor U15991 (N_15991,N_14496,N_13691);
nor U15992 (N_15992,N_13128,N_13291);
nand U15993 (N_15993,N_13716,N_13703);
or U15994 (N_15994,N_14979,N_13021);
xor U15995 (N_15995,N_12851,N_14999);
xor U15996 (N_15996,N_14252,N_13531);
xnor U15997 (N_15997,N_13579,N_14433);
nor U15998 (N_15998,N_14244,N_12885);
nor U15999 (N_15999,N_12801,N_13551);
nand U16000 (N_16000,N_13647,N_14420);
nand U16001 (N_16001,N_14055,N_13012);
xor U16002 (N_16002,N_13116,N_12948);
nand U16003 (N_16003,N_12936,N_14354);
nand U16004 (N_16004,N_13161,N_12554);
nor U16005 (N_16005,N_12930,N_14090);
and U16006 (N_16006,N_13166,N_13492);
or U16007 (N_16007,N_13648,N_13908);
and U16008 (N_16008,N_12932,N_13311);
and U16009 (N_16009,N_14762,N_14883);
nand U16010 (N_16010,N_14123,N_14242);
and U16011 (N_16011,N_13722,N_13221);
nor U16012 (N_16012,N_14718,N_14721);
and U16013 (N_16013,N_12500,N_13115);
xnor U16014 (N_16014,N_13218,N_14906);
nor U16015 (N_16015,N_13290,N_13446);
nor U16016 (N_16016,N_14698,N_13724);
xnor U16017 (N_16017,N_14857,N_14100);
or U16018 (N_16018,N_14389,N_13536);
and U16019 (N_16019,N_12845,N_13666);
nand U16020 (N_16020,N_14065,N_14682);
and U16021 (N_16021,N_14243,N_13947);
nand U16022 (N_16022,N_13849,N_14079);
nor U16023 (N_16023,N_14371,N_13177);
nor U16024 (N_16024,N_14453,N_13985);
nor U16025 (N_16025,N_14312,N_13751);
nand U16026 (N_16026,N_14886,N_14628);
xnor U16027 (N_16027,N_13409,N_14826);
xnor U16028 (N_16028,N_14885,N_13936);
nor U16029 (N_16029,N_14742,N_14882);
or U16030 (N_16030,N_13663,N_13623);
nand U16031 (N_16031,N_12544,N_13719);
nand U16032 (N_16032,N_13505,N_14495);
nor U16033 (N_16033,N_14049,N_13774);
and U16034 (N_16034,N_14874,N_13077);
and U16035 (N_16035,N_12982,N_14227);
or U16036 (N_16036,N_14578,N_13459);
and U16037 (N_16037,N_14740,N_13046);
or U16038 (N_16038,N_13204,N_14172);
and U16039 (N_16039,N_14404,N_14573);
or U16040 (N_16040,N_13026,N_13268);
and U16041 (N_16041,N_14822,N_12745);
nand U16042 (N_16042,N_13555,N_13777);
xor U16043 (N_16043,N_12597,N_14836);
nor U16044 (N_16044,N_12970,N_14477);
and U16045 (N_16045,N_13682,N_13527);
nand U16046 (N_16046,N_13139,N_13501);
and U16047 (N_16047,N_14706,N_13904);
or U16048 (N_16048,N_14014,N_14228);
nor U16049 (N_16049,N_14931,N_14613);
or U16050 (N_16050,N_14160,N_13373);
and U16051 (N_16051,N_14502,N_14853);
or U16052 (N_16052,N_13574,N_14287);
nor U16053 (N_16053,N_14535,N_13993);
or U16054 (N_16054,N_13866,N_13770);
and U16055 (N_16055,N_13982,N_13425);
and U16056 (N_16056,N_12939,N_14047);
xnor U16057 (N_16057,N_13922,N_14533);
xnor U16058 (N_16058,N_12567,N_14705);
nand U16059 (N_16059,N_14435,N_14541);
nand U16060 (N_16060,N_12952,N_12878);
xor U16061 (N_16061,N_14031,N_14311);
and U16062 (N_16062,N_13635,N_12980);
xor U16063 (N_16063,N_14363,N_13498);
xnor U16064 (N_16064,N_13735,N_12731);
and U16065 (N_16065,N_13310,N_14421);
xnor U16066 (N_16066,N_14292,N_13687);
nor U16067 (N_16067,N_12774,N_12675);
and U16068 (N_16068,N_12706,N_14523);
nand U16069 (N_16069,N_14713,N_14793);
and U16070 (N_16070,N_13195,N_13488);
nor U16071 (N_16071,N_12698,N_14559);
xnor U16072 (N_16072,N_13382,N_14870);
nand U16073 (N_16073,N_14133,N_12912);
or U16074 (N_16074,N_14337,N_12576);
or U16075 (N_16075,N_14571,N_12743);
nand U16076 (N_16076,N_14099,N_14930);
nor U16077 (N_16077,N_14582,N_14660);
and U16078 (N_16078,N_14472,N_13622);
and U16079 (N_16079,N_13965,N_14813);
and U16080 (N_16080,N_12886,N_14612);
xor U16081 (N_16081,N_13651,N_12837);
or U16082 (N_16082,N_14610,N_14654);
or U16083 (N_16083,N_13036,N_13237);
nor U16084 (N_16084,N_14996,N_13159);
and U16085 (N_16085,N_13895,N_14537);
or U16086 (N_16086,N_13813,N_14513);
or U16087 (N_16087,N_14482,N_14918);
xnor U16088 (N_16088,N_14008,N_12521);
nand U16089 (N_16089,N_13134,N_13919);
nor U16090 (N_16090,N_13759,N_13899);
nor U16091 (N_16091,N_14827,N_14916);
and U16092 (N_16092,N_13730,N_13522);
and U16093 (N_16093,N_13440,N_14687);
and U16094 (N_16094,N_14777,N_14985);
nor U16095 (N_16095,N_13172,N_13892);
xor U16096 (N_16096,N_14282,N_13833);
and U16097 (N_16097,N_13749,N_13616);
or U16098 (N_16098,N_13258,N_14692);
nand U16099 (N_16099,N_13700,N_12691);
and U16100 (N_16100,N_13608,N_13073);
and U16101 (N_16101,N_12705,N_12532);
or U16102 (N_16102,N_14149,N_14723);
nor U16103 (N_16103,N_14105,N_14413);
or U16104 (N_16104,N_14938,N_13084);
nor U16105 (N_16105,N_12910,N_13558);
and U16106 (N_16106,N_13080,N_14468);
and U16107 (N_16107,N_13067,N_12969);
and U16108 (N_16108,N_13188,N_13030);
or U16109 (N_16109,N_12665,N_13029);
xor U16110 (N_16110,N_14026,N_14318);
and U16111 (N_16111,N_13893,N_12909);
xor U16112 (N_16112,N_13479,N_13677);
and U16113 (N_16113,N_14368,N_14804);
nor U16114 (N_16114,N_13537,N_14209);
and U16115 (N_16115,N_13494,N_14506);
and U16116 (N_16116,N_13775,N_13717);
or U16117 (N_16117,N_13394,N_12589);
xnor U16118 (N_16118,N_14028,N_14254);
or U16119 (N_16119,N_14954,N_12513);
nor U16120 (N_16120,N_14976,N_14210);
nand U16121 (N_16121,N_12650,N_12946);
nand U16122 (N_16122,N_12540,N_13518);
xor U16123 (N_16123,N_13185,N_13875);
nand U16124 (N_16124,N_13676,N_13845);
nor U16125 (N_16125,N_13885,N_13120);
or U16126 (N_16126,N_14751,N_14370);
nand U16127 (N_16127,N_12937,N_13432);
xnor U16128 (N_16128,N_14250,N_14233);
nand U16129 (N_16129,N_14840,N_12582);
nor U16130 (N_16130,N_13031,N_13171);
nand U16131 (N_16131,N_13913,N_14818);
and U16132 (N_16132,N_12652,N_14972);
or U16133 (N_16133,N_13772,N_13883);
nor U16134 (N_16134,N_14321,N_13971);
xor U16135 (N_16135,N_13043,N_12802);
and U16136 (N_16136,N_14214,N_12713);
or U16137 (N_16137,N_13152,N_13672);
nand U16138 (N_16138,N_13933,N_13805);
xor U16139 (N_16139,N_12830,N_13324);
or U16140 (N_16140,N_12655,N_12901);
or U16141 (N_16141,N_13793,N_14832);
nor U16142 (N_16142,N_12668,N_12790);
or U16143 (N_16143,N_13146,N_14658);
or U16144 (N_16144,N_13856,N_13199);
xor U16145 (N_16145,N_14393,N_14802);
nand U16146 (N_16146,N_13151,N_14092);
xnor U16147 (N_16147,N_13930,N_12993);
and U16148 (N_16148,N_13226,N_13508);
nand U16149 (N_16149,N_12908,N_13804);
nand U16150 (N_16150,N_12503,N_13778);
nand U16151 (N_16151,N_14278,N_13103);
nand U16152 (N_16152,N_12649,N_13946);
nand U16153 (N_16153,N_13213,N_12766);
nand U16154 (N_16154,N_13071,N_13270);
nor U16155 (N_16155,N_12583,N_14298);
nor U16156 (N_16156,N_13113,N_14965);
nand U16157 (N_16157,N_13827,N_14774);
nor U16158 (N_16158,N_12627,N_13619);
and U16159 (N_16159,N_14782,N_14643);
nand U16160 (N_16160,N_13418,N_13405);
xor U16161 (N_16161,N_13605,N_13764);
nor U16162 (N_16162,N_13024,N_12639);
nor U16163 (N_16163,N_14867,N_13173);
nor U16164 (N_16164,N_12610,N_13050);
nor U16165 (N_16165,N_13732,N_13194);
nand U16166 (N_16166,N_14974,N_14923);
and U16167 (N_16167,N_12913,N_13260);
nand U16168 (N_16168,N_12671,N_13060);
nand U16169 (N_16169,N_13203,N_12720);
or U16170 (N_16170,N_13671,N_13696);
or U16171 (N_16171,N_13223,N_12869);
and U16172 (N_16172,N_13157,N_14245);
nor U16173 (N_16173,N_14336,N_14728);
nand U16174 (N_16174,N_13573,N_14588);
xor U16175 (N_16175,N_13013,N_14779);
and U16176 (N_16176,N_14061,N_14135);
and U16177 (N_16177,N_13088,N_14868);
nor U16178 (N_16178,N_14221,N_14585);
and U16179 (N_16179,N_14216,N_13621);
nor U16180 (N_16180,N_13884,N_14157);
nor U16181 (N_16181,N_13859,N_13822);
and U16182 (N_16182,N_14476,N_12560);
xnor U16183 (N_16183,N_14143,N_12873);
nand U16184 (N_16184,N_13530,N_14637);
or U16185 (N_16185,N_12659,N_13086);
and U16186 (N_16186,N_14789,N_14375);
xnor U16187 (N_16187,N_13481,N_12918);
nand U16188 (N_16188,N_14232,N_14647);
nor U16189 (N_16189,N_13970,N_13889);
nand U16190 (N_16190,N_12849,N_12987);
and U16191 (N_16191,N_14323,N_14479);
nand U16192 (N_16192,N_13842,N_13920);
nand U16193 (N_16193,N_13407,N_14290);
and U16194 (N_16194,N_13958,N_12739);
or U16195 (N_16195,N_13316,N_14036);
xnor U16196 (N_16196,N_13454,N_12758);
and U16197 (N_16197,N_12832,N_13265);
nand U16198 (N_16198,N_12833,N_13153);
nand U16199 (N_16199,N_14275,N_13880);
or U16200 (N_16200,N_13613,N_13474);
nand U16201 (N_16201,N_14921,N_13484);
xor U16202 (N_16202,N_12753,N_14120);
nor U16203 (N_16203,N_14842,N_13132);
and U16204 (N_16204,N_13301,N_13236);
or U16205 (N_16205,N_13499,N_13646);
xor U16206 (N_16206,N_14500,N_14520);
or U16207 (N_16207,N_13543,N_12876);
and U16208 (N_16208,N_14241,N_13546);
xor U16209 (N_16209,N_13726,N_13785);
xor U16210 (N_16210,N_14068,N_13385);
nor U16211 (N_16211,N_12535,N_13910);
nand U16212 (N_16212,N_14284,N_14642);
nand U16213 (N_16213,N_13638,N_14866);
xor U16214 (N_16214,N_13353,N_13176);
and U16215 (N_16215,N_14211,N_13294);
xnor U16216 (N_16216,N_13587,N_13800);
nor U16217 (N_16217,N_13253,N_14325);
or U16218 (N_16218,N_13990,N_14678);
and U16219 (N_16219,N_12957,N_13607);
and U16220 (N_16220,N_13267,N_12699);
nand U16221 (N_16221,N_12531,N_13964);
nand U16222 (N_16222,N_13960,N_14661);
and U16223 (N_16223,N_13091,N_12994);
nand U16224 (N_16224,N_14843,N_14604);
xnor U16225 (N_16225,N_13792,N_13525);
nor U16226 (N_16226,N_14398,N_14584);
and U16227 (N_16227,N_12796,N_13538);
nor U16228 (N_16228,N_13811,N_14620);
nor U16229 (N_16229,N_13564,N_12747);
nor U16230 (N_16230,N_13371,N_13873);
xor U16231 (N_16231,N_14494,N_12895);
xor U16232 (N_16232,N_12585,N_12813);
or U16233 (N_16233,N_14810,N_12590);
xnor U16234 (N_16234,N_14878,N_13661);
nor U16235 (N_16235,N_13837,N_14944);
nor U16236 (N_16236,N_14056,N_14432);
or U16237 (N_16237,N_12509,N_14970);
xor U16238 (N_16238,N_14457,N_12508);
or U16239 (N_16239,N_13821,N_14710);
xnor U16240 (N_16240,N_14850,N_14234);
nand U16241 (N_16241,N_14828,N_14665);
or U16242 (N_16242,N_12683,N_13178);
xnor U16243 (N_16243,N_14772,N_12519);
or U16244 (N_16244,N_12515,N_14992);
nor U16245 (N_16245,N_14145,N_13255);
and U16246 (N_16246,N_13609,N_13707);
or U16247 (N_16247,N_12890,N_12685);
nand U16248 (N_16248,N_13517,N_14270);
and U16249 (N_16249,N_14884,N_14914);
or U16250 (N_16250,N_13920,N_13023);
or U16251 (N_16251,N_13160,N_13652);
and U16252 (N_16252,N_14726,N_14634);
and U16253 (N_16253,N_12848,N_12798);
or U16254 (N_16254,N_14629,N_14712);
and U16255 (N_16255,N_12717,N_12883);
xnor U16256 (N_16256,N_14862,N_13051);
and U16257 (N_16257,N_13256,N_14018);
nand U16258 (N_16258,N_14206,N_13376);
nand U16259 (N_16259,N_12582,N_12872);
and U16260 (N_16260,N_14761,N_12933);
xnor U16261 (N_16261,N_12747,N_14316);
xnor U16262 (N_16262,N_12658,N_13887);
and U16263 (N_16263,N_13954,N_13968);
or U16264 (N_16264,N_12867,N_13220);
and U16265 (N_16265,N_13760,N_14746);
or U16266 (N_16266,N_12513,N_13717);
and U16267 (N_16267,N_12553,N_12732);
nor U16268 (N_16268,N_13243,N_14239);
or U16269 (N_16269,N_14936,N_13959);
nand U16270 (N_16270,N_14468,N_13573);
xor U16271 (N_16271,N_14860,N_13456);
xor U16272 (N_16272,N_14584,N_14230);
and U16273 (N_16273,N_13335,N_13489);
nand U16274 (N_16274,N_13166,N_13653);
and U16275 (N_16275,N_13676,N_13147);
or U16276 (N_16276,N_14200,N_12988);
nor U16277 (N_16277,N_13263,N_14690);
or U16278 (N_16278,N_12531,N_12757);
nor U16279 (N_16279,N_14338,N_12738);
and U16280 (N_16280,N_14685,N_12803);
and U16281 (N_16281,N_13149,N_14040);
nand U16282 (N_16282,N_14913,N_14218);
nand U16283 (N_16283,N_13939,N_13501);
xnor U16284 (N_16284,N_13417,N_14235);
or U16285 (N_16285,N_14558,N_13370);
and U16286 (N_16286,N_13601,N_14390);
or U16287 (N_16287,N_12533,N_13170);
nand U16288 (N_16288,N_14101,N_12716);
and U16289 (N_16289,N_13808,N_14524);
and U16290 (N_16290,N_12512,N_12604);
nor U16291 (N_16291,N_14971,N_13488);
or U16292 (N_16292,N_12915,N_13781);
nand U16293 (N_16293,N_14081,N_14194);
or U16294 (N_16294,N_12657,N_14565);
or U16295 (N_16295,N_14133,N_12501);
and U16296 (N_16296,N_14379,N_13251);
and U16297 (N_16297,N_14227,N_14053);
xor U16298 (N_16298,N_13490,N_14670);
nand U16299 (N_16299,N_12617,N_13324);
nand U16300 (N_16300,N_13890,N_14112);
and U16301 (N_16301,N_12725,N_14960);
nand U16302 (N_16302,N_12758,N_13164);
nand U16303 (N_16303,N_14906,N_14827);
nand U16304 (N_16304,N_12811,N_13046);
and U16305 (N_16305,N_14250,N_14830);
or U16306 (N_16306,N_13675,N_12946);
nor U16307 (N_16307,N_14271,N_13559);
or U16308 (N_16308,N_13802,N_14807);
or U16309 (N_16309,N_13480,N_14389);
nor U16310 (N_16310,N_13579,N_14351);
nor U16311 (N_16311,N_14335,N_13159);
and U16312 (N_16312,N_14627,N_14690);
or U16313 (N_16313,N_13995,N_12568);
nor U16314 (N_16314,N_13960,N_14791);
and U16315 (N_16315,N_13362,N_12985);
nor U16316 (N_16316,N_14972,N_13603);
and U16317 (N_16317,N_14927,N_12987);
or U16318 (N_16318,N_12525,N_13544);
nor U16319 (N_16319,N_13690,N_13485);
xor U16320 (N_16320,N_13204,N_12522);
nor U16321 (N_16321,N_13070,N_12982);
and U16322 (N_16322,N_14302,N_12808);
and U16323 (N_16323,N_12777,N_14686);
nor U16324 (N_16324,N_14507,N_14591);
nand U16325 (N_16325,N_14091,N_13583);
and U16326 (N_16326,N_12632,N_14563);
nand U16327 (N_16327,N_13125,N_14682);
nand U16328 (N_16328,N_13524,N_14048);
nand U16329 (N_16329,N_13010,N_12987);
and U16330 (N_16330,N_12974,N_14799);
xor U16331 (N_16331,N_14504,N_14554);
xor U16332 (N_16332,N_12744,N_13050);
xnor U16333 (N_16333,N_13784,N_14729);
nor U16334 (N_16334,N_13811,N_12942);
and U16335 (N_16335,N_12517,N_13733);
and U16336 (N_16336,N_13546,N_14348);
xnor U16337 (N_16337,N_13587,N_13919);
and U16338 (N_16338,N_13562,N_14196);
or U16339 (N_16339,N_14736,N_14236);
and U16340 (N_16340,N_14313,N_14687);
nor U16341 (N_16341,N_14165,N_13736);
and U16342 (N_16342,N_12612,N_13333);
nor U16343 (N_16343,N_14917,N_14850);
or U16344 (N_16344,N_12667,N_13172);
xor U16345 (N_16345,N_14658,N_14389);
xor U16346 (N_16346,N_13523,N_14833);
or U16347 (N_16347,N_13818,N_13006);
xor U16348 (N_16348,N_14539,N_14752);
nor U16349 (N_16349,N_14127,N_14225);
and U16350 (N_16350,N_12663,N_13703);
nand U16351 (N_16351,N_13085,N_12955);
and U16352 (N_16352,N_14755,N_14319);
nor U16353 (N_16353,N_13862,N_14285);
nor U16354 (N_16354,N_13629,N_14357);
xor U16355 (N_16355,N_14059,N_13769);
nand U16356 (N_16356,N_13977,N_12786);
or U16357 (N_16357,N_12679,N_13756);
or U16358 (N_16358,N_12744,N_13502);
and U16359 (N_16359,N_14091,N_14580);
or U16360 (N_16360,N_13546,N_12555);
nand U16361 (N_16361,N_13695,N_14336);
xnor U16362 (N_16362,N_14723,N_12744);
and U16363 (N_16363,N_14135,N_13212);
and U16364 (N_16364,N_14556,N_13505);
and U16365 (N_16365,N_13265,N_13046);
and U16366 (N_16366,N_13440,N_14252);
nand U16367 (N_16367,N_12537,N_14745);
nand U16368 (N_16368,N_13598,N_13261);
nor U16369 (N_16369,N_13355,N_13655);
xnor U16370 (N_16370,N_14111,N_14983);
nand U16371 (N_16371,N_14734,N_13199);
nor U16372 (N_16372,N_13776,N_12552);
or U16373 (N_16373,N_13601,N_13616);
and U16374 (N_16374,N_14082,N_14765);
or U16375 (N_16375,N_13941,N_13613);
or U16376 (N_16376,N_13388,N_14991);
xnor U16377 (N_16377,N_14747,N_14930);
xor U16378 (N_16378,N_14541,N_14692);
xnor U16379 (N_16379,N_12590,N_13208);
or U16380 (N_16380,N_13050,N_13515);
nand U16381 (N_16381,N_13908,N_12606);
and U16382 (N_16382,N_13897,N_13494);
nor U16383 (N_16383,N_14384,N_14727);
or U16384 (N_16384,N_13078,N_13783);
nand U16385 (N_16385,N_13680,N_13797);
nor U16386 (N_16386,N_14123,N_13511);
nand U16387 (N_16387,N_14809,N_14866);
and U16388 (N_16388,N_14143,N_13809);
and U16389 (N_16389,N_13200,N_13551);
nand U16390 (N_16390,N_14794,N_12779);
nand U16391 (N_16391,N_14807,N_13501);
or U16392 (N_16392,N_14221,N_13619);
nor U16393 (N_16393,N_14080,N_14818);
nor U16394 (N_16394,N_13923,N_13461);
nor U16395 (N_16395,N_13544,N_13629);
and U16396 (N_16396,N_14024,N_13159);
nand U16397 (N_16397,N_12629,N_13247);
xnor U16398 (N_16398,N_12829,N_13361);
or U16399 (N_16399,N_13366,N_14229);
nor U16400 (N_16400,N_14673,N_13895);
nor U16401 (N_16401,N_12604,N_14974);
and U16402 (N_16402,N_13404,N_14739);
or U16403 (N_16403,N_14112,N_12701);
nand U16404 (N_16404,N_14030,N_12548);
nand U16405 (N_16405,N_14310,N_14462);
or U16406 (N_16406,N_14901,N_14208);
or U16407 (N_16407,N_14983,N_12953);
xnor U16408 (N_16408,N_14918,N_14152);
xor U16409 (N_16409,N_13813,N_12762);
and U16410 (N_16410,N_13480,N_12838);
and U16411 (N_16411,N_12641,N_14541);
xor U16412 (N_16412,N_13290,N_13091);
xnor U16413 (N_16413,N_14566,N_14021);
nor U16414 (N_16414,N_13817,N_14325);
xnor U16415 (N_16415,N_12818,N_14353);
nor U16416 (N_16416,N_12891,N_13463);
nand U16417 (N_16417,N_13163,N_12571);
and U16418 (N_16418,N_12556,N_13913);
xnor U16419 (N_16419,N_12712,N_14614);
nand U16420 (N_16420,N_14093,N_14673);
nand U16421 (N_16421,N_12572,N_14042);
and U16422 (N_16422,N_13474,N_13639);
xnor U16423 (N_16423,N_13148,N_12766);
or U16424 (N_16424,N_13541,N_13704);
xor U16425 (N_16425,N_14348,N_14629);
nor U16426 (N_16426,N_14669,N_13109);
or U16427 (N_16427,N_14816,N_12516);
or U16428 (N_16428,N_14885,N_13410);
nor U16429 (N_16429,N_14531,N_13354);
xnor U16430 (N_16430,N_14687,N_14438);
or U16431 (N_16431,N_14574,N_14283);
nand U16432 (N_16432,N_13689,N_13764);
nand U16433 (N_16433,N_14560,N_14323);
xnor U16434 (N_16434,N_12913,N_13290);
xor U16435 (N_16435,N_12531,N_13075);
nand U16436 (N_16436,N_14685,N_13883);
xnor U16437 (N_16437,N_14593,N_13642);
and U16438 (N_16438,N_14992,N_12994);
xnor U16439 (N_16439,N_12692,N_14213);
xnor U16440 (N_16440,N_14824,N_14459);
and U16441 (N_16441,N_14522,N_14681);
or U16442 (N_16442,N_12596,N_14777);
xnor U16443 (N_16443,N_14373,N_12893);
nor U16444 (N_16444,N_13955,N_13935);
xor U16445 (N_16445,N_12968,N_12516);
and U16446 (N_16446,N_12746,N_14932);
nor U16447 (N_16447,N_14408,N_14235);
and U16448 (N_16448,N_14981,N_13211);
or U16449 (N_16449,N_13566,N_14336);
nor U16450 (N_16450,N_12573,N_13443);
xnor U16451 (N_16451,N_14485,N_13441);
nor U16452 (N_16452,N_14895,N_14934);
and U16453 (N_16453,N_12860,N_12967);
or U16454 (N_16454,N_13740,N_14187);
xnor U16455 (N_16455,N_13959,N_13948);
nand U16456 (N_16456,N_12993,N_13068);
xnor U16457 (N_16457,N_14793,N_14169);
xor U16458 (N_16458,N_12796,N_12795);
and U16459 (N_16459,N_14703,N_14741);
nand U16460 (N_16460,N_13067,N_13824);
and U16461 (N_16461,N_13752,N_13189);
and U16462 (N_16462,N_13999,N_13268);
nand U16463 (N_16463,N_12611,N_14235);
or U16464 (N_16464,N_14053,N_13658);
or U16465 (N_16465,N_12544,N_14876);
and U16466 (N_16466,N_14048,N_12605);
nand U16467 (N_16467,N_14569,N_12600);
and U16468 (N_16468,N_12631,N_14886);
and U16469 (N_16469,N_13793,N_14424);
or U16470 (N_16470,N_12790,N_14353);
or U16471 (N_16471,N_14325,N_12547);
nand U16472 (N_16472,N_14122,N_14758);
nor U16473 (N_16473,N_12825,N_12725);
nand U16474 (N_16474,N_13127,N_12623);
nor U16475 (N_16475,N_14121,N_13538);
xnor U16476 (N_16476,N_12958,N_13752);
nand U16477 (N_16477,N_13470,N_14717);
xnor U16478 (N_16478,N_14552,N_14824);
nand U16479 (N_16479,N_14988,N_12519);
and U16480 (N_16480,N_14231,N_14550);
xor U16481 (N_16481,N_13909,N_14168);
and U16482 (N_16482,N_12861,N_12548);
xor U16483 (N_16483,N_12742,N_14829);
or U16484 (N_16484,N_14869,N_14844);
xnor U16485 (N_16485,N_13583,N_14529);
and U16486 (N_16486,N_14428,N_14328);
and U16487 (N_16487,N_13839,N_14241);
nand U16488 (N_16488,N_14306,N_13671);
nor U16489 (N_16489,N_14297,N_13316);
nor U16490 (N_16490,N_14784,N_14968);
or U16491 (N_16491,N_12813,N_14961);
and U16492 (N_16492,N_14782,N_14179);
and U16493 (N_16493,N_12570,N_12876);
nand U16494 (N_16494,N_14692,N_14611);
nor U16495 (N_16495,N_12612,N_13397);
nor U16496 (N_16496,N_14328,N_13692);
xor U16497 (N_16497,N_14120,N_13880);
or U16498 (N_16498,N_14423,N_14643);
or U16499 (N_16499,N_14202,N_13574);
and U16500 (N_16500,N_13324,N_13470);
and U16501 (N_16501,N_14069,N_13871);
and U16502 (N_16502,N_14070,N_13068);
and U16503 (N_16503,N_13438,N_13228);
nor U16504 (N_16504,N_13096,N_12638);
xor U16505 (N_16505,N_13416,N_14112);
nand U16506 (N_16506,N_12586,N_14341);
nand U16507 (N_16507,N_13082,N_14250);
nor U16508 (N_16508,N_14541,N_14873);
nor U16509 (N_16509,N_13628,N_14770);
nand U16510 (N_16510,N_14030,N_13840);
and U16511 (N_16511,N_12899,N_13998);
nand U16512 (N_16512,N_12535,N_14347);
xor U16513 (N_16513,N_14329,N_14098);
xor U16514 (N_16514,N_13805,N_13153);
or U16515 (N_16515,N_14742,N_12900);
xor U16516 (N_16516,N_13254,N_13757);
or U16517 (N_16517,N_12822,N_14727);
nor U16518 (N_16518,N_12734,N_14175);
nand U16519 (N_16519,N_12679,N_13305);
xor U16520 (N_16520,N_14296,N_13582);
and U16521 (N_16521,N_14593,N_13985);
or U16522 (N_16522,N_14883,N_12622);
nand U16523 (N_16523,N_14822,N_14234);
or U16524 (N_16524,N_14065,N_14639);
xnor U16525 (N_16525,N_12814,N_14477);
or U16526 (N_16526,N_13005,N_14714);
nor U16527 (N_16527,N_14264,N_14806);
nand U16528 (N_16528,N_14602,N_14269);
or U16529 (N_16529,N_13685,N_12961);
and U16530 (N_16530,N_13987,N_12982);
nor U16531 (N_16531,N_14942,N_14644);
xor U16532 (N_16532,N_13681,N_13860);
nor U16533 (N_16533,N_12570,N_14106);
nand U16534 (N_16534,N_14776,N_14069);
nand U16535 (N_16535,N_14071,N_14188);
nand U16536 (N_16536,N_14929,N_12611);
or U16537 (N_16537,N_12816,N_12559);
nand U16538 (N_16538,N_13201,N_14272);
xnor U16539 (N_16539,N_12992,N_12644);
nor U16540 (N_16540,N_13407,N_12680);
nand U16541 (N_16541,N_14344,N_13187);
xnor U16542 (N_16542,N_13449,N_12640);
or U16543 (N_16543,N_13005,N_12893);
or U16544 (N_16544,N_14472,N_14303);
nor U16545 (N_16545,N_14403,N_13364);
nand U16546 (N_16546,N_13422,N_13311);
xnor U16547 (N_16547,N_13221,N_13651);
and U16548 (N_16548,N_13081,N_14382);
and U16549 (N_16549,N_14188,N_13575);
or U16550 (N_16550,N_14254,N_13297);
and U16551 (N_16551,N_14034,N_14450);
xnor U16552 (N_16552,N_13222,N_13646);
or U16553 (N_16553,N_14741,N_13525);
and U16554 (N_16554,N_14448,N_13495);
xor U16555 (N_16555,N_14211,N_14666);
nor U16556 (N_16556,N_13530,N_13521);
nand U16557 (N_16557,N_12827,N_12707);
or U16558 (N_16558,N_13704,N_14265);
and U16559 (N_16559,N_14634,N_14308);
nand U16560 (N_16560,N_14552,N_14177);
or U16561 (N_16561,N_12956,N_13845);
nand U16562 (N_16562,N_13518,N_13250);
or U16563 (N_16563,N_13363,N_12727);
nand U16564 (N_16564,N_12956,N_13332);
nor U16565 (N_16565,N_13542,N_14213);
nor U16566 (N_16566,N_12969,N_14531);
and U16567 (N_16567,N_14743,N_13891);
nor U16568 (N_16568,N_14357,N_12986);
nor U16569 (N_16569,N_14635,N_14314);
or U16570 (N_16570,N_13425,N_14102);
nand U16571 (N_16571,N_13699,N_14484);
xor U16572 (N_16572,N_12746,N_13686);
xnor U16573 (N_16573,N_12868,N_13047);
nand U16574 (N_16574,N_14615,N_14555);
or U16575 (N_16575,N_12652,N_13384);
nand U16576 (N_16576,N_13447,N_13006);
and U16577 (N_16577,N_12997,N_14626);
nor U16578 (N_16578,N_12945,N_13039);
xor U16579 (N_16579,N_14067,N_14705);
nand U16580 (N_16580,N_13613,N_13670);
xnor U16581 (N_16581,N_14504,N_12706);
xor U16582 (N_16582,N_14110,N_13863);
nand U16583 (N_16583,N_13437,N_13519);
xor U16584 (N_16584,N_12906,N_14573);
xnor U16585 (N_16585,N_14869,N_13965);
nor U16586 (N_16586,N_13187,N_14614);
or U16587 (N_16587,N_13944,N_14377);
nor U16588 (N_16588,N_14800,N_12827);
nor U16589 (N_16589,N_14411,N_14670);
xnor U16590 (N_16590,N_13817,N_14852);
or U16591 (N_16591,N_14840,N_12951);
or U16592 (N_16592,N_14609,N_13588);
xor U16593 (N_16593,N_13733,N_12835);
nor U16594 (N_16594,N_13554,N_12872);
nor U16595 (N_16595,N_14813,N_14489);
nand U16596 (N_16596,N_14313,N_14497);
and U16597 (N_16597,N_14339,N_13815);
and U16598 (N_16598,N_14119,N_13294);
or U16599 (N_16599,N_13016,N_14236);
and U16600 (N_16600,N_14912,N_13500);
nand U16601 (N_16601,N_12736,N_13371);
xor U16602 (N_16602,N_13108,N_14450);
nor U16603 (N_16603,N_13234,N_13677);
or U16604 (N_16604,N_14970,N_13623);
nand U16605 (N_16605,N_13184,N_14580);
or U16606 (N_16606,N_13852,N_13251);
or U16607 (N_16607,N_14028,N_13318);
xnor U16608 (N_16608,N_13084,N_14648);
xnor U16609 (N_16609,N_12525,N_14479);
or U16610 (N_16610,N_14041,N_14459);
xor U16611 (N_16611,N_13281,N_13769);
or U16612 (N_16612,N_12802,N_13277);
or U16613 (N_16613,N_14605,N_13186);
and U16614 (N_16614,N_13488,N_13017);
nand U16615 (N_16615,N_13367,N_13944);
or U16616 (N_16616,N_14764,N_14495);
or U16617 (N_16617,N_12701,N_14162);
and U16618 (N_16618,N_14939,N_12716);
or U16619 (N_16619,N_14039,N_13070);
xnor U16620 (N_16620,N_14421,N_13848);
and U16621 (N_16621,N_14998,N_12595);
or U16622 (N_16622,N_12767,N_14068);
and U16623 (N_16623,N_13314,N_12633);
nand U16624 (N_16624,N_13491,N_13829);
or U16625 (N_16625,N_12814,N_13658);
nor U16626 (N_16626,N_14392,N_12565);
xor U16627 (N_16627,N_13456,N_14531);
xnor U16628 (N_16628,N_13073,N_14730);
and U16629 (N_16629,N_14933,N_13120);
or U16630 (N_16630,N_14906,N_13536);
and U16631 (N_16631,N_14631,N_13004);
xor U16632 (N_16632,N_12733,N_12514);
and U16633 (N_16633,N_12743,N_13545);
or U16634 (N_16634,N_13548,N_12869);
and U16635 (N_16635,N_14640,N_12798);
or U16636 (N_16636,N_13905,N_14183);
and U16637 (N_16637,N_13854,N_14424);
or U16638 (N_16638,N_14970,N_14611);
and U16639 (N_16639,N_14798,N_13988);
nor U16640 (N_16640,N_14601,N_14340);
nor U16641 (N_16641,N_14211,N_12683);
xnor U16642 (N_16642,N_13028,N_14319);
nor U16643 (N_16643,N_12759,N_13478);
nor U16644 (N_16644,N_13409,N_13602);
and U16645 (N_16645,N_14764,N_14909);
nor U16646 (N_16646,N_14287,N_12737);
or U16647 (N_16647,N_14220,N_12885);
and U16648 (N_16648,N_14712,N_14182);
nor U16649 (N_16649,N_12617,N_13352);
xnor U16650 (N_16650,N_13285,N_14414);
nor U16651 (N_16651,N_13025,N_12701);
and U16652 (N_16652,N_13334,N_13971);
nand U16653 (N_16653,N_13822,N_13987);
nand U16654 (N_16654,N_14353,N_13742);
or U16655 (N_16655,N_12734,N_13167);
nand U16656 (N_16656,N_13524,N_13283);
and U16657 (N_16657,N_12921,N_13124);
or U16658 (N_16658,N_12599,N_14051);
or U16659 (N_16659,N_14546,N_14313);
xor U16660 (N_16660,N_14884,N_12545);
nand U16661 (N_16661,N_13438,N_12788);
xor U16662 (N_16662,N_14306,N_14274);
nor U16663 (N_16663,N_14292,N_14970);
nor U16664 (N_16664,N_13080,N_12801);
nor U16665 (N_16665,N_12804,N_14257);
nor U16666 (N_16666,N_13756,N_12569);
or U16667 (N_16667,N_13580,N_13792);
and U16668 (N_16668,N_13230,N_13396);
nor U16669 (N_16669,N_13827,N_14010);
nand U16670 (N_16670,N_13519,N_14472);
xnor U16671 (N_16671,N_14086,N_13569);
nor U16672 (N_16672,N_14516,N_14265);
xnor U16673 (N_16673,N_14281,N_12522);
nor U16674 (N_16674,N_14667,N_13977);
and U16675 (N_16675,N_14319,N_13260);
xnor U16676 (N_16676,N_12844,N_13279);
xor U16677 (N_16677,N_14913,N_13166);
or U16678 (N_16678,N_14175,N_12910);
nand U16679 (N_16679,N_14600,N_12979);
nand U16680 (N_16680,N_13619,N_14749);
xnor U16681 (N_16681,N_14127,N_14765);
xor U16682 (N_16682,N_13370,N_14206);
and U16683 (N_16683,N_12893,N_13454);
nand U16684 (N_16684,N_14928,N_14169);
nor U16685 (N_16685,N_13879,N_13099);
and U16686 (N_16686,N_13564,N_13556);
and U16687 (N_16687,N_13155,N_13195);
and U16688 (N_16688,N_13538,N_13554);
nor U16689 (N_16689,N_13222,N_14950);
or U16690 (N_16690,N_13263,N_12965);
xnor U16691 (N_16691,N_14742,N_13484);
nand U16692 (N_16692,N_12760,N_14589);
nor U16693 (N_16693,N_14609,N_13039);
or U16694 (N_16694,N_12982,N_14095);
nand U16695 (N_16695,N_14263,N_14978);
xor U16696 (N_16696,N_13010,N_13414);
and U16697 (N_16697,N_14828,N_14939);
or U16698 (N_16698,N_14285,N_14543);
and U16699 (N_16699,N_13930,N_13657);
and U16700 (N_16700,N_13200,N_14048);
nor U16701 (N_16701,N_14714,N_14264);
nand U16702 (N_16702,N_14480,N_14295);
xnor U16703 (N_16703,N_14897,N_14889);
and U16704 (N_16704,N_13911,N_12655);
and U16705 (N_16705,N_14697,N_14245);
or U16706 (N_16706,N_13015,N_12753);
xnor U16707 (N_16707,N_12562,N_13920);
or U16708 (N_16708,N_14320,N_14875);
and U16709 (N_16709,N_14137,N_13454);
and U16710 (N_16710,N_13921,N_14259);
nand U16711 (N_16711,N_13994,N_13956);
xnor U16712 (N_16712,N_14272,N_12838);
and U16713 (N_16713,N_13972,N_13163);
or U16714 (N_16714,N_14475,N_14678);
or U16715 (N_16715,N_12625,N_13002);
nor U16716 (N_16716,N_12799,N_14285);
or U16717 (N_16717,N_13098,N_14159);
and U16718 (N_16718,N_14870,N_12716);
and U16719 (N_16719,N_13893,N_13954);
or U16720 (N_16720,N_12652,N_14599);
and U16721 (N_16721,N_14598,N_13054);
nand U16722 (N_16722,N_13793,N_14706);
xor U16723 (N_16723,N_13301,N_13300);
nor U16724 (N_16724,N_13613,N_14604);
or U16725 (N_16725,N_14444,N_12830);
or U16726 (N_16726,N_14186,N_14165);
and U16727 (N_16727,N_14176,N_12829);
and U16728 (N_16728,N_12830,N_14149);
nor U16729 (N_16729,N_13109,N_14699);
nor U16730 (N_16730,N_14564,N_13314);
nand U16731 (N_16731,N_13863,N_14804);
xnor U16732 (N_16732,N_14307,N_13556);
nand U16733 (N_16733,N_14908,N_14010);
xnor U16734 (N_16734,N_12861,N_13890);
nor U16735 (N_16735,N_14780,N_14441);
or U16736 (N_16736,N_13363,N_14499);
nor U16737 (N_16737,N_12678,N_13933);
or U16738 (N_16738,N_14666,N_13050);
nor U16739 (N_16739,N_12874,N_14053);
and U16740 (N_16740,N_14873,N_13613);
nor U16741 (N_16741,N_13013,N_14836);
nor U16742 (N_16742,N_13137,N_13553);
nand U16743 (N_16743,N_12656,N_14657);
nor U16744 (N_16744,N_14639,N_14990);
nor U16745 (N_16745,N_13074,N_13322);
and U16746 (N_16746,N_13085,N_14397);
nor U16747 (N_16747,N_13871,N_14494);
xor U16748 (N_16748,N_14475,N_13556);
and U16749 (N_16749,N_14208,N_12914);
or U16750 (N_16750,N_14850,N_13207);
and U16751 (N_16751,N_12949,N_13385);
or U16752 (N_16752,N_13872,N_13631);
xor U16753 (N_16753,N_13471,N_14508);
xnor U16754 (N_16754,N_12815,N_13618);
or U16755 (N_16755,N_12723,N_14628);
xor U16756 (N_16756,N_13972,N_14600);
nor U16757 (N_16757,N_14778,N_13330);
nor U16758 (N_16758,N_12698,N_14006);
or U16759 (N_16759,N_14935,N_13625);
nand U16760 (N_16760,N_13401,N_14053);
and U16761 (N_16761,N_12977,N_13464);
and U16762 (N_16762,N_14532,N_13888);
nor U16763 (N_16763,N_14016,N_14082);
and U16764 (N_16764,N_14732,N_14329);
or U16765 (N_16765,N_14803,N_14887);
nor U16766 (N_16766,N_13691,N_13474);
nand U16767 (N_16767,N_12650,N_12921);
nor U16768 (N_16768,N_13271,N_14556);
and U16769 (N_16769,N_14449,N_12509);
and U16770 (N_16770,N_12617,N_12609);
xnor U16771 (N_16771,N_13205,N_13359);
and U16772 (N_16772,N_14956,N_12930);
and U16773 (N_16773,N_14773,N_14120);
and U16774 (N_16774,N_14500,N_13328);
nand U16775 (N_16775,N_13913,N_14904);
and U16776 (N_16776,N_12711,N_13683);
and U16777 (N_16777,N_14870,N_14101);
nor U16778 (N_16778,N_14792,N_14483);
nor U16779 (N_16779,N_13598,N_14569);
or U16780 (N_16780,N_14016,N_14424);
nand U16781 (N_16781,N_13752,N_12780);
nor U16782 (N_16782,N_14880,N_13907);
xor U16783 (N_16783,N_13341,N_13622);
or U16784 (N_16784,N_12645,N_13295);
and U16785 (N_16785,N_14559,N_14652);
or U16786 (N_16786,N_14932,N_14690);
nand U16787 (N_16787,N_14529,N_13571);
nor U16788 (N_16788,N_12508,N_14600);
xor U16789 (N_16789,N_13730,N_14944);
or U16790 (N_16790,N_14937,N_12887);
xor U16791 (N_16791,N_13172,N_12962);
or U16792 (N_16792,N_14584,N_12722);
and U16793 (N_16793,N_12815,N_14857);
or U16794 (N_16794,N_14175,N_14719);
and U16795 (N_16795,N_13469,N_14123);
or U16796 (N_16796,N_13517,N_12623);
or U16797 (N_16797,N_12979,N_13815);
or U16798 (N_16798,N_14545,N_13819);
nand U16799 (N_16799,N_13244,N_13860);
nand U16800 (N_16800,N_13222,N_14033);
or U16801 (N_16801,N_13340,N_12858);
nand U16802 (N_16802,N_14276,N_14182);
nand U16803 (N_16803,N_13972,N_14375);
xnor U16804 (N_16804,N_12771,N_14332);
and U16805 (N_16805,N_12954,N_14551);
nor U16806 (N_16806,N_12698,N_13727);
or U16807 (N_16807,N_12994,N_14570);
xor U16808 (N_16808,N_13081,N_13817);
or U16809 (N_16809,N_13175,N_13440);
nor U16810 (N_16810,N_13542,N_12512);
or U16811 (N_16811,N_13199,N_12852);
and U16812 (N_16812,N_12542,N_14025);
and U16813 (N_16813,N_12819,N_12615);
and U16814 (N_16814,N_13203,N_14766);
nand U16815 (N_16815,N_12891,N_12551);
and U16816 (N_16816,N_14432,N_13522);
nor U16817 (N_16817,N_14590,N_13874);
nor U16818 (N_16818,N_12692,N_14402);
and U16819 (N_16819,N_13025,N_14952);
and U16820 (N_16820,N_14141,N_14281);
nand U16821 (N_16821,N_14460,N_13878);
or U16822 (N_16822,N_13842,N_14753);
and U16823 (N_16823,N_13055,N_13426);
nand U16824 (N_16824,N_12668,N_13796);
nor U16825 (N_16825,N_13820,N_14488);
nand U16826 (N_16826,N_12798,N_13104);
nand U16827 (N_16827,N_12864,N_14091);
and U16828 (N_16828,N_13399,N_13407);
nand U16829 (N_16829,N_13496,N_13945);
and U16830 (N_16830,N_14825,N_13696);
xnor U16831 (N_16831,N_14163,N_14863);
nand U16832 (N_16832,N_13805,N_13972);
nor U16833 (N_16833,N_13502,N_13812);
and U16834 (N_16834,N_12976,N_14967);
or U16835 (N_16835,N_13286,N_13633);
nor U16836 (N_16836,N_13336,N_12741);
nand U16837 (N_16837,N_12694,N_13848);
nand U16838 (N_16838,N_12867,N_12667);
xor U16839 (N_16839,N_14890,N_13705);
and U16840 (N_16840,N_14592,N_12809);
and U16841 (N_16841,N_14872,N_13605);
nor U16842 (N_16842,N_14261,N_13128);
xnor U16843 (N_16843,N_14997,N_12726);
xor U16844 (N_16844,N_14615,N_14278);
nand U16845 (N_16845,N_14943,N_14010);
xor U16846 (N_16846,N_14433,N_14409);
and U16847 (N_16847,N_13025,N_14346);
and U16848 (N_16848,N_14297,N_14799);
xnor U16849 (N_16849,N_13116,N_13137);
nand U16850 (N_16850,N_14624,N_13236);
nor U16851 (N_16851,N_14482,N_13263);
and U16852 (N_16852,N_14554,N_12675);
or U16853 (N_16853,N_13534,N_14486);
or U16854 (N_16854,N_13585,N_13149);
xnor U16855 (N_16855,N_12749,N_12949);
nand U16856 (N_16856,N_13854,N_14241);
nor U16857 (N_16857,N_13022,N_14834);
nor U16858 (N_16858,N_14652,N_14218);
and U16859 (N_16859,N_14619,N_14012);
xor U16860 (N_16860,N_12850,N_14932);
or U16861 (N_16861,N_13003,N_13972);
xor U16862 (N_16862,N_14455,N_13149);
or U16863 (N_16863,N_13277,N_14642);
nand U16864 (N_16864,N_13619,N_13362);
nor U16865 (N_16865,N_12554,N_13727);
nand U16866 (N_16866,N_12591,N_13344);
xor U16867 (N_16867,N_12577,N_13562);
nor U16868 (N_16868,N_13138,N_13442);
xnor U16869 (N_16869,N_13922,N_12775);
xor U16870 (N_16870,N_14763,N_13299);
nor U16871 (N_16871,N_13409,N_14753);
and U16872 (N_16872,N_12908,N_13196);
xor U16873 (N_16873,N_13531,N_14572);
and U16874 (N_16874,N_14709,N_14355);
and U16875 (N_16875,N_12562,N_13115);
xor U16876 (N_16876,N_13121,N_14509);
nand U16877 (N_16877,N_12631,N_13706);
or U16878 (N_16878,N_13188,N_13032);
nor U16879 (N_16879,N_12609,N_13474);
nand U16880 (N_16880,N_13248,N_13890);
nor U16881 (N_16881,N_14779,N_13166);
xor U16882 (N_16882,N_12835,N_12816);
xor U16883 (N_16883,N_14933,N_13253);
or U16884 (N_16884,N_13662,N_12897);
xor U16885 (N_16885,N_14168,N_14447);
nor U16886 (N_16886,N_14149,N_14260);
or U16887 (N_16887,N_14469,N_14976);
or U16888 (N_16888,N_13875,N_13611);
nand U16889 (N_16889,N_14316,N_14857);
or U16890 (N_16890,N_13948,N_13563);
and U16891 (N_16891,N_14389,N_12988);
nor U16892 (N_16892,N_14259,N_14468);
nand U16893 (N_16893,N_14022,N_12942);
nor U16894 (N_16894,N_13199,N_14584);
or U16895 (N_16895,N_13512,N_14280);
xnor U16896 (N_16896,N_13090,N_13223);
nor U16897 (N_16897,N_13765,N_12714);
or U16898 (N_16898,N_13921,N_13749);
xnor U16899 (N_16899,N_13718,N_14791);
and U16900 (N_16900,N_14415,N_13687);
or U16901 (N_16901,N_14008,N_12723);
or U16902 (N_16902,N_14837,N_14241);
and U16903 (N_16903,N_14959,N_14482);
or U16904 (N_16904,N_12562,N_13655);
xor U16905 (N_16905,N_12798,N_13498);
and U16906 (N_16906,N_13257,N_13596);
nand U16907 (N_16907,N_13939,N_13532);
and U16908 (N_16908,N_14581,N_12611);
and U16909 (N_16909,N_14591,N_14631);
or U16910 (N_16910,N_14222,N_13357);
or U16911 (N_16911,N_12738,N_13445);
nor U16912 (N_16912,N_13669,N_13119);
nor U16913 (N_16913,N_12704,N_12621);
xnor U16914 (N_16914,N_13700,N_14491);
or U16915 (N_16915,N_13831,N_14258);
or U16916 (N_16916,N_14252,N_13626);
nand U16917 (N_16917,N_14441,N_14369);
nand U16918 (N_16918,N_14248,N_13684);
nand U16919 (N_16919,N_14641,N_12698);
or U16920 (N_16920,N_14834,N_14399);
xnor U16921 (N_16921,N_14869,N_13964);
xnor U16922 (N_16922,N_14651,N_14759);
nand U16923 (N_16923,N_14395,N_13720);
nand U16924 (N_16924,N_14218,N_12707);
or U16925 (N_16925,N_13781,N_12994);
or U16926 (N_16926,N_14628,N_14868);
or U16927 (N_16927,N_13630,N_14381);
nor U16928 (N_16928,N_14495,N_14285);
or U16929 (N_16929,N_12963,N_13596);
and U16930 (N_16930,N_14611,N_14071);
and U16931 (N_16931,N_14704,N_14980);
or U16932 (N_16932,N_13371,N_12979);
and U16933 (N_16933,N_13319,N_12845);
xnor U16934 (N_16934,N_12870,N_13037);
nand U16935 (N_16935,N_14189,N_14102);
and U16936 (N_16936,N_12748,N_13495);
and U16937 (N_16937,N_12685,N_14173);
and U16938 (N_16938,N_14257,N_12977);
nand U16939 (N_16939,N_12625,N_13754);
or U16940 (N_16940,N_13509,N_14176);
or U16941 (N_16941,N_14607,N_14045);
xor U16942 (N_16942,N_13080,N_13744);
and U16943 (N_16943,N_13077,N_14860);
or U16944 (N_16944,N_12877,N_14937);
nor U16945 (N_16945,N_13333,N_14407);
and U16946 (N_16946,N_12605,N_13920);
and U16947 (N_16947,N_13163,N_14428);
and U16948 (N_16948,N_13710,N_12615);
nor U16949 (N_16949,N_14559,N_14535);
nand U16950 (N_16950,N_13963,N_14708);
and U16951 (N_16951,N_12981,N_13973);
or U16952 (N_16952,N_13736,N_13307);
nand U16953 (N_16953,N_12543,N_12542);
nor U16954 (N_16954,N_13517,N_14842);
or U16955 (N_16955,N_14365,N_13139);
nand U16956 (N_16956,N_12857,N_14369);
and U16957 (N_16957,N_13381,N_13473);
and U16958 (N_16958,N_14795,N_13140);
nand U16959 (N_16959,N_13163,N_13670);
nand U16960 (N_16960,N_12617,N_12829);
xnor U16961 (N_16961,N_14631,N_12621);
and U16962 (N_16962,N_14347,N_12908);
or U16963 (N_16963,N_14098,N_12586);
nand U16964 (N_16964,N_13674,N_12828);
nand U16965 (N_16965,N_14134,N_12714);
and U16966 (N_16966,N_14329,N_14315);
nand U16967 (N_16967,N_12623,N_13031);
and U16968 (N_16968,N_14608,N_14243);
nor U16969 (N_16969,N_13173,N_14144);
or U16970 (N_16970,N_14901,N_14480);
nor U16971 (N_16971,N_14515,N_13176);
nand U16972 (N_16972,N_14662,N_14294);
nor U16973 (N_16973,N_13515,N_14029);
nor U16974 (N_16974,N_12538,N_12950);
and U16975 (N_16975,N_13839,N_13430);
nor U16976 (N_16976,N_12740,N_13285);
and U16977 (N_16977,N_13751,N_13798);
nand U16978 (N_16978,N_14000,N_14367);
xnor U16979 (N_16979,N_14026,N_14861);
or U16980 (N_16980,N_13684,N_13853);
nor U16981 (N_16981,N_13739,N_12904);
nor U16982 (N_16982,N_14254,N_14215);
nor U16983 (N_16983,N_13434,N_14410);
and U16984 (N_16984,N_14849,N_14128);
nand U16985 (N_16985,N_14970,N_12876);
nand U16986 (N_16986,N_14435,N_13773);
nor U16987 (N_16987,N_13495,N_13839);
nor U16988 (N_16988,N_14313,N_14770);
xor U16989 (N_16989,N_13224,N_14532);
nand U16990 (N_16990,N_14229,N_13869);
nand U16991 (N_16991,N_14370,N_12691);
nand U16992 (N_16992,N_14016,N_14905);
or U16993 (N_16993,N_12872,N_14825);
xor U16994 (N_16994,N_13116,N_13866);
and U16995 (N_16995,N_14060,N_14001);
xnor U16996 (N_16996,N_13404,N_14784);
xnor U16997 (N_16997,N_13209,N_12578);
nand U16998 (N_16998,N_13730,N_13687);
or U16999 (N_16999,N_14496,N_12993);
xnor U17000 (N_17000,N_13750,N_13716);
and U17001 (N_17001,N_13420,N_14664);
nor U17002 (N_17002,N_14550,N_13374);
and U17003 (N_17003,N_13459,N_12961);
and U17004 (N_17004,N_13555,N_12751);
or U17005 (N_17005,N_13416,N_12910);
or U17006 (N_17006,N_14954,N_14351);
nand U17007 (N_17007,N_13697,N_13731);
and U17008 (N_17008,N_12505,N_14126);
and U17009 (N_17009,N_13151,N_14873);
xor U17010 (N_17010,N_13856,N_14931);
xor U17011 (N_17011,N_14122,N_13168);
and U17012 (N_17012,N_13404,N_13521);
nor U17013 (N_17013,N_14235,N_13319);
and U17014 (N_17014,N_13468,N_13784);
or U17015 (N_17015,N_14508,N_13604);
and U17016 (N_17016,N_14278,N_13260);
xor U17017 (N_17017,N_14214,N_14104);
and U17018 (N_17018,N_13619,N_13038);
nor U17019 (N_17019,N_13083,N_12572);
nor U17020 (N_17020,N_12662,N_12508);
or U17021 (N_17021,N_14258,N_14462);
xor U17022 (N_17022,N_12552,N_13901);
and U17023 (N_17023,N_13578,N_12902);
or U17024 (N_17024,N_14174,N_13279);
nand U17025 (N_17025,N_12786,N_13557);
nand U17026 (N_17026,N_12757,N_12745);
and U17027 (N_17027,N_13607,N_14412);
xnor U17028 (N_17028,N_13381,N_13138);
and U17029 (N_17029,N_14202,N_12691);
or U17030 (N_17030,N_14797,N_14295);
nor U17031 (N_17031,N_14068,N_13925);
and U17032 (N_17032,N_13447,N_12700);
nor U17033 (N_17033,N_14049,N_12897);
or U17034 (N_17034,N_12737,N_14617);
or U17035 (N_17035,N_14974,N_12648);
nor U17036 (N_17036,N_12600,N_12787);
nor U17037 (N_17037,N_13682,N_13832);
and U17038 (N_17038,N_14123,N_13096);
xnor U17039 (N_17039,N_13802,N_13026);
and U17040 (N_17040,N_13153,N_14132);
and U17041 (N_17041,N_13798,N_12693);
xnor U17042 (N_17042,N_13650,N_14153);
nor U17043 (N_17043,N_13069,N_12671);
xor U17044 (N_17044,N_13046,N_12930);
or U17045 (N_17045,N_12706,N_14412);
and U17046 (N_17046,N_12515,N_14248);
xnor U17047 (N_17047,N_12731,N_14858);
nand U17048 (N_17048,N_13672,N_12622);
or U17049 (N_17049,N_13222,N_12940);
nand U17050 (N_17050,N_13403,N_14513);
and U17051 (N_17051,N_12542,N_13029);
and U17052 (N_17052,N_13112,N_12531);
nor U17053 (N_17053,N_14598,N_13056);
or U17054 (N_17054,N_12689,N_14803);
or U17055 (N_17055,N_14250,N_13151);
nand U17056 (N_17056,N_14515,N_14219);
xnor U17057 (N_17057,N_13948,N_14178);
or U17058 (N_17058,N_14063,N_14363);
and U17059 (N_17059,N_14955,N_13580);
or U17060 (N_17060,N_14336,N_14578);
and U17061 (N_17061,N_14590,N_14713);
nor U17062 (N_17062,N_14928,N_13658);
nor U17063 (N_17063,N_12505,N_13283);
and U17064 (N_17064,N_12801,N_14923);
or U17065 (N_17065,N_13405,N_12517);
and U17066 (N_17066,N_14457,N_12876);
or U17067 (N_17067,N_12789,N_13206);
nand U17068 (N_17068,N_12565,N_13282);
xnor U17069 (N_17069,N_13618,N_12670);
nor U17070 (N_17070,N_12740,N_14404);
nor U17071 (N_17071,N_12725,N_13613);
nor U17072 (N_17072,N_12575,N_13427);
nand U17073 (N_17073,N_13976,N_13266);
xnor U17074 (N_17074,N_14885,N_13558);
and U17075 (N_17075,N_13662,N_13430);
and U17076 (N_17076,N_14518,N_13513);
nor U17077 (N_17077,N_14570,N_12963);
xnor U17078 (N_17078,N_14835,N_12958);
nand U17079 (N_17079,N_13328,N_13064);
xnor U17080 (N_17080,N_13610,N_12982);
or U17081 (N_17081,N_14891,N_14324);
nor U17082 (N_17082,N_14107,N_13777);
or U17083 (N_17083,N_13299,N_13381);
nor U17084 (N_17084,N_14636,N_13747);
and U17085 (N_17085,N_12734,N_12880);
or U17086 (N_17086,N_14770,N_14112);
nor U17087 (N_17087,N_14393,N_13908);
nor U17088 (N_17088,N_12709,N_14930);
nand U17089 (N_17089,N_14744,N_12931);
xor U17090 (N_17090,N_13100,N_14404);
nand U17091 (N_17091,N_12634,N_12966);
and U17092 (N_17092,N_12679,N_14376);
nand U17093 (N_17093,N_14120,N_14050);
nand U17094 (N_17094,N_14234,N_14895);
and U17095 (N_17095,N_13402,N_14797);
nand U17096 (N_17096,N_14056,N_13615);
xor U17097 (N_17097,N_13510,N_12573);
nand U17098 (N_17098,N_13399,N_13699);
and U17099 (N_17099,N_12591,N_12626);
nand U17100 (N_17100,N_13649,N_14449);
or U17101 (N_17101,N_12809,N_14650);
xnor U17102 (N_17102,N_14527,N_13557);
or U17103 (N_17103,N_14917,N_12911);
or U17104 (N_17104,N_14427,N_13790);
and U17105 (N_17105,N_14777,N_13352);
and U17106 (N_17106,N_12732,N_14464);
and U17107 (N_17107,N_13548,N_12655);
or U17108 (N_17108,N_12643,N_14045);
nor U17109 (N_17109,N_13342,N_14446);
or U17110 (N_17110,N_13536,N_14586);
nand U17111 (N_17111,N_14628,N_14570);
nor U17112 (N_17112,N_13143,N_13610);
and U17113 (N_17113,N_13718,N_12840);
nand U17114 (N_17114,N_14217,N_14075);
xor U17115 (N_17115,N_14525,N_14060);
or U17116 (N_17116,N_14559,N_14940);
nor U17117 (N_17117,N_14911,N_14337);
nor U17118 (N_17118,N_14899,N_13702);
xor U17119 (N_17119,N_14768,N_13766);
xor U17120 (N_17120,N_12886,N_13547);
and U17121 (N_17121,N_13166,N_14856);
and U17122 (N_17122,N_14691,N_13835);
or U17123 (N_17123,N_12709,N_14239);
and U17124 (N_17124,N_13665,N_14743);
nand U17125 (N_17125,N_14583,N_13925);
nand U17126 (N_17126,N_12876,N_13730);
xnor U17127 (N_17127,N_13103,N_14135);
nand U17128 (N_17128,N_13031,N_12530);
nor U17129 (N_17129,N_12799,N_13874);
nor U17130 (N_17130,N_14867,N_14356);
nor U17131 (N_17131,N_13761,N_14850);
and U17132 (N_17132,N_13904,N_13252);
nand U17133 (N_17133,N_13378,N_13087);
xnor U17134 (N_17134,N_12711,N_13780);
xor U17135 (N_17135,N_13079,N_13876);
or U17136 (N_17136,N_13954,N_14267);
xor U17137 (N_17137,N_13873,N_14235);
or U17138 (N_17138,N_13760,N_14251);
or U17139 (N_17139,N_14943,N_14840);
or U17140 (N_17140,N_14768,N_12865);
and U17141 (N_17141,N_13617,N_13572);
or U17142 (N_17142,N_14355,N_14551);
xnor U17143 (N_17143,N_14810,N_12974);
nor U17144 (N_17144,N_14368,N_14025);
nor U17145 (N_17145,N_14714,N_13713);
and U17146 (N_17146,N_14405,N_13190);
or U17147 (N_17147,N_14907,N_13666);
nor U17148 (N_17148,N_13679,N_13371);
xnor U17149 (N_17149,N_14002,N_14479);
nor U17150 (N_17150,N_14682,N_14481);
and U17151 (N_17151,N_14259,N_14789);
xnor U17152 (N_17152,N_13214,N_13907);
xnor U17153 (N_17153,N_14739,N_12762);
xnor U17154 (N_17154,N_14707,N_13242);
and U17155 (N_17155,N_12594,N_13612);
or U17156 (N_17156,N_12846,N_14113);
nand U17157 (N_17157,N_12957,N_14995);
or U17158 (N_17158,N_12926,N_12519);
or U17159 (N_17159,N_14353,N_13274);
or U17160 (N_17160,N_14548,N_12595);
nand U17161 (N_17161,N_14642,N_13589);
nor U17162 (N_17162,N_13118,N_13631);
nand U17163 (N_17163,N_14992,N_13335);
nand U17164 (N_17164,N_13824,N_13358);
xor U17165 (N_17165,N_13855,N_14457);
nand U17166 (N_17166,N_13927,N_13836);
xor U17167 (N_17167,N_12962,N_13980);
xnor U17168 (N_17168,N_13317,N_12766);
xor U17169 (N_17169,N_13701,N_14691);
nand U17170 (N_17170,N_13888,N_12691);
nand U17171 (N_17171,N_13829,N_14876);
or U17172 (N_17172,N_14134,N_13945);
xnor U17173 (N_17173,N_14802,N_12729);
or U17174 (N_17174,N_13517,N_13846);
nand U17175 (N_17175,N_14388,N_14566);
or U17176 (N_17176,N_13012,N_14938);
nor U17177 (N_17177,N_13811,N_13991);
or U17178 (N_17178,N_14891,N_13639);
or U17179 (N_17179,N_14000,N_12618);
and U17180 (N_17180,N_12621,N_13627);
and U17181 (N_17181,N_13202,N_13260);
nor U17182 (N_17182,N_13242,N_14159);
nand U17183 (N_17183,N_14747,N_14474);
or U17184 (N_17184,N_14003,N_14369);
and U17185 (N_17185,N_13448,N_12696);
nand U17186 (N_17186,N_13041,N_14842);
nor U17187 (N_17187,N_14929,N_13972);
and U17188 (N_17188,N_12886,N_14870);
xor U17189 (N_17189,N_14117,N_14993);
or U17190 (N_17190,N_14797,N_14371);
nand U17191 (N_17191,N_14363,N_13603);
or U17192 (N_17192,N_13093,N_14847);
xnor U17193 (N_17193,N_14773,N_13181);
xor U17194 (N_17194,N_13259,N_14625);
and U17195 (N_17195,N_13156,N_13316);
nand U17196 (N_17196,N_13704,N_14132);
or U17197 (N_17197,N_13004,N_13233);
xnor U17198 (N_17198,N_13703,N_12566);
nor U17199 (N_17199,N_14363,N_14502);
xnor U17200 (N_17200,N_14631,N_12626);
xnor U17201 (N_17201,N_14311,N_13436);
xnor U17202 (N_17202,N_12630,N_12907);
and U17203 (N_17203,N_14873,N_13257);
nor U17204 (N_17204,N_13471,N_12847);
nor U17205 (N_17205,N_13604,N_13709);
and U17206 (N_17206,N_13792,N_14939);
nor U17207 (N_17207,N_12840,N_14430);
xor U17208 (N_17208,N_13535,N_13377);
xnor U17209 (N_17209,N_12909,N_13208);
nor U17210 (N_17210,N_14067,N_13650);
xnor U17211 (N_17211,N_14083,N_13469);
and U17212 (N_17212,N_12535,N_13162);
and U17213 (N_17213,N_13486,N_12730);
xor U17214 (N_17214,N_13649,N_14975);
nand U17215 (N_17215,N_13690,N_14692);
xnor U17216 (N_17216,N_13854,N_13937);
or U17217 (N_17217,N_13583,N_12534);
xor U17218 (N_17218,N_12521,N_13377);
nand U17219 (N_17219,N_13011,N_14364);
xor U17220 (N_17220,N_14059,N_13982);
xor U17221 (N_17221,N_12528,N_14675);
xnor U17222 (N_17222,N_13519,N_12566);
xor U17223 (N_17223,N_14818,N_12909);
nor U17224 (N_17224,N_14172,N_13501);
xor U17225 (N_17225,N_14920,N_13539);
and U17226 (N_17226,N_14583,N_14442);
nand U17227 (N_17227,N_14705,N_13932);
and U17228 (N_17228,N_13246,N_14211);
or U17229 (N_17229,N_13791,N_13348);
xnor U17230 (N_17230,N_14679,N_13522);
and U17231 (N_17231,N_13843,N_12559);
nand U17232 (N_17232,N_13366,N_12751);
nor U17233 (N_17233,N_13290,N_13749);
nor U17234 (N_17234,N_14549,N_12629);
nand U17235 (N_17235,N_13953,N_14835);
or U17236 (N_17236,N_12627,N_14785);
xor U17237 (N_17237,N_12772,N_12665);
xor U17238 (N_17238,N_13168,N_14413);
or U17239 (N_17239,N_14595,N_12507);
nor U17240 (N_17240,N_14097,N_12658);
nor U17241 (N_17241,N_13202,N_12747);
or U17242 (N_17242,N_12517,N_13181);
xnor U17243 (N_17243,N_13984,N_13291);
nand U17244 (N_17244,N_13585,N_13446);
or U17245 (N_17245,N_14895,N_12701);
nor U17246 (N_17246,N_14738,N_14442);
nand U17247 (N_17247,N_13081,N_14177);
and U17248 (N_17248,N_14332,N_14167);
nor U17249 (N_17249,N_13552,N_14801);
xor U17250 (N_17250,N_12850,N_14123);
or U17251 (N_17251,N_12525,N_13994);
xnor U17252 (N_17252,N_12895,N_13241);
nor U17253 (N_17253,N_14918,N_14007);
or U17254 (N_17254,N_13837,N_13513);
nand U17255 (N_17255,N_13113,N_14471);
or U17256 (N_17256,N_14568,N_13233);
nand U17257 (N_17257,N_14492,N_14506);
nor U17258 (N_17258,N_13586,N_13380);
nor U17259 (N_17259,N_13321,N_14478);
xor U17260 (N_17260,N_14737,N_14682);
or U17261 (N_17261,N_13574,N_13727);
nor U17262 (N_17262,N_14212,N_14513);
and U17263 (N_17263,N_13813,N_13261);
nor U17264 (N_17264,N_14334,N_13272);
xor U17265 (N_17265,N_13134,N_14876);
or U17266 (N_17266,N_14429,N_13352);
xnor U17267 (N_17267,N_13773,N_13102);
nand U17268 (N_17268,N_14424,N_14761);
or U17269 (N_17269,N_13891,N_13569);
and U17270 (N_17270,N_13986,N_12895);
nand U17271 (N_17271,N_13806,N_14034);
and U17272 (N_17272,N_13299,N_13470);
nand U17273 (N_17273,N_14387,N_13069);
nor U17274 (N_17274,N_12790,N_14212);
and U17275 (N_17275,N_14827,N_14223);
nor U17276 (N_17276,N_13614,N_13509);
nand U17277 (N_17277,N_13875,N_14588);
xnor U17278 (N_17278,N_14596,N_13696);
or U17279 (N_17279,N_13972,N_13613);
nor U17280 (N_17280,N_13233,N_14254);
nor U17281 (N_17281,N_14244,N_13502);
xor U17282 (N_17282,N_14399,N_12901);
or U17283 (N_17283,N_13210,N_14519);
nor U17284 (N_17284,N_12764,N_14994);
nand U17285 (N_17285,N_12522,N_14088);
or U17286 (N_17286,N_12709,N_14807);
xor U17287 (N_17287,N_14867,N_13006);
nor U17288 (N_17288,N_13309,N_14485);
and U17289 (N_17289,N_14387,N_14510);
and U17290 (N_17290,N_13583,N_13838);
xnor U17291 (N_17291,N_14153,N_13857);
and U17292 (N_17292,N_13785,N_14793);
nor U17293 (N_17293,N_13316,N_12545);
or U17294 (N_17294,N_14190,N_12641);
nor U17295 (N_17295,N_13306,N_14395);
nand U17296 (N_17296,N_14777,N_12618);
nor U17297 (N_17297,N_14349,N_12724);
or U17298 (N_17298,N_13965,N_13598);
and U17299 (N_17299,N_12620,N_13333);
nor U17300 (N_17300,N_14738,N_13030);
and U17301 (N_17301,N_12521,N_12682);
or U17302 (N_17302,N_14807,N_12710);
nor U17303 (N_17303,N_14799,N_13264);
nor U17304 (N_17304,N_13256,N_14702);
nand U17305 (N_17305,N_14921,N_12963);
nand U17306 (N_17306,N_13096,N_13693);
and U17307 (N_17307,N_14824,N_14943);
and U17308 (N_17308,N_13063,N_13603);
xor U17309 (N_17309,N_13071,N_12878);
nor U17310 (N_17310,N_12955,N_14034);
and U17311 (N_17311,N_14900,N_14301);
nor U17312 (N_17312,N_13063,N_13031);
xor U17313 (N_17313,N_13140,N_14217);
or U17314 (N_17314,N_14406,N_14561);
nor U17315 (N_17315,N_13239,N_13816);
nand U17316 (N_17316,N_13010,N_14940);
or U17317 (N_17317,N_13959,N_13191);
nor U17318 (N_17318,N_14865,N_14151);
and U17319 (N_17319,N_12702,N_14693);
or U17320 (N_17320,N_13266,N_14151);
nand U17321 (N_17321,N_13326,N_13942);
and U17322 (N_17322,N_14468,N_12831);
nand U17323 (N_17323,N_14149,N_13559);
nor U17324 (N_17324,N_14929,N_13661);
nand U17325 (N_17325,N_14384,N_13235);
or U17326 (N_17326,N_14227,N_14421);
and U17327 (N_17327,N_13625,N_13875);
or U17328 (N_17328,N_13585,N_14036);
nand U17329 (N_17329,N_14573,N_13994);
xnor U17330 (N_17330,N_13972,N_14372);
nor U17331 (N_17331,N_13246,N_13362);
xnor U17332 (N_17332,N_14618,N_14418);
or U17333 (N_17333,N_12555,N_14864);
nand U17334 (N_17334,N_13213,N_14306);
xnor U17335 (N_17335,N_14242,N_14133);
or U17336 (N_17336,N_13864,N_13476);
xnor U17337 (N_17337,N_13418,N_13822);
nand U17338 (N_17338,N_14580,N_14776);
and U17339 (N_17339,N_13300,N_14090);
nor U17340 (N_17340,N_14354,N_14820);
and U17341 (N_17341,N_14851,N_14368);
and U17342 (N_17342,N_13549,N_14459);
nand U17343 (N_17343,N_14961,N_14926);
nor U17344 (N_17344,N_12868,N_13464);
or U17345 (N_17345,N_13717,N_13591);
nor U17346 (N_17346,N_13019,N_14240);
xnor U17347 (N_17347,N_14123,N_14138);
nand U17348 (N_17348,N_13045,N_13566);
or U17349 (N_17349,N_14027,N_14720);
xnor U17350 (N_17350,N_14207,N_13846);
or U17351 (N_17351,N_14877,N_12637);
xnor U17352 (N_17352,N_13036,N_13091);
xnor U17353 (N_17353,N_12515,N_13889);
or U17354 (N_17354,N_14553,N_12673);
or U17355 (N_17355,N_12910,N_14154);
nor U17356 (N_17356,N_14635,N_13487);
xor U17357 (N_17357,N_13240,N_13578);
nor U17358 (N_17358,N_13267,N_14290);
xor U17359 (N_17359,N_12893,N_13913);
or U17360 (N_17360,N_14064,N_14844);
nand U17361 (N_17361,N_12909,N_14058);
xnor U17362 (N_17362,N_13366,N_13055);
or U17363 (N_17363,N_13151,N_12957);
and U17364 (N_17364,N_13866,N_12766);
nor U17365 (N_17365,N_14432,N_13862);
and U17366 (N_17366,N_14115,N_14595);
xor U17367 (N_17367,N_14418,N_13516);
xnor U17368 (N_17368,N_12730,N_13621);
or U17369 (N_17369,N_12785,N_13022);
and U17370 (N_17370,N_12914,N_13527);
xor U17371 (N_17371,N_14489,N_13295);
xnor U17372 (N_17372,N_12534,N_14817);
nor U17373 (N_17373,N_14642,N_12683);
nand U17374 (N_17374,N_14743,N_14253);
nand U17375 (N_17375,N_13574,N_14312);
nor U17376 (N_17376,N_14945,N_13512);
nor U17377 (N_17377,N_12779,N_14818);
nand U17378 (N_17378,N_12798,N_13402);
nor U17379 (N_17379,N_13669,N_12554);
xnor U17380 (N_17380,N_13068,N_12504);
nand U17381 (N_17381,N_14393,N_13696);
nand U17382 (N_17382,N_12890,N_13998);
nor U17383 (N_17383,N_12777,N_12769);
xor U17384 (N_17384,N_14272,N_14385);
nor U17385 (N_17385,N_13923,N_14597);
nor U17386 (N_17386,N_14950,N_13082);
xor U17387 (N_17387,N_14060,N_12849);
and U17388 (N_17388,N_13653,N_14680);
or U17389 (N_17389,N_13221,N_13400);
nand U17390 (N_17390,N_14534,N_14008);
nand U17391 (N_17391,N_14243,N_13117);
xor U17392 (N_17392,N_14263,N_13428);
and U17393 (N_17393,N_12837,N_14936);
and U17394 (N_17394,N_14707,N_13891);
nor U17395 (N_17395,N_14003,N_14664);
xor U17396 (N_17396,N_14241,N_14322);
and U17397 (N_17397,N_14171,N_13871);
nand U17398 (N_17398,N_14426,N_13128);
or U17399 (N_17399,N_13938,N_13061);
nand U17400 (N_17400,N_14481,N_13638);
or U17401 (N_17401,N_12845,N_14973);
xor U17402 (N_17402,N_13571,N_14976);
xor U17403 (N_17403,N_13472,N_12728);
nand U17404 (N_17404,N_14893,N_12606);
xor U17405 (N_17405,N_14670,N_14357);
or U17406 (N_17406,N_14614,N_13529);
nor U17407 (N_17407,N_14668,N_12759);
nor U17408 (N_17408,N_14091,N_12843);
nand U17409 (N_17409,N_14905,N_14191);
nor U17410 (N_17410,N_14480,N_13896);
or U17411 (N_17411,N_12956,N_14354);
or U17412 (N_17412,N_14850,N_13217);
xor U17413 (N_17413,N_13013,N_14700);
nand U17414 (N_17414,N_13059,N_12830);
nand U17415 (N_17415,N_14451,N_12606);
and U17416 (N_17416,N_14823,N_14859);
nor U17417 (N_17417,N_14771,N_12594);
xnor U17418 (N_17418,N_14790,N_13145);
nor U17419 (N_17419,N_14074,N_14715);
or U17420 (N_17420,N_13509,N_14340);
and U17421 (N_17421,N_13906,N_12787);
nand U17422 (N_17422,N_13547,N_14974);
nand U17423 (N_17423,N_12655,N_13744);
xnor U17424 (N_17424,N_14018,N_14056);
and U17425 (N_17425,N_12531,N_14108);
nor U17426 (N_17426,N_13814,N_12651);
xnor U17427 (N_17427,N_14499,N_14453);
or U17428 (N_17428,N_14927,N_13285);
xnor U17429 (N_17429,N_14096,N_14522);
xnor U17430 (N_17430,N_13568,N_12931);
xnor U17431 (N_17431,N_14994,N_14646);
nand U17432 (N_17432,N_12810,N_13109);
or U17433 (N_17433,N_13517,N_14584);
nand U17434 (N_17434,N_13075,N_12673);
nor U17435 (N_17435,N_14703,N_14808);
nor U17436 (N_17436,N_14150,N_13047);
nor U17437 (N_17437,N_14456,N_14605);
or U17438 (N_17438,N_13259,N_14342);
or U17439 (N_17439,N_14896,N_13157);
and U17440 (N_17440,N_14427,N_12984);
nor U17441 (N_17441,N_14968,N_14947);
xnor U17442 (N_17442,N_13480,N_13916);
nor U17443 (N_17443,N_14237,N_13647);
nor U17444 (N_17444,N_14720,N_13987);
or U17445 (N_17445,N_14701,N_14452);
xnor U17446 (N_17446,N_13511,N_14032);
nor U17447 (N_17447,N_13340,N_13646);
or U17448 (N_17448,N_14422,N_14233);
nand U17449 (N_17449,N_13598,N_14067);
nor U17450 (N_17450,N_13489,N_14239);
and U17451 (N_17451,N_14773,N_14926);
and U17452 (N_17452,N_13607,N_14696);
xor U17453 (N_17453,N_14956,N_12555);
xnor U17454 (N_17454,N_13145,N_12938);
nor U17455 (N_17455,N_12603,N_14307);
nor U17456 (N_17456,N_14736,N_13934);
nand U17457 (N_17457,N_14489,N_13671);
xnor U17458 (N_17458,N_13643,N_14307);
and U17459 (N_17459,N_14431,N_13003);
nand U17460 (N_17460,N_13335,N_13114);
nor U17461 (N_17461,N_12722,N_14713);
nor U17462 (N_17462,N_13211,N_14995);
nor U17463 (N_17463,N_14627,N_12997);
nand U17464 (N_17464,N_14861,N_14453);
xnor U17465 (N_17465,N_14394,N_14856);
nand U17466 (N_17466,N_13618,N_14147);
nor U17467 (N_17467,N_12700,N_14713);
nand U17468 (N_17468,N_14586,N_14905);
xor U17469 (N_17469,N_13330,N_13103);
xnor U17470 (N_17470,N_13637,N_13133);
or U17471 (N_17471,N_13536,N_14198);
or U17472 (N_17472,N_13618,N_14056);
or U17473 (N_17473,N_12767,N_13522);
nor U17474 (N_17474,N_12559,N_12500);
xor U17475 (N_17475,N_13738,N_12556);
nand U17476 (N_17476,N_14407,N_14593);
and U17477 (N_17477,N_13797,N_14136);
or U17478 (N_17478,N_14931,N_14585);
or U17479 (N_17479,N_14135,N_13114);
xor U17480 (N_17480,N_12697,N_14239);
nand U17481 (N_17481,N_13890,N_13413);
and U17482 (N_17482,N_12904,N_13019);
nand U17483 (N_17483,N_13161,N_14342);
nand U17484 (N_17484,N_14781,N_12703);
nand U17485 (N_17485,N_14310,N_14093);
xnor U17486 (N_17486,N_13217,N_14649);
nor U17487 (N_17487,N_13903,N_14240);
xnor U17488 (N_17488,N_14023,N_12708);
nor U17489 (N_17489,N_14224,N_13459);
nor U17490 (N_17490,N_12519,N_12790);
nand U17491 (N_17491,N_13121,N_14685);
or U17492 (N_17492,N_14196,N_14614);
and U17493 (N_17493,N_13124,N_13120);
xnor U17494 (N_17494,N_12618,N_13299);
nand U17495 (N_17495,N_12538,N_14991);
or U17496 (N_17496,N_13449,N_13130);
or U17497 (N_17497,N_14908,N_13319);
or U17498 (N_17498,N_13303,N_12504);
nor U17499 (N_17499,N_14281,N_14946);
xor U17500 (N_17500,N_15112,N_16005);
xor U17501 (N_17501,N_15658,N_16408);
nand U17502 (N_17502,N_15134,N_17390);
or U17503 (N_17503,N_16645,N_16304);
or U17504 (N_17504,N_16729,N_16558);
nor U17505 (N_17505,N_16765,N_16837);
and U17506 (N_17506,N_15542,N_16014);
nor U17507 (N_17507,N_15297,N_15373);
nand U17508 (N_17508,N_16263,N_16887);
or U17509 (N_17509,N_15771,N_15032);
or U17510 (N_17510,N_16816,N_15946);
and U17511 (N_17511,N_17014,N_16423);
or U17512 (N_17512,N_16984,N_15507);
nor U17513 (N_17513,N_15033,N_15943);
xnor U17514 (N_17514,N_17017,N_17070);
nand U17515 (N_17515,N_15058,N_16202);
nand U17516 (N_17516,N_16495,N_15192);
xor U17517 (N_17517,N_15569,N_17009);
and U17518 (N_17518,N_15038,N_15661);
nand U17519 (N_17519,N_17444,N_17322);
and U17520 (N_17520,N_17059,N_16950);
nor U17521 (N_17521,N_17032,N_15017);
nor U17522 (N_17522,N_17026,N_15419);
nor U17523 (N_17523,N_16438,N_17308);
nor U17524 (N_17524,N_16492,N_16930);
nor U17525 (N_17525,N_17073,N_15921);
nor U17526 (N_17526,N_15422,N_15647);
and U17527 (N_17527,N_15166,N_16908);
and U17528 (N_17528,N_16786,N_16214);
xnor U17529 (N_17529,N_17450,N_17168);
xnor U17530 (N_17530,N_15342,N_15809);
nand U17531 (N_17531,N_16650,N_15572);
nor U17532 (N_17532,N_16971,N_17145);
nor U17533 (N_17533,N_16413,N_15235);
or U17534 (N_17534,N_16711,N_16384);
nand U17535 (N_17535,N_15355,N_15001);
nand U17536 (N_17536,N_16524,N_15805);
xnor U17537 (N_17537,N_15654,N_15836);
nand U17538 (N_17538,N_15552,N_16293);
nor U17539 (N_17539,N_16692,N_16195);
nand U17540 (N_17540,N_15719,N_16483);
xor U17541 (N_17541,N_15413,N_15434);
and U17542 (N_17542,N_15279,N_16493);
nand U17543 (N_17543,N_15894,N_16654);
and U17544 (N_17544,N_17021,N_15679);
xnor U17545 (N_17545,N_16453,N_16512);
nand U17546 (N_17546,N_15494,N_15837);
or U17547 (N_17547,N_15278,N_15874);
xor U17548 (N_17548,N_16457,N_16734);
nor U17549 (N_17549,N_16844,N_17300);
and U17550 (N_17550,N_15453,N_16383);
xor U17551 (N_17551,N_15315,N_15633);
nor U17552 (N_17552,N_15343,N_15376);
or U17553 (N_17553,N_15987,N_16078);
and U17554 (N_17554,N_15187,N_17056);
nor U17555 (N_17555,N_15920,N_16503);
xor U17556 (N_17556,N_16001,N_16600);
or U17557 (N_17557,N_16207,N_17051);
or U17558 (N_17558,N_17196,N_15349);
or U17559 (N_17559,N_17359,N_15902);
nor U17560 (N_17560,N_16802,N_15547);
xnor U17561 (N_17561,N_16647,N_16193);
nor U17562 (N_17562,N_17002,N_15834);
xnor U17563 (N_17563,N_17298,N_15177);
nor U17564 (N_17564,N_16069,N_16016);
and U17565 (N_17565,N_16003,N_16159);
xnor U17566 (N_17566,N_15175,N_16536);
nor U17567 (N_17567,N_16914,N_17183);
nand U17568 (N_17568,N_17116,N_17370);
xor U17569 (N_17569,N_15220,N_16220);
nor U17570 (N_17570,N_15872,N_16843);
xor U17571 (N_17571,N_16864,N_16826);
xor U17572 (N_17572,N_16993,N_15710);
nand U17573 (N_17573,N_16142,N_16222);
nand U17574 (N_17574,N_15833,N_15416);
xnor U17575 (N_17575,N_15474,N_15446);
xnor U17576 (N_17576,N_16388,N_16247);
xor U17577 (N_17577,N_16534,N_15986);
nor U17578 (N_17578,N_15445,N_15178);
xnor U17579 (N_17579,N_15682,N_15160);
nor U17580 (N_17580,N_15308,N_17166);
nand U17581 (N_17581,N_15319,N_15199);
nand U17582 (N_17582,N_16450,N_15486);
nor U17583 (N_17583,N_17256,N_17023);
nand U17584 (N_17584,N_16616,N_15736);
and U17585 (N_17585,N_16023,N_16559);
xnor U17586 (N_17586,N_15994,N_17352);
xnor U17587 (N_17587,N_16801,N_15966);
nor U17588 (N_17588,N_16609,N_15483);
xor U17589 (N_17589,N_15609,N_16302);
or U17590 (N_17590,N_16305,N_16259);
or U17591 (N_17591,N_15357,N_15176);
xor U17592 (N_17592,N_15251,N_17001);
nor U17593 (N_17593,N_17355,N_16225);
nand U17594 (N_17594,N_17197,N_17101);
nand U17595 (N_17595,N_16145,N_17118);
nor U17596 (N_17596,N_15972,N_17003);
nand U17597 (N_17597,N_16052,N_15186);
and U17598 (N_17598,N_16219,N_16319);
xnor U17599 (N_17599,N_15604,N_16648);
xnor U17600 (N_17600,N_16507,N_17195);
nor U17601 (N_17601,N_16596,N_17131);
nor U17602 (N_17602,N_17386,N_16925);
and U17603 (N_17603,N_17278,N_17123);
xor U17604 (N_17604,N_16015,N_16291);
or U17605 (N_17605,N_15583,N_17206);
or U17606 (N_17606,N_15551,N_15287);
and U17607 (N_17607,N_15888,N_15195);
nand U17608 (N_17608,N_16968,N_15852);
nor U17609 (N_17609,N_15523,N_17072);
and U17610 (N_17610,N_15020,N_16190);
or U17611 (N_17611,N_17012,N_15348);
nor U17612 (N_17612,N_17143,N_16352);
or U17613 (N_17613,N_15640,N_15580);
xor U17614 (N_17614,N_15992,N_16415);
and U17615 (N_17615,N_15127,N_17043);
nand U17616 (N_17616,N_15889,N_16687);
and U17617 (N_17617,N_15293,N_16212);
or U17618 (N_17618,N_16924,N_16994);
nor U17619 (N_17619,N_15900,N_15923);
xor U17620 (N_17620,N_16331,N_16748);
or U17621 (N_17621,N_15708,N_15141);
xnor U17622 (N_17622,N_15075,N_16674);
nand U17623 (N_17623,N_16206,N_16705);
nor U17624 (N_17624,N_16235,N_15189);
or U17625 (N_17625,N_16424,N_16763);
or U17626 (N_17626,N_15694,N_15487);
nand U17627 (N_17627,N_15937,N_16497);
nand U17628 (N_17628,N_16550,N_15490);
nor U17629 (N_17629,N_16511,N_17063);
xor U17630 (N_17630,N_15709,N_16970);
nand U17631 (N_17631,N_15263,N_15458);
nand U17632 (N_17632,N_16253,N_16165);
xor U17633 (N_17633,N_16975,N_15745);
and U17634 (N_17634,N_15047,N_15121);
or U17635 (N_17635,N_15575,N_15151);
nand U17636 (N_17636,N_17328,N_15859);
nor U17637 (N_17637,N_16756,N_15299);
nand U17638 (N_17638,N_16552,N_15678);
xor U17639 (N_17639,N_15261,N_15692);
or U17640 (N_17640,N_15835,N_16642);
xor U17641 (N_17641,N_16619,N_17269);
and U17642 (N_17642,N_16731,N_15497);
or U17643 (N_17643,N_16137,N_16876);
xor U17644 (N_17644,N_17453,N_15450);
or U17645 (N_17645,N_17204,N_15699);
and U17646 (N_17646,N_16581,N_17120);
or U17647 (N_17647,N_16272,N_15147);
or U17648 (N_17648,N_15431,N_15945);
xor U17649 (N_17649,N_15275,N_16443);
nor U17650 (N_17650,N_15788,N_15706);
and U17651 (N_17651,N_17011,N_17376);
xnor U17652 (N_17652,N_15179,N_16761);
xnor U17653 (N_17653,N_17398,N_15049);
and U17654 (N_17654,N_16894,N_15008);
or U17655 (N_17655,N_16872,N_15707);
nand U17656 (N_17656,N_16258,N_16999);
and U17657 (N_17657,N_16656,N_17348);
or U17658 (N_17658,N_15917,N_16744);
and U17659 (N_17659,N_17454,N_16580);
and U17660 (N_17660,N_16311,N_17046);
xor U17661 (N_17661,N_16560,N_15417);
and U17662 (N_17662,N_17329,N_17174);
nor U17663 (N_17663,N_17024,N_16615);
nor U17664 (N_17664,N_16431,N_15755);
xor U17665 (N_17665,N_15282,N_15798);
nand U17666 (N_17666,N_16152,N_15104);
xor U17667 (N_17667,N_15120,N_15886);
nand U17668 (N_17668,N_17165,N_15356);
or U17669 (N_17669,N_15586,N_17483);
or U17670 (N_17670,N_17281,N_15555);
and U17671 (N_17671,N_17464,N_16860);
and U17672 (N_17672,N_16898,N_15584);
nor U17673 (N_17673,N_17122,N_15562);
and U17674 (N_17674,N_15600,N_15242);
and U17675 (N_17675,N_16261,N_16625);
and U17676 (N_17676,N_15864,N_17288);
or U17677 (N_17677,N_16481,N_15934);
nand U17678 (N_17678,N_17147,N_15025);
xnor U17679 (N_17679,N_15044,N_15098);
nand U17680 (N_17680,N_16835,N_16571);
nand U17681 (N_17681,N_15004,N_17305);
xnor U17682 (N_17682,N_15146,N_15782);
nor U17683 (N_17683,N_15757,N_15062);
xor U17684 (N_17684,N_16449,N_15061);
or U17685 (N_17685,N_15642,N_16301);
nand U17686 (N_17686,N_15607,N_15068);
or U17687 (N_17687,N_15082,N_15789);
xor U17688 (N_17688,N_16125,N_17261);
nand U17689 (N_17689,N_16593,N_17358);
nor U17690 (N_17690,N_16646,N_16082);
nand U17691 (N_17691,N_17069,N_16274);
nand U17692 (N_17692,N_15720,N_17282);
or U17693 (N_17693,N_17339,N_15631);
nand U17694 (N_17694,N_15423,N_15333);
xor U17695 (N_17695,N_17130,N_16962);
or U17696 (N_17696,N_15262,N_17470);
nor U17697 (N_17697,N_16653,N_15103);
xor U17698 (N_17698,N_17285,N_15668);
xnor U17699 (N_17699,N_17488,N_17252);
and U17700 (N_17700,N_17462,N_16127);
nor U17701 (N_17701,N_15123,N_17277);
xnor U17702 (N_17702,N_16547,N_16806);
xor U17703 (N_17703,N_15245,N_15997);
nor U17704 (N_17704,N_15045,N_16979);
nor U17705 (N_17705,N_17193,N_15639);
or U17706 (N_17706,N_16102,N_17140);
xor U17707 (N_17707,N_17409,N_15398);
xor U17708 (N_17708,N_16562,N_15036);
nor U17709 (N_17709,N_15107,N_15421);
and U17710 (N_17710,N_16330,N_15233);
nor U17711 (N_17711,N_15399,N_15167);
xor U17712 (N_17712,N_17034,N_16861);
nor U17713 (N_17713,N_16484,N_16364);
or U17714 (N_17714,N_15406,N_15999);
and U17715 (N_17715,N_16267,N_16807);
nor U17716 (N_17716,N_16133,N_16009);
xnor U17717 (N_17717,N_17227,N_17031);
xor U17718 (N_17718,N_16838,N_15887);
xor U17719 (N_17719,N_16480,N_15521);
or U17720 (N_17720,N_15460,N_16162);
nor U17721 (N_17721,N_16945,N_16264);
nand U17722 (N_17722,N_15285,N_16168);
nor U17723 (N_17723,N_15741,N_16537);
xnor U17724 (N_17724,N_16758,N_15689);
nand U17725 (N_17725,N_17461,N_16915);
xor U17726 (N_17726,N_16521,N_15129);
nand U17727 (N_17727,N_16266,N_15813);
or U17728 (N_17728,N_16494,N_15526);
nor U17729 (N_17729,N_15392,N_17138);
or U17730 (N_17730,N_15983,N_15196);
or U17731 (N_17731,N_15725,N_16691);
nand U17732 (N_17732,N_15630,N_17291);
or U17733 (N_17733,N_16077,N_15394);
and U17734 (N_17734,N_15712,N_16396);
or U17735 (N_17735,N_16848,N_15185);
or U17736 (N_17736,N_16324,N_16091);
xnor U17737 (N_17737,N_16004,N_17267);
xnor U17738 (N_17738,N_16759,N_17296);
nor U17739 (N_17739,N_15685,N_15014);
and U17740 (N_17740,N_15467,N_16607);
or U17741 (N_17741,N_16671,N_16868);
nor U17742 (N_17742,N_16446,N_16502);
nor U17743 (N_17743,N_16587,N_16632);
nand U17744 (N_17744,N_16878,N_15778);
nand U17745 (N_17745,N_17452,N_16695);
or U17746 (N_17746,N_16961,N_15231);
nand U17747 (N_17747,N_16386,N_16948);
and U17748 (N_17748,N_16238,N_17090);
nor U17749 (N_17749,N_16939,N_16474);
xnor U17750 (N_17750,N_16467,N_16518);
or U17751 (N_17751,N_16044,N_16049);
nor U17752 (N_17752,N_16066,N_16074);
nor U17753 (N_17753,N_16509,N_16278);
nand U17754 (N_17754,N_16942,N_15982);
nand U17755 (N_17755,N_15686,N_16972);
nand U17756 (N_17756,N_16046,N_16076);
nand U17757 (N_17757,N_16956,N_15544);
nand U17758 (N_17758,N_15078,N_16753);
and U17759 (N_17759,N_16505,N_17173);
nand U17760 (N_17760,N_16895,N_15165);
nor U17761 (N_17761,N_17037,N_16870);
nor U17762 (N_17762,N_16426,N_17455);
nor U17763 (N_17763,N_15265,N_17498);
and U17764 (N_17764,N_16556,N_16842);
nor U17765 (N_17765,N_16444,N_16136);
and U17766 (N_17766,N_16730,N_16809);
or U17767 (N_17767,N_15664,N_15126);
or U17768 (N_17768,N_15746,N_17445);
xor U17769 (N_17769,N_16209,N_15698);
xnor U17770 (N_17770,N_15320,N_16610);
nand U17771 (N_17771,N_15635,N_16766);
or U17772 (N_17772,N_16201,N_15227);
and U17773 (N_17773,N_15158,N_15800);
nand U17774 (N_17774,N_17020,N_16935);
xnor U17775 (N_17775,N_15198,N_15236);
xor U17776 (N_17776,N_15095,N_16223);
nand U17777 (N_17777,N_15200,N_16134);
nand U17778 (N_17778,N_16932,N_16789);
nand U17779 (N_17779,N_16416,N_15878);
or U17780 (N_17780,N_15202,N_15513);
nand U17781 (N_17781,N_17071,N_16108);
nand U17782 (N_17782,N_16146,N_17229);
xor U17783 (N_17783,N_17345,N_16670);
nor U17784 (N_17784,N_15850,N_17133);
or U17785 (N_17785,N_17258,N_15340);
nand U17786 (N_17786,N_15271,N_17319);
nand U17787 (N_17787,N_15669,N_15159);
xor U17788 (N_17788,N_17436,N_16829);
xor U17789 (N_17789,N_15076,N_15305);
and U17790 (N_17790,N_16831,N_17373);
nor U17791 (N_17791,N_16815,N_15776);
nor U17792 (N_17792,N_16114,N_17030);
xor U17793 (N_17793,N_16353,N_15915);
or U17794 (N_17794,N_16459,N_16469);
xnor U17795 (N_17795,N_15660,N_16166);
nand U17796 (N_17796,N_15870,N_16812);
nor U17797 (N_17797,N_15286,N_17112);
or U17798 (N_17798,N_15335,N_15479);
xor U17799 (N_17799,N_16439,N_16900);
nor U17800 (N_17800,N_16197,N_15223);
nand U17801 (N_17801,N_15313,N_15307);
xnor U17802 (N_17802,N_15732,N_15737);
and U17803 (N_17803,N_16393,N_16362);
nor U17804 (N_17804,N_15426,N_15388);
nor U17805 (N_17805,N_15904,N_16406);
nand U17806 (N_17806,N_15488,N_15442);
or U17807 (N_17807,N_15427,N_15688);
or U17808 (N_17808,N_17045,N_16629);
nor U17809 (N_17809,N_15056,N_15430);
nand U17810 (N_17810,N_16740,N_15046);
nor U17811 (N_17811,N_17110,N_16681);
xor U17812 (N_17812,N_15701,N_17437);
nor U17813 (N_17813,N_15255,N_16840);
or U17814 (N_17814,N_16434,N_17270);
xor U17815 (N_17815,N_17055,N_16138);
xor U17816 (N_17816,N_16564,N_15081);
or U17817 (N_17817,N_16401,N_15256);
nand U17818 (N_17818,N_16392,N_16982);
and U17819 (N_17819,N_15324,N_15283);
and U17820 (N_17820,N_17401,N_16087);
nand U17821 (N_17821,N_16067,N_17154);
nand U17822 (N_17822,N_16240,N_15473);
xor U17823 (N_17823,N_16095,N_17367);
xnor U17824 (N_17824,N_16333,N_16429);
and U17825 (N_17825,N_16030,N_15155);
or U17826 (N_17826,N_16965,N_15854);
and U17827 (N_17827,N_16940,N_16833);
or U17828 (N_17828,N_15024,N_17335);
xnor U17829 (N_17829,N_15140,N_16698);
xor U17830 (N_17830,N_15119,N_15139);
nor U17831 (N_17831,N_16187,N_17006);
or U17832 (N_17832,N_17205,N_17054);
or U17833 (N_17833,N_15469,N_15926);
nand U17834 (N_17834,N_17244,N_15270);
nor U17835 (N_17835,N_16199,N_15527);
xnor U17836 (N_17836,N_17363,N_15462);
xnor U17837 (N_17837,N_16725,N_15363);
nand U17838 (N_17838,N_16182,N_17231);
xor U17839 (N_17839,N_16832,N_16776);
nand U17840 (N_17840,N_16425,N_15791);
or U17841 (N_17841,N_17389,N_16022);
nor U17842 (N_17842,N_16418,N_15831);
nor U17843 (N_17843,N_16501,N_16839);
nand U17844 (N_17844,N_15978,N_15705);
nor U17845 (N_17845,N_16751,N_15832);
xor U17846 (N_17846,N_16042,N_17347);
or U17847 (N_17847,N_16229,N_15211);
or U17848 (N_17848,N_16255,N_16144);
or U17849 (N_17849,N_15425,N_17114);
nor U17850 (N_17850,N_16419,N_16120);
and U17851 (N_17851,N_16797,N_16539);
or U17852 (N_17852,N_16742,N_17167);
and U17853 (N_17853,N_16281,N_16499);
nand U17854 (N_17854,N_16325,N_15637);
or U17855 (N_17855,N_16340,N_16334);
nor U17856 (N_17856,N_16399,N_15499);
xnor U17857 (N_17857,N_15015,N_15949);
xor U17858 (N_17858,N_17218,N_16923);
nand U17859 (N_17859,N_17184,N_15135);
nor U17860 (N_17860,N_16586,N_15821);
and U17861 (N_17861,N_16062,N_15232);
or U17862 (N_17862,N_16111,N_16527);
xor U17863 (N_17863,N_15128,N_16997);
nand U17864 (N_17864,N_15704,N_15644);
or U17865 (N_17865,N_16055,N_16496);
xnor U17866 (N_17866,N_16465,N_17253);
nand U17867 (N_17867,N_17465,N_15131);
or U17868 (N_17868,N_16880,N_17463);
or U17869 (N_17869,N_15492,N_15407);
or U17870 (N_17870,N_15762,N_15013);
nor U17871 (N_17871,N_17257,N_15226);
nand U17872 (N_17872,N_16327,N_15601);
and U17873 (N_17873,N_17460,N_17326);
and U17874 (N_17874,N_17128,N_16471);
xnor U17875 (N_17875,N_17321,N_16661);
nor U17876 (N_17876,N_16828,N_15659);
or U17877 (N_17877,N_16799,N_16929);
nand U17878 (N_17878,N_16792,N_16633);
xor U17879 (N_17879,N_15561,N_16658);
nor U17880 (N_17880,N_15006,N_15498);
nand U17881 (N_17881,N_15344,N_15770);
and U17882 (N_17882,N_17216,N_15329);
nand U17883 (N_17883,N_16462,N_17259);
nand U17884 (N_17884,N_16227,N_15893);
and U17885 (N_17885,N_15534,N_15804);
xor U17886 (N_17886,N_15898,N_15616);
nor U17887 (N_17887,N_15774,N_15351);
nand U17888 (N_17888,N_17094,N_15034);
nor U17889 (N_17889,N_16978,N_15420);
nand U17890 (N_17890,N_16315,N_16251);
and U17891 (N_17891,N_15424,N_17384);
and U17892 (N_17892,N_16904,N_17236);
and U17893 (N_17893,N_17406,N_16375);
nand U17894 (N_17894,N_17481,N_16702);
and U17895 (N_17895,N_17357,N_16037);
or U17896 (N_17896,N_15519,N_16871);
nand U17897 (N_17897,N_15009,N_15817);
and U17898 (N_17898,N_15368,N_16321);
and U17899 (N_17899,N_16184,N_17303);
nand U17900 (N_17900,N_16105,N_16522);
nor U17901 (N_17901,N_16475,N_16176);
and U17902 (N_17902,N_17441,N_16417);
nand U17903 (N_17903,N_16139,N_16714);
nand U17904 (N_17904,N_15309,N_17474);
nor U17905 (N_17905,N_17198,N_17180);
and U17906 (N_17906,N_16525,N_15750);
nand U17907 (N_17907,N_16360,N_15086);
or U17908 (N_17908,N_16047,N_15827);
xnor U17909 (N_17909,N_16541,N_15883);
nor U17910 (N_17910,N_17005,N_16048);
nand U17911 (N_17911,N_15629,N_15026);
and U17912 (N_17912,N_17405,N_16174);
nor U17913 (N_17913,N_17410,N_15259);
or U17914 (N_17914,N_15288,N_16208);
xor U17915 (N_17915,N_15191,N_15919);
nand U17916 (N_17916,N_16680,N_15622);
xnor U17917 (N_17917,N_15332,N_16421);
or U17918 (N_17918,N_15518,N_17274);
nor U17919 (N_17919,N_17113,N_16218);
nand U17920 (N_17920,N_16099,N_17325);
or U17921 (N_17921,N_15336,N_15744);
nor U17922 (N_17922,N_15645,N_15302);
nor U17923 (N_17923,N_16020,N_15940);
nand U17924 (N_17924,N_17098,N_15150);
nor U17925 (N_17925,N_15760,N_17052);
xnor U17926 (N_17926,N_15216,N_16036);
nor U17927 (N_17927,N_15448,N_16735);
xor U17928 (N_17928,N_16365,N_16628);
nor U17929 (N_17929,N_16988,N_16779);
and U17930 (N_17930,N_16545,N_16154);
nor U17931 (N_17931,N_16707,N_17310);
and U17932 (N_17932,N_16025,N_16370);
or U17933 (N_17933,N_15385,N_15478);
nand U17934 (N_17934,N_15632,N_15005);
nor U17935 (N_17935,N_15577,N_16685);
xor U17936 (N_17936,N_16463,N_16589);
or U17937 (N_17937,N_16081,N_16853);
and U17938 (N_17938,N_17396,N_15454);
nand U17939 (N_17939,N_15249,N_15892);
or U17940 (N_17940,N_15048,N_17142);
and U17941 (N_17941,N_15144,N_16158);
or U17942 (N_17942,N_16299,N_15266);
nor U17943 (N_17943,N_17019,N_16411);
xor U17944 (N_17944,N_15721,N_15390);
or U17945 (N_17945,N_16189,N_16712);
nand U17946 (N_17946,N_15443,N_15316);
nand U17947 (N_17947,N_15794,N_15436);
nand U17948 (N_17948,N_15754,N_15053);
xor U17949 (N_17949,N_17179,N_16204);
nand U17950 (N_17950,N_16745,N_17399);
and U17951 (N_17951,N_16599,N_16122);
or U17952 (N_17952,N_17082,N_15927);
nor U17953 (N_17953,N_15525,N_17178);
nand U17954 (N_17954,N_15444,N_15291);
nand U17955 (N_17955,N_15565,N_15793);
nand U17956 (N_17956,N_16132,N_17353);
or U17957 (N_17957,N_15868,N_17459);
or U17958 (N_17958,N_16770,N_16285);
or U17959 (N_17959,N_15952,N_16768);
or U17960 (N_17960,N_16862,N_15801);
nor U17961 (N_17961,N_16310,N_16841);
nor U17962 (N_17962,N_15403,N_15603);
xnor U17963 (N_17963,N_16228,N_15579);
xnor U17964 (N_17964,N_17234,N_15856);
or U17965 (N_17965,N_15244,N_17286);
xnor U17966 (N_17966,N_15021,N_15779);
or U17967 (N_17967,N_16675,N_15825);
nand U17968 (N_17968,N_17170,N_15914);
nor U17969 (N_17969,N_16913,N_16949);
nor U17970 (N_17970,N_15085,N_15570);
nand U17971 (N_17971,N_15785,N_16135);
nand U17972 (N_17972,N_17172,N_16983);
and U17973 (N_17973,N_15558,N_16306);
xnor U17974 (N_17974,N_16821,N_15777);
xor U17975 (N_17975,N_16919,N_15596);
nor U17976 (N_17976,N_16641,N_17414);
and U17977 (N_17977,N_16854,N_16275);
and U17978 (N_17978,N_16173,N_15132);
and U17979 (N_17979,N_15480,N_15060);
xnor U17980 (N_17980,N_16367,N_17490);
or U17981 (N_17981,N_15163,N_15371);
nand U17982 (N_17982,N_16314,N_16447);
and U17983 (N_17983,N_15472,N_17494);
or U17984 (N_17984,N_17327,N_16164);
and U17985 (N_17985,N_15387,N_17155);
or U17986 (N_17986,N_17217,N_17187);
and U17987 (N_17987,N_16963,N_16409);
nor U17988 (N_17988,N_16644,N_15676);
xnor U17989 (N_17989,N_17027,N_17408);
nand U17990 (N_17990,N_15840,N_17323);
xnor U17991 (N_17991,N_15331,N_17220);
nand U17992 (N_17992,N_17162,N_16412);
or U17993 (N_17993,N_16252,N_15369);
or U17994 (N_17994,N_15208,N_15374);
xor U17995 (N_17995,N_15602,N_15181);
nor U17996 (N_17996,N_17320,N_16798);
and U17997 (N_17997,N_15411,N_17480);
and U17998 (N_17998,N_17421,N_15576);
nor U17999 (N_17999,N_15384,N_17158);
and U18000 (N_18000,N_16764,N_15941);
xor U18001 (N_18001,N_15317,N_16205);
xor U18002 (N_18002,N_15590,N_17139);
nand U18003 (N_18003,N_16976,N_16995);
nor U18004 (N_18004,N_16116,N_16323);
xnor U18005 (N_18005,N_17395,N_16198);
xor U18006 (N_18006,N_16400,N_16454);
nor U18007 (N_18007,N_16638,N_16941);
nand U18008 (N_18008,N_16410,N_15361);
xnor U18009 (N_18009,N_16808,N_16130);
xor U18010 (N_18010,N_17275,N_15441);
and U18011 (N_18011,N_15965,N_16194);
nor U18012 (N_18012,N_16473,N_16103);
or U18013 (N_18013,N_16933,N_15433);
and U18014 (N_18014,N_15554,N_15830);
nor U18015 (N_18015,N_15161,N_15734);
or U18016 (N_18016,N_15197,N_17191);
nor U18017 (N_18017,N_15587,N_15470);
and U18018 (N_18018,N_15960,N_16109);
and U18019 (N_18019,N_16749,N_15752);
nor U18020 (N_18020,N_17010,N_15295);
or U18021 (N_18021,N_17495,N_16572);
nor U18022 (N_18022,N_17473,N_15037);
nor U18023 (N_18023,N_17251,N_16554);
and U18024 (N_18024,N_15067,N_16804);
nor U18025 (N_18025,N_17416,N_16397);
nand U18026 (N_18026,N_16244,N_16260);
nor U18027 (N_18027,N_17062,N_16300);
and U18028 (N_18028,N_17482,N_15861);
or U18029 (N_18029,N_15810,N_17456);
xnor U18030 (N_18030,N_15842,N_16989);
nand U18031 (N_18031,N_16543,N_17000);
nor U18032 (N_18032,N_15506,N_17232);
nor U18033 (N_18033,N_15323,N_16874);
or U18034 (N_18034,N_16881,N_15449);
nor U18035 (N_18035,N_15327,N_17276);
or U18036 (N_18036,N_16879,N_15612);
nand U18037 (N_18037,N_16072,N_17117);
xor U18038 (N_18038,N_15970,N_15906);
xor U18039 (N_18039,N_15643,N_16357);
or U18040 (N_18040,N_15386,N_17126);
nor U18041 (N_18041,N_15520,N_16775);
nor U18042 (N_18042,N_16901,N_17092);
nand U18043 (N_18043,N_16533,N_16582);
nor U18044 (N_18044,N_16100,N_16373);
nor U18045 (N_18045,N_15040,N_15027);
and U18046 (N_18046,N_15768,N_15593);
or U18047 (N_18047,N_16337,N_16237);
xor U18048 (N_18048,N_15533,N_17304);
and U18049 (N_18049,N_15581,N_17487);
nor U18050 (N_18050,N_15124,N_15964);
or U18051 (N_18051,N_15435,N_17302);
nor U18052 (N_18052,N_15096,N_16309);
nor U18053 (N_18053,N_16601,N_17271);
nand U18054 (N_18054,N_16875,N_15239);
nand U18055 (N_18055,N_15414,N_16574);
nand U18056 (N_18056,N_17210,N_16456);
or U18057 (N_18057,N_16350,N_16669);
and U18058 (N_18058,N_17351,N_15334);
xor U18059 (N_18059,N_16246,N_15879);
xnor U18060 (N_18060,N_15362,N_15799);
or U18061 (N_18061,N_16430,N_16243);
or U18062 (N_18062,N_16245,N_16478);
nor U18063 (N_18063,N_16858,N_15860);
xnor U18064 (N_18064,N_15050,N_16317);
nor U18065 (N_18065,N_16905,N_16391);
xnor U18066 (N_18066,N_15838,N_17039);
nor U18067 (N_18067,N_16882,N_16964);
xnor U18068 (N_18068,N_15464,N_15775);
or U18069 (N_18069,N_16703,N_15740);
and U18070 (N_18070,N_16909,N_15796);
or U18071 (N_18071,N_15863,N_15477);
nor U18072 (N_18072,N_15380,N_16322);
nand U18073 (N_18073,N_17076,N_15792);
nor U18074 (N_18074,N_15290,N_17313);
and U18075 (N_18075,N_16126,N_15911);
xor U18076 (N_18076,N_17004,N_17427);
nand U18077 (N_18077,N_16200,N_15869);
and U18078 (N_18078,N_15549,N_17466);
nor U18079 (N_18079,N_15984,N_16348);
xnor U18080 (N_18080,N_15452,N_16402);
and U18081 (N_18081,N_16690,N_15364);
nor U18082 (N_18082,N_16038,N_15370);
nand U18083 (N_18083,N_16795,N_15666);
and U18084 (N_18084,N_17447,N_15795);
xnor U18085 (N_18085,N_16555,N_16850);
xnor U18086 (N_18086,N_15665,N_15070);
xnor U18087 (N_18087,N_15405,N_15007);
or U18088 (N_18088,N_15925,N_15432);
xnor U18089 (N_18089,N_15206,N_16701);
nand U18090 (N_18090,N_15148,N_15820);
and U18091 (N_18091,N_17181,N_15988);
nand U18092 (N_18092,N_17289,N_15000);
and U18093 (N_18093,N_16668,N_16631);
xor U18094 (N_18094,N_16918,N_16959);
nand U18095 (N_18095,N_15350,N_17360);
nand U18096 (N_18096,N_16231,N_16316);
xor U18097 (N_18097,N_16170,N_16031);
or U18098 (N_18098,N_17121,N_16476);
or U18099 (N_18099,N_17429,N_15471);
nor U18100 (N_18100,N_16233,N_15193);
or U18101 (N_18101,N_15229,N_17222);
and U18102 (N_18102,N_15613,N_15677);
or U18103 (N_18103,N_16303,N_16010);
and U18104 (N_18104,N_17297,N_16257);
or U18105 (N_18105,N_16825,N_15410);
nand U18106 (N_18106,N_15944,N_16563);
or U18107 (N_18107,N_16140,N_15212);
xor U18108 (N_18108,N_16630,N_15039);
nor U18109 (N_18109,N_16351,N_15300);
and U18110 (N_18110,N_17160,N_17280);
and U18111 (N_18111,N_15065,N_15932);
nand U18112 (N_18112,N_16813,N_16663);
or U18113 (N_18113,N_15722,N_15314);
nor U18114 (N_18114,N_17486,N_15383);
xor U18115 (N_18115,N_16678,N_15267);
nand U18116 (N_18116,N_15002,N_15154);
or U18117 (N_18117,N_16277,N_15947);
or U18118 (N_18118,N_15171,N_15330);
nor U18119 (N_18119,N_15130,N_15876);
xnor U18120 (N_18120,N_16684,N_16510);
or U18121 (N_18121,N_16332,N_16382);
and U18122 (N_18122,N_16292,N_15808);
xnor U18123 (N_18123,N_16342,N_15072);
xor U18124 (N_18124,N_15322,N_17240);
or U18125 (N_18125,N_17068,N_16955);
and U18126 (N_18126,N_15354,N_16724);
xnor U18127 (N_18127,N_16472,N_16626);
nand U18128 (N_18128,N_17467,N_16041);
nor U18129 (N_18129,N_16163,N_15891);
nand U18130 (N_18130,N_16594,N_16893);
nand U18131 (N_18131,N_16376,N_17007);
xnor U18132 (N_18132,N_15234,N_16436);
xor U18133 (N_18133,N_17176,N_15657);
nor U18134 (N_18134,N_16516,N_15714);
xnor U18135 (N_18135,N_15183,N_16934);
and U18136 (N_18136,N_17424,N_16746);
nor U18137 (N_18137,N_16883,N_15230);
nor U18138 (N_18138,N_17361,N_17371);
xor U18139 (N_18139,N_16377,N_16161);
xor U18140 (N_18140,N_16782,N_16221);
xor U18141 (N_18141,N_15951,N_16602);
xnor U18142 (N_18142,N_16611,N_15684);
and U18143 (N_18143,N_16911,N_17124);
nand U18144 (N_18144,N_15041,N_15950);
nand U18145 (N_18145,N_15401,N_16694);
and U18146 (N_18146,N_17407,N_17479);
nor U18147 (N_18147,N_16298,N_17393);
or U18148 (N_18148,N_16800,N_15772);
nand U18149 (N_18149,N_16012,N_17493);
or U18150 (N_18150,N_17383,N_17132);
and U18151 (N_18151,N_17478,N_17430);
nor U18152 (N_18152,N_15802,N_17088);
xor U18153 (N_18153,N_16617,N_16033);
or U18154 (N_18154,N_16928,N_16297);
nor U18155 (N_18155,N_16649,N_15168);
nor U18156 (N_18156,N_16805,N_16270);
nor U18157 (N_18157,N_15928,N_15881);
or U18158 (N_18158,N_15680,N_15382);
or U18159 (N_18159,N_16803,N_15913);
nor U18160 (N_18160,N_15138,N_17161);
nand U18161 (N_18161,N_15393,N_16791);
or U18162 (N_18162,N_16479,N_16750);
xnor U18163 (N_18163,N_15560,N_17433);
and U18164 (N_18164,N_16060,N_16271);
xor U18165 (N_18165,N_16294,N_17301);
nand U18166 (N_18166,N_15738,N_17332);
and U18167 (N_18167,N_16977,N_16773);
or U18168 (N_18168,N_16059,N_17175);
xnor U18169 (N_18169,N_15092,N_16035);
xnor U18170 (N_18170,N_15289,N_17471);
nor U18171 (N_18171,N_15877,N_16788);
or U18172 (N_18172,N_15909,N_16500);
or U18173 (N_18173,N_17404,N_16575);
xnor U18174 (N_18174,N_16992,N_15851);
xnor U18175 (N_18175,N_15969,N_15638);
nor U18176 (N_18176,N_17028,N_16865);
or U18177 (N_18177,N_17188,N_17066);
or U18178 (N_18178,N_16973,N_16485);
nor U18179 (N_18179,N_15621,N_17391);
xnor U18180 (N_18180,N_17243,N_15998);
and U18181 (N_18181,N_16343,N_15258);
nand U18182 (N_18182,N_17485,N_17242);
nand U18183 (N_18183,N_17458,N_16877);
or U18184 (N_18184,N_16531,N_16546);
nand U18185 (N_18185,N_16084,N_15597);
nor U18186 (N_18186,N_16112,N_15543);
xor U18187 (N_18187,N_16903,N_15346);
xnor U18188 (N_18188,N_15573,N_16057);
or U18189 (N_18189,N_17263,N_15646);
and U18190 (N_18190,N_15592,N_16051);
nor U18191 (N_18191,N_16627,N_16178);
xor U18192 (N_18192,N_15528,N_15274);
nor U18193 (N_18193,N_15149,N_16709);
or U18194 (N_18194,N_15459,N_17089);
xnor U18195 (N_18195,N_16369,N_17202);
nor U18196 (N_18196,N_16947,N_16290);
xnor U18197 (N_18197,N_17338,N_15218);
and U18198 (N_18198,N_15277,N_15381);
and U18199 (N_18199,N_16591,N_15537);
nor U18200 (N_18200,N_17144,N_15412);
or U18201 (N_18201,N_16590,N_15652);
nand U18202 (N_18202,N_16643,N_15751);
and U18203 (N_18203,N_15938,N_17091);
and U18204 (N_18204,N_15803,N_15481);
nor U18205 (N_18205,N_15634,N_16050);
and U18206 (N_18206,N_16445,N_17164);
xor U18207 (N_18207,N_17125,N_16508);
and U18208 (N_18208,N_16054,N_16943);
xor U18209 (N_18209,N_16514,N_16584);
xnor U18210 (N_18210,N_17103,N_15993);
or U18211 (N_18211,N_15503,N_17201);
nor U18212 (N_18212,N_16836,N_15568);
nand U18213 (N_18213,N_15089,N_16980);
and U18214 (N_18214,N_16000,N_15016);
nor U18215 (N_18215,N_17077,N_16723);
or U18216 (N_18216,N_17084,N_15559);
and U18217 (N_18217,N_16922,N_17448);
xor U18218 (N_18218,N_15977,N_17307);
xnor U18219 (N_18219,N_15353,N_16747);
xnor U18220 (N_18220,N_16899,N_15097);
nor U18221 (N_18221,N_16592,N_17403);
xor U18222 (N_18222,N_16468,N_16073);
xor U18223 (N_18223,N_15326,N_15194);
or U18224 (N_18224,N_15958,N_16576);
xor U18225 (N_18225,N_17013,N_17266);
nor U18226 (N_18226,N_15748,N_15910);
xnor U18227 (N_18227,N_17292,N_15011);
or U18228 (N_18228,N_16385,N_16338);
nor U18229 (N_18229,N_17246,N_16824);
or U18230 (N_18230,N_15939,N_16867);
xnor U18231 (N_18231,N_16249,N_15787);
nor U18232 (N_18232,N_15182,N_17369);
or U18233 (N_18233,N_15404,N_16098);
xor U18234 (N_18234,N_15276,N_16998);
xnor U18235 (N_18235,N_16210,N_16622);
nand U18236 (N_18236,N_16239,N_15156);
xor U18237 (N_18237,N_16532,N_15524);
and U18238 (N_18238,N_17223,N_16215);
xnor U18239 (N_18239,N_15764,N_17141);
xnor U18240 (N_18240,N_16990,N_16693);
nand U18241 (N_18241,N_15090,N_16513);
and U18242 (N_18242,N_15365,N_17362);
nand U18243 (N_18243,N_15606,N_15611);
xor U18244 (N_18244,N_16986,N_15954);
nor U18245 (N_18245,N_17273,N_16295);
xnor U18246 (N_18246,N_16068,N_15115);
nor U18247 (N_18247,N_16623,N_15585);
or U18248 (N_18248,N_16640,N_16347);
nor U18249 (N_18249,N_15615,N_15083);
or U18250 (N_18250,N_17299,N_15605);
nor U18251 (N_18251,N_16981,N_15485);
xor U18252 (N_18252,N_17337,N_15674);
nor U18253 (N_18253,N_16715,N_16167);
xor U18254 (N_18254,N_15961,N_17374);
nor U18255 (N_18255,N_15057,N_15756);
and U18256 (N_18256,N_16034,N_15971);
or U18257 (N_18257,N_17016,N_15824);
or U18258 (N_18258,N_17213,N_15636);
xor U18259 (N_18259,N_15428,N_15651);
and U18260 (N_18260,N_16614,N_15599);
nor U18261 (N_18261,N_17431,N_16728);
nand U18262 (N_18262,N_15713,N_16772);
xor U18263 (N_18263,N_16762,N_17425);
or U18264 (N_18264,N_15933,N_15397);
xnor U18265 (N_18265,N_16760,N_16958);
or U18266 (N_18266,N_15858,N_16757);
nand U18267 (N_18267,N_15221,N_15747);
and U18268 (N_18268,N_16869,N_15571);
xnor U18269 (N_18269,N_17492,N_17293);
nor U18270 (N_18270,N_17469,N_15379);
and U18271 (N_18271,N_15510,N_17035);
xnor U18272 (N_18272,N_15169,N_16783);
and U18273 (N_18273,N_17226,N_16719);
xor U18274 (N_18274,N_16224,N_15209);
nor U18275 (N_18275,N_15439,N_17237);
or U18276 (N_18276,N_16845,N_16790);
nand U18277 (N_18277,N_17060,N_15109);
or U18278 (N_18278,N_16183,N_17081);
and U18279 (N_18279,N_16557,N_15991);
and U18280 (N_18280,N_17476,N_17350);
nand U18281 (N_18281,N_17209,N_15511);
nor U18282 (N_18282,N_15215,N_16486);
xnor U18283 (N_18283,N_15930,N_16179);
xnor U18284 (N_18284,N_15884,N_16372);
or U18285 (N_18285,N_15753,N_16606);
xnor U18286 (N_18286,N_16079,N_15461);
or U18287 (N_18287,N_15935,N_17083);
xor U18288 (N_18288,N_16394,N_16652);
or U18289 (N_18289,N_16780,N_17364);
nor U18290 (N_18290,N_15042,N_16931);
xor U18291 (N_18291,N_17238,N_16318);
nand U18292 (N_18292,N_16185,N_17354);
nand U18293 (N_18293,N_16280,N_17484);
and U18294 (N_18294,N_15908,N_16101);
and U18295 (N_18295,N_15248,N_17477);
nor U18296 (N_18296,N_15693,N_15328);
and U18297 (N_18297,N_17022,N_16075);
nor U18298 (N_18298,N_15702,N_15823);
nand U18299 (N_18299,N_16689,N_15784);
or U18300 (N_18300,N_16211,N_16708);
nand U18301 (N_18301,N_15670,N_16733);
xnor U18302 (N_18302,N_16389,N_16086);
nand U18303 (N_18303,N_16155,N_15990);
nor U18304 (N_18304,N_16506,N_15563);
xnor U18305 (N_18305,N_15681,N_16673);
or U18306 (N_18306,N_17440,N_17290);
xnor U18307 (N_18307,N_15916,N_16188);
nor U18308 (N_18308,N_15272,N_16686);
xnor U18309 (N_18309,N_16381,N_16477);
xnor U18310 (N_18310,N_16784,N_17041);
nand U18311 (N_18311,N_17111,N_15084);
xnor U18312 (N_18312,N_17426,N_15318);
nor U18313 (N_18313,N_17311,N_15051);
nor U18314 (N_18314,N_16856,N_17432);
or U18315 (N_18315,N_17316,N_16061);
or U18316 (N_18316,N_16129,N_15345);
nand U18317 (N_18317,N_17208,N_15766);
nand U18318 (N_18318,N_16063,N_17341);
xnor U18319 (N_18319,N_17134,N_16657);
nor U18320 (N_18320,N_15922,N_15122);
nand U18321 (N_18321,N_15773,N_15224);
nor U18322 (N_18322,N_17499,N_16857);
nand U18323 (N_18323,N_15055,N_16849);
nand U18324 (N_18324,N_16566,N_16636);
and U18325 (N_18325,N_16498,N_16884);
or U18326 (N_18326,N_17260,N_15204);
or U18327 (N_18327,N_17438,N_16637);
nor U18328 (N_18328,N_15358,N_16936);
and U18329 (N_18329,N_15143,N_16608);
and U18330 (N_18330,N_15594,N_15626);
nor U18331 (N_18331,N_16141,N_15377);
and U18332 (N_18332,N_15247,N_16006);
nor U18333 (N_18333,N_16991,N_15819);
or U18334 (N_18334,N_15574,N_17385);
xor U18335 (N_18335,N_17097,N_15540);
or U18336 (N_18336,N_17356,N_15531);
nor U18337 (N_18337,N_15582,N_16358);
xor U18338 (N_18338,N_16885,N_15493);
nand U18339 (N_18339,N_15257,N_17392);
and U18340 (N_18340,N_16254,N_17036);
or U18341 (N_18341,N_16573,N_17199);
xor U18342 (N_18342,N_16954,N_15866);
xor U18343 (N_18343,N_15400,N_16696);
and U18344 (N_18344,N_16053,N_16027);
nor U18345 (N_18345,N_16320,N_17079);
or U18346 (N_18346,N_16700,N_15241);
xnor U18347 (N_18347,N_15695,N_17272);
nor U18348 (N_18348,N_16567,N_16827);
and U18349 (N_18349,N_16276,N_16639);
xnor U18350 (N_18350,N_15767,N_17149);
xnor U18351 (N_18351,N_16461,N_15491);
nor U18352 (N_18352,N_16064,N_15298);
or U18353 (N_18353,N_15529,N_17015);
nand U18354 (N_18354,N_16515,N_17047);
nor U18355 (N_18355,N_15828,N_17233);
xnor U18356 (N_18356,N_16967,N_15203);
nand U18357 (N_18357,N_15901,N_15967);
or U18358 (N_18358,N_15723,N_15862);
and U18359 (N_18359,N_16181,N_16561);
xor U18360 (N_18360,N_17366,N_15974);
xnor U18361 (N_18361,N_15214,N_16096);
and U18362 (N_18362,N_15142,N_16455);
or U18363 (N_18363,N_16045,N_16177);
or U18364 (N_18364,N_16013,N_16957);
nor U18365 (N_18365,N_15545,N_15595);
nand U18366 (N_18366,N_15683,N_16262);
nor U18367 (N_18367,N_16926,N_17497);
xor U18368 (N_18368,N_16917,N_15222);
and U18369 (N_18369,N_15281,N_15589);
nor U18370 (N_18370,N_15857,N_16944);
or U18371 (N_18371,N_15201,N_16568);
nand U18372 (N_18372,N_16530,N_15164);
or U18373 (N_18373,N_15253,N_17312);
or U18374 (N_18374,N_16118,N_16440);
and U18375 (N_18375,N_15059,N_16697);
and U18376 (N_18376,N_15848,N_17451);
and U18377 (N_18377,N_15210,N_16996);
nor U18378 (N_18378,N_16032,N_15246);
nor U18379 (N_18379,N_16308,N_15790);
and U18380 (N_18380,N_16288,N_17157);
nand U18381 (N_18381,N_16366,N_16818);
nand U18382 (N_18382,N_17102,N_15567);
nor U18383 (N_18383,N_15136,N_15895);
nand U18384 (N_18384,N_16570,N_17185);
or U18385 (N_18385,N_17067,N_17375);
nand U18386 (N_18386,N_15463,N_17446);
nor U18387 (N_18387,N_15687,N_15924);
or U18388 (N_18388,N_16387,N_15268);
xnor U18389 (N_18389,N_16175,N_17435);
or U18390 (N_18390,N_15170,N_16585);
xor U18391 (N_18391,N_16716,N_16578);
nand U18392 (N_18392,N_17241,N_17150);
nor U18393 (N_18393,N_16927,N_17309);
nand U18394 (N_18394,N_15063,N_17344);
nand U18395 (N_18395,N_15614,N_16487);
nand U18396 (N_18396,N_15093,N_15672);
or U18397 (N_18397,N_16093,N_15325);
xor U18398 (N_18398,N_17074,N_16727);
nor U18399 (N_18399,N_15173,N_16737);
xnor U18400 (N_18400,N_15811,N_16169);
nand U18401 (N_18401,N_15814,N_16710);
nor U18402 (N_18402,N_16404,N_16916);
nor U18403 (N_18403,N_17255,N_15618);
nand U18404 (N_18404,N_16739,N_17330);
and U18405 (N_18405,N_16085,N_16987);
xnor U18406 (N_18406,N_15031,N_16660);
nor U18407 (N_18407,N_17008,N_15012);
or U18408 (N_18408,N_16124,N_15468);
or U18409 (N_18409,N_16405,N_15375);
xnor U18410 (N_18410,N_16726,N_16528);
nor U18411 (N_18411,N_16886,N_15675);
and U18412 (N_18412,N_15347,N_17058);
xnor U18413 (N_18413,N_17224,N_16230);
xor U18414 (N_18414,N_15066,N_16699);
or U18415 (N_18415,N_17228,N_15240);
nand U18416 (N_18416,N_15301,N_15726);
nor U18417 (N_18417,N_15269,N_16796);
xor U18418 (N_18418,N_15957,N_15628);
and U18419 (N_18419,N_15591,N_16242);
and U18420 (N_18420,N_16192,N_16665);
nor U18421 (N_18421,N_15989,N_17109);
nand U18422 (N_18422,N_17472,N_17115);
xor U18423 (N_18423,N_17317,N_16851);
and U18424 (N_18424,N_16540,N_17402);
nor U18425 (N_18425,N_15455,N_15207);
xnor U18426 (N_18426,N_16058,N_16966);
and U18427 (N_18427,N_15145,N_15690);
or U18428 (N_18428,N_15043,N_17349);
nor U18429 (N_18429,N_15213,N_16677);
nor U18430 (N_18430,N_17342,N_16529);
and U18431 (N_18431,N_15780,N_15996);
and U18432 (N_18432,N_15378,N_15880);
nand U18433 (N_18433,N_15656,N_16428);
and U18434 (N_18434,N_16717,N_16659);
or U18435 (N_18435,N_17400,N_15476);
or U18436 (N_18436,N_17239,N_17107);
or U18437 (N_18437,N_16452,N_17053);
xor U18438 (N_18438,N_15496,N_15304);
or U18439 (N_18439,N_15111,N_17189);
xor U18440 (N_18440,N_15564,N_16888);
and U18441 (N_18441,N_16115,N_16283);
nor U18442 (N_18442,N_15649,N_16834);
xor U18443 (N_18443,N_16938,N_15761);
xor U18444 (N_18444,N_17248,N_15541);
or U18445 (N_18445,N_16326,N_16354);
nand U18446 (N_18446,N_16160,N_17294);
or U18447 (N_18447,N_16307,N_15717);
or U18448 (N_18448,N_17318,N_16618);
nor U18449 (N_18449,N_16040,N_17264);
nand U18450 (N_18450,N_16113,N_17211);
and U18451 (N_18451,N_15306,N_15010);
nand U18452 (N_18452,N_15457,N_16889);
or U18453 (N_18453,N_17379,N_15292);
nand U18454 (N_18454,N_17343,N_16441);
nor U18455 (N_18455,N_16489,N_17085);
nor U18456 (N_18456,N_17331,N_17418);
xor U18457 (N_18457,N_17148,N_16718);
and U18458 (N_18458,N_16312,N_17428);
nor U18459 (N_18459,N_15366,N_16451);
or U18460 (N_18460,N_16148,N_16846);
xor U18461 (N_18461,N_15625,N_16906);
xnor U18462 (N_18462,N_16284,N_15912);
or U18463 (N_18463,N_16713,N_16655);
or U18464 (N_18464,N_16008,N_16186);
or U18465 (N_18465,N_15284,N_16920);
or U18466 (N_18466,N_16672,N_15237);
nand U18467 (N_18467,N_16548,N_16603);
and U18468 (N_18468,N_17108,N_17096);
and U18469 (N_18469,N_16595,N_16781);
xnor U18470 (N_18470,N_16551,N_15408);
and U18471 (N_18471,N_15273,N_15153);
or U18472 (N_18472,N_15550,N_16104);
and U18473 (N_18473,N_16080,N_17152);
or U18474 (N_18474,N_16241,N_15280);
xnor U18475 (N_18475,N_16196,N_16019);
or U18476 (N_18476,N_16043,N_16634);
and U18477 (N_18477,N_15539,N_16738);
nor U18478 (N_18478,N_16544,N_15311);
and U18479 (N_18479,N_17219,N_16621);
nand U18480 (N_18480,N_15118,N_17468);
xor U18481 (N_18481,N_16847,N_15337);
nand U18482 (N_18482,N_15653,N_16722);
nand U18483 (N_18483,N_16432,N_16150);
and U18484 (N_18484,N_17324,N_16896);
and U18485 (N_18485,N_17443,N_15114);
nand U18486 (N_18486,N_15447,N_15673);
nand U18487 (N_18487,N_16613,N_16065);
and U18488 (N_18488,N_15849,N_15023);
and U18489 (N_18489,N_16217,N_16328);
nand U18490 (N_18490,N_16704,N_17457);
xnor U18491 (N_18491,N_15105,N_16953);
nand U18492 (N_18492,N_16460,N_15339);
and U18493 (N_18493,N_16810,N_15536);
or U18494 (N_18494,N_16070,N_16488);
nand U18495 (N_18495,N_15077,N_15252);
xnor U18496 (N_18496,N_15359,N_16355);
nand U18497 (N_18497,N_16736,N_15663);
or U18498 (N_18498,N_16427,N_16482);
and U18499 (N_18499,N_16265,N_16526);
and U18500 (N_18500,N_15296,N_16156);
nor U18501 (N_18501,N_15608,N_17284);
xor U18502 (N_18502,N_17040,N_16598);
or U18503 (N_18503,N_17129,N_16785);
or U18504 (N_18504,N_15054,N_16612);
nor U18505 (N_18505,N_15438,N_16123);
nand U18506 (N_18506,N_16089,N_17415);
xor U18507 (N_18507,N_17449,N_16863);
nand U18508 (N_18508,N_16368,N_16248);
xor U18509 (N_18509,N_16028,N_17340);
or U18510 (N_18510,N_16088,N_16119);
nand U18511 (N_18511,N_16907,N_15956);
nand U18512 (N_18512,N_16339,N_16157);
nor U18513 (N_18513,N_16269,N_15896);
or U18514 (N_18514,N_16688,N_15865);
nor U18515 (N_18515,N_16021,N_16910);
xor U18516 (N_18516,N_15873,N_16213);
xnor U18517 (N_18517,N_17186,N_15071);
nor U18518 (N_18518,N_15953,N_16029);
or U18519 (N_18519,N_16131,N_15019);
nor U18520 (N_18520,N_16666,N_16852);
xnor U18521 (N_18521,N_15718,N_15980);
and U18522 (N_18522,N_15087,N_16679);
or U18523 (N_18523,N_15716,N_15514);
nand U18524 (N_18524,N_16793,N_15264);
nor U18525 (N_18525,N_17368,N_16007);
and U18526 (N_18526,N_16952,N_15338);
nand U18527 (N_18527,N_17100,N_15113);
xnor U18528 (N_18528,N_15028,N_15871);
xor U18529 (N_18529,N_15578,N_16951);
or U18530 (N_18530,N_15968,N_17412);
xnor U18531 (N_18531,N_15749,N_15882);
xor U18532 (N_18532,N_15402,N_16448);
and U18533 (N_18533,N_16380,N_16682);
xnor U18534 (N_18534,N_16289,N_16097);
and U18535 (N_18535,N_16147,N_17420);
or U18536 (N_18536,N_15080,N_17491);
nor U18537 (N_18537,N_15088,N_15553);
xnor U18538 (N_18538,N_15655,N_15429);
nand U18539 (N_18539,N_15064,N_16094);
nor U18540 (N_18540,N_16721,N_17397);
nor U18541 (N_18541,N_16769,N_16577);
nor U18542 (N_18542,N_15619,N_15184);
and U18543 (N_18543,N_17434,N_15500);
and U18544 (N_18544,N_17333,N_17105);
xnor U18545 (N_18545,N_15391,N_16897);
nor U18546 (N_18546,N_15003,N_16787);
nor U18547 (N_18547,N_17018,N_15759);
nand U18548 (N_18548,N_15786,N_15515);
or U18549 (N_18549,N_17442,N_15162);
xor U18550 (N_18550,N_15758,N_16830);
nor U18551 (N_18551,N_15225,N_17093);
and U18552 (N_18552,N_15697,N_15502);
xor U18553 (N_18553,N_17475,N_15532);
xnor U18554 (N_18554,N_15035,N_16026);
and U18555 (N_18555,N_15018,N_15846);
and U18556 (N_18556,N_16822,N_15117);
and U18557 (N_18557,N_16523,N_15566);
and U18558 (N_18558,N_16985,N_15855);
nand U18559 (N_18559,N_15598,N_15372);
and U18560 (N_18560,N_17151,N_15501);
and U18561 (N_18561,N_15341,N_15504);
nand U18562 (N_18562,N_16286,N_15781);
and U18563 (N_18563,N_17254,N_16361);
nand U18564 (N_18564,N_15116,N_16892);
nand U18565 (N_18565,N_15094,N_15942);
nor U18566 (N_18566,N_17137,N_16662);
and U18567 (N_18567,N_16855,N_15671);
xor U18568 (N_18568,N_15959,N_15729);
nand U18569 (N_18569,N_15437,N_15743);
and U18570 (N_18570,N_17171,N_16720);
nand U18571 (N_18571,N_15973,N_15955);
and U18572 (N_18572,N_16741,N_17215);
xor U18573 (N_18573,N_16273,N_16341);
or U18574 (N_18574,N_17489,N_17279);
nand U18575 (N_18575,N_17394,N_17306);
or U18576 (N_18576,N_17080,N_16090);
xnor U18577 (N_18577,N_17044,N_15508);
and U18578 (N_18578,N_16921,N_17163);
nand U18579 (N_18579,N_17177,N_15905);
and U18580 (N_18580,N_16470,N_16974);
or U18581 (N_18581,N_16774,N_17136);
xor U18582 (N_18582,N_16635,N_16466);
xor U18583 (N_18583,N_16403,N_16820);
nor U18584 (N_18584,N_15321,N_16172);
nor U18585 (N_18585,N_16588,N_17087);
and U18586 (N_18586,N_16143,N_15696);
nor U18587 (N_18587,N_15839,N_15029);
and U18588 (N_18588,N_16433,N_17095);
or U18589 (N_18589,N_15188,N_17413);
nor U18590 (N_18590,N_16891,N_16356);
xor U18591 (N_18591,N_15110,N_15899);
nand U18592 (N_18592,N_16794,N_15312);
or U18593 (N_18593,N_16538,N_16491);
xor U18594 (N_18594,N_16407,N_16017);
nor U18595 (N_18595,N_16778,N_17221);
and U18596 (N_18596,N_16814,N_15620);
nor U18597 (N_18597,N_15052,N_15440);
nor U18598 (N_18598,N_15396,N_15546);
nor U18599 (N_18599,N_16149,N_16676);
nor U18600 (N_18600,N_15963,N_17042);
and U18601 (N_18601,N_16121,N_16565);
or U18602 (N_18602,N_15091,N_15489);
nand U18603 (N_18603,N_16732,N_15557);
nand U18604 (N_18604,N_15623,N_15829);
xnor U18605 (N_18605,N_16553,N_16203);
nor U18606 (N_18606,N_17182,N_16039);
xor U18607 (N_18607,N_15238,N_15733);
nand U18608 (N_18608,N_15641,N_15985);
and U18609 (N_18609,N_16866,N_17381);
nand U18610 (N_18610,N_16024,N_15108);
and U18611 (N_18611,N_15867,N_16344);
or U18612 (N_18612,N_15516,N_17050);
xor U18613 (N_18613,N_17235,N_15106);
and U18614 (N_18614,N_16106,N_15174);
or U18615 (N_18615,N_15509,N_16583);
xnor U18616 (N_18616,N_16651,N_17230);
and U18617 (N_18617,N_16667,N_15995);
and U18618 (N_18618,N_16755,N_15588);
xnor U18619 (N_18619,N_15627,N_16442);
and U18620 (N_18620,N_17200,N_16549);
nand U18621 (N_18621,N_15217,N_15074);
nor U18622 (N_18622,N_16395,N_17061);
xnor U18623 (N_18623,N_16216,N_17387);
nor U18624 (N_18624,N_15765,N_16011);
or U18625 (N_18625,N_15648,N_15815);
nand U18626 (N_18626,N_15180,N_17250);
nand U18627 (N_18627,N_16151,N_15818);
and U18628 (N_18628,N_17212,N_16777);
nor U18629 (N_18629,N_17086,N_15903);
and U18630 (N_18630,N_16683,N_16250);
and U18631 (N_18631,N_16859,N_15711);
xnor U18632 (N_18632,N_15517,N_16056);
nor U18633 (N_18633,N_15797,N_16234);
and U18634 (N_18634,N_16937,N_16180);
nand U18635 (N_18635,N_17135,N_15157);
or U18636 (N_18636,N_16313,N_17295);
nand U18637 (N_18637,N_17048,N_15482);
and U18638 (N_18638,N_16604,N_17417);
or U18639 (N_18639,N_17075,N_16390);
nand U18640 (N_18640,N_15100,N_16706);
or U18641 (N_18641,N_15703,N_15152);
or U18642 (N_18642,N_17262,N_16226);
or U18643 (N_18643,N_15418,N_16371);
or U18644 (N_18644,N_15667,N_15806);
or U18645 (N_18645,N_15826,N_15885);
or U18646 (N_18646,N_15022,N_17377);
or U18647 (N_18647,N_15073,N_15538);
or U18648 (N_18648,N_16346,N_15724);
nor U18649 (N_18649,N_16268,N_17247);
xor U18650 (N_18650,N_15079,N_17159);
xor U18651 (N_18651,N_16153,N_17169);
and U18652 (N_18652,N_17372,N_16819);
or U18653 (N_18653,N_17268,N_17336);
or U18654 (N_18654,N_17214,N_16398);
nand U18655 (N_18655,N_16435,N_16890);
nand U18656 (N_18656,N_17245,N_15730);
nand U18657 (N_18657,N_15548,N_16329);
nand U18658 (N_18658,N_15125,N_15310);
xnor U18659 (N_18659,N_15847,N_16083);
and U18660 (N_18660,N_16437,N_16754);
nor U18661 (N_18661,N_17346,N_16817);
nand U18662 (N_18662,N_15807,N_17057);
nor U18663 (N_18663,N_16420,N_16282);
xnor U18664 (N_18664,N_16002,N_16110);
xor U18665 (N_18665,N_17225,N_15395);
and U18666 (N_18666,N_15981,N_17192);
or U18667 (N_18667,N_17423,N_16379);
nand U18668 (N_18668,N_16520,N_15763);
or U18669 (N_18669,N_15530,N_16363);
nor U18670 (N_18670,N_16374,N_16279);
xor U18671 (N_18671,N_15069,N_16579);
and U18672 (N_18672,N_16349,N_15475);
nor U18673 (N_18673,N_15466,N_15465);
xnor U18674 (N_18674,N_17078,N_17146);
and U18675 (N_18675,N_16743,N_16287);
nand U18676 (N_18676,N_17249,N_15617);
xor U18677 (N_18677,N_15731,N_15228);
nand U18678 (N_18678,N_17378,N_16902);
nand U18679 (N_18679,N_15219,N_15250);
xor U18680 (N_18680,N_15456,N_16542);
or U18681 (N_18681,N_16414,N_15389);
xnor U18682 (N_18682,N_17411,N_15495);
and U18683 (N_18683,N_15172,N_16335);
nor U18684 (N_18684,N_16107,N_16232);
xor U18685 (N_18685,N_17153,N_16771);
and U18686 (N_18686,N_15735,N_17315);
xor U18687 (N_18687,N_15260,N_15875);
nand U18688 (N_18688,N_15303,N_17049);
and U18689 (N_18689,N_15816,N_17065);
nand U18690 (N_18690,N_16752,N_15522);
xnor U18691 (N_18691,N_16946,N_17388);
nor U18692 (N_18692,N_17283,N_16071);
and U18693 (N_18693,N_15742,N_16811);
xnor U18694 (N_18694,N_15360,N_15451);
and U18695 (N_18695,N_17422,N_16535);
and U18696 (N_18696,N_17099,N_16873);
nand U18697 (N_18697,N_15853,N_16345);
xor U18698 (N_18698,N_15505,N_15610);
and U18699 (N_18699,N_16517,N_15691);
xor U18700 (N_18700,N_16296,N_15556);
or U18701 (N_18701,N_17419,N_17064);
and U18702 (N_18702,N_16117,N_16569);
nor U18703 (N_18703,N_15948,N_17106);
and U18704 (N_18704,N_15727,N_16092);
xor U18705 (N_18705,N_15484,N_15650);
nor U18706 (N_18706,N_16912,N_17207);
and U18707 (N_18707,N_15409,N_17025);
or U18708 (N_18708,N_15822,N_16823);
or U18709 (N_18709,N_15254,N_17156);
nand U18710 (N_18710,N_16128,N_15841);
xnor U18711 (N_18711,N_17104,N_15190);
and U18712 (N_18712,N_16767,N_16458);
or U18713 (N_18713,N_17365,N_15783);
or U18714 (N_18714,N_15929,N_17439);
or U18715 (N_18715,N_15907,N_15739);
or U18716 (N_18716,N_17287,N_16171);
and U18717 (N_18717,N_16378,N_16256);
xnor U18718 (N_18718,N_15367,N_16336);
and U18719 (N_18719,N_15976,N_17203);
nand U18720 (N_18720,N_15897,N_15962);
nor U18721 (N_18721,N_15030,N_17334);
and U18722 (N_18722,N_17265,N_17029);
and U18723 (N_18723,N_16359,N_15936);
xnor U18724 (N_18724,N_16519,N_15812);
or U18725 (N_18725,N_16422,N_16504);
nand U18726 (N_18726,N_15099,N_16597);
nor U18727 (N_18727,N_15535,N_16969);
nor U18728 (N_18728,N_17382,N_15243);
xor U18729 (N_18729,N_15728,N_15700);
and U18730 (N_18730,N_15512,N_16018);
nand U18731 (N_18731,N_16490,N_15715);
xnor U18732 (N_18732,N_15890,N_16664);
xnor U18733 (N_18733,N_15662,N_15294);
xor U18734 (N_18734,N_16624,N_16464);
nand U18735 (N_18735,N_17033,N_15133);
nor U18736 (N_18736,N_15205,N_16236);
or U18737 (N_18737,N_17380,N_15415);
or U18738 (N_18738,N_17127,N_16605);
nor U18739 (N_18739,N_17496,N_15101);
or U18740 (N_18740,N_15979,N_15845);
nand U18741 (N_18741,N_15769,N_17194);
and U18742 (N_18742,N_16960,N_17190);
or U18743 (N_18743,N_15931,N_15352);
nor U18744 (N_18744,N_15844,N_17038);
nor U18745 (N_18745,N_15918,N_17119);
or U18746 (N_18746,N_16191,N_17314);
xnor U18747 (N_18747,N_15102,N_15137);
nor U18748 (N_18748,N_15624,N_16620);
and U18749 (N_18749,N_15843,N_15975);
xnor U18750 (N_18750,N_16097,N_16380);
xor U18751 (N_18751,N_16306,N_16816);
nor U18752 (N_18752,N_16354,N_16184);
nor U18753 (N_18753,N_16745,N_17047);
nand U18754 (N_18754,N_16598,N_16448);
and U18755 (N_18755,N_15175,N_16243);
nand U18756 (N_18756,N_17469,N_17154);
nand U18757 (N_18757,N_16912,N_16355);
xnor U18758 (N_18758,N_15447,N_16901);
and U18759 (N_18759,N_16041,N_15757);
nor U18760 (N_18760,N_16140,N_17045);
xor U18761 (N_18761,N_15719,N_15040);
nand U18762 (N_18762,N_15224,N_16618);
and U18763 (N_18763,N_16899,N_17273);
or U18764 (N_18764,N_16336,N_17127);
and U18765 (N_18765,N_15545,N_15238);
nand U18766 (N_18766,N_16391,N_15025);
and U18767 (N_18767,N_16409,N_16010);
nand U18768 (N_18768,N_17090,N_15645);
nor U18769 (N_18769,N_17317,N_16112);
nand U18770 (N_18770,N_16594,N_17215);
nor U18771 (N_18771,N_15964,N_16102);
nor U18772 (N_18772,N_16135,N_16056);
nor U18773 (N_18773,N_16859,N_16232);
nor U18774 (N_18774,N_17407,N_15087);
and U18775 (N_18775,N_16893,N_15681);
xor U18776 (N_18776,N_16896,N_17043);
xnor U18777 (N_18777,N_17237,N_15460);
or U18778 (N_18778,N_15886,N_15282);
nor U18779 (N_18779,N_16901,N_16424);
or U18780 (N_18780,N_15885,N_15782);
and U18781 (N_18781,N_15882,N_16409);
and U18782 (N_18782,N_16820,N_16121);
or U18783 (N_18783,N_15829,N_16652);
nor U18784 (N_18784,N_16921,N_17448);
nand U18785 (N_18785,N_15816,N_17478);
xor U18786 (N_18786,N_15619,N_16178);
or U18787 (N_18787,N_15446,N_16041);
or U18788 (N_18788,N_15352,N_16165);
and U18789 (N_18789,N_15982,N_17414);
nor U18790 (N_18790,N_16656,N_15966);
xnor U18791 (N_18791,N_16004,N_15522);
xor U18792 (N_18792,N_15533,N_16929);
or U18793 (N_18793,N_16821,N_16679);
and U18794 (N_18794,N_17080,N_16247);
xnor U18795 (N_18795,N_15865,N_15160);
nand U18796 (N_18796,N_16344,N_17192);
and U18797 (N_18797,N_16786,N_15720);
nand U18798 (N_18798,N_16902,N_15375);
nor U18799 (N_18799,N_15842,N_17209);
or U18800 (N_18800,N_17142,N_16651);
or U18801 (N_18801,N_16860,N_16465);
and U18802 (N_18802,N_15078,N_15180);
and U18803 (N_18803,N_16553,N_15794);
xor U18804 (N_18804,N_16704,N_15867);
and U18805 (N_18805,N_16532,N_15800);
or U18806 (N_18806,N_16266,N_15455);
nor U18807 (N_18807,N_15878,N_16785);
and U18808 (N_18808,N_16553,N_16159);
or U18809 (N_18809,N_16547,N_15957);
xor U18810 (N_18810,N_17240,N_17392);
nor U18811 (N_18811,N_16941,N_17118);
or U18812 (N_18812,N_15720,N_17315);
nand U18813 (N_18813,N_16452,N_16287);
xnor U18814 (N_18814,N_17380,N_16166);
or U18815 (N_18815,N_16868,N_16684);
or U18816 (N_18816,N_15305,N_15265);
nand U18817 (N_18817,N_16695,N_17411);
or U18818 (N_18818,N_16036,N_17086);
xor U18819 (N_18819,N_15579,N_16521);
xor U18820 (N_18820,N_15610,N_15237);
or U18821 (N_18821,N_16027,N_16770);
xor U18822 (N_18822,N_16831,N_17288);
nand U18823 (N_18823,N_17131,N_16942);
or U18824 (N_18824,N_15491,N_15621);
nor U18825 (N_18825,N_16477,N_17173);
nor U18826 (N_18826,N_15146,N_17083);
and U18827 (N_18827,N_15689,N_15261);
nor U18828 (N_18828,N_16139,N_17296);
nor U18829 (N_18829,N_15283,N_15943);
xor U18830 (N_18830,N_16548,N_16894);
nand U18831 (N_18831,N_15367,N_15820);
nor U18832 (N_18832,N_15837,N_15637);
or U18833 (N_18833,N_16206,N_16848);
nand U18834 (N_18834,N_16694,N_15585);
or U18835 (N_18835,N_17394,N_16049);
nand U18836 (N_18836,N_17325,N_15743);
and U18837 (N_18837,N_17050,N_16729);
or U18838 (N_18838,N_17042,N_15204);
xor U18839 (N_18839,N_17333,N_15886);
and U18840 (N_18840,N_15306,N_15831);
and U18841 (N_18841,N_15661,N_17044);
or U18842 (N_18842,N_15672,N_16473);
and U18843 (N_18843,N_16741,N_15370);
xnor U18844 (N_18844,N_16218,N_15814);
nor U18845 (N_18845,N_17099,N_15912);
nor U18846 (N_18846,N_16384,N_16327);
or U18847 (N_18847,N_16862,N_16543);
or U18848 (N_18848,N_17434,N_16950);
nor U18849 (N_18849,N_17335,N_16058);
nor U18850 (N_18850,N_15052,N_15282);
and U18851 (N_18851,N_17245,N_15455);
xor U18852 (N_18852,N_16771,N_17455);
and U18853 (N_18853,N_15715,N_15792);
and U18854 (N_18854,N_15610,N_16731);
nand U18855 (N_18855,N_16442,N_17393);
or U18856 (N_18856,N_17311,N_17086);
xor U18857 (N_18857,N_16092,N_15791);
or U18858 (N_18858,N_15862,N_15014);
nor U18859 (N_18859,N_17098,N_16291);
or U18860 (N_18860,N_16504,N_17353);
or U18861 (N_18861,N_15246,N_15227);
or U18862 (N_18862,N_15715,N_17330);
and U18863 (N_18863,N_16302,N_16376);
nor U18864 (N_18864,N_15387,N_16886);
and U18865 (N_18865,N_17162,N_15418);
xnor U18866 (N_18866,N_16609,N_16131);
xor U18867 (N_18867,N_15425,N_15857);
xnor U18868 (N_18868,N_16467,N_16171);
nor U18869 (N_18869,N_17408,N_15094);
nor U18870 (N_18870,N_17414,N_16552);
nor U18871 (N_18871,N_17026,N_15400);
and U18872 (N_18872,N_16154,N_15174);
and U18873 (N_18873,N_15057,N_16615);
nand U18874 (N_18874,N_17139,N_17446);
and U18875 (N_18875,N_15612,N_16446);
and U18876 (N_18876,N_17205,N_17140);
or U18877 (N_18877,N_16970,N_16845);
nand U18878 (N_18878,N_16582,N_15669);
and U18879 (N_18879,N_15575,N_15568);
and U18880 (N_18880,N_16041,N_15204);
or U18881 (N_18881,N_15846,N_16912);
nor U18882 (N_18882,N_17316,N_15952);
and U18883 (N_18883,N_15180,N_15293);
nand U18884 (N_18884,N_15105,N_16758);
nand U18885 (N_18885,N_15250,N_15357);
nor U18886 (N_18886,N_15256,N_16753);
xnor U18887 (N_18887,N_15524,N_15610);
nand U18888 (N_18888,N_15372,N_16647);
or U18889 (N_18889,N_16250,N_17171);
or U18890 (N_18890,N_16664,N_15147);
or U18891 (N_18891,N_16021,N_17213);
nand U18892 (N_18892,N_17293,N_15341);
or U18893 (N_18893,N_15075,N_15623);
nor U18894 (N_18894,N_16732,N_16837);
xor U18895 (N_18895,N_16355,N_15104);
nor U18896 (N_18896,N_17418,N_16334);
xor U18897 (N_18897,N_16857,N_15457);
or U18898 (N_18898,N_16105,N_15698);
nor U18899 (N_18899,N_15624,N_16173);
xnor U18900 (N_18900,N_17236,N_15791);
and U18901 (N_18901,N_16852,N_15947);
or U18902 (N_18902,N_17481,N_15132);
nand U18903 (N_18903,N_16714,N_17116);
nor U18904 (N_18904,N_16867,N_15637);
nand U18905 (N_18905,N_15154,N_17097);
nand U18906 (N_18906,N_16456,N_15868);
or U18907 (N_18907,N_15267,N_16203);
xor U18908 (N_18908,N_17188,N_17111);
xnor U18909 (N_18909,N_17024,N_17094);
and U18910 (N_18910,N_16802,N_15906);
or U18911 (N_18911,N_15542,N_15360);
nand U18912 (N_18912,N_17417,N_16059);
nand U18913 (N_18913,N_15810,N_16306);
nand U18914 (N_18914,N_15186,N_16875);
and U18915 (N_18915,N_17415,N_16755);
nand U18916 (N_18916,N_16916,N_16712);
xnor U18917 (N_18917,N_15233,N_16160);
or U18918 (N_18918,N_16155,N_15143);
nor U18919 (N_18919,N_16924,N_16221);
xnor U18920 (N_18920,N_16911,N_15890);
and U18921 (N_18921,N_15231,N_15057);
nand U18922 (N_18922,N_16671,N_15323);
xnor U18923 (N_18923,N_15173,N_16102);
or U18924 (N_18924,N_17111,N_15475);
xnor U18925 (N_18925,N_17029,N_16840);
xor U18926 (N_18926,N_15392,N_17454);
or U18927 (N_18927,N_16292,N_15583);
and U18928 (N_18928,N_15123,N_16620);
nor U18929 (N_18929,N_17019,N_15747);
and U18930 (N_18930,N_15847,N_17419);
and U18931 (N_18931,N_15063,N_16909);
or U18932 (N_18932,N_17147,N_16206);
xor U18933 (N_18933,N_15523,N_16671);
or U18934 (N_18934,N_16590,N_16365);
nand U18935 (N_18935,N_17323,N_15780);
nor U18936 (N_18936,N_15308,N_15739);
nand U18937 (N_18937,N_15889,N_16732);
and U18938 (N_18938,N_17276,N_15823);
or U18939 (N_18939,N_15213,N_16412);
nor U18940 (N_18940,N_15596,N_16364);
nor U18941 (N_18941,N_15787,N_16054);
and U18942 (N_18942,N_16583,N_15289);
or U18943 (N_18943,N_15080,N_15240);
or U18944 (N_18944,N_16257,N_17302);
and U18945 (N_18945,N_15512,N_15452);
and U18946 (N_18946,N_16505,N_17148);
nor U18947 (N_18947,N_15943,N_17166);
and U18948 (N_18948,N_16254,N_15537);
or U18949 (N_18949,N_16538,N_16581);
nor U18950 (N_18950,N_15707,N_15164);
and U18951 (N_18951,N_16983,N_15715);
xnor U18952 (N_18952,N_15381,N_16268);
xnor U18953 (N_18953,N_15940,N_16948);
xor U18954 (N_18954,N_16646,N_17181);
nor U18955 (N_18955,N_16055,N_15685);
nor U18956 (N_18956,N_16927,N_16314);
nand U18957 (N_18957,N_16525,N_15721);
nor U18958 (N_18958,N_17187,N_15041);
nor U18959 (N_18959,N_15818,N_17392);
nor U18960 (N_18960,N_17267,N_16097);
nand U18961 (N_18961,N_17131,N_15911);
xnor U18962 (N_18962,N_17252,N_15184);
nor U18963 (N_18963,N_16756,N_15353);
xor U18964 (N_18964,N_16431,N_16975);
nor U18965 (N_18965,N_16900,N_16764);
nor U18966 (N_18966,N_15671,N_16581);
xor U18967 (N_18967,N_15657,N_17183);
and U18968 (N_18968,N_16540,N_15224);
and U18969 (N_18969,N_16308,N_17171);
and U18970 (N_18970,N_15338,N_15885);
nand U18971 (N_18971,N_15967,N_15238);
nand U18972 (N_18972,N_17368,N_16812);
and U18973 (N_18973,N_16282,N_15048);
and U18974 (N_18974,N_15122,N_15055);
and U18975 (N_18975,N_17248,N_16078);
and U18976 (N_18976,N_16780,N_15985);
xnor U18977 (N_18977,N_17092,N_17449);
and U18978 (N_18978,N_16735,N_15653);
nor U18979 (N_18979,N_16176,N_15717);
xnor U18980 (N_18980,N_16141,N_15454);
nor U18981 (N_18981,N_17134,N_15933);
xnor U18982 (N_18982,N_15136,N_16828);
nor U18983 (N_18983,N_15029,N_15107);
nand U18984 (N_18984,N_16399,N_15972);
xnor U18985 (N_18985,N_15773,N_15522);
and U18986 (N_18986,N_15763,N_15884);
nor U18987 (N_18987,N_16189,N_16629);
nor U18988 (N_18988,N_15695,N_16105);
xnor U18989 (N_18989,N_15670,N_16509);
or U18990 (N_18990,N_17272,N_17328);
and U18991 (N_18991,N_17465,N_16705);
and U18992 (N_18992,N_17045,N_17281);
xnor U18993 (N_18993,N_15986,N_16154);
and U18994 (N_18994,N_16606,N_16796);
xnor U18995 (N_18995,N_17033,N_15628);
nand U18996 (N_18996,N_16951,N_16243);
or U18997 (N_18997,N_17023,N_16546);
or U18998 (N_18998,N_16740,N_17091);
nor U18999 (N_18999,N_16075,N_16146);
xor U19000 (N_19000,N_16204,N_15861);
nand U19001 (N_19001,N_15245,N_16767);
xor U19002 (N_19002,N_17089,N_15619);
nand U19003 (N_19003,N_16260,N_15064);
nor U19004 (N_19004,N_16040,N_15694);
or U19005 (N_19005,N_16651,N_16433);
xnor U19006 (N_19006,N_16846,N_16330);
nor U19007 (N_19007,N_15613,N_16779);
xor U19008 (N_19008,N_15532,N_15965);
and U19009 (N_19009,N_15369,N_16932);
and U19010 (N_19010,N_15395,N_16166);
nand U19011 (N_19011,N_16036,N_15534);
or U19012 (N_19012,N_16819,N_15541);
or U19013 (N_19013,N_17090,N_15994);
or U19014 (N_19014,N_17021,N_16583);
or U19015 (N_19015,N_16720,N_16511);
nor U19016 (N_19016,N_15881,N_17144);
or U19017 (N_19017,N_16573,N_16865);
or U19018 (N_19018,N_15015,N_15233);
or U19019 (N_19019,N_16610,N_17178);
and U19020 (N_19020,N_15349,N_15224);
xor U19021 (N_19021,N_16712,N_17136);
or U19022 (N_19022,N_15790,N_16168);
or U19023 (N_19023,N_16925,N_15170);
or U19024 (N_19024,N_17049,N_15713);
or U19025 (N_19025,N_15041,N_15663);
or U19026 (N_19026,N_16120,N_15932);
nand U19027 (N_19027,N_16691,N_16543);
nor U19028 (N_19028,N_15713,N_17199);
nand U19029 (N_19029,N_15015,N_17105);
nor U19030 (N_19030,N_16874,N_16786);
xnor U19031 (N_19031,N_16232,N_15032);
and U19032 (N_19032,N_15130,N_15790);
and U19033 (N_19033,N_15104,N_15560);
xnor U19034 (N_19034,N_16858,N_15074);
xnor U19035 (N_19035,N_15739,N_15633);
nor U19036 (N_19036,N_16791,N_15440);
or U19037 (N_19037,N_15327,N_16256);
xor U19038 (N_19038,N_16291,N_17315);
nand U19039 (N_19039,N_15721,N_15031);
or U19040 (N_19040,N_17484,N_15128);
xnor U19041 (N_19041,N_17069,N_16759);
nand U19042 (N_19042,N_15508,N_16571);
xnor U19043 (N_19043,N_16777,N_16125);
nand U19044 (N_19044,N_17077,N_15222);
and U19045 (N_19045,N_16050,N_16500);
nand U19046 (N_19046,N_16999,N_15635);
xnor U19047 (N_19047,N_16039,N_16504);
nor U19048 (N_19048,N_15258,N_15407);
nand U19049 (N_19049,N_17002,N_16541);
or U19050 (N_19050,N_16166,N_16521);
or U19051 (N_19051,N_15807,N_15094);
and U19052 (N_19052,N_15310,N_17060);
and U19053 (N_19053,N_16838,N_16141);
or U19054 (N_19054,N_15164,N_16470);
nor U19055 (N_19055,N_15044,N_16917);
and U19056 (N_19056,N_15742,N_16849);
xor U19057 (N_19057,N_15800,N_15379);
nand U19058 (N_19058,N_15126,N_16335);
and U19059 (N_19059,N_16572,N_16578);
and U19060 (N_19060,N_16634,N_17323);
nand U19061 (N_19061,N_15781,N_16089);
xor U19062 (N_19062,N_16356,N_15011);
and U19063 (N_19063,N_17087,N_15061);
or U19064 (N_19064,N_16046,N_15942);
or U19065 (N_19065,N_17213,N_17283);
nand U19066 (N_19066,N_17017,N_16075);
and U19067 (N_19067,N_16354,N_17116);
nor U19068 (N_19068,N_16160,N_15941);
nor U19069 (N_19069,N_16373,N_17161);
nand U19070 (N_19070,N_15122,N_17326);
nand U19071 (N_19071,N_15516,N_15758);
nor U19072 (N_19072,N_16349,N_16868);
and U19073 (N_19073,N_15294,N_15156);
xnor U19074 (N_19074,N_17081,N_15334);
xnor U19075 (N_19075,N_16801,N_16354);
and U19076 (N_19076,N_15646,N_17426);
and U19077 (N_19077,N_17286,N_15848);
xor U19078 (N_19078,N_15162,N_16395);
nor U19079 (N_19079,N_16909,N_16206);
or U19080 (N_19080,N_17230,N_16299);
nor U19081 (N_19081,N_16227,N_15133);
or U19082 (N_19082,N_16292,N_16119);
or U19083 (N_19083,N_16945,N_16409);
xnor U19084 (N_19084,N_16220,N_15244);
and U19085 (N_19085,N_15361,N_16880);
and U19086 (N_19086,N_16985,N_16672);
nor U19087 (N_19087,N_15841,N_16648);
nor U19088 (N_19088,N_15229,N_16931);
nand U19089 (N_19089,N_15859,N_16808);
nand U19090 (N_19090,N_17104,N_15070);
nand U19091 (N_19091,N_15871,N_17183);
xor U19092 (N_19092,N_16200,N_17183);
xor U19093 (N_19093,N_15119,N_15663);
xor U19094 (N_19094,N_16646,N_15971);
nand U19095 (N_19095,N_15149,N_17025);
nor U19096 (N_19096,N_17389,N_17138);
xnor U19097 (N_19097,N_16599,N_15315);
xnor U19098 (N_19098,N_17036,N_16117);
and U19099 (N_19099,N_17443,N_15638);
xor U19100 (N_19100,N_16369,N_15517);
and U19101 (N_19101,N_15568,N_15336);
nand U19102 (N_19102,N_15345,N_15082);
nor U19103 (N_19103,N_15885,N_16594);
nand U19104 (N_19104,N_16161,N_16910);
nand U19105 (N_19105,N_15071,N_15825);
or U19106 (N_19106,N_15221,N_16543);
xnor U19107 (N_19107,N_17072,N_16837);
nor U19108 (N_19108,N_16425,N_16666);
xnor U19109 (N_19109,N_17086,N_15920);
nor U19110 (N_19110,N_15340,N_15634);
and U19111 (N_19111,N_16820,N_17310);
nor U19112 (N_19112,N_16559,N_17441);
nand U19113 (N_19113,N_17381,N_15321);
and U19114 (N_19114,N_16575,N_16051);
xor U19115 (N_19115,N_16936,N_15031);
and U19116 (N_19116,N_15816,N_15076);
or U19117 (N_19117,N_15566,N_15318);
xnor U19118 (N_19118,N_17409,N_16368);
nand U19119 (N_19119,N_15561,N_17366);
or U19120 (N_19120,N_16875,N_15724);
nand U19121 (N_19121,N_17266,N_16288);
nand U19122 (N_19122,N_15065,N_15425);
and U19123 (N_19123,N_16323,N_17215);
nand U19124 (N_19124,N_16287,N_17424);
or U19125 (N_19125,N_15131,N_16558);
xor U19126 (N_19126,N_15726,N_15163);
or U19127 (N_19127,N_15702,N_15907);
or U19128 (N_19128,N_16473,N_15169);
nand U19129 (N_19129,N_16668,N_16727);
and U19130 (N_19130,N_15464,N_15615);
nor U19131 (N_19131,N_15281,N_17059);
and U19132 (N_19132,N_16023,N_17467);
nor U19133 (N_19133,N_16367,N_15339);
or U19134 (N_19134,N_16618,N_15974);
or U19135 (N_19135,N_16136,N_17166);
xor U19136 (N_19136,N_15817,N_15295);
xnor U19137 (N_19137,N_15727,N_15590);
xor U19138 (N_19138,N_15258,N_15496);
nor U19139 (N_19139,N_15388,N_17264);
and U19140 (N_19140,N_15174,N_17130);
xnor U19141 (N_19141,N_15286,N_15073);
or U19142 (N_19142,N_15704,N_15086);
nor U19143 (N_19143,N_15591,N_16467);
nor U19144 (N_19144,N_16322,N_17463);
nand U19145 (N_19145,N_16359,N_17320);
nor U19146 (N_19146,N_15752,N_15461);
xor U19147 (N_19147,N_16530,N_15107);
nor U19148 (N_19148,N_15527,N_16228);
nor U19149 (N_19149,N_15230,N_15173);
nand U19150 (N_19150,N_15010,N_15972);
and U19151 (N_19151,N_16240,N_16258);
nor U19152 (N_19152,N_16156,N_15629);
nor U19153 (N_19153,N_17351,N_16546);
or U19154 (N_19154,N_15785,N_17404);
nand U19155 (N_19155,N_16595,N_15049);
nand U19156 (N_19156,N_16026,N_17307);
nand U19157 (N_19157,N_15066,N_16333);
or U19158 (N_19158,N_16014,N_16690);
nand U19159 (N_19159,N_15744,N_15870);
nor U19160 (N_19160,N_15942,N_16937);
or U19161 (N_19161,N_16889,N_15512);
nor U19162 (N_19162,N_16693,N_15726);
nand U19163 (N_19163,N_16429,N_17171);
or U19164 (N_19164,N_15024,N_16399);
and U19165 (N_19165,N_16225,N_16854);
or U19166 (N_19166,N_16294,N_16816);
nor U19167 (N_19167,N_17085,N_15962);
nand U19168 (N_19168,N_15731,N_15014);
or U19169 (N_19169,N_17135,N_15534);
nor U19170 (N_19170,N_17352,N_16977);
nor U19171 (N_19171,N_16375,N_16102);
and U19172 (N_19172,N_15396,N_16371);
or U19173 (N_19173,N_17493,N_15967);
or U19174 (N_19174,N_17114,N_15868);
nand U19175 (N_19175,N_15119,N_16972);
nand U19176 (N_19176,N_15701,N_16458);
nand U19177 (N_19177,N_15845,N_16233);
or U19178 (N_19178,N_17088,N_15498);
nor U19179 (N_19179,N_17264,N_16932);
nand U19180 (N_19180,N_17248,N_15609);
nand U19181 (N_19181,N_15772,N_16234);
or U19182 (N_19182,N_16388,N_15756);
and U19183 (N_19183,N_16615,N_15499);
and U19184 (N_19184,N_16526,N_16611);
and U19185 (N_19185,N_15555,N_16823);
and U19186 (N_19186,N_15424,N_16606);
and U19187 (N_19187,N_15178,N_17339);
nor U19188 (N_19188,N_16974,N_16175);
xor U19189 (N_19189,N_15397,N_17253);
xor U19190 (N_19190,N_15578,N_16737);
or U19191 (N_19191,N_16255,N_16160);
nor U19192 (N_19192,N_15930,N_16574);
and U19193 (N_19193,N_17016,N_17011);
nor U19194 (N_19194,N_15124,N_17210);
nor U19195 (N_19195,N_15625,N_17481);
or U19196 (N_19196,N_17294,N_17132);
or U19197 (N_19197,N_16836,N_15917);
nor U19198 (N_19198,N_16663,N_16595);
xor U19199 (N_19199,N_17218,N_16215);
nor U19200 (N_19200,N_15511,N_17238);
or U19201 (N_19201,N_15228,N_16879);
or U19202 (N_19202,N_15445,N_15509);
or U19203 (N_19203,N_16181,N_15178);
nand U19204 (N_19204,N_16826,N_17457);
and U19205 (N_19205,N_16508,N_15088);
xnor U19206 (N_19206,N_15539,N_15492);
or U19207 (N_19207,N_17345,N_16471);
and U19208 (N_19208,N_17130,N_15346);
nand U19209 (N_19209,N_15521,N_15054);
or U19210 (N_19210,N_17167,N_15793);
nand U19211 (N_19211,N_15000,N_17191);
or U19212 (N_19212,N_16092,N_15145);
xnor U19213 (N_19213,N_15694,N_16024);
nor U19214 (N_19214,N_17048,N_16763);
xnor U19215 (N_19215,N_15721,N_15909);
or U19216 (N_19216,N_16674,N_15751);
and U19217 (N_19217,N_16758,N_16063);
xnor U19218 (N_19218,N_15558,N_16440);
nor U19219 (N_19219,N_15780,N_16306);
and U19220 (N_19220,N_15234,N_15412);
xor U19221 (N_19221,N_16223,N_15738);
xor U19222 (N_19222,N_16046,N_17027);
xnor U19223 (N_19223,N_17489,N_16788);
nand U19224 (N_19224,N_17493,N_15811);
xnor U19225 (N_19225,N_15420,N_16287);
and U19226 (N_19226,N_16363,N_16992);
and U19227 (N_19227,N_16094,N_15359);
xor U19228 (N_19228,N_15884,N_17115);
nand U19229 (N_19229,N_17128,N_17230);
nor U19230 (N_19230,N_16890,N_17007);
nand U19231 (N_19231,N_15332,N_16272);
xor U19232 (N_19232,N_16152,N_15522);
xnor U19233 (N_19233,N_15789,N_17464);
and U19234 (N_19234,N_16056,N_17273);
nand U19235 (N_19235,N_15858,N_15982);
and U19236 (N_19236,N_15498,N_16411);
and U19237 (N_19237,N_16932,N_17057);
and U19238 (N_19238,N_15808,N_16582);
xnor U19239 (N_19239,N_17023,N_15038);
and U19240 (N_19240,N_17481,N_15379);
xnor U19241 (N_19241,N_17044,N_15758);
and U19242 (N_19242,N_17456,N_16086);
nand U19243 (N_19243,N_15258,N_16568);
and U19244 (N_19244,N_15139,N_17227);
and U19245 (N_19245,N_16511,N_15656);
nor U19246 (N_19246,N_16278,N_15985);
xnor U19247 (N_19247,N_15445,N_15821);
or U19248 (N_19248,N_15597,N_15982);
xor U19249 (N_19249,N_15295,N_15788);
nor U19250 (N_19250,N_15684,N_16958);
nor U19251 (N_19251,N_16328,N_15804);
nor U19252 (N_19252,N_15904,N_17096);
nor U19253 (N_19253,N_16846,N_15979);
nor U19254 (N_19254,N_16856,N_15291);
or U19255 (N_19255,N_16449,N_15823);
nor U19256 (N_19256,N_16020,N_15903);
xor U19257 (N_19257,N_15221,N_15940);
xor U19258 (N_19258,N_15102,N_16278);
or U19259 (N_19259,N_15079,N_16046);
xor U19260 (N_19260,N_17183,N_15899);
xnor U19261 (N_19261,N_17107,N_17442);
or U19262 (N_19262,N_16450,N_15476);
nor U19263 (N_19263,N_15067,N_16036);
xnor U19264 (N_19264,N_15760,N_17459);
nand U19265 (N_19265,N_17402,N_16528);
and U19266 (N_19266,N_16970,N_16835);
and U19267 (N_19267,N_16434,N_16124);
or U19268 (N_19268,N_17320,N_15877);
or U19269 (N_19269,N_16564,N_17027);
nand U19270 (N_19270,N_16545,N_17032);
nand U19271 (N_19271,N_15909,N_15529);
nor U19272 (N_19272,N_15306,N_15709);
and U19273 (N_19273,N_15883,N_16091);
nand U19274 (N_19274,N_16556,N_15938);
xnor U19275 (N_19275,N_16029,N_15058);
nand U19276 (N_19276,N_15515,N_16238);
nand U19277 (N_19277,N_17138,N_15985);
and U19278 (N_19278,N_16983,N_16484);
and U19279 (N_19279,N_15917,N_15738);
and U19280 (N_19280,N_16809,N_15854);
and U19281 (N_19281,N_17275,N_15966);
nand U19282 (N_19282,N_15760,N_16909);
xor U19283 (N_19283,N_17385,N_16151);
xnor U19284 (N_19284,N_16805,N_15720);
xnor U19285 (N_19285,N_16523,N_16026);
or U19286 (N_19286,N_16077,N_15318);
xor U19287 (N_19287,N_16334,N_16023);
nor U19288 (N_19288,N_15389,N_17052);
nand U19289 (N_19289,N_15846,N_17052);
nor U19290 (N_19290,N_16436,N_16229);
and U19291 (N_19291,N_16914,N_17046);
and U19292 (N_19292,N_17245,N_15388);
nand U19293 (N_19293,N_16494,N_16284);
xnor U19294 (N_19294,N_16182,N_15312);
nand U19295 (N_19295,N_16515,N_16699);
nand U19296 (N_19296,N_17252,N_15214);
nand U19297 (N_19297,N_15794,N_15899);
xnor U19298 (N_19298,N_15119,N_15595);
and U19299 (N_19299,N_15903,N_15529);
nand U19300 (N_19300,N_15579,N_16774);
xor U19301 (N_19301,N_16882,N_17258);
nand U19302 (N_19302,N_15779,N_15222);
and U19303 (N_19303,N_15986,N_15797);
or U19304 (N_19304,N_16889,N_15704);
and U19305 (N_19305,N_17014,N_17243);
nor U19306 (N_19306,N_15212,N_15220);
nand U19307 (N_19307,N_16626,N_15999);
nand U19308 (N_19308,N_15410,N_15821);
or U19309 (N_19309,N_17048,N_16821);
and U19310 (N_19310,N_15257,N_16910);
nor U19311 (N_19311,N_16298,N_16431);
nor U19312 (N_19312,N_15381,N_17462);
or U19313 (N_19313,N_16693,N_15767);
nand U19314 (N_19314,N_15231,N_17209);
nor U19315 (N_19315,N_15984,N_16180);
and U19316 (N_19316,N_15774,N_15175);
and U19317 (N_19317,N_16158,N_15853);
xnor U19318 (N_19318,N_17068,N_16098);
or U19319 (N_19319,N_15984,N_16636);
xor U19320 (N_19320,N_16739,N_17486);
xor U19321 (N_19321,N_15750,N_17438);
nor U19322 (N_19322,N_17361,N_15036);
nand U19323 (N_19323,N_15589,N_16982);
nand U19324 (N_19324,N_16272,N_17324);
and U19325 (N_19325,N_16712,N_16785);
and U19326 (N_19326,N_16586,N_15842);
or U19327 (N_19327,N_15545,N_17190);
and U19328 (N_19328,N_16290,N_15572);
and U19329 (N_19329,N_15263,N_16546);
or U19330 (N_19330,N_15110,N_15550);
and U19331 (N_19331,N_15846,N_16628);
xor U19332 (N_19332,N_15141,N_17159);
xor U19333 (N_19333,N_15539,N_17079);
or U19334 (N_19334,N_17397,N_15400);
or U19335 (N_19335,N_15657,N_16427);
nand U19336 (N_19336,N_15416,N_16752);
xnor U19337 (N_19337,N_15026,N_15110);
or U19338 (N_19338,N_16270,N_15466);
xnor U19339 (N_19339,N_16894,N_17456);
xnor U19340 (N_19340,N_17215,N_15043);
and U19341 (N_19341,N_15075,N_15131);
and U19342 (N_19342,N_15778,N_15060);
or U19343 (N_19343,N_15670,N_17195);
nor U19344 (N_19344,N_17072,N_16208);
nand U19345 (N_19345,N_17077,N_15898);
and U19346 (N_19346,N_15304,N_15524);
nand U19347 (N_19347,N_16846,N_17036);
nand U19348 (N_19348,N_16872,N_16369);
or U19349 (N_19349,N_17037,N_15302);
or U19350 (N_19350,N_15506,N_15182);
and U19351 (N_19351,N_17263,N_16096);
or U19352 (N_19352,N_15486,N_15534);
or U19353 (N_19353,N_15356,N_16495);
nand U19354 (N_19354,N_15434,N_15749);
or U19355 (N_19355,N_15614,N_17155);
or U19356 (N_19356,N_15271,N_16150);
xor U19357 (N_19357,N_17237,N_15810);
nand U19358 (N_19358,N_17132,N_15367);
and U19359 (N_19359,N_16073,N_15228);
nand U19360 (N_19360,N_16826,N_15980);
and U19361 (N_19361,N_17496,N_17439);
nor U19362 (N_19362,N_16259,N_15099);
nor U19363 (N_19363,N_15635,N_15254);
nor U19364 (N_19364,N_16719,N_15535);
nor U19365 (N_19365,N_15814,N_15212);
or U19366 (N_19366,N_15491,N_16642);
xnor U19367 (N_19367,N_16637,N_15055);
nand U19368 (N_19368,N_15066,N_16032);
xnor U19369 (N_19369,N_16019,N_16200);
xnor U19370 (N_19370,N_17441,N_16083);
or U19371 (N_19371,N_16616,N_15285);
and U19372 (N_19372,N_16995,N_16988);
nand U19373 (N_19373,N_17016,N_16892);
nand U19374 (N_19374,N_17412,N_17469);
xor U19375 (N_19375,N_15339,N_15112);
or U19376 (N_19376,N_16522,N_16165);
nand U19377 (N_19377,N_16562,N_15420);
nor U19378 (N_19378,N_17439,N_15955);
or U19379 (N_19379,N_15583,N_17493);
or U19380 (N_19380,N_17361,N_16521);
nand U19381 (N_19381,N_16143,N_15884);
xor U19382 (N_19382,N_15125,N_16763);
nand U19383 (N_19383,N_17399,N_17321);
and U19384 (N_19384,N_15597,N_17110);
nor U19385 (N_19385,N_17044,N_15695);
nor U19386 (N_19386,N_16122,N_17080);
xnor U19387 (N_19387,N_15222,N_16511);
nand U19388 (N_19388,N_16189,N_16356);
xnor U19389 (N_19389,N_16376,N_16198);
xnor U19390 (N_19390,N_16133,N_15641);
nor U19391 (N_19391,N_17356,N_15218);
nand U19392 (N_19392,N_16364,N_16850);
and U19393 (N_19393,N_16675,N_16195);
or U19394 (N_19394,N_15924,N_15821);
and U19395 (N_19395,N_17403,N_15183);
or U19396 (N_19396,N_17313,N_16850);
and U19397 (N_19397,N_17001,N_17483);
xnor U19398 (N_19398,N_16648,N_17068);
and U19399 (N_19399,N_16239,N_16867);
and U19400 (N_19400,N_16960,N_16685);
nor U19401 (N_19401,N_15485,N_16157);
xnor U19402 (N_19402,N_17347,N_15017);
and U19403 (N_19403,N_16708,N_15487);
nand U19404 (N_19404,N_15068,N_16582);
or U19405 (N_19405,N_16632,N_16655);
and U19406 (N_19406,N_16699,N_15963);
nand U19407 (N_19407,N_16492,N_17034);
or U19408 (N_19408,N_16746,N_15276);
or U19409 (N_19409,N_15922,N_17499);
nand U19410 (N_19410,N_16317,N_15068);
nor U19411 (N_19411,N_17429,N_15036);
nor U19412 (N_19412,N_17478,N_16662);
xnor U19413 (N_19413,N_15494,N_16584);
nor U19414 (N_19414,N_15328,N_16644);
and U19415 (N_19415,N_15231,N_15657);
or U19416 (N_19416,N_15039,N_17438);
nand U19417 (N_19417,N_15970,N_17484);
nand U19418 (N_19418,N_17358,N_15620);
nor U19419 (N_19419,N_15812,N_17289);
or U19420 (N_19420,N_17260,N_16184);
nand U19421 (N_19421,N_16554,N_15785);
and U19422 (N_19422,N_16664,N_17002);
nor U19423 (N_19423,N_15792,N_17219);
nand U19424 (N_19424,N_15585,N_15216);
nor U19425 (N_19425,N_15850,N_15392);
and U19426 (N_19426,N_16014,N_15979);
and U19427 (N_19427,N_15275,N_16684);
xnor U19428 (N_19428,N_16077,N_16124);
nand U19429 (N_19429,N_16812,N_16049);
nor U19430 (N_19430,N_17173,N_16753);
or U19431 (N_19431,N_15673,N_17207);
nor U19432 (N_19432,N_16515,N_15684);
nand U19433 (N_19433,N_15934,N_17406);
nand U19434 (N_19434,N_15696,N_16492);
nor U19435 (N_19435,N_16214,N_15984);
nor U19436 (N_19436,N_15892,N_16178);
xnor U19437 (N_19437,N_16640,N_15027);
and U19438 (N_19438,N_16848,N_16711);
or U19439 (N_19439,N_16722,N_15336);
nor U19440 (N_19440,N_16758,N_17451);
nor U19441 (N_19441,N_15070,N_15190);
and U19442 (N_19442,N_15006,N_16190);
nand U19443 (N_19443,N_17027,N_16911);
and U19444 (N_19444,N_15371,N_15828);
or U19445 (N_19445,N_16003,N_15202);
nor U19446 (N_19446,N_17432,N_16000);
nand U19447 (N_19447,N_15875,N_16955);
or U19448 (N_19448,N_17141,N_16540);
and U19449 (N_19449,N_15380,N_17419);
nand U19450 (N_19450,N_16001,N_17307);
nand U19451 (N_19451,N_16762,N_15586);
nand U19452 (N_19452,N_16747,N_15698);
nand U19453 (N_19453,N_17288,N_15262);
nand U19454 (N_19454,N_16788,N_17378);
nand U19455 (N_19455,N_17357,N_15052);
nor U19456 (N_19456,N_17317,N_15990);
or U19457 (N_19457,N_15730,N_17039);
and U19458 (N_19458,N_16750,N_16749);
or U19459 (N_19459,N_15791,N_16403);
nor U19460 (N_19460,N_15716,N_16802);
nor U19461 (N_19461,N_15571,N_16446);
or U19462 (N_19462,N_16397,N_16314);
or U19463 (N_19463,N_16157,N_16978);
xor U19464 (N_19464,N_15334,N_17007);
nor U19465 (N_19465,N_15541,N_15106);
or U19466 (N_19466,N_16801,N_16426);
or U19467 (N_19467,N_17055,N_16103);
xnor U19468 (N_19468,N_16200,N_16503);
xor U19469 (N_19469,N_15954,N_16230);
xnor U19470 (N_19470,N_17339,N_15177);
and U19471 (N_19471,N_17222,N_16137);
nor U19472 (N_19472,N_15134,N_16394);
nand U19473 (N_19473,N_15346,N_16667);
and U19474 (N_19474,N_16933,N_17296);
nand U19475 (N_19475,N_16328,N_16268);
nand U19476 (N_19476,N_16344,N_15556);
and U19477 (N_19477,N_15614,N_16922);
nor U19478 (N_19478,N_16225,N_16276);
or U19479 (N_19479,N_16995,N_17017);
nand U19480 (N_19480,N_17209,N_17445);
nand U19481 (N_19481,N_16021,N_16186);
xor U19482 (N_19482,N_16900,N_15058);
or U19483 (N_19483,N_15961,N_16924);
nor U19484 (N_19484,N_15903,N_17455);
nor U19485 (N_19485,N_17404,N_17345);
nor U19486 (N_19486,N_17069,N_16580);
nor U19487 (N_19487,N_16863,N_16985);
or U19488 (N_19488,N_16467,N_16507);
or U19489 (N_19489,N_15148,N_17499);
nor U19490 (N_19490,N_15463,N_15773);
nand U19491 (N_19491,N_15962,N_17262);
nor U19492 (N_19492,N_15328,N_15602);
nand U19493 (N_19493,N_17211,N_16492);
and U19494 (N_19494,N_17496,N_15864);
nand U19495 (N_19495,N_16666,N_16450);
or U19496 (N_19496,N_15581,N_17333);
nand U19497 (N_19497,N_16832,N_16548);
nor U19498 (N_19498,N_15189,N_16022);
and U19499 (N_19499,N_15321,N_15854);
nor U19500 (N_19500,N_17453,N_15841);
xnor U19501 (N_19501,N_17299,N_15356);
or U19502 (N_19502,N_15237,N_17277);
or U19503 (N_19503,N_16688,N_17056);
or U19504 (N_19504,N_15198,N_15689);
xor U19505 (N_19505,N_16525,N_16632);
nor U19506 (N_19506,N_17211,N_16896);
and U19507 (N_19507,N_15865,N_17167);
nor U19508 (N_19508,N_15426,N_16711);
or U19509 (N_19509,N_16152,N_16222);
nand U19510 (N_19510,N_17329,N_15692);
nor U19511 (N_19511,N_15383,N_16770);
nor U19512 (N_19512,N_15611,N_17074);
and U19513 (N_19513,N_16464,N_15153);
and U19514 (N_19514,N_15602,N_17317);
and U19515 (N_19515,N_16276,N_16221);
and U19516 (N_19516,N_16807,N_16959);
and U19517 (N_19517,N_17218,N_16552);
or U19518 (N_19518,N_16054,N_16994);
nor U19519 (N_19519,N_15130,N_15604);
nor U19520 (N_19520,N_16101,N_15923);
or U19521 (N_19521,N_15226,N_15301);
or U19522 (N_19522,N_16852,N_15437);
and U19523 (N_19523,N_16974,N_17155);
nor U19524 (N_19524,N_16074,N_15880);
xnor U19525 (N_19525,N_17233,N_16554);
xor U19526 (N_19526,N_15023,N_17388);
and U19527 (N_19527,N_16431,N_16573);
or U19528 (N_19528,N_17071,N_15451);
nand U19529 (N_19529,N_15216,N_17273);
or U19530 (N_19530,N_15606,N_16966);
xnor U19531 (N_19531,N_15154,N_15586);
xnor U19532 (N_19532,N_15982,N_17431);
nor U19533 (N_19533,N_16006,N_16098);
or U19534 (N_19534,N_17170,N_15118);
xor U19535 (N_19535,N_16651,N_15052);
nand U19536 (N_19536,N_16257,N_16041);
xnor U19537 (N_19537,N_17436,N_15092);
or U19538 (N_19538,N_17017,N_16150);
or U19539 (N_19539,N_15011,N_15606);
nand U19540 (N_19540,N_15049,N_15207);
xor U19541 (N_19541,N_16918,N_16144);
xor U19542 (N_19542,N_16653,N_17020);
nor U19543 (N_19543,N_17419,N_16681);
nor U19544 (N_19544,N_16447,N_15261);
xnor U19545 (N_19545,N_15084,N_16845);
nand U19546 (N_19546,N_17160,N_16723);
and U19547 (N_19547,N_16462,N_16482);
nor U19548 (N_19548,N_16686,N_15425);
nor U19549 (N_19549,N_16724,N_15530);
nand U19550 (N_19550,N_17344,N_15814);
xor U19551 (N_19551,N_16122,N_16771);
xnor U19552 (N_19552,N_16938,N_17111);
and U19553 (N_19553,N_15553,N_15776);
or U19554 (N_19554,N_15249,N_15570);
and U19555 (N_19555,N_16836,N_15878);
nor U19556 (N_19556,N_15805,N_15382);
or U19557 (N_19557,N_16001,N_16586);
nand U19558 (N_19558,N_15383,N_16005);
and U19559 (N_19559,N_15874,N_17463);
nand U19560 (N_19560,N_17390,N_16377);
nand U19561 (N_19561,N_15145,N_16010);
nand U19562 (N_19562,N_16666,N_17217);
nor U19563 (N_19563,N_15528,N_17050);
and U19564 (N_19564,N_15157,N_15900);
or U19565 (N_19565,N_16806,N_17393);
xnor U19566 (N_19566,N_17363,N_16571);
or U19567 (N_19567,N_16640,N_16931);
nand U19568 (N_19568,N_15327,N_15357);
nor U19569 (N_19569,N_16094,N_17142);
xor U19570 (N_19570,N_15813,N_16407);
nand U19571 (N_19571,N_15543,N_15074);
nor U19572 (N_19572,N_16414,N_16486);
or U19573 (N_19573,N_15796,N_16064);
or U19574 (N_19574,N_16405,N_16365);
and U19575 (N_19575,N_17357,N_16053);
nor U19576 (N_19576,N_17208,N_16668);
or U19577 (N_19577,N_17178,N_16951);
and U19578 (N_19578,N_17234,N_15703);
nand U19579 (N_19579,N_16740,N_15138);
xor U19580 (N_19580,N_17109,N_15258);
and U19581 (N_19581,N_15905,N_17419);
nand U19582 (N_19582,N_15631,N_17372);
and U19583 (N_19583,N_17284,N_16876);
nand U19584 (N_19584,N_17102,N_15742);
xor U19585 (N_19585,N_15978,N_17043);
or U19586 (N_19586,N_15433,N_17441);
or U19587 (N_19587,N_15080,N_17225);
xor U19588 (N_19588,N_17381,N_16405);
nor U19589 (N_19589,N_15030,N_15788);
nor U19590 (N_19590,N_16560,N_15664);
xnor U19591 (N_19591,N_15433,N_16467);
nor U19592 (N_19592,N_17348,N_16535);
nor U19593 (N_19593,N_17208,N_17369);
nand U19594 (N_19594,N_16224,N_16588);
nand U19595 (N_19595,N_16321,N_15469);
xnor U19596 (N_19596,N_16817,N_15578);
nor U19597 (N_19597,N_16568,N_16984);
nand U19598 (N_19598,N_17068,N_15269);
nand U19599 (N_19599,N_15306,N_15824);
nor U19600 (N_19600,N_17351,N_16492);
nor U19601 (N_19601,N_16317,N_15709);
xor U19602 (N_19602,N_17365,N_16274);
nor U19603 (N_19603,N_17426,N_16850);
nand U19604 (N_19604,N_17166,N_16725);
nor U19605 (N_19605,N_15608,N_16580);
or U19606 (N_19606,N_16870,N_17234);
nand U19607 (N_19607,N_16984,N_15734);
nand U19608 (N_19608,N_16914,N_16816);
or U19609 (N_19609,N_17105,N_15025);
nor U19610 (N_19610,N_16879,N_16843);
xor U19611 (N_19611,N_15326,N_15539);
nand U19612 (N_19612,N_15135,N_16393);
nor U19613 (N_19613,N_17438,N_15152);
or U19614 (N_19614,N_16297,N_16405);
or U19615 (N_19615,N_17472,N_16100);
nor U19616 (N_19616,N_16545,N_15556);
nand U19617 (N_19617,N_16716,N_16451);
nor U19618 (N_19618,N_15629,N_15432);
nand U19619 (N_19619,N_16602,N_15258);
nor U19620 (N_19620,N_15043,N_15324);
and U19621 (N_19621,N_15433,N_16721);
or U19622 (N_19622,N_16754,N_16043);
or U19623 (N_19623,N_15163,N_15293);
xnor U19624 (N_19624,N_16235,N_15961);
and U19625 (N_19625,N_17052,N_17046);
or U19626 (N_19626,N_16259,N_15906);
and U19627 (N_19627,N_16848,N_16047);
xnor U19628 (N_19628,N_16091,N_15836);
xnor U19629 (N_19629,N_15517,N_15025);
or U19630 (N_19630,N_17213,N_16306);
xnor U19631 (N_19631,N_15647,N_16837);
or U19632 (N_19632,N_17070,N_15696);
and U19633 (N_19633,N_17444,N_15641);
or U19634 (N_19634,N_16296,N_17170);
xor U19635 (N_19635,N_16675,N_17354);
nand U19636 (N_19636,N_16214,N_17407);
and U19637 (N_19637,N_16430,N_15468);
nor U19638 (N_19638,N_15746,N_15220);
xnor U19639 (N_19639,N_17019,N_17176);
nor U19640 (N_19640,N_16509,N_15457);
xor U19641 (N_19641,N_17195,N_17253);
and U19642 (N_19642,N_16067,N_16624);
nand U19643 (N_19643,N_16098,N_16737);
or U19644 (N_19644,N_15483,N_15787);
or U19645 (N_19645,N_15948,N_16613);
xnor U19646 (N_19646,N_15284,N_15331);
or U19647 (N_19647,N_17032,N_16819);
nand U19648 (N_19648,N_16234,N_17100);
xnor U19649 (N_19649,N_16888,N_15551);
nand U19650 (N_19650,N_16217,N_15526);
and U19651 (N_19651,N_16389,N_15146);
nor U19652 (N_19652,N_15826,N_16135);
nor U19653 (N_19653,N_16468,N_17480);
xor U19654 (N_19654,N_16298,N_17061);
nand U19655 (N_19655,N_16782,N_15996);
nand U19656 (N_19656,N_17020,N_15880);
and U19657 (N_19657,N_16562,N_16913);
nor U19658 (N_19658,N_17117,N_16012);
nor U19659 (N_19659,N_16704,N_17070);
or U19660 (N_19660,N_15963,N_15240);
nand U19661 (N_19661,N_16288,N_17475);
nand U19662 (N_19662,N_15618,N_15550);
and U19663 (N_19663,N_16727,N_15360);
and U19664 (N_19664,N_17491,N_17381);
nand U19665 (N_19665,N_17465,N_16219);
or U19666 (N_19666,N_17427,N_17014);
or U19667 (N_19667,N_15534,N_15666);
and U19668 (N_19668,N_17030,N_15776);
and U19669 (N_19669,N_16358,N_15728);
nand U19670 (N_19670,N_15499,N_17487);
xnor U19671 (N_19671,N_17173,N_16489);
nor U19672 (N_19672,N_16058,N_15402);
or U19673 (N_19673,N_16243,N_16923);
nor U19674 (N_19674,N_16068,N_17168);
xnor U19675 (N_19675,N_15878,N_16246);
and U19676 (N_19676,N_16770,N_15152);
or U19677 (N_19677,N_16652,N_17385);
nor U19678 (N_19678,N_17220,N_15195);
nor U19679 (N_19679,N_16187,N_16162);
xnor U19680 (N_19680,N_15734,N_15752);
or U19681 (N_19681,N_16806,N_15581);
nor U19682 (N_19682,N_16145,N_15922);
and U19683 (N_19683,N_17340,N_15147);
nand U19684 (N_19684,N_15886,N_15563);
and U19685 (N_19685,N_16336,N_16810);
and U19686 (N_19686,N_16467,N_16721);
or U19687 (N_19687,N_15786,N_16283);
nor U19688 (N_19688,N_15331,N_15806);
nand U19689 (N_19689,N_17443,N_16032);
or U19690 (N_19690,N_17469,N_15996);
xor U19691 (N_19691,N_17037,N_15989);
nand U19692 (N_19692,N_15131,N_15722);
and U19693 (N_19693,N_16804,N_16576);
and U19694 (N_19694,N_16828,N_15509);
and U19695 (N_19695,N_16336,N_15659);
nand U19696 (N_19696,N_16364,N_17276);
xnor U19697 (N_19697,N_16252,N_15069);
nor U19698 (N_19698,N_15355,N_15075);
or U19699 (N_19699,N_17253,N_15619);
nand U19700 (N_19700,N_16680,N_16001);
nor U19701 (N_19701,N_16448,N_17009);
and U19702 (N_19702,N_17169,N_17287);
and U19703 (N_19703,N_16139,N_15133);
and U19704 (N_19704,N_17392,N_15221);
nor U19705 (N_19705,N_16748,N_16502);
nand U19706 (N_19706,N_15115,N_16327);
nand U19707 (N_19707,N_16037,N_15266);
nand U19708 (N_19708,N_16694,N_16797);
or U19709 (N_19709,N_16785,N_15176);
nor U19710 (N_19710,N_17293,N_16144);
nand U19711 (N_19711,N_15441,N_15631);
nor U19712 (N_19712,N_17296,N_15833);
and U19713 (N_19713,N_16016,N_15301);
or U19714 (N_19714,N_16426,N_15072);
and U19715 (N_19715,N_16781,N_16765);
xor U19716 (N_19716,N_16335,N_15862);
and U19717 (N_19717,N_16993,N_15914);
nand U19718 (N_19718,N_16515,N_16610);
or U19719 (N_19719,N_15765,N_16248);
nand U19720 (N_19720,N_16469,N_16463);
or U19721 (N_19721,N_15852,N_15183);
or U19722 (N_19722,N_15964,N_16379);
or U19723 (N_19723,N_15991,N_17267);
or U19724 (N_19724,N_16930,N_17271);
and U19725 (N_19725,N_16579,N_16645);
and U19726 (N_19726,N_16286,N_16519);
nor U19727 (N_19727,N_16052,N_15317);
nor U19728 (N_19728,N_15365,N_15190);
nand U19729 (N_19729,N_16963,N_17350);
nand U19730 (N_19730,N_16392,N_17388);
and U19731 (N_19731,N_15739,N_16700);
and U19732 (N_19732,N_16689,N_16565);
xor U19733 (N_19733,N_16869,N_17115);
and U19734 (N_19734,N_16280,N_17268);
nand U19735 (N_19735,N_16866,N_16572);
xnor U19736 (N_19736,N_17399,N_17384);
nand U19737 (N_19737,N_16245,N_16162);
nor U19738 (N_19738,N_16947,N_17394);
and U19739 (N_19739,N_16936,N_15534);
and U19740 (N_19740,N_16440,N_16946);
or U19741 (N_19741,N_15318,N_15284);
xor U19742 (N_19742,N_15489,N_15088);
xnor U19743 (N_19743,N_15765,N_15729);
xnor U19744 (N_19744,N_15881,N_15988);
or U19745 (N_19745,N_17118,N_16951);
nand U19746 (N_19746,N_16522,N_15031);
and U19747 (N_19747,N_16360,N_17275);
nand U19748 (N_19748,N_16132,N_16198);
and U19749 (N_19749,N_16813,N_15076);
xnor U19750 (N_19750,N_16111,N_15690);
or U19751 (N_19751,N_17044,N_17249);
and U19752 (N_19752,N_16374,N_16487);
xnor U19753 (N_19753,N_16949,N_17362);
nand U19754 (N_19754,N_17356,N_16520);
nor U19755 (N_19755,N_15264,N_15164);
and U19756 (N_19756,N_15887,N_15444);
nor U19757 (N_19757,N_17496,N_15910);
nor U19758 (N_19758,N_15897,N_15892);
nand U19759 (N_19759,N_15022,N_16460);
or U19760 (N_19760,N_16516,N_16289);
nor U19761 (N_19761,N_16694,N_15606);
xor U19762 (N_19762,N_16642,N_16426);
or U19763 (N_19763,N_16900,N_16774);
nor U19764 (N_19764,N_17020,N_17123);
and U19765 (N_19765,N_15461,N_16995);
nand U19766 (N_19766,N_16269,N_17162);
nand U19767 (N_19767,N_16800,N_16216);
and U19768 (N_19768,N_15507,N_17004);
or U19769 (N_19769,N_17142,N_15886);
nand U19770 (N_19770,N_15574,N_16386);
nor U19771 (N_19771,N_15913,N_16823);
and U19772 (N_19772,N_15534,N_16753);
and U19773 (N_19773,N_15349,N_16137);
or U19774 (N_19774,N_15681,N_15706);
nor U19775 (N_19775,N_15844,N_17318);
or U19776 (N_19776,N_17165,N_16012);
and U19777 (N_19777,N_16418,N_16469);
xnor U19778 (N_19778,N_16797,N_15316);
and U19779 (N_19779,N_15422,N_16846);
and U19780 (N_19780,N_15957,N_17052);
nand U19781 (N_19781,N_16419,N_15584);
xnor U19782 (N_19782,N_16813,N_16043);
and U19783 (N_19783,N_15767,N_16784);
and U19784 (N_19784,N_16321,N_15665);
and U19785 (N_19785,N_16879,N_17190);
nand U19786 (N_19786,N_15044,N_17231);
or U19787 (N_19787,N_17441,N_16972);
nor U19788 (N_19788,N_16189,N_17306);
nand U19789 (N_19789,N_16087,N_15099);
nand U19790 (N_19790,N_15715,N_15142);
or U19791 (N_19791,N_17253,N_16799);
xnor U19792 (N_19792,N_15555,N_16953);
xor U19793 (N_19793,N_17376,N_15267);
xor U19794 (N_19794,N_15093,N_17139);
xnor U19795 (N_19795,N_15690,N_16544);
nor U19796 (N_19796,N_15009,N_16402);
nand U19797 (N_19797,N_16232,N_15386);
or U19798 (N_19798,N_17217,N_15232);
and U19799 (N_19799,N_15026,N_15060);
and U19800 (N_19800,N_17307,N_17164);
or U19801 (N_19801,N_16934,N_17302);
or U19802 (N_19802,N_16322,N_15041);
nand U19803 (N_19803,N_16637,N_17427);
xor U19804 (N_19804,N_16401,N_16789);
and U19805 (N_19805,N_15902,N_15221);
nor U19806 (N_19806,N_15312,N_16293);
nand U19807 (N_19807,N_15966,N_16660);
xor U19808 (N_19808,N_16803,N_15400);
xor U19809 (N_19809,N_17022,N_15064);
and U19810 (N_19810,N_15482,N_16600);
nand U19811 (N_19811,N_16706,N_16565);
and U19812 (N_19812,N_16240,N_15780);
nor U19813 (N_19813,N_16589,N_16276);
xnor U19814 (N_19814,N_15568,N_16164);
nor U19815 (N_19815,N_16642,N_15698);
nand U19816 (N_19816,N_16777,N_15600);
xor U19817 (N_19817,N_15146,N_16040);
and U19818 (N_19818,N_15509,N_15728);
or U19819 (N_19819,N_15625,N_16798);
xnor U19820 (N_19820,N_16188,N_16457);
nand U19821 (N_19821,N_15569,N_15005);
nand U19822 (N_19822,N_15575,N_17131);
and U19823 (N_19823,N_17365,N_15216);
xnor U19824 (N_19824,N_15104,N_16958);
nor U19825 (N_19825,N_16024,N_15598);
nor U19826 (N_19826,N_15832,N_16155);
or U19827 (N_19827,N_17048,N_15061);
nand U19828 (N_19828,N_16573,N_16498);
and U19829 (N_19829,N_15960,N_16870);
or U19830 (N_19830,N_15464,N_16885);
nand U19831 (N_19831,N_16141,N_15146);
and U19832 (N_19832,N_15519,N_16359);
and U19833 (N_19833,N_15208,N_16972);
nor U19834 (N_19834,N_15090,N_16031);
nand U19835 (N_19835,N_15685,N_16261);
nor U19836 (N_19836,N_15108,N_16399);
xnor U19837 (N_19837,N_16805,N_17453);
or U19838 (N_19838,N_16619,N_15349);
nand U19839 (N_19839,N_15538,N_16074);
nand U19840 (N_19840,N_16933,N_16275);
and U19841 (N_19841,N_15450,N_16009);
or U19842 (N_19842,N_17418,N_15350);
nand U19843 (N_19843,N_17450,N_15011);
and U19844 (N_19844,N_16563,N_15491);
xor U19845 (N_19845,N_17051,N_17496);
xor U19846 (N_19846,N_16341,N_16332);
xor U19847 (N_19847,N_16420,N_16626);
xnor U19848 (N_19848,N_15884,N_15887);
xor U19849 (N_19849,N_17432,N_15829);
or U19850 (N_19850,N_16788,N_15659);
and U19851 (N_19851,N_15261,N_16338);
or U19852 (N_19852,N_16784,N_16067);
nor U19853 (N_19853,N_15576,N_15545);
and U19854 (N_19854,N_17158,N_16412);
and U19855 (N_19855,N_15349,N_16882);
or U19856 (N_19856,N_16787,N_16211);
xnor U19857 (N_19857,N_16652,N_15978);
xnor U19858 (N_19858,N_15183,N_15752);
nand U19859 (N_19859,N_16990,N_15908);
or U19860 (N_19860,N_16815,N_16746);
xor U19861 (N_19861,N_15320,N_15865);
and U19862 (N_19862,N_16903,N_17044);
and U19863 (N_19863,N_15131,N_16122);
nand U19864 (N_19864,N_16145,N_16812);
and U19865 (N_19865,N_15520,N_15160);
nor U19866 (N_19866,N_15747,N_16594);
nand U19867 (N_19867,N_15855,N_15592);
nand U19868 (N_19868,N_17337,N_17233);
or U19869 (N_19869,N_15630,N_16207);
nor U19870 (N_19870,N_17072,N_16080);
nor U19871 (N_19871,N_16032,N_17340);
or U19872 (N_19872,N_17023,N_15546);
xnor U19873 (N_19873,N_15189,N_15739);
nor U19874 (N_19874,N_17016,N_17493);
nand U19875 (N_19875,N_16562,N_15344);
nand U19876 (N_19876,N_17025,N_16457);
nand U19877 (N_19877,N_16188,N_17142);
nor U19878 (N_19878,N_15015,N_15490);
nand U19879 (N_19879,N_17044,N_16077);
xor U19880 (N_19880,N_17246,N_15439);
and U19881 (N_19881,N_16553,N_15487);
xor U19882 (N_19882,N_16591,N_17318);
or U19883 (N_19883,N_16214,N_15145);
nand U19884 (N_19884,N_15751,N_16682);
nor U19885 (N_19885,N_16842,N_16788);
xnor U19886 (N_19886,N_16419,N_16277);
or U19887 (N_19887,N_17024,N_16244);
xor U19888 (N_19888,N_16703,N_17215);
nand U19889 (N_19889,N_16091,N_16514);
nand U19890 (N_19890,N_17439,N_17049);
or U19891 (N_19891,N_17156,N_17097);
or U19892 (N_19892,N_16875,N_16580);
xnor U19893 (N_19893,N_15624,N_16887);
xor U19894 (N_19894,N_15160,N_16805);
nor U19895 (N_19895,N_16055,N_17491);
xnor U19896 (N_19896,N_16627,N_15594);
nand U19897 (N_19897,N_16306,N_17277);
nand U19898 (N_19898,N_17198,N_16412);
nand U19899 (N_19899,N_17169,N_15491);
and U19900 (N_19900,N_15709,N_15804);
nand U19901 (N_19901,N_17399,N_17190);
or U19902 (N_19902,N_16646,N_16642);
nor U19903 (N_19903,N_15694,N_15281);
nor U19904 (N_19904,N_15421,N_16667);
xor U19905 (N_19905,N_16999,N_15759);
nand U19906 (N_19906,N_15959,N_15136);
or U19907 (N_19907,N_16975,N_15506);
nand U19908 (N_19908,N_15704,N_15572);
and U19909 (N_19909,N_15500,N_16253);
nand U19910 (N_19910,N_16647,N_15403);
xnor U19911 (N_19911,N_15770,N_15907);
and U19912 (N_19912,N_16934,N_16048);
and U19913 (N_19913,N_16593,N_17263);
and U19914 (N_19914,N_15092,N_16728);
and U19915 (N_19915,N_15393,N_16014);
or U19916 (N_19916,N_17356,N_16120);
and U19917 (N_19917,N_15556,N_15870);
nand U19918 (N_19918,N_15567,N_16434);
or U19919 (N_19919,N_17442,N_16453);
xnor U19920 (N_19920,N_17267,N_17025);
or U19921 (N_19921,N_15045,N_16888);
or U19922 (N_19922,N_16363,N_16662);
or U19923 (N_19923,N_16639,N_16105);
xor U19924 (N_19924,N_16902,N_15027);
nand U19925 (N_19925,N_15093,N_15603);
and U19926 (N_19926,N_15166,N_15817);
nand U19927 (N_19927,N_16424,N_17375);
and U19928 (N_19928,N_16912,N_16294);
or U19929 (N_19929,N_16846,N_17249);
xor U19930 (N_19930,N_15954,N_15235);
nand U19931 (N_19931,N_16302,N_16798);
or U19932 (N_19932,N_16841,N_16785);
and U19933 (N_19933,N_16515,N_15201);
nand U19934 (N_19934,N_15821,N_16699);
or U19935 (N_19935,N_15486,N_16945);
nor U19936 (N_19936,N_17469,N_15263);
nor U19937 (N_19937,N_15264,N_17242);
or U19938 (N_19938,N_17315,N_15191);
and U19939 (N_19939,N_15872,N_15561);
xor U19940 (N_19940,N_16780,N_16421);
nor U19941 (N_19941,N_16142,N_16374);
and U19942 (N_19942,N_15943,N_16078);
nor U19943 (N_19943,N_15813,N_15493);
nor U19944 (N_19944,N_17330,N_16097);
nand U19945 (N_19945,N_17138,N_16901);
or U19946 (N_19946,N_16102,N_16357);
or U19947 (N_19947,N_16292,N_15833);
xnor U19948 (N_19948,N_16874,N_16017);
and U19949 (N_19949,N_15501,N_15937);
or U19950 (N_19950,N_16666,N_16292);
nor U19951 (N_19951,N_17363,N_15184);
nor U19952 (N_19952,N_17079,N_16831);
or U19953 (N_19953,N_15644,N_17406);
nor U19954 (N_19954,N_15652,N_15014);
or U19955 (N_19955,N_17370,N_15644);
xor U19956 (N_19956,N_15058,N_16787);
nand U19957 (N_19957,N_17359,N_15795);
nand U19958 (N_19958,N_16250,N_16913);
nor U19959 (N_19959,N_16743,N_16523);
xor U19960 (N_19960,N_17363,N_15783);
nor U19961 (N_19961,N_16995,N_17153);
xor U19962 (N_19962,N_15001,N_17031);
nand U19963 (N_19963,N_16693,N_17351);
or U19964 (N_19964,N_15439,N_17470);
and U19965 (N_19965,N_15489,N_17074);
nand U19966 (N_19966,N_15186,N_16525);
nor U19967 (N_19967,N_16928,N_15807);
or U19968 (N_19968,N_17176,N_16254);
and U19969 (N_19969,N_16492,N_17384);
nand U19970 (N_19970,N_17037,N_16723);
or U19971 (N_19971,N_15550,N_16053);
or U19972 (N_19972,N_17389,N_16991);
and U19973 (N_19973,N_16389,N_15691);
and U19974 (N_19974,N_16494,N_15621);
or U19975 (N_19975,N_17245,N_15613);
nor U19976 (N_19976,N_16713,N_16720);
and U19977 (N_19977,N_17223,N_15445);
and U19978 (N_19978,N_16597,N_16474);
and U19979 (N_19979,N_15740,N_15806);
xnor U19980 (N_19980,N_17129,N_17100);
nand U19981 (N_19981,N_17413,N_16742);
xnor U19982 (N_19982,N_15973,N_15818);
xnor U19983 (N_19983,N_16563,N_16623);
and U19984 (N_19984,N_17130,N_17224);
and U19985 (N_19985,N_16694,N_16946);
nand U19986 (N_19986,N_15197,N_15621);
nor U19987 (N_19987,N_15533,N_15637);
nand U19988 (N_19988,N_16470,N_16397);
xor U19989 (N_19989,N_15133,N_15090);
nand U19990 (N_19990,N_15576,N_16169);
xor U19991 (N_19991,N_16778,N_15750);
xor U19992 (N_19992,N_17110,N_15651);
and U19993 (N_19993,N_16866,N_16190);
or U19994 (N_19994,N_15615,N_16978);
nor U19995 (N_19995,N_15014,N_15400);
or U19996 (N_19996,N_15832,N_15161);
xor U19997 (N_19997,N_16637,N_15280);
xor U19998 (N_19998,N_16863,N_15504);
nor U19999 (N_19999,N_17303,N_16904);
xnor U20000 (N_20000,N_19033,N_19111);
and U20001 (N_20001,N_19044,N_17965);
and U20002 (N_20002,N_18434,N_17755);
nor U20003 (N_20003,N_18675,N_19160);
and U20004 (N_20004,N_19161,N_19934);
or U20005 (N_20005,N_19723,N_18062);
and U20006 (N_20006,N_18588,N_19418);
nor U20007 (N_20007,N_18228,N_18332);
and U20008 (N_20008,N_19185,N_18641);
and U20009 (N_20009,N_19046,N_19110);
nand U20010 (N_20010,N_18803,N_19606);
nand U20011 (N_20011,N_17563,N_19931);
nor U20012 (N_20012,N_18432,N_18320);
or U20013 (N_20013,N_19688,N_18623);
or U20014 (N_20014,N_19247,N_19602);
xnor U20015 (N_20015,N_19375,N_19292);
xnor U20016 (N_20016,N_18405,N_19305);
xor U20017 (N_20017,N_17623,N_19576);
and U20018 (N_20018,N_18037,N_19995);
and U20019 (N_20019,N_19999,N_19028);
or U20020 (N_20020,N_18582,N_19861);
and U20021 (N_20021,N_17818,N_18518);
nor U20022 (N_20022,N_19960,N_18970);
xnor U20023 (N_20023,N_18289,N_18239);
nand U20024 (N_20024,N_19821,N_17997);
nor U20025 (N_20025,N_17947,N_19684);
nand U20026 (N_20026,N_17772,N_18330);
and U20027 (N_20027,N_19683,N_17726);
or U20028 (N_20028,N_19729,N_17658);
and U20029 (N_20029,N_17595,N_18103);
and U20030 (N_20030,N_17695,N_18761);
or U20031 (N_20031,N_17647,N_17979);
and U20032 (N_20032,N_18942,N_18141);
and U20033 (N_20033,N_18387,N_19912);
or U20034 (N_20034,N_18012,N_19433);
nor U20035 (N_20035,N_18030,N_19014);
xor U20036 (N_20036,N_18350,N_17984);
xor U20037 (N_20037,N_19484,N_19927);
nand U20038 (N_20038,N_19508,N_19012);
nor U20039 (N_20039,N_18979,N_19826);
xor U20040 (N_20040,N_18143,N_18581);
nand U20041 (N_20041,N_17787,N_18776);
or U20042 (N_20042,N_18064,N_17759);
nand U20043 (N_20043,N_18634,N_19444);
and U20044 (N_20044,N_19517,N_17580);
or U20045 (N_20045,N_19037,N_17769);
nor U20046 (N_20046,N_18895,N_19806);
nand U20047 (N_20047,N_19896,N_19592);
and U20048 (N_20048,N_17817,N_18295);
and U20049 (N_20049,N_19794,N_19678);
and U20050 (N_20050,N_17604,N_18080);
nor U20051 (N_20051,N_18626,N_17730);
and U20052 (N_20052,N_18782,N_18959);
nand U20053 (N_20053,N_19890,N_17971);
or U20054 (N_20054,N_18002,N_18000);
nor U20055 (N_20055,N_18251,N_19768);
or U20056 (N_20056,N_19724,N_19280);
and U20057 (N_20057,N_19289,N_19608);
or U20058 (N_20058,N_19139,N_19385);
nand U20059 (N_20059,N_19184,N_19051);
nand U20060 (N_20060,N_17662,N_19640);
and U20061 (N_20061,N_18740,N_17773);
nor U20062 (N_20062,N_18887,N_19257);
nand U20063 (N_20063,N_17812,N_19879);
or U20064 (N_20064,N_18913,N_18372);
or U20065 (N_20065,N_18953,N_18880);
xor U20066 (N_20066,N_18016,N_19963);
or U20067 (N_20067,N_19035,N_17807);
xnor U20068 (N_20068,N_17879,N_19314);
or U20069 (N_20069,N_17919,N_17592);
and U20070 (N_20070,N_19760,N_18408);
or U20071 (N_20071,N_18273,N_18778);
or U20072 (N_20072,N_17705,N_17936);
and U20073 (N_20073,N_18791,N_17878);
nor U20074 (N_20074,N_19603,N_17646);
and U20075 (N_20075,N_19326,N_19453);
nand U20076 (N_20076,N_17915,N_18823);
nand U20077 (N_20077,N_19054,N_18863);
or U20078 (N_20078,N_18858,N_19210);
nand U20079 (N_20079,N_17576,N_18629);
nor U20080 (N_20080,N_18914,N_19565);
and U20081 (N_20081,N_19932,N_18697);
nand U20082 (N_20082,N_17959,N_17678);
or U20083 (N_20083,N_18991,N_19483);
nor U20084 (N_20084,N_19168,N_18255);
xnor U20085 (N_20085,N_19798,N_18241);
and U20086 (N_20086,N_18671,N_17581);
nand U20087 (N_20087,N_19598,N_18260);
nor U20088 (N_20088,N_18958,N_19228);
and U20089 (N_20089,N_18083,N_19884);
and U20090 (N_20090,N_19980,N_19062);
nor U20091 (N_20091,N_19425,N_19911);
or U20092 (N_20092,N_19260,N_18164);
or U20093 (N_20093,N_18476,N_18804);
and U20094 (N_20094,N_18053,N_19659);
xnor U20095 (N_20095,N_19795,N_19836);
nand U20096 (N_20096,N_18955,N_18221);
or U20097 (N_20097,N_18178,N_18345);
nor U20098 (N_20098,N_19880,N_19384);
and U20099 (N_20099,N_18940,N_18192);
nor U20100 (N_20100,N_19163,N_19616);
xor U20101 (N_20101,N_18831,N_17501);
nor U20102 (N_20102,N_17949,N_17672);
nor U20103 (N_20103,N_18682,N_17731);
nand U20104 (N_20104,N_18988,N_19923);
or U20105 (N_20105,N_18878,N_18706);
and U20106 (N_20106,N_19154,N_19547);
and U20107 (N_20107,N_17738,N_18833);
nand U20108 (N_20108,N_19568,N_18166);
nand U20109 (N_20109,N_19601,N_18355);
nor U20110 (N_20110,N_17920,N_19561);
nand U20111 (N_20111,N_18751,N_19859);
or U20112 (N_20112,N_18034,N_19221);
or U20113 (N_20113,N_18743,N_17846);
nor U20114 (N_20114,N_17703,N_19446);
and U20115 (N_20115,N_18898,N_18720);
and U20116 (N_20116,N_18153,N_19588);
nand U20117 (N_20117,N_17924,N_19709);
nand U20118 (N_20118,N_19748,N_19593);
nand U20119 (N_20119,N_18247,N_18750);
xor U20120 (N_20120,N_17578,N_19081);
and U20121 (N_20121,N_18191,N_18733);
nand U20122 (N_20122,N_18280,N_18516);
xnor U20123 (N_20123,N_17607,N_19549);
nor U20124 (N_20124,N_17736,N_18386);
nand U20125 (N_20125,N_19829,N_19582);
and U20126 (N_20126,N_18445,N_19432);
nor U20127 (N_20127,N_19079,N_19716);
nand U20128 (N_20128,N_18099,N_18648);
xnor U20129 (N_20129,N_19658,N_19265);
or U20130 (N_20130,N_19735,N_17859);
nor U20131 (N_20131,N_18362,N_18088);
or U20132 (N_20132,N_19973,N_18526);
nand U20133 (N_20133,N_19355,N_19774);
and U20134 (N_20134,N_19909,N_17781);
xnor U20135 (N_20135,N_17668,N_18598);
nor U20136 (N_20136,N_19071,N_18723);
nor U20137 (N_20137,N_18091,N_17778);
and U20138 (N_20138,N_19645,N_19142);
nor U20139 (N_20139,N_18071,N_18054);
nor U20140 (N_20140,N_18111,N_18756);
xor U20141 (N_20141,N_19984,N_18356);
and U20142 (N_20142,N_17680,N_19604);
nand U20143 (N_20143,N_18729,N_19104);
nor U20144 (N_20144,N_18699,N_19178);
xor U20145 (N_20145,N_19443,N_19620);
xor U20146 (N_20146,N_19192,N_19701);
nand U20147 (N_20147,N_19136,N_17621);
xor U20148 (N_20148,N_18413,N_19531);
nand U20149 (N_20149,N_18748,N_19840);
and U20150 (N_20150,N_18998,N_18254);
and U20151 (N_20151,N_19449,N_19556);
nand U20152 (N_20152,N_19341,N_18822);
or U20153 (N_20153,N_18686,N_19962);
xnor U20154 (N_20154,N_18707,N_19697);
and U20155 (N_20155,N_17752,N_18231);
nor U20156 (N_20156,N_17877,N_19475);
and U20157 (N_20157,N_19343,N_17655);
or U20158 (N_20158,N_19030,N_19170);
nand U20159 (N_20159,N_18522,N_19162);
nor U20160 (N_20160,N_19413,N_17692);
xor U20161 (N_20161,N_19311,N_19405);
nand U20162 (N_20162,N_18041,N_19631);
or U20163 (N_20163,N_19010,N_17847);
or U20164 (N_20164,N_17996,N_18379);
and U20165 (N_20165,N_18856,N_19954);
nand U20166 (N_20166,N_17845,N_18754);
xnor U20167 (N_20167,N_17721,N_18291);
and U20168 (N_20168,N_19476,N_19644);
nand U20169 (N_20169,N_19074,N_19525);
or U20170 (N_20170,N_17914,N_19374);
xor U20171 (N_20171,N_17627,N_19898);
nor U20172 (N_20172,N_19916,N_18187);
nor U20173 (N_20173,N_18121,N_17753);
or U20174 (N_20174,N_18227,N_19526);
xnor U20175 (N_20175,N_18825,N_18601);
nand U20176 (N_20176,N_18836,N_17746);
nand U20177 (N_20177,N_18923,N_18044);
and U20178 (N_20178,N_19087,N_19481);
nand U20179 (N_20179,N_18534,N_18252);
nand U20180 (N_20180,N_18486,N_18029);
and U20181 (N_20181,N_17739,N_19072);
or U20182 (N_20182,N_18349,N_18632);
nand U20183 (N_20183,N_19302,N_17701);
xnor U20184 (N_20184,N_17614,N_18642);
xor U20185 (N_20185,N_18020,N_17968);
or U20186 (N_20186,N_17970,N_17694);
and U20187 (N_20187,N_19656,N_18385);
nor U20188 (N_20188,N_17923,N_17814);
xnor U20189 (N_20189,N_19654,N_19031);
and U20190 (N_20190,N_19940,N_18689);
nand U20191 (N_20191,N_19465,N_18446);
xor U20192 (N_20192,N_19507,N_19667);
nand U20193 (N_20193,N_17888,N_19987);
nand U20194 (N_20194,N_18541,N_18725);
xnor U20195 (N_20195,N_19267,N_17515);
or U20196 (N_20196,N_17600,N_18232);
or U20197 (N_20197,N_18899,N_19005);
and U20198 (N_20198,N_19849,N_18691);
or U20199 (N_20199,N_17619,N_18996);
xor U20200 (N_20200,N_18838,N_19417);
or U20201 (N_20201,N_19918,N_19632);
and U20202 (N_20202,N_19590,N_18563);
nand U20203 (N_20203,N_18416,N_17679);
and U20204 (N_20204,N_19562,N_19240);
and U20205 (N_20205,N_19863,N_17560);
nor U20206 (N_20206,N_18087,N_17798);
xor U20207 (N_20207,N_18673,N_19287);
xor U20208 (N_20208,N_17842,N_17744);
nor U20209 (N_20209,N_19874,N_18311);
and U20210 (N_20210,N_17556,N_19926);
nor U20211 (N_20211,N_19822,N_18834);
nand U20212 (N_20212,N_19943,N_17551);
and U20213 (N_20213,N_18764,N_17535);
and U20214 (N_20214,N_18014,N_18657);
nand U20215 (N_20215,N_18558,N_18709);
nor U20216 (N_20216,N_19583,N_19494);
xnor U20217 (N_20217,N_19278,N_18982);
xnor U20218 (N_20218,N_18901,N_18464);
or U20219 (N_20219,N_17543,N_18716);
nor U20220 (N_20220,N_19720,N_17579);
xor U20221 (N_20221,N_17999,N_18637);
nor U20222 (N_20222,N_17916,N_17605);
or U20223 (N_20223,N_18907,N_17972);
nor U20224 (N_20224,N_18656,N_19502);
nor U20225 (N_20225,N_18467,N_19004);
or U20226 (N_20226,N_18779,N_18501);
nand U20227 (N_20227,N_17566,N_18158);
nor U20228 (N_20228,N_17756,N_19368);
nand U20229 (N_20229,N_18867,N_19824);
xnor U20230 (N_20230,N_19778,N_19770);
nand U20231 (N_20231,N_17760,N_17597);
nand U20232 (N_20232,N_18316,N_17506);
and U20233 (N_20233,N_19817,N_19133);
xnor U20234 (N_20234,N_18908,N_18175);
nor U20235 (N_20235,N_18393,N_19749);
nand U20236 (N_20236,N_18207,N_18028);
xnor U20237 (N_20237,N_18995,N_18555);
or U20238 (N_20238,N_19633,N_18573);
or U20239 (N_20239,N_17861,N_19304);
or U20240 (N_20240,N_18814,N_18668);
nand U20241 (N_20241,N_19864,N_18425);
and U20242 (N_20242,N_18329,N_18314);
and U20243 (N_20243,N_18935,N_18595);
and U20244 (N_20244,N_18337,N_18375);
xor U20245 (N_20245,N_18564,N_19796);
or U20246 (N_20246,N_19239,N_18552);
xor U20247 (N_20247,N_18698,N_17673);
or U20248 (N_20248,N_18036,N_17735);
or U20249 (N_20249,N_18104,N_18447);
xor U20250 (N_20250,N_19691,N_17706);
nor U20251 (N_20251,N_19389,N_17674);
nor U20252 (N_20252,N_19485,N_17624);
and U20253 (N_20253,N_18902,N_18131);
xor U20254 (N_20254,N_17553,N_17856);
or U20255 (N_20255,N_18947,N_17704);
xor U20256 (N_20256,N_18897,N_18710);
xnor U20257 (N_20257,N_18489,N_19668);
nor U20258 (N_20258,N_18139,N_18497);
or U20259 (N_20259,N_18061,N_19319);
or U20260 (N_20260,N_19811,N_19313);
or U20261 (N_20261,N_19140,N_18620);
xnor U20262 (N_20262,N_19991,N_19263);
nand U20263 (N_20263,N_18218,N_19600);
or U20264 (N_20264,N_19513,N_18868);
or U20265 (N_20265,N_17832,N_19186);
nor U20266 (N_20266,N_19312,N_19804);
nor U20267 (N_20267,N_18453,N_18205);
xor U20268 (N_20268,N_18883,N_19361);
nand U20269 (N_20269,N_18060,N_19297);
and U20270 (N_20270,N_18410,N_18211);
xor U20271 (N_20271,N_19090,N_18336);
xor U20272 (N_20272,N_18742,N_18571);
nand U20273 (N_20273,N_18735,N_18796);
nand U20274 (N_20274,N_17945,N_18565);
nand U20275 (N_20275,N_19555,N_18313);
or U20276 (N_20276,N_17745,N_19096);
or U20277 (N_20277,N_18070,N_18543);
or U20278 (N_20278,N_18357,N_18859);
or U20279 (N_20279,N_18891,N_18325);
or U20280 (N_20280,N_18593,N_18266);
nor U20281 (N_20281,N_18592,N_19345);
and U20282 (N_20282,N_17880,N_19646);
or U20283 (N_20283,N_18059,N_18046);
nor U20284 (N_20284,N_19295,N_18661);
or U20285 (N_20285,N_17711,N_18638);
nor U20286 (N_20286,N_18370,N_17631);
xnor U20287 (N_20287,N_18879,N_19611);
or U20288 (N_20288,N_18793,N_19381);
nand U20289 (N_20289,N_19179,N_19856);
xnor U20290 (N_20290,N_18458,N_19091);
nor U20291 (N_20291,N_19773,N_19949);
nand U20292 (N_20292,N_18816,N_18161);
nand U20293 (N_20293,N_18392,N_17791);
xor U20294 (N_20294,N_19441,N_17659);
or U20295 (N_20295,N_19342,N_18738);
nor U20296 (N_20296,N_18098,N_18505);
nor U20297 (N_20297,N_19928,N_17713);
nand U20298 (N_20298,N_19883,N_19365);
xor U20299 (N_20299,N_17653,N_18346);
or U20300 (N_20300,N_18442,N_18465);
nor U20301 (N_20301,N_19628,N_17536);
or U20302 (N_20302,N_19805,N_17849);
xnor U20303 (N_20303,N_19205,N_17795);
xor U20304 (N_20304,N_19333,N_19043);
xor U20305 (N_20305,N_18631,N_18524);
and U20306 (N_20306,N_17656,N_18212);
or U20307 (N_20307,N_19666,N_17748);
or U20308 (N_20308,N_18096,N_18499);
nand U20309 (N_20309,N_18845,N_19147);
nand U20310 (N_20310,N_19948,N_18075);
and U20311 (N_20311,N_19438,N_18310);
xnor U20312 (N_20312,N_19388,N_18240);
nand U20313 (N_20313,N_18702,N_18767);
nor U20314 (N_20314,N_18052,N_19873);
or U20315 (N_20315,N_19236,N_19581);
nor U20316 (N_20316,N_19414,N_19218);
or U20317 (N_20317,N_19634,N_17629);
nor U20318 (N_20318,N_19938,N_17797);
xor U20319 (N_20319,N_18230,N_19842);
or U20320 (N_20320,N_18797,N_19651);
nand U20321 (N_20321,N_18123,N_19690);
xor U20322 (N_20322,N_18269,N_18084);
xnor U20323 (N_20323,N_19956,N_18679);
xor U20324 (N_20324,N_18114,N_18688);
and U20325 (N_20325,N_19857,N_17723);
nor U20326 (N_20326,N_17998,N_19976);
and U20327 (N_20327,N_19925,N_18630);
and U20328 (N_20328,N_17890,N_17718);
and U20329 (N_20329,N_19885,N_17574);
nand U20330 (N_20330,N_18484,N_18922);
nand U20331 (N_20331,N_17691,N_19225);
nand U20332 (N_20332,N_19895,N_17689);
xor U20333 (N_20333,N_19370,N_18561);
and U20334 (N_20334,N_18643,N_18426);
or U20335 (N_20335,N_19718,N_19887);
nor U20336 (N_20336,N_18611,N_17869);
or U20337 (N_20337,N_18628,N_17643);
or U20338 (N_20338,N_19870,N_18951);
nand U20339 (N_20339,N_18250,N_19093);
and U20340 (N_20340,N_17805,N_17858);
xor U20341 (N_20341,N_18435,N_19586);
and U20342 (N_20342,N_19964,N_19145);
nand U20343 (N_20343,N_19950,N_19636);
nand U20344 (N_20344,N_19195,N_17505);
and U20345 (N_20345,N_18335,N_19216);
nand U20346 (N_20346,N_19695,N_17808);
xor U20347 (N_20347,N_18423,N_17918);
nor U20348 (N_20348,N_17826,N_18170);
and U20349 (N_20349,N_18390,N_19396);
nor U20350 (N_20350,N_19700,N_17725);
xor U20351 (N_20351,N_18896,N_19635);
nor U20352 (N_20352,N_18333,N_17940);
nand U20353 (N_20353,N_19906,N_17944);
nand U20354 (N_20354,N_19784,N_19164);
and U20355 (N_20355,N_17635,N_19942);
xor U20356 (N_20356,N_17820,N_17520);
xor U20357 (N_20357,N_18430,N_19983);
xnor U20358 (N_20358,N_19440,N_17702);
xor U20359 (N_20359,N_18406,N_19120);
nor U20360 (N_20360,N_18961,N_18140);
nor U20361 (N_20361,N_18461,N_18606);
nand U20362 (N_20362,N_18011,N_19613);
xor U20363 (N_20363,N_19569,N_19233);
or U20364 (N_20364,N_19436,N_19614);
nor U20365 (N_20365,N_19273,N_19467);
or U20366 (N_20366,N_19017,N_17555);
and U20367 (N_20367,N_18929,N_18490);
xor U20368 (N_20368,N_18815,N_18627);
nand U20369 (N_20369,N_19809,N_19944);
xor U20370 (N_20370,N_17874,N_19534);
or U20371 (N_20371,N_17722,N_19532);
and U20372 (N_20372,N_17978,N_19522);
nand U20373 (N_20373,N_19982,N_19011);
or U20374 (N_20374,N_17942,N_19673);
nor U20375 (N_20375,N_17591,N_17765);
and U20376 (N_20376,N_18302,N_19308);
nor U20377 (N_20377,N_19194,N_19994);
and U20378 (N_20378,N_17909,N_19281);
or U20379 (N_20379,N_17603,N_17740);
or U20380 (N_20380,N_18705,N_19722);
and U20381 (N_20381,N_19336,N_19223);
nand U20382 (N_20382,N_19627,N_19913);
nand U20383 (N_20383,N_18214,N_19903);
xnor U20384 (N_20384,N_18235,N_18460);
nand U20385 (N_20385,N_19758,N_18033);
xor U20386 (N_20386,N_18342,N_19769);
nor U20387 (N_20387,N_18529,N_18910);
xnor U20388 (N_20388,N_19128,N_18696);
nor U20389 (N_20389,N_19830,N_18024);
nor U20390 (N_20390,N_19785,N_17962);
or U20391 (N_20391,N_18568,N_18801);
and U20392 (N_20392,N_19026,N_17893);
or U20393 (N_20393,N_18437,N_17608);
xnor U20394 (N_20394,N_17786,N_18136);
and U20395 (N_20395,N_18219,N_17836);
or U20396 (N_20396,N_19439,N_19789);
xor U20397 (N_20397,N_18527,N_18719);
nand U20398 (N_20398,N_19241,N_19053);
nand U20399 (N_20399,N_17626,N_18157);
nor U20400 (N_20400,N_19733,N_17911);
nor U20401 (N_20401,N_19781,N_18126);
nor U20402 (N_20402,N_18520,N_18596);
nand U20403 (N_20403,N_18636,N_19032);
and U20404 (N_20404,N_18206,N_18993);
nand U20405 (N_20405,N_19109,N_18297);
nor U20406 (N_20406,N_19571,N_17754);
and U20407 (N_20407,N_18428,N_18894);
or U20408 (N_20408,N_17552,N_18286);
xnor U20409 (N_20409,N_17686,N_19480);
and U20410 (N_20410,N_17640,N_18690);
or U20411 (N_20411,N_18659,N_17710);
nor U20412 (N_20412,N_17601,N_18517);
nand U20413 (N_20413,N_18197,N_18188);
xor U20414 (N_20414,N_18456,N_17810);
nand U20415 (N_20415,N_19825,N_18889);
nor U20416 (N_20416,N_19082,N_18770);
xnor U20417 (N_20417,N_18234,N_19892);
nand U20418 (N_20418,N_17670,N_18492);
and U20419 (N_20419,N_18132,N_17677);
xor U20420 (N_20420,N_18693,N_19001);
or U20421 (N_20421,N_18479,N_19981);
or U20422 (N_20422,N_18348,N_18293);
xnor U20423 (N_20423,N_19828,N_17539);
nor U20424 (N_20424,N_17696,N_17866);
nand U20425 (N_20425,N_19554,N_19196);
nor U20426 (N_20426,N_18722,N_18339);
and U20427 (N_20427,N_19726,N_18391);
or U20428 (N_20428,N_18967,N_19854);
xor U20429 (N_20429,N_18713,N_19208);
xor U20430 (N_20430,N_19166,N_18806);
xnor U20431 (N_20431,N_19129,N_19334);
nor U20432 (N_20432,N_18583,N_17850);
or U20433 (N_20433,N_17665,N_17796);
nor U20434 (N_20434,N_17546,N_18537);
xnor U20435 (N_20435,N_19957,N_17525);
nand U20436 (N_20436,N_19843,N_18704);
nand U20437 (N_20437,N_18554,N_19966);
or U20438 (N_20438,N_19738,N_18560);
xnor U20439 (N_20439,N_18545,N_18354);
or U20440 (N_20440,N_19056,N_17953);
and U20441 (N_20441,N_19754,N_19296);
xnor U20442 (N_20442,N_18535,N_17898);
or U20443 (N_20443,N_19533,N_18684);
or U20444 (N_20444,N_18790,N_17799);
nor U20445 (N_20445,N_18575,N_18288);
or U20446 (N_20446,N_17868,N_19114);
or U20447 (N_20447,N_19224,N_19034);
or U20448 (N_20448,N_18201,N_19585);
and U20449 (N_20449,N_18222,N_17774);
nor U20450 (N_20450,N_19776,N_18378);
nor U20451 (N_20451,N_18546,N_18022);
nand U20452 (N_20452,N_17862,N_17606);
xor U20453 (N_20453,N_18768,N_19434);
nor U20454 (N_20454,N_17632,N_17707);
xor U20455 (N_20455,N_18411,N_17975);
and U20456 (N_20456,N_19605,N_17699);
nor U20457 (N_20457,N_19577,N_17573);
or U20458 (N_20458,N_19860,N_19687);
nand U20459 (N_20459,N_19524,N_17676);
and U20460 (N_20460,N_18507,N_17612);
and U20461 (N_20461,N_19491,N_19403);
and U20462 (N_20462,N_18414,N_19177);
nor U20463 (N_20463,N_18213,N_18292);
nand U20464 (N_20464,N_17887,N_18275);
nor U20465 (N_20465,N_18892,N_18371);
nor U20466 (N_20466,N_18352,N_19535);
or U20467 (N_20467,N_18652,N_17848);
xor U20468 (N_20468,N_17986,N_19702);
nor U20469 (N_20469,N_19648,N_19219);
nor U20470 (N_20470,N_19521,N_19222);
or U20471 (N_20471,N_19573,N_17681);
nand U20472 (N_20472,N_18299,N_18736);
and U20473 (N_20473,N_19430,N_19268);
xor U20474 (N_20474,N_18116,N_19550);
nor U20475 (N_20475,N_19807,N_18759);
xnor U20476 (N_20476,N_19252,N_19841);
nand U20477 (N_20477,N_17568,N_18076);
xnor U20478 (N_20478,N_17819,N_19169);
xnor U20479 (N_20479,N_18672,N_18369);
nand U20480 (N_20480,N_18938,N_17860);
nor U20481 (N_20481,N_19039,N_19641);
or U20482 (N_20482,N_18994,N_19454);
or U20483 (N_20483,N_17709,N_18513);
xnor U20484 (N_20484,N_18270,N_19902);
or U20485 (N_20485,N_18703,N_18451);
nor U20486 (N_20486,N_19915,N_19068);
nand U20487 (N_20487,N_18849,N_18805);
nand U20488 (N_20488,N_19286,N_19327);
nand U20489 (N_20489,N_18331,N_19352);
nand U20490 (N_20490,N_17875,N_19346);
and U20491 (N_20491,N_17766,N_19952);
or U20492 (N_20492,N_19595,N_18477);
nor U20493 (N_20493,N_18242,N_18482);
nand U20494 (N_20494,N_17751,N_18918);
and U20495 (N_20495,N_17895,N_18962);
nor U20496 (N_20496,N_18068,N_17941);
and U20497 (N_20497,N_19411,N_18256);
nand U20498 (N_20498,N_19515,N_19699);
and U20499 (N_20499,N_19881,N_17728);
nand U20500 (N_20500,N_19041,N_19706);
or U20501 (N_20501,N_19941,N_18326);
xor U20502 (N_20502,N_19493,N_19775);
xor U20503 (N_20503,N_19558,N_17800);
and U20504 (N_20504,N_19126,N_17789);
or U20505 (N_20505,N_19423,N_19642);
xor U20506 (N_20506,N_18566,N_19246);
xor U20507 (N_20507,N_18309,N_18972);
nor U20508 (N_20508,N_17533,N_18058);
nand U20509 (N_20509,N_17851,N_18419);
and U20510 (N_20510,N_18556,N_18980);
and U20511 (N_20511,N_18559,N_18347);
and U20512 (N_20512,N_18400,N_18973);
and U20513 (N_20513,N_18666,N_17987);
and U20514 (N_20514,N_18876,N_19047);
xor U20515 (N_20515,N_19002,N_17717);
xor U20516 (N_20516,N_18574,N_17572);
xor U20517 (N_20517,N_19061,N_17811);
nor U20518 (N_20518,N_19894,N_19693);
nand U20519 (N_20519,N_19564,N_18404);
nand U20520 (N_20520,N_17864,N_17779);
or U20521 (N_20521,N_18843,N_19335);
nor U20522 (N_20522,N_19134,N_19901);
nor U20523 (N_20523,N_19839,N_17886);
and U20524 (N_20524,N_17682,N_19251);
or U20525 (N_20525,N_19649,N_19269);
nor U20526 (N_20526,N_17963,N_18787);
nor U20527 (N_20527,N_17687,N_19123);
xnor U20528 (N_20528,N_18757,N_17943);
nor U20529 (N_20529,N_19108,N_19477);
nand U20530 (N_20530,N_17645,N_17825);
xnor U20531 (N_20531,N_18683,N_19567);
nand U20532 (N_20532,N_17788,N_18015);
and U20533 (N_20533,N_19827,N_19152);
nor U20534 (N_20534,N_19202,N_18609);
xnor U20535 (N_20535,N_19029,N_18579);
nor U20536 (N_20536,N_17813,N_19993);
xor U20537 (N_20537,N_19459,N_17995);
nor U20538 (N_20538,N_18457,N_17598);
or U20539 (N_20539,N_18312,N_19528);
nand U20540 (N_20540,N_19922,N_19350);
nor U20541 (N_20541,N_19408,N_19392);
and U20542 (N_20542,N_17542,N_19783);
xor U20543 (N_20543,N_19538,N_19727);
nand U20544 (N_20544,N_17537,N_19988);
xnor U20545 (N_20545,N_18605,N_19509);
nand U20546 (N_20546,N_19121,N_18093);
xor U20547 (N_20547,N_18480,N_18956);
nand U20548 (N_20548,N_19848,N_17654);
nor U20549 (N_20549,N_19739,N_17716);
xnor U20550 (N_20550,N_19998,N_19933);
nor U20551 (N_20551,N_19763,N_19969);
nand U20552 (N_20552,N_19360,N_18997);
xor U20553 (N_20553,N_17990,N_19529);
or U20554 (N_20554,N_19371,N_18200);
or U20555 (N_20555,N_17732,N_18043);
xnor U20556 (N_20556,N_18162,N_19316);
nand U20557 (N_20557,N_17917,N_19974);
xor U20558 (N_20558,N_18338,N_17749);
xnor U20559 (N_20559,N_19955,N_19207);
or U20560 (N_20560,N_18008,N_17641);
nor U20561 (N_20561,N_18650,N_18622);
nand U20562 (N_20562,N_19801,N_19230);
or U20563 (N_20563,N_19959,N_17514);
or U20564 (N_20564,N_18021,N_17526);
or U20565 (N_20565,N_19020,N_19105);
and U20566 (N_20566,N_19622,N_18773);
nand U20567 (N_20567,N_19100,N_18921);
nor U20568 (N_20568,N_19871,N_17639);
xnor U20569 (N_20569,N_18042,N_17913);
or U20570 (N_20570,N_18117,N_18730);
nor U20571 (N_20571,N_17742,N_17531);
nor U20572 (N_20572,N_19888,N_18882);
nor U20573 (N_20573,N_19158,N_18133);
nor U20574 (N_20574,N_18548,N_18999);
and U20575 (N_20575,N_17652,N_17884);
nand U20576 (N_20576,N_17666,N_18100);
and U20577 (N_20577,N_19665,N_19175);
nand U20578 (N_20578,N_19536,N_18557);
nor U20579 (N_20579,N_18888,N_17928);
xnor U20580 (N_20580,N_18937,N_19492);
xor U20581 (N_20581,N_17946,N_18209);
nand U20582 (N_20582,N_19624,N_17609);
and U20583 (N_20583,N_19852,N_19171);
and U20584 (N_20584,N_19908,N_19989);
nor U20585 (N_20585,N_18824,N_18259);
nor U20586 (N_20586,N_19652,N_19946);
or U20587 (N_20587,N_18491,N_18813);
nor U20588 (N_20588,N_18645,N_17823);
and U20589 (N_20589,N_18472,N_18909);
nor U20590 (N_20590,N_18173,N_18726);
nor U20591 (N_20591,N_19975,N_19422);
or U20592 (N_20592,N_17554,N_17981);
or U20593 (N_20593,N_18984,N_17519);
nor U20594 (N_20594,N_17758,N_17839);
nand U20595 (N_20595,N_19596,N_19189);
or U20596 (N_20596,N_18229,N_17853);
nor U20597 (N_20597,N_17910,N_18306);
xnor U20598 (N_20598,N_17507,N_18613);
nand U20599 (N_20599,N_19650,N_18495);
and U20600 (N_20600,N_18992,N_18057);
xor U20601 (N_20601,N_19356,N_17693);
nor U20602 (N_20602,N_19782,N_18865);
or U20603 (N_20603,N_17615,N_19679);
or U20604 (N_20604,N_19711,N_18160);
xor U20605 (N_20605,N_18496,N_18189);
nor U20606 (N_20606,N_18939,N_19328);
or U20607 (N_20607,N_17571,N_18744);
xnor U20608 (N_20608,N_18268,N_18974);
nor U20609 (N_20609,N_19643,N_19141);
nand U20610 (N_20610,N_18468,N_18025);
and U20611 (N_20611,N_18124,N_19505);
xnor U20612 (N_20612,N_19244,N_18128);
xor U20613 (N_20613,N_18086,N_19073);
xor U20614 (N_20614,N_18176,N_19972);
xor U20615 (N_20615,N_19415,N_18818);
nand U20616 (N_20616,N_18819,N_19463);
nand U20617 (N_20617,N_19275,N_18635);
xnor U20618 (N_20618,N_18741,N_19248);
xnor U20619 (N_20619,N_18590,N_17529);
nand U20620 (N_20620,N_19905,N_18409);
xnor U20621 (N_20621,N_17871,N_18353);
xor U20622 (N_20622,N_19845,N_18862);
nand U20623 (N_20623,N_17785,N_18066);
nand U20624 (N_20624,N_19619,N_19914);
nand U20625 (N_20625,N_19394,N_18577);
or U20626 (N_20626,N_18978,N_18092);
nor U20627 (N_20627,N_19021,N_18586);
xor U20628 (N_20628,N_19174,N_19539);
or U20629 (N_20629,N_19968,N_17806);
nand U20630 (N_20630,N_18789,N_19182);
xor U20631 (N_20631,N_17741,N_18263);
nand U20632 (N_20632,N_17530,N_18665);
nor U20633 (N_20633,N_17977,N_19187);
or U20634 (N_20634,N_18454,N_17782);
or U20635 (N_20635,N_19055,N_19036);
xnor U20636 (N_20636,N_17865,N_19457);
xnor U20637 (N_20637,N_17802,N_19024);
nor U20638 (N_20638,N_18307,N_17617);
nand U20639 (N_20639,N_18243,N_17584);
and U20640 (N_20640,N_18835,N_17637);
and U20641 (N_20641,N_17931,N_17618);
xnor U20642 (N_20642,N_18224,N_19324);
nand U20643 (N_20643,N_18752,N_18144);
nand U20644 (N_20644,N_17570,N_18853);
or U20645 (N_20645,N_18463,N_19510);
and U20646 (N_20646,N_19173,N_18917);
nor U20647 (N_20647,N_18179,N_18504);
xor U20648 (N_20648,N_17583,N_19800);
and U20649 (N_20649,N_18448,N_18708);
and U20650 (N_20650,N_19897,N_17590);
nand U20651 (N_20651,N_19469,N_18035);
xor U20652 (N_20652,N_19965,N_19929);
or U20653 (N_20653,N_19387,N_18957);
nor U20654 (N_20654,N_18225,N_18199);
nand U20655 (N_20655,N_17545,N_19331);
and U20656 (N_20656,N_19663,N_18360);
and U20657 (N_20657,N_19402,N_19728);
or U20658 (N_20658,N_17771,N_19682);
nand U20659 (N_20659,N_19877,N_19788);
and U20660 (N_20660,N_19285,N_18544);
nor U20661 (N_20661,N_18784,N_19318);
and U20662 (N_20662,N_19732,N_18315);
nand U20663 (N_20663,N_17727,N_18807);
and U20664 (N_20664,N_19437,N_18125);
xnor U20665 (N_20665,N_18023,N_19391);
and U20666 (N_20666,N_18380,N_19756);
nor U20667 (N_20667,N_19198,N_19506);
xor U20668 (N_20668,N_19837,N_17611);
or U20669 (N_20669,N_18264,N_18968);
nor U20670 (N_20670,N_18134,N_18949);
nand U20671 (N_20671,N_18049,N_18459);
or U20672 (N_20672,N_18389,N_17780);
and U20673 (N_20673,N_19471,N_17500);
nor U20674 (N_20674,N_17902,N_17870);
xnor U20675 (N_20675,N_18296,N_18478);
or U20676 (N_20676,N_17518,N_17969);
nor U20677 (N_20677,N_17638,N_18498);
xnor U20678 (N_20678,N_17883,N_19717);
nand U20679 (N_20679,N_17528,N_18159);
nor U20680 (N_20680,N_17538,N_17956);
xnor U20681 (N_20681,N_18562,N_18438);
or U20682 (N_20682,N_19373,N_18402);
nor U20683 (N_20683,N_19745,N_19653);
nand U20684 (N_20684,N_18576,N_19676);
xnor U20685 (N_20685,N_19803,N_19270);
nor U20686 (N_20686,N_18530,N_18983);
or U20687 (N_20687,N_17991,N_18233);
or U20688 (N_20688,N_18415,N_19985);
nor U20689 (N_20689,N_19380,N_18137);
or U20690 (N_20690,N_19713,N_18639);
xnor U20691 (N_20691,N_19566,N_18599);
or U20692 (N_20692,N_18149,N_19671);
xor U20693 (N_20693,N_17548,N_19719);
nand U20694 (N_20694,N_18852,N_19802);
or U20695 (N_20695,N_18261,N_17575);
or U20696 (N_20696,N_19570,N_18283);
xnor U20697 (N_20697,N_18662,N_18321);
nor U20698 (N_20698,N_18749,N_19226);
and U20699 (N_20699,N_18327,N_19199);
nand U20700 (N_20700,N_17937,N_19548);
xor U20701 (N_20701,N_17715,N_17667);
nand U20702 (N_20702,N_18067,N_18500);
or U20703 (N_20703,N_17983,N_19855);
and U20704 (N_20704,N_19704,N_17793);
and U20705 (N_20705,N_18532,N_19579);
or U20706 (N_20706,N_17958,N_19125);
or U20707 (N_20707,N_19271,N_18097);
and U20708 (N_20708,N_18271,N_19615);
xor U20709 (N_20709,N_19953,N_19869);
nor U20710 (N_20710,N_17675,N_17559);
and U20711 (N_20711,N_17510,N_19022);
and U20712 (N_20712,N_19088,N_19705);
and U20713 (N_20713,N_18195,N_19503);
nor U20714 (N_20714,N_18919,N_18169);
and U20715 (N_20715,N_19958,N_19250);
or U20716 (N_20716,N_18864,N_17830);
or U20717 (N_20717,N_18528,N_18511);
and U20718 (N_20718,N_18640,N_18146);
or U20719 (N_20719,N_18506,N_18963);
nand U20720 (N_20720,N_17834,N_18065);
nand U20721 (N_20721,N_19818,N_18226);
nand U20722 (N_20722,N_18077,N_19468);
or U20723 (N_20723,N_18475,N_18829);
xnor U20724 (N_20724,N_17719,N_18069);
and U20725 (N_20725,N_19618,N_18215);
or U20726 (N_20726,N_17540,N_19066);
or U20727 (N_20727,N_19686,N_17894);
xnor U20728 (N_20728,N_17762,N_18948);
nand U20729 (N_20729,N_19366,N_18017);
and U20730 (N_20730,N_18920,N_17669);
nor U20731 (N_20731,N_19089,N_18578);
and U20732 (N_20732,N_18653,N_18078);
nor U20733 (N_20733,N_19594,N_19675);
nand U20734 (N_20734,N_18005,N_19878);
nor U20735 (N_20735,N_19113,N_19237);
xor U20736 (N_20736,N_18514,N_18322);
and U20737 (N_20737,N_18536,N_18090);
xnor U20738 (N_20738,N_19689,N_18018);
xor U20739 (N_20739,N_17541,N_18323);
nand U20740 (N_20740,N_19541,N_18990);
or U20741 (N_20741,N_19144,N_19919);
nor U20742 (N_20742,N_17900,N_19747);
or U20743 (N_20743,N_17967,N_18050);
xnor U20744 (N_20744,N_18775,N_19447);
or U20745 (N_20745,N_19132,N_19301);
nor U20746 (N_20746,N_19050,N_19630);
or U20747 (N_20747,N_19112,N_18614);
or U20748 (N_20748,N_19574,N_19084);
or U20749 (N_20749,N_17863,N_18798);
xor U20750 (N_20750,N_19213,N_18711);
nand U20751 (N_20751,N_18600,N_19262);
and U20752 (N_20752,N_19730,N_17891);
or U20753 (N_20753,N_17938,N_19347);
and U20754 (N_20754,N_17777,N_19847);
nor U20755 (N_20755,N_19409,N_19487);
or U20756 (N_20756,N_19461,N_19460);
or U20757 (N_20757,N_17948,N_18359);
or U20758 (N_20758,N_19910,N_19337);
or U20759 (N_20759,N_17596,N_18772);
nor U20760 (N_20760,N_18685,N_18663);
or U20761 (N_20761,N_17783,N_19322);
nand U20762 (N_20762,N_19462,N_18837);
or U20763 (N_20763,N_17955,N_19978);
or U20764 (N_20764,N_19846,N_18734);
nand U20765 (N_20765,N_19063,N_17838);
and U20766 (N_20766,N_17922,N_19217);
nor U20767 (N_20767,N_19424,N_18223);
nor U20768 (N_20768,N_18130,N_18930);
xnor U20769 (N_20769,N_18427,N_19891);
nor U20770 (N_20770,N_18502,N_18318);
nand U20771 (N_20771,N_18924,N_18481);
nand U20772 (N_20772,N_19464,N_19793);
nor U20773 (N_20773,N_18553,N_18869);
nor U20774 (N_20774,N_19122,N_17664);
nor U20775 (N_20775,N_19235,N_19359);
and U20776 (N_20776,N_19694,N_18680);
and U20777 (N_20777,N_19234,N_19393);
nand U20778 (N_20778,N_18249,N_17602);
nor U20779 (N_20779,N_18246,N_19734);
or U20780 (N_20780,N_19329,N_18279);
xor U20781 (N_20781,N_18981,N_19766);
xnor U20782 (N_20782,N_18625,N_17757);
and U20783 (N_20783,N_18202,N_19736);
nand U20784 (N_20784,N_19692,N_18424);
nand U20785 (N_20785,N_18580,N_17521);
xor U20786 (N_20786,N_18452,N_17794);
or U20787 (N_20787,N_18760,N_19703);
or U20788 (N_20788,N_18431,N_19920);
nand U20789 (N_20789,N_19591,N_19996);
xor U20790 (N_20790,N_19095,N_17829);
nand U20791 (N_20791,N_18943,N_19298);
nor U20792 (N_20792,N_17831,N_18550);
or U20793 (N_20793,N_17564,N_19815);
nor U20794 (N_20794,N_18687,N_18521);
nand U20795 (N_20795,N_19172,N_19572);
nor U20796 (N_20796,N_19813,N_19452);
nand U20797 (N_20797,N_19354,N_19330);
xnor U20798 (N_20798,N_19741,N_19255);
xor U20799 (N_20799,N_19917,N_19791);
xnor U20800 (N_20800,N_19814,N_19256);
xor U20801 (N_20801,N_19274,N_18792);
or U20802 (N_20802,N_18674,N_19714);
or U20803 (N_20803,N_17982,N_17873);
nor U20804 (N_20804,N_17985,N_17589);
nor U20805 (N_20805,N_19156,N_19077);
nand U20806 (N_20806,N_19779,N_18512);
nor U20807 (N_20807,N_17927,N_19560);
xnor U20808 (N_20808,N_17743,N_18916);
or U20809 (N_20809,N_19623,N_19655);
nand U20810 (N_20810,N_19348,N_18934);
or U20811 (N_20811,N_17828,N_18538);
nor U20812 (N_20812,N_18110,N_18106);
nand U20813 (N_20813,N_19395,N_19015);
or U20814 (N_20814,N_18113,N_18470);
nor U20815 (N_20815,N_18395,N_19587);
xor U20816 (N_20816,N_18945,N_18594);
and U20817 (N_20817,N_17961,N_18063);
xor U20818 (N_20818,N_18875,N_17815);
and U20819 (N_20819,N_18821,N_18572);
or U20820 (N_20820,N_19599,N_18633);
nor U20821 (N_20821,N_17522,N_18154);
or U20822 (N_20822,N_19951,N_17934);
and U20823 (N_20823,N_19442,N_19155);
and U20824 (N_20824,N_18193,N_17974);
or U20825 (N_20825,N_18519,N_19563);
and U20826 (N_20826,N_18651,N_19868);
xor U20827 (N_20827,N_19992,N_18115);
and U20828 (N_20828,N_19637,N_19742);
or U20829 (N_20829,N_19190,N_18989);
and U20830 (N_20830,N_18851,N_18436);
nand U20831 (N_20831,N_19412,N_18163);
nand U20832 (N_20832,N_19119,N_18074);
xor U20833 (N_20833,N_19206,N_19399);
nor U20834 (N_20834,N_19009,N_18547);
or U20835 (N_20835,N_19283,N_17881);
and U20836 (N_20836,N_19889,N_18341);
nand U20837 (N_20837,N_19369,N_18281);
nor U20838 (N_20838,N_17822,N_19488);
nor U20839 (N_20839,N_18731,N_18278);
nand U20840 (N_20840,N_18262,N_18717);
nand U20841 (N_20841,N_17776,N_19882);
or U20842 (N_20842,N_18072,N_19743);
nand U20843 (N_20843,N_19907,N_19661);
nor U20844 (N_20844,N_19003,N_19886);
and U20845 (N_20845,N_19578,N_17663);
nand U20846 (N_20846,N_18493,N_19127);
or U20847 (N_20847,N_18952,N_19986);
nor U20848 (N_20848,N_18081,N_19504);
or U20849 (N_20849,N_17593,N_17912);
nor U20850 (N_20850,N_19138,N_19294);
nor U20851 (N_20851,N_18842,N_19500);
and U20852 (N_20852,N_19698,N_19307);
nor U20853 (N_20853,N_18433,N_19746);
and U20854 (N_20854,N_19191,N_19936);
or U20855 (N_20855,N_18727,N_19771);
nand U20856 (N_20856,N_18398,N_18658);
nand U20857 (N_20857,N_19543,N_18351);
nor U20858 (N_20858,N_19584,N_19518);
nand U20859 (N_20859,N_17988,N_18455);
nand U20860 (N_20860,N_17960,N_17550);
nand U20861 (N_20861,N_18399,N_19150);
nor U20862 (N_20862,N_18245,N_19450);
nor U20863 (N_20863,N_18755,N_18860);
nor U20864 (N_20864,N_18971,N_18870);
nand U20865 (N_20865,N_17688,N_18101);
nand U20866 (N_20866,N_19456,N_19060);
xor U20867 (N_20867,N_18237,N_17976);
or U20868 (N_20868,N_18183,N_18403);
nand U20869 (N_20869,N_19231,N_17708);
nand U20870 (N_20870,N_18604,N_19258);
nand U20871 (N_20871,N_17903,N_18724);
nand U20872 (N_20872,N_19085,N_18364);
or U20873 (N_20873,N_18248,N_19939);
and U20874 (N_20874,N_17622,N_18152);
and U20875 (N_20875,N_19261,N_17821);
nor U20876 (N_20876,N_19851,N_18343);
nor U20877 (N_20877,N_19612,N_19961);
xnor U20878 (N_20878,N_19013,N_19272);
nor U20879 (N_20879,N_19725,N_18771);
xor U20880 (N_20880,N_18244,N_19277);
nor U20881 (N_20881,N_18960,N_18361);
nor U20882 (N_20882,N_17582,N_19924);
and U20883 (N_20883,N_19288,N_18969);
or U20884 (N_20884,N_18129,N_18216);
nand U20885 (N_20885,N_19007,N_18396);
nand U20886 (N_20886,N_17561,N_18107);
or U20887 (N_20887,N_17503,N_19382);
xnor U20888 (N_20888,N_19243,N_17840);
and U20889 (N_20889,N_19744,N_18365);
nand U20890 (N_20890,N_18946,N_19364);
and U20891 (N_20891,N_18839,N_19455);
xor U20892 (N_20892,N_18089,N_19107);
nor U20893 (N_20893,N_18794,N_19406);
and U20894 (N_20894,N_19023,N_18094);
and U20895 (N_20895,N_19157,N_18608);
nand U20896 (N_20896,N_17905,N_19486);
and U20897 (N_20897,N_19511,N_19358);
nor U20898 (N_20898,N_19401,N_17661);
xnor U20899 (N_20899,N_17636,N_17932);
or U20900 (N_20900,N_18324,N_17734);
or U20901 (N_20901,N_17827,N_19780);
xnor U20902 (N_20902,N_18108,N_19398);
nand U20903 (N_20903,N_17733,N_19647);
or U20904 (N_20904,N_17801,N_19816);
or U20905 (N_20905,N_19478,N_18840);
xor U20906 (N_20906,N_19629,N_19537);
xor U20907 (N_20907,N_18165,N_19721);
and U20908 (N_20908,N_19967,N_18150);
nor U20909 (N_20909,N_19935,N_18844);
and U20910 (N_20910,N_19420,N_18148);
and U20911 (N_20911,N_18138,N_18095);
or U20912 (N_20912,N_17750,N_18655);
nand U20913 (N_20913,N_19428,N_19772);
or U20914 (N_20914,N_17833,N_18857);
or U20915 (N_20915,N_19833,N_18795);
nor U20916 (N_20916,N_18985,N_17616);
nand U20917 (N_20917,N_17586,N_18401);
nand U20918 (N_20918,N_18388,N_19340);
or U20919 (N_20919,N_19193,N_17939);
or U20920 (N_20920,N_19786,N_18276);
xor U20921 (N_20921,N_18298,N_19151);
nand U20922 (N_20922,N_17950,N_18282);
nor U20923 (N_20923,N_17837,N_18319);
and U20924 (N_20924,N_19979,N_17897);
nand U20925 (N_20925,N_19075,N_17790);
nor U20926 (N_20926,N_18120,N_19971);
and U20927 (N_20927,N_17906,N_18762);
nor U20928 (N_20928,N_19740,N_18766);
and U20929 (N_20929,N_18407,N_19496);
and U20930 (N_20930,N_19259,N_18373);
and U20931 (N_20931,N_17562,N_19850);
xnor U20932 (N_20932,N_19131,N_18585);
nand U20933 (N_20933,N_19445,N_18700);
xor U20934 (N_20934,N_17577,N_19519);
or U20935 (N_20935,N_19094,N_18285);
nor U20936 (N_20936,N_19552,N_19997);
xor U20937 (N_20937,N_19019,N_18660);
or U20938 (N_20938,N_18471,N_18569);
nand U20939 (N_20939,N_18551,N_19872);
nor U20940 (N_20940,N_19377,N_19254);
nor U20941 (N_20941,N_18142,N_18487);
xnor U20942 (N_20942,N_18190,N_19421);
or U20943 (N_20943,N_19597,N_19310);
or U20944 (N_20944,N_19400,N_18418);
and U20945 (N_20945,N_18809,N_18872);
and U20946 (N_20946,N_19639,N_19076);
nand U20947 (N_20947,N_19070,N_17613);
or U20948 (N_20948,N_17594,N_17775);
or U20949 (N_20949,N_18850,N_18303);
and U20950 (N_20950,N_19372,N_19086);
nand U20951 (N_20951,N_19715,N_19710);
or U20952 (N_20952,N_19242,N_18287);
nor U20953 (N_20953,N_18344,N_18208);
and U20954 (N_20954,N_17511,N_19101);
nor U20955 (N_20955,N_18884,N_17648);
nand U20956 (N_20956,N_17892,N_19832);
xor U20957 (N_20957,N_19609,N_18987);
xnor U20958 (N_20958,N_17567,N_17904);
xor U20959 (N_20959,N_18647,N_18846);
and U20960 (N_20960,N_19000,N_17671);
nand U20961 (N_20961,N_17517,N_19299);
xnor U20962 (N_20962,N_19426,N_18676);
and U20963 (N_20963,N_18681,N_19353);
and U20964 (N_20964,N_18589,N_18172);
nand U20965 (N_20965,N_19937,N_19542);
and U20966 (N_20966,N_19069,N_19712);
xor U20967 (N_20967,N_18367,N_18903);
and U20968 (N_20968,N_19559,N_19067);
nor U20969 (N_20969,N_18450,N_18510);
nand U20970 (N_20970,N_18412,N_19812);
nor U20971 (N_20971,N_19799,N_18429);
xnor U20972 (N_20972,N_19670,N_18182);
nor U20973 (N_20973,N_18290,N_17835);
xnor U20974 (N_20974,N_18944,N_19495);
or U20975 (N_20975,N_17610,N_19520);
nor U20976 (N_20976,N_18488,N_18485);
nand U20977 (N_20977,N_19831,N_17907);
and U20978 (N_20978,N_17620,N_17901);
and U20979 (N_20979,N_18587,N_19204);
or U20980 (N_20980,N_19344,N_19284);
nor U20981 (N_20981,N_19188,N_19238);
xnor U20982 (N_20982,N_19052,N_19448);
nor U20983 (N_20983,N_19279,N_19672);
or U20984 (N_20984,N_18439,N_17885);
or U20985 (N_20985,N_18654,N_18737);
and U20986 (N_20986,N_17993,N_18384);
xor U20987 (N_20987,N_19866,N_18032);
and U20988 (N_20988,N_19451,N_19575);
nand U20989 (N_20989,N_18677,N_18220);
nand U20990 (N_20990,N_18186,N_18925);
and U20991 (N_20991,N_17973,N_17803);
or U20992 (N_20992,N_18013,N_18469);
xnor U20993 (N_20993,N_18462,N_19253);
or U20994 (N_20994,N_17516,N_18026);
nand U20995 (N_20995,N_18847,N_19853);
and U20996 (N_20996,N_18185,N_19390);
nor U20997 (N_20997,N_19764,N_18927);
xnor U20998 (N_20998,N_19220,N_19006);
and U20999 (N_20999,N_18692,N_17852);
xnor U21000 (N_21000,N_18777,N_19546);
and U21001 (N_21001,N_18007,N_18466);
xor U21002 (N_21002,N_19149,N_19367);
or U21003 (N_21003,N_19790,N_17523);
nor U21004 (N_21004,N_17630,N_18194);
xor U21005 (N_21005,N_17899,N_18474);
nand U21006 (N_21006,N_19180,N_17657);
xnor U21007 (N_21007,N_18417,N_18542);
xnor U21008 (N_21008,N_17547,N_18174);
or U21009 (N_21009,N_18047,N_19977);
xnor U21010 (N_21010,N_19309,N_17700);
and U21011 (N_21011,N_18483,N_19203);
and U21012 (N_21012,N_18539,N_18965);
nand U21013 (N_21013,N_19058,N_18027);
and U21014 (N_21014,N_19249,N_19098);
xor U21015 (N_21015,N_18786,N_19490);
and U21016 (N_21016,N_18383,N_18210);
xor U21017 (N_21017,N_19276,N_18911);
nand U21018 (N_21018,N_17642,N_18874);
xnor U21019 (N_21019,N_17683,N_18900);
nand U21020 (N_21020,N_19610,N_19153);
xor U21021 (N_21021,N_17720,N_18881);
nand U21022 (N_21022,N_19470,N_17504);
or U21023 (N_21023,N_18533,N_17957);
xor U21024 (N_21024,N_19048,N_19765);
xor U21025 (N_21025,N_19893,N_19115);
xnor U21026 (N_21026,N_18905,N_18258);
xnor U21027 (N_21027,N_19167,N_19875);
nor U21028 (N_21028,N_19945,N_19970);
xor U21029 (N_21029,N_19482,N_18003);
or U21030 (N_21030,N_18105,N_18616);
xor U21031 (N_21031,N_19135,N_18774);
nand U21032 (N_21032,N_19016,N_19737);
nor U21033 (N_21033,N_19083,N_18217);
nand U21034 (N_21034,N_18799,N_18567);
xor U21035 (N_21035,N_18612,N_18509);
and U21036 (N_21036,N_18038,N_19229);
xnor U21037 (N_21037,N_18817,N_19130);
and U21038 (N_21038,N_19215,N_19092);
nand U21039 (N_21039,N_18010,N_19544);
nor U21040 (N_21040,N_19212,N_19820);
nor U21041 (N_21041,N_18155,N_19681);
xnor U21042 (N_21042,N_17908,N_18828);
xnor U21043 (N_21043,N_17633,N_19458);
nand U21044 (N_21044,N_19357,N_19808);
nand U21045 (N_21045,N_18531,N_18381);
nand U21046 (N_21046,N_18866,N_19363);
nor U21047 (N_21047,N_17763,N_19696);
and U21048 (N_21048,N_17954,N_19685);
or U21049 (N_21049,N_19792,N_18826);
nor U21050 (N_21050,N_17513,N_18841);
and U21051 (N_21051,N_19499,N_17770);
nand U21052 (N_21052,N_19755,N_19589);
nand U21053 (N_21053,N_18503,N_19750);
nor U21054 (N_21054,N_17929,N_19497);
nor U21055 (N_21055,N_18933,N_19580);
or U21056 (N_21056,N_19858,N_19835);
and U21057 (N_21057,N_18886,N_19621);
and U21058 (N_21058,N_18928,N_18602);
nand U21059 (N_21059,N_19674,N_19752);
nand U21060 (N_21060,N_18694,N_19106);
nor U21061 (N_21061,N_17930,N_17921);
nand U21062 (N_21062,N_18334,N_17896);
or U21063 (N_21063,N_19293,N_18085);
and U21064 (N_21064,N_19245,N_18715);
and U21065 (N_21065,N_18394,N_18265);
and U21066 (N_21066,N_19810,N_17690);
xnor U21067 (N_21067,N_18912,N_18753);
nand U21068 (N_21068,N_19797,N_17714);
nor U21069 (N_21069,N_18610,N_18494);
or U21070 (N_21070,N_17824,N_19466);
or U21071 (N_21071,N_18893,N_18718);
and U21072 (N_21072,N_18977,N_17651);
nand U21073 (N_21073,N_18871,N_19282);
and U21074 (N_21074,N_18986,N_17650);
nand U21075 (N_21075,N_18926,N_18366);
or U21076 (N_21076,N_18284,N_19819);
or U21077 (N_21077,N_18272,N_19038);
nor U21078 (N_21078,N_19378,N_18739);
nand U21079 (N_21079,N_19664,N_17966);
or U21080 (N_21080,N_17747,N_19431);
xnor U21081 (N_21081,N_18830,N_18274);
xnor U21082 (N_21082,N_18964,N_19266);
xnor U21083 (N_21083,N_17844,N_19183);
nor U21084 (N_21084,N_18649,N_19660);
nand U21085 (N_21085,N_19823,N_18305);
xor U21086 (N_21086,N_19899,N_17925);
or U21087 (N_21087,N_18783,N_18119);
xnor U21088 (N_21088,N_18854,N_19419);
and U21089 (N_21089,N_19315,N_17697);
nor U21090 (N_21090,N_18294,N_19025);
nand U21091 (N_21091,N_19042,N_18549);
nor U21092 (N_21092,N_19523,N_17544);
nand U21093 (N_21093,N_18540,N_17549);
and U21094 (N_21094,N_19159,N_18603);
or U21095 (N_21095,N_17502,N_17599);
nor U21096 (N_21096,N_18932,N_18135);
or U21097 (N_21097,N_19321,N_17951);
xnor U21098 (N_21098,N_18196,N_17649);
and U21099 (N_21099,N_19638,N_18127);
or U21100 (N_21100,N_18377,N_19777);
nor U21101 (N_21101,N_19753,N_17872);
or U21102 (N_21102,N_18669,N_18936);
and U21103 (N_21103,N_19551,N_19040);
or U21104 (N_21104,N_18171,N_18763);
or U21105 (N_21105,N_18045,N_17729);
or U21106 (N_21106,N_19767,N_17724);
or U21107 (N_21107,N_17994,N_18040);
and U21108 (N_21108,N_19059,N_19397);
nor U21109 (N_21109,N_19512,N_18382);
or U21110 (N_21110,N_17876,N_18203);
nand U21111 (N_21111,N_18820,N_19349);
and U21112 (N_21112,N_18695,N_18954);
nor U21113 (N_21113,N_19844,N_19876);
nand U21114 (N_21114,N_19102,N_19214);
xor U21115 (N_21115,N_19376,N_19404);
nor U21116 (N_21116,N_18728,N_19416);
or U21117 (N_21117,N_17532,N_19834);
and U21118 (N_21118,N_17855,N_18397);
xor U21119 (N_21119,N_19708,N_18328);
or U21120 (N_21120,N_19306,N_19787);
and U21121 (N_21121,N_17964,N_18732);
xnor U21122 (N_21122,N_18802,N_19662);
nand U21123 (N_21123,N_19607,N_17952);
nand U21124 (N_21124,N_17527,N_18019);
and U21125 (N_21125,N_18808,N_18615);
or U21126 (N_21126,N_18877,N_18827);
nand U21127 (N_21127,N_18931,N_19553);
nor U21128 (N_21128,N_17585,N_19557);
and U21129 (N_21129,N_19930,N_18678);
or U21130 (N_21130,N_18368,N_19176);
or U21131 (N_21131,N_18421,N_18975);
nor U21132 (N_21132,N_19947,N_18765);
nor U21133 (N_21133,N_18525,N_18721);
nor U21134 (N_21134,N_19118,N_19080);
xnor U21135 (N_21135,N_19317,N_19117);
or U21136 (N_21136,N_17587,N_18607);
nor U21137 (N_21137,N_19514,N_18810);
xor U21138 (N_21138,N_19435,N_19291);
xnor U21139 (N_21139,N_19197,N_19516);
xor U21140 (N_21140,N_18950,N_17625);
nor U21141 (N_21141,N_18848,N_17933);
xnor U21142 (N_21142,N_19862,N_18523);
xor U21143 (N_21143,N_19867,N_17737);
nor U21144 (N_21144,N_18597,N_17512);
xor U21145 (N_21145,N_17792,N_19209);
nand U21146 (N_21146,N_18122,N_18758);
and U21147 (N_21147,N_17557,N_18109);
or U21148 (N_21148,N_19657,N_18667);
nor U21149 (N_21149,N_19707,N_18591);
xnor U21150 (N_21150,N_17558,N_18812);
nor U21151 (N_21151,N_17854,N_19362);
nand U21152 (N_21152,N_18267,N_17804);
xor U21153 (N_21153,N_18181,N_18769);
or U21154 (N_21154,N_17989,N_19227);
and U21155 (N_21155,N_18340,N_18184);
or U21156 (N_21156,N_19008,N_17768);
nand U21157 (N_21157,N_17816,N_18253);
nand U21158 (N_21158,N_19303,N_18701);
or U21159 (N_21159,N_18941,N_18238);
xor U21160 (N_21160,N_18073,N_18714);
and U21161 (N_21161,N_17565,N_18277);
nand U21162 (N_21162,N_18304,N_17926);
nor U21163 (N_21163,N_17761,N_19211);
or U21164 (N_21164,N_18800,N_18082);
or U21165 (N_21165,N_18873,N_18156);
and U21166 (N_21166,N_19472,N_19300);
or U21167 (N_21167,N_18422,N_18624);
or U21168 (N_21168,N_19429,N_18363);
and U21169 (N_21169,N_17809,N_19143);
nor U21170 (N_21170,N_18745,N_18976);
xor U21171 (N_21171,N_17767,N_19097);
xor U21172 (N_21172,N_18112,N_18746);
or U21173 (N_21173,N_19078,N_18781);
xnor U21174 (N_21174,N_18257,N_17712);
nor U21175 (N_21175,N_18449,N_17660);
or U21176 (N_21176,N_18376,N_18048);
or U21177 (N_21177,N_18358,N_17843);
or U21178 (N_21178,N_18167,N_19264);
nand U21179 (N_21179,N_18308,N_18855);
xnor U21180 (N_21180,N_18619,N_18039);
nand U21181 (N_21181,N_17569,N_19427);
and U21182 (N_21182,N_17857,N_18009);
xnor U21183 (N_21183,N_17634,N_19669);
or U21184 (N_21184,N_19049,N_19625);
xnor U21185 (N_21185,N_18861,N_19617);
xor U21186 (N_21186,N_17935,N_19838);
and U21187 (N_21187,N_19165,N_19018);
and U21188 (N_21188,N_19545,N_18198);
nor U21189 (N_21189,N_19410,N_17992);
nand U21190 (N_21190,N_18788,N_18004);
xnor U21191 (N_21191,N_19320,N_17882);
nand U21192 (N_21192,N_17889,N_19383);
nand U21193 (N_21193,N_18118,N_18473);
and U21194 (N_21194,N_17867,N_18180);
or U21195 (N_21195,N_18006,N_19540);
nand U21196 (N_21196,N_18055,N_18441);
nor U21197 (N_21197,N_18145,N_17588);
and U21198 (N_21198,N_19181,N_19498);
and U21199 (N_21199,N_19762,N_18617);
or U21200 (N_21200,N_19677,N_17628);
nand U21201 (N_21201,N_19904,N_19045);
xnor U21202 (N_21202,N_19527,N_18747);
or U21203 (N_21203,N_18147,N_19325);
nor U21204 (N_21204,N_18236,N_19065);
xor U21205 (N_21205,N_19099,N_19990);
nand U21206 (N_21206,N_18915,N_18031);
or U21207 (N_21207,N_19489,N_19351);
nor U21208 (N_21208,N_19626,N_18621);
xnor U21209 (N_21209,N_18712,N_19759);
nand U21210 (N_21210,N_17685,N_19338);
nand U21211 (N_21211,N_17841,N_19027);
or U21212 (N_21212,N_18151,N_18420);
xor U21213 (N_21213,N_18508,N_17764);
nand U21214 (N_21214,N_19290,N_18832);
and U21215 (N_21215,N_17784,N_18646);
xnor U21216 (N_21216,N_18890,N_18001);
and U21217 (N_21217,N_19731,N_18102);
nand U21218 (N_21218,N_19407,N_19761);
xor U21219 (N_21219,N_18317,N_17698);
nor U21220 (N_21220,N_19339,N_17980);
or U21221 (N_21221,N_18644,N_19323);
xnor U21222 (N_21222,N_18570,N_19474);
xor U21223 (N_21223,N_18618,N_18785);
nor U21224 (N_21224,N_18966,N_17508);
or U21225 (N_21225,N_18664,N_18374);
and U21226 (N_21226,N_19116,N_19103);
nand U21227 (N_21227,N_19757,N_19057);
xnor U21228 (N_21228,N_19379,N_19530);
xnor U21229 (N_21229,N_19921,N_19332);
xor U21230 (N_21230,N_18440,N_17509);
or U21231 (N_21231,N_17644,N_19137);
xnor U21232 (N_21232,N_18177,N_18056);
and U21233 (N_21233,N_18079,N_19751);
or U21234 (N_21234,N_19501,N_19865);
or U21235 (N_21235,N_18780,N_19148);
and U21236 (N_21236,N_17524,N_18515);
xnor U21237 (N_21237,N_18444,N_17534);
and U21238 (N_21238,N_17684,N_18670);
xnor U21239 (N_21239,N_19900,N_19680);
or U21240 (N_21240,N_18885,N_18584);
and U21241 (N_21241,N_18300,N_18301);
xor U21242 (N_21242,N_19479,N_18443);
and U21243 (N_21243,N_18811,N_18168);
xnor U21244 (N_21244,N_19473,N_18204);
nand U21245 (N_21245,N_18906,N_19064);
and U21246 (N_21246,N_19200,N_18904);
xor U21247 (N_21247,N_19201,N_19124);
nand U21248 (N_21248,N_19386,N_19232);
nand U21249 (N_21249,N_19146,N_18051);
xnor U21250 (N_21250,N_18549,N_17665);
and U21251 (N_21251,N_19893,N_17939);
or U21252 (N_21252,N_18228,N_18137);
nor U21253 (N_21253,N_19849,N_18748);
or U21254 (N_21254,N_19796,N_19676);
and U21255 (N_21255,N_17946,N_18677);
xnor U21256 (N_21256,N_17974,N_18309);
or U21257 (N_21257,N_17897,N_19762);
and U21258 (N_21258,N_18501,N_17550);
or U21259 (N_21259,N_18473,N_17932);
and U21260 (N_21260,N_19126,N_18912);
xor U21261 (N_21261,N_19657,N_19986);
xnor U21262 (N_21262,N_19040,N_18329);
xnor U21263 (N_21263,N_19844,N_19557);
xor U21264 (N_21264,N_17758,N_19451);
nand U21265 (N_21265,N_19627,N_19530);
nor U21266 (N_21266,N_18618,N_17663);
nor U21267 (N_21267,N_17861,N_18041);
nand U21268 (N_21268,N_19660,N_18711);
nor U21269 (N_21269,N_18008,N_17748);
nor U21270 (N_21270,N_18046,N_18978);
xor U21271 (N_21271,N_19666,N_19942);
nand U21272 (N_21272,N_17583,N_18655);
or U21273 (N_21273,N_18575,N_19246);
and U21274 (N_21274,N_19116,N_19702);
xor U21275 (N_21275,N_17896,N_18839);
nor U21276 (N_21276,N_19970,N_19068);
xor U21277 (N_21277,N_18889,N_17917);
nor U21278 (N_21278,N_19673,N_19757);
nor U21279 (N_21279,N_18510,N_19189);
nor U21280 (N_21280,N_17942,N_19288);
and U21281 (N_21281,N_19683,N_18692);
xor U21282 (N_21282,N_18558,N_19764);
xnor U21283 (N_21283,N_18453,N_18988);
nor U21284 (N_21284,N_18152,N_19127);
xor U21285 (N_21285,N_17775,N_17651);
xor U21286 (N_21286,N_19468,N_17613);
or U21287 (N_21287,N_19027,N_18640);
nor U21288 (N_21288,N_19602,N_17955);
nor U21289 (N_21289,N_17833,N_17538);
nand U21290 (N_21290,N_19572,N_17823);
nor U21291 (N_21291,N_18699,N_18402);
xnor U21292 (N_21292,N_19176,N_18594);
and U21293 (N_21293,N_17751,N_19503);
and U21294 (N_21294,N_19125,N_18454);
nor U21295 (N_21295,N_18525,N_17625);
xor U21296 (N_21296,N_18399,N_17508);
xor U21297 (N_21297,N_19189,N_19113);
nor U21298 (N_21298,N_19355,N_17892);
nor U21299 (N_21299,N_17925,N_18473);
nand U21300 (N_21300,N_18471,N_17905);
or U21301 (N_21301,N_19936,N_17932);
xor U21302 (N_21302,N_18699,N_18714);
and U21303 (N_21303,N_17881,N_18367);
xnor U21304 (N_21304,N_18268,N_19750);
xnor U21305 (N_21305,N_18320,N_17696);
and U21306 (N_21306,N_18032,N_17524);
nor U21307 (N_21307,N_18072,N_18458);
nand U21308 (N_21308,N_19972,N_17939);
and U21309 (N_21309,N_18542,N_17533);
and U21310 (N_21310,N_18190,N_19295);
nand U21311 (N_21311,N_18605,N_19842);
nand U21312 (N_21312,N_19066,N_17500);
nand U21313 (N_21313,N_17730,N_18181);
and U21314 (N_21314,N_18589,N_19123);
or U21315 (N_21315,N_19311,N_18905);
and U21316 (N_21316,N_18716,N_18897);
nor U21317 (N_21317,N_18822,N_17628);
or U21318 (N_21318,N_18238,N_19630);
nand U21319 (N_21319,N_19597,N_18097);
or U21320 (N_21320,N_19487,N_19506);
nor U21321 (N_21321,N_19667,N_17735);
xnor U21322 (N_21322,N_19443,N_18986);
nand U21323 (N_21323,N_19676,N_18651);
nor U21324 (N_21324,N_17657,N_19901);
nor U21325 (N_21325,N_19292,N_19422);
nand U21326 (N_21326,N_18163,N_17513);
nor U21327 (N_21327,N_18096,N_17603);
or U21328 (N_21328,N_18601,N_17954);
nand U21329 (N_21329,N_17978,N_18916);
nor U21330 (N_21330,N_18427,N_19655);
nor U21331 (N_21331,N_18080,N_19660);
or U21332 (N_21332,N_18395,N_17790);
nor U21333 (N_21333,N_17647,N_19994);
xnor U21334 (N_21334,N_19594,N_18855);
or U21335 (N_21335,N_19485,N_18019);
xnor U21336 (N_21336,N_18683,N_17998);
nand U21337 (N_21337,N_19521,N_19052);
nor U21338 (N_21338,N_18899,N_17945);
xor U21339 (N_21339,N_18290,N_18926);
nand U21340 (N_21340,N_18241,N_17856);
xor U21341 (N_21341,N_17819,N_19492);
nor U21342 (N_21342,N_17635,N_19122);
and U21343 (N_21343,N_18720,N_19345);
and U21344 (N_21344,N_18462,N_18653);
or U21345 (N_21345,N_19518,N_19184);
xnor U21346 (N_21346,N_18593,N_18363);
nand U21347 (N_21347,N_18763,N_18646);
or U21348 (N_21348,N_19673,N_17997);
nand U21349 (N_21349,N_17959,N_19816);
and U21350 (N_21350,N_19140,N_18229);
nor U21351 (N_21351,N_18775,N_19195);
and U21352 (N_21352,N_17822,N_18491);
xnor U21353 (N_21353,N_18319,N_18445);
nor U21354 (N_21354,N_17773,N_18138);
nor U21355 (N_21355,N_19364,N_19502);
and U21356 (N_21356,N_17628,N_18927);
xnor U21357 (N_21357,N_18767,N_18709);
and U21358 (N_21358,N_19926,N_19352);
nand U21359 (N_21359,N_18855,N_18475);
xor U21360 (N_21360,N_19873,N_17929);
xor U21361 (N_21361,N_18031,N_19557);
or U21362 (N_21362,N_18573,N_18820);
or U21363 (N_21363,N_17820,N_19165);
xnor U21364 (N_21364,N_18810,N_18859);
xnor U21365 (N_21365,N_19624,N_17549);
and U21366 (N_21366,N_19641,N_18120);
or U21367 (N_21367,N_18683,N_18311);
or U21368 (N_21368,N_18804,N_19211);
xnor U21369 (N_21369,N_18220,N_19170);
or U21370 (N_21370,N_19495,N_17868);
nor U21371 (N_21371,N_19585,N_17668);
nor U21372 (N_21372,N_17820,N_19463);
nor U21373 (N_21373,N_18726,N_17823);
or U21374 (N_21374,N_17855,N_17661);
nand U21375 (N_21375,N_19328,N_18690);
nand U21376 (N_21376,N_18482,N_17852);
nor U21377 (N_21377,N_19265,N_19145);
xnor U21378 (N_21378,N_19851,N_18601);
and U21379 (N_21379,N_19645,N_17820);
and U21380 (N_21380,N_18612,N_19074);
xnor U21381 (N_21381,N_19307,N_18156);
nor U21382 (N_21382,N_17746,N_19269);
nand U21383 (N_21383,N_18671,N_19923);
or U21384 (N_21384,N_18927,N_18382);
xor U21385 (N_21385,N_18542,N_19253);
or U21386 (N_21386,N_19915,N_19091);
nand U21387 (N_21387,N_18260,N_17950);
xnor U21388 (N_21388,N_18863,N_17746);
nor U21389 (N_21389,N_19196,N_18425);
nor U21390 (N_21390,N_18759,N_17501);
nand U21391 (N_21391,N_19409,N_17979);
nand U21392 (N_21392,N_18310,N_18541);
or U21393 (N_21393,N_18918,N_17542);
xnor U21394 (N_21394,N_19549,N_18904);
nor U21395 (N_21395,N_17950,N_18389);
nand U21396 (N_21396,N_17659,N_19458);
nand U21397 (N_21397,N_18449,N_17931);
and U21398 (N_21398,N_19250,N_19129);
xor U21399 (N_21399,N_19183,N_18377);
nor U21400 (N_21400,N_18207,N_18856);
and U21401 (N_21401,N_19267,N_17666);
and U21402 (N_21402,N_19082,N_18427);
or U21403 (N_21403,N_18637,N_18009);
and U21404 (N_21404,N_18696,N_19412);
nor U21405 (N_21405,N_18537,N_19426);
or U21406 (N_21406,N_19267,N_17858);
and U21407 (N_21407,N_19431,N_19481);
nand U21408 (N_21408,N_18625,N_18386);
or U21409 (N_21409,N_19871,N_19812);
and U21410 (N_21410,N_19365,N_19630);
nor U21411 (N_21411,N_18559,N_18254);
and U21412 (N_21412,N_19751,N_19155);
xor U21413 (N_21413,N_18536,N_19350);
nand U21414 (N_21414,N_19742,N_19772);
and U21415 (N_21415,N_18683,N_18417);
or U21416 (N_21416,N_19129,N_19614);
or U21417 (N_21417,N_17567,N_18141);
nand U21418 (N_21418,N_18165,N_18423);
and U21419 (N_21419,N_19989,N_17756);
nand U21420 (N_21420,N_19788,N_17813);
nor U21421 (N_21421,N_18496,N_18826);
xnor U21422 (N_21422,N_19871,N_19545);
and U21423 (N_21423,N_19751,N_17685);
xor U21424 (N_21424,N_19882,N_19430);
and U21425 (N_21425,N_18259,N_19106);
nor U21426 (N_21426,N_18189,N_19924);
nand U21427 (N_21427,N_19230,N_19091);
and U21428 (N_21428,N_19462,N_19482);
xnor U21429 (N_21429,N_17967,N_18668);
nand U21430 (N_21430,N_17526,N_19089);
xnor U21431 (N_21431,N_18840,N_19460);
nor U21432 (N_21432,N_18397,N_19021);
nand U21433 (N_21433,N_18707,N_18693);
nand U21434 (N_21434,N_19514,N_19840);
nand U21435 (N_21435,N_19710,N_19432);
nand U21436 (N_21436,N_19313,N_19696);
xor U21437 (N_21437,N_17525,N_17559);
nand U21438 (N_21438,N_19729,N_18151);
nand U21439 (N_21439,N_19713,N_18202);
and U21440 (N_21440,N_18596,N_18553);
or U21441 (N_21441,N_18906,N_18486);
xor U21442 (N_21442,N_18680,N_19949);
or U21443 (N_21443,N_17520,N_17759);
or U21444 (N_21444,N_18495,N_18981);
or U21445 (N_21445,N_17908,N_18296);
xor U21446 (N_21446,N_19800,N_19412);
and U21447 (N_21447,N_18889,N_18863);
or U21448 (N_21448,N_18622,N_19500);
or U21449 (N_21449,N_18531,N_17853);
or U21450 (N_21450,N_19332,N_18535);
or U21451 (N_21451,N_18749,N_19168);
nor U21452 (N_21452,N_17639,N_18988);
nor U21453 (N_21453,N_19103,N_18843);
nor U21454 (N_21454,N_19834,N_19082);
and U21455 (N_21455,N_18693,N_17883);
or U21456 (N_21456,N_19810,N_17805);
xnor U21457 (N_21457,N_19122,N_18565);
and U21458 (N_21458,N_19139,N_17825);
and U21459 (N_21459,N_18167,N_19128);
or U21460 (N_21460,N_19228,N_18769);
or U21461 (N_21461,N_18484,N_18455);
nand U21462 (N_21462,N_18038,N_18508);
xor U21463 (N_21463,N_18312,N_17709);
and U21464 (N_21464,N_18191,N_18801);
nor U21465 (N_21465,N_19566,N_19621);
or U21466 (N_21466,N_19254,N_18475);
nor U21467 (N_21467,N_19681,N_19990);
or U21468 (N_21468,N_19048,N_18309);
nor U21469 (N_21469,N_18545,N_19322);
nor U21470 (N_21470,N_18514,N_18395);
or U21471 (N_21471,N_19848,N_18193);
xnor U21472 (N_21472,N_18251,N_17516);
and U21473 (N_21473,N_19299,N_19300);
nand U21474 (N_21474,N_18472,N_18106);
and U21475 (N_21475,N_19736,N_19384);
nor U21476 (N_21476,N_19193,N_19047);
or U21477 (N_21477,N_18202,N_18050);
nor U21478 (N_21478,N_18366,N_19460);
nand U21479 (N_21479,N_18138,N_19801);
xnor U21480 (N_21480,N_18168,N_17690);
and U21481 (N_21481,N_19963,N_18850);
xor U21482 (N_21482,N_18369,N_17557);
or U21483 (N_21483,N_19931,N_18536);
and U21484 (N_21484,N_18002,N_19587);
nand U21485 (N_21485,N_19959,N_19444);
nand U21486 (N_21486,N_18035,N_18782);
and U21487 (N_21487,N_19918,N_18425);
nand U21488 (N_21488,N_19675,N_18935);
and U21489 (N_21489,N_19713,N_18804);
nand U21490 (N_21490,N_17896,N_18595);
nand U21491 (N_21491,N_18978,N_19247);
and U21492 (N_21492,N_19729,N_19074);
nor U21493 (N_21493,N_19381,N_17889);
xnor U21494 (N_21494,N_17549,N_17659);
and U21495 (N_21495,N_19833,N_18559);
nand U21496 (N_21496,N_19231,N_19114);
and U21497 (N_21497,N_19618,N_17598);
nand U21498 (N_21498,N_17866,N_19347);
and U21499 (N_21499,N_18351,N_19118);
nand U21500 (N_21500,N_18699,N_18627);
nor U21501 (N_21501,N_18350,N_18248);
nand U21502 (N_21502,N_19870,N_18578);
nand U21503 (N_21503,N_18593,N_17744);
or U21504 (N_21504,N_18397,N_18553);
or U21505 (N_21505,N_17966,N_17947);
nor U21506 (N_21506,N_19671,N_17765);
and U21507 (N_21507,N_18031,N_18441);
nand U21508 (N_21508,N_19384,N_19716);
xor U21509 (N_21509,N_19648,N_19080);
or U21510 (N_21510,N_19689,N_17525);
xor U21511 (N_21511,N_18382,N_19987);
nor U21512 (N_21512,N_18454,N_17504);
nand U21513 (N_21513,N_17974,N_19122);
xnor U21514 (N_21514,N_19534,N_19912);
nor U21515 (N_21515,N_18544,N_18801);
nor U21516 (N_21516,N_18223,N_19906);
nor U21517 (N_21517,N_18607,N_18937);
xor U21518 (N_21518,N_18123,N_18778);
or U21519 (N_21519,N_19914,N_18310);
and U21520 (N_21520,N_19204,N_19564);
and U21521 (N_21521,N_19438,N_19727);
or U21522 (N_21522,N_19206,N_19761);
and U21523 (N_21523,N_17766,N_17660);
nand U21524 (N_21524,N_19781,N_19901);
or U21525 (N_21525,N_18447,N_19142);
nand U21526 (N_21526,N_18011,N_18266);
nand U21527 (N_21527,N_18827,N_18699);
xnor U21528 (N_21528,N_18129,N_17714);
or U21529 (N_21529,N_19338,N_19861);
and U21530 (N_21530,N_17846,N_18605);
or U21531 (N_21531,N_17553,N_19193);
nor U21532 (N_21532,N_19666,N_19262);
and U21533 (N_21533,N_18064,N_19111);
and U21534 (N_21534,N_19305,N_19393);
or U21535 (N_21535,N_18835,N_19183);
or U21536 (N_21536,N_19917,N_18367);
and U21537 (N_21537,N_17700,N_17601);
nor U21538 (N_21538,N_17980,N_17762);
and U21539 (N_21539,N_18348,N_18154);
nor U21540 (N_21540,N_19059,N_19980);
and U21541 (N_21541,N_18137,N_19268);
xor U21542 (N_21542,N_18147,N_17599);
or U21543 (N_21543,N_19939,N_18404);
xnor U21544 (N_21544,N_18346,N_18919);
nor U21545 (N_21545,N_17579,N_17589);
or U21546 (N_21546,N_18820,N_18570);
nand U21547 (N_21547,N_19825,N_19926);
and U21548 (N_21548,N_19012,N_18226);
or U21549 (N_21549,N_19494,N_18321);
xnor U21550 (N_21550,N_18526,N_19641);
and U21551 (N_21551,N_19726,N_17945);
xor U21552 (N_21552,N_18300,N_19711);
or U21553 (N_21553,N_18848,N_18122);
or U21554 (N_21554,N_18645,N_17839);
nand U21555 (N_21555,N_18912,N_19828);
nor U21556 (N_21556,N_18658,N_17987);
and U21557 (N_21557,N_19947,N_19524);
or U21558 (N_21558,N_19723,N_18334);
and U21559 (N_21559,N_18122,N_19481);
nor U21560 (N_21560,N_18301,N_18654);
nand U21561 (N_21561,N_18360,N_18340);
xnor U21562 (N_21562,N_19444,N_18564);
xnor U21563 (N_21563,N_19581,N_19742);
nor U21564 (N_21564,N_18591,N_18951);
xor U21565 (N_21565,N_19787,N_19891);
nor U21566 (N_21566,N_19688,N_18742);
or U21567 (N_21567,N_18446,N_19844);
xnor U21568 (N_21568,N_19341,N_19610);
nor U21569 (N_21569,N_19893,N_18238);
nand U21570 (N_21570,N_17938,N_18063);
nor U21571 (N_21571,N_17621,N_19610);
nand U21572 (N_21572,N_18243,N_19017);
nand U21573 (N_21573,N_17873,N_19994);
xor U21574 (N_21574,N_17975,N_17657);
and U21575 (N_21575,N_18844,N_19366);
nor U21576 (N_21576,N_18740,N_18269);
xor U21577 (N_21577,N_18291,N_19665);
or U21578 (N_21578,N_19296,N_19383);
nor U21579 (N_21579,N_17701,N_19192);
or U21580 (N_21580,N_19187,N_19848);
nor U21581 (N_21581,N_19244,N_19222);
nand U21582 (N_21582,N_18015,N_19504);
or U21583 (N_21583,N_17625,N_18070);
xor U21584 (N_21584,N_18924,N_19680);
and U21585 (N_21585,N_18202,N_19290);
xor U21586 (N_21586,N_17563,N_18830);
and U21587 (N_21587,N_17841,N_18544);
or U21588 (N_21588,N_19295,N_17731);
nand U21589 (N_21589,N_18553,N_17993);
xnor U21590 (N_21590,N_19979,N_18594);
nor U21591 (N_21591,N_18746,N_19039);
nand U21592 (N_21592,N_19880,N_18164);
or U21593 (N_21593,N_19396,N_17800);
nand U21594 (N_21594,N_19624,N_19893);
and U21595 (N_21595,N_19322,N_18541);
and U21596 (N_21596,N_18964,N_19764);
nor U21597 (N_21597,N_17650,N_19294);
xnor U21598 (N_21598,N_19676,N_17858);
nand U21599 (N_21599,N_17739,N_18600);
nor U21600 (N_21600,N_18051,N_18280);
and U21601 (N_21601,N_19547,N_19086);
xnor U21602 (N_21602,N_17667,N_18717);
nor U21603 (N_21603,N_17651,N_19927);
and U21604 (N_21604,N_18269,N_19794);
nor U21605 (N_21605,N_19869,N_19601);
nor U21606 (N_21606,N_19482,N_17634);
and U21607 (N_21607,N_19604,N_17855);
nor U21608 (N_21608,N_19041,N_18859);
nor U21609 (N_21609,N_19078,N_17741);
xnor U21610 (N_21610,N_17929,N_18177);
and U21611 (N_21611,N_18091,N_19567);
xnor U21612 (N_21612,N_18106,N_17538);
nor U21613 (N_21613,N_19093,N_18881);
nand U21614 (N_21614,N_17848,N_18886);
nor U21615 (N_21615,N_17966,N_19032);
nand U21616 (N_21616,N_18012,N_18204);
and U21617 (N_21617,N_19357,N_18228);
nand U21618 (N_21618,N_18306,N_18380);
xor U21619 (N_21619,N_19605,N_19802);
nor U21620 (N_21620,N_17678,N_18594);
nor U21621 (N_21621,N_19326,N_18519);
xor U21622 (N_21622,N_19268,N_17839);
and U21623 (N_21623,N_19928,N_19626);
nand U21624 (N_21624,N_18530,N_17868);
nand U21625 (N_21625,N_17713,N_18251);
xor U21626 (N_21626,N_18838,N_19998);
nand U21627 (N_21627,N_17691,N_19479);
nand U21628 (N_21628,N_17954,N_18879);
xor U21629 (N_21629,N_19462,N_19903);
or U21630 (N_21630,N_17864,N_19377);
xor U21631 (N_21631,N_19468,N_19250);
and U21632 (N_21632,N_18344,N_18028);
xor U21633 (N_21633,N_19898,N_18438);
or U21634 (N_21634,N_17617,N_19749);
nor U21635 (N_21635,N_19325,N_17633);
and U21636 (N_21636,N_18184,N_17917);
xor U21637 (N_21637,N_18361,N_18010);
or U21638 (N_21638,N_18818,N_17983);
and U21639 (N_21639,N_19841,N_17841);
or U21640 (N_21640,N_19063,N_19553);
nor U21641 (N_21641,N_17697,N_18060);
nand U21642 (N_21642,N_17616,N_19397);
nor U21643 (N_21643,N_19196,N_18212);
or U21644 (N_21644,N_18316,N_19124);
xor U21645 (N_21645,N_19671,N_19096);
nor U21646 (N_21646,N_18200,N_19609);
or U21647 (N_21647,N_19841,N_19523);
xor U21648 (N_21648,N_18827,N_19667);
nand U21649 (N_21649,N_18146,N_19242);
and U21650 (N_21650,N_19157,N_19912);
and U21651 (N_21651,N_19212,N_19558);
nand U21652 (N_21652,N_18469,N_19353);
or U21653 (N_21653,N_19212,N_18000);
xor U21654 (N_21654,N_18359,N_18673);
xnor U21655 (N_21655,N_19123,N_18050);
nor U21656 (N_21656,N_18196,N_17717);
nand U21657 (N_21657,N_18708,N_18639);
or U21658 (N_21658,N_19285,N_17531);
xnor U21659 (N_21659,N_18610,N_19978);
nand U21660 (N_21660,N_18240,N_17898);
nand U21661 (N_21661,N_19969,N_18272);
xnor U21662 (N_21662,N_19544,N_19838);
xnor U21663 (N_21663,N_19367,N_17938);
nor U21664 (N_21664,N_17830,N_19198);
nand U21665 (N_21665,N_18361,N_17899);
or U21666 (N_21666,N_18809,N_19274);
xnor U21667 (N_21667,N_17918,N_18892);
xor U21668 (N_21668,N_17881,N_19852);
nand U21669 (N_21669,N_18184,N_18074);
and U21670 (N_21670,N_17517,N_19564);
xor U21671 (N_21671,N_18357,N_18556);
xnor U21672 (N_21672,N_17830,N_19635);
or U21673 (N_21673,N_19776,N_18968);
or U21674 (N_21674,N_17599,N_18382);
nand U21675 (N_21675,N_18303,N_19580);
nor U21676 (N_21676,N_18592,N_19650);
nor U21677 (N_21677,N_18929,N_18168);
xnor U21678 (N_21678,N_18552,N_18927);
xnor U21679 (N_21679,N_17923,N_18991);
nor U21680 (N_21680,N_19295,N_19932);
nand U21681 (N_21681,N_18875,N_17520);
nand U21682 (N_21682,N_18711,N_19418);
and U21683 (N_21683,N_17533,N_17506);
or U21684 (N_21684,N_18403,N_17608);
xnor U21685 (N_21685,N_19923,N_18748);
and U21686 (N_21686,N_17584,N_19214);
or U21687 (N_21687,N_17997,N_17534);
xor U21688 (N_21688,N_18099,N_19912);
nor U21689 (N_21689,N_19897,N_18793);
or U21690 (N_21690,N_19922,N_17892);
nor U21691 (N_21691,N_17892,N_19050);
or U21692 (N_21692,N_17635,N_19462);
xnor U21693 (N_21693,N_18751,N_17665);
and U21694 (N_21694,N_19340,N_19143);
nor U21695 (N_21695,N_18460,N_17993);
xor U21696 (N_21696,N_19746,N_19092);
and U21697 (N_21697,N_19796,N_17798);
nor U21698 (N_21698,N_19118,N_18559);
nor U21699 (N_21699,N_18161,N_18924);
nor U21700 (N_21700,N_19827,N_19378);
xor U21701 (N_21701,N_18351,N_19385);
xnor U21702 (N_21702,N_18408,N_19821);
xor U21703 (N_21703,N_17816,N_18176);
xor U21704 (N_21704,N_19462,N_19761);
nor U21705 (N_21705,N_19096,N_19684);
nand U21706 (N_21706,N_18292,N_18467);
nand U21707 (N_21707,N_19539,N_19037);
xor U21708 (N_21708,N_19679,N_19441);
nand U21709 (N_21709,N_18128,N_18493);
nor U21710 (N_21710,N_19276,N_19079);
xnor U21711 (N_21711,N_18349,N_19498);
xnor U21712 (N_21712,N_17665,N_19991);
nand U21713 (N_21713,N_19008,N_19150);
and U21714 (N_21714,N_19125,N_19810);
nor U21715 (N_21715,N_18234,N_19168);
or U21716 (N_21716,N_19272,N_17622);
nand U21717 (N_21717,N_19483,N_18612);
nor U21718 (N_21718,N_18843,N_18252);
xnor U21719 (N_21719,N_19880,N_19887);
nand U21720 (N_21720,N_17795,N_18825);
and U21721 (N_21721,N_17575,N_17993);
xnor U21722 (N_21722,N_19580,N_19884);
and U21723 (N_21723,N_19630,N_18804);
or U21724 (N_21724,N_19820,N_17782);
nor U21725 (N_21725,N_19745,N_18401);
and U21726 (N_21726,N_18114,N_17741);
xor U21727 (N_21727,N_17902,N_18744);
and U21728 (N_21728,N_19821,N_18024);
nand U21729 (N_21729,N_19953,N_17898);
or U21730 (N_21730,N_18079,N_19638);
or U21731 (N_21731,N_17676,N_17719);
nand U21732 (N_21732,N_19878,N_19507);
xnor U21733 (N_21733,N_18876,N_19401);
xor U21734 (N_21734,N_17504,N_18994);
nand U21735 (N_21735,N_19252,N_17743);
and U21736 (N_21736,N_18153,N_17590);
xnor U21737 (N_21737,N_18975,N_19279);
nor U21738 (N_21738,N_18706,N_17553);
or U21739 (N_21739,N_18115,N_17602);
or U21740 (N_21740,N_17845,N_18608);
nor U21741 (N_21741,N_18327,N_19933);
xnor U21742 (N_21742,N_17899,N_18093);
or U21743 (N_21743,N_18766,N_19196);
xor U21744 (N_21744,N_19502,N_19990);
or U21745 (N_21745,N_17823,N_19133);
and U21746 (N_21746,N_19617,N_17635);
nand U21747 (N_21747,N_17608,N_18318);
and U21748 (N_21748,N_19248,N_19240);
and U21749 (N_21749,N_19084,N_18685);
and U21750 (N_21750,N_18346,N_19749);
and U21751 (N_21751,N_18196,N_18950);
nand U21752 (N_21752,N_19007,N_17646);
nand U21753 (N_21753,N_18172,N_17602);
nand U21754 (N_21754,N_18059,N_18562);
nor U21755 (N_21755,N_18643,N_18908);
and U21756 (N_21756,N_18141,N_17834);
xor U21757 (N_21757,N_18857,N_17847);
and U21758 (N_21758,N_19454,N_18465);
nand U21759 (N_21759,N_19170,N_18571);
and U21760 (N_21760,N_18655,N_19397);
xnor U21761 (N_21761,N_18988,N_18150);
or U21762 (N_21762,N_17967,N_18632);
nand U21763 (N_21763,N_18351,N_18517);
and U21764 (N_21764,N_18113,N_19695);
nand U21765 (N_21765,N_18134,N_18765);
and U21766 (N_21766,N_19399,N_17835);
nand U21767 (N_21767,N_18290,N_17524);
nor U21768 (N_21768,N_19182,N_17930);
xnor U21769 (N_21769,N_19984,N_17935);
nand U21770 (N_21770,N_17675,N_17728);
xnor U21771 (N_21771,N_19516,N_18416);
nor U21772 (N_21772,N_18883,N_19829);
nor U21773 (N_21773,N_17977,N_17912);
nand U21774 (N_21774,N_18562,N_17685);
or U21775 (N_21775,N_19132,N_19277);
xnor U21776 (N_21776,N_18574,N_17525);
and U21777 (N_21777,N_19990,N_19697);
xor U21778 (N_21778,N_18780,N_18481);
and U21779 (N_21779,N_17679,N_18247);
and U21780 (N_21780,N_17611,N_19548);
or U21781 (N_21781,N_19641,N_19626);
xor U21782 (N_21782,N_18201,N_19235);
or U21783 (N_21783,N_19895,N_19207);
nand U21784 (N_21784,N_19543,N_19005);
nor U21785 (N_21785,N_18145,N_19610);
and U21786 (N_21786,N_17539,N_17754);
xor U21787 (N_21787,N_18189,N_18908);
nor U21788 (N_21788,N_19319,N_17644);
xor U21789 (N_21789,N_17695,N_18807);
nor U21790 (N_21790,N_18762,N_19913);
or U21791 (N_21791,N_19073,N_18732);
or U21792 (N_21792,N_19037,N_18799);
nor U21793 (N_21793,N_19254,N_19766);
nand U21794 (N_21794,N_18981,N_19045);
or U21795 (N_21795,N_19423,N_17819);
xnor U21796 (N_21796,N_17869,N_18912);
or U21797 (N_21797,N_18837,N_19304);
nand U21798 (N_21798,N_18857,N_17937);
nor U21799 (N_21799,N_17997,N_19052);
nand U21800 (N_21800,N_18063,N_19350);
nor U21801 (N_21801,N_18615,N_18884);
and U21802 (N_21802,N_18713,N_19393);
nor U21803 (N_21803,N_18899,N_19869);
xnor U21804 (N_21804,N_18693,N_19829);
nand U21805 (N_21805,N_19250,N_18802);
xor U21806 (N_21806,N_18354,N_17915);
nand U21807 (N_21807,N_19117,N_19767);
xor U21808 (N_21808,N_19416,N_17946);
nand U21809 (N_21809,N_17906,N_18081);
or U21810 (N_21810,N_18909,N_17639);
or U21811 (N_21811,N_18856,N_19979);
or U21812 (N_21812,N_19248,N_18127);
nor U21813 (N_21813,N_18156,N_19251);
xor U21814 (N_21814,N_18606,N_19513);
or U21815 (N_21815,N_19706,N_17617);
xnor U21816 (N_21816,N_18754,N_18862);
nor U21817 (N_21817,N_17764,N_18853);
nand U21818 (N_21818,N_18955,N_19443);
and U21819 (N_21819,N_18004,N_18428);
xnor U21820 (N_21820,N_18405,N_18010);
and U21821 (N_21821,N_19747,N_17904);
nand U21822 (N_21822,N_18059,N_18556);
xnor U21823 (N_21823,N_19766,N_19941);
xnor U21824 (N_21824,N_18798,N_18792);
xnor U21825 (N_21825,N_18457,N_19579);
xnor U21826 (N_21826,N_17548,N_17920);
or U21827 (N_21827,N_18196,N_19259);
or U21828 (N_21828,N_19414,N_18708);
and U21829 (N_21829,N_19223,N_17692);
nand U21830 (N_21830,N_18170,N_19656);
nand U21831 (N_21831,N_19549,N_18502);
nand U21832 (N_21832,N_17799,N_18617);
or U21833 (N_21833,N_18764,N_18544);
or U21834 (N_21834,N_19910,N_17663);
or U21835 (N_21835,N_18585,N_18451);
or U21836 (N_21836,N_19883,N_18678);
nor U21837 (N_21837,N_17965,N_18251);
nor U21838 (N_21838,N_17529,N_19758);
or U21839 (N_21839,N_19750,N_18738);
or U21840 (N_21840,N_18206,N_19397);
xnor U21841 (N_21841,N_19639,N_17894);
and U21842 (N_21842,N_18981,N_19334);
xor U21843 (N_21843,N_18268,N_19869);
or U21844 (N_21844,N_18427,N_19562);
xor U21845 (N_21845,N_18517,N_19974);
nor U21846 (N_21846,N_19780,N_18161);
xor U21847 (N_21847,N_18404,N_18767);
or U21848 (N_21848,N_19486,N_18327);
or U21849 (N_21849,N_17691,N_19498);
xor U21850 (N_21850,N_19954,N_19526);
xnor U21851 (N_21851,N_19323,N_19941);
nand U21852 (N_21852,N_19804,N_19627);
or U21853 (N_21853,N_17771,N_18782);
xnor U21854 (N_21854,N_19961,N_18326);
and U21855 (N_21855,N_18122,N_17726);
and U21856 (N_21856,N_17849,N_19972);
or U21857 (N_21857,N_17691,N_19025);
xnor U21858 (N_21858,N_19426,N_18281);
xnor U21859 (N_21859,N_19844,N_19622);
and U21860 (N_21860,N_18489,N_17526);
or U21861 (N_21861,N_19675,N_18833);
xor U21862 (N_21862,N_18969,N_19378);
or U21863 (N_21863,N_18387,N_17914);
nor U21864 (N_21864,N_19379,N_18664);
nor U21865 (N_21865,N_19247,N_19022);
nand U21866 (N_21866,N_18547,N_19153);
nor U21867 (N_21867,N_18878,N_18626);
and U21868 (N_21868,N_18601,N_18051);
nand U21869 (N_21869,N_18695,N_19651);
and U21870 (N_21870,N_19898,N_18383);
and U21871 (N_21871,N_19161,N_18457);
xnor U21872 (N_21872,N_17772,N_19730);
xor U21873 (N_21873,N_18111,N_17530);
and U21874 (N_21874,N_19924,N_19556);
or U21875 (N_21875,N_19556,N_17987);
nand U21876 (N_21876,N_19362,N_19142);
and U21877 (N_21877,N_18792,N_18512);
or U21878 (N_21878,N_18584,N_18512);
nand U21879 (N_21879,N_18756,N_19451);
nor U21880 (N_21880,N_19824,N_19895);
nand U21881 (N_21881,N_18876,N_18733);
or U21882 (N_21882,N_19892,N_19207);
xor U21883 (N_21883,N_18320,N_18746);
or U21884 (N_21884,N_17890,N_18962);
xor U21885 (N_21885,N_19329,N_17997);
xor U21886 (N_21886,N_17844,N_18342);
xor U21887 (N_21887,N_18856,N_19116);
or U21888 (N_21888,N_18696,N_18321);
xnor U21889 (N_21889,N_18107,N_19491);
and U21890 (N_21890,N_18239,N_19332);
xnor U21891 (N_21891,N_18441,N_18086);
and U21892 (N_21892,N_17541,N_19271);
xnor U21893 (N_21893,N_18297,N_19405);
and U21894 (N_21894,N_19965,N_18794);
nor U21895 (N_21895,N_19260,N_18444);
and U21896 (N_21896,N_17750,N_19123);
nor U21897 (N_21897,N_17567,N_18580);
nor U21898 (N_21898,N_19371,N_19061);
xnor U21899 (N_21899,N_17955,N_19266);
nor U21900 (N_21900,N_19204,N_18919);
and U21901 (N_21901,N_18362,N_17627);
or U21902 (N_21902,N_19199,N_19253);
or U21903 (N_21903,N_17749,N_19509);
xnor U21904 (N_21904,N_19827,N_19607);
nand U21905 (N_21905,N_17809,N_17944);
and U21906 (N_21906,N_18155,N_18896);
nor U21907 (N_21907,N_18567,N_17623);
nand U21908 (N_21908,N_18374,N_19272);
and U21909 (N_21909,N_19636,N_19952);
or U21910 (N_21910,N_18067,N_18000);
xor U21911 (N_21911,N_19225,N_18980);
and U21912 (N_21912,N_18085,N_19835);
and U21913 (N_21913,N_18018,N_18228);
xor U21914 (N_21914,N_19425,N_18928);
nand U21915 (N_21915,N_19759,N_18195);
and U21916 (N_21916,N_18353,N_18456);
and U21917 (N_21917,N_19784,N_19851);
or U21918 (N_21918,N_19030,N_18920);
xnor U21919 (N_21919,N_19475,N_17880);
or U21920 (N_21920,N_17864,N_19198);
or U21921 (N_21921,N_18930,N_19650);
xnor U21922 (N_21922,N_19487,N_19220);
and U21923 (N_21923,N_18066,N_19725);
nand U21924 (N_21924,N_18920,N_19440);
or U21925 (N_21925,N_17955,N_18881);
nand U21926 (N_21926,N_18097,N_18222);
nand U21927 (N_21927,N_18982,N_18995);
xnor U21928 (N_21928,N_19945,N_18918);
or U21929 (N_21929,N_19071,N_18774);
and U21930 (N_21930,N_18861,N_19370);
and U21931 (N_21931,N_18149,N_18935);
or U21932 (N_21932,N_18742,N_19731);
and U21933 (N_21933,N_17710,N_18061);
xor U21934 (N_21934,N_17580,N_18323);
and U21935 (N_21935,N_18807,N_18554);
nand U21936 (N_21936,N_17597,N_18067);
nor U21937 (N_21937,N_19444,N_19401);
nor U21938 (N_21938,N_19230,N_19094);
xnor U21939 (N_21939,N_19294,N_19243);
nor U21940 (N_21940,N_19286,N_19203);
and U21941 (N_21941,N_19459,N_19851);
xnor U21942 (N_21942,N_18803,N_18238);
and U21943 (N_21943,N_18134,N_17702);
or U21944 (N_21944,N_17956,N_19711);
and U21945 (N_21945,N_18857,N_18825);
nand U21946 (N_21946,N_19953,N_19574);
or U21947 (N_21947,N_18718,N_17640);
and U21948 (N_21948,N_17619,N_17916);
or U21949 (N_21949,N_18126,N_18461);
xnor U21950 (N_21950,N_18093,N_17946);
and U21951 (N_21951,N_17715,N_19918);
and U21952 (N_21952,N_17599,N_19705);
xnor U21953 (N_21953,N_18464,N_18103);
or U21954 (N_21954,N_18034,N_19305);
xor U21955 (N_21955,N_19366,N_18000);
or U21956 (N_21956,N_19198,N_18133);
or U21957 (N_21957,N_18898,N_19877);
or U21958 (N_21958,N_17915,N_19175);
nor U21959 (N_21959,N_18852,N_19394);
or U21960 (N_21960,N_17859,N_17847);
or U21961 (N_21961,N_18635,N_19678);
nor U21962 (N_21962,N_19030,N_19588);
and U21963 (N_21963,N_18948,N_18475);
and U21964 (N_21964,N_19233,N_17815);
nor U21965 (N_21965,N_18081,N_19778);
or U21966 (N_21966,N_17543,N_19989);
and U21967 (N_21967,N_18149,N_19178);
xor U21968 (N_21968,N_17625,N_19538);
nor U21969 (N_21969,N_18324,N_19535);
or U21970 (N_21970,N_17929,N_19680);
xor U21971 (N_21971,N_19651,N_19767);
xnor U21972 (N_21972,N_19963,N_19337);
xor U21973 (N_21973,N_19716,N_18413);
and U21974 (N_21974,N_18434,N_18430);
or U21975 (N_21975,N_19470,N_18657);
or U21976 (N_21976,N_18998,N_19563);
and U21977 (N_21977,N_19162,N_18898);
and U21978 (N_21978,N_17899,N_19203);
and U21979 (N_21979,N_19905,N_19276);
nor U21980 (N_21980,N_19111,N_18096);
and U21981 (N_21981,N_18223,N_18785);
xor U21982 (N_21982,N_18112,N_19243);
nor U21983 (N_21983,N_18718,N_17687);
and U21984 (N_21984,N_19525,N_17615);
nor U21985 (N_21985,N_19047,N_18496);
and U21986 (N_21986,N_18310,N_18404);
xnor U21987 (N_21987,N_18711,N_19566);
nor U21988 (N_21988,N_19919,N_19239);
or U21989 (N_21989,N_19719,N_18793);
or U21990 (N_21990,N_19598,N_19176);
xnor U21991 (N_21991,N_19133,N_18881);
or U21992 (N_21992,N_18296,N_17568);
or U21993 (N_21993,N_19231,N_18747);
or U21994 (N_21994,N_19344,N_18567);
or U21995 (N_21995,N_17871,N_18516);
nor U21996 (N_21996,N_18025,N_18304);
nand U21997 (N_21997,N_19730,N_19567);
nor U21998 (N_21998,N_18131,N_19656);
xor U21999 (N_21999,N_19794,N_18746);
or U22000 (N_22000,N_19893,N_18419);
xor U22001 (N_22001,N_19637,N_18268);
nand U22002 (N_22002,N_19602,N_17974);
or U22003 (N_22003,N_17831,N_17871);
and U22004 (N_22004,N_19177,N_19666);
or U22005 (N_22005,N_18179,N_19366);
xor U22006 (N_22006,N_19739,N_19091);
nand U22007 (N_22007,N_18775,N_17815);
nand U22008 (N_22008,N_18601,N_18925);
nand U22009 (N_22009,N_19879,N_19023);
nand U22010 (N_22010,N_18455,N_18735);
xor U22011 (N_22011,N_19726,N_18360);
nand U22012 (N_22012,N_18740,N_17699);
or U22013 (N_22013,N_19977,N_19791);
nand U22014 (N_22014,N_18830,N_19587);
nor U22015 (N_22015,N_18279,N_18156);
nor U22016 (N_22016,N_17668,N_18247);
nand U22017 (N_22017,N_17969,N_19904);
nand U22018 (N_22018,N_19167,N_19700);
xnor U22019 (N_22019,N_18648,N_17799);
or U22020 (N_22020,N_18584,N_17981);
nor U22021 (N_22021,N_18150,N_18475);
and U22022 (N_22022,N_18304,N_19994);
or U22023 (N_22023,N_19592,N_18109);
or U22024 (N_22024,N_17740,N_19723);
xor U22025 (N_22025,N_19335,N_18849);
nor U22026 (N_22026,N_17744,N_19617);
nand U22027 (N_22027,N_17543,N_18539);
xor U22028 (N_22028,N_17935,N_19274);
nand U22029 (N_22029,N_17654,N_19668);
xor U22030 (N_22030,N_17507,N_19598);
nand U22031 (N_22031,N_19343,N_19860);
nor U22032 (N_22032,N_19663,N_19564);
or U22033 (N_22033,N_18102,N_17533);
xor U22034 (N_22034,N_19734,N_18527);
and U22035 (N_22035,N_17644,N_17914);
nor U22036 (N_22036,N_18953,N_18534);
or U22037 (N_22037,N_17827,N_17970);
or U22038 (N_22038,N_17994,N_18749);
or U22039 (N_22039,N_17648,N_17633);
and U22040 (N_22040,N_17607,N_17684);
or U22041 (N_22041,N_17719,N_18266);
and U22042 (N_22042,N_17735,N_17535);
xnor U22043 (N_22043,N_19000,N_17850);
nand U22044 (N_22044,N_17933,N_19997);
nand U22045 (N_22045,N_17640,N_17541);
or U22046 (N_22046,N_18335,N_19598);
or U22047 (N_22047,N_18418,N_18137);
nand U22048 (N_22048,N_19674,N_18747);
or U22049 (N_22049,N_18474,N_17547);
nor U22050 (N_22050,N_19703,N_17714);
or U22051 (N_22051,N_17602,N_19213);
or U22052 (N_22052,N_17700,N_18347);
and U22053 (N_22053,N_18187,N_17971);
nand U22054 (N_22054,N_19809,N_19090);
nor U22055 (N_22055,N_18688,N_19876);
nor U22056 (N_22056,N_17882,N_19702);
nand U22057 (N_22057,N_18482,N_18898);
or U22058 (N_22058,N_17838,N_19841);
nand U22059 (N_22059,N_17862,N_18363);
or U22060 (N_22060,N_19161,N_17781);
xor U22061 (N_22061,N_19828,N_17694);
and U22062 (N_22062,N_19737,N_19884);
xor U22063 (N_22063,N_18962,N_18720);
nor U22064 (N_22064,N_19211,N_19075);
nor U22065 (N_22065,N_18476,N_18648);
nand U22066 (N_22066,N_19631,N_19264);
or U22067 (N_22067,N_19555,N_19539);
nor U22068 (N_22068,N_18016,N_18856);
xor U22069 (N_22069,N_18588,N_17751);
xnor U22070 (N_22070,N_18096,N_18394);
nand U22071 (N_22071,N_19383,N_18228);
xor U22072 (N_22072,N_18025,N_19245);
nor U22073 (N_22073,N_18517,N_18820);
and U22074 (N_22074,N_19671,N_18753);
nand U22075 (N_22075,N_18078,N_18838);
or U22076 (N_22076,N_18681,N_19323);
and U22077 (N_22077,N_17893,N_19592);
nor U22078 (N_22078,N_19259,N_18720);
xor U22079 (N_22079,N_19058,N_19078);
xnor U22080 (N_22080,N_19491,N_19024);
or U22081 (N_22081,N_19060,N_19357);
or U22082 (N_22082,N_17520,N_18627);
xnor U22083 (N_22083,N_19564,N_19333);
nand U22084 (N_22084,N_19869,N_18224);
nor U22085 (N_22085,N_18433,N_18261);
nor U22086 (N_22086,N_19963,N_18107);
and U22087 (N_22087,N_19221,N_18989);
nor U22088 (N_22088,N_19377,N_19663);
xor U22089 (N_22089,N_19935,N_18291);
xor U22090 (N_22090,N_17729,N_19990);
or U22091 (N_22091,N_19920,N_19148);
nor U22092 (N_22092,N_17819,N_18038);
nand U22093 (N_22093,N_17667,N_18471);
nor U22094 (N_22094,N_18207,N_18474);
xor U22095 (N_22095,N_18731,N_17702);
nor U22096 (N_22096,N_19452,N_17503);
and U22097 (N_22097,N_17686,N_19452);
xor U22098 (N_22098,N_18522,N_19185);
and U22099 (N_22099,N_18001,N_19223);
or U22100 (N_22100,N_19476,N_19141);
and U22101 (N_22101,N_18798,N_17551);
or U22102 (N_22102,N_18024,N_17928);
xor U22103 (N_22103,N_19640,N_19004);
nand U22104 (N_22104,N_19451,N_18829);
nor U22105 (N_22105,N_18404,N_17677);
nand U22106 (N_22106,N_19487,N_17593);
nand U22107 (N_22107,N_19807,N_19044);
nand U22108 (N_22108,N_19947,N_17773);
nand U22109 (N_22109,N_17577,N_17586);
nand U22110 (N_22110,N_19805,N_19824);
and U22111 (N_22111,N_18301,N_19986);
and U22112 (N_22112,N_19368,N_19714);
xnor U22113 (N_22113,N_19705,N_18420);
nand U22114 (N_22114,N_19172,N_18340);
xor U22115 (N_22115,N_19723,N_19637);
nor U22116 (N_22116,N_17720,N_19442);
nor U22117 (N_22117,N_18141,N_19792);
xnor U22118 (N_22118,N_18423,N_19956);
nor U22119 (N_22119,N_18632,N_18707);
and U22120 (N_22120,N_19700,N_18630);
nand U22121 (N_22121,N_17918,N_19380);
xnor U22122 (N_22122,N_17501,N_18257);
nor U22123 (N_22123,N_19298,N_19837);
nor U22124 (N_22124,N_18649,N_18078);
nand U22125 (N_22125,N_18196,N_18471);
or U22126 (N_22126,N_19394,N_19653);
or U22127 (N_22127,N_18306,N_18588);
or U22128 (N_22128,N_19273,N_17938);
nor U22129 (N_22129,N_19885,N_19896);
or U22130 (N_22130,N_19332,N_18569);
nor U22131 (N_22131,N_19847,N_19564);
or U22132 (N_22132,N_19313,N_18650);
nor U22133 (N_22133,N_18901,N_17851);
xnor U22134 (N_22134,N_19579,N_19520);
nor U22135 (N_22135,N_19790,N_19297);
nor U22136 (N_22136,N_18944,N_19362);
nor U22137 (N_22137,N_17588,N_19445);
xor U22138 (N_22138,N_18306,N_17949);
and U22139 (N_22139,N_19267,N_17577);
xor U22140 (N_22140,N_18615,N_19339);
nand U22141 (N_22141,N_17507,N_19091);
nand U22142 (N_22142,N_19065,N_19352);
nand U22143 (N_22143,N_18126,N_18125);
nand U22144 (N_22144,N_18256,N_17916);
or U22145 (N_22145,N_17923,N_19826);
nand U22146 (N_22146,N_17611,N_19718);
and U22147 (N_22147,N_17839,N_18046);
xnor U22148 (N_22148,N_17825,N_18750);
xnor U22149 (N_22149,N_19374,N_18659);
xnor U22150 (N_22150,N_18598,N_19903);
or U22151 (N_22151,N_19124,N_19415);
or U22152 (N_22152,N_17511,N_18943);
nand U22153 (N_22153,N_19470,N_18618);
xor U22154 (N_22154,N_18838,N_18088);
nor U22155 (N_22155,N_18443,N_19085);
xnor U22156 (N_22156,N_19227,N_19266);
or U22157 (N_22157,N_19588,N_19389);
nand U22158 (N_22158,N_18774,N_18745);
or U22159 (N_22159,N_19838,N_19318);
nand U22160 (N_22160,N_18485,N_19754);
or U22161 (N_22161,N_19060,N_18149);
and U22162 (N_22162,N_19214,N_18506);
nor U22163 (N_22163,N_17748,N_18763);
or U22164 (N_22164,N_19502,N_18867);
nand U22165 (N_22165,N_19206,N_18497);
or U22166 (N_22166,N_18283,N_18413);
nor U22167 (N_22167,N_18528,N_18208);
xnor U22168 (N_22168,N_18579,N_19339);
nor U22169 (N_22169,N_18829,N_18093);
and U22170 (N_22170,N_18854,N_19384);
xor U22171 (N_22171,N_19131,N_18977);
and U22172 (N_22172,N_17750,N_18194);
xor U22173 (N_22173,N_17790,N_18398);
or U22174 (N_22174,N_17973,N_18542);
nor U22175 (N_22175,N_18176,N_17636);
or U22176 (N_22176,N_18946,N_17961);
nand U22177 (N_22177,N_17937,N_18324);
or U22178 (N_22178,N_18214,N_17761);
or U22179 (N_22179,N_19575,N_19507);
and U22180 (N_22180,N_17707,N_18317);
xor U22181 (N_22181,N_17592,N_18048);
xor U22182 (N_22182,N_17897,N_17576);
and U22183 (N_22183,N_17696,N_18882);
or U22184 (N_22184,N_18600,N_19734);
nand U22185 (N_22185,N_18327,N_19127);
nor U22186 (N_22186,N_19099,N_19809);
and U22187 (N_22187,N_19960,N_17902);
and U22188 (N_22188,N_19781,N_19973);
nand U22189 (N_22189,N_18954,N_17587);
xnor U22190 (N_22190,N_17502,N_19953);
or U22191 (N_22191,N_19895,N_18216);
xnor U22192 (N_22192,N_17720,N_18044);
xor U22193 (N_22193,N_17799,N_19634);
nor U22194 (N_22194,N_19692,N_18292);
and U22195 (N_22195,N_19763,N_17677);
nor U22196 (N_22196,N_18321,N_18472);
nor U22197 (N_22197,N_19267,N_18133);
and U22198 (N_22198,N_19186,N_18775);
and U22199 (N_22199,N_17900,N_19916);
and U22200 (N_22200,N_19835,N_18878);
and U22201 (N_22201,N_18241,N_18900);
and U22202 (N_22202,N_19693,N_18934);
nand U22203 (N_22203,N_19508,N_18524);
and U22204 (N_22204,N_18355,N_19514);
nor U22205 (N_22205,N_19026,N_18468);
nand U22206 (N_22206,N_18105,N_19359);
and U22207 (N_22207,N_17844,N_18767);
nand U22208 (N_22208,N_18463,N_18390);
xnor U22209 (N_22209,N_17874,N_19917);
and U22210 (N_22210,N_19662,N_18921);
or U22211 (N_22211,N_19154,N_19102);
and U22212 (N_22212,N_19597,N_19260);
or U22213 (N_22213,N_19349,N_17695);
nor U22214 (N_22214,N_18132,N_18235);
xor U22215 (N_22215,N_18377,N_19108);
or U22216 (N_22216,N_18258,N_19969);
or U22217 (N_22217,N_18465,N_19165);
xor U22218 (N_22218,N_19847,N_18596);
nor U22219 (N_22219,N_17835,N_17672);
nand U22220 (N_22220,N_18795,N_19316);
or U22221 (N_22221,N_17716,N_17527);
xnor U22222 (N_22222,N_19571,N_19393);
nand U22223 (N_22223,N_17813,N_18107);
nand U22224 (N_22224,N_18258,N_18540);
nor U22225 (N_22225,N_19042,N_17660);
or U22226 (N_22226,N_18873,N_18929);
nand U22227 (N_22227,N_19111,N_19104);
or U22228 (N_22228,N_17929,N_18341);
nor U22229 (N_22229,N_18756,N_18647);
nand U22230 (N_22230,N_18395,N_19044);
nand U22231 (N_22231,N_19836,N_19227);
xnor U22232 (N_22232,N_19406,N_19021);
and U22233 (N_22233,N_18044,N_18602);
xnor U22234 (N_22234,N_18362,N_19882);
nor U22235 (N_22235,N_18521,N_18168);
nor U22236 (N_22236,N_19557,N_18909);
xor U22237 (N_22237,N_17666,N_19447);
xor U22238 (N_22238,N_17563,N_18470);
and U22239 (N_22239,N_18777,N_17833);
nand U22240 (N_22240,N_18319,N_19116);
nand U22241 (N_22241,N_19643,N_18529);
or U22242 (N_22242,N_18703,N_18824);
nand U22243 (N_22243,N_18662,N_18132);
nor U22244 (N_22244,N_17747,N_18405);
or U22245 (N_22245,N_18828,N_18879);
or U22246 (N_22246,N_19755,N_17985);
nand U22247 (N_22247,N_18835,N_18322);
and U22248 (N_22248,N_18210,N_19326);
xnor U22249 (N_22249,N_18790,N_19679);
nand U22250 (N_22250,N_18493,N_19775);
nor U22251 (N_22251,N_17622,N_17796);
nor U22252 (N_22252,N_17999,N_18965);
nor U22253 (N_22253,N_19882,N_18459);
nor U22254 (N_22254,N_18581,N_19921);
or U22255 (N_22255,N_19872,N_19597);
or U22256 (N_22256,N_18932,N_19098);
and U22257 (N_22257,N_19349,N_18319);
nand U22258 (N_22258,N_18012,N_19225);
and U22259 (N_22259,N_19984,N_19318);
and U22260 (N_22260,N_17567,N_18375);
and U22261 (N_22261,N_19579,N_18433);
and U22262 (N_22262,N_17678,N_19162);
xnor U22263 (N_22263,N_19950,N_17907);
xnor U22264 (N_22264,N_17814,N_17801);
nor U22265 (N_22265,N_18307,N_18261);
or U22266 (N_22266,N_18284,N_18763);
nor U22267 (N_22267,N_17875,N_18015);
or U22268 (N_22268,N_17738,N_18642);
nor U22269 (N_22269,N_19280,N_18992);
nor U22270 (N_22270,N_19463,N_19946);
xor U22271 (N_22271,N_19007,N_18622);
or U22272 (N_22272,N_18264,N_18656);
xor U22273 (N_22273,N_19662,N_18125);
or U22274 (N_22274,N_18778,N_17612);
nand U22275 (N_22275,N_18076,N_17661);
and U22276 (N_22276,N_19265,N_18027);
nand U22277 (N_22277,N_17747,N_17830);
or U22278 (N_22278,N_18196,N_19476);
xor U22279 (N_22279,N_18594,N_19030);
or U22280 (N_22280,N_17529,N_19690);
nand U22281 (N_22281,N_17899,N_19104);
or U22282 (N_22282,N_19826,N_18195);
or U22283 (N_22283,N_17579,N_19471);
and U22284 (N_22284,N_19216,N_19235);
xor U22285 (N_22285,N_17554,N_18880);
nor U22286 (N_22286,N_19871,N_19803);
nand U22287 (N_22287,N_18055,N_18924);
xor U22288 (N_22288,N_18653,N_18164);
and U22289 (N_22289,N_18173,N_18076);
and U22290 (N_22290,N_18410,N_18916);
nand U22291 (N_22291,N_19651,N_18125);
and U22292 (N_22292,N_17809,N_19610);
or U22293 (N_22293,N_19738,N_17972);
xnor U22294 (N_22294,N_19825,N_17960);
nand U22295 (N_22295,N_18903,N_18093);
or U22296 (N_22296,N_19808,N_17723);
and U22297 (N_22297,N_18435,N_19775);
nand U22298 (N_22298,N_18094,N_18196);
xor U22299 (N_22299,N_19344,N_19721);
or U22300 (N_22300,N_18445,N_18014);
xor U22301 (N_22301,N_17985,N_19252);
nand U22302 (N_22302,N_19091,N_18910);
nor U22303 (N_22303,N_18510,N_17703);
xnor U22304 (N_22304,N_19227,N_19994);
nor U22305 (N_22305,N_18299,N_19809);
xor U22306 (N_22306,N_19891,N_18810);
or U22307 (N_22307,N_19140,N_17611);
nor U22308 (N_22308,N_18723,N_17501);
and U22309 (N_22309,N_19248,N_19500);
or U22310 (N_22310,N_17873,N_19242);
nand U22311 (N_22311,N_18896,N_19744);
xnor U22312 (N_22312,N_17658,N_18431);
nand U22313 (N_22313,N_17961,N_18121);
nand U22314 (N_22314,N_18976,N_19005);
xor U22315 (N_22315,N_18622,N_17721);
nor U22316 (N_22316,N_17514,N_18376);
nor U22317 (N_22317,N_19516,N_18190);
nand U22318 (N_22318,N_18308,N_18279);
xor U22319 (N_22319,N_19055,N_18959);
nor U22320 (N_22320,N_18469,N_18295);
nand U22321 (N_22321,N_18458,N_17571);
nand U22322 (N_22322,N_19826,N_19422);
and U22323 (N_22323,N_19344,N_18819);
nand U22324 (N_22324,N_18879,N_18840);
or U22325 (N_22325,N_18310,N_19342);
nor U22326 (N_22326,N_19327,N_17785);
and U22327 (N_22327,N_18434,N_19248);
or U22328 (N_22328,N_18094,N_19912);
nor U22329 (N_22329,N_18125,N_19643);
xor U22330 (N_22330,N_18761,N_18417);
xnor U22331 (N_22331,N_19111,N_18326);
xor U22332 (N_22332,N_19823,N_19214);
nor U22333 (N_22333,N_17726,N_19996);
xor U22334 (N_22334,N_18784,N_19513);
nor U22335 (N_22335,N_19858,N_18314);
nor U22336 (N_22336,N_18189,N_18784);
nor U22337 (N_22337,N_19370,N_18928);
and U22338 (N_22338,N_18079,N_19365);
and U22339 (N_22339,N_19745,N_19524);
nor U22340 (N_22340,N_18579,N_18678);
nand U22341 (N_22341,N_19644,N_19945);
nand U22342 (N_22342,N_18792,N_17632);
nand U22343 (N_22343,N_19228,N_19841);
and U22344 (N_22344,N_18977,N_17612);
and U22345 (N_22345,N_19940,N_18091);
and U22346 (N_22346,N_19166,N_19616);
or U22347 (N_22347,N_18496,N_18594);
nand U22348 (N_22348,N_18315,N_19958);
nor U22349 (N_22349,N_18752,N_17933);
nand U22350 (N_22350,N_18185,N_17821);
nor U22351 (N_22351,N_19130,N_19610);
and U22352 (N_22352,N_19675,N_18574);
or U22353 (N_22353,N_18929,N_19064);
and U22354 (N_22354,N_17766,N_19078);
or U22355 (N_22355,N_17994,N_19240);
or U22356 (N_22356,N_19407,N_17886);
and U22357 (N_22357,N_18377,N_17992);
nand U22358 (N_22358,N_18015,N_17828);
or U22359 (N_22359,N_17957,N_17583);
nand U22360 (N_22360,N_18171,N_18005);
xor U22361 (N_22361,N_19698,N_18893);
xnor U22362 (N_22362,N_18513,N_17632);
nor U22363 (N_22363,N_18794,N_19391);
xnor U22364 (N_22364,N_18544,N_19859);
nand U22365 (N_22365,N_17714,N_19458);
xnor U22366 (N_22366,N_17652,N_19817);
or U22367 (N_22367,N_18377,N_18283);
nand U22368 (N_22368,N_18534,N_19042);
and U22369 (N_22369,N_17580,N_19022);
nor U22370 (N_22370,N_19847,N_18817);
nand U22371 (N_22371,N_18456,N_18669);
or U22372 (N_22372,N_17683,N_18383);
xnor U22373 (N_22373,N_19551,N_19120);
nor U22374 (N_22374,N_18496,N_18958);
xor U22375 (N_22375,N_18621,N_18348);
nand U22376 (N_22376,N_19283,N_18007);
nor U22377 (N_22377,N_19355,N_18884);
nand U22378 (N_22378,N_19524,N_17696);
xnor U22379 (N_22379,N_18391,N_18878);
xor U22380 (N_22380,N_18725,N_19207);
nand U22381 (N_22381,N_19011,N_17786);
nand U22382 (N_22382,N_18289,N_19690);
nor U22383 (N_22383,N_19909,N_18357);
xnor U22384 (N_22384,N_19884,N_18691);
and U22385 (N_22385,N_19513,N_18496);
nor U22386 (N_22386,N_18346,N_19485);
and U22387 (N_22387,N_19221,N_19021);
xor U22388 (N_22388,N_19451,N_18347);
or U22389 (N_22389,N_19599,N_18531);
nor U22390 (N_22390,N_18147,N_18997);
nor U22391 (N_22391,N_18923,N_19673);
or U22392 (N_22392,N_19353,N_17885);
or U22393 (N_22393,N_19702,N_19233);
or U22394 (N_22394,N_18666,N_19955);
nor U22395 (N_22395,N_19668,N_18097);
or U22396 (N_22396,N_18131,N_17649);
and U22397 (N_22397,N_18398,N_19058);
nand U22398 (N_22398,N_18017,N_18844);
or U22399 (N_22399,N_18152,N_17776);
xnor U22400 (N_22400,N_18793,N_18535);
nor U22401 (N_22401,N_17784,N_19564);
and U22402 (N_22402,N_18311,N_17778);
and U22403 (N_22403,N_18688,N_18037);
xor U22404 (N_22404,N_19781,N_17692);
or U22405 (N_22405,N_17751,N_19549);
or U22406 (N_22406,N_18821,N_18382);
or U22407 (N_22407,N_18748,N_19906);
or U22408 (N_22408,N_17917,N_17519);
xor U22409 (N_22409,N_18199,N_18267);
nand U22410 (N_22410,N_19673,N_18694);
nand U22411 (N_22411,N_19496,N_18337);
nor U22412 (N_22412,N_18003,N_19212);
nand U22413 (N_22413,N_19345,N_17507);
nand U22414 (N_22414,N_18765,N_18882);
nand U22415 (N_22415,N_18490,N_17621);
nand U22416 (N_22416,N_18595,N_17553);
and U22417 (N_22417,N_19200,N_19345);
xor U22418 (N_22418,N_19122,N_19105);
and U22419 (N_22419,N_17906,N_19670);
nand U22420 (N_22420,N_18973,N_18011);
or U22421 (N_22421,N_19044,N_19814);
nand U22422 (N_22422,N_17782,N_19682);
nand U22423 (N_22423,N_18390,N_19881);
xnor U22424 (N_22424,N_19716,N_18364);
nand U22425 (N_22425,N_19371,N_17923);
and U22426 (N_22426,N_18579,N_19522);
xor U22427 (N_22427,N_19412,N_18367);
or U22428 (N_22428,N_17891,N_18232);
and U22429 (N_22429,N_19493,N_19514);
and U22430 (N_22430,N_18530,N_18750);
xnor U22431 (N_22431,N_19199,N_18939);
nand U22432 (N_22432,N_19238,N_19565);
nand U22433 (N_22433,N_17820,N_18614);
and U22434 (N_22434,N_17747,N_18942);
nand U22435 (N_22435,N_19458,N_17761);
xor U22436 (N_22436,N_19206,N_18147);
nand U22437 (N_22437,N_17702,N_17995);
or U22438 (N_22438,N_18668,N_19309);
nor U22439 (N_22439,N_18540,N_18927);
or U22440 (N_22440,N_17679,N_19074);
or U22441 (N_22441,N_19984,N_18303);
xnor U22442 (N_22442,N_19815,N_19240);
xor U22443 (N_22443,N_19368,N_18197);
nor U22444 (N_22444,N_19234,N_19232);
or U22445 (N_22445,N_19860,N_18974);
nand U22446 (N_22446,N_18055,N_18017);
or U22447 (N_22447,N_17698,N_19375);
and U22448 (N_22448,N_17902,N_19041);
and U22449 (N_22449,N_19989,N_18141);
or U22450 (N_22450,N_17560,N_17656);
xor U22451 (N_22451,N_18357,N_18962);
or U22452 (N_22452,N_19310,N_18270);
nand U22453 (N_22453,N_18025,N_18108);
or U22454 (N_22454,N_18689,N_18929);
or U22455 (N_22455,N_18794,N_18670);
nor U22456 (N_22456,N_17633,N_17854);
nand U22457 (N_22457,N_18322,N_18847);
nand U22458 (N_22458,N_18030,N_19650);
nand U22459 (N_22459,N_18011,N_18946);
xor U22460 (N_22460,N_18399,N_19836);
xor U22461 (N_22461,N_19373,N_19414);
or U22462 (N_22462,N_17542,N_18758);
or U22463 (N_22463,N_17759,N_19140);
nand U22464 (N_22464,N_18090,N_19489);
or U22465 (N_22465,N_17838,N_17819);
nand U22466 (N_22466,N_17514,N_19584);
and U22467 (N_22467,N_19132,N_19883);
nand U22468 (N_22468,N_18247,N_17792);
or U22469 (N_22469,N_19467,N_19987);
nand U22470 (N_22470,N_18454,N_17607);
and U22471 (N_22471,N_19902,N_18029);
nor U22472 (N_22472,N_17742,N_18833);
or U22473 (N_22473,N_19196,N_18414);
or U22474 (N_22474,N_17613,N_19968);
nand U22475 (N_22475,N_19075,N_18818);
xor U22476 (N_22476,N_18474,N_19725);
nand U22477 (N_22477,N_18509,N_18132);
and U22478 (N_22478,N_17576,N_18490);
nand U22479 (N_22479,N_18421,N_19533);
xnor U22480 (N_22480,N_19691,N_18943);
and U22481 (N_22481,N_18222,N_19079);
xnor U22482 (N_22482,N_18829,N_19060);
nand U22483 (N_22483,N_18575,N_19986);
nor U22484 (N_22484,N_17582,N_19763);
xnor U22485 (N_22485,N_19062,N_17788);
xor U22486 (N_22486,N_17640,N_17963);
nor U22487 (N_22487,N_17613,N_18670);
or U22488 (N_22488,N_18535,N_19059);
and U22489 (N_22489,N_18637,N_19285);
nor U22490 (N_22490,N_19325,N_19333);
or U22491 (N_22491,N_17716,N_19271);
nand U22492 (N_22492,N_19280,N_18946);
nand U22493 (N_22493,N_18100,N_19699);
nand U22494 (N_22494,N_17890,N_19310);
nand U22495 (N_22495,N_18927,N_19526);
xor U22496 (N_22496,N_17969,N_19799);
and U22497 (N_22497,N_19079,N_19525);
nand U22498 (N_22498,N_19307,N_18314);
nand U22499 (N_22499,N_19740,N_17670);
nand U22500 (N_22500,N_21770,N_20352);
and U22501 (N_22501,N_22132,N_20966);
nand U22502 (N_22502,N_20892,N_20686);
xor U22503 (N_22503,N_21864,N_21161);
xnor U22504 (N_22504,N_21254,N_21337);
or U22505 (N_22505,N_21899,N_20429);
and U22506 (N_22506,N_21904,N_22306);
nand U22507 (N_22507,N_20244,N_21397);
nor U22508 (N_22508,N_21614,N_21643);
and U22509 (N_22509,N_22287,N_22234);
or U22510 (N_22510,N_21192,N_22101);
or U22511 (N_22511,N_21407,N_20665);
nor U22512 (N_22512,N_20375,N_20838);
and U22513 (N_22513,N_21937,N_21227);
or U22514 (N_22514,N_20197,N_20868);
and U22515 (N_22515,N_21394,N_20062);
nand U22516 (N_22516,N_21859,N_21135);
and U22517 (N_22517,N_21054,N_22353);
xor U22518 (N_22518,N_22417,N_21076);
xor U22519 (N_22519,N_20130,N_21528);
or U22520 (N_22520,N_22313,N_21431);
nand U22521 (N_22521,N_22424,N_20186);
and U22522 (N_22522,N_20345,N_22314);
nor U22523 (N_22523,N_20199,N_20543);
xnor U22524 (N_22524,N_21711,N_21312);
xor U22525 (N_22525,N_21663,N_21068);
nand U22526 (N_22526,N_22401,N_20024);
or U22527 (N_22527,N_21748,N_21629);
nor U22528 (N_22528,N_20235,N_20783);
and U22529 (N_22529,N_20029,N_21644);
and U22530 (N_22530,N_22474,N_20627);
nand U22531 (N_22531,N_20717,N_20081);
and U22532 (N_22532,N_21561,N_21522);
nand U22533 (N_22533,N_21044,N_21707);
nor U22534 (N_22534,N_20516,N_20467);
nand U22535 (N_22535,N_21545,N_20877);
and U22536 (N_22536,N_20441,N_20419);
nand U22537 (N_22537,N_20159,N_20573);
xnor U22538 (N_22538,N_22260,N_20597);
and U22539 (N_22539,N_20889,N_21700);
nand U22540 (N_22540,N_20472,N_20263);
xor U22541 (N_22541,N_21300,N_20378);
xnor U22542 (N_22542,N_20604,N_20797);
and U22543 (N_22543,N_20387,N_22099);
nand U22544 (N_22544,N_21327,N_21040);
xor U22545 (N_22545,N_21001,N_20401);
nor U22546 (N_22546,N_21553,N_21396);
or U22547 (N_22547,N_20363,N_21325);
xnor U22548 (N_22548,N_20914,N_20567);
xnor U22549 (N_22549,N_22043,N_20924);
and U22550 (N_22550,N_22094,N_20121);
nor U22551 (N_22551,N_21087,N_22255);
or U22552 (N_22552,N_21538,N_20246);
or U22553 (N_22553,N_21977,N_20942);
and U22554 (N_22554,N_21334,N_21570);
nand U22555 (N_22555,N_20257,N_20476);
nand U22556 (N_22556,N_22139,N_20430);
or U22557 (N_22557,N_20652,N_22217);
nor U22558 (N_22558,N_22237,N_22449);
nand U22559 (N_22559,N_20954,N_20997);
and U22560 (N_22560,N_21143,N_21437);
nand U22561 (N_22561,N_21781,N_21563);
nor U22562 (N_22562,N_20798,N_20007);
nor U22563 (N_22563,N_20591,N_21210);
and U22564 (N_22564,N_20465,N_21406);
and U22565 (N_22565,N_22177,N_20583);
and U22566 (N_22566,N_20044,N_22366);
xor U22567 (N_22567,N_20497,N_21526);
xor U22568 (N_22568,N_20642,N_22315);
nor U22569 (N_22569,N_21595,N_20564);
xnor U22570 (N_22570,N_21688,N_20874);
nor U22571 (N_22571,N_21322,N_21400);
or U22572 (N_22572,N_22161,N_21024);
or U22573 (N_22573,N_22453,N_20643);
and U22574 (N_22574,N_22076,N_20850);
or U22575 (N_22575,N_21370,N_20648);
and U22576 (N_22576,N_21666,N_21647);
nor U22577 (N_22577,N_22324,N_21673);
and U22578 (N_22578,N_20177,N_21232);
or U22579 (N_22579,N_20766,N_20703);
xnor U22580 (N_22580,N_20618,N_21457);
nand U22581 (N_22581,N_20106,N_21415);
xor U22582 (N_22582,N_20391,N_22395);
or U22583 (N_22583,N_21664,N_21131);
xor U22584 (N_22584,N_21788,N_21336);
nor U22585 (N_22585,N_21785,N_21980);
nor U22586 (N_22586,N_21955,N_21819);
nand U22587 (N_22587,N_22320,N_20948);
or U22588 (N_22588,N_20520,N_22151);
nor U22589 (N_22589,N_20833,N_21361);
nand U22590 (N_22590,N_20771,N_21066);
xnor U22591 (N_22591,N_20861,N_22272);
nand U22592 (N_22592,N_22096,N_22204);
and U22593 (N_22593,N_20899,N_20370);
and U22594 (N_22594,N_20041,N_20935);
nand U22595 (N_22595,N_20851,N_20232);
xnor U22596 (N_22596,N_20316,N_21467);
or U22597 (N_22597,N_22201,N_22456);
and U22598 (N_22598,N_21963,N_21498);
nor U22599 (N_22599,N_22238,N_21591);
or U22600 (N_22600,N_20545,N_20014);
nor U22601 (N_22601,N_21418,N_20485);
nor U22602 (N_22602,N_21543,N_20949);
xor U22603 (N_22603,N_22061,N_22082);
xnor U22604 (N_22604,N_21836,N_20112);
and U22605 (N_22605,N_20353,N_22390);
and U22606 (N_22606,N_22239,N_20697);
nor U22607 (N_22607,N_21927,N_22440);
nor U22608 (N_22608,N_20416,N_22023);
or U22609 (N_22609,N_21912,N_20158);
and U22610 (N_22610,N_21520,N_21913);
nand U22611 (N_22611,N_20625,N_20817);
nand U22612 (N_22612,N_20418,N_22307);
nor U22613 (N_22613,N_22131,N_20253);
nand U22614 (N_22614,N_21798,N_22466);
nor U22615 (N_22615,N_20623,N_21569);
nor U22616 (N_22616,N_20547,N_22142);
xor U22617 (N_22617,N_21975,N_21189);
nor U22618 (N_22618,N_20038,N_20068);
nand U22619 (N_22619,N_21659,N_20109);
nand U22620 (N_22620,N_20426,N_20488);
and U22621 (N_22621,N_20337,N_22229);
and U22622 (N_22622,N_20349,N_20801);
nor U22623 (N_22623,N_20982,N_20367);
xor U22624 (N_22624,N_21079,N_20614);
nor U22625 (N_22625,N_20981,N_20331);
nand U22626 (N_22626,N_22304,N_21309);
and U22627 (N_22627,N_21314,N_22410);
nor U22628 (N_22628,N_22167,N_22492);
or U22629 (N_22629,N_21324,N_22310);
nor U22630 (N_22630,N_21482,N_20509);
nand U22631 (N_22631,N_21206,N_21814);
and U22632 (N_22632,N_21170,N_22067);
and U22633 (N_22633,N_22467,N_21662);
and U22634 (N_22634,N_22357,N_20167);
nand U22635 (N_22635,N_20905,N_20763);
or U22636 (N_22636,N_20513,N_22035);
xor U22637 (N_22637,N_20818,N_21514);
nand U22638 (N_22638,N_21136,N_21997);
nor U22639 (N_22639,N_20535,N_21989);
and U22640 (N_22640,N_20983,N_20538);
or U22641 (N_22641,N_21637,N_22233);
nor U22642 (N_22642,N_21320,N_21617);
and U22643 (N_22643,N_20719,N_21758);
and U22644 (N_22644,N_22321,N_20428);
nor U22645 (N_22645,N_20596,N_20380);
and U22646 (N_22646,N_21171,N_21871);
xnor U22647 (N_22647,N_21439,N_22258);
nor U22648 (N_22648,N_21884,N_20501);
or U22649 (N_22649,N_21472,N_20593);
nand U22650 (N_22650,N_21088,N_20313);
nor U22651 (N_22651,N_22343,N_22044);
nor U22652 (N_22652,N_21133,N_20289);
or U22653 (N_22653,N_22352,N_20929);
nor U22654 (N_22654,N_22015,N_22326);
and U22655 (N_22655,N_20631,N_22499);
nand U22656 (N_22656,N_21845,N_20694);
nor U22657 (N_22657,N_20031,N_20863);
nand U22658 (N_22658,N_21060,N_21897);
nand U22659 (N_22659,N_20039,N_20339);
and U22660 (N_22660,N_22460,N_20882);
or U22661 (N_22661,N_21584,N_22316);
xnor U22662 (N_22662,N_20640,N_20032);
xnor U22663 (N_22663,N_20052,N_21960);
nor U22664 (N_22664,N_20125,N_20386);
xnor U22665 (N_22665,N_21841,N_20055);
or U22666 (N_22666,N_20434,N_20579);
and U22667 (N_22667,N_21110,N_22379);
nor U22668 (N_22668,N_20210,N_22329);
xnor U22669 (N_22669,N_22104,N_20563);
and U22670 (N_22670,N_21012,N_20713);
xnor U22671 (N_22671,N_22214,N_22488);
xnor U22672 (N_22672,N_21120,N_21633);
or U22673 (N_22673,N_20211,N_21154);
nor U22674 (N_22674,N_20710,N_20938);
xor U22675 (N_22675,N_20169,N_20328);
nor U22676 (N_22676,N_20736,N_20468);
xor U22677 (N_22677,N_20036,N_22108);
and U22678 (N_22678,N_21441,N_21548);
xor U22679 (N_22679,N_20973,N_21657);
or U22680 (N_22680,N_20681,N_22382);
and U22681 (N_22681,N_20421,N_20928);
and U22682 (N_22682,N_21346,N_22374);
nand U22683 (N_22683,N_20553,N_21566);
or U22684 (N_22684,N_22309,N_22236);
and U22685 (N_22685,N_20699,N_22259);
nand U22686 (N_22686,N_21444,N_21501);
nor U22687 (N_22687,N_20012,N_20056);
and U22688 (N_22688,N_22001,N_20084);
or U22689 (N_22689,N_20306,N_22019);
or U22690 (N_22690,N_21075,N_20654);
xor U22691 (N_22691,N_21261,N_20342);
or U22692 (N_22692,N_21687,N_21646);
and U22693 (N_22693,N_22426,N_22286);
or U22694 (N_22694,N_22459,N_20915);
nand U22695 (N_22695,N_21275,N_22418);
and U22696 (N_22696,N_21486,N_21402);
nor U22697 (N_22697,N_20389,N_20114);
nor U22698 (N_22698,N_21703,N_20296);
or U22699 (N_22699,N_20941,N_21029);
xor U22700 (N_22700,N_22389,N_20198);
xor U22701 (N_22701,N_22271,N_21847);
and U22702 (N_22702,N_21768,N_21696);
and U22703 (N_22703,N_21948,N_21456);
nand U22704 (N_22704,N_21806,N_20303);
or U22705 (N_22705,N_20178,N_22435);
xnor U22706 (N_22706,N_21235,N_21010);
nor U22707 (N_22707,N_21055,N_21086);
and U22708 (N_22708,N_21215,N_21429);
xnor U22709 (N_22709,N_21592,N_20063);
nand U22710 (N_22710,N_21984,N_22241);
xor U22711 (N_22711,N_20917,N_21926);
and U22712 (N_22712,N_21811,N_21541);
xor U22713 (N_22713,N_21784,N_21670);
nand U22714 (N_22714,N_21917,N_21253);
nand U22715 (N_22715,N_21698,N_21350);
nor U22716 (N_22716,N_21554,N_20976);
and U22717 (N_22717,N_20778,N_21160);
or U22718 (N_22718,N_20858,N_20165);
nor U22719 (N_22719,N_20500,N_22288);
or U22720 (N_22720,N_20598,N_21387);
or U22721 (N_22721,N_22039,N_20629);
and U22722 (N_22722,N_20011,N_20463);
nand U22723 (N_22723,N_20536,N_21114);
and U22724 (N_22724,N_21578,N_22185);
and U22725 (N_22725,N_20191,N_21523);
or U22726 (N_22726,N_20558,N_21477);
or U22727 (N_22727,N_20984,N_21460);
and U22728 (N_22728,N_20700,N_20279);
and U22729 (N_22729,N_22330,N_21855);
and U22730 (N_22730,N_22191,N_21985);
and U22731 (N_22731,N_20883,N_20462);
and U22732 (N_22732,N_20847,N_20385);
nand U22733 (N_22733,N_20330,N_21945);
xnor U22734 (N_22734,N_20124,N_21550);
nand U22735 (N_22735,N_21485,N_20921);
nand U22736 (N_22736,N_21064,N_22432);
xor U22737 (N_22737,N_20885,N_22222);
xor U22738 (N_22738,N_20131,N_21179);
xnor U22739 (N_22739,N_21159,N_21112);
nor U22740 (N_22740,N_20264,N_21347);
xor U22741 (N_22741,N_20356,N_21838);
and U22742 (N_22742,N_21727,N_22494);
xnor U22743 (N_22743,N_21676,N_21842);
nand U22744 (N_22744,N_20927,N_21108);
and U22745 (N_22745,N_20280,N_21279);
nand U22746 (N_22746,N_20317,N_21754);
and U22747 (N_22747,N_20826,N_21729);
nand U22748 (N_22748,N_21900,N_21500);
xnor U22749 (N_22749,N_20967,N_20053);
or U22750 (N_22750,N_21983,N_20205);
and U22751 (N_22751,N_20533,N_20823);
xnor U22752 (N_22752,N_21411,N_22053);
xor U22753 (N_22753,N_20361,N_21893);
or U22754 (N_22754,N_20276,N_22373);
or U22755 (N_22755,N_22136,N_21326);
and U22756 (N_22756,N_20379,N_21533);
and U22757 (N_22757,N_21162,N_20423);
and U22758 (N_22758,N_22468,N_20212);
nand U22759 (N_22759,N_21011,N_21311);
nand U22760 (N_22760,N_22338,N_20852);
nor U22761 (N_22761,N_20947,N_21328);
nor U22762 (N_22762,N_20505,N_21780);
nand U22763 (N_22763,N_21084,N_20839);
nand U22764 (N_22764,N_21832,N_22482);
or U22765 (N_22765,N_22034,N_20599);
or U22766 (N_22766,N_20682,N_20138);
and U22767 (N_22767,N_22486,N_21146);
or U22768 (N_22768,N_20644,N_21709);
xnor U22769 (N_22769,N_20206,N_21127);
nand U22770 (N_22770,N_21021,N_20845);
or U22771 (N_22771,N_20201,N_20857);
or U22772 (N_22772,N_20932,N_21534);
and U22773 (N_22773,N_20245,N_21471);
nor U22774 (N_22774,N_20677,N_20098);
xor U22775 (N_22775,N_21680,N_22109);
and U22776 (N_22776,N_20872,N_22248);
xor U22777 (N_22777,N_22380,N_20616);
and U22778 (N_22778,N_21905,N_22478);
and U22779 (N_22779,N_20712,N_20884);
and U22780 (N_22780,N_21623,N_21061);
nor U22781 (N_22781,N_21735,N_21405);
xnor U22782 (N_22782,N_21095,N_22428);
nor U22783 (N_22783,N_21892,N_20534);
or U22784 (N_22784,N_21372,N_21737);
xor U22785 (N_22785,N_21734,N_21318);
xor U22786 (N_22786,N_20359,N_20443);
and U22787 (N_22787,N_21902,N_21940);
nor U22788 (N_22788,N_20003,N_20190);
xor U22789 (N_22789,N_21258,N_21713);
nor U22790 (N_22790,N_20061,N_20707);
nand U22791 (N_22791,N_20213,N_20447);
nand U22792 (N_22792,N_20701,N_20026);
or U22793 (N_22793,N_21217,N_20128);
xor U22794 (N_22794,N_22022,N_21593);
or U22795 (N_22795,N_20164,N_21956);
nand U22796 (N_22796,N_21419,N_20726);
or U22797 (N_22797,N_21865,N_22408);
or U22798 (N_22798,N_20115,N_21052);
nor U22799 (N_22799,N_20556,N_22293);
nand U22800 (N_22800,N_21882,N_20148);
or U22801 (N_22801,N_20828,N_21805);
xnor U22802 (N_22802,N_22202,N_21357);
and U22803 (N_22803,N_20249,N_21317);
nor U22804 (N_22804,N_20412,N_22154);
or U22805 (N_22805,N_22350,N_22302);
nand U22806 (N_22806,N_22419,N_20469);
or U22807 (N_22807,N_21993,N_21015);
or U22808 (N_22808,N_20365,N_20247);
xnor U22809 (N_22809,N_22045,N_21990);
nand U22810 (N_22810,N_22105,N_20168);
and U22811 (N_22811,N_21180,N_21421);
nor U22812 (N_22812,N_22425,N_20269);
nor U22813 (N_22813,N_20824,N_20998);
and U22814 (N_22814,N_22384,N_22146);
or U22815 (N_22815,N_21188,N_21582);
xor U22816 (N_22816,N_21555,N_22273);
nor U22817 (N_22817,N_20528,N_22180);
nor U22818 (N_22818,N_21213,N_21894);
or U22819 (N_22819,N_21186,N_21436);
or U22820 (N_22820,N_20077,N_21374);
nand U22821 (N_22821,N_21725,N_21315);
nand U22822 (N_22822,N_20594,N_22059);
nor U22823 (N_22823,N_20294,N_20435);
nand U22824 (N_22824,N_20795,N_21660);
or U22825 (N_22825,N_20819,N_21209);
and U22826 (N_22826,N_20590,N_21720);
nand U22827 (N_22827,N_20173,N_22403);
xnor U22828 (N_22828,N_20971,N_21605);
nor U22829 (N_22829,N_21490,N_21779);
or U22830 (N_22830,N_21961,N_21539);
nor U22831 (N_22831,N_20894,N_21603);
and U22832 (N_22832,N_22125,N_21013);
xnor U22833 (N_22833,N_22444,N_21577);
xor U22834 (N_22834,N_20153,N_20806);
nor U22835 (N_22835,N_20521,N_20405);
and U22836 (N_22836,N_20561,N_20776);
nor U22837 (N_22837,N_20072,N_21398);
and U22838 (N_22838,N_21041,N_21417);
or U22839 (N_22839,N_20940,N_22294);
and U22840 (N_22840,N_20143,N_21009);
nand U22841 (N_22841,N_20271,N_21829);
xor U22842 (N_22842,N_21246,N_20110);
nand U22843 (N_22843,N_20895,N_20102);
and U22844 (N_22844,N_21560,N_20876);
nand U22845 (N_22845,N_20309,N_22476);
and U22846 (N_22846,N_20481,N_20893);
or U22847 (N_22847,N_20891,N_21916);
xor U22848 (N_22848,N_22358,N_21494);
or U22849 (N_22849,N_20887,N_21033);
and U22850 (N_22850,N_22469,N_21218);
xnor U22851 (N_22851,N_22381,N_20849);
or U22852 (N_22852,N_21104,N_21694);
xnor U22853 (N_22853,N_20046,N_20791);
xor U22854 (N_22854,N_20672,N_20986);
and U22855 (N_22855,N_20835,N_21777);
or U22856 (N_22856,N_21744,N_20531);
xnor U22857 (N_22857,N_21484,N_20262);
xnor U22858 (N_22858,N_20348,N_20720);
nor U22859 (N_22859,N_20293,N_21969);
nand U22860 (N_22860,N_21668,N_21330);
and U22861 (N_22861,N_21265,N_22195);
or U22862 (N_22862,N_22348,N_21478);
and U22863 (N_22863,N_21365,N_20413);
nor U22864 (N_22864,N_20242,N_20445);
nand U22865 (N_22865,N_21307,N_20010);
and U22866 (N_22866,N_21003,N_20827);
xnor U22867 (N_22867,N_20484,N_22495);
and U22868 (N_22868,N_20865,N_21693);
or U22869 (N_22869,N_20716,N_20602);
nand U22870 (N_22870,N_22113,N_22489);
nor U22871 (N_22871,N_21291,N_20193);
nor U22872 (N_22872,N_20515,N_21778);
or U22873 (N_22873,N_21240,N_20721);
or U22874 (N_22874,N_22032,N_21177);
xnor U22875 (N_22875,N_20376,N_22206);
nor U22876 (N_22876,N_22479,N_20285);
xnor U22877 (N_22877,N_20808,N_21840);
xor U22878 (N_22878,N_21020,N_20562);
xor U22879 (N_22879,N_21071,N_21966);
or U22880 (N_22880,N_22030,N_21914);
nor U22881 (N_22881,N_21236,N_22264);
nand U22882 (N_22882,N_20661,N_21126);
nor U22883 (N_22883,N_21764,N_20911);
or U22884 (N_22884,N_20494,N_22496);
or U22885 (N_22885,N_21877,N_22118);
nor U22886 (N_22886,N_21699,N_20393);
nand U22887 (N_22887,N_21808,N_22198);
and U22888 (N_22888,N_22477,N_21762);
and U22889 (N_22889,N_20035,N_21399);
nor U22890 (N_22890,N_20344,N_21214);
nand U22891 (N_22891,N_21107,N_21717);
or U22892 (N_22892,N_20299,N_20295);
and U22893 (N_22893,N_20220,N_20334);
xor U22894 (N_22894,N_21890,N_20291);
and U22895 (N_22895,N_20107,N_21796);
or U22896 (N_22896,N_21625,N_22416);
or U22897 (N_22897,N_21817,N_21986);
nand U22898 (N_22898,N_20120,N_21641);
or U22899 (N_22899,N_20491,N_20048);
or U22900 (N_22900,N_20160,N_20105);
nor U22901 (N_22901,N_22078,N_21671);
xor U22902 (N_22902,N_20088,N_21244);
nand U22903 (N_22903,N_21723,N_21163);
nand U22904 (N_22904,N_21093,N_21512);
or U22905 (N_22905,N_20837,N_20358);
xnor U22906 (N_22906,N_20338,N_20094);
or U22907 (N_22907,N_22010,N_21342);
or U22908 (N_22908,N_21587,N_20754);
xnor U22909 (N_22909,N_21981,N_21816);
xor U22910 (N_22910,N_20912,N_20111);
or U22911 (N_22911,N_20779,N_21930);
nand U22912 (N_22912,N_21351,N_20715);
nor U22913 (N_22913,N_21954,N_21081);
and U22914 (N_22914,N_20532,N_20377);
and U22915 (N_22915,N_21004,N_20527);
xnor U22916 (N_22916,N_22150,N_21970);
nor U22917 (N_22917,N_22050,N_20607);
xnor U22918 (N_22918,N_21656,N_20829);
xor U22919 (N_22919,N_20222,N_20318);
and U22920 (N_22920,N_21036,N_21257);
nand U22921 (N_22921,N_22075,N_20224);
or U22922 (N_22922,N_22356,N_20504);
nor U22923 (N_22923,N_22332,N_21726);
xnor U22924 (N_22924,N_21822,N_21354);
nor U22925 (N_22925,N_21583,N_21072);
or U22926 (N_22926,N_21287,N_20250);
or U22927 (N_22927,N_20335,N_22054);
xnor U22928 (N_22928,N_21519,N_22085);
nor U22929 (N_22929,N_21476,N_21856);
xor U22930 (N_22930,N_22111,N_21952);
and U22931 (N_22931,N_20962,N_20846);
or U22932 (N_22932,N_20970,N_20187);
nor U22933 (N_22933,N_20651,N_21332);
or U22934 (N_22934,N_20675,N_20812);
nor U22935 (N_22935,N_22196,N_21911);
nor U22936 (N_22936,N_21607,N_21496);
and U22937 (N_22937,N_21156,N_21065);
xnor U22938 (N_22938,N_20820,N_21366);
or U22939 (N_22939,N_21741,N_21048);
or U22940 (N_22940,N_22203,N_21812);
nand U22941 (N_22941,N_20961,N_20388);
or U22942 (N_22942,N_22292,N_22210);
and U22943 (N_22943,N_21367,N_21589);
nand U22944 (N_22944,N_22156,N_21043);
xor U22945 (N_22945,N_20156,N_20569);
xor U22946 (N_22946,N_22098,N_22345);
nand U22947 (N_22947,N_21957,N_21844);
nor U22948 (N_22948,N_20283,N_22016);
and U22949 (N_22949,N_20231,N_21843);
and U22950 (N_22950,N_21443,N_21141);
nor U22951 (N_22951,N_21750,N_21573);
nand U22952 (N_22952,N_22405,N_21090);
nor U22953 (N_22953,N_21225,N_21031);
or U22954 (N_22954,N_20004,N_21958);
or U22955 (N_22955,N_20953,N_22213);
xor U22956 (N_22956,N_21831,N_22254);
xor U22957 (N_22957,N_20790,N_20226);
nand U22958 (N_22958,N_20147,N_21568);
and U22959 (N_22959,N_21705,N_20900);
or U22960 (N_22960,N_21773,N_21827);
nand U22961 (N_22961,N_20658,N_22277);
nor U22962 (N_22962,N_22297,N_20693);
or U22963 (N_22963,N_21557,N_21995);
or U22964 (N_22964,N_22354,N_20343);
and U22965 (N_22965,N_20748,N_22089);
and U22966 (N_22966,N_20455,N_22436);
or U22967 (N_22967,N_22144,N_21462);
or U22968 (N_22968,N_22126,N_21259);
or U22969 (N_22969,N_20633,N_22083);
and U22970 (N_22970,N_20646,N_21820);
xor U22971 (N_22971,N_20794,N_20480);
nor U22972 (N_22972,N_22064,N_21147);
nand U22973 (N_22973,N_20807,N_21268);
xor U22974 (N_22974,N_20951,N_22231);
xor U22975 (N_22975,N_21771,N_22005);
nand U22976 (N_22976,N_20079,N_22137);
nand U22977 (N_22977,N_22448,N_21907);
and U22978 (N_22978,N_21313,N_22145);
nand U22979 (N_22979,N_20645,N_20456);
nand U22980 (N_22980,N_21378,N_20685);
xnor U22981 (N_22981,N_21035,N_20321);
nor U22982 (N_22982,N_20133,N_22328);
or U22983 (N_22983,N_21283,N_21182);
xnor U22984 (N_22984,N_20433,N_20304);
nand U22985 (N_22985,N_21998,N_22285);
and U22986 (N_22986,N_20896,N_22412);
nor U22987 (N_22987,N_21263,N_21999);
or U22988 (N_22988,N_22429,N_21994);
and U22989 (N_22989,N_21248,N_20727);
nand U22990 (N_22990,N_20965,N_21801);
nand U22991 (N_22991,N_21070,N_21222);
or U22992 (N_22992,N_21719,N_21155);
or U22993 (N_22993,N_21118,N_20000);
nor U22994 (N_22994,N_20274,N_20653);
and U22995 (N_22995,N_20383,N_21876);
and U22996 (N_22996,N_21951,N_21588);
nand U22997 (N_22997,N_21527,N_21947);
or U22998 (N_22998,N_21851,N_21140);
or U22999 (N_22999,N_20759,N_22107);
xnor U23000 (N_23000,N_21005,N_21708);
and U23001 (N_23001,N_20215,N_22462);
or U23002 (N_23002,N_20867,N_21349);
xnor U23003 (N_23003,N_21340,N_22014);
nor U23004 (N_23004,N_21886,N_20906);
nand U23005 (N_23005,N_20006,N_20760);
or U23006 (N_23006,N_22394,N_21804);
nor U23007 (N_23007,N_20964,N_21933);
xnor U23008 (N_23008,N_21608,N_21772);
nand U23009 (N_23009,N_21026,N_21124);
nand U23010 (N_23010,N_21692,N_22414);
and U23011 (N_23011,N_20514,N_20415);
and U23012 (N_23012,N_21207,N_21123);
xor U23013 (N_23013,N_20608,N_22205);
or U23014 (N_23014,N_20396,N_21464);
nand U23015 (N_23015,N_22153,N_21377);
nor U23016 (N_23016,N_21793,N_21078);
nor U23017 (N_23017,N_21731,N_21416);
nor U23018 (N_23018,N_20448,N_20251);
nor U23019 (N_23019,N_20074,N_22159);
and U23020 (N_23020,N_22402,N_20639);
or U23021 (N_23021,N_20990,N_21839);
nand U23022 (N_23022,N_20483,N_21630);
xor U23023 (N_23023,N_20605,N_22069);
nand U23024 (N_23024,N_21282,N_21872);
xnor U23025 (N_23025,N_21901,N_22188);
and U23026 (N_23026,N_20873,N_21706);
and U23027 (N_23027,N_22228,N_21461);
or U23028 (N_23028,N_21059,N_21506);
nand U23029 (N_23029,N_22281,N_21386);
xor U23030 (N_23030,N_21624,N_21867);
xnor U23031 (N_23031,N_21269,N_20793);
xor U23032 (N_23032,N_22391,N_22100);
nand U23033 (N_23033,N_22447,N_20792);
xor U23034 (N_23034,N_21423,N_20813);
nor U23035 (N_23035,N_20319,N_21513);
nand U23036 (N_23036,N_20910,N_20972);
nor U23037 (N_23037,N_22155,N_21113);
nor U23038 (N_23038,N_21508,N_21728);
nor U23039 (N_23039,N_21648,N_21364);
nand U23040 (N_23040,N_20270,N_21362);
or U23041 (N_23041,N_21524,N_21861);
nor U23042 (N_23042,N_20968,N_20040);
or U23043 (N_23043,N_20009,N_20637);
or U23044 (N_23044,N_20758,N_21164);
nand U23045 (N_23045,N_20134,N_22422);
and U23046 (N_23046,N_22006,N_20442);
and U23047 (N_23047,N_20286,N_21968);
nand U23048 (N_23048,N_22450,N_22470);
or U23049 (N_23049,N_21835,N_20816);
or U23050 (N_23050,N_21925,N_21601);
nand U23051 (N_23051,N_21194,N_20228);
and U23052 (N_23052,N_20750,N_21106);
nand U23053 (N_23053,N_20802,N_21432);
xnor U23054 (N_23054,N_21949,N_21286);
nor U23055 (N_23055,N_20522,N_22296);
and U23056 (N_23056,N_21922,N_21174);
nand U23057 (N_23057,N_20157,N_21776);
xor U23058 (N_23058,N_21455,N_22257);
and U23059 (N_23059,N_21233,N_22335);
nand U23060 (N_23060,N_20332,N_21338);
xor U23061 (N_23061,N_20493,N_20933);
and U23062 (N_23062,N_20129,N_22179);
nor U23063 (N_23063,N_22218,N_21252);
and U23064 (N_23064,N_22183,N_21795);
or U23065 (N_23065,N_22128,N_20324);
xor U23066 (N_23066,N_20449,N_21602);
nand U23067 (N_23067,N_20136,N_20298);
nor U23068 (N_23068,N_20174,N_20075);
nor U23069 (N_23069,N_20587,N_21618);
nor U23070 (N_23070,N_21037,N_21691);
or U23071 (N_23071,N_20765,N_20702);
xnor U23072 (N_23072,N_21069,N_21738);
and U23073 (N_23073,N_22219,N_20636);
or U23074 (N_23074,N_21220,N_20530);
or U23075 (N_23075,N_22346,N_22127);
xor U23076 (N_23076,N_20668,N_21888);
nor U23077 (N_23077,N_22147,N_21101);
nor U23078 (N_23078,N_21604,N_20630);
nor U23079 (N_23079,N_20752,N_20034);
nor U23080 (N_23080,N_20696,N_21532);
nor U23081 (N_23081,N_20116,N_20179);
xor U23082 (N_23082,N_20071,N_22186);
or U23083 (N_23083,N_20132,N_20634);
nor U23084 (N_23084,N_21451,N_20329);
and U23085 (N_23085,N_21885,N_20184);
or U23086 (N_23086,N_21381,N_20773);
or U23087 (N_23087,N_20015,N_22168);
nor U23088 (N_23088,N_20649,N_21492);
nor U23089 (N_23089,N_21938,N_20753);
nor U23090 (N_23090,N_20880,N_20749);
and U23091 (N_23091,N_20273,N_20825);
nor U23092 (N_23092,N_21567,N_20768);
nand U23093 (N_23093,N_22025,N_20821);
or U23094 (N_23094,N_21746,N_20473);
nor U23095 (N_23095,N_21967,N_20486);
or U23096 (N_23096,N_20113,N_21290);
or U23097 (N_23097,N_21339,N_20650);
and U23098 (N_23098,N_21837,N_22452);
nor U23099 (N_23099,N_21449,N_20281);
and U23100 (N_23100,N_20659,N_21383);
nor U23101 (N_23101,N_21757,N_21531);
nor U23102 (N_23102,N_21978,N_21145);
and U23103 (N_23103,N_22166,N_20875);
or U23104 (N_23104,N_21303,N_20742);
and U23105 (N_23105,N_22245,N_21828);
nand U23106 (N_23106,N_21296,N_22095);
and U23107 (N_23107,N_20236,N_20871);
or U23108 (N_23108,N_21424,N_20384);
nand U23109 (N_23109,N_22457,N_21200);
or U23110 (N_23110,N_20781,N_21518);
or U23111 (N_23111,N_21655,N_22404);
or U23112 (N_23112,N_21946,N_20524);
nor U23113 (N_23113,N_21830,N_22369);
nor U23114 (N_23114,N_20678,N_20777);
or U23115 (N_23115,N_20844,N_22256);
nand U23116 (N_23116,N_20302,N_20994);
xor U23117 (N_23117,N_22340,N_21853);
and U23118 (N_23118,N_21628,N_21669);
nor U23119 (N_23119,N_20454,N_21288);
and U23120 (N_23120,N_20541,N_22192);
or U23121 (N_23121,N_21117,N_22170);
and U23122 (N_23122,N_20679,N_21150);
xnor U23123 (N_23123,N_21950,N_22498);
xor U23124 (N_23124,N_21178,N_20422);
or U23125 (N_23125,N_20918,N_20788);
and U23126 (N_23126,N_20764,N_22220);
xor U23127 (N_23127,N_21992,N_22208);
or U23128 (N_23128,N_21142,N_22124);
nand U23129 (N_23129,N_20549,N_22000);
xor U23130 (N_23130,N_21488,N_21103);
xnor U23131 (N_23131,N_20622,N_21493);
and U23132 (N_23132,N_20657,N_21761);
or U23133 (N_23133,N_20021,N_20691);
and U23134 (N_23134,N_22398,N_20706);
or U23135 (N_23135,N_20687,N_21857);
nor U23136 (N_23136,N_21341,N_20225);
and U23137 (N_23137,N_21241,N_21564);
and U23138 (N_23138,N_20848,N_20560);
and U23139 (N_23139,N_21359,N_21308);
and U23140 (N_23140,N_20118,N_20586);
xor U23141 (N_23141,N_21547,N_21759);
nand U23142 (N_23142,N_22276,N_22483);
nor U23143 (N_23143,N_20624,N_21428);
nor U23144 (N_23144,N_21109,N_21204);
or U23145 (N_23145,N_20325,N_20680);
nand U23146 (N_23146,N_20297,N_21447);
nor U23147 (N_23147,N_20203,N_21918);
nor U23148 (N_23148,N_22033,N_21736);
nor U23149 (N_23149,N_21923,N_22041);
xnor U23150 (N_23150,N_22224,N_22007);
and U23151 (N_23151,N_20371,N_21475);
xor U23152 (N_23152,N_20866,N_21430);
and U23153 (N_23153,N_22349,N_20725);
and U23154 (N_23154,N_21025,N_20577);
nor U23155 (N_23155,N_21574,N_21237);
xor U23156 (N_23156,N_22121,N_20830);
nor U23157 (N_23157,N_22002,N_21809);
xor U23158 (N_23158,N_21409,N_21504);
xor U23159 (N_23159,N_22011,N_21008);
nand U23160 (N_23160,N_21787,N_20671);
xor U23161 (N_23161,N_21634,N_20978);
and U23162 (N_23162,N_22427,N_20221);
and U23163 (N_23163,N_22251,N_21682);
xnor U23164 (N_23164,N_20571,N_22484);
and U23165 (N_23165,N_21414,N_20517);
xor U23166 (N_23166,N_20508,N_21273);
and U23167 (N_23167,N_21863,N_22431);
nand U23168 (N_23168,N_20595,N_21854);
or U23169 (N_23169,N_21739,N_22164);
xnor U23170 (N_23170,N_20739,N_21208);
or U23171 (N_23171,N_20898,N_21929);
or U23172 (N_23172,N_22056,N_21874);
xnor U23173 (N_23173,N_20937,N_20070);
and U23174 (N_23174,N_20453,N_21860);
nor U23175 (N_23175,N_20234,N_21404);
and U23176 (N_23176,N_22140,N_22318);
nand U23177 (N_23177,N_22344,N_21858);
and U23178 (N_23178,N_20955,N_20565);
nand U23179 (N_23179,N_20087,N_20399);
nor U23180 (N_23180,N_22308,N_20341);
and U23181 (N_23181,N_22365,N_20002);
nor U23182 (N_23182,N_22062,N_21251);
xnor U23183 (N_23183,N_21267,N_22003);
or U23184 (N_23184,N_20336,N_22441);
nor U23185 (N_23185,N_20458,N_20323);
nor U23186 (N_23186,N_20440,N_21091);
and U23187 (N_23187,N_20351,N_20150);
and U23188 (N_23188,N_20860,N_20619);
and U23189 (N_23189,N_22181,N_22465);
or U23190 (N_23190,N_22143,N_22333);
and U23191 (N_23191,N_21195,N_20402);
xor U23192 (N_23192,N_21639,N_22130);
nor U23193 (N_23193,N_20090,N_21502);
and U23194 (N_23194,N_20049,N_22079);
or U23195 (N_23195,N_21964,N_21797);
nor U23196 (N_23196,N_20258,N_20814);
xor U23197 (N_23197,N_20444,N_20746);
nor U23198 (N_23198,N_20864,N_20089);
and U23199 (N_23199,N_20214,N_21974);
and U23200 (N_23200,N_21745,N_20022);
or U23201 (N_23201,N_22138,N_20738);
or U23202 (N_23202,N_20101,N_22230);
or U23203 (N_23203,N_21335,N_21606);
nand U23204 (N_23204,N_20320,N_20638);
and U23205 (N_23205,N_22172,N_21384);
and U23206 (N_23206,N_22102,N_21304);
nand U23207 (N_23207,N_21014,N_20417);
nand U23208 (N_23208,N_22312,N_20392);
nor U23209 (N_23209,N_20901,N_20019);
and U23210 (N_23210,N_21306,N_21074);
nand U23211 (N_23211,N_21658,N_22226);
or U23212 (N_23212,N_21943,N_21580);
or U23213 (N_23213,N_20420,N_21683);
nor U23214 (N_23214,N_21873,N_22037);
and U23215 (N_23215,N_20362,N_21260);
xor U23216 (N_23216,N_21247,N_21953);
xnor U23217 (N_23217,N_20047,N_21343);
xor U23218 (N_23218,N_21826,N_22148);
and U23219 (N_23219,N_20229,N_21242);
xnor U23220 (N_23220,N_22024,N_20670);
and U23221 (N_23221,N_22009,N_21480);
or U23222 (N_23222,N_20692,N_21941);
or U23223 (N_23223,N_20208,N_21264);
and U23224 (N_23224,N_20350,N_20067);
nor U23225 (N_23225,N_20663,N_21783);
xnor U23226 (N_23226,N_22266,N_21205);
xor U23227 (N_23227,N_20688,N_20252);
nand U23228 (N_23228,N_21285,N_22135);
xor U23229 (N_23229,N_20711,N_20123);
nor U23230 (N_23230,N_20890,N_20732);
nand U23231 (N_23231,N_21653,N_20254);
nor U23232 (N_23232,N_21165,N_22406);
and U23233 (N_23233,N_21371,N_20406);
xnor U23234 (N_23234,N_21733,N_22103);
nor U23235 (N_23235,N_21944,N_22383);
nor U23236 (N_23236,N_21181,N_21799);
or U23237 (N_23237,N_21473,N_20008);
xnor U23238 (N_23238,N_21710,N_20620);
xor U23239 (N_23239,N_21212,N_22473);
nand U23240 (N_23240,N_20728,N_22243);
xnor U23241 (N_23241,N_21316,N_21450);
nand U23242 (N_23242,N_21878,N_21053);
and U23243 (N_23243,N_21881,N_20992);
or U23244 (N_23244,N_20119,N_21067);
nand U23245 (N_23245,N_21250,N_22421);
nand U23246 (N_23246,N_20869,N_20064);
nand U23247 (N_23247,N_21469,N_22097);
nand U23248 (N_23248,N_20667,N_20969);
and U23249 (N_23249,N_21495,N_21846);
and U23250 (N_23250,N_21049,N_21299);
and U23251 (N_23251,N_20288,N_21276);
xor U23252 (N_23252,N_20809,N_20043);
xor U23253 (N_23253,N_20195,N_20568);
xnor U23254 (N_23254,N_20267,N_21266);
nand U23255 (N_23255,N_20916,N_20144);
and U23256 (N_23256,N_21979,N_20248);
or U23257 (N_23257,N_20407,N_21685);
xnor U23258 (N_23258,N_20374,N_21426);
nand U23259 (N_23259,N_22223,N_21598);
or U23260 (N_23260,N_20277,N_22430);
nand U23261 (N_23261,N_22413,N_22269);
or U23262 (N_23262,N_21689,N_21167);
xnor U23263 (N_23263,N_20626,N_20733);
xnor U23264 (N_23264,N_21128,N_20772);
or U23265 (N_23265,N_21298,N_21497);
nand U23266 (N_23266,N_20369,N_20576);
xnor U23267 (N_23267,N_22122,N_20438);
nor U23268 (N_23268,N_20853,N_22472);
nand U23269 (N_23269,N_21971,N_21732);
xnor U23270 (N_23270,N_21517,N_21448);
nand U23271 (N_23271,N_21535,N_20542);
and U23272 (N_23272,N_22040,N_21230);
or U23273 (N_23273,N_21360,N_22018);
nand U23274 (N_23274,N_22086,N_21825);
nor U23275 (N_23275,N_21996,N_21184);
or U23276 (N_23276,N_21452,N_21883);
or U23277 (N_23277,N_22253,N_22013);
xnor U23278 (N_23278,N_22178,N_22433);
xor U23279 (N_23279,N_21909,N_20958);
xor U23280 (N_23280,N_22446,N_21849);
or U23281 (N_23281,N_22376,N_21774);
xnor U23282 (N_23282,N_21521,N_21479);
and U23283 (N_23283,N_20870,N_20945);
or U23284 (N_23284,N_22163,N_21721);
xor U23285 (N_23285,N_21813,N_20897);
and U23286 (N_23286,N_20730,N_20632);
or U23287 (N_23287,N_20284,N_21891);
or U23288 (N_23288,N_20326,N_21898);
nand U23289 (N_23289,N_20611,N_20305);
nor U23290 (N_23290,N_20466,N_20537);
or U23291 (N_23291,N_20360,N_20993);
nor U23292 (N_23292,N_21379,N_20695);
nand U23293 (N_23293,N_21243,N_21201);
nor U23294 (N_23294,N_22268,N_20729);
xor U23295 (N_23295,N_20588,N_21445);
nor U23296 (N_23296,N_21231,N_20146);
nand U23297 (N_23297,N_20139,N_21852);
nand U23298 (N_23298,N_21818,N_20987);
or U23299 (N_23299,N_21505,N_21224);
nand U23300 (N_23300,N_22038,N_20909);
or U23301 (N_23301,N_20811,N_21295);
or U23302 (N_23302,N_20878,N_21042);
nor U23303 (N_23303,N_21099,N_22129);
nand U23304 (N_23304,N_20724,N_21649);
nor U23305 (N_23305,N_21747,N_20189);
nand U23306 (N_23306,N_22263,N_20903);
or U23307 (N_23307,N_20315,N_21546);
nand U23308 (N_23308,N_20239,N_22091);
nor U23309 (N_23309,N_22197,N_22359);
and U23310 (N_23310,N_20745,N_20656);
nand U23311 (N_23311,N_20307,N_20815);
nor U23312 (N_23312,N_20936,N_21919);
nand U23313 (N_23313,N_21046,N_22409);
or U23314 (N_23314,N_20919,N_20097);
nor U23315 (N_23315,N_21824,N_21596);
xor U23316 (N_23316,N_21509,N_22322);
or U23317 (N_23317,N_22280,N_21991);
and U23318 (N_23318,N_21302,N_20836);
nand U23319 (N_23319,N_20785,N_20574);
xnor U23320 (N_23320,N_20770,N_21132);
xor U23321 (N_23321,N_20183,N_21677);
and U23322 (N_23322,N_22157,N_22060);
or U23323 (N_23323,N_21866,N_21636);
and U23324 (N_23324,N_20127,N_20735);
or U23325 (N_23325,N_20856,N_22165);
xor U23326 (N_23326,N_20314,N_22372);
or U23327 (N_23327,N_21096,N_21791);
xor U23328 (N_23328,N_22116,N_21810);
nor U23329 (N_23329,N_20557,N_22289);
xor U23330 (N_23330,N_21089,N_21058);
and U23331 (N_23331,N_21915,N_20357);
and U23332 (N_23332,N_20555,N_21355);
nand U23333 (N_23333,N_20073,N_21080);
nand U23334 (N_23334,N_20581,N_20261);
xor U23335 (N_23335,N_20354,N_21051);
nor U23336 (N_23336,N_21211,N_21875);
or U23337 (N_23337,N_20425,N_20931);
or U23338 (N_23338,N_21092,N_20584);
nor U23339 (N_23339,N_22200,N_20001);
nor U23340 (N_23340,N_22407,N_22036);
or U23341 (N_23341,N_22485,N_21226);
nand U23342 (N_23342,N_21007,N_20999);
or U23343 (N_23343,N_22262,N_21006);
nand U23344 (N_23344,N_20037,N_21740);
nand U23345 (N_23345,N_21712,N_22169);
and U23346 (N_23346,N_21198,N_22068);
and U23347 (N_23347,N_22199,N_20355);
nor U23348 (N_23348,N_20030,N_20554);
nor U23349 (N_23349,N_20519,N_21579);
or U23350 (N_23350,N_21722,N_20959);
nand U23351 (N_23351,N_21197,N_20427);
and U23352 (N_23352,N_21190,N_20464);
nor U23353 (N_23353,N_20511,N_22028);
or U23354 (N_23354,N_20171,N_20741);
nor U23355 (N_23355,N_22027,N_20227);
xor U23356 (N_23356,N_21767,N_21934);
and U23357 (N_23357,N_20841,N_20592);
or U23358 (N_23358,N_20409,N_21196);
xnor U23359 (N_23359,N_20723,N_20690);
or U23360 (N_23360,N_20471,N_22370);
or U23361 (N_23361,N_22187,N_22301);
nor U23362 (N_23362,N_21000,N_22493);
xnor U23363 (N_23363,N_21438,N_21565);
nand U23364 (N_23364,N_21530,N_21895);
nand U23365 (N_23365,N_22184,N_22212);
nand U23366 (N_23366,N_20859,N_22261);
nand U23367 (N_23367,N_21613,N_20666);
nor U23368 (N_23368,N_22221,N_20609);
and U23369 (N_23369,N_21255,N_20989);
xnor U23370 (N_23370,N_21032,N_21503);
nor U23371 (N_23371,N_22411,N_21632);
or U23372 (N_23372,N_20439,N_21752);
xor U23373 (N_23373,N_20718,N_20292);
and U23374 (N_23374,N_20172,N_20676);
nand U23375 (N_23375,N_21672,N_21679);
and U23376 (N_23376,N_21369,N_21834);
or U23377 (N_23377,N_22497,N_20470);
nor U23378 (N_23378,N_21412,N_21556);
xnor U23379 (N_23379,N_20149,N_21572);
nand U23380 (N_23380,N_21594,N_22115);
nor U23381 (N_23381,N_21622,N_20382);
and U23382 (N_23382,N_22305,N_21645);
or U23383 (N_23383,N_20582,N_22057);
nand U23384 (N_23384,N_21921,N_22377);
nor U23385 (N_23385,N_21510,N_21760);
xor U23386 (N_23386,N_21870,N_21789);
xor U23387 (N_23387,N_20398,N_20734);
xor U23388 (N_23388,N_22339,N_21908);
and U23389 (N_23389,N_21499,N_20613);
nand U23390 (N_23390,N_20460,N_22341);
nor U23391 (N_23391,N_21686,N_22387);
xnor U23392 (N_23392,N_20180,N_22216);
xor U23393 (N_23393,N_21782,N_20016);
and U23394 (N_23394,N_21640,N_20058);
nor U23395 (N_23395,N_21724,N_20570);
xnor U23396 (N_23396,N_20282,N_21022);
and U23397 (N_23397,N_20540,N_20996);
nand U23398 (N_23398,N_22189,N_22282);
nand U23399 (N_23399,N_22046,N_21803);
nor U23400 (N_23400,N_21098,N_22475);
nor U23401 (N_23401,N_21755,N_20496);
nor U23402 (N_23402,N_21329,N_20093);
or U23403 (N_23403,N_20017,N_20991);
xnor U23404 (N_23404,N_20782,N_20769);
nand U23405 (N_23405,N_21050,N_20684);
xnor U23406 (N_23406,N_21924,N_20140);
and U23407 (N_23407,N_22090,N_21702);
nand U23408 (N_23408,N_21380,N_20737);
nand U23409 (N_23409,N_22278,N_20310);
and U23410 (N_23410,N_20957,N_22246);
nand U23411 (N_23411,N_20977,N_20780);
xor U23412 (N_23412,N_20925,N_21245);
or U23413 (N_23413,N_20142,N_20137);
nor U23414 (N_23414,N_21742,N_21576);
xor U23415 (N_23415,N_20974,N_20946);
and U23416 (N_23416,N_21684,N_20051);
xnor U23417 (N_23417,N_20550,N_21620);
or U23418 (N_23418,N_22351,N_21039);
and U23419 (N_23419,N_22284,N_21038);
nor U23420 (N_23420,N_20240,N_20489);
nand U23421 (N_23421,N_20122,N_21599);
and U23422 (N_23422,N_20025,N_21869);
or U23423 (N_23423,N_21016,N_21166);
nand U23424 (N_23424,N_21427,N_21228);
xor U23425 (N_23425,N_21559,N_21621);
nand U23426 (N_23426,N_22160,N_20223);
xor U23427 (N_23427,N_21390,N_20477);
nor U23428 (N_23428,N_22319,N_21615);
or U23429 (N_23429,N_20888,N_21363);
nand U23430 (N_23430,N_21749,N_22400);
xor U23431 (N_23431,N_22334,N_21959);
nor U23432 (N_23432,N_22337,N_21115);
nor U23433 (N_23433,N_20163,N_21753);
nand U23434 (N_23434,N_20069,N_20503);
nand U23435 (N_23435,N_21609,N_22491);
or U23436 (N_23436,N_22106,N_22267);
nor U23437 (N_23437,N_22242,N_20060);
xor U23438 (N_23438,N_22173,N_20799);
and U23439 (N_23439,N_20862,N_21256);
xnor U23440 (N_23440,N_20832,N_21935);
or U23441 (N_23441,N_20800,N_20810);
nor U23442 (N_23442,N_20395,N_21121);
nand U23443 (N_23443,N_20879,N_21463);
nand U23444 (N_23444,N_22175,N_20886);
or U23445 (N_23445,N_20192,N_22445);
xor U23446 (N_23446,N_20099,N_21017);
xnor U23447 (N_23447,N_21442,N_22397);
and U23448 (N_23448,N_21681,N_22317);
xor U23449 (N_23449,N_20461,N_21368);
and U23450 (N_23450,N_20755,N_21833);
xor U23451 (N_23451,N_22004,N_21292);
or U23452 (N_23452,N_22463,N_21552);
or U23453 (N_23453,N_20066,N_21807);
nor U23454 (N_23454,N_21470,N_22141);
nor U23455 (N_23455,N_20709,N_21149);
xnor U23456 (N_23456,N_21389,N_22439);
nand U23457 (N_23457,N_21540,N_21187);
xor U23458 (N_23458,N_22162,N_20255);
or U23459 (N_23459,N_20381,N_22008);
or U23460 (N_23460,N_21169,N_21249);
nor U23461 (N_23461,N_21408,N_21175);
and U23462 (N_23462,N_22058,N_20506);
and U23463 (N_23463,N_21823,N_20641);
xor U23464 (N_23464,N_22052,N_20647);
or U23465 (N_23465,N_20743,N_21597);
nor U23466 (N_23466,N_20145,N_20698);
or U23467 (N_23467,N_21122,N_21551);
nor U23468 (N_23468,N_21151,N_22134);
xnor U23469 (N_23469,N_22388,N_20786);
and U23470 (N_23470,N_21321,N_21661);
nand U23471 (N_23471,N_21172,N_20078);
nor U23472 (N_23472,N_20446,N_20621);
or U23473 (N_23473,N_21942,N_21391);
nor U23474 (N_23474,N_21982,N_21697);
nand U23475 (N_23475,N_22051,N_22291);
nand U23476 (N_23476,N_21715,N_20083);
nand U23477 (N_23477,N_22371,N_21375);
nor U23478 (N_23478,N_22193,N_21323);
or U23479 (N_23479,N_21765,N_21152);
nor U23480 (N_23480,N_20831,N_20260);
nand U23481 (N_23481,N_22443,N_20664);
or U23482 (N_23482,N_20085,N_21792);
or U23483 (N_23483,N_21987,N_22065);
xnor U23484 (N_23484,N_22149,N_21116);
or U23485 (N_23485,N_21094,N_20474);
or U23486 (N_23486,N_20042,N_20259);
xnor U23487 (N_23487,N_21454,N_20539);
or U23488 (N_23488,N_21769,N_21453);
and U23489 (N_23489,N_21650,N_21868);
nand U23490 (N_23490,N_20217,N_21333);
nand U23491 (N_23491,N_20404,N_21790);
or U23492 (N_23492,N_20479,N_21848);
nand U23493 (N_23493,N_21393,N_22182);
xnor U23494 (N_23494,N_21403,N_21880);
or U23495 (N_23495,N_21420,N_20204);
nand U23496 (N_23496,N_20525,N_20020);
nor U23497 (N_23497,N_22209,N_21491);
xor U23498 (N_23498,N_20512,N_20076);
nand U23499 (N_23499,N_21130,N_22283);
nand U23500 (N_23500,N_22211,N_21111);
nand U23501 (N_23501,N_21119,N_22290);
xnor U23502 (N_23502,N_20207,N_22327);
or U23503 (N_23503,N_20411,N_20662);
nand U23504 (N_23504,N_20926,N_20154);
xnor U23505 (N_23505,N_20459,N_20502);
nand U23506 (N_23506,N_22235,N_20475);
or U23507 (N_23507,N_21988,N_21931);
nand U23508 (N_23508,N_21665,N_21238);
xnor U23509 (N_23509,N_20200,N_21433);
or U23510 (N_23510,N_20373,N_20995);
nand U23511 (N_23511,N_21191,N_20432);
or U23512 (N_23512,N_22215,N_21278);
or U23513 (N_23513,N_21487,N_20194);
and U23514 (N_23514,N_21766,N_22355);
xnor U23515 (N_23515,N_21219,N_22367);
nor U23516 (N_23516,N_21085,N_22420);
and U23517 (N_23517,N_21270,N_20490);
and U23518 (N_23518,N_20546,N_21887);
nor U23519 (N_23519,N_21425,N_21544);
xnor U23520 (N_23520,N_22299,N_20400);
and U23521 (N_23521,N_21786,N_20775);
xnor U23522 (N_23522,N_22194,N_21458);
and U23523 (N_23523,N_21274,N_21410);
and U23524 (N_23524,N_21468,N_21920);
xor U23525 (N_23525,N_21229,N_20414);
or U23526 (N_23526,N_22250,N_21105);
nand U23527 (N_23527,N_20908,N_21973);
and U23528 (N_23528,N_22451,N_22252);
xnor U23529 (N_23529,N_21896,N_22295);
xnor U23530 (N_23530,N_21932,N_20266);
nand U23531 (N_23531,N_21199,N_20347);
xor U23532 (N_23532,N_22385,N_21821);
or U23533 (N_23533,N_22087,N_22152);
or U23534 (N_23534,N_20740,N_22119);
or U23535 (N_23535,N_22077,N_21611);
and U23536 (N_23536,N_20268,N_20673);
xor U23537 (N_23537,N_22092,N_20410);
xor U23538 (N_23538,N_20126,N_22120);
or U23539 (N_23539,N_21889,N_22074);
nor U23540 (N_23540,N_21082,N_21144);
nand U23541 (N_23541,N_21138,N_20589);
nor U23542 (N_23542,N_20722,N_21616);
nor U23543 (N_23543,N_21345,N_21936);
nor U23544 (N_23544,N_21097,N_20219);
nand U23545 (N_23545,N_21481,N_22455);
or U23546 (N_23546,N_22133,N_21575);
or U23547 (N_23547,N_20287,N_20390);
nand U23548 (N_23548,N_20057,N_21704);
and U23549 (N_23549,N_20854,N_20960);
nor U23550 (N_23550,N_20050,N_20237);
nor U23551 (N_23551,N_21281,N_22362);
or U23552 (N_23552,N_22363,N_22331);
or U23553 (N_23553,N_21600,N_21284);
nand U23554 (N_23554,N_20095,N_22093);
and U23555 (N_23555,N_20290,N_21906);
nor U23556 (N_23556,N_22114,N_21373);
and U23557 (N_23557,N_20181,N_20091);
or U23558 (N_23558,N_20364,N_21382);
nor U23559 (N_23559,N_20796,N_21763);
and U23560 (N_23560,N_22012,N_20188);
nor U23561 (N_23561,N_20552,N_20518);
nand U23562 (N_23562,N_20762,N_21018);
or U23563 (N_23563,N_20902,N_20843);
or U23564 (N_23564,N_21356,N_20548);
nand U23565 (N_23565,N_21775,N_20272);
nor U23566 (N_23566,N_22240,N_21903);
and U23567 (N_23567,N_22434,N_21862);
nand U23568 (N_23568,N_20457,N_20907);
nor U23569 (N_23569,N_20575,N_21202);
xnor U23570 (N_23570,N_20635,N_21137);
or U23571 (N_23571,N_20834,N_21185);
nand U23572 (N_23572,N_22270,N_21294);
nand U23573 (N_23573,N_21610,N_20920);
nand U23574 (N_23574,N_22399,N_21586);
or U23575 (N_23575,N_22336,N_21401);
xnor U23576 (N_23576,N_21695,N_21507);
or U23577 (N_23577,N_20855,N_20610);
and U23578 (N_23578,N_20196,N_21571);
and U23579 (N_23579,N_21234,N_21536);
and U23580 (N_23580,N_20492,N_20155);
xor U23581 (N_23581,N_21529,N_21459);
xor U23582 (N_23582,N_22274,N_21674);
xor U23583 (N_23583,N_21730,N_22368);
nand U23584 (N_23584,N_22300,N_21139);
xor U23585 (N_23585,N_21352,N_20487);
xnor U23586 (N_23586,N_22049,N_20585);
nand U23587 (N_23587,N_20059,N_20804);
or U23588 (N_23588,N_20744,N_20151);
and U23589 (N_23589,N_20963,N_21344);
xnor U23590 (N_23590,N_22361,N_22232);
or U23591 (N_23591,N_20301,N_21626);
and U23592 (N_23592,N_20603,N_21297);
xor U23593 (N_23593,N_21483,N_22279);
nor U23594 (N_23594,N_20767,N_21654);
nor U23595 (N_23595,N_20842,N_20615);
nand U23596 (N_23596,N_21516,N_21581);
xor U23597 (N_23597,N_22323,N_20979);
or U23598 (N_23598,N_20394,N_21675);
xor U23599 (N_23599,N_20922,N_20789);
and U23600 (N_23600,N_21289,N_20135);
nand U23601 (N_23601,N_20086,N_22360);
and U23602 (N_23602,N_22438,N_21422);
nor U23603 (N_23603,N_21153,N_21511);
nor U23604 (N_23604,N_20202,N_20617);
and U23605 (N_23605,N_22487,N_21239);
nand U23606 (N_23606,N_22110,N_21358);
nand U23607 (N_23607,N_21125,N_22042);
nor U23608 (N_23608,N_21562,N_21701);
and U23609 (N_23609,N_20322,N_21203);
or U23610 (N_23610,N_20108,N_20166);
nand U23611 (N_23611,N_20660,N_21102);
nand U23612 (N_23612,N_22298,N_21928);
nand U23613 (N_23613,N_21413,N_22442);
nand U23614 (N_23614,N_22084,N_21910);
xor U23615 (N_23615,N_21073,N_20822);
xor U23616 (N_23616,N_20572,N_22437);
nor U23617 (N_23617,N_21489,N_20152);
nand U23618 (N_23618,N_20141,N_22031);
nand U23619 (N_23619,N_20705,N_20980);
nor U23620 (N_23620,N_21280,N_22080);
and U23621 (N_23621,N_20499,N_21392);
and U23622 (N_23622,N_22275,N_21271);
or U23623 (N_23623,N_21223,N_20170);
or U23624 (N_23624,N_21277,N_20033);
or U23625 (N_23625,N_21158,N_22471);
nand U23626 (N_23626,N_20950,N_20424);
and U23627 (N_23627,N_20100,N_20162);
nor U23628 (N_23628,N_20104,N_21627);
xnor U23629 (N_23629,N_20452,N_20774);
nor U23630 (N_23630,N_21148,N_22158);
nand U23631 (N_23631,N_22171,N_20930);
and U23632 (N_23632,N_21800,N_21466);
xor U23633 (N_23633,N_22423,N_20495);
and U23634 (N_23634,N_22247,N_20327);
nor U23635 (N_23635,N_22123,N_20628);
or U23636 (N_23636,N_20451,N_20510);
or U23637 (N_23637,N_21815,N_20498);
and U23638 (N_23638,N_21751,N_22375);
nand U23639 (N_23639,N_21716,N_21976);
and U23640 (N_23640,N_20683,N_21794);
xnor U23641 (N_23641,N_22396,N_21585);
and U23642 (N_23642,N_22071,N_20674);
xor U23643 (N_23643,N_20988,N_21651);
xor U23644 (N_23644,N_21542,N_20241);
nor U23645 (N_23645,N_22227,N_20065);
and U23646 (N_23646,N_20787,N_20176);
xnor U23647 (N_23647,N_21034,N_22303);
or U23648 (N_23648,N_22048,N_22225);
and U23649 (N_23649,N_20185,N_20551);
xnor U23650 (N_23650,N_21376,N_20714);
xor U23651 (N_23651,N_21440,N_20096);
nor U23652 (N_23652,N_21129,N_20027);
nor U23653 (N_23653,N_21047,N_20233);
or U23654 (N_23654,N_21027,N_20578);
and U23655 (N_23655,N_21590,N_20985);
and U23656 (N_23656,N_21023,N_20013);
nor U23657 (N_23657,N_20028,N_20952);
and U23658 (N_23658,N_21652,N_20403);
nand U23659 (N_23659,N_21030,N_20689);
nor U23660 (N_23660,N_21100,N_22017);
and U23661 (N_23661,N_20275,N_21348);
nand U23662 (N_23662,N_22311,N_20600);
nand U23663 (N_23663,N_21293,N_20230);
and U23664 (N_23664,N_21435,N_22072);
or U23665 (N_23665,N_20523,N_20756);
nand U23666 (N_23666,N_20580,N_20431);
nand U23667 (N_23667,N_21319,N_20529);
and U23668 (N_23668,N_21019,N_21045);
nor U23669 (N_23669,N_22342,N_22066);
nand U23670 (N_23670,N_21718,N_20478);
and U23671 (N_23671,N_20218,N_22364);
and U23672 (N_23672,N_20238,N_21193);
or U23673 (N_23673,N_20045,N_20840);
nor U23674 (N_23674,N_21395,N_20103);
xnor U23675 (N_23675,N_20265,N_22490);
or U23676 (N_23676,N_22244,N_20436);
nand U23677 (N_23677,N_22073,N_20278);
xnor U23678 (N_23678,N_20805,N_22392);
nor U23679 (N_23679,N_21446,N_21310);
and U23680 (N_23680,N_20333,N_20092);
nand U23681 (N_23681,N_20300,N_21965);
xnor U23682 (N_23682,N_20708,N_20944);
and U23683 (N_23683,N_22415,N_22063);
nor U23684 (N_23684,N_20312,N_21850);
or U23685 (N_23685,N_21028,N_20669);
nand U23686 (N_23686,N_20117,N_21962);
xor U23687 (N_23687,N_21388,N_22458);
nor U23688 (N_23688,N_20803,N_20757);
or U23689 (N_23689,N_21972,N_20956);
or U23690 (N_23690,N_22461,N_21063);
nor U23691 (N_23691,N_21134,N_22055);
or U23692 (N_23692,N_20082,N_20913);
and U23693 (N_23693,N_20612,N_22081);
and U23694 (N_23694,N_20182,N_20054);
nand U23695 (N_23695,N_21465,N_20601);
nand U23696 (N_23696,N_20761,N_22026);
nor U23697 (N_23697,N_21619,N_21635);
xnor U23698 (N_23698,N_22112,N_21678);
and U23699 (N_23699,N_20751,N_22454);
nand U23700 (N_23700,N_22020,N_21802);
nand U23701 (N_23701,N_21690,N_21558);
and U23702 (N_23702,N_21631,N_22393);
xor U23703 (N_23703,N_20437,N_20526);
xnor U23704 (N_23704,N_20606,N_21939);
and U23705 (N_23705,N_20507,N_20308);
nor U23706 (N_23706,N_20372,N_22176);
or U23707 (N_23707,N_21077,N_20566);
and U23708 (N_23708,N_20408,N_20975);
and U23709 (N_23709,N_21176,N_21879);
xor U23710 (N_23710,N_21515,N_20482);
and U23711 (N_23711,N_21525,N_22481);
xor U23712 (N_23712,N_21168,N_21434);
xnor U23713 (N_23713,N_20080,N_20366);
nand U23714 (N_23714,N_21474,N_21756);
and U23715 (N_23715,N_20731,N_22325);
and U23716 (N_23716,N_20005,N_21221);
or U23717 (N_23717,N_22480,N_21612);
and U23718 (N_23718,N_20018,N_20161);
and U23719 (N_23719,N_20209,N_20784);
xnor U23720 (N_23720,N_22070,N_22464);
or U23721 (N_23721,N_21272,N_20216);
nand U23722 (N_23722,N_21083,N_22174);
nor U23723 (N_23723,N_21642,N_21183);
or U23724 (N_23724,N_22021,N_20340);
nand U23725 (N_23725,N_20256,N_20450);
and U23726 (N_23726,N_21262,N_21549);
or U23727 (N_23727,N_22386,N_21353);
or U23728 (N_23728,N_22265,N_21157);
nor U23729 (N_23729,N_20934,N_20544);
or U23730 (N_23730,N_22347,N_21667);
nand U23731 (N_23731,N_21537,N_20175);
nand U23732 (N_23732,N_21331,N_21638);
nor U23733 (N_23733,N_20704,N_20923);
nor U23734 (N_23734,N_20311,N_21301);
nand U23735 (N_23735,N_22249,N_20904);
or U23736 (N_23736,N_20559,N_20397);
or U23737 (N_23737,N_20243,N_22378);
xor U23738 (N_23738,N_20655,N_22190);
or U23739 (N_23739,N_21714,N_20939);
or U23740 (N_23740,N_21057,N_21216);
nand U23741 (N_23741,N_22207,N_21062);
xor U23742 (N_23742,N_20368,N_20346);
nor U23743 (N_23743,N_20747,N_22117);
or U23744 (N_23744,N_21002,N_22088);
xor U23745 (N_23745,N_20943,N_21305);
nand U23746 (N_23746,N_22029,N_21743);
and U23747 (N_23747,N_21173,N_21385);
nor U23748 (N_23748,N_20023,N_22047);
and U23749 (N_23749,N_21056,N_20881);
xnor U23750 (N_23750,N_20168,N_20972);
nor U23751 (N_23751,N_20983,N_21127);
xor U23752 (N_23752,N_21456,N_21743);
nor U23753 (N_23753,N_21256,N_22130);
and U23754 (N_23754,N_21352,N_20179);
or U23755 (N_23755,N_21872,N_21418);
or U23756 (N_23756,N_20102,N_21687);
nand U23757 (N_23757,N_20172,N_21696);
and U23758 (N_23758,N_22230,N_20804);
nand U23759 (N_23759,N_21539,N_20080);
and U23760 (N_23760,N_20817,N_22270);
nor U23761 (N_23761,N_22400,N_21467);
nor U23762 (N_23762,N_22449,N_21340);
or U23763 (N_23763,N_21001,N_21290);
nand U23764 (N_23764,N_20076,N_21930);
nand U23765 (N_23765,N_20758,N_21847);
or U23766 (N_23766,N_21077,N_21178);
nand U23767 (N_23767,N_20135,N_21594);
nand U23768 (N_23768,N_21289,N_20055);
nand U23769 (N_23769,N_20161,N_20805);
xor U23770 (N_23770,N_21964,N_21378);
and U23771 (N_23771,N_21592,N_21049);
and U23772 (N_23772,N_21198,N_21716);
nand U23773 (N_23773,N_21542,N_22485);
nor U23774 (N_23774,N_22029,N_20753);
nor U23775 (N_23775,N_20470,N_20163);
nor U23776 (N_23776,N_21461,N_20094);
xor U23777 (N_23777,N_21785,N_22246);
or U23778 (N_23778,N_21596,N_20854);
nand U23779 (N_23779,N_21505,N_20709);
xor U23780 (N_23780,N_21835,N_21209);
and U23781 (N_23781,N_20985,N_20633);
nand U23782 (N_23782,N_21523,N_20163);
or U23783 (N_23783,N_20643,N_21141);
nand U23784 (N_23784,N_20282,N_21618);
xnor U23785 (N_23785,N_22482,N_20610);
or U23786 (N_23786,N_20935,N_21126);
xor U23787 (N_23787,N_21027,N_21276);
nor U23788 (N_23788,N_22472,N_21653);
nand U23789 (N_23789,N_21354,N_20827);
nor U23790 (N_23790,N_20003,N_21484);
or U23791 (N_23791,N_21787,N_21666);
or U23792 (N_23792,N_20403,N_21635);
nor U23793 (N_23793,N_21408,N_20989);
nor U23794 (N_23794,N_21938,N_20452);
nand U23795 (N_23795,N_21456,N_20275);
xor U23796 (N_23796,N_20764,N_20307);
xnor U23797 (N_23797,N_21284,N_21707);
or U23798 (N_23798,N_20698,N_20827);
xor U23799 (N_23799,N_21883,N_21835);
nor U23800 (N_23800,N_22161,N_22249);
xor U23801 (N_23801,N_21173,N_21764);
and U23802 (N_23802,N_20875,N_20129);
nand U23803 (N_23803,N_20932,N_22310);
nor U23804 (N_23804,N_21680,N_20767);
nand U23805 (N_23805,N_21683,N_22156);
and U23806 (N_23806,N_21236,N_21096);
nand U23807 (N_23807,N_22092,N_20086);
nand U23808 (N_23808,N_21571,N_21558);
nor U23809 (N_23809,N_21720,N_21997);
nor U23810 (N_23810,N_20700,N_20397);
or U23811 (N_23811,N_20568,N_20627);
nor U23812 (N_23812,N_20641,N_22443);
xor U23813 (N_23813,N_20516,N_21900);
and U23814 (N_23814,N_21042,N_20452);
or U23815 (N_23815,N_20913,N_21587);
xor U23816 (N_23816,N_21202,N_20028);
nand U23817 (N_23817,N_22401,N_22480);
xnor U23818 (N_23818,N_20039,N_21050);
nand U23819 (N_23819,N_21783,N_22186);
nor U23820 (N_23820,N_21222,N_21166);
nand U23821 (N_23821,N_21560,N_21880);
nor U23822 (N_23822,N_22265,N_20633);
nor U23823 (N_23823,N_21761,N_21252);
nand U23824 (N_23824,N_20375,N_21238);
or U23825 (N_23825,N_20826,N_21372);
nand U23826 (N_23826,N_20541,N_21904);
xnor U23827 (N_23827,N_21501,N_20500);
nor U23828 (N_23828,N_20405,N_22324);
or U23829 (N_23829,N_20926,N_22299);
nor U23830 (N_23830,N_20374,N_20062);
xnor U23831 (N_23831,N_20290,N_21315);
and U23832 (N_23832,N_20853,N_21987);
and U23833 (N_23833,N_22479,N_21641);
or U23834 (N_23834,N_21760,N_22013);
nor U23835 (N_23835,N_20381,N_21432);
xor U23836 (N_23836,N_20559,N_22235);
xor U23837 (N_23837,N_21719,N_22348);
nand U23838 (N_23838,N_22120,N_21195);
xor U23839 (N_23839,N_22459,N_20213);
nor U23840 (N_23840,N_20791,N_20749);
nand U23841 (N_23841,N_20911,N_20954);
nor U23842 (N_23842,N_20378,N_20831);
nor U23843 (N_23843,N_21424,N_21442);
xnor U23844 (N_23844,N_21258,N_21554);
or U23845 (N_23845,N_20826,N_21462);
and U23846 (N_23846,N_21915,N_21628);
nor U23847 (N_23847,N_21372,N_21826);
nor U23848 (N_23848,N_20859,N_22071);
or U23849 (N_23849,N_22234,N_22011);
nand U23850 (N_23850,N_22109,N_22014);
nand U23851 (N_23851,N_21709,N_21281);
and U23852 (N_23852,N_21700,N_20719);
and U23853 (N_23853,N_21933,N_21673);
nand U23854 (N_23854,N_21500,N_22106);
and U23855 (N_23855,N_22030,N_22368);
xor U23856 (N_23856,N_21285,N_21543);
or U23857 (N_23857,N_20280,N_20923);
nand U23858 (N_23858,N_20742,N_21788);
nand U23859 (N_23859,N_21896,N_20330);
nor U23860 (N_23860,N_22496,N_22127);
or U23861 (N_23861,N_20462,N_22105);
nor U23862 (N_23862,N_20838,N_21930);
xnor U23863 (N_23863,N_21047,N_20000);
nand U23864 (N_23864,N_21333,N_20906);
and U23865 (N_23865,N_20900,N_21912);
nand U23866 (N_23866,N_20286,N_21460);
and U23867 (N_23867,N_20481,N_22091);
or U23868 (N_23868,N_20042,N_20844);
or U23869 (N_23869,N_20662,N_21328);
xor U23870 (N_23870,N_22392,N_21127);
or U23871 (N_23871,N_20643,N_20606);
xnor U23872 (N_23872,N_20581,N_22445);
or U23873 (N_23873,N_22281,N_22242);
or U23874 (N_23874,N_21183,N_20429);
and U23875 (N_23875,N_22179,N_21446);
or U23876 (N_23876,N_20799,N_20475);
nand U23877 (N_23877,N_21097,N_20002);
and U23878 (N_23878,N_21336,N_22324);
or U23879 (N_23879,N_22333,N_21378);
nand U23880 (N_23880,N_22199,N_20730);
xor U23881 (N_23881,N_20888,N_20220);
or U23882 (N_23882,N_20292,N_21742);
or U23883 (N_23883,N_20093,N_21248);
nand U23884 (N_23884,N_20732,N_21921);
nor U23885 (N_23885,N_21433,N_22270);
or U23886 (N_23886,N_21261,N_20322);
nor U23887 (N_23887,N_21606,N_20667);
and U23888 (N_23888,N_20395,N_22172);
nand U23889 (N_23889,N_20843,N_22495);
or U23890 (N_23890,N_22493,N_20465);
xnor U23891 (N_23891,N_21416,N_21334);
xor U23892 (N_23892,N_22050,N_20093);
nand U23893 (N_23893,N_20385,N_21015);
nor U23894 (N_23894,N_21921,N_22276);
nand U23895 (N_23895,N_20949,N_20768);
or U23896 (N_23896,N_21647,N_21733);
nand U23897 (N_23897,N_21369,N_20863);
xnor U23898 (N_23898,N_20404,N_22117);
xnor U23899 (N_23899,N_22127,N_21047);
or U23900 (N_23900,N_21741,N_22285);
and U23901 (N_23901,N_21199,N_21523);
nor U23902 (N_23902,N_22461,N_21069);
or U23903 (N_23903,N_21805,N_20854);
nand U23904 (N_23904,N_20348,N_20899);
or U23905 (N_23905,N_20414,N_20702);
nor U23906 (N_23906,N_20241,N_20039);
nand U23907 (N_23907,N_22017,N_21832);
and U23908 (N_23908,N_20139,N_21346);
nor U23909 (N_23909,N_21335,N_21256);
nor U23910 (N_23910,N_20953,N_22339);
xnor U23911 (N_23911,N_20827,N_20050);
nor U23912 (N_23912,N_21768,N_22490);
and U23913 (N_23913,N_20259,N_20841);
or U23914 (N_23914,N_21189,N_21180);
xnor U23915 (N_23915,N_20991,N_20934);
nor U23916 (N_23916,N_20596,N_21059);
nand U23917 (N_23917,N_20309,N_20099);
or U23918 (N_23918,N_21982,N_21904);
nand U23919 (N_23919,N_20572,N_22438);
nand U23920 (N_23920,N_22457,N_20171);
xor U23921 (N_23921,N_21675,N_21313);
nand U23922 (N_23922,N_21661,N_20549);
nand U23923 (N_23923,N_21195,N_20381);
nand U23924 (N_23924,N_21690,N_20037);
and U23925 (N_23925,N_21654,N_20279);
nor U23926 (N_23926,N_22318,N_21438);
xnor U23927 (N_23927,N_21857,N_21936);
nor U23928 (N_23928,N_21610,N_22039);
nor U23929 (N_23929,N_20953,N_22398);
or U23930 (N_23930,N_20473,N_21190);
nand U23931 (N_23931,N_22119,N_21816);
or U23932 (N_23932,N_21915,N_21652);
nor U23933 (N_23933,N_20479,N_20039);
xor U23934 (N_23934,N_20772,N_21299);
or U23935 (N_23935,N_21923,N_22438);
xnor U23936 (N_23936,N_21850,N_21006);
nor U23937 (N_23937,N_20153,N_21772);
nor U23938 (N_23938,N_21483,N_20989);
nor U23939 (N_23939,N_20862,N_21547);
or U23940 (N_23940,N_20409,N_21130);
nor U23941 (N_23941,N_20689,N_20467);
or U23942 (N_23942,N_22314,N_21001);
or U23943 (N_23943,N_20567,N_22329);
xor U23944 (N_23944,N_22171,N_20130);
and U23945 (N_23945,N_22029,N_21152);
nand U23946 (N_23946,N_20552,N_21231);
xor U23947 (N_23947,N_20421,N_20129);
nand U23948 (N_23948,N_22418,N_22128);
nand U23949 (N_23949,N_21328,N_20648);
and U23950 (N_23950,N_21149,N_22315);
or U23951 (N_23951,N_21297,N_20877);
xnor U23952 (N_23952,N_20673,N_21046);
nand U23953 (N_23953,N_21497,N_20060);
and U23954 (N_23954,N_22390,N_20873);
xnor U23955 (N_23955,N_20900,N_20120);
xor U23956 (N_23956,N_21093,N_20988);
nand U23957 (N_23957,N_21828,N_20876);
and U23958 (N_23958,N_22422,N_20639);
or U23959 (N_23959,N_21376,N_20405);
and U23960 (N_23960,N_20231,N_21334);
nand U23961 (N_23961,N_22020,N_22117);
xnor U23962 (N_23962,N_21048,N_22478);
xnor U23963 (N_23963,N_21802,N_20408);
nand U23964 (N_23964,N_20001,N_21116);
nor U23965 (N_23965,N_20886,N_21825);
xnor U23966 (N_23966,N_20198,N_20880);
or U23967 (N_23967,N_22391,N_20887);
nor U23968 (N_23968,N_20037,N_20276);
or U23969 (N_23969,N_22240,N_20061);
and U23970 (N_23970,N_21948,N_21159);
and U23971 (N_23971,N_20627,N_22437);
or U23972 (N_23972,N_21940,N_20977);
xnor U23973 (N_23973,N_21763,N_21604);
nand U23974 (N_23974,N_20700,N_20073);
and U23975 (N_23975,N_22030,N_20059);
nand U23976 (N_23976,N_21482,N_22445);
nand U23977 (N_23977,N_20366,N_22357);
xnor U23978 (N_23978,N_21373,N_21265);
xor U23979 (N_23979,N_20430,N_21400);
xor U23980 (N_23980,N_22282,N_21288);
nor U23981 (N_23981,N_21050,N_21437);
nand U23982 (N_23982,N_22153,N_22184);
xnor U23983 (N_23983,N_20297,N_20203);
xnor U23984 (N_23984,N_20486,N_20065);
xor U23985 (N_23985,N_22287,N_20192);
and U23986 (N_23986,N_20344,N_22115);
and U23987 (N_23987,N_22486,N_20846);
nor U23988 (N_23988,N_20834,N_22294);
or U23989 (N_23989,N_21654,N_20722);
nand U23990 (N_23990,N_22054,N_21228);
xor U23991 (N_23991,N_22400,N_21961);
nor U23992 (N_23992,N_22474,N_20771);
or U23993 (N_23993,N_20754,N_22158);
nand U23994 (N_23994,N_21051,N_20253);
xor U23995 (N_23995,N_21394,N_21617);
nor U23996 (N_23996,N_21308,N_21819);
or U23997 (N_23997,N_20462,N_20798);
nand U23998 (N_23998,N_20260,N_21055);
and U23999 (N_23999,N_20732,N_20917);
nand U24000 (N_24000,N_20597,N_20418);
or U24001 (N_24001,N_20697,N_22373);
and U24002 (N_24002,N_21862,N_20749);
xnor U24003 (N_24003,N_20709,N_21243);
or U24004 (N_24004,N_21029,N_20257);
nand U24005 (N_24005,N_21251,N_20052);
nand U24006 (N_24006,N_21744,N_20348);
nand U24007 (N_24007,N_21486,N_20410);
nand U24008 (N_24008,N_20826,N_22456);
nand U24009 (N_24009,N_21499,N_20911);
nand U24010 (N_24010,N_21456,N_22212);
or U24011 (N_24011,N_20907,N_20643);
nand U24012 (N_24012,N_21507,N_21128);
nand U24013 (N_24013,N_20466,N_22167);
and U24014 (N_24014,N_22375,N_20454);
xnor U24015 (N_24015,N_21462,N_20945);
nand U24016 (N_24016,N_21785,N_21903);
and U24017 (N_24017,N_21532,N_21237);
and U24018 (N_24018,N_21528,N_20665);
xor U24019 (N_24019,N_21589,N_22306);
nor U24020 (N_24020,N_21922,N_20155);
xor U24021 (N_24021,N_21904,N_20089);
xor U24022 (N_24022,N_20514,N_20506);
nor U24023 (N_24023,N_20426,N_20849);
xnor U24024 (N_24024,N_22447,N_21714);
nand U24025 (N_24025,N_22135,N_21789);
or U24026 (N_24026,N_21400,N_20078);
and U24027 (N_24027,N_22095,N_21876);
or U24028 (N_24028,N_21200,N_20463);
xnor U24029 (N_24029,N_20089,N_21721);
xnor U24030 (N_24030,N_21723,N_20712);
nand U24031 (N_24031,N_21594,N_21150);
nor U24032 (N_24032,N_21568,N_21497);
xnor U24033 (N_24033,N_21593,N_21057);
nor U24034 (N_24034,N_20769,N_21370);
and U24035 (N_24035,N_20588,N_21047);
xnor U24036 (N_24036,N_20978,N_22269);
xnor U24037 (N_24037,N_21843,N_22471);
or U24038 (N_24038,N_20392,N_21426);
or U24039 (N_24039,N_22060,N_22022);
nand U24040 (N_24040,N_22183,N_21431);
xor U24041 (N_24041,N_21518,N_21983);
nand U24042 (N_24042,N_21492,N_21337);
nand U24043 (N_24043,N_20505,N_20394);
xnor U24044 (N_24044,N_21320,N_21176);
nor U24045 (N_24045,N_20259,N_21144);
xnor U24046 (N_24046,N_20392,N_21894);
xor U24047 (N_24047,N_21447,N_22200);
xor U24048 (N_24048,N_21176,N_21890);
nand U24049 (N_24049,N_21089,N_20054);
nor U24050 (N_24050,N_20125,N_22026);
nand U24051 (N_24051,N_22460,N_22408);
and U24052 (N_24052,N_20887,N_22133);
and U24053 (N_24053,N_20007,N_21941);
or U24054 (N_24054,N_20437,N_20223);
xor U24055 (N_24055,N_21354,N_20763);
or U24056 (N_24056,N_21963,N_20648);
xor U24057 (N_24057,N_21383,N_20190);
nor U24058 (N_24058,N_20516,N_20545);
nor U24059 (N_24059,N_21087,N_20018);
nand U24060 (N_24060,N_20356,N_21199);
and U24061 (N_24061,N_21749,N_21165);
nand U24062 (N_24062,N_21527,N_21875);
nor U24063 (N_24063,N_21277,N_21683);
and U24064 (N_24064,N_22404,N_21886);
and U24065 (N_24065,N_22048,N_20661);
nand U24066 (N_24066,N_21310,N_21176);
nor U24067 (N_24067,N_21391,N_21580);
or U24068 (N_24068,N_20157,N_21069);
or U24069 (N_24069,N_21924,N_21943);
or U24070 (N_24070,N_22335,N_20953);
nand U24071 (N_24071,N_20645,N_20163);
and U24072 (N_24072,N_20493,N_20571);
nand U24073 (N_24073,N_22219,N_22376);
nor U24074 (N_24074,N_21495,N_20650);
nand U24075 (N_24075,N_21801,N_20851);
xor U24076 (N_24076,N_21009,N_22317);
nor U24077 (N_24077,N_20442,N_20608);
xnor U24078 (N_24078,N_20449,N_21416);
xor U24079 (N_24079,N_21651,N_20990);
xnor U24080 (N_24080,N_22012,N_20187);
or U24081 (N_24081,N_21218,N_21536);
nand U24082 (N_24082,N_20676,N_21718);
nor U24083 (N_24083,N_20023,N_21749);
and U24084 (N_24084,N_21966,N_20401);
and U24085 (N_24085,N_21799,N_21179);
nand U24086 (N_24086,N_21646,N_20217);
xnor U24087 (N_24087,N_20124,N_20243);
and U24088 (N_24088,N_22403,N_21752);
nand U24089 (N_24089,N_21176,N_20874);
and U24090 (N_24090,N_20223,N_21248);
or U24091 (N_24091,N_20644,N_21282);
xnor U24092 (N_24092,N_21751,N_20609);
and U24093 (N_24093,N_22212,N_20049);
xnor U24094 (N_24094,N_22486,N_21323);
nand U24095 (N_24095,N_20920,N_20645);
xor U24096 (N_24096,N_21208,N_20290);
nor U24097 (N_24097,N_20851,N_20366);
nand U24098 (N_24098,N_20679,N_20240);
and U24099 (N_24099,N_21967,N_21900);
nand U24100 (N_24100,N_22238,N_20205);
nand U24101 (N_24101,N_21573,N_21925);
and U24102 (N_24102,N_20541,N_21523);
or U24103 (N_24103,N_21143,N_20752);
nor U24104 (N_24104,N_22005,N_20090);
xnor U24105 (N_24105,N_22368,N_21653);
nor U24106 (N_24106,N_21660,N_21909);
or U24107 (N_24107,N_20029,N_21432);
and U24108 (N_24108,N_21030,N_20235);
xnor U24109 (N_24109,N_21507,N_21732);
nor U24110 (N_24110,N_21557,N_20550);
or U24111 (N_24111,N_21062,N_20420);
and U24112 (N_24112,N_20342,N_20743);
or U24113 (N_24113,N_20385,N_20974);
and U24114 (N_24114,N_21722,N_20368);
or U24115 (N_24115,N_20648,N_22115);
nand U24116 (N_24116,N_22452,N_20028);
nand U24117 (N_24117,N_20884,N_21103);
xor U24118 (N_24118,N_20997,N_21214);
or U24119 (N_24119,N_21303,N_20833);
nor U24120 (N_24120,N_20581,N_20011);
nand U24121 (N_24121,N_20183,N_22283);
nand U24122 (N_24122,N_20066,N_20377);
nand U24123 (N_24123,N_22256,N_21456);
and U24124 (N_24124,N_21070,N_20303);
and U24125 (N_24125,N_21737,N_20637);
and U24126 (N_24126,N_20263,N_20482);
nand U24127 (N_24127,N_21051,N_20545);
nor U24128 (N_24128,N_20976,N_20566);
xnor U24129 (N_24129,N_21170,N_21176);
and U24130 (N_24130,N_21051,N_22496);
xor U24131 (N_24131,N_20281,N_20059);
nor U24132 (N_24132,N_22440,N_21192);
nor U24133 (N_24133,N_22088,N_21556);
nand U24134 (N_24134,N_21826,N_20736);
nor U24135 (N_24135,N_20918,N_20069);
or U24136 (N_24136,N_20792,N_22384);
or U24137 (N_24137,N_22330,N_21157);
nand U24138 (N_24138,N_21054,N_21028);
nand U24139 (N_24139,N_20441,N_21909);
xor U24140 (N_24140,N_20702,N_20829);
nor U24141 (N_24141,N_21699,N_21785);
or U24142 (N_24142,N_22313,N_22255);
and U24143 (N_24143,N_20516,N_20895);
nor U24144 (N_24144,N_22497,N_21313);
nand U24145 (N_24145,N_20989,N_22235);
and U24146 (N_24146,N_20048,N_20419);
nor U24147 (N_24147,N_22112,N_21724);
and U24148 (N_24148,N_21571,N_20859);
nand U24149 (N_24149,N_21652,N_22031);
or U24150 (N_24150,N_20125,N_20365);
xnor U24151 (N_24151,N_21062,N_21772);
nor U24152 (N_24152,N_20278,N_22206);
xor U24153 (N_24153,N_21574,N_21011);
and U24154 (N_24154,N_21615,N_22371);
and U24155 (N_24155,N_21783,N_20558);
nand U24156 (N_24156,N_20641,N_22364);
xor U24157 (N_24157,N_20857,N_21506);
xor U24158 (N_24158,N_21368,N_21893);
xnor U24159 (N_24159,N_22234,N_22332);
or U24160 (N_24160,N_21415,N_22298);
or U24161 (N_24161,N_20000,N_20617);
xnor U24162 (N_24162,N_21791,N_21196);
nor U24163 (N_24163,N_21042,N_20290);
or U24164 (N_24164,N_21232,N_20044);
nor U24165 (N_24165,N_21495,N_22283);
xor U24166 (N_24166,N_21822,N_21557);
xnor U24167 (N_24167,N_21934,N_21741);
or U24168 (N_24168,N_21401,N_22311);
or U24169 (N_24169,N_21064,N_20514);
xnor U24170 (N_24170,N_20769,N_20971);
xnor U24171 (N_24171,N_21947,N_21903);
nand U24172 (N_24172,N_20882,N_22109);
or U24173 (N_24173,N_22035,N_20506);
or U24174 (N_24174,N_21048,N_21432);
and U24175 (N_24175,N_21018,N_20752);
nand U24176 (N_24176,N_21330,N_21996);
nor U24177 (N_24177,N_20373,N_20504);
xor U24178 (N_24178,N_22382,N_22483);
or U24179 (N_24179,N_20218,N_22223);
nand U24180 (N_24180,N_20668,N_21993);
or U24181 (N_24181,N_22071,N_22279);
nand U24182 (N_24182,N_21126,N_22486);
or U24183 (N_24183,N_20781,N_21912);
nor U24184 (N_24184,N_21689,N_21814);
xnor U24185 (N_24185,N_20572,N_20743);
nand U24186 (N_24186,N_22144,N_20883);
nand U24187 (N_24187,N_21502,N_20047);
and U24188 (N_24188,N_20006,N_20435);
nand U24189 (N_24189,N_21953,N_20126);
nand U24190 (N_24190,N_21801,N_21630);
and U24191 (N_24191,N_20813,N_20007);
and U24192 (N_24192,N_21373,N_22261);
or U24193 (N_24193,N_20295,N_21822);
xor U24194 (N_24194,N_21177,N_21564);
xnor U24195 (N_24195,N_20307,N_22015);
and U24196 (N_24196,N_20990,N_22051);
nor U24197 (N_24197,N_20080,N_20352);
and U24198 (N_24198,N_22034,N_21820);
xor U24199 (N_24199,N_21931,N_21947);
nand U24200 (N_24200,N_20684,N_20635);
xnor U24201 (N_24201,N_20626,N_20214);
nand U24202 (N_24202,N_22188,N_21295);
and U24203 (N_24203,N_20293,N_21467);
nand U24204 (N_24204,N_20957,N_21822);
or U24205 (N_24205,N_21923,N_22290);
xor U24206 (N_24206,N_20654,N_20667);
xnor U24207 (N_24207,N_21666,N_21804);
nand U24208 (N_24208,N_21755,N_21053);
or U24209 (N_24209,N_21247,N_21634);
nand U24210 (N_24210,N_21321,N_20354);
nand U24211 (N_24211,N_21974,N_21118);
xnor U24212 (N_24212,N_22442,N_21788);
or U24213 (N_24213,N_20853,N_20465);
or U24214 (N_24214,N_21100,N_21017);
or U24215 (N_24215,N_20722,N_21197);
and U24216 (N_24216,N_21939,N_22485);
xor U24217 (N_24217,N_21314,N_20889);
xnor U24218 (N_24218,N_22381,N_21289);
or U24219 (N_24219,N_21456,N_20187);
xnor U24220 (N_24220,N_22342,N_22293);
nor U24221 (N_24221,N_20444,N_21079);
and U24222 (N_24222,N_20862,N_20103);
xor U24223 (N_24223,N_21740,N_20384);
and U24224 (N_24224,N_20344,N_22202);
nand U24225 (N_24225,N_22150,N_21248);
nand U24226 (N_24226,N_20999,N_22481);
xor U24227 (N_24227,N_21164,N_21497);
nor U24228 (N_24228,N_22325,N_20396);
xor U24229 (N_24229,N_21683,N_20362);
nor U24230 (N_24230,N_20435,N_20317);
and U24231 (N_24231,N_20473,N_21505);
and U24232 (N_24232,N_20469,N_21797);
or U24233 (N_24233,N_21003,N_20833);
and U24234 (N_24234,N_20500,N_22428);
or U24235 (N_24235,N_22232,N_22077);
or U24236 (N_24236,N_21770,N_20490);
and U24237 (N_24237,N_20739,N_22143);
and U24238 (N_24238,N_22046,N_21694);
or U24239 (N_24239,N_21322,N_21791);
and U24240 (N_24240,N_20744,N_20722);
or U24241 (N_24241,N_20391,N_20115);
and U24242 (N_24242,N_20041,N_20986);
xor U24243 (N_24243,N_21801,N_20218);
and U24244 (N_24244,N_20065,N_20191);
or U24245 (N_24245,N_20287,N_20669);
nand U24246 (N_24246,N_21204,N_20520);
xor U24247 (N_24247,N_21027,N_20033);
or U24248 (N_24248,N_20539,N_20100);
nor U24249 (N_24249,N_21982,N_20196);
nand U24250 (N_24250,N_20615,N_20366);
and U24251 (N_24251,N_21053,N_20071);
or U24252 (N_24252,N_21510,N_20380);
or U24253 (N_24253,N_21515,N_22475);
nand U24254 (N_24254,N_20511,N_20161);
nand U24255 (N_24255,N_20908,N_21379);
nand U24256 (N_24256,N_21255,N_21962);
nor U24257 (N_24257,N_20530,N_20570);
nand U24258 (N_24258,N_20443,N_20821);
and U24259 (N_24259,N_20251,N_21978);
or U24260 (N_24260,N_20185,N_21544);
or U24261 (N_24261,N_22393,N_20711);
nand U24262 (N_24262,N_22014,N_20792);
nand U24263 (N_24263,N_21643,N_21386);
and U24264 (N_24264,N_20913,N_21258);
and U24265 (N_24265,N_20127,N_21048);
or U24266 (N_24266,N_20145,N_22482);
xor U24267 (N_24267,N_21076,N_22034);
and U24268 (N_24268,N_22228,N_20448);
xnor U24269 (N_24269,N_21284,N_21877);
or U24270 (N_24270,N_22358,N_21986);
or U24271 (N_24271,N_20855,N_20302);
xnor U24272 (N_24272,N_21895,N_22341);
xnor U24273 (N_24273,N_21477,N_21135);
nor U24274 (N_24274,N_20642,N_20640);
xnor U24275 (N_24275,N_21291,N_20237);
or U24276 (N_24276,N_21624,N_21779);
nor U24277 (N_24277,N_22221,N_20174);
or U24278 (N_24278,N_22494,N_20708);
and U24279 (N_24279,N_20910,N_21104);
nand U24280 (N_24280,N_21222,N_21483);
or U24281 (N_24281,N_21603,N_22166);
nand U24282 (N_24282,N_21165,N_20992);
nor U24283 (N_24283,N_20021,N_20967);
or U24284 (N_24284,N_21023,N_22290);
nand U24285 (N_24285,N_21083,N_20491);
or U24286 (N_24286,N_20113,N_20691);
nand U24287 (N_24287,N_21471,N_20847);
and U24288 (N_24288,N_22233,N_20585);
xor U24289 (N_24289,N_21468,N_20996);
or U24290 (N_24290,N_20646,N_20434);
xnor U24291 (N_24291,N_20971,N_21784);
and U24292 (N_24292,N_21361,N_21443);
or U24293 (N_24293,N_21945,N_22427);
xor U24294 (N_24294,N_20177,N_21946);
nand U24295 (N_24295,N_21435,N_20944);
nor U24296 (N_24296,N_22192,N_22077);
xor U24297 (N_24297,N_20314,N_22204);
nor U24298 (N_24298,N_22163,N_21478);
nand U24299 (N_24299,N_22263,N_20301);
xnor U24300 (N_24300,N_21137,N_21913);
nand U24301 (N_24301,N_21506,N_20624);
nor U24302 (N_24302,N_21738,N_21579);
nand U24303 (N_24303,N_21156,N_22461);
or U24304 (N_24304,N_20322,N_21836);
nand U24305 (N_24305,N_21271,N_20662);
nor U24306 (N_24306,N_21255,N_20662);
or U24307 (N_24307,N_20041,N_22389);
and U24308 (N_24308,N_21000,N_20825);
nand U24309 (N_24309,N_22392,N_20849);
nand U24310 (N_24310,N_21140,N_21959);
or U24311 (N_24311,N_20826,N_20126);
xor U24312 (N_24312,N_21720,N_22000);
nor U24313 (N_24313,N_21128,N_20169);
nand U24314 (N_24314,N_21182,N_21353);
xor U24315 (N_24315,N_22301,N_21013);
xnor U24316 (N_24316,N_22087,N_20342);
nand U24317 (N_24317,N_21608,N_21733);
nand U24318 (N_24318,N_22327,N_21730);
nand U24319 (N_24319,N_21179,N_20908);
and U24320 (N_24320,N_22293,N_21468);
and U24321 (N_24321,N_21178,N_20458);
nand U24322 (N_24322,N_20200,N_20056);
xor U24323 (N_24323,N_21994,N_20061);
xnor U24324 (N_24324,N_21938,N_21452);
nand U24325 (N_24325,N_21807,N_22278);
and U24326 (N_24326,N_20725,N_21527);
nor U24327 (N_24327,N_20394,N_20198);
and U24328 (N_24328,N_20160,N_22218);
nand U24329 (N_24329,N_22281,N_22245);
and U24330 (N_24330,N_22419,N_20299);
xor U24331 (N_24331,N_21039,N_22153);
nor U24332 (N_24332,N_20902,N_20707);
and U24333 (N_24333,N_22357,N_20526);
xor U24334 (N_24334,N_21773,N_21187);
nor U24335 (N_24335,N_21942,N_21474);
or U24336 (N_24336,N_22237,N_21941);
xor U24337 (N_24337,N_20102,N_20175);
xnor U24338 (N_24338,N_21007,N_21029);
or U24339 (N_24339,N_21610,N_21055);
xnor U24340 (N_24340,N_20047,N_20422);
and U24341 (N_24341,N_22200,N_20647);
or U24342 (N_24342,N_22265,N_20878);
nor U24343 (N_24343,N_20855,N_20356);
nand U24344 (N_24344,N_20806,N_21432);
nand U24345 (N_24345,N_21722,N_21303);
or U24346 (N_24346,N_22138,N_21481);
nand U24347 (N_24347,N_22028,N_20506);
nand U24348 (N_24348,N_22219,N_21540);
nor U24349 (N_24349,N_21250,N_21886);
nand U24350 (N_24350,N_20083,N_20535);
xor U24351 (N_24351,N_22418,N_21558);
and U24352 (N_24352,N_22364,N_22160);
and U24353 (N_24353,N_20597,N_20543);
and U24354 (N_24354,N_21301,N_22306);
or U24355 (N_24355,N_21913,N_21124);
and U24356 (N_24356,N_21951,N_22237);
nand U24357 (N_24357,N_20895,N_22276);
or U24358 (N_24358,N_20330,N_21093);
nor U24359 (N_24359,N_20476,N_21410);
xor U24360 (N_24360,N_22306,N_20693);
or U24361 (N_24361,N_20779,N_20654);
or U24362 (N_24362,N_20682,N_22473);
and U24363 (N_24363,N_22322,N_21791);
nand U24364 (N_24364,N_22219,N_21380);
nor U24365 (N_24365,N_22285,N_20715);
nor U24366 (N_24366,N_22040,N_21277);
xor U24367 (N_24367,N_21534,N_22241);
xor U24368 (N_24368,N_20239,N_21008);
nand U24369 (N_24369,N_22386,N_21164);
nor U24370 (N_24370,N_22423,N_20237);
or U24371 (N_24371,N_22125,N_21884);
or U24372 (N_24372,N_22462,N_20151);
nor U24373 (N_24373,N_21923,N_21776);
nor U24374 (N_24374,N_22156,N_21073);
xor U24375 (N_24375,N_20082,N_21962);
or U24376 (N_24376,N_20991,N_20310);
xnor U24377 (N_24377,N_22101,N_20158);
nand U24378 (N_24378,N_20712,N_20834);
xor U24379 (N_24379,N_21313,N_21497);
nand U24380 (N_24380,N_21881,N_21657);
and U24381 (N_24381,N_21170,N_20850);
nand U24382 (N_24382,N_21879,N_22339);
nand U24383 (N_24383,N_20970,N_20353);
xnor U24384 (N_24384,N_20537,N_20039);
and U24385 (N_24385,N_20072,N_22203);
nor U24386 (N_24386,N_20408,N_20222);
or U24387 (N_24387,N_20387,N_21471);
and U24388 (N_24388,N_20934,N_20572);
or U24389 (N_24389,N_21886,N_20763);
nor U24390 (N_24390,N_20327,N_21259);
and U24391 (N_24391,N_21791,N_21983);
or U24392 (N_24392,N_20619,N_22417);
xor U24393 (N_24393,N_20845,N_21680);
nand U24394 (N_24394,N_20290,N_20616);
or U24395 (N_24395,N_22418,N_21601);
and U24396 (N_24396,N_22120,N_20776);
or U24397 (N_24397,N_20210,N_21099);
xnor U24398 (N_24398,N_22050,N_21623);
nor U24399 (N_24399,N_22134,N_20523);
nor U24400 (N_24400,N_20369,N_20990);
or U24401 (N_24401,N_21771,N_21323);
nor U24402 (N_24402,N_22206,N_21690);
nand U24403 (N_24403,N_22411,N_22021);
xnor U24404 (N_24404,N_20829,N_22327);
nor U24405 (N_24405,N_22312,N_22300);
or U24406 (N_24406,N_20592,N_20394);
nand U24407 (N_24407,N_20702,N_20508);
nor U24408 (N_24408,N_21004,N_20818);
xnor U24409 (N_24409,N_22156,N_21719);
nor U24410 (N_24410,N_20918,N_20690);
or U24411 (N_24411,N_20938,N_20746);
nor U24412 (N_24412,N_20084,N_22209);
nor U24413 (N_24413,N_22236,N_20340);
xor U24414 (N_24414,N_21780,N_20571);
xor U24415 (N_24415,N_20893,N_20320);
xnor U24416 (N_24416,N_20547,N_21344);
nor U24417 (N_24417,N_20905,N_21824);
and U24418 (N_24418,N_22273,N_21262);
xor U24419 (N_24419,N_22344,N_21027);
xor U24420 (N_24420,N_21003,N_22137);
xor U24421 (N_24421,N_20051,N_22030);
or U24422 (N_24422,N_20807,N_20238);
nor U24423 (N_24423,N_20908,N_21966);
nand U24424 (N_24424,N_20791,N_21105);
xor U24425 (N_24425,N_22346,N_20562);
nor U24426 (N_24426,N_20324,N_21390);
and U24427 (N_24427,N_21473,N_20534);
nor U24428 (N_24428,N_21402,N_21315);
and U24429 (N_24429,N_20607,N_22072);
and U24430 (N_24430,N_20077,N_21318);
nor U24431 (N_24431,N_20251,N_20332);
or U24432 (N_24432,N_21387,N_20407);
nor U24433 (N_24433,N_20983,N_21648);
nand U24434 (N_24434,N_22388,N_22351);
and U24435 (N_24435,N_20344,N_20859);
and U24436 (N_24436,N_21558,N_20749);
nand U24437 (N_24437,N_21985,N_21847);
xor U24438 (N_24438,N_20436,N_21505);
or U24439 (N_24439,N_22475,N_20090);
xnor U24440 (N_24440,N_21569,N_20713);
or U24441 (N_24441,N_21266,N_21905);
nor U24442 (N_24442,N_21997,N_22322);
and U24443 (N_24443,N_20964,N_21372);
and U24444 (N_24444,N_20095,N_21698);
nor U24445 (N_24445,N_22133,N_21381);
xor U24446 (N_24446,N_21813,N_21957);
and U24447 (N_24447,N_20128,N_21471);
nand U24448 (N_24448,N_20477,N_21174);
nand U24449 (N_24449,N_20939,N_21033);
or U24450 (N_24450,N_20665,N_22268);
xor U24451 (N_24451,N_21108,N_22250);
or U24452 (N_24452,N_21508,N_22473);
and U24453 (N_24453,N_20730,N_21314);
nor U24454 (N_24454,N_21019,N_20800);
nand U24455 (N_24455,N_21656,N_21992);
and U24456 (N_24456,N_20156,N_20321);
nand U24457 (N_24457,N_20201,N_21817);
nor U24458 (N_24458,N_21371,N_20298);
or U24459 (N_24459,N_20825,N_20502);
or U24460 (N_24460,N_20996,N_20723);
xnor U24461 (N_24461,N_22385,N_22401);
nand U24462 (N_24462,N_20287,N_21338);
or U24463 (N_24463,N_20401,N_20440);
or U24464 (N_24464,N_22392,N_21648);
xor U24465 (N_24465,N_22028,N_21385);
xor U24466 (N_24466,N_21978,N_20717);
xnor U24467 (N_24467,N_21361,N_20852);
and U24468 (N_24468,N_22385,N_22272);
and U24469 (N_24469,N_20537,N_21670);
xnor U24470 (N_24470,N_20530,N_21765);
xnor U24471 (N_24471,N_20004,N_22374);
xnor U24472 (N_24472,N_21588,N_21248);
nor U24473 (N_24473,N_20156,N_21157);
and U24474 (N_24474,N_20911,N_22032);
nand U24475 (N_24475,N_21577,N_20137);
or U24476 (N_24476,N_20891,N_20186);
xor U24477 (N_24477,N_21766,N_22206);
nor U24478 (N_24478,N_20657,N_20922);
or U24479 (N_24479,N_21186,N_21860);
xor U24480 (N_24480,N_20999,N_21163);
or U24481 (N_24481,N_21232,N_21364);
and U24482 (N_24482,N_22301,N_21086);
or U24483 (N_24483,N_20782,N_21114);
xor U24484 (N_24484,N_22295,N_20339);
nor U24485 (N_24485,N_20137,N_20915);
xnor U24486 (N_24486,N_21122,N_21387);
nand U24487 (N_24487,N_22063,N_20175);
nor U24488 (N_24488,N_21213,N_22216);
nor U24489 (N_24489,N_20125,N_21544);
xnor U24490 (N_24490,N_20158,N_22271);
nand U24491 (N_24491,N_21184,N_21579);
nor U24492 (N_24492,N_20881,N_21822);
nor U24493 (N_24493,N_21259,N_22156);
or U24494 (N_24494,N_22483,N_20999);
nor U24495 (N_24495,N_21659,N_22478);
nor U24496 (N_24496,N_20274,N_20756);
xnor U24497 (N_24497,N_22185,N_21437);
nor U24498 (N_24498,N_21545,N_21962);
and U24499 (N_24499,N_20631,N_21265);
nand U24500 (N_24500,N_21181,N_20810);
xnor U24501 (N_24501,N_20655,N_21301);
xnor U24502 (N_24502,N_20052,N_22306);
nor U24503 (N_24503,N_21416,N_22032);
xor U24504 (N_24504,N_20454,N_20169);
and U24505 (N_24505,N_22224,N_20637);
nand U24506 (N_24506,N_20386,N_21434);
nand U24507 (N_24507,N_22154,N_22378);
and U24508 (N_24508,N_20863,N_21615);
xor U24509 (N_24509,N_22315,N_20190);
xor U24510 (N_24510,N_20739,N_20938);
and U24511 (N_24511,N_21365,N_21268);
and U24512 (N_24512,N_21444,N_20747);
nor U24513 (N_24513,N_21208,N_21242);
nand U24514 (N_24514,N_21312,N_22168);
nor U24515 (N_24515,N_20849,N_20972);
nor U24516 (N_24516,N_21452,N_21236);
or U24517 (N_24517,N_21564,N_20809);
nand U24518 (N_24518,N_21937,N_21311);
and U24519 (N_24519,N_20612,N_20582);
nand U24520 (N_24520,N_22456,N_22129);
and U24521 (N_24521,N_22024,N_20986);
xnor U24522 (N_24522,N_20641,N_20475);
nand U24523 (N_24523,N_20675,N_22176);
or U24524 (N_24524,N_20857,N_21193);
or U24525 (N_24525,N_20922,N_22273);
nor U24526 (N_24526,N_21655,N_20579);
nand U24527 (N_24527,N_22112,N_22458);
nand U24528 (N_24528,N_21364,N_22244);
xnor U24529 (N_24529,N_20533,N_20940);
nand U24530 (N_24530,N_22271,N_22163);
xor U24531 (N_24531,N_20910,N_22470);
nand U24532 (N_24532,N_21592,N_21561);
or U24533 (N_24533,N_21268,N_20884);
nor U24534 (N_24534,N_21782,N_21921);
or U24535 (N_24535,N_21084,N_21337);
and U24536 (N_24536,N_21988,N_20670);
xor U24537 (N_24537,N_20697,N_21056);
and U24538 (N_24538,N_21851,N_22211);
nor U24539 (N_24539,N_21084,N_20011);
and U24540 (N_24540,N_20069,N_21803);
nand U24541 (N_24541,N_21966,N_20032);
or U24542 (N_24542,N_21808,N_20333);
or U24543 (N_24543,N_21345,N_20924);
nor U24544 (N_24544,N_20311,N_20913);
or U24545 (N_24545,N_20482,N_22469);
nor U24546 (N_24546,N_21075,N_21301);
nand U24547 (N_24547,N_21413,N_22266);
and U24548 (N_24548,N_20023,N_20589);
xnor U24549 (N_24549,N_22060,N_21855);
or U24550 (N_24550,N_21373,N_21949);
nor U24551 (N_24551,N_21266,N_21691);
nand U24552 (N_24552,N_20047,N_21569);
and U24553 (N_24553,N_20553,N_20118);
nor U24554 (N_24554,N_20972,N_22116);
nor U24555 (N_24555,N_20390,N_21543);
xor U24556 (N_24556,N_21806,N_20581);
xor U24557 (N_24557,N_21752,N_21568);
and U24558 (N_24558,N_20881,N_22012);
nor U24559 (N_24559,N_21962,N_21425);
or U24560 (N_24560,N_20959,N_20644);
nor U24561 (N_24561,N_20014,N_22365);
and U24562 (N_24562,N_20107,N_21861);
or U24563 (N_24563,N_22462,N_20783);
or U24564 (N_24564,N_21954,N_21331);
nand U24565 (N_24565,N_20914,N_20113);
nand U24566 (N_24566,N_20510,N_21428);
and U24567 (N_24567,N_22181,N_21478);
nand U24568 (N_24568,N_21347,N_21324);
nor U24569 (N_24569,N_21033,N_21401);
nand U24570 (N_24570,N_20674,N_21827);
or U24571 (N_24571,N_20435,N_21072);
or U24572 (N_24572,N_21180,N_22004);
and U24573 (N_24573,N_20979,N_20192);
xnor U24574 (N_24574,N_20793,N_20011);
xor U24575 (N_24575,N_20756,N_20765);
nand U24576 (N_24576,N_21969,N_22189);
nand U24577 (N_24577,N_22214,N_20671);
and U24578 (N_24578,N_20670,N_22314);
xnor U24579 (N_24579,N_22462,N_22051);
or U24580 (N_24580,N_20322,N_20297);
or U24581 (N_24581,N_21268,N_22213);
or U24582 (N_24582,N_21781,N_21467);
nand U24583 (N_24583,N_20086,N_22026);
xor U24584 (N_24584,N_21949,N_21832);
and U24585 (N_24585,N_20063,N_22080);
or U24586 (N_24586,N_20745,N_20407);
xnor U24587 (N_24587,N_20262,N_21138);
xnor U24588 (N_24588,N_20053,N_20822);
or U24589 (N_24589,N_21990,N_22364);
nor U24590 (N_24590,N_21951,N_20905);
nand U24591 (N_24591,N_21690,N_20225);
xnor U24592 (N_24592,N_20987,N_22432);
nand U24593 (N_24593,N_22338,N_20981);
nand U24594 (N_24594,N_21681,N_22220);
nor U24595 (N_24595,N_22064,N_20416);
or U24596 (N_24596,N_20933,N_20405);
xnor U24597 (N_24597,N_22173,N_21596);
nor U24598 (N_24598,N_21211,N_22051);
or U24599 (N_24599,N_21892,N_22172);
nor U24600 (N_24600,N_22210,N_22004);
xor U24601 (N_24601,N_20548,N_21164);
nand U24602 (N_24602,N_21257,N_21449);
nand U24603 (N_24603,N_21998,N_20508);
or U24604 (N_24604,N_20122,N_20085);
and U24605 (N_24605,N_20773,N_22302);
xnor U24606 (N_24606,N_22439,N_20331);
and U24607 (N_24607,N_20701,N_21307);
and U24608 (N_24608,N_21134,N_20962);
nor U24609 (N_24609,N_20758,N_20131);
and U24610 (N_24610,N_21442,N_20011);
nor U24611 (N_24611,N_21162,N_22228);
nand U24612 (N_24612,N_21328,N_21776);
xor U24613 (N_24613,N_22320,N_20549);
and U24614 (N_24614,N_21441,N_20006);
or U24615 (N_24615,N_20806,N_21534);
nor U24616 (N_24616,N_22486,N_21357);
and U24617 (N_24617,N_21336,N_20969);
nor U24618 (N_24618,N_21096,N_21460);
nor U24619 (N_24619,N_20547,N_22002);
and U24620 (N_24620,N_21255,N_22455);
nor U24621 (N_24621,N_22334,N_21754);
or U24622 (N_24622,N_20841,N_20975);
xnor U24623 (N_24623,N_22093,N_21766);
xor U24624 (N_24624,N_21847,N_21120);
and U24625 (N_24625,N_20739,N_20301);
xnor U24626 (N_24626,N_21897,N_20816);
or U24627 (N_24627,N_20277,N_22139);
nand U24628 (N_24628,N_20618,N_20809);
xnor U24629 (N_24629,N_20165,N_20299);
nand U24630 (N_24630,N_20005,N_21479);
and U24631 (N_24631,N_21108,N_21078);
nor U24632 (N_24632,N_20299,N_21706);
nor U24633 (N_24633,N_21549,N_22187);
nand U24634 (N_24634,N_21195,N_20455);
nor U24635 (N_24635,N_21684,N_20158);
nor U24636 (N_24636,N_22438,N_21169);
nand U24637 (N_24637,N_20185,N_20248);
nor U24638 (N_24638,N_21603,N_21895);
and U24639 (N_24639,N_20424,N_21013);
nor U24640 (N_24640,N_21314,N_20871);
and U24641 (N_24641,N_21585,N_22045);
nand U24642 (N_24642,N_20859,N_20201);
xor U24643 (N_24643,N_20320,N_20279);
nor U24644 (N_24644,N_20635,N_21308);
or U24645 (N_24645,N_22475,N_21947);
and U24646 (N_24646,N_21550,N_20053);
nand U24647 (N_24647,N_21344,N_21089);
and U24648 (N_24648,N_20018,N_21268);
and U24649 (N_24649,N_21449,N_21249);
or U24650 (N_24650,N_20214,N_20902);
nand U24651 (N_24651,N_21700,N_22362);
nand U24652 (N_24652,N_21513,N_22189);
or U24653 (N_24653,N_21311,N_20528);
xor U24654 (N_24654,N_22432,N_21523);
or U24655 (N_24655,N_21087,N_22111);
xor U24656 (N_24656,N_21699,N_20628);
and U24657 (N_24657,N_21614,N_20616);
and U24658 (N_24658,N_21097,N_21285);
and U24659 (N_24659,N_22335,N_20837);
or U24660 (N_24660,N_21647,N_20001);
nor U24661 (N_24661,N_20053,N_22099);
nor U24662 (N_24662,N_20613,N_21816);
nand U24663 (N_24663,N_20415,N_20238);
or U24664 (N_24664,N_21343,N_22202);
or U24665 (N_24665,N_20270,N_20117);
nor U24666 (N_24666,N_22241,N_21834);
xor U24667 (N_24667,N_21824,N_21647);
nor U24668 (N_24668,N_22483,N_20809);
nand U24669 (N_24669,N_20906,N_20593);
nand U24670 (N_24670,N_22300,N_21257);
nor U24671 (N_24671,N_21513,N_20287);
nor U24672 (N_24672,N_20871,N_21087);
and U24673 (N_24673,N_20111,N_21397);
nor U24674 (N_24674,N_21174,N_20734);
nand U24675 (N_24675,N_21179,N_20994);
nand U24676 (N_24676,N_21359,N_22325);
nand U24677 (N_24677,N_21921,N_20130);
or U24678 (N_24678,N_20163,N_22370);
xor U24679 (N_24679,N_21850,N_21054);
nor U24680 (N_24680,N_20186,N_20685);
nor U24681 (N_24681,N_21921,N_20380);
nand U24682 (N_24682,N_22391,N_22129);
nand U24683 (N_24683,N_20640,N_21477);
nand U24684 (N_24684,N_20317,N_20324);
xnor U24685 (N_24685,N_22421,N_21994);
or U24686 (N_24686,N_21341,N_21545);
nand U24687 (N_24687,N_22319,N_21030);
nor U24688 (N_24688,N_21818,N_22140);
nor U24689 (N_24689,N_21992,N_20467);
nand U24690 (N_24690,N_21817,N_21576);
xor U24691 (N_24691,N_20328,N_22381);
and U24692 (N_24692,N_20107,N_20410);
xor U24693 (N_24693,N_22247,N_21778);
and U24694 (N_24694,N_20315,N_21329);
and U24695 (N_24695,N_20556,N_20636);
or U24696 (N_24696,N_21790,N_20242);
and U24697 (N_24697,N_21175,N_20524);
xnor U24698 (N_24698,N_21793,N_22476);
and U24699 (N_24699,N_22157,N_22138);
and U24700 (N_24700,N_21170,N_21539);
xor U24701 (N_24701,N_20476,N_22162);
xor U24702 (N_24702,N_21245,N_20147);
or U24703 (N_24703,N_20235,N_22148);
nand U24704 (N_24704,N_21268,N_20307);
and U24705 (N_24705,N_21202,N_20474);
or U24706 (N_24706,N_20153,N_21902);
nand U24707 (N_24707,N_22469,N_20410);
xnor U24708 (N_24708,N_21903,N_20716);
or U24709 (N_24709,N_20987,N_20511);
nand U24710 (N_24710,N_20155,N_20293);
or U24711 (N_24711,N_21082,N_22031);
or U24712 (N_24712,N_20712,N_21083);
nand U24713 (N_24713,N_22469,N_21794);
xnor U24714 (N_24714,N_20608,N_20954);
nand U24715 (N_24715,N_20927,N_21780);
nor U24716 (N_24716,N_20700,N_20378);
and U24717 (N_24717,N_22241,N_20001);
nand U24718 (N_24718,N_22416,N_21823);
and U24719 (N_24719,N_21962,N_21523);
or U24720 (N_24720,N_20834,N_22067);
nor U24721 (N_24721,N_21458,N_20463);
nor U24722 (N_24722,N_20934,N_20075);
nor U24723 (N_24723,N_20020,N_21721);
nor U24724 (N_24724,N_21203,N_22367);
xnor U24725 (N_24725,N_21919,N_21896);
nor U24726 (N_24726,N_20141,N_21560);
or U24727 (N_24727,N_20021,N_22213);
nand U24728 (N_24728,N_20755,N_22198);
nor U24729 (N_24729,N_20221,N_21907);
and U24730 (N_24730,N_21514,N_21433);
xor U24731 (N_24731,N_21786,N_20092);
xor U24732 (N_24732,N_20498,N_21872);
and U24733 (N_24733,N_21150,N_20114);
nand U24734 (N_24734,N_21866,N_20972);
or U24735 (N_24735,N_20854,N_20380);
nand U24736 (N_24736,N_21276,N_20353);
and U24737 (N_24737,N_20961,N_22392);
nand U24738 (N_24738,N_20865,N_22431);
or U24739 (N_24739,N_21279,N_21186);
nand U24740 (N_24740,N_20059,N_21348);
or U24741 (N_24741,N_20771,N_20478);
nor U24742 (N_24742,N_21989,N_21045);
nor U24743 (N_24743,N_21628,N_20202);
nor U24744 (N_24744,N_21435,N_21523);
nand U24745 (N_24745,N_21604,N_22459);
nor U24746 (N_24746,N_21207,N_21893);
or U24747 (N_24747,N_22497,N_20018);
and U24748 (N_24748,N_21425,N_20673);
or U24749 (N_24749,N_21402,N_20236);
and U24750 (N_24750,N_21310,N_20514);
xnor U24751 (N_24751,N_21146,N_20642);
and U24752 (N_24752,N_20086,N_21922);
xnor U24753 (N_24753,N_20594,N_21255);
nand U24754 (N_24754,N_21838,N_22279);
nand U24755 (N_24755,N_20974,N_20656);
xnor U24756 (N_24756,N_22279,N_20798);
nand U24757 (N_24757,N_21560,N_20084);
xor U24758 (N_24758,N_20864,N_20984);
nand U24759 (N_24759,N_21718,N_21074);
and U24760 (N_24760,N_22313,N_21459);
nand U24761 (N_24761,N_20899,N_21071);
or U24762 (N_24762,N_21263,N_20566);
and U24763 (N_24763,N_21610,N_21363);
nand U24764 (N_24764,N_21877,N_21854);
or U24765 (N_24765,N_22046,N_20219);
and U24766 (N_24766,N_22077,N_21320);
or U24767 (N_24767,N_20846,N_21935);
xnor U24768 (N_24768,N_20354,N_21974);
and U24769 (N_24769,N_20811,N_21453);
and U24770 (N_24770,N_20339,N_21569);
or U24771 (N_24771,N_20836,N_20413);
or U24772 (N_24772,N_20429,N_21014);
nor U24773 (N_24773,N_20082,N_22343);
nand U24774 (N_24774,N_20258,N_22393);
nand U24775 (N_24775,N_22474,N_20582);
and U24776 (N_24776,N_22476,N_20258);
and U24777 (N_24777,N_21533,N_22322);
and U24778 (N_24778,N_22300,N_22233);
or U24779 (N_24779,N_22112,N_20531);
xor U24780 (N_24780,N_22148,N_22421);
nand U24781 (N_24781,N_21679,N_22481);
or U24782 (N_24782,N_20732,N_20010);
nand U24783 (N_24783,N_21097,N_20042);
nand U24784 (N_24784,N_22000,N_22492);
xnor U24785 (N_24785,N_21348,N_22001);
or U24786 (N_24786,N_20668,N_20059);
xnor U24787 (N_24787,N_21170,N_20595);
and U24788 (N_24788,N_22268,N_20866);
and U24789 (N_24789,N_20409,N_21955);
and U24790 (N_24790,N_21044,N_22095);
xor U24791 (N_24791,N_21410,N_20229);
nand U24792 (N_24792,N_21740,N_20957);
xnor U24793 (N_24793,N_21154,N_20109);
nor U24794 (N_24794,N_22136,N_20085);
nor U24795 (N_24795,N_20601,N_20797);
and U24796 (N_24796,N_22424,N_20946);
and U24797 (N_24797,N_22431,N_20605);
or U24798 (N_24798,N_21730,N_21512);
xnor U24799 (N_24799,N_20486,N_22178);
and U24800 (N_24800,N_22068,N_20667);
nor U24801 (N_24801,N_20063,N_20431);
or U24802 (N_24802,N_20866,N_20447);
xor U24803 (N_24803,N_22027,N_20876);
xnor U24804 (N_24804,N_20105,N_20801);
or U24805 (N_24805,N_20411,N_20277);
nor U24806 (N_24806,N_21336,N_21238);
xnor U24807 (N_24807,N_20571,N_22494);
nor U24808 (N_24808,N_21448,N_20126);
nor U24809 (N_24809,N_21027,N_21311);
nand U24810 (N_24810,N_20413,N_21713);
or U24811 (N_24811,N_22055,N_20766);
nor U24812 (N_24812,N_21766,N_20538);
nor U24813 (N_24813,N_22239,N_20164);
nand U24814 (N_24814,N_21611,N_21170);
or U24815 (N_24815,N_20417,N_21417);
xor U24816 (N_24816,N_22129,N_21807);
nand U24817 (N_24817,N_21479,N_20285);
nor U24818 (N_24818,N_20799,N_22413);
xor U24819 (N_24819,N_22063,N_22460);
xor U24820 (N_24820,N_22186,N_21478);
or U24821 (N_24821,N_20043,N_21270);
xnor U24822 (N_24822,N_21043,N_20161);
nand U24823 (N_24823,N_22168,N_20498);
nor U24824 (N_24824,N_21286,N_20765);
and U24825 (N_24825,N_21870,N_22315);
nand U24826 (N_24826,N_21865,N_20236);
nand U24827 (N_24827,N_21234,N_22282);
xor U24828 (N_24828,N_22358,N_20316);
xor U24829 (N_24829,N_21667,N_21524);
nor U24830 (N_24830,N_21870,N_20791);
and U24831 (N_24831,N_20669,N_20530);
nand U24832 (N_24832,N_20005,N_20833);
nand U24833 (N_24833,N_20362,N_22098);
or U24834 (N_24834,N_20434,N_22407);
xnor U24835 (N_24835,N_22221,N_21858);
nor U24836 (N_24836,N_21882,N_21919);
xor U24837 (N_24837,N_21163,N_20615);
nand U24838 (N_24838,N_21658,N_21042);
and U24839 (N_24839,N_21969,N_21527);
nor U24840 (N_24840,N_22158,N_21047);
xnor U24841 (N_24841,N_20152,N_21808);
nand U24842 (N_24842,N_21705,N_21638);
nor U24843 (N_24843,N_21497,N_21013);
or U24844 (N_24844,N_22055,N_20145);
and U24845 (N_24845,N_21493,N_21896);
nand U24846 (N_24846,N_21273,N_21511);
nor U24847 (N_24847,N_21039,N_21296);
nor U24848 (N_24848,N_20426,N_20265);
nand U24849 (N_24849,N_22133,N_20253);
and U24850 (N_24850,N_21195,N_21262);
and U24851 (N_24851,N_22048,N_21140);
xnor U24852 (N_24852,N_20893,N_22338);
nor U24853 (N_24853,N_22420,N_21276);
and U24854 (N_24854,N_21921,N_20929);
and U24855 (N_24855,N_21067,N_20022);
nor U24856 (N_24856,N_21631,N_22436);
and U24857 (N_24857,N_20923,N_21125);
xnor U24858 (N_24858,N_20875,N_22167);
nor U24859 (N_24859,N_21541,N_22341);
or U24860 (N_24860,N_20349,N_20537);
xnor U24861 (N_24861,N_21260,N_21398);
xor U24862 (N_24862,N_21485,N_21075);
or U24863 (N_24863,N_20549,N_21927);
xor U24864 (N_24864,N_21070,N_20426);
nor U24865 (N_24865,N_21314,N_21024);
and U24866 (N_24866,N_20524,N_21133);
xnor U24867 (N_24867,N_20354,N_20451);
or U24868 (N_24868,N_20125,N_20694);
nand U24869 (N_24869,N_20163,N_22317);
and U24870 (N_24870,N_21846,N_22146);
xor U24871 (N_24871,N_21970,N_20384);
nor U24872 (N_24872,N_22233,N_21651);
and U24873 (N_24873,N_20659,N_20824);
or U24874 (N_24874,N_21532,N_20487);
xor U24875 (N_24875,N_21489,N_22203);
nor U24876 (N_24876,N_20399,N_20306);
or U24877 (N_24877,N_22399,N_20730);
or U24878 (N_24878,N_20683,N_22244);
nor U24879 (N_24879,N_20791,N_21165);
xnor U24880 (N_24880,N_20765,N_22260);
nand U24881 (N_24881,N_20420,N_21811);
nor U24882 (N_24882,N_20033,N_21689);
xor U24883 (N_24883,N_21338,N_20463);
and U24884 (N_24884,N_20196,N_21478);
or U24885 (N_24885,N_20309,N_21969);
and U24886 (N_24886,N_22054,N_21736);
nor U24887 (N_24887,N_20505,N_20466);
nand U24888 (N_24888,N_21226,N_20370);
and U24889 (N_24889,N_22097,N_21051);
and U24890 (N_24890,N_20850,N_20470);
nand U24891 (N_24891,N_21935,N_22475);
nand U24892 (N_24892,N_21569,N_21031);
and U24893 (N_24893,N_20579,N_20761);
xnor U24894 (N_24894,N_21702,N_21204);
nand U24895 (N_24895,N_21510,N_21755);
xnor U24896 (N_24896,N_21635,N_20209);
and U24897 (N_24897,N_22228,N_21347);
nor U24898 (N_24898,N_21528,N_20429);
xor U24899 (N_24899,N_21402,N_20617);
xnor U24900 (N_24900,N_21593,N_20842);
or U24901 (N_24901,N_20431,N_22017);
xnor U24902 (N_24902,N_20184,N_21552);
or U24903 (N_24903,N_20815,N_20101);
nor U24904 (N_24904,N_20500,N_20962);
or U24905 (N_24905,N_20599,N_21247);
xnor U24906 (N_24906,N_21636,N_21274);
nand U24907 (N_24907,N_22277,N_20066);
xnor U24908 (N_24908,N_21503,N_22049);
xor U24909 (N_24909,N_22234,N_20102);
xnor U24910 (N_24910,N_20421,N_20150);
nor U24911 (N_24911,N_21657,N_20358);
xnor U24912 (N_24912,N_21519,N_22404);
or U24913 (N_24913,N_21452,N_21323);
nor U24914 (N_24914,N_20326,N_20229);
xnor U24915 (N_24915,N_20524,N_21750);
xor U24916 (N_24916,N_20609,N_21402);
nor U24917 (N_24917,N_21425,N_22479);
xnor U24918 (N_24918,N_20621,N_20892);
and U24919 (N_24919,N_20266,N_20942);
and U24920 (N_24920,N_20296,N_21394);
nor U24921 (N_24921,N_20697,N_20885);
nand U24922 (N_24922,N_21096,N_20250);
or U24923 (N_24923,N_20091,N_22006);
and U24924 (N_24924,N_21186,N_20863);
or U24925 (N_24925,N_21541,N_20244);
nor U24926 (N_24926,N_20147,N_21359);
xnor U24927 (N_24927,N_21677,N_22127);
nor U24928 (N_24928,N_21946,N_22072);
or U24929 (N_24929,N_21206,N_20393);
or U24930 (N_24930,N_20223,N_22404);
and U24931 (N_24931,N_21855,N_21872);
xnor U24932 (N_24932,N_20886,N_21292);
nand U24933 (N_24933,N_21879,N_20494);
or U24934 (N_24934,N_20488,N_22350);
and U24935 (N_24935,N_20522,N_21058);
and U24936 (N_24936,N_21706,N_21701);
xnor U24937 (N_24937,N_21618,N_22176);
nand U24938 (N_24938,N_21521,N_20847);
nor U24939 (N_24939,N_20015,N_21259);
or U24940 (N_24940,N_20001,N_22092);
nand U24941 (N_24941,N_21568,N_21857);
and U24942 (N_24942,N_22391,N_20243);
nand U24943 (N_24943,N_20689,N_22353);
xor U24944 (N_24944,N_22430,N_22159);
nor U24945 (N_24945,N_21034,N_20333);
and U24946 (N_24946,N_22230,N_20923);
or U24947 (N_24947,N_22050,N_20690);
and U24948 (N_24948,N_20539,N_21627);
or U24949 (N_24949,N_20903,N_21769);
xnor U24950 (N_24950,N_21813,N_20040);
nor U24951 (N_24951,N_21284,N_22389);
and U24952 (N_24952,N_22105,N_20232);
nand U24953 (N_24953,N_22109,N_21475);
nand U24954 (N_24954,N_21565,N_20697);
xor U24955 (N_24955,N_21153,N_20944);
xnor U24956 (N_24956,N_21335,N_22024);
xnor U24957 (N_24957,N_21626,N_22242);
nand U24958 (N_24958,N_20096,N_21754);
and U24959 (N_24959,N_21721,N_20762);
nand U24960 (N_24960,N_20147,N_21556);
nand U24961 (N_24961,N_21004,N_22452);
or U24962 (N_24962,N_20375,N_20708);
or U24963 (N_24963,N_21010,N_22324);
xor U24964 (N_24964,N_21185,N_21759);
nand U24965 (N_24965,N_22177,N_20735);
and U24966 (N_24966,N_20220,N_20321);
or U24967 (N_24967,N_20146,N_20468);
nand U24968 (N_24968,N_21098,N_20237);
nor U24969 (N_24969,N_22097,N_22421);
or U24970 (N_24970,N_21294,N_22175);
and U24971 (N_24971,N_22048,N_20276);
or U24972 (N_24972,N_21818,N_20754);
xnor U24973 (N_24973,N_21915,N_21461);
nor U24974 (N_24974,N_20746,N_20951);
xnor U24975 (N_24975,N_21904,N_21896);
and U24976 (N_24976,N_20079,N_21355);
or U24977 (N_24977,N_21879,N_20442);
or U24978 (N_24978,N_21717,N_22069);
xnor U24979 (N_24979,N_21190,N_21286);
nand U24980 (N_24980,N_21486,N_21569);
or U24981 (N_24981,N_22077,N_21266);
nand U24982 (N_24982,N_21834,N_20028);
nor U24983 (N_24983,N_20366,N_21375);
nand U24984 (N_24984,N_22411,N_20227);
xnor U24985 (N_24985,N_20630,N_22209);
nor U24986 (N_24986,N_21857,N_22102);
xnor U24987 (N_24987,N_20044,N_20287);
and U24988 (N_24988,N_20045,N_22273);
xnor U24989 (N_24989,N_21210,N_21104);
nor U24990 (N_24990,N_21782,N_22341);
nand U24991 (N_24991,N_20922,N_20647);
nor U24992 (N_24992,N_20106,N_21924);
xor U24993 (N_24993,N_22283,N_21120);
nor U24994 (N_24994,N_21636,N_21140);
xor U24995 (N_24995,N_21476,N_20781);
or U24996 (N_24996,N_22497,N_21998);
or U24997 (N_24997,N_20801,N_20568);
nor U24998 (N_24998,N_22120,N_20666);
nor U24999 (N_24999,N_22380,N_22379);
nand U25000 (N_25000,N_24451,N_23480);
xor U25001 (N_25001,N_23290,N_22636);
nand U25002 (N_25002,N_24879,N_24005);
and U25003 (N_25003,N_24209,N_24499);
nand U25004 (N_25004,N_24321,N_22568);
or U25005 (N_25005,N_23139,N_23012);
nor U25006 (N_25006,N_22877,N_23934);
and U25007 (N_25007,N_24516,N_23774);
nor U25008 (N_25008,N_23600,N_23104);
xnor U25009 (N_25009,N_23944,N_23911);
or U25010 (N_25010,N_23834,N_23639);
nor U25011 (N_25011,N_23202,N_22508);
or U25012 (N_25012,N_24160,N_24827);
and U25013 (N_25013,N_23625,N_22555);
nor U25014 (N_25014,N_23133,N_23341);
xor U25015 (N_25015,N_24779,N_24784);
xor U25016 (N_25016,N_24269,N_22738);
nand U25017 (N_25017,N_23673,N_23888);
or U25018 (N_25018,N_24541,N_23142);
nor U25019 (N_25019,N_23090,N_23984);
nand U25020 (N_25020,N_23242,N_24057);
nor U25021 (N_25021,N_24168,N_23602);
xor U25022 (N_25022,N_24098,N_22548);
or U25023 (N_25023,N_24865,N_23508);
or U25024 (N_25024,N_23114,N_22980);
nor U25025 (N_25025,N_23676,N_24909);
or U25026 (N_25026,N_23475,N_23688);
nand U25027 (N_25027,N_24186,N_24976);
nand U25028 (N_25028,N_24034,N_24935);
nor U25029 (N_25029,N_24037,N_22930);
nor U25030 (N_25030,N_22707,N_22810);
xor U25031 (N_25031,N_24312,N_23775);
xnor U25032 (N_25032,N_24617,N_23649);
nor U25033 (N_25033,N_24855,N_22733);
xor U25034 (N_25034,N_24553,N_23029);
or U25035 (N_25035,N_24573,N_24838);
or U25036 (N_25036,N_23216,N_23608);
xor U25037 (N_25037,N_22895,N_23221);
nor U25038 (N_25038,N_22634,N_24635);
nor U25039 (N_25039,N_23179,N_23623);
and U25040 (N_25040,N_23906,N_23154);
nand U25041 (N_25041,N_24698,N_22604);
or U25042 (N_25042,N_23809,N_23177);
or U25043 (N_25043,N_22708,N_24226);
nand U25044 (N_25044,N_23359,N_23690);
nor U25045 (N_25045,N_23886,N_23778);
or U25046 (N_25046,N_22748,N_22745);
or U25047 (N_25047,N_23421,N_24352);
nand U25048 (N_25048,N_23605,N_23237);
xor U25049 (N_25049,N_23245,N_23067);
nor U25050 (N_25050,N_23721,N_22857);
or U25051 (N_25051,N_23529,N_24257);
xor U25052 (N_25052,N_23921,N_23742);
and U25053 (N_25053,N_22759,N_22608);
and U25054 (N_25054,N_22900,N_23940);
nand U25055 (N_25055,N_24601,N_24810);
nor U25056 (N_25056,N_24000,N_23042);
xor U25057 (N_25057,N_23483,N_24609);
nor U25058 (N_25058,N_24164,N_24863);
nand U25059 (N_25059,N_22963,N_23233);
and U25060 (N_25060,N_24822,N_22528);
xor U25061 (N_25061,N_22815,N_24272);
nor U25062 (N_25062,N_24254,N_24276);
xor U25063 (N_25063,N_24705,N_22909);
xnor U25064 (N_25064,N_24154,N_23334);
nand U25065 (N_25065,N_23008,N_23293);
xnor U25066 (N_25066,N_24859,N_24889);
nand U25067 (N_25067,N_24809,N_23800);
xor U25068 (N_25068,N_23776,N_22560);
xnor U25069 (N_25069,N_23770,N_24943);
nand U25070 (N_25070,N_24593,N_24237);
nand U25071 (N_25071,N_23590,N_24500);
xnor U25072 (N_25072,N_24509,N_23871);
nor U25073 (N_25073,N_23604,N_23016);
and U25074 (N_25074,N_23661,N_23342);
nand U25075 (N_25075,N_23626,N_24120);
nor U25076 (N_25076,N_24216,N_23683);
and U25077 (N_25077,N_24688,N_22673);
and U25078 (N_25078,N_24159,N_23203);
xnor U25079 (N_25079,N_23534,N_24256);
xor U25080 (N_25080,N_23085,N_23611);
nand U25081 (N_25081,N_23632,N_24800);
nor U25082 (N_25082,N_23348,N_23808);
and U25083 (N_25083,N_24316,N_24268);
xnor U25084 (N_25084,N_24129,N_22841);
xor U25085 (N_25085,N_24040,N_23303);
or U25086 (N_25086,N_23244,N_24108);
or U25087 (N_25087,N_22535,N_24939);
or U25088 (N_25088,N_24244,N_24818);
nor U25089 (N_25089,N_23382,N_23589);
nand U25090 (N_25090,N_23120,N_24437);
and U25091 (N_25091,N_24984,N_22739);
nand U25092 (N_25092,N_24602,N_22975);
nand U25093 (N_25093,N_24556,N_23436);
nor U25094 (N_25094,N_22536,N_23681);
or U25095 (N_25095,N_23282,N_23259);
or U25096 (N_25096,N_23748,N_24068);
nand U25097 (N_25097,N_23469,N_24724);
nor U25098 (N_25098,N_23034,N_23655);
and U25099 (N_25099,N_24368,N_22646);
xor U25100 (N_25100,N_24551,N_22515);
xnor U25101 (N_25101,N_23209,N_24049);
nand U25102 (N_25102,N_24929,N_22684);
and U25103 (N_25103,N_23642,N_24622);
nor U25104 (N_25104,N_24170,N_23430);
xnor U25105 (N_25105,N_23507,N_24107);
nor U25106 (N_25106,N_24557,N_22717);
nand U25107 (N_25107,N_22920,N_24858);
nor U25108 (N_25108,N_23722,N_24860);
nor U25109 (N_25109,N_23183,N_23163);
nand U25110 (N_25110,N_23361,N_24053);
or U25111 (N_25111,N_22959,N_24836);
xnor U25112 (N_25112,N_23738,N_24462);
and U25113 (N_25113,N_23620,N_22613);
and U25114 (N_25114,N_24751,N_23207);
and U25115 (N_25115,N_22782,N_24760);
nor U25116 (N_25116,N_24910,N_23696);
nor U25117 (N_25117,N_22922,N_24522);
and U25118 (N_25118,N_23110,N_24737);
xor U25119 (N_25119,N_24139,N_24283);
or U25120 (N_25120,N_22872,N_23520);
nor U25121 (N_25121,N_23297,N_24421);
and U25122 (N_25122,N_22763,N_23252);
and U25123 (N_25123,N_24231,N_24264);
and U25124 (N_25124,N_23771,N_22934);
or U25125 (N_25125,N_24355,N_22750);
nor U25126 (N_25126,N_24333,N_23652);
nor U25127 (N_25127,N_23556,N_22721);
nor U25128 (N_25128,N_23176,N_23964);
nor U25129 (N_25129,N_23923,N_24937);
and U25130 (N_25130,N_24900,N_23599);
nor U25131 (N_25131,N_22846,N_24851);
and U25132 (N_25132,N_22631,N_24917);
and U25133 (N_25133,N_23580,N_23331);
xor U25134 (N_25134,N_23879,N_23129);
and U25135 (N_25135,N_23052,N_23284);
nand U25136 (N_25136,N_23300,N_22714);
nand U25137 (N_25137,N_23811,N_23723);
nand U25138 (N_25138,N_24391,N_23093);
or U25139 (N_25139,N_24629,N_24665);
nand U25140 (N_25140,N_24744,N_24988);
and U25141 (N_25141,N_24440,N_24728);
and U25142 (N_25142,N_23253,N_23489);
xor U25143 (N_25143,N_24326,N_22858);
or U25144 (N_25144,N_23422,N_22789);
and U25145 (N_25145,N_24510,N_23858);
xor U25146 (N_25146,N_23118,N_23666);
nor U25147 (N_25147,N_22772,N_23967);
nand U25148 (N_25148,N_23558,N_24069);
nor U25149 (N_25149,N_24971,N_22741);
and U25150 (N_25150,N_22942,N_22812);
xnor U25151 (N_25151,N_24439,N_22776);
or U25152 (N_25152,N_23470,N_24203);
or U25153 (N_25153,N_24852,N_23610);
nor U25154 (N_25154,N_24627,N_24741);
and U25155 (N_25155,N_24786,N_23866);
or U25156 (N_25156,N_23979,N_22578);
or U25157 (N_25157,N_22790,N_24947);
or U25158 (N_25158,N_23930,N_24794);
and U25159 (N_25159,N_23555,N_23582);
nand U25160 (N_25160,N_23499,N_24038);
nor U25161 (N_25161,N_23783,N_24133);
xor U25162 (N_25162,N_24528,N_23103);
xor U25163 (N_25163,N_24403,N_24271);
nor U25164 (N_25164,N_23780,N_24389);
nand U25165 (N_25165,N_24790,N_23710);
and U25166 (N_25166,N_23365,N_24134);
or U25167 (N_25167,N_22711,N_23719);
nand U25168 (N_25168,N_23338,N_22754);
and U25169 (N_25169,N_23889,N_24762);
and U25170 (N_25170,N_23119,N_24384);
and U25171 (N_25171,N_24835,N_23003);
nand U25172 (N_25172,N_24619,N_23272);
xnor U25173 (N_25173,N_24405,N_24798);
nand U25174 (N_25174,N_24513,N_23640);
nand U25175 (N_25175,N_24346,N_22887);
and U25176 (N_25176,N_23168,N_23459);
and U25177 (N_25177,N_24088,N_22585);
and U25178 (N_25178,N_24493,N_22556);
or U25179 (N_25179,N_24165,N_24309);
or U25180 (N_25180,N_22979,N_24595);
and U25181 (N_25181,N_23020,N_23403);
xnor U25182 (N_25182,N_23588,N_24162);
nand U25183 (N_25183,N_23201,N_23862);
nand U25184 (N_25184,N_24207,N_24075);
nor U25185 (N_25185,N_23569,N_23954);
nand U25186 (N_25186,N_23148,N_23966);
nor U25187 (N_25187,N_24306,N_23420);
and U25188 (N_25188,N_22944,N_23087);
and U25189 (N_25189,N_24892,N_23375);
or U25190 (N_25190,N_22521,N_23318);
nand U25191 (N_25191,N_23302,N_23400);
xor U25192 (N_25192,N_23224,N_24985);
and U25193 (N_25193,N_22814,N_23464);
xor U25194 (N_25194,N_23397,N_24660);
or U25195 (N_25195,N_24432,N_23404);
or U25196 (N_25196,N_23200,N_23474);
nor U25197 (N_25197,N_23152,N_24248);
nand U25198 (N_25198,N_24518,N_22986);
xnor U25199 (N_25199,N_24716,N_23584);
and U25200 (N_25200,N_22677,N_23901);
and U25201 (N_25201,N_24621,N_23398);
and U25202 (N_25202,N_22725,N_24912);
nand U25203 (N_25203,N_24769,N_24696);
nand U25204 (N_25204,N_24184,N_23689);
or U25205 (N_25205,N_23065,N_24533);
xnor U25206 (N_25206,N_23706,N_24419);
or U25207 (N_25207,N_24146,N_22875);
nand U25208 (N_25208,N_23585,N_24630);
or U25209 (N_25209,N_24375,N_23601);
nand U25210 (N_25210,N_24546,N_23873);
and U25211 (N_25211,N_23231,N_23477);
nor U25212 (N_25212,N_24914,N_22893);
nor U25213 (N_25213,N_23098,N_23002);
or U25214 (N_25214,N_24549,N_24356);
nor U25215 (N_25215,N_24147,N_22913);
nand U25216 (N_25216,N_22925,N_23150);
and U25217 (N_25217,N_23344,N_23881);
and U25218 (N_25218,N_23454,N_24957);
or U25219 (N_25219,N_22784,N_24888);
or U25220 (N_25220,N_24076,N_23513);
nor U25221 (N_25221,N_24480,N_23432);
nand U25222 (N_25222,N_24915,N_23543);
xnor U25223 (N_25223,N_23294,N_24592);
nand U25224 (N_25224,N_23535,N_23532);
nor U25225 (N_25225,N_24583,N_23646);
xnor U25226 (N_25226,N_24830,N_24561);
nand U25227 (N_25227,N_22924,N_23312);
xnor U25228 (N_25228,N_24763,N_22757);
xor U25229 (N_25229,N_22502,N_23996);
or U25230 (N_25230,N_23055,N_23405);
nand U25231 (N_25231,N_23726,N_23968);
nor U25232 (N_25232,N_23144,N_24931);
or U25233 (N_25233,N_24580,N_24670);
xnor U25234 (N_25234,N_24459,N_24789);
nor U25235 (N_25235,N_23899,N_22670);
and U25236 (N_25236,N_24447,N_23806);
or U25237 (N_25237,N_22679,N_24575);
or U25238 (N_25238,N_23542,N_24065);
or U25239 (N_25239,N_23388,N_23686);
xor U25240 (N_25240,N_22598,N_24853);
nand U25241 (N_25241,N_23794,N_23606);
nand U25242 (N_25242,N_23143,N_23305);
nand U25243 (N_25243,N_24456,N_24785);
nor U25244 (N_25244,N_22962,N_23113);
nand U25245 (N_25245,N_22623,N_24024);
or U25246 (N_25246,N_24708,N_23735);
nor U25247 (N_25247,N_23512,N_22907);
nor U25248 (N_25248,N_23024,N_24274);
nor U25249 (N_25249,N_24436,N_24179);
xnor U25250 (N_25250,N_22947,N_23586);
nor U25251 (N_25251,N_24072,N_24093);
xor U25252 (N_25252,N_23492,N_23737);
or U25253 (N_25253,N_24647,N_24542);
or U25254 (N_25254,N_24396,N_24358);
and U25255 (N_25255,N_24449,N_23160);
or U25256 (N_25256,N_24702,N_24267);
nor U25257 (N_25257,N_22523,N_22654);
nor U25258 (N_25258,N_23406,N_24119);
nor U25259 (N_25259,N_23059,N_23978);
nor U25260 (N_25260,N_22614,N_24350);
nand U25261 (N_25261,N_24197,N_24987);
and U25262 (N_25262,N_24265,N_23347);
and U25263 (N_25263,N_24567,N_23634);
or U25264 (N_25264,N_24472,N_24523);
nor U25265 (N_25265,N_23078,N_22829);
or U25266 (N_25266,N_22870,N_24110);
and U25267 (N_25267,N_22565,N_23596);
and U25268 (N_25268,N_23579,N_23720);
nand U25269 (N_25269,N_24903,N_23465);
nand U25270 (N_25270,N_22674,N_23815);
and U25271 (N_25271,N_24840,N_24298);
and U25272 (N_25272,N_23725,N_23839);
and U25273 (N_25273,N_24156,N_22593);
and U25274 (N_25274,N_24047,N_22530);
xnor U25275 (N_25275,N_23445,N_23446);
nand U25276 (N_25276,N_23656,N_24682);
nor U25277 (N_25277,N_24579,N_23461);
nand U25278 (N_25278,N_23048,N_23731);
nand U25279 (N_25279,N_24431,N_23316);
or U25280 (N_25280,N_23266,N_22974);
and U25281 (N_25281,N_23644,N_24711);
and U25282 (N_25282,N_23473,N_23732);
nor U25283 (N_25283,N_24486,N_23145);
xnor U25284 (N_25284,N_24543,N_24981);
and U25285 (N_25285,N_22540,N_23935);
xnor U25286 (N_25286,N_22561,N_22939);
nand U25287 (N_25287,N_24923,N_24726);
xnor U25288 (N_25288,N_24877,N_24811);
xnor U25289 (N_25289,N_22764,N_23790);
or U25290 (N_25290,N_24948,N_22830);
xnor U25291 (N_25291,N_23685,N_24521);
nand U25292 (N_25292,N_22847,N_22647);
nor U25293 (N_25293,N_24752,N_23414);
nor U25294 (N_25294,N_22891,N_24189);
nand U25295 (N_25295,N_23332,N_23208);
nand U25296 (N_25296,N_24875,N_22943);
or U25297 (N_25297,N_22576,N_24640);
or U25298 (N_25298,N_23467,N_24232);
or U25299 (N_25299,N_23917,N_22538);
nor U25300 (N_25300,N_22849,N_23415);
nor U25301 (N_25301,N_23823,N_24911);
nand U25302 (N_25302,N_22729,N_24713);
xnor U25303 (N_25303,N_24245,N_24293);
nor U25304 (N_25304,N_24428,N_23945);
and U25305 (N_25305,N_23418,N_24690);
xor U25306 (N_25306,N_24791,N_22620);
xor U25307 (N_25307,N_24089,N_23924);
and U25308 (N_25308,N_22518,N_23817);
or U25309 (N_25309,N_24902,N_23670);
nor U25310 (N_25310,N_23974,N_23962);
and U25311 (N_25311,N_22886,N_23928);
and U25312 (N_25312,N_22510,N_24031);
or U25313 (N_25313,N_22899,N_23040);
xor U25314 (N_25314,N_22558,N_23758);
and U25315 (N_25315,N_23616,N_23619);
or U25316 (N_25316,N_22685,N_23759);
and U25317 (N_25317,N_22831,N_23158);
and U25318 (N_25318,N_22881,N_24259);
nor U25319 (N_25319,N_23883,N_23025);
or U25320 (N_25320,N_24961,N_24322);
xnor U25321 (N_25321,N_24394,N_24078);
nor U25322 (N_25322,N_24183,N_23907);
or U25323 (N_25323,N_24550,N_24132);
nand U25324 (N_25324,N_22906,N_22611);
or U25325 (N_25325,N_22588,N_24867);
or U25326 (N_25326,N_23522,N_23864);
nand U25327 (N_25327,N_22932,N_22501);
nor U25328 (N_25328,N_23615,N_23677);
or U25329 (N_25329,N_22767,N_23867);
nand U25330 (N_25330,N_22919,N_22534);
nand U25331 (N_25331,N_24152,N_23927);
or U25332 (N_25332,N_24974,N_22753);
or U25333 (N_25333,N_24768,N_23292);
xnor U25334 (N_25334,N_23963,N_23672);
xor U25335 (N_25335,N_22675,N_23653);
or U25336 (N_25336,N_23314,N_23607);
nand U25337 (N_25337,N_24534,N_23969);
and U25338 (N_25338,N_22823,N_24932);
or U25339 (N_25339,N_23383,N_23628);
nor U25340 (N_25340,N_24895,N_22871);
nand U25341 (N_25341,N_23339,N_23565);
nor U25342 (N_25342,N_24668,N_23280);
and U25343 (N_25343,N_22522,N_23086);
nand U25344 (N_25344,N_24692,N_23835);
and U25345 (N_25345,N_23659,N_23880);
xor U25346 (N_25346,N_23578,N_24275);
or U25347 (N_25347,N_24217,N_23358);
nand U25348 (N_25348,N_23976,N_22701);
or U25349 (N_25349,N_23852,N_22574);
xnor U25350 (N_25350,N_24699,N_24778);
or U25351 (N_25351,N_23301,N_24641);
nor U25352 (N_25352,N_23490,N_23320);
or U25353 (N_25353,N_22583,N_23495);
or U25354 (N_25354,N_23180,N_23981);
xor U25355 (N_25355,N_24829,N_23028);
nor U25356 (N_25356,N_24055,N_22559);
xnor U25357 (N_25357,N_24027,N_23570);
and U25358 (N_25358,N_24938,N_24648);
and U25359 (N_25359,N_24643,N_24176);
and U25360 (N_25360,N_24328,N_22539);
or U25361 (N_25361,N_24874,N_24584);
and U25362 (N_25362,N_24331,N_23286);
nand U25363 (N_25363,N_24504,N_22769);
and U25364 (N_25364,N_23088,N_23526);
or U25365 (N_25365,N_22743,N_23682);
xnor U25366 (N_25366,N_23360,N_24631);
or U25367 (N_25367,N_22520,N_24190);
or U25368 (N_25368,N_24524,N_22665);
or U25369 (N_25369,N_24153,N_24834);
and U25370 (N_25370,N_24986,N_23986);
xor U25371 (N_25371,N_24876,N_24940);
or U25372 (N_25372,N_23697,N_23931);
nor U25373 (N_25373,N_24291,N_22969);
and U25374 (N_25374,N_24680,N_24299);
and U25375 (N_25375,N_24393,N_22742);
nand U25376 (N_25376,N_24382,N_24497);
and U25377 (N_25377,N_22519,N_23549);
or U25378 (N_25378,N_23551,N_23396);
or U25379 (N_25379,N_24594,N_24701);
xor U25380 (N_25380,N_22809,N_22710);
nand U25381 (N_25381,N_22972,N_24857);
nand U25382 (N_25382,N_23226,N_22662);
and U25383 (N_25383,N_24882,N_22688);
and U25384 (N_25384,N_23271,N_23457);
or U25385 (N_25385,N_24843,N_22572);
nand U25386 (N_25386,N_23741,N_23739);
xnor U25387 (N_25387,N_24199,N_23898);
or U25388 (N_25388,N_24205,N_22822);
nand U25389 (N_25389,N_22640,N_22956);
or U25390 (N_25390,N_23516,N_23583);
and U25391 (N_25391,N_24126,N_23069);
nand U25392 (N_25392,N_23349,N_24715);
xor U25393 (N_25393,N_24413,N_23576);
and U25394 (N_25394,N_22587,N_23043);
and U25395 (N_25395,N_23929,N_22988);
or U25396 (N_25396,N_23437,N_24936);
or U25397 (N_25397,N_22938,N_24386);
nor U25398 (N_25398,N_23117,N_22946);
nand U25399 (N_25399,N_24343,N_23836);
or U25400 (N_25400,N_24022,N_23749);
and U25401 (N_25401,N_22514,N_23902);
and U25402 (N_25402,N_22866,N_24030);
xnor U25403 (N_25403,N_22616,N_24079);
and U25404 (N_25404,N_24097,N_23255);
nor U25405 (N_25405,N_22801,N_23251);
xnor U25406 (N_25406,N_24679,N_22724);
nand U25407 (N_25407,N_23536,N_22850);
and U25408 (N_25408,N_23204,N_24864);
xnor U25409 (N_25409,N_24397,N_24765);
nor U25410 (N_25410,N_23693,N_24211);
or U25411 (N_25411,N_24505,N_22880);
xor U25412 (N_25412,N_22595,N_23441);
xnor U25413 (N_25413,N_22723,N_24520);
nor U25414 (N_25414,N_24674,N_24388);
and U25415 (N_25415,N_24026,N_24337);
or U25416 (N_25416,N_23357,N_23667);
and U25417 (N_25417,N_23130,N_24560);
and U25418 (N_25418,N_23453,N_22702);
xnor U25419 (N_25419,N_24136,N_23840);
nand U25420 (N_25420,N_22612,N_23428);
or U25421 (N_25421,N_23376,N_24642);
xor U25422 (N_25422,N_24653,N_22781);
xnor U25423 (N_25423,N_23493,N_22639);
or U25424 (N_25424,N_24746,N_22885);
xor U25425 (N_25425,N_24967,N_24919);
nor U25426 (N_25426,N_23633,N_24399);
and U25427 (N_25427,N_24434,N_23949);
nor U25428 (N_25428,N_24001,N_24219);
or U25429 (N_25429,N_24398,N_23250);
nor U25430 (N_25430,N_24234,N_24458);
nand U25431 (N_25431,N_23031,N_22532);
and U25432 (N_25432,N_22936,N_22660);
nor U25433 (N_25433,N_24954,N_24354);
xor U25434 (N_25434,N_24638,N_22888);
nor U25435 (N_25435,N_22550,N_24086);
nand U25436 (N_25436,N_23149,N_23447);
nand U25437 (N_25437,N_24481,N_24793);
or U25438 (N_25438,N_23240,N_23997);
xnor U25439 (N_25439,N_22806,N_23472);
nand U25440 (N_25440,N_23784,N_24872);
xor U25441 (N_25441,N_24969,N_23765);
nand U25442 (N_25442,N_24982,N_24979);
and U25443 (N_25443,N_23621,N_23194);
nor U25444 (N_25444,N_24527,N_22989);
xor U25445 (N_25445,N_23393,N_23229);
or U25446 (N_25446,N_22599,N_23843);
or U25447 (N_25447,N_24347,N_24661);
nand U25448 (N_25448,N_23135,N_24624);
nor U25449 (N_25449,N_24103,N_23426);
nand U25450 (N_25450,N_23869,N_23351);
nor U25451 (N_25451,N_24395,N_23018);
xnor U25452 (N_25452,N_24406,N_24689);
nor U25453 (N_25453,N_23736,N_24048);
xor U25454 (N_25454,N_24130,N_23482);
or U25455 (N_25455,N_24066,N_22878);
and U25456 (N_25456,N_24144,N_24109);
and U25457 (N_25457,N_24727,N_24894);
nor U25458 (N_25458,N_24616,N_24059);
or U25459 (N_25459,N_24906,N_23392);
or U25460 (N_25460,N_23861,N_23548);
and U25461 (N_25461,N_24515,N_24576);
xnor U25462 (N_25462,N_23239,N_24342);
xor U25463 (N_25463,N_22577,N_23013);
nor U25464 (N_25464,N_24461,N_24297);
nor U25465 (N_25465,N_23826,N_24465);
nand U25466 (N_25466,N_23868,N_23322);
or U25467 (N_25467,N_23687,N_23313);
or U25468 (N_25468,N_23729,N_24060);
nand U25469 (N_25469,N_24927,N_24315);
and U25470 (N_25470,N_23246,N_24443);
xnor U25471 (N_25471,N_24250,N_22517);
and U25472 (N_25472,N_24883,N_23566);
and U25473 (N_25473,N_24673,N_22978);
nor U25474 (N_25474,N_24896,N_23989);
and U25475 (N_25475,N_24815,N_24280);
nand U25476 (N_25476,N_24823,N_24819);
and U25477 (N_25477,N_23236,N_22869);
and U25478 (N_25478,N_22626,N_23920);
xnor U25479 (N_25479,N_22797,N_24494);
nor U25480 (N_25480,N_23704,N_23744);
and U25481 (N_25481,N_24100,N_22964);
nor U25482 (N_25482,N_23166,N_24942);
xor U25483 (N_25483,N_23395,N_24817);
nand U25484 (N_25484,N_24338,N_24623);
nand U25485 (N_25485,N_23573,N_23264);
nor U25486 (N_25486,N_22821,N_23431);
or U25487 (N_25487,N_22622,N_24045);
nand U25488 (N_25488,N_22905,N_23530);
nand U25489 (N_25489,N_23010,N_23387);
and U25490 (N_25490,N_24169,N_23764);
xor U25491 (N_25491,N_23015,N_23455);
and U25492 (N_25492,N_24474,N_22633);
or U25493 (N_25493,N_24191,N_22828);
nor U25494 (N_25494,N_22526,N_24131);
xnor U25495 (N_25495,N_23401,N_24628);
xor U25496 (N_25496,N_24214,N_24087);
nor U25497 (N_25497,N_22715,N_24138);
nor U25498 (N_25498,N_24473,N_23485);
or U25499 (N_25499,N_23092,N_23014);
or U25500 (N_25500,N_22712,N_22661);
and U25501 (N_25501,N_24118,N_22752);
nor U25502 (N_25502,N_23064,N_23356);
or U25503 (N_25503,N_24198,N_23199);
nor U25504 (N_25504,N_24562,N_22504);
nor U25505 (N_25505,N_22923,N_22546);
and U25506 (N_25506,N_24904,N_23366);
or U25507 (N_25507,N_23631,N_24535);
xnor U25508 (N_25508,N_24841,N_24525);
nor U25509 (N_25509,N_23699,N_22687);
xnor U25510 (N_25510,N_24754,N_23757);
nor U25511 (N_25511,N_23218,N_23991);
nor U25512 (N_25512,N_24410,N_23848);
or U25513 (N_25513,N_23434,N_23756);
or U25514 (N_25514,N_24517,N_24539);
nor U25515 (N_25515,N_22896,N_22719);
nor U25516 (N_25516,N_24610,N_22512);
nand U25517 (N_25517,N_23123,N_23256);
nor U25518 (N_25518,N_24651,N_22503);
or U25519 (N_25519,N_23805,N_24907);
nor U25520 (N_25520,N_22590,N_23263);
xnor U25521 (N_25521,N_24412,N_23941);
and U25522 (N_25522,N_24869,N_23371);
or U25523 (N_25523,N_23335,N_23896);
nor U25524 (N_25524,N_24788,N_23503);
nand U25525 (N_25525,N_23115,N_23724);
nand U25526 (N_25526,N_22513,N_24700);
or U25527 (N_25527,N_23061,N_22579);
and U25528 (N_25528,N_23597,N_24901);
nor U25529 (N_25529,N_23279,N_24420);
xnor U25530 (N_25530,N_22537,N_24848);
or U25531 (N_25531,N_24009,N_24783);
or U25532 (N_25532,N_23527,N_22820);
xnor U25533 (N_25533,N_23851,N_23708);
xor U25534 (N_25534,N_23915,N_23101);
and U25535 (N_25535,N_24471,N_23125);
xor U25536 (N_25536,N_23175,N_24825);
nand U25537 (N_25537,N_22793,N_22985);
xnor U25538 (N_25538,N_23982,N_24757);
xor U25539 (N_25539,N_23773,N_24341);
or U25540 (N_25540,N_23450,N_23822);
nor U25541 (N_25541,N_24409,N_24884);
nand U25542 (N_25542,N_22791,N_22807);
xnor U25543 (N_25543,N_23916,N_23629);
and U25544 (N_25544,N_23959,N_23384);
xor U25545 (N_25545,N_24383,N_23701);
and U25546 (N_25546,N_24587,N_22529);
or U25547 (N_25547,N_23933,N_24284);
xnor U25548 (N_25548,N_24828,N_24324);
or U25549 (N_25549,N_22894,N_23062);
nor U25550 (N_25550,N_23813,N_24697);
nand U25551 (N_25551,N_22921,N_23700);
nand U25552 (N_25552,N_22663,N_24090);
nor U25553 (N_25553,N_24577,N_22580);
nor U25554 (N_25554,N_24508,N_24693);
and U25555 (N_25555,N_24287,N_23213);
or U25556 (N_25556,N_24028,N_23833);
or U25557 (N_25557,N_23821,N_23801);
nand U25558 (N_25558,N_23679,N_24099);
nand U25559 (N_25559,N_22861,N_22958);
nor U25560 (N_25560,N_24112,N_24304);
and U25561 (N_25561,N_24201,N_23487);
xor U25562 (N_25562,N_24224,N_24457);
or U25563 (N_25563,N_22904,N_22817);
nand U25564 (N_25564,N_23791,N_22606);
xnor U25565 (N_25565,N_24890,N_24188);
xnor U25566 (N_25566,N_24735,N_24430);
and U25567 (N_25567,N_24980,N_24253);
nor U25568 (N_25568,N_23641,N_23692);
and U25569 (N_25569,N_23402,N_24885);
and U25570 (N_25570,N_24320,N_24652);
nand U25571 (N_25571,N_23788,N_24196);
xnor U25572 (N_25572,N_24019,N_24373);
and U25573 (N_25573,N_24569,N_23798);
xnor U25574 (N_25574,N_23456,N_24334);
nand U25575 (N_25575,N_23273,N_22940);
nand U25576 (N_25576,N_22678,N_22668);
nor U25577 (N_25577,N_23021,N_23011);
nor U25578 (N_25578,N_24116,N_22569);
nand U25579 (N_25579,N_23391,N_23772);
nand U25580 (N_25580,N_24029,N_23705);
nor U25581 (N_25581,N_23367,N_22833);
and U25582 (N_25582,N_23539,N_24709);
nor U25583 (N_25583,N_22760,N_23324);
nand U25584 (N_25584,N_24739,N_24288);
or U25585 (N_25585,N_24808,N_24074);
nor U25586 (N_25586,N_24239,N_23241);
or U25587 (N_25587,N_24482,N_22770);
nor U25588 (N_25588,N_23892,N_24128);
nor U25589 (N_25589,N_23635,N_23460);
and U25590 (N_25590,N_24854,N_24096);
xor U25591 (N_25591,N_22856,N_24319);
or U25592 (N_25592,N_22970,N_22838);
and U25593 (N_25593,N_24532,N_23174);
nor U25594 (N_25594,N_23855,N_23545);
or U25595 (N_25595,N_23053,N_23664);
and U25596 (N_25596,N_24175,N_23519);
or U25597 (N_25597,N_23463,N_24366);
nor U25598 (N_25598,N_23462,N_23380);
or U25599 (N_25599,N_24318,N_24695);
xor U25600 (N_25600,N_23319,N_24991);
nand U25601 (N_25601,N_23567,N_23346);
and U25602 (N_25602,N_23745,N_22992);
nand U25603 (N_25603,N_22664,N_24844);
and U25604 (N_25604,N_23591,N_23425);
nand U25605 (N_25605,N_24033,N_24492);
nand U25606 (N_25606,N_24258,N_24155);
or U25607 (N_25607,N_23762,N_23734);
nor U25608 (N_25608,N_24983,N_23423);
xnor U25609 (N_25609,N_23825,N_23095);
xnor U25610 (N_25610,N_23691,N_24555);
or U25611 (N_25611,N_23270,N_24041);
nor U25612 (N_25612,N_24905,N_23197);
nor U25613 (N_25613,N_22656,N_24085);
nor U25614 (N_25614,N_23099,N_23173);
nand U25615 (N_25615,N_23364,N_24662);
xor U25616 (N_25616,N_23523,N_22744);
nor U25617 (N_25617,N_22780,N_23947);
xor U25618 (N_25618,N_22783,N_24977);
nor U25619 (N_25619,N_23538,N_23925);
nor U25620 (N_25620,N_24545,N_23560);
and U25621 (N_25621,N_23956,N_23777);
nand U25622 (N_25622,N_24913,N_22731);
and U25623 (N_25623,N_24285,N_23006);
nand U25624 (N_25624,N_24251,N_24633);
or U25625 (N_25625,N_22686,N_24442);
nand U25626 (N_25626,N_23466,N_24018);
and U25627 (N_25627,N_24672,N_23922);
nand U25628 (N_25628,N_24677,N_23045);
or U25629 (N_25629,N_24227,N_23853);
and U25630 (N_25630,N_24755,N_24174);
nand U25631 (N_25631,N_24770,N_24797);
xnor U25632 (N_25632,N_24742,N_24307);
or U25633 (N_25633,N_24934,N_24564);
and U25634 (N_25634,N_22728,N_22968);
nand U25635 (N_25635,N_23452,N_23496);
xnor U25636 (N_25636,N_24080,N_24998);
and U25637 (N_25637,N_23792,N_24776);
xor U25638 (N_25638,N_24740,N_23760);
nor U25639 (N_25639,N_23389,N_23486);
xnor U25640 (N_25640,N_23897,N_23715);
xnor U25641 (N_25641,N_22804,N_23448);
xor U25642 (N_25642,N_24946,N_24645);
and U25643 (N_25643,N_22657,N_24502);
xnor U25644 (N_25644,N_22736,N_24064);
nor U25645 (N_25645,N_24993,N_24956);
xor U25646 (N_25646,N_22643,N_24487);
nand U25647 (N_25647,N_24011,N_24747);
nand U25648 (N_25648,N_22683,N_24407);
nor U25649 (N_25649,N_23167,N_24092);
nand U25650 (N_25650,N_24290,N_23063);
nand U25651 (N_25651,N_24501,N_24833);
nand U25652 (N_25652,N_22799,N_22982);
or U25653 (N_25653,N_24611,N_23674);
nand U25654 (N_25654,N_23957,N_24476);
xnor U25655 (N_25655,N_23235,N_24454);
nor U25656 (N_25656,N_24469,N_24758);
xnor U25657 (N_25657,N_23830,N_24847);
and U25658 (N_25658,N_23872,N_22527);
xor U25659 (N_25659,N_22787,N_24636);
nand U25660 (N_25660,N_22645,N_24816);
or U25661 (N_25661,N_24866,N_23262);
and U25662 (N_25662,N_24590,N_23958);
nand U25663 (N_25663,N_23803,N_23654);
nand U25664 (N_25664,N_24016,N_23484);
xnor U25665 (N_25665,N_23254,N_23122);
nor U25666 (N_25666,N_23857,N_24141);
xnor U25667 (N_25667,N_23926,N_23521);
and U25668 (N_25668,N_23709,N_23295);
nor U25669 (N_25669,N_24111,N_24598);
nand U25670 (N_25670,N_23439,N_24200);
nand U25671 (N_25671,N_22773,N_22890);
nand U25672 (N_25672,N_24962,N_23531);
or U25673 (N_25673,N_22607,N_24764);
or U25674 (N_25674,N_24371,N_24423);
or U25675 (N_25675,N_22835,N_23444);
and U25676 (N_25676,N_24260,N_24717);
and U25677 (N_25677,N_24292,N_23315);
nor U25678 (N_25678,N_24361,N_23820);
nand U25679 (N_25679,N_22591,N_24731);
nor U25680 (N_25680,N_24380,N_23598);
and U25681 (N_25681,N_22884,N_23903);
nor U25682 (N_25682,N_24143,N_23651);
nand U25683 (N_25683,N_22573,N_22650);
xnor U25684 (N_25684,N_24363,N_24246);
or U25685 (N_25685,N_22624,N_23993);
nor U25686 (N_25686,N_23593,N_24970);
nor U25687 (N_25687,N_23504,N_24123);
and U25688 (N_25688,N_22629,N_22843);
xor U25689 (N_25689,N_24639,N_24221);
and U25690 (N_25690,N_24351,N_22563);
nand U25691 (N_25691,N_23665,N_22926);
and U25692 (N_25692,N_24964,N_23937);
or U25693 (N_25693,N_24344,N_23107);
nor U25694 (N_25694,N_24429,N_24687);
nand U25695 (N_25695,N_24773,N_23278);
and U25696 (N_25696,N_23952,N_22722);
xor U25697 (N_25697,N_23429,N_23763);
nand U25698 (N_25698,N_23362,N_24707);
nor U25699 (N_25699,N_23786,N_23106);
or U25700 (N_25700,N_22691,N_24925);
nor U25701 (N_25701,N_23054,N_24955);
and U25702 (N_25702,N_22911,N_24308);
nor U25703 (N_25703,N_23189,N_23819);
and U25704 (N_25704,N_24262,N_24704);
nor U25705 (N_25705,N_23230,N_22796);
or U25706 (N_25706,N_24761,N_23073);
nor U25707 (N_25707,N_22965,N_24418);
nand U25708 (N_25708,N_24336,N_22740);
and U25709 (N_25709,N_22732,N_24738);
xor U25710 (N_25710,N_23260,N_23837);
nand U25711 (N_25711,N_23828,N_24124);
nand U25712 (N_25712,N_23277,N_23577);
and U25713 (N_25713,N_22889,N_23355);
nor U25714 (N_25714,N_23609,N_23592);
nand U25715 (N_25715,N_23544,N_22993);
nand U25716 (N_25716,N_24416,N_23097);
and U25717 (N_25717,N_23678,N_22990);
nor U25718 (N_25718,N_23938,N_24973);
nand U25719 (N_25719,N_22848,N_23849);
nand U25720 (N_25720,N_23283,N_24182);
nand U25721 (N_25721,N_23443,N_24488);
and U25722 (N_25722,N_23793,N_23386);
nor U25723 (N_25723,N_24374,N_22954);
nand U25724 (N_25724,N_22862,N_24812);
xor U25725 (N_25725,N_24020,N_23035);
xor U25726 (N_25726,N_24604,N_23041);
nor U25727 (N_25727,N_23071,N_22998);
nor U25728 (N_25728,N_22692,N_24782);
or U25729 (N_25729,N_23091,N_23658);
or U25730 (N_25730,N_22589,N_23990);
xor U25731 (N_25731,N_23850,N_23156);
or U25732 (N_25732,N_23195,N_23227);
or U25733 (N_25733,N_22601,N_23860);
nor U25734 (N_25734,N_22690,N_24222);
nand U25735 (N_25735,N_24614,N_24233);
nand U25736 (N_25736,N_22933,N_23111);
and U25737 (N_25737,N_24489,N_22524);
xor U25738 (N_25738,N_22805,N_23217);
nor U25739 (N_25739,N_24511,N_24496);
or U25740 (N_25740,N_22638,N_24270);
xor U25741 (N_25741,N_22818,N_22533);
nand U25742 (N_25742,N_22726,N_24255);
and U25743 (N_25743,N_22666,N_23269);
nor U25744 (N_25744,N_24151,N_23912);
or U25745 (N_25745,N_23712,N_24591);
nor U25746 (N_25746,N_24228,N_24479);
xor U25747 (N_25747,N_24603,N_23904);
nand U25748 (N_25748,N_24411,N_23942);
xor U25749 (N_25749,N_23752,N_23128);
nor U25750 (N_25750,N_23970,N_22525);
nor U25751 (N_25751,N_24166,N_24478);
and U25752 (N_25752,N_22581,N_24725);
nand U25753 (N_25753,N_24050,N_23219);
xnor U25754 (N_25754,N_23228,N_23352);
or U25755 (N_25755,N_24404,N_23707);
xnor U25756 (N_25756,N_23971,N_23036);
and U25757 (N_25757,N_24625,N_24637);
and U25758 (N_25758,N_24862,N_24252);
and U25759 (N_25759,N_23797,N_22718);
xor U25760 (N_25760,N_23648,N_24873);
and U25761 (N_25761,N_23076,N_23182);
and U25762 (N_25762,N_23481,N_23824);
or U25763 (N_25763,N_22854,N_22778);
xnor U25764 (N_25764,N_23755,N_24718);
or U25765 (N_25765,N_23274,N_22615);
and U25766 (N_25766,N_22751,N_24194);
or U25767 (N_25767,N_24278,N_23618);
nor U25768 (N_25768,N_23876,N_24994);
xor U25769 (N_25769,N_22935,N_23554);
or U25770 (N_25770,N_22617,N_23435);
and U25771 (N_25771,N_23992,N_23141);
nand U25772 (N_25772,N_23716,N_23753);
xor U25773 (N_25773,N_24563,N_23847);
and U25774 (N_25774,N_23878,N_23131);
nand U25775 (N_25775,N_23802,N_23308);
and U25776 (N_25776,N_22816,N_23385);
and U25777 (N_25777,N_23243,N_24323);
and U25778 (N_25778,N_24753,N_24348);
and U25779 (N_25779,N_24477,N_23146);
or U25780 (N_25780,N_24613,N_22775);
xnor U25781 (N_25781,N_22570,N_24849);
or U25782 (N_25782,N_22937,N_22758);
nand U25783 (N_25783,N_22651,N_24172);
nor U25784 (N_25784,N_23727,N_24667);
nand U25785 (N_25785,N_22803,N_22542);
nand U25786 (N_25786,N_23795,N_22950);
nor U25787 (N_25787,N_24588,N_22826);
nor U25788 (N_25788,N_23787,N_23698);
or U25789 (N_25789,N_23804,N_23563);
nor U25790 (N_25790,N_24918,N_23624);
and U25791 (N_25791,N_24002,N_22541);
nand U25792 (N_25792,N_22506,N_22669);
nor U25793 (N_25793,N_24710,N_23877);
xnor U25794 (N_25794,N_24792,N_24659);
xnor U25795 (N_25795,N_23442,N_23440);
nor U25796 (N_25796,N_22705,N_22766);
nand U25797 (N_25797,N_24846,N_24723);
nor U25798 (N_25798,N_24279,N_22774);
nand U25799 (N_25799,N_23185,N_23309);
nor U25800 (N_25800,N_24538,N_22682);
and U25801 (N_25801,N_24332,N_24444);
and U25802 (N_25802,N_24070,N_23663);
nand U25803 (N_25803,N_23136,N_22859);
xnor U25804 (N_25804,N_24073,N_24922);
and U25805 (N_25805,N_24756,N_24826);
or U25806 (N_25806,N_23537,N_23740);
xor U25807 (N_25807,N_23169,N_24999);
xor U25808 (N_25808,N_22908,N_24295);
or U25809 (N_25809,N_23424,N_23026);
or U25810 (N_25810,N_24325,N_22844);
or U25811 (N_25811,N_23502,N_22798);
nor U25812 (N_25812,N_23854,N_24150);
xnor U25813 (N_25813,N_23094,N_24898);
nand U25814 (N_25814,N_24435,N_24015);
nand U25815 (N_25815,N_24056,N_24046);
nor U25816 (N_25816,N_24114,N_23438);
nor U25817 (N_25817,N_23234,N_24750);
nand U25818 (N_25818,N_22627,N_22961);
and U25819 (N_25819,N_23550,N_24805);
and U25820 (N_25820,N_23188,N_22973);
nand U25821 (N_25821,N_24061,N_23785);
or U25822 (N_25822,N_23181,N_23162);
nand U25823 (N_25823,N_23000,N_24335);
nor U25824 (N_25824,N_23409,N_23033);
xnor U25825 (N_25825,N_23680,N_23998);
or U25826 (N_25826,N_23410,N_23399);
nand U25827 (N_25827,N_24814,N_24626);
nor U25828 (N_25828,N_23751,N_22777);
nand U25829 (N_25829,N_24212,N_24968);
nor U25830 (N_25830,N_23865,N_23225);
nand U25831 (N_25831,N_23275,N_22505);
or U25832 (N_25832,N_24657,N_23810);
nor U25833 (N_25833,N_23032,N_23750);
xor U25834 (N_25834,N_24506,N_23614);
or U25835 (N_25835,N_23863,N_24035);
nor U25836 (N_25836,N_24730,N_22852);
nor U25837 (N_25837,N_23050,N_24039);
xnor U25838 (N_25838,N_23695,N_22873);
xnor U25839 (N_25839,N_24425,N_23468);
nor U25840 (N_25840,N_23172,N_24365);
nand U25841 (N_25841,N_23408,N_23814);
or U25842 (N_25842,N_22704,N_24161);
nand U25843 (N_25843,N_23210,N_24081);
nor U25844 (N_25844,N_23728,N_23215);
nand U25845 (N_25845,N_23547,N_23296);
and U25846 (N_25846,N_23844,N_24058);
nor U25847 (N_25847,N_24837,N_22902);
and U25848 (N_25848,N_23381,N_24303);
nand U25849 (N_25849,N_24377,N_24158);
and U25850 (N_25850,N_23505,N_24552);
nand U25851 (N_25851,N_24536,N_24051);
or U25852 (N_25852,N_24286,N_22910);
or U25853 (N_25853,N_24281,N_24658);
nor U25854 (N_25854,N_24930,N_24597);
nand U25855 (N_25855,N_22600,N_22901);
nor U25856 (N_25856,N_23044,N_24663);
or U25857 (N_25857,N_24992,N_23630);
or U25858 (N_25858,N_23572,N_24554);
xnor U25859 (N_25859,N_23761,N_23192);
xor U25860 (N_25860,N_23528,N_23330);
nor U25861 (N_25861,N_23211,N_22952);
nand U25862 (N_25862,N_24145,N_23882);
nand U25863 (N_25863,N_23184,N_24581);
nor U25864 (N_25864,N_24678,N_23557);
nor U25865 (N_25865,N_24113,N_23782);
nand U25866 (N_25866,N_24868,N_23575);
xor U25867 (N_25867,N_23498,N_23205);
and U25868 (N_25868,N_23307,N_24122);
and U25869 (N_25869,N_24438,N_24607);
nor U25870 (N_25870,N_22916,N_22971);
and U25871 (N_25871,N_23132,N_23413);
xnor U25872 (N_25872,N_22699,N_24054);
nand U25873 (N_25873,N_23500,N_24787);
nand U25874 (N_25874,N_23953,N_23887);
and U25875 (N_25875,N_24213,N_22696);
and U25876 (N_25876,N_24296,N_23747);
and U25877 (N_25877,N_24586,N_22941);
and U25878 (N_25878,N_24427,N_24599);
and U25879 (N_25879,N_23378,N_24490);
nor U25880 (N_25880,N_24007,N_24767);
xnor U25881 (N_25881,N_24548,N_23799);
nor U25882 (N_25882,N_22592,N_24605);
nor U25883 (N_25883,N_23343,N_24340);
nor U25884 (N_25884,N_23874,N_23645);
and U25885 (N_25885,N_24734,N_24148);
nand U25886 (N_25886,N_24157,N_24101);
and U25887 (N_25887,N_24367,N_23746);
nor U25888 (N_25888,N_24450,N_23553);
nand U25889 (N_25889,N_23121,N_23612);
xor U25890 (N_25890,N_22749,N_22957);
xnor U25891 (N_25891,N_22547,N_23975);
and U25892 (N_25892,N_24446,N_24242);
or U25893 (N_25893,N_24719,N_24247);
and U25894 (N_25894,N_24305,N_23509);
or U25895 (N_25895,N_22659,N_24052);
nor U25896 (N_25896,N_23258,N_23327);
nor U25897 (N_25897,N_24989,N_22516);
xor U25898 (N_25898,N_22903,N_24390);
nor U25899 (N_25899,N_23987,N_24289);
nor U25900 (N_25900,N_24571,N_23829);
xnor U25901 (N_25901,N_22735,N_24417);
or U25902 (N_25902,N_22557,N_22765);
nand U25903 (N_25903,N_23476,N_24796);
and U25904 (N_25904,N_23248,N_23198);
nand U25905 (N_25905,N_24928,N_23994);
xor U25906 (N_25906,N_23574,N_24240);
xnor U25907 (N_25907,N_23304,N_24951);
nor U25908 (N_25908,N_24722,N_23832);
or U25909 (N_25909,N_22644,N_23291);
and U25910 (N_25910,N_22876,N_24241);
and U25911 (N_25911,N_24683,N_24733);
xnor U25912 (N_25912,N_23345,N_23265);
xnor U25913 (N_25913,N_23070,N_22883);
nand U25914 (N_25914,N_24484,N_24831);
xnor U25915 (N_25915,N_22655,N_23427);
xnor U25916 (N_25916,N_22983,N_22918);
xor U25917 (N_25917,N_23116,N_24300);
and U25918 (N_25918,N_23187,N_24317);
and U25919 (N_25919,N_24558,N_24220);
nor U25920 (N_25920,N_22619,N_23005);
nand U25921 (N_25921,N_23058,N_24042);
nor U25922 (N_25922,N_23066,N_24071);
or U25923 (N_25923,N_24426,N_24574);
and U25924 (N_25924,N_22981,N_24589);
nand U25925 (N_25925,N_24424,N_23261);
nand U25926 (N_25926,N_24014,N_24063);
or U25927 (N_25927,N_24357,N_22955);
nand U25928 (N_25928,N_22794,N_22855);
nand U25929 (N_25929,N_22845,N_24339);
and U25930 (N_25930,N_22602,N_24966);
or U25931 (N_25931,N_24329,N_23138);
and U25932 (N_25932,N_22892,N_24950);
nor U25933 (N_25933,N_24415,N_23713);
xor U25934 (N_25934,N_23662,N_24615);
nand U25935 (N_25935,N_24933,N_24330);
or U25936 (N_25936,N_22681,N_22867);
or U25937 (N_25937,N_23323,N_23084);
xnor U25938 (N_25938,N_23845,N_23299);
or U25939 (N_25939,N_23961,N_24491);
and U25940 (N_25940,N_23105,N_23370);
nor U25941 (N_25941,N_22716,N_23223);
nand U25942 (N_25942,N_22996,N_23222);
or U25943 (N_25943,N_23766,N_23743);
nor U25944 (N_25944,N_23306,N_23046);
and U25945 (N_25945,N_24230,N_24466);
and U25946 (N_25946,N_24173,N_23004);
nor U25947 (N_25947,N_24378,N_23433);
nand U25948 (N_25948,N_24777,N_22756);
xnor U25949 (N_25949,N_23511,N_24171);
xor U25950 (N_25950,N_24210,N_24972);
nand U25951 (N_25951,N_23170,N_24686);
and U25952 (N_25952,N_24023,N_22977);
xnor U25953 (N_25953,N_24807,N_23096);
or U25954 (N_25954,N_24685,N_22567);
nand U25955 (N_25955,N_24531,N_24870);
xor U25956 (N_25956,N_24414,N_23276);
and U25957 (N_25957,N_24944,N_23711);
and U25958 (N_25958,N_23908,N_23326);
nand U25959 (N_25959,N_23374,N_24507);
or U25960 (N_25960,N_22994,N_24802);
xor U25961 (N_25961,N_22792,N_22915);
and U25962 (N_25962,N_23909,N_22551);
nand U25963 (N_25963,N_24675,N_23079);
and U25964 (N_25964,N_23017,N_23089);
and U25965 (N_25965,N_23077,N_22637);
nor U25966 (N_25966,N_23100,N_23491);
and U25967 (N_25967,N_24978,N_22507);
nor U25968 (N_25968,N_22698,N_23220);
nor U25969 (N_25969,N_22734,N_24202);
and U25970 (N_25970,N_22694,N_23702);
xor U25971 (N_25971,N_24712,N_24578);
xnor U25972 (N_25972,N_24498,N_22995);
nand U25973 (N_25973,N_23451,N_24400);
and U25974 (N_25974,N_24804,N_24408);
and U25975 (N_25975,N_23965,N_24311);
xor U25976 (N_25976,N_24495,N_24077);
nor U25977 (N_25977,N_23671,N_24839);
nor U25978 (N_25978,N_22999,N_23675);
or U25979 (N_25979,N_22874,N_22700);
and U25980 (N_25980,N_23478,N_22582);
or U25981 (N_25981,N_24891,N_22618);
xnor U25982 (N_25982,N_24780,N_24514);
nor U25983 (N_25983,N_23807,N_24163);
nor U25984 (N_25984,N_23009,N_24084);
xor U25985 (N_25985,N_22610,N_24036);
and U25986 (N_25986,N_24945,N_22808);
or U25987 (N_25987,N_24485,N_22545);
nor U25988 (N_25988,N_23134,N_24083);
xor U25989 (N_25989,N_22597,N_22649);
and U25990 (N_25990,N_22706,N_22951);
xnor U25991 (N_25991,N_23552,N_23980);
or U25992 (N_25992,N_24899,N_22813);
nand U25993 (N_25993,N_23894,N_23249);
nor U25994 (N_25994,N_22827,N_24596);
xnor U25995 (N_25995,N_23562,N_22648);
xor U25996 (N_25996,N_23419,N_24091);
nand U25997 (N_25997,N_24464,N_24483);
nand U25998 (N_25998,N_22839,N_22860);
or U25999 (N_25999,N_22966,N_23019);
nand U26000 (N_26000,N_23369,N_23796);
and U26001 (N_26001,N_24671,N_23524);
and U26002 (N_26002,N_23140,N_22596);
xnor U26003 (N_26003,N_23684,N_24729);
or U26004 (N_26004,N_24082,N_22621);
or U26005 (N_26005,N_22991,N_24381);
and U26006 (N_26006,N_24463,N_24345);
xor U26007 (N_26007,N_24387,N_22531);
nor U26008 (N_26008,N_23075,N_23001);
xnor U26009 (N_26009,N_24650,N_24392);
or U26010 (N_26010,N_23186,N_23694);
or U26011 (N_26011,N_24960,N_24582);
nand U26012 (N_26012,N_24908,N_23082);
or U26013 (N_26013,N_23068,N_24547);
and U26014 (N_26014,N_22553,N_22762);
or U26015 (N_26015,N_23350,N_23449);
and U26016 (N_26016,N_24106,N_22897);
or U26017 (N_26017,N_23595,N_22713);
nand U26018 (N_26018,N_23060,N_23153);
and U26019 (N_26019,N_22746,N_23960);
or U26020 (N_26020,N_24568,N_23212);
nand U26021 (N_26021,N_23885,N_23056);
nor U26022 (N_26022,N_22562,N_24952);
xor U26023 (N_26023,N_23841,N_22737);
nor U26024 (N_26024,N_23257,N_22953);
and U26025 (N_26025,N_22967,N_24142);
nand U26026 (N_26026,N_23074,N_24475);
nor U26027 (N_26027,N_23587,N_22834);
nand U26028 (N_26028,N_24453,N_23875);
and U26029 (N_26029,N_23471,N_23972);
xnor U26030 (N_26030,N_23714,N_22575);
or U26031 (N_26031,N_23411,N_24691);
xnor U26032 (N_26032,N_24012,N_24277);
xnor U26033 (N_26033,N_24608,N_23285);
nor U26034 (N_26034,N_23730,N_22697);
nor U26035 (N_26035,N_24401,N_23950);
and U26036 (N_26036,N_23647,N_24537);
nand U26037 (N_26037,N_24360,N_23072);
or U26038 (N_26038,N_23581,N_22603);
xor U26039 (N_26039,N_22586,N_23948);
or U26040 (N_26040,N_24634,N_23372);
and U26041 (N_26041,N_24249,N_24104);
and U26042 (N_26042,N_23109,N_23157);
nor U26043 (N_26043,N_23859,N_22800);
xor U26044 (N_26044,N_24887,N_24620);
nand U26045 (N_26045,N_22945,N_24310);
xnor U26046 (N_26046,N_22931,N_24654);
xor U26047 (N_26047,N_23458,N_23768);
or U26048 (N_26048,N_24115,N_24379);
and U26049 (N_26049,N_23407,N_22863);
or U26050 (N_26050,N_24195,N_23638);
nor U26051 (N_26051,N_23905,N_23893);
xnor U26052 (N_26052,N_23057,N_24646);
nor U26053 (N_26053,N_22549,N_24470);
nand U26054 (N_26054,N_22584,N_24540);
nand U26055 (N_26055,N_24206,N_24021);
nand U26056 (N_26056,N_24871,N_23178);
xnor U26057 (N_26057,N_22652,N_22914);
or U26058 (N_26058,N_24881,N_23910);
nand U26059 (N_26059,N_23870,N_23946);
nand U26060 (N_26060,N_24010,N_23533);
nor U26061 (N_26061,N_22795,N_23884);
xnor U26062 (N_26062,N_24714,N_23703);
or U26063 (N_26063,N_22693,N_23943);
nor U26064 (N_26064,N_24095,N_23317);
and U26065 (N_26065,N_22976,N_22785);
nor U26066 (N_26066,N_24649,N_24125);
nand U26067 (N_26067,N_22544,N_24460);
nand U26068 (N_26068,N_23494,N_23417);
nor U26069 (N_26069,N_24920,N_24208);
xor U26070 (N_26070,N_24223,N_23999);
nor U26071 (N_26071,N_22635,N_23669);
nand U26072 (N_26072,N_23081,N_23027);
nor U26073 (N_26073,N_24953,N_24585);
nor U26074 (N_26074,N_23767,N_22882);
nand U26075 (N_26075,N_23779,N_23900);
and U26076 (N_26076,N_24570,N_24529);
and U26077 (N_26077,N_23127,N_22802);
or U26078 (N_26078,N_23287,N_23781);
xnor U26079 (N_26079,N_23165,N_24813);
nand U26080 (N_26080,N_24799,N_24949);
nand U26081 (N_26081,N_22837,N_23514);
xnor U26082 (N_26082,N_24235,N_22695);
xor U26083 (N_26083,N_24448,N_23561);
nand U26084 (N_26084,N_22825,N_24861);
nor U26085 (N_26085,N_24236,N_24455);
nor U26086 (N_26086,N_22779,N_24105);
or U26087 (N_26087,N_24795,N_24736);
nor U26088 (N_26088,N_24301,N_24821);
or U26089 (N_26089,N_23818,N_23939);
nor U26090 (N_26090,N_24385,N_23617);
nor U26091 (N_26091,N_22511,N_23718);
and U26092 (N_26092,N_23919,N_24774);
nand U26093 (N_26093,N_23657,N_23789);
xor U26094 (N_26094,N_24032,N_23337);
and U26095 (N_26095,N_23333,N_22771);
or U26096 (N_26096,N_22566,N_24921);
or U26097 (N_26097,N_22709,N_24926);
or U26098 (N_26098,N_24897,N_23102);
nor U26099 (N_26099,N_22672,N_24263);
and U26100 (N_26100,N_24618,N_24732);
nand U26101 (N_26101,N_24990,N_24362);
nand U26102 (N_26102,N_22609,N_24273);
xnor U26103 (N_26103,N_22929,N_24766);
nand U26104 (N_26104,N_23022,N_24544);
or U26105 (N_26105,N_24748,N_23353);
and U26106 (N_26106,N_24721,N_23636);
and U26107 (N_26107,N_22879,N_24192);
nor U26108 (N_26108,N_24468,N_24565);
or U26109 (N_26109,N_23037,N_24238);
and U26110 (N_26110,N_24017,N_23080);
nand U26111 (N_26111,N_24094,N_24327);
xnor U26112 (N_26112,N_24149,N_23827);
nor U26113 (N_26113,N_23977,N_24806);
nand U26114 (N_26114,N_22927,N_24218);
and U26115 (N_26115,N_24941,N_23564);
or U26116 (N_26116,N_22671,N_23340);
and U26117 (N_26117,N_24243,N_22625);
or U26118 (N_26118,N_24452,N_24370);
or U26119 (N_26119,N_23660,N_22509);
xnor U26120 (N_26120,N_22948,N_24043);
and U26121 (N_26121,N_23108,N_24215);
nand U26122 (N_26122,N_23030,N_22594);
nand U26123 (N_26123,N_24959,N_23518);
xnor U26124 (N_26124,N_24566,N_23831);
and U26125 (N_26125,N_24880,N_23190);
xnor U26126 (N_26126,N_22768,N_24004);
xor U26127 (N_26127,N_23488,N_24025);
nand U26128 (N_26128,N_24749,N_23546);
nand U26129 (N_26129,N_23298,N_23891);
and U26130 (N_26130,N_22864,N_23047);
nor U26131 (N_26131,N_22632,N_23196);
xor U26132 (N_26132,N_24775,N_23206);
and U26133 (N_26133,N_24121,N_23594);
nor U26134 (N_26134,N_24655,N_23049);
and U26135 (N_26135,N_23268,N_24669);
and U26136 (N_26136,N_24684,N_22987);
xnor U26137 (N_26137,N_23321,N_23985);
nor U26138 (N_26138,N_24666,N_24916);
nand U26139 (N_26139,N_24137,N_22689);
nand U26140 (N_26140,N_24102,N_24167);
or U26141 (N_26141,N_23151,N_22543);
nand U26142 (N_26142,N_23501,N_24187);
nor U26143 (N_26143,N_24656,N_23394);
and U26144 (N_26144,N_24359,N_23124);
xnor U26145 (N_26145,N_23668,N_23247);
nand U26146 (N_26146,N_24140,N_24266);
nand U26147 (N_26147,N_24294,N_22761);
or U26148 (N_26148,N_23515,N_24771);
or U26149 (N_26149,N_23506,N_23913);
xor U26150 (N_26150,N_22667,N_22997);
or U26151 (N_26151,N_24759,N_23238);
or U26152 (N_26152,N_22571,N_23988);
nand U26153 (N_26153,N_23379,N_24062);
and U26154 (N_26154,N_24376,N_24676);
xor U26155 (N_26155,N_22658,N_24644);
and U26156 (N_26156,N_24364,N_23232);
nor U26157 (N_26157,N_22630,N_23613);
or U26158 (N_26158,N_24632,N_23416);
or U26159 (N_26159,N_24832,N_23479);
xnor U26160 (N_26160,N_23932,N_24177);
and U26161 (N_26161,N_24781,N_22730);
nand U26162 (N_26162,N_23325,N_24445);
nand U26163 (N_26163,N_22898,N_22865);
or U26164 (N_26164,N_22786,N_23568);
and U26165 (N_26165,N_23267,N_24842);
nand U26166 (N_26166,N_24706,N_24606);
and U26167 (N_26167,N_23622,N_23769);
nand U26168 (N_26168,N_23846,N_22832);
nand U26169 (N_26169,N_24067,N_24572);
and U26170 (N_26170,N_24559,N_24530);
xor U26171 (N_26171,N_23973,N_23754);
xor U26172 (N_26172,N_24824,N_23637);
nand U26173 (N_26173,N_24720,N_24261);
or U26174 (N_26174,N_24703,N_22868);
xor U26175 (N_26175,N_23541,N_23354);
or U26176 (N_26176,N_24850,N_24745);
or U26177 (N_26177,N_23159,N_24694);
xnor U26178 (N_26178,N_24503,N_22836);
nand U26179 (N_26179,N_24975,N_23147);
or U26180 (N_26180,N_22628,N_23171);
nor U26181 (N_26181,N_22853,N_23838);
nand U26182 (N_26182,N_23164,N_24225);
and U26183 (N_26183,N_23112,N_24743);
nand U26184 (N_26184,N_24044,N_23717);
xor U26185 (N_26185,N_24349,N_23191);
nor U26186 (N_26186,N_23193,N_24965);
nor U26187 (N_26187,N_23914,N_23038);
nand U26188 (N_26188,N_23288,N_23816);
or U26189 (N_26189,N_23895,N_22949);
or U26190 (N_26190,N_24845,N_22851);
xnor U26191 (N_26191,N_24801,N_22500);
nand U26192 (N_26192,N_23918,N_23368);
and U26193 (N_26193,N_24313,N_23842);
and U26194 (N_26194,N_23983,N_23281);
and U26195 (N_26195,N_23329,N_23517);
and U26196 (N_26196,N_24117,N_23733);
xor U26197 (N_26197,N_24803,N_24996);
or U26198 (N_26198,N_23603,N_24314);
and U26199 (N_26199,N_23812,N_22676);
nand U26200 (N_26200,N_22747,N_22960);
or U26201 (N_26201,N_24441,N_23627);
nor U26202 (N_26202,N_22912,N_23155);
nand U26203 (N_26203,N_23890,N_23083);
nand U26204 (N_26204,N_23559,N_24193);
and U26205 (N_26205,N_23161,N_23936);
xor U26206 (N_26206,N_24924,N_23023);
and U26207 (N_26207,N_23497,N_23363);
nand U26208 (N_26208,N_24681,N_24772);
nor U26209 (N_26209,N_22840,N_24372);
and U26210 (N_26210,N_23310,N_24003);
and U26211 (N_26211,N_22641,N_22984);
nand U26212 (N_26212,N_23137,N_22703);
nand U26213 (N_26213,N_23311,N_23051);
nor U26214 (N_26214,N_22727,N_24433);
nor U26215 (N_26215,N_22811,N_24178);
or U26216 (N_26216,N_24013,N_22788);
or U26217 (N_26217,N_24856,N_24402);
nor U26218 (N_26218,N_23007,N_24369);
and U26219 (N_26219,N_24008,N_24353);
nand U26220 (N_26220,N_24526,N_23373);
or U26221 (N_26221,N_23289,N_22842);
xnor U26222 (N_26222,N_24467,N_23336);
nand U26223 (N_26223,N_23510,N_23412);
nor U26224 (N_26224,N_24893,N_24963);
and U26225 (N_26225,N_24512,N_24181);
xor U26226 (N_26226,N_23650,N_24600);
nor U26227 (N_26227,N_24422,N_24204);
and U26228 (N_26228,N_24229,N_22755);
nand U26229 (N_26229,N_23377,N_24995);
or U26230 (N_26230,N_22554,N_23856);
nor U26231 (N_26231,N_22824,N_22642);
xor U26232 (N_26232,N_23126,N_24006);
nand U26233 (N_26233,N_22680,N_23955);
nor U26234 (N_26234,N_23995,N_24878);
nand U26235 (N_26235,N_24185,N_23571);
xnor U26236 (N_26236,N_22917,N_23214);
or U26237 (N_26237,N_24664,N_24612);
or U26238 (N_26238,N_22720,N_24127);
xnor U26239 (N_26239,N_24135,N_22819);
xor U26240 (N_26240,N_22653,N_23525);
nand U26241 (N_26241,N_24886,N_24820);
xor U26242 (N_26242,N_23540,N_23039);
nor U26243 (N_26243,N_23328,N_23643);
or U26244 (N_26244,N_22552,N_24519);
or U26245 (N_26245,N_24958,N_22928);
xor U26246 (N_26246,N_23951,N_24997);
and U26247 (N_26247,N_24302,N_24180);
xor U26248 (N_26248,N_24282,N_22605);
or U26249 (N_26249,N_22564,N_23390);
or U26250 (N_26250,N_24544,N_23954);
and U26251 (N_26251,N_23069,N_24318);
nand U26252 (N_26252,N_23793,N_23532);
or U26253 (N_26253,N_24093,N_23512);
nor U26254 (N_26254,N_24675,N_22902);
or U26255 (N_26255,N_23766,N_22622);
xor U26256 (N_26256,N_22526,N_23816);
and U26257 (N_26257,N_23308,N_23503);
nand U26258 (N_26258,N_23626,N_23920);
nor U26259 (N_26259,N_24356,N_24308);
or U26260 (N_26260,N_22546,N_23331);
xnor U26261 (N_26261,N_24410,N_23135);
xnor U26262 (N_26262,N_22637,N_22607);
nor U26263 (N_26263,N_24852,N_23930);
nor U26264 (N_26264,N_23759,N_24379);
nand U26265 (N_26265,N_24121,N_23961);
or U26266 (N_26266,N_23946,N_24893);
xnor U26267 (N_26267,N_23587,N_22593);
nor U26268 (N_26268,N_23521,N_22991);
nand U26269 (N_26269,N_23347,N_23859);
xor U26270 (N_26270,N_24412,N_23875);
xnor U26271 (N_26271,N_24233,N_23612);
and U26272 (N_26272,N_23145,N_22595);
nand U26273 (N_26273,N_23918,N_23486);
nand U26274 (N_26274,N_24611,N_24444);
nand U26275 (N_26275,N_22508,N_23561);
and U26276 (N_26276,N_23478,N_24061);
nand U26277 (N_26277,N_23402,N_23758);
or U26278 (N_26278,N_24157,N_23291);
nand U26279 (N_26279,N_24955,N_23202);
and U26280 (N_26280,N_23490,N_23802);
nand U26281 (N_26281,N_22711,N_23052);
or U26282 (N_26282,N_23092,N_24061);
and U26283 (N_26283,N_23297,N_24903);
or U26284 (N_26284,N_24849,N_24952);
nor U26285 (N_26285,N_24787,N_22812);
xnor U26286 (N_26286,N_22572,N_23773);
or U26287 (N_26287,N_22532,N_24390);
or U26288 (N_26288,N_24828,N_23411);
xnor U26289 (N_26289,N_23589,N_23629);
nor U26290 (N_26290,N_24686,N_24850);
nand U26291 (N_26291,N_24263,N_23261);
nor U26292 (N_26292,N_22643,N_23465);
nand U26293 (N_26293,N_22527,N_22790);
nand U26294 (N_26294,N_24330,N_22894);
and U26295 (N_26295,N_23418,N_22756);
nand U26296 (N_26296,N_22815,N_23197);
nor U26297 (N_26297,N_24381,N_24508);
nand U26298 (N_26298,N_22723,N_23115);
and U26299 (N_26299,N_24093,N_23622);
and U26300 (N_26300,N_23077,N_24612);
and U26301 (N_26301,N_24179,N_23330);
or U26302 (N_26302,N_23521,N_23692);
xnor U26303 (N_26303,N_22944,N_24287);
nand U26304 (N_26304,N_23925,N_24661);
and U26305 (N_26305,N_24349,N_23027);
and U26306 (N_26306,N_24624,N_24057);
xor U26307 (N_26307,N_22571,N_23386);
xor U26308 (N_26308,N_24677,N_24685);
or U26309 (N_26309,N_22615,N_24354);
nor U26310 (N_26310,N_22806,N_24880);
or U26311 (N_26311,N_24304,N_24392);
and U26312 (N_26312,N_24059,N_24225);
xnor U26313 (N_26313,N_23754,N_24366);
nor U26314 (N_26314,N_23450,N_24566);
xor U26315 (N_26315,N_22624,N_24045);
and U26316 (N_26316,N_23493,N_23649);
and U26317 (N_26317,N_23743,N_23964);
nand U26318 (N_26318,N_23978,N_23357);
nor U26319 (N_26319,N_23141,N_24136);
or U26320 (N_26320,N_23811,N_24798);
nand U26321 (N_26321,N_24983,N_22668);
xnor U26322 (N_26322,N_24696,N_23386);
or U26323 (N_26323,N_24870,N_22669);
nor U26324 (N_26324,N_22978,N_24622);
and U26325 (N_26325,N_23121,N_23461);
or U26326 (N_26326,N_24402,N_23409);
and U26327 (N_26327,N_24727,N_24581);
nand U26328 (N_26328,N_23623,N_24180);
nor U26329 (N_26329,N_23927,N_24472);
nand U26330 (N_26330,N_24364,N_22625);
or U26331 (N_26331,N_24366,N_23285);
nand U26332 (N_26332,N_22833,N_23027);
or U26333 (N_26333,N_23216,N_24249);
nor U26334 (N_26334,N_23442,N_23055);
xnor U26335 (N_26335,N_24394,N_23887);
nand U26336 (N_26336,N_24004,N_24233);
xnor U26337 (N_26337,N_23699,N_24356);
or U26338 (N_26338,N_23737,N_23491);
or U26339 (N_26339,N_23746,N_24302);
nand U26340 (N_26340,N_23456,N_23514);
xor U26341 (N_26341,N_22918,N_23948);
or U26342 (N_26342,N_24332,N_23783);
nand U26343 (N_26343,N_24650,N_24230);
nor U26344 (N_26344,N_22840,N_23873);
xnor U26345 (N_26345,N_23153,N_23305);
or U26346 (N_26346,N_23555,N_23258);
nor U26347 (N_26347,N_23529,N_24294);
nand U26348 (N_26348,N_23239,N_22958);
xnor U26349 (N_26349,N_23361,N_23862);
or U26350 (N_26350,N_23772,N_24735);
and U26351 (N_26351,N_24727,N_24987);
or U26352 (N_26352,N_23408,N_24873);
or U26353 (N_26353,N_23009,N_24568);
or U26354 (N_26354,N_23924,N_23374);
xor U26355 (N_26355,N_22970,N_23898);
nand U26356 (N_26356,N_23554,N_23508);
nand U26357 (N_26357,N_22578,N_24265);
xnor U26358 (N_26358,N_22786,N_24309);
xor U26359 (N_26359,N_24705,N_24717);
nand U26360 (N_26360,N_24035,N_22704);
and U26361 (N_26361,N_24387,N_23686);
or U26362 (N_26362,N_24486,N_24776);
or U26363 (N_26363,N_24133,N_24519);
and U26364 (N_26364,N_22663,N_24484);
nand U26365 (N_26365,N_22850,N_24240);
nor U26366 (N_26366,N_23797,N_23046);
xnor U26367 (N_26367,N_24036,N_23604);
and U26368 (N_26368,N_23849,N_22893);
or U26369 (N_26369,N_23834,N_23626);
nand U26370 (N_26370,N_22511,N_22931);
or U26371 (N_26371,N_23663,N_23729);
and U26372 (N_26372,N_23490,N_24348);
and U26373 (N_26373,N_24594,N_24017);
xor U26374 (N_26374,N_24250,N_23237);
or U26375 (N_26375,N_24815,N_22702);
nand U26376 (N_26376,N_24845,N_23950);
and U26377 (N_26377,N_23579,N_24887);
and U26378 (N_26378,N_24124,N_24683);
nor U26379 (N_26379,N_23945,N_22575);
or U26380 (N_26380,N_23393,N_22598);
and U26381 (N_26381,N_24416,N_22981);
xnor U26382 (N_26382,N_22978,N_23230);
and U26383 (N_26383,N_24305,N_24264);
and U26384 (N_26384,N_24093,N_23828);
or U26385 (N_26385,N_24264,N_24687);
or U26386 (N_26386,N_24985,N_23749);
and U26387 (N_26387,N_24428,N_22821);
nand U26388 (N_26388,N_23837,N_24281);
and U26389 (N_26389,N_24532,N_22562);
xnor U26390 (N_26390,N_23265,N_22909);
and U26391 (N_26391,N_22914,N_23601);
nand U26392 (N_26392,N_22679,N_23706);
and U26393 (N_26393,N_24737,N_23016);
nor U26394 (N_26394,N_24175,N_24552);
or U26395 (N_26395,N_22955,N_24909);
nand U26396 (N_26396,N_24640,N_23331);
nand U26397 (N_26397,N_24501,N_23419);
nand U26398 (N_26398,N_23405,N_23295);
or U26399 (N_26399,N_24902,N_24509);
nor U26400 (N_26400,N_24253,N_22719);
nand U26401 (N_26401,N_23976,N_22641);
nand U26402 (N_26402,N_24778,N_22643);
or U26403 (N_26403,N_22855,N_23773);
nor U26404 (N_26404,N_24268,N_23038);
nand U26405 (N_26405,N_22661,N_22606);
nor U26406 (N_26406,N_24838,N_22964);
nand U26407 (N_26407,N_24104,N_24101);
xnor U26408 (N_26408,N_23723,N_23270);
or U26409 (N_26409,N_24213,N_23708);
and U26410 (N_26410,N_24338,N_23133);
nand U26411 (N_26411,N_24849,N_24174);
nor U26412 (N_26412,N_24548,N_23331);
nand U26413 (N_26413,N_23689,N_24358);
or U26414 (N_26414,N_23354,N_23410);
and U26415 (N_26415,N_23604,N_24930);
xnor U26416 (N_26416,N_24791,N_23812);
nand U26417 (N_26417,N_22765,N_24505);
or U26418 (N_26418,N_22535,N_22590);
nor U26419 (N_26419,N_24295,N_23774);
or U26420 (N_26420,N_24592,N_22842);
or U26421 (N_26421,N_23926,N_24131);
xnor U26422 (N_26422,N_24860,N_24831);
nand U26423 (N_26423,N_22575,N_24705);
or U26424 (N_26424,N_24533,N_24708);
or U26425 (N_26425,N_23029,N_23099);
and U26426 (N_26426,N_24240,N_23312);
xnor U26427 (N_26427,N_22842,N_23977);
or U26428 (N_26428,N_22747,N_22557);
or U26429 (N_26429,N_22700,N_23855);
nor U26430 (N_26430,N_23393,N_22945);
nor U26431 (N_26431,N_23432,N_23965);
xor U26432 (N_26432,N_24104,N_23274);
xnor U26433 (N_26433,N_23766,N_24936);
or U26434 (N_26434,N_23446,N_23526);
nand U26435 (N_26435,N_24214,N_23405);
and U26436 (N_26436,N_23892,N_24822);
and U26437 (N_26437,N_22773,N_23668);
xnor U26438 (N_26438,N_24077,N_24070);
and U26439 (N_26439,N_22788,N_23503);
nand U26440 (N_26440,N_23513,N_24492);
nor U26441 (N_26441,N_23610,N_23383);
nor U26442 (N_26442,N_23914,N_23516);
nor U26443 (N_26443,N_24789,N_23533);
nor U26444 (N_26444,N_23164,N_23502);
nand U26445 (N_26445,N_22621,N_24348);
xnor U26446 (N_26446,N_24553,N_24525);
nand U26447 (N_26447,N_22756,N_23380);
xnor U26448 (N_26448,N_24611,N_24936);
xnor U26449 (N_26449,N_23876,N_24306);
and U26450 (N_26450,N_22634,N_23337);
and U26451 (N_26451,N_23301,N_24046);
or U26452 (N_26452,N_23349,N_23185);
xor U26453 (N_26453,N_24053,N_23356);
and U26454 (N_26454,N_24063,N_24837);
nand U26455 (N_26455,N_23720,N_24744);
and U26456 (N_26456,N_24024,N_23361);
nor U26457 (N_26457,N_24605,N_23195);
xnor U26458 (N_26458,N_23493,N_23880);
and U26459 (N_26459,N_23172,N_22929);
xnor U26460 (N_26460,N_22899,N_23986);
or U26461 (N_26461,N_23397,N_23702);
or U26462 (N_26462,N_23542,N_23793);
xnor U26463 (N_26463,N_23341,N_22896);
nand U26464 (N_26464,N_23677,N_24430);
nand U26465 (N_26465,N_24349,N_22729);
and U26466 (N_26466,N_24597,N_24744);
xor U26467 (N_26467,N_22661,N_24714);
nor U26468 (N_26468,N_24771,N_24337);
xnor U26469 (N_26469,N_22673,N_24216);
or U26470 (N_26470,N_23152,N_22553);
nand U26471 (N_26471,N_24471,N_23894);
xnor U26472 (N_26472,N_24160,N_24081);
and U26473 (N_26473,N_24003,N_24701);
xnor U26474 (N_26474,N_23035,N_24056);
nor U26475 (N_26475,N_22904,N_22650);
nor U26476 (N_26476,N_23312,N_23431);
or U26477 (N_26477,N_24908,N_22778);
nand U26478 (N_26478,N_23144,N_23759);
nor U26479 (N_26479,N_23794,N_24105);
xor U26480 (N_26480,N_23300,N_24716);
nor U26481 (N_26481,N_22695,N_24662);
nor U26482 (N_26482,N_24410,N_23535);
or U26483 (N_26483,N_23348,N_24796);
or U26484 (N_26484,N_23597,N_24045);
and U26485 (N_26485,N_22962,N_24263);
and U26486 (N_26486,N_24861,N_23840);
xnor U26487 (N_26487,N_23901,N_24002);
or U26488 (N_26488,N_23227,N_23880);
or U26489 (N_26489,N_23401,N_23871);
xor U26490 (N_26490,N_23657,N_24104);
nor U26491 (N_26491,N_23383,N_24423);
xor U26492 (N_26492,N_24519,N_23962);
nor U26493 (N_26493,N_22617,N_22817);
or U26494 (N_26494,N_24389,N_24665);
or U26495 (N_26495,N_24024,N_24628);
nand U26496 (N_26496,N_24187,N_23356);
nor U26497 (N_26497,N_22782,N_24279);
or U26498 (N_26498,N_23795,N_24350);
and U26499 (N_26499,N_22692,N_24070);
or U26500 (N_26500,N_22715,N_23905);
or U26501 (N_26501,N_23358,N_22976);
nand U26502 (N_26502,N_23139,N_23109);
nand U26503 (N_26503,N_22911,N_24637);
and U26504 (N_26504,N_24588,N_22796);
or U26505 (N_26505,N_24644,N_24346);
and U26506 (N_26506,N_24802,N_24770);
nand U26507 (N_26507,N_23261,N_24726);
nor U26508 (N_26508,N_22691,N_22850);
or U26509 (N_26509,N_23747,N_24148);
nand U26510 (N_26510,N_23303,N_23654);
xor U26511 (N_26511,N_24337,N_23118);
and U26512 (N_26512,N_23302,N_24397);
xor U26513 (N_26513,N_24360,N_24562);
and U26514 (N_26514,N_23469,N_23448);
xor U26515 (N_26515,N_23386,N_24744);
nand U26516 (N_26516,N_23244,N_24074);
and U26517 (N_26517,N_24311,N_23381);
nand U26518 (N_26518,N_23989,N_22697);
and U26519 (N_26519,N_24471,N_24973);
nor U26520 (N_26520,N_22857,N_24364);
xnor U26521 (N_26521,N_24934,N_23985);
nor U26522 (N_26522,N_22589,N_24661);
nand U26523 (N_26523,N_24994,N_22802);
or U26524 (N_26524,N_23230,N_23563);
or U26525 (N_26525,N_24839,N_24345);
xor U26526 (N_26526,N_24087,N_24967);
nand U26527 (N_26527,N_22541,N_23897);
or U26528 (N_26528,N_23662,N_22722);
nor U26529 (N_26529,N_23746,N_24524);
or U26530 (N_26530,N_24738,N_23600);
or U26531 (N_26531,N_24320,N_23099);
nor U26532 (N_26532,N_23487,N_23395);
or U26533 (N_26533,N_23395,N_23799);
nor U26534 (N_26534,N_23797,N_22972);
or U26535 (N_26535,N_23365,N_22544);
xnor U26536 (N_26536,N_22721,N_24822);
xor U26537 (N_26537,N_22872,N_24650);
or U26538 (N_26538,N_24595,N_23856);
or U26539 (N_26539,N_23061,N_22618);
xor U26540 (N_26540,N_23501,N_23074);
nand U26541 (N_26541,N_23606,N_22869);
nor U26542 (N_26542,N_24465,N_23569);
or U26543 (N_26543,N_23209,N_22691);
nor U26544 (N_26544,N_24687,N_24884);
xor U26545 (N_26545,N_24738,N_24207);
nand U26546 (N_26546,N_23130,N_22820);
nor U26547 (N_26547,N_22634,N_23232);
or U26548 (N_26548,N_23883,N_23106);
or U26549 (N_26549,N_24503,N_23610);
nand U26550 (N_26550,N_24472,N_23413);
nand U26551 (N_26551,N_23149,N_24819);
nand U26552 (N_26552,N_24870,N_22784);
xor U26553 (N_26553,N_22953,N_22647);
or U26554 (N_26554,N_22610,N_23926);
and U26555 (N_26555,N_24448,N_22581);
nand U26556 (N_26556,N_22702,N_23041);
nor U26557 (N_26557,N_23209,N_24139);
or U26558 (N_26558,N_23541,N_24405);
or U26559 (N_26559,N_24021,N_24269);
nand U26560 (N_26560,N_23386,N_24995);
and U26561 (N_26561,N_24957,N_22532);
nand U26562 (N_26562,N_22605,N_24513);
and U26563 (N_26563,N_22858,N_22933);
and U26564 (N_26564,N_24941,N_22856);
nor U26565 (N_26565,N_24285,N_24267);
nand U26566 (N_26566,N_22672,N_23462);
and U26567 (N_26567,N_23621,N_23397);
nor U26568 (N_26568,N_23428,N_23491);
and U26569 (N_26569,N_24410,N_24764);
or U26570 (N_26570,N_23869,N_24173);
nor U26571 (N_26571,N_23403,N_23901);
nor U26572 (N_26572,N_23913,N_23236);
nor U26573 (N_26573,N_22771,N_23457);
xor U26574 (N_26574,N_22783,N_24885);
or U26575 (N_26575,N_24793,N_24895);
nand U26576 (N_26576,N_22900,N_24345);
or U26577 (N_26577,N_22787,N_22559);
nand U26578 (N_26578,N_23025,N_24941);
nand U26579 (N_26579,N_23970,N_23713);
and U26580 (N_26580,N_23300,N_23051);
nor U26581 (N_26581,N_23608,N_24484);
nor U26582 (N_26582,N_22754,N_24213);
xor U26583 (N_26583,N_24568,N_23675);
nor U26584 (N_26584,N_23431,N_24870);
or U26585 (N_26585,N_23447,N_23122);
or U26586 (N_26586,N_23713,N_23212);
nand U26587 (N_26587,N_24794,N_24472);
xor U26588 (N_26588,N_24826,N_24955);
xor U26589 (N_26589,N_24199,N_23241);
or U26590 (N_26590,N_24415,N_23617);
or U26591 (N_26591,N_24981,N_22551);
and U26592 (N_26592,N_22937,N_24315);
or U26593 (N_26593,N_23512,N_24929);
and U26594 (N_26594,N_24710,N_24458);
or U26595 (N_26595,N_24691,N_23422);
and U26596 (N_26596,N_24421,N_23425);
or U26597 (N_26597,N_23920,N_23715);
and U26598 (N_26598,N_23217,N_24808);
and U26599 (N_26599,N_22577,N_24111);
nor U26600 (N_26600,N_23350,N_24574);
nand U26601 (N_26601,N_24678,N_23206);
xor U26602 (N_26602,N_23730,N_24396);
or U26603 (N_26603,N_23072,N_22533);
or U26604 (N_26604,N_22944,N_23194);
nand U26605 (N_26605,N_24795,N_22988);
and U26606 (N_26606,N_24105,N_23632);
xnor U26607 (N_26607,N_22572,N_24761);
nand U26608 (N_26608,N_24173,N_23998);
nand U26609 (N_26609,N_23844,N_23023);
nor U26610 (N_26610,N_24771,N_23854);
xnor U26611 (N_26611,N_23891,N_22781);
nor U26612 (N_26612,N_23384,N_23467);
nor U26613 (N_26613,N_24093,N_24183);
or U26614 (N_26614,N_23314,N_24435);
nand U26615 (N_26615,N_23197,N_24105);
nand U26616 (N_26616,N_24955,N_23722);
or U26617 (N_26617,N_22708,N_23951);
or U26618 (N_26618,N_23163,N_23168);
nor U26619 (N_26619,N_23096,N_24166);
nor U26620 (N_26620,N_24415,N_24106);
or U26621 (N_26621,N_23364,N_23147);
or U26622 (N_26622,N_24536,N_24335);
or U26623 (N_26623,N_24704,N_23037);
nor U26624 (N_26624,N_24374,N_23819);
nor U26625 (N_26625,N_23200,N_24623);
or U26626 (N_26626,N_22646,N_22689);
nand U26627 (N_26627,N_23047,N_24561);
and U26628 (N_26628,N_22737,N_24784);
nand U26629 (N_26629,N_23708,N_24748);
and U26630 (N_26630,N_23125,N_23041);
or U26631 (N_26631,N_22703,N_23274);
nand U26632 (N_26632,N_23191,N_22649);
or U26633 (N_26633,N_23712,N_23937);
nand U26634 (N_26634,N_23562,N_24880);
and U26635 (N_26635,N_23751,N_24783);
or U26636 (N_26636,N_22535,N_24477);
nand U26637 (N_26637,N_24992,N_24817);
nand U26638 (N_26638,N_23346,N_24374);
nand U26639 (N_26639,N_22878,N_22640);
nor U26640 (N_26640,N_24744,N_24159);
and U26641 (N_26641,N_22787,N_23576);
or U26642 (N_26642,N_24331,N_22728);
xnor U26643 (N_26643,N_22821,N_23251);
or U26644 (N_26644,N_24693,N_22915);
and U26645 (N_26645,N_22622,N_24862);
xor U26646 (N_26646,N_22985,N_23114);
and U26647 (N_26647,N_24582,N_23811);
nand U26648 (N_26648,N_23526,N_24472);
xnor U26649 (N_26649,N_24248,N_22581);
or U26650 (N_26650,N_22995,N_24966);
and U26651 (N_26651,N_24924,N_22554);
nand U26652 (N_26652,N_24991,N_24759);
and U26653 (N_26653,N_23649,N_24449);
or U26654 (N_26654,N_24697,N_23040);
xnor U26655 (N_26655,N_23130,N_23132);
nor U26656 (N_26656,N_24650,N_24426);
nor U26657 (N_26657,N_23105,N_23051);
and U26658 (N_26658,N_24080,N_22732);
xnor U26659 (N_26659,N_24565,N_22986);
nor U26660 (N_26660,N_23665,N_24400);
or U26661 (N_26661,N_22505,N_22830);
xnor U26662 (N_26662,N_23547,N_23379);
xor U26663 (N_26663,N_23494,N_23584);
and U26664 (N_26664,N_22508,N_24080);
or U26665 (N_26665,N_23655,N_22833);
nand U26666 (N_26666,N_23609,N_23719);
nor U26667 (N_26667,N_22546,N_24573);
and U26668 (N_26668,N_23584,N_23860);
xnor U26669 (N_26669,N_24930,N_23072);
nand U26670 (N_26670,N_23734,N_24768);
nand U26671 (N_26671,N_23158,N_24705);
or U26672 (N_26672,N_23353,N_24223);
xor U26673 (N_26673,N_23904,N_24473);
nor U26674 (N_26674,N_22581,N_24707);
xor U26675 (N_26675,N_23218,N_24213);
or U26676 (N_26676,N_23891,N_24539);
nor U26677 (N_26677,N_24793,N_24746);
and U26678 (N_26678,N_22879,N_23463);
nor U26679 (N_26679,N_22829,N_24541);
nand U26680 (N_26680,N_23732,N_23780);
or U26681 (N_26681,N_23308,N_24908);
nand U26682 (N_26682,N_24444,N_22721);
and U26683 (N_26683,N_24708,N_23001);
xor U26684 (N_26684,N_24070,N_22622);
xnor U26685 (N_26685,N_23262,N_24524);
and U26686 (N_26686,N_23782,N_24329);
nor U26687 (N_26687,N_22520,N_23130);
nor U26688 (N_26688,N_22806,N_23286);
or U26689 (N_26689,N_23950,N_23130);
nor U26690 (N_26690,N_23302,N_24251);
xnor U26691 (N_26691,N_23941,N_23328);
xor U26692 (N_26692,N_23829,N_23261);
nor U26693 (N_26693,N_22989,N_23449);
or U26694 (N_26694,N_23477,N_23276);
xnor U26695 (N_26695,N_23839,N_23776);
xor U26696 (N_26696,N_23786,N_22736);
and U26697 (N_26697,N_23425,N_24911);
nor U26698 (N_26698,N_23701,N_24613);
or U26699 (N_26699,N_23629,N_23579);
xnor U26700 (N_26700,N_23943,N_22597);
nand U26701 (N_26701,N_22625,N_23152);
and U26702 (N_26702,N_24366,N_23840);
and U26703 (N_26703,N_24120,N_24166);
nand U26704 (N_26704,N_22800,N_24343);
nand U26705 (N_26705,N_24544,N_23058);
and U26706 (N_26706,N_23041,N_24766);
and U26707 (N_26707,N_22813,N_23193);
nor U26708 (N_26708,N_24930,N_23469);
and U26709 (N_26709,N_24615,N_24367);
nor U26710 (N_26710,N_23390,N_24164);
or U26711 (N_26711,N_23563,N_24035);
nor U26712 (N_26712,N_24109,N_22746);
nand U26713 (N_26713,N_23491,N_22507);
xor U26714 (N_26714,N_22676,N_23594);
nor U26715 (N_26715,N_24430,N_23315);
nor U26716 (N_26716,N_24143,N_24416);
and U26717 (N_26717,N_22541,N_24419);
nand U26718 (N_26718,N_23596,N_22839);
or U26719 (N_26719,N_23366,N_24665);
nand U26720 (N_26720,N_24687,N_24815);
nand U26721 (N_26721,N_23142,N_23148);
nor U26722 (N_26722,N_23638,N_23072);
or U26723 (N_26723,N_24851,N_24636);
and U26724 (N_26724,N_24020,N_24829);
or U26725 (N_26725,N_24709,N_23854);
nor U26726 (N_26726,N_23604,N_23156);
and U26727 (N_26727,N_22878,N_24336);
nand U26728 (N_26728,N_22658,N_24593);
and U26729 (N_26729,N_24096,N_24004);
nand U26730 (N_26730,N_22820,N_22572);
nand U26731 (N_26731,N_23358,N_24331);
xnor U26732 (N_26732,N_22563,N_24066);
xor U26733 (N_26733,N_23253,N_22731);
or U26734 (N_26734,N_23562,N_23838);
or U26735 (N_26735,N_24626,N_23968);
nor U26736 (N_26736,N_24134,N_23297);
and U26737 (N_26737,N_24734,N_24871);
and U26738 (N_26738,N_23670,N_24746);
nand U26739 (N_26739,N_24398,N_24633);
xor U26740 (N_26740,N_23222,N_23198);
and U26741 (N_26741,N_22670,N_24307);
or U26742 (N_26742,N_24753,N_22700);
nor U26743 (N_26743,N_24026,N_24070);
or U26744 (N_26744,N_24171,N_24490);
and U26745 (N_26745,N_23559,N_23637);
and U26746 (N_26746,N_23678,N_23469);
xnor U26747 (N_26747,N_23705,N_24134);
nand U26748 (N_26748,N_22553,N_24212);
nand U26749 (N_26749,N_24824,N_22949);
or U26750 (N_26750,N_23307,N_23057);
xor U26751 (N_26751,N_23223,N_22708);
nand U26752 (N_26752,N_24071,N_24877);
nor U26753 (N_26753,N_22548,N_24301);
and U26754 (N_26754,N_23474,N_23549);
or U26755 (N_26755,N_22853,N_22730);
xor U26756 (N_26756,N_22686,N_22993);
xnor U26757 (N_26757,N_24636,N_22780);
and U26758 (N_26758,N_24873,N_23778);
and U26759 (N_26759,N_24839,N_23352);
nor U26760 (N_26760,N_24644,N_23047);
and U26761 (N_26761,N_23272,N_24551);
xnor U26762 (N_26762,N_24672,N_24854);
xnor U26763 (N_26763,N_23258,N_22605);
xnor U26764 (N_26764,N_24548,N_24241);
nor U26765 (N_26765,N_22982,N_24442);
nand U26766 (N_26766,N_23098,N_24489);
xor U26767 (N_26767,N_24171,N_22922);
nor U26768 (N_26768,N_24145,N_23537);
xor U26769 (N_26769,N_24808,N_22961);
or U26770 (N_26770,N_24215,N_22750);
and U26771 (N_26771,N_22653,N_24255);
xnor U26772 (N_26772,N_23631,N_23126);
xnor U26773 (N_26773,N_22896,N_23610);
nor U26774 (N_26774,N_23964,N_24985);
nor U26775 (N_26775,N_23811,N_24436);
nor U26776 (N_26776,N_23513,N_23017);
xor U26777 (N_26777,N_24160,N_23615);
or U26778 (N_26778,N_22692,N_24799);
nand U26779 (N_26779,N_22728,N_23596);
nand U26780 (N_26780,N_23012,N_23153);
nand U26781 (N_26781,N_24628,N_24701);
and U26782 (N_26782,N_24456,N_24743);
nand U26783 (N_26783,N_24992,N_23309);
or U26784 (N_26784,N_23191,N_23973);
xnor U26785 (N_26785,N_24455,N_23699);
or U26786 (N_26786,N_24674,N_22510);
nor U26787 (N_26787,N_22520,N_23690);
nor U26788 (N_26788,N_23044,N_24733);
nor U26789 (N_26789,N_24558,N_23331);
xnor U26790 (N_26790,N_24545,N_23295);
nand U26791 (N_26791,N_22761,N_24607);
nor U26792 (N_26792,N_24897,N_22930);
or U26793 (N_26793,N_23357,N_24428);
nand U26794 (N_26794,N_22651,N_24310);
nand U26795 (N_26795,N_23716,N_24583);
xnor U26796 (N_26796,N_22835,N_22944);
or U26797 (N_26797,N_23530,N_23207);
xor U26798 (N_26798,N_23753,N_24896);
xor U26799 (N_26799,N_23727,N_22592);
or U26800 (N_26800,N_24128,N_23052);
nor U26801 (N_26801,N_23886,N_24081);
or U26802 (N_26802,N_22994,N_24196);
xnor U26803 (N_26803,N_24976,N_24319);
and U26804 (N_26804,N_23431,N_24224);
or U26805 (N_26805,N_23336,N_24777);
nand U26806 (N_26806,N_23586,N_24856);
xor U26807 (N_26807,N_24139,N_23286);
and U26808 (N_26808,N_24498,N_23863);
nand U26809 (N_26809,N_23353,N_23028);
nand U26810 (N_26810,N_23222,N_23914);
or U26811 (N_26811,N_23778,N_24572);
nand U26812 (N_26812,N_24213,N_22701);
or U26813 (N_26813,N_23944,N_23951);
nand U26814 (N_26814,N_22663,N_23455);
nand U26815 (N_26815,N_23815,N_22941);
nand U26816 (N_26816,N_23050,N_23065);
nor U26817 (N_26817,N_23909,N_24053);
or U26818 (N_26818,N_22785,N_24306);
or U26819 (N_26819,N_23036,N_24124);
or U26820 (N_26820,N_24118,N_24611);
and U26821 (N_26821,N_24321,N_24106);
and U26822 (N_26822,N_22901,N_22597);
or U26823 (N_26823,N_23970,N_24647);
nor U26824 (N_26824,N_23654,N_22735);
and U26825 (N_26825,N_24683,N_22585);
nor U26826 (N_26826,N_24717,N_24096);
or U26827 (N_26827,N_23895,N_24775);
nand U26828 (N_26828,N_24514,N_24884);
xor U26829 (N_26829,N_24848,N_24076);
and U26830 (N_26830,N_23267,N_22662);
xnor U26831 (N_26831,N_22761,N_22884);
nand U26832 (N_26832,N_24786,N_24870);
or U26833 (N_26833,N_24416,N_24285);
nand U26834 (N_26834,N_22834,N_23695);
nand U26835 (N_26835,N_23051,N_23587);
xnor U26836 (N_26836,N_22816,N_22545);
nor U26837 (N_26837,N_22906,N_23854);
xnor U26838 (N_26838,N_23800,N_24988);
nand U26839 (N_26839,N_24411,N_24398);
nor U26840 (N_26840,N_22713,N_24313);
nand U26841 (N_26841,N_24686,N_24736);
or U26842 (N_26842,N_23787,N_23920);
xnor U26843 (N_26843,N_23512,N_23324);
nand U26844 (N_26844,N_23601,N_23806);
nor U26845 (N_26845,N_24413,N_22692);
xnor U26846 (N_26846,N_23521,N_24814);
nand U26847 (N_26847,N_24437,N_23279);
or U26848 (N_26848,N_24585,N_24636);
or U26849 (N_26849,N_24049,N_23408);
or U26850 (N_26850,N_22980,N_24726);
or U26851 (N_26851,N_23372,N_23640);
and U26852 (N_26852,N_24770,N_23635);
and U26853 (N_26853,N_22720,N_24268);
xnor U26854 (N_26854,N_23192,N_23522);
nand U26855 (N_26855,N_24204,N_23071);
xnor U26856 (N_26856,N_23141,N_24101);
and U26857 (N_26857,N_23753,N_22863);
or U26858 (N_26858,N_24906,N_23580);
xnor U26859 (N_26859,N_24535,N_24293);
or U26860 (N_26860,N_23921,N_23722);
nand U26861 (N_26861,N_23800,N_23633);
xor U26862 (N_26862,N_24544,N_24340);
nor U26863 (N_26863,N_22918,N_24187);
and U26864 (N_26864,N_24637,N_23524);
xnor U26865 (N_26865,N_24414,N_24235);
or U26866 (N_26866,N_24502,N_22628);
nand U26867 (N_26867,N_24912,N_24548);
nor U26868 (N_26868,N_23160,N_23295);
or U26869 (N_26869,N_24687,N_24980);
or U26870 (N_26870,N_23610,N_23317);
or U26871 (N_26871,N_23770,N_23526);
nor U26872 (N_26872,N_22555,N_24948);
nand U26873 (N_26873,N_22610,N_24881);
nor U26874 (N_26874,N_24924,N_24950);
xnor U26875 (N_26875,N_23745,N_23085);
nand U26876 (N_26876,N_23698,N_23464);
nor U26877 (N_26877,N_24985,N_23306);
or U26878 (N_26878,N_24755,N_23381);
nand U26879 (N_26879,N_23058,N_24469);
nor U26880 (N_26880,N_22772,N_23607);
nor U26881 (N_26881,N_23976,N_24708);
and U26882 (N_26882,N_24824,N_23027);
xor U26883 (N_26883,N_23775,N_22985);
nand U26884 (N_26884,N_22978,N_23897);
or U26885 (N_26885,N_23429,N_22693);
xnor U26886 (N_26886,N_24433,N_23316);
or U26887 (N_26887,N_23354,N_22605);
nor U26888 (N_26888,N_24658,N_24553);
nor U26889 (N_26889,N_23745,N_23879);
xor U26890 (N_26890,N_24625,N_23510);
nor U26891 (N_26891,N_23705,N_23917);
nand U26892 (N_26892,N_23775,N_23191);
xnor U26893 (N_26893,N_24130,N_24050);
xnor U26894 (N_26894,N_24773,N_22683);
nand U26895 (N_26895,N_24203,N_23048);
nor U26896 (N_26896,N_23429,N_24927);
nor U26897 (N_26897,N_24983,N_23775);
nor U26898 (N_26898,N_22746,N_23526);
nor U26899 (N_26899,N_23731,N_23042);
nor U26900 (N_26900,N_24687,N_24978);
and U26901 (N_26901,N_24755,N_23526);
and U26902 (N_26902,N_24271,N_23431);
or U26903 (N_26903,N_23112,N_22767);
or U26904 (N_26904,N_22617,N_24904);
xnor U26905 (N_26905,N_23829,N_23925);
nand U26906 (N_26906,N_24204,N_23747);
nor U26907 (N_26907,N_24265,N_24315);
or U26908 (N_26908,N_24810,N_23743);
nand U26909 (N_26909,N_24268,N_24500);
or U26910 (N_26910,N_23371,N_24895);
and U26911 (N_26911,N_23918,N_23406);
or U26912 (N_26912,N_24378,N_24301);
xnor U26913 (N_26913,N_24751,N_24750);
nand U26914 (N_26914,N_23318,N_24870);
xnor U26915 (N_26915,N_22737,N_24370);
xor U26916 (N_26916,N_24959,N_23180);
nor U26917 (N_26917,N_24848,N_24267);
and U26918 (N_26918,N_24826,N_24339);
nand U26919 (N_26919,N_22897,N_22591);
or U26920 (N_26920,N_22663,N_22808);
nand U26921 (N_26921,N_24394,N_24634);
nor U26922 (N_26922,N_23819,N_23296);
nor U26923 (N_26923,N_23404,N_24752);
nand U26924 (N_26924,N_23037,N_23220);
nand U26925 (N_26925,N_23981,N_24021);
xnor U26926 (N_26926,N_22881,N_24340);
xnor U26927 (N_26927,N_22936,N_23211);
or U26928 (N_26928,N_22991,N_24257);
and U26929 (N_26929,N_22906,N_23449);
and U26930 (N_26930,N_23792,N_23370);
nand U26931 (N_26931,N_23024,N_24916);
nor U26932 (N_26932,N_24801,N_22585);
or U26933 (N_26933,N_22551,N_24915);
and U26934 (N_26934,N_23795,N_23710);
nor U26935 (N_26935,N_24090,N_23048);
xnor U26936 (N_26936,N_24873,N_23271);
nand U26937 (N_26937,N_24741,N_23830);
nor U26938 (N_26938,N_23354,N_24981);
nand U26939 (N_26939,N_23932,N_23614);
and U26940 (N_26940,N_24839,N_24712);
nand U26941 (N_26941,N_24067,N_24324);
and U26942 (N_26942,N_24776,N_23461);
nor U26943 (N_26943,N_24059,N_24479);
nand U26944 (N_26944,N_23168,N_23312);
xor U26945 (N_26945,N_23387,N_24220);
nor U26946 (N_26946,N_22865,N_24004);
or U26947 (N_26947,N_24969,N_23337);
nand U26948 (N_26948,N_23637,N_23682);
xnor U26949 (N_26949,N_24086,N_23826);
and U26950 (N_26950,N_22842,N_23303);
nand U26951 (N_26951,N_23909,N_23627);
or U26952 (N_26952,N_23986,N_22841);
and U26953 (N_26953,N_24350,N_23205);
and U26954 (N_26954,N_24913,N_22578);
nor U26955 (N_26955,N_24057,N_22850);
xnor U26956 (N_26956,N_23055,N_22974);
nor U26957 (N_26957,N_23995,N_22666);
nand U26958 (N_26958,N_22571,N_23590);
xnor U26959 (N_26959,N_22841,N_23482);
xnor U26960 (N_26960,N_24682,N_23255);
nand U26961 (N_26961,N_23633,N_22788);
nor U26962 (N_26962,N_24544,N_23355);
nor U26963 (N_26963,N_23802,N_24745);
and U26964 (N_26964,N_22815,N_23838);
or U26965 (N_26965,N_23105,N_23758);
and U26966 (N_26966,N_24794,N_24481);
or U26967 (N_26967,N_24378,N_24197);
nand U26968 (N_26968,N_23417,N_22956);
xor U26969 (N_26969,N_22851,N_22703);
nor U26970 (N_26970,N_24643,N_24642);
or U26971 (N_26971,N_23648,N_24026);
and U26972 (N_26972,N_22889,N_24850);
nor U26973 (N_26973,N_24332,N_24175);
or U26974 (N_26974,N_22735,N_24400);
or U26975 (N_26975,N_22803,N_24815);
nor U26976 (N_26976,N_24993,N_23644);
or U26977 (N_26977,N_24399,N_23564);
nand U26978 (N_26978,N_24817,N_24041);
or U26979 (N_26979,N_23357,N_22930);
nor U26980 (N_26980,N_24084,N_23642);
or U26981 (N_26981,N_23493,N_23710);
and U26982 (N_26982,N_24254,N_24243);
nor U26983 (N_26983,N_24961,N_23660);
and U26984 (N_26984,N_22911,N_23730);
nand U26985 (N_26985,N_24545,N_24893);
and U26986 (N_26986,N_24163,N_23803);
and U26987 (N_26987,N_23486,N_23143);
nand U26988 (N_26988,N_23161,N_23477);
xor U26989 (N_26989,N_23040,N_24725);
or U26990 (N_26990,N_23694,N_24386);
nor U26991 (N_26991,N_22606,N_24735);
nand U26992 (N_26992,N_22669,N_23306);
nand U26993 (N_26993,N_23226,N_23625);
nand U26994 (N_26994,N_24824,N_23403);
or U26995 (N_26995,N_24288,N_23635);
nor U26996 (N_26996,N_24537,N_23070);
nand U26997 (N_26997,N_24598,N_24287);
and U26998 (N_26998,N_23221,N_24577);
nor U26999 (N_26999,N_24825,N_23474);
and U27000 (N_27000,N_24059,N_23405);
xnor U27001 (N_27001,N_23485,N_24798);
and U27002 (N_27002,N_23979,N_24477);
or U27003 (N_27003,N_23494,N_22858);
and U27004 (N_27004,N_24856,N_22631);
and U27005 (N_27005,N_22841,N_24726);
nand U27006 (N_27006,N_24044,N_22502);
and U27007 (N_27007,N_24403,N_24514);
nor U27008 (N_27008,N_22974,N_24521);
nor U27009 (N_27009,N_23344,N_23425);
xnor U27010 (N_27010,N_22953,N_24393);
nand U27011 (N_27011,N_24678,N_24931);
nand U27012 (N_27012,N_23662,N_24089);
and U27013 (N_27013,N_22735,N_24927);
or U27014 (N_27014,N_23151,N_24428);
nand U27015 (N_27015,N_23191,N_23460);
nand U27016 (N_27016,N_22737,N_23584);
or U27017 (N_27017,N_23044,N_22529);
xor U27018 (N_27018,N_24569,N_23327);
nand U27019 (N_27019,N_22878,N_24947);
nor U27020 (N_27020,N_22743,N_24082);
nand U27021 (N_27021,N_23335,N_23297);
nor U27022 (N_27022,N_23001,N_23221);
or U27023 (N_27023,N_23900,N_24948);
nand U27024 (N_27024,N_23880,N_24936);
xnor U27025 (N_27025,N_24938,N_22540);
nand U27026 (N_27026,N_22953,N_23270);
nand U27027 (N_27027,N_23839,N_24292);
or U27028 (N_27028,N_23404,N_24628);
and U27029 (N_27029,N_24349,N_22630);
xor U27030 (N_27030,N_24841,N_24707);
nor U27031 (N_27031,N_23300,N_23934);
or U27032 (N_27032,N_24920,N_23220);
nor U27033 (N_27033,N_24841,N_24987);
and U27034 (N_27034,N_23812,N_23890);
xnor U27035 (N_27035,N_23746,N_24658);
nor U27036 (N_27036,N_24394,N_23360);
nor U27037 (N_27037,N_24412,N_23688);
xnor U27038 (N_27038,N_24402,N_24221);
nand U27039 (N_27039,N_23355,N_22917);
xor U27040 (N_27040,N_23023,N_22681);
and U27041 (N_27041,N_24916,N_22643);
nand U27042 (N_27042,N_24448,N_24855);
and U27043 (N_27043,N_22848,N_23946);
or U27044 (N_27044,N_24343,N_23711);
nor U27045 (N_27045,N_22968,N_23340);
nor U27046 (N_27046,N_24050,N_24771);
and U27047 (N_27047,N_24585,N_24827);
nand U27048 (N_27048,N_24637,N_23339);
xnor U27049 (N_27049,N_24821,N_24534);
nor U27050 (N_27050,N_23969,N_23943);
and U27051 (N_27051,N_24049,N_23330);
nand U27052 (N_27052,N_24768,N_23883);
xor U27053 (N_27053,N_23450,N_24249);
and U27054 (N_27054,N_24133,N_23134);
nor U27055 (N_27055,N_24124,N_24290);
or U27056 (N_27056,N_24236,N_23886);
xor U27057 (N_27057,N_24757,N_23205);
xnor U27058 (N_27058,N_23189,N_22570);
nand U27059 (N_27059,N_24560,N_22906);
nor U27060 (N_27060,N_22546,N_22739);
and U27061 (N_27061,N_23933,N_24854);
and U27062 (N_27062,N_22907,N_22991);
nor U27063 (N_27063,N_24043,N_23225);
and U27064 (N_27064,N_22933,N_24111);
or U27065 (N_27065,N_23105,N_24285);
xnor U27066 (N_27066,N_24648,N_24053);
xor U27067 (N_27067,N_23048,N_23332);
nor U27068 (N_27068,N_24730,N_23051);
or U27069 (N_27069,N_23092,N_24527);
and U27070 (N_27070,N_23844,N_24394);
and U27071 (N_27071,N_22505,N_23658);
xnor U27072 (N_27072,N_23985,N_23045);
and U27073 (N_27073,N_24586,N_23338);
nand U27074 (N_27074,N_24275,N_23476);
or U27075 (N_27075,N_22961,N_24302);
xor U27076 (N_27076,N_23667,N_22671);
and U27077 (N_27077,N_24425,N_24900);
or U27078 (N_27078,N_23673,N_23837);
or U27079 (N_27079,N_23932,N_23129);
nor U27080 (N_27080,N_23930,N_23260);
and U27081 (N_27081,N_23027,N_24959);
xor U27082 (N_27082,N_23033,N_23436);
xnor U27083 (N_27083,N_24584,N_24451);
nor U27084 (N_27084,N_23908,N_24072);
xor U27085 (N_27085,N_23097,N_23280);
nand U27086 (N_27086,N_23195,N_23369);
or U27087 (N_27087,N_22538,N_23257);
nor U27088 (N_27088,N_24821,N_22935);
and U27089 (N_27089,N_22911,N_23311);
and U27090 (N_27090,N_24151,N_23663);
or U27091 (N_27091,N_23994,N_24501);
or U27092 (N_27092,N_23654,N_23044);
nand U27093 (N_27093,N_24958,N_22940);
nor U27094 (N_27094,N_23986,N_24116);
nor U27095 (N_27095,N_24166,N_24144);
xor U27096 (N_27096,N_24093,N_23798);
and U27097 (N_27097,N_24837,N_24586);
nand U27098 (N_27098,N_23271,N_24443);
and U27099 (N_27099,N_23035,N_24647);
or U27100 (N_27100,N_23577,N_22834);
nand U27101 (N_27101,N_23348,N_23068);
xor U27102 (N_27102,N_24996,N_24974);
xor U27103 (N_27103,N_23851,N_23029);
or U27104 (N_27104,N_24152,N_22809);
or U27105 (N_27105,N_22875,N_22652);
nor U27106 (N_27106,N_23484,N_24059);
or U27107 (N_27107,N_23857,N_24490);
xnor U27108 (N_27108,N_23654,N_23707);
nor U27109 (N_27109,N_24664,N_24275);
or U27110 (N_27110,N_24571,N_24907);
nand U27111 (N_27111,N_24998,N_23828);
and U27112 (N_27112,N_23871,N_22689);
xor U27113 (N_27113,N_23473,N_22591);
nor U27114 (N_27114,N_22785,N_24075);
and U27115 (N_27115,N_24001,N_22653);
nor U27116 (N_27116,N_22836,N_24348);
and U27117 (N_27117,N_23276,N_22668);
xor U27118 (N_27118,N_23314,N_23153);
or U27119 (N_27119,N_22535,N_24787);
and U27120 (N_27120,N_23064,N_23142);
xor U27121 (N_27121,N_22745,N_22855);
or U27122 (N_27122,N_24431,N_24269);
and U27123 (N_27123,N_24457,N_24287);
and U27124 (N_27124,N_24297,N_24827);
and U27125 (N_27125,N_24854,N_24391);
xor U27126 (N_27126,N_23202,N_23670);
xnor U27127 (N_27127,N_24839,N_22619);
nor U27128 (N_27128,N_22526,N_23919);
nor U27129 (N_27129,N_23073,N_23112);
or U27130 (N_27130,N_22885,N_23030);
nor U27131 (N_27131,N_24227,N_24222);
xnor U27132 (N_27132,N_23800,N_24216);
xor U27133 (N_27133,N_23252,N_22718);
xnor U27134 (N_27134,N_23089,N_23237);
or U27135 (N_27135,N_22583,N_22520);
xor U27136 (N_27136,N_23784,N_23907);
nor U27137 (N_27137,N_24626,N_24942);
xor U27138 (N_27138,N_23383,N_22577);
nor U27139 (N_27139,N_24304,N_22748);
and U27140 (N_27140,N_24182,N_24126);
nand U27141 (N_27141,N_24035,N_23274);
or U27142 (N_27142,N_24619,N_23196);
xnor U27143 (N_27143,N_22871,N_23512);
nand U27144 (N_27144,N_22704,N_24618);
nor U27145 (N_27145,N_23533,N_24513);
xor U27146 (N_27146,N_24501,N_23861);
xnor U27147 (N_27147,N_22983,N_24549);
nand U27148 (N_27148,N_24735,N_23312);
and U27149 (N_27149,N_24048,N_23760);
and U27150 (N_27150,N_23467,N_23129);
nor U27151 (N_27151,N_23926,N_23597);
or U27152 (N_27152,N_23518,N_24255);
and U27153 (N_27153,N_23373,N_22667);
nor U27154 (N_27154,N_23722,N_24198);
nor U27155 (N_27155,N_22652,N_22832);
nor U27156 (N_27156,N_24546,N_23618);
nor U27157 (N_27157,N_23530,N_24034);
nor U27158 (N_27158,N_24087,N_24206);
nor U27159 (N_27159,N_24596,N_23697);
nand U27160 (N_27160,N_22657,N_23724);
xor U27161 (N_27161,N_24634,N_23906);
nand U27162 (N_27162,N_24547,N_23506);
and U27163 (N_27163,N_24186,N_24658);
or U27164 (N_27164,N_23492,N_23926);
xnor U27165 (N_27165,N_24283,N_23140);
and U27166 (N_27166,N_22575,N_22569);
nor U27167 (N_27167,N_22864,N_24613);
or U27168 (N_27168,N_23531,N_22633);
and U27169 (N_27169,N_22733,N_23827);
xor U27170 (N_27170,N_24793,N_24777);
or U27171 (N_27171,N_23931,N_23727);
nand U27172 (N_27172,N_24465,N_22711);
nand U27173 (N_27173,N_22777,N_23563);
nor U27174 (N_27174,N_24458,N_23785);
nor U27175 (N_27175,N_24776,N_24627);
nand U27176 (N_27176,N_22941,N_24599);
xnor U27177 (N_27177,N_22553,N_24504);
xor U27178 (N_27178,N_23241,N_24818);
nor U27179 (N_27179,N_22615,N_24371);
or U27180 (N_27180,N_23751,N_24377);
nor U27181 (N_27181,N_23290,N_22865);
or U27182 (N_27182,N_24439,N_22826);
xnor U27183 (N_27183,N_23372,N_23194);
or U27184 (N_27184,N_22849,N_24848);
nor U27185 (N_27185,N_22559,N_24581);
or U27186 (N_27186,N_23626,N_24442);
or U27187 (N_27187,N_23560,N_23815);
and U27188 (N_27188,N_24198,N_24247);
nor U27189 (N_27189,N_23113,N_24149);
nor U27190 (N_27190,N_23841,N_24589);
and U27191 (N_27191,N_23040,N_24925);
or U27192 (N_27192,N_23640,N_24504);
nor U27193 (N_27193,N_23715,N_23175);
nor U27194 (N_27194,N_24310,N_23909);
and U27195 (N_27195,N_22959,N_24716);
and U27196 (N_27196,N_23879,N_23045);
and U27197 (N_27197,N_22738,N_24724);
nand U27198 (N_27198,N_23889,N_23816);
xor U27199 (N_27199,N_24303,N_23557);
or U27200 (N_27200,N_22823,N_24759);
nand U27201 (N_27201,N_24922,N_22726);
or U27202 (N_27202,N_22739,N_24541);
and U27203 (N_27203,N_22670,N_23537);
nor U27204 (N_27204,N_23085,N_23620);
or U27205 (N_27205,N_24938,N_24656);
nor U27206 (N_27206,N_23188,N_24139);
or U27207 (N_27207,N_23123,N_24459);
and U27208 (N_27208,N_22791,N_23864);
or U27209 (N_27209,N_23678,N_23736);
or U27210 (N_27210,N_23398,N_24140);
nor U27211 (N_27211,N_24082,N_22774);
nor U27212 (N_27212,N_24688,N_24725);
and U27213 (N_27213,N_24098,N_22783);
xor U27214 (N_27214,N_23088,N_24340);
nor U27215 (N_27215,N_23918,N_22861);
nor U27216 (N_27216,N_23950,N_23192);
nor U27217 (N_27217,N_23305,N_23001);
or U27218 (N_27218,N_22595,N_23056);
and U27219 (N_27219,N_23191,N_23236);
nor U27220 (N_27220,N_24963,N_24569);
nor U27221 (N_27221,N_24939,N_22778);
nand U27222 (N_27222,N_23477,N_23737);
xnor U27223 (N_27223,N_22620,N_24189);
nor U27224 (N_27224,N_23920,N_24183);
or U27225 (N_27225,N_22752,N_23856);
nor U27226 (N_27226,N_23044,N_23163);
or U27227 (N_27227,N_22892,N_24087);
or U27228 (N_27228,N_24237,N_23414);
or U27229 (N_27229,N_23117,N_23864);
nand U27230 (N_27230,N_24314,N_23894);
nor U27231 (N_27231,N_24735,N_24481);
nand U27232 (N_27232,N_24745,N_24699);
nand U27233 (N_27233,N_23439,N_22947);
and U27234 (N_27234,N_24118,N_24397);
or U27235 (N_27235,N_22507,N_23324);
xnor U27236 (N_27236,N_22646,N_23317);
nor U27237 (N_27237,N_23050,N_24454);
and U27238 (N_27238,N_23772,N_24855);
xor U27239 (N_27239,N_24106,N_24716);
xnor U27240 (N_27240,N_23337,N_23903);
xnor U27241 (N_27241,N_24577,N_24718);
xor U27242 (N_27242,N_24430,N_23641);
nor U27243 (N_27243,N_23683,N_24040);
or U27244 (N_27244,N_24630,N_23140);
and U27245 (N_27245,N_23650,N_24704);
or U27246 (N_27246,N_23460,N_23956);
xnor U27247 (N_27247,N_24665,N_24860);
nand U27248 (N_27248,N_23118,N_22535);
and U27249 (N_27249,N_24862,N_24784);
xor U27250 (N_27250,N_23549,N_23065);
or U27251 (N_27251,N_23838,N_22553);
xor U27252 (N_27252,N_23400,N_23791);
nand U27253 (N_27253,N_24337,N_23762);
nand U27254 (N_27254,N_22920,N_24740);
xnor U27255 (N_27255,N_24836,N_22694);
nand U27256 (N_27256,N_24025,N_23962);
or U27257 (N_27257,N_23397,N_22516);
and U27258 (N_27258,N_22962,N_22641);
or U27259 (N_27259,N_23505,N_23433);
or U27260 (N_27260,N_24579,N_24042);
nor U27261 (N_27261,N_23505,N_24203);
and U27262 (N_27262,N_24064,N_24243);
or U27263 (N_27263,N_22660,N_23928);
and U27264 (N_27264,N_22917,N_23325);
nor U27265 (N_27265,N_22597,N_23944);
and U27266 (N_27266,N_23195,N_22759);
xor U27267 (N_27267,N_23227,N_22819);
nand U27268 (N_27268,N_22553,N_22544);
or U27269 (N_27269,N_23768,N_22851);
nor U27270 (N_27270,N_24900,N_24228);
xnor U27271 (N_27271,N_24123,N_24278);
xnor U27272 (N_27272,N_23366,N_24129);
nand U27273 (N_27273,N_22508,N_24003);
nand U27274 (N_27274,N_24735,N_24154);
and U27275 (N_27275,N_22846,N_22857);
and U27276 (N_27276,N_22927,N_23191);
xor U27277 (N_27277,N_24248,N_23002);
xor U27278 (N_27278,N_24456,N_23966);
and U27279 (N_27279,N_22517,N_24609);
nand U27280 (N_27280,N_22561,N_24344);
nor U27281 (N_27281,N_24880,N_24607);
nand U27282 (N_27282,N_22971,N_24900);
and U27283 (N_27283,N_24868,N_24809);
nand U27284 (N_27284,N_24541,N_24226);
xnor U27285 (N_27285,N_24791,N_23830);
or U27286 (N_27286,N_22854,N_22790);
xnor U27287 (N_27287,N_23431,N_24478);
and U27288 (N_27288,N_23937,N_22844);
and U27289 (N_27289,N_23322,N_22630);
xnor U27290 (N_27290,N_24083,N_22827);
nor U27291 (N_27291,N_23706,N_22718);
xor U27292 (N_27292,N_24030,N_24007);
nor U27293 (N_27293,N_23166,N_22721);
nor U27294 (N_27294,N_22928,N_23649);
or U27295 (N_27295,N_23092,N_22728);
or U27296 (N_27296,N_22709,N_23368);
nor U27297 (N_27297,N_22530,N_23727);
and U27298 (N_27298,N_24375,N_23842);
or U27299 (N_27299,N_22771,N_23275);
nor U27300 (N_27300,N_24702,N_24220);
xor U27301 (N_27301,N_22813,N_23816);
nor U27302 (N_27302,N_22626,N_23553);
or U27303 (N_27303,N_22745,N_22661);
and U27304 (N_27304,N_23688,N_23903);
nand U27305 (N_27305,N_22878,N_23161);
xnor U27306 (N_27306,N_23205,N_22506);
and U27307 (N_27307,N_23676,N_23366);
nor U27308 (N_27308,N_23529,N_23611);
and U27309 (N_27309,N_23305,N_24458);
nand U27310 (N_27310,N_24413,N_23956);
nor U27311 (N_27311,N_23732,N_24363);
nor U27312 (N_27312,N_23444,N_23378);
xnor U27313 (N_27313,N_24976,N_23890);
or U27314 (N_27314,N_23432,N_22862);
and U27315 (N_27315,N_24738,N_23956);
and U27316 (N_27316,N_24133,N_22570);
or U27317 (N_27317,N_24760,N_23508);
nand U27318 (N_27318,N_24187,N_23875);
or U27319 (N_27319,N_24233,N_23697);
or U27320 (N_27320,N_24724,N_23738);
or U27321 (N_27321,N_22524,N_23328);
or U27322 (N_27322,N_23627,N_24149);
or U27323 (N_27323,N_23635,N_24106);
nand U27324 (N_27324,N_23817,N_24583);
xor U27325 (N_27325,N_22861,N_23110);
and U27326 (N_27326,N_23322,N_23546);
or U27327 (N_27327,N_23824,N_24727);
xnor U27328 (N_27328,N_23217,N_23883);
nor U27329 (N_27329,N_24305,N_22736);
or U27330 (N_27330,N_24636,N_22818);
xor U27331 (N_27331,N_24497,N_23071);
nor U27332 (N_27332,N_23828,N_24880);
or U27333 (N_27333,N_23471,N_22638);
and U27334 (N_27334,N_24383,N_24143);
nor U27335 (N_27335,N_24039,N_24414);
xor U27336 (N_27336,N_24599,N_24424);
and U27337 (N_27337,N_23536,N_22603);
nand U27338 (N_27338,N_24567,N_24547);
nand U27339 (N_27339,N_24635,N_24625);
nor U27340 (N_27340,N_24411,N_23805);
and U27341 (N_27341,N_22728,N_24122);
and U27342 (N_27342,N_22976,N_23837);
or U27343 (N_27343,N_23518,N_22683);
xnor U27344 (N_27344,N_23396,N_24024);
nor U27345 (N_27345,N_23171,N_24725);
and U27346 (N_27346,N_24011,N_22806);
nand U27347 (N_27347,N_24488,N_24286);
or U27348 (N_27348,N_23666,N_22694);
xnor U27349 (N_27349,N_23361,N_23982);
and U27350 (N_27350,N_22812,N_23366);
xnor U27351 (N_27351,N_22699,N_22843);
or U27352 (N_27352,N_22754,N_22853);
nand U27353 (N_27353,N_24462,N_24613);
nor U27354 (N_27354,N_24308,N_22527);
nor U27355 (N_27355,N_22978,N_24432);
xor U27356 (N_27356,N_23428,N_24095);
nor U27357 (N_27357,N_24024,N_24110);
nor U27358 (N_27358,N_24163,N_22941);
nand U27359 (N_27359,N_24820,N_23512);
xor U27360 (N_27360,N_23528,N_24210);
nand U27361 (N_27361,N_24743,N_24599);
nor U27362 (N_27362,N_22612,N_22545);
and U27363 (N_27363,N_23119,N_24476);
xnor U27364 (N_27364,N_22804,N_24598);
xor U27365 (N_27365,N_23411,N_23174);
xnor U27366 (N_27366,N_22682,N_23256);
and U27367 (N_27367,N_23247,N_23642);
nand U27368 (N_27368,N_24387,N_23283);
and U27369 (N_27369,N_23410,N_24185);
nand U27370 (N_27370,N_24124,N_23796);
nand U27371 (N_27371,N_24718,N_23153);
nand U27372 (N_27372,N_24521,N_23853);
nor U27373 (N_27373,N_24309,N_23831);
xor U27374 (N_27374,N_24126,N_24936);
and U27375 (N_27375,N_24075,N_24564);
or U27376 (N_27376,N_24099,N_23497);
or U27377 (N_27377,N_23204,N_23091);
nand U27378 (N_27378,N_23198,N_24071);
xor U27379 (N_27379,N_22634,N_23940);
nand U27380 (N_27380,N_24125,N_24772);
or U27381 (N_27381,N_23722,N_24528);
nor U27382 (N_27382,N_23141,N_24617);
and U27383 (N_27383,N_22790,N_23921);
xnor U27384 (N_27384,N_24997,N_24656);
and U27385 (N_27385,N_24405,N_23426);
nand U27386 (N_27386,N_23508,N_24779);
and U27387 (N_27387,N_22666,N_24766);
nor U27388 (N_27388,N_24938,N_24333);
nand U27389 (N_27389,N_23757,N_24077);
xnor U27390 (N_27390,N_24504,N_24980);
nand U27391 (N_27391,N_24309,N_23978);
and U27392 (N_27392,N_22533,N_24356);
and U27393 (N_27393,N_24747,N_23950);
nand U27394 (N_27394,N_23003,N_23341);
and U27395 (N_27395,N_24392,N_22765);
or U27396 (N_27396,N_24531,N_22669);
nand U27397 (N_27397,N_24400,N_24068);
nand U27398 (N_27398,N_24259,N_24761);
nand U27399 (N_27399,N_23873,N_23722);
nor U27400 (N_27400,N_24207,N_23740);
and U27401 (N_27401,N_24524,N_24963);
or U27402 (N_27402,N_22722,N_24045);
or U27403 (N_27403,N_24519,N_24092);
nand U27404 (N_27404,N_24890,N_22671);
or U27405 (N_27405,N_24530,N_24597);
nand U27406 (N_27406,N_23525,N_23531);
or U27407 (N_27407,N_22976,N_22614);
nand U27408 (N_27408,N_23271,N_24744);
and U27409 (N_27409,N_24866,N_22624);
and U27410 (N_27410,N_24716,N_22927);
and U27411 (N_27411,N_24513,N_23419);
or U27412 (N_27412,N_22652,N_24098);
or U27413 (N_27413,N_23110,N_24177);
and U27414 (N_27414,N_24600,N_24263);
and U27415 (N_27415,N_22722,N_22684);
xor U27416 (N_27416,N_23836,N_22653);
and U27417 (N_27417,N_24696,N_22721);
nor U27418 (N_27418,N_23627,N_24986);
xnor U27419 (N_27419,N_24731,N_24415);
or U27420 (N_27420,N_23490,N_23495);
or U27421 (N_27421,N_23333,N_23498);
and U27422 (N_27422,N_22587,N_23756);
xnor U27423 (N_27423,N_24907,N_23847);
and U27424 (N_27424,N_22997,N_22633);
or U27425 (N_27425,N_24114,N_24837);
nand U27426 (N_27426,N_23031,N_24609);
and U27427 (N_27427,N_23638,N_22985);
and U27428 (N_27428,N_23336,N_23250);
or U27429 (N_27429,N_23294,N_23578);
nand U27430 (N_27430,N_22617,N_24490);
and U27431 (N_27431,N_24272,N_24187);
nand U27432 (N_27432,N_24555,N_22855);
nand U27433 (N_27433,N_24449,N_22807);
or U27434 (N_27434,N_23609,N_23853);
and U27435 (N_27435,N_23607,N_24186);
nand U27436 (N_27436,N_22828,N_23779);
or U27437 (N_27437,N_23384,N_22591);
nand U27438 (N_27438,N_24561,N_22845);
or U27439 (N_27439,N_22785,N_24363);
nor U27440 (N_27440,N_23945,N_24743);
nand U27441 (N_27441,N_22785,N_23795);
or U27442 (N_27442,N_23114,N_22676);
xor U27443 (N_27443,N_22663,N_24325);
or U27444 (N_27444,N_24538,N_24916);
xnor U27445 (N_27445,N_23465,N_23648);
and U27446 (N_27446,N_24337,N_24230);
xor U27447 (N_27447,N_22786,N_24715);
or U27448 (N_27448,N_23411,N_24713);
nor U27449 (N_27449,N_22779,N_24169);
and U27450 (N_27450,N_24958,N_23118);
and U27451 (N_27451,N_23487,N_22562);
nand U27452 (N_27452,N_22933,N_24478);
or U27453 (N_27453,N_23882,N_24005);
xor U27454 (N_27454,N_22849,N_23128);
and U27455 (N_27455,N_22836,N_23211);
nand U27456 (N_27456,N_23246,N_23026);
xor U27457 (N_27457,N_23861,N_24496);
nand U27458 (N_27458,N_22507,N_23564);
nand U27459 (N_27459,N_24333,N_24745);
and U27460 (N_27460,N_24102,N_24374);
nor U27461 (N_27461,N_23841,N_24656);
xnor U27462 (N_27462,N_23213,N_22805);
nand U27463 (N_27463,N_23910,N_23100);
or U27464 (N_27464,N_23276,N_23448);
and U27465 (N_27465,N_23458,N_22920);
and U27466 (N_27466,N_24180,N_22773);
or U27467 (N_27467,N_24310,N_23640);
xnor U27468 (N_27468,N_22713,N_22662);
nor U27469 (N_27469,N_23932,N_24222);
xnor U27470 (N_27470,N_23327,N_23473);
xnor U27471 (N_27471,N_22607,N_22515);
or U27472 (N_27472,N_24406,N_24139);
and U27473 (N_27473,N_24799,N_24318);
xnor U27474 (N_27474,N_23098,N_22872);
or U27475 (N_27475,N_23589,N_24744);
nand U27476 (N_27476,N_22885,N_23792);
xor U27477 (N_27477,N_23033,N_22910);
nor U27478 (N_27478,N_22633,N_22817);
nand U27479 (N_27479,N_23747,N_23831);
xor U27480 (N_27480,N_22852,N_23970);
or U27481 (N_27481,N_23192,N_23301);
or U27482 (N_27482,N_24045,N_23267);
and U27483 (N_27483,N_24920,N_24571);
nor U27484 (N_27484,N_24553,N_24247);
nor U27485 (N_27485,N_24833,N_23056);
and U27486 (N_27486,N_22701,N_23250);
xnor U27487 (N_27487,N_24535,N_23545);
nor U27488 (N_27488,N_22508,N_24014);
or U27489 (N_27489,N_23677,N_22832);
or U27490 (N_27490,N_22541,N_24748);
nor U27491 (N_27491,N_23929,N_24849);
and U27492 (N_27492,N_24124,N_23657);
and U27493 (N_27493,N_24126,N_23434);
nand U27494 (N_27494,N_23051,N_23327);
xnor U27495 (N_27495,N_22858,N_24745);
xor U27496 (N_27496,N_23681,N_23323);
or U27497 (N_27497,N_22674,N_24841);
and U27498 (N_27498,N_22700,N_23591);
nand U27499 (N_27499,N_24246,N_22595);
and U27500 (N_27500,N_26442,N_26226);
xor U27501 (N_27501,N_27256,N_25397);
xor U27502 (N_27502,N_25608,N_25075);
xnor U27503 (N_27503,N_25305,N_25371);
or U27504 (N_27504,N_26394,N_25805);
and U27505 (N_27505,N_27282,N_27244);
nor U27506 (N_27506,N_25641,N_27238);
or U27507 (N_27507,N_27200,N_25786);
xnor U27508 (N_27508,N_25538,N_25960);
nand U27509 (N_27509,N_27320,N_25071);
xnor U27510 (N_27510,N_25540,N_26834);
nand U27511 (N_27511,N_26152,N_25217);
nand U27512 (N_27512,N_26204,N_25949);
nor U27513 (N_27513,N_25324,N_26883);
xor U27514 (N_27514,N_26037,N_27471);
nand U27515 (N_27515,N_27129,N_26523);
nand U27516 (N_27516,N_26386,N_25828);
xor U27517 (N_27517,N_27472,N_26746);
nand U27518 (N_27518,N_26137,N_26635);
nor U27519 (N_27519,N_25160,N_26965);
nand U27520 (N_27520,N_26822,N_26168);
xor U27521 (N_27521,N_25045,N_25588);
xor U27522 (N_27522,N_27105,N_26871);
nor U27523 (N_27523,N_25335,N_25103);
and U27524 (N_27524,N_26842,N_26653);
xnor U27525 (N_27525,N_27036,N_26351);
or U27526 (N_27526,N_27075,N_27057);
nand U27527 (N_27527,N_27398,N_26547);
nor U27528 (N_27528,N_25696,N_27035);
nor U27529 (N_27529,N_25237,N_25395);
nor U27530 (N_27530,N_27215,N_25593);
xor U27531 (N_27531,N_27302,N_26165);
or U27532 (N_27532,N_26967,N_26030);
nand U27533 (N_27533,N_25746,N_25547);
and U27534 (N_27534,N_26040,N_25282);
xnor U27535 (N_27535,N_26280,N_27182);
xor U27536 (N_27536,N_25627,N_26320);
and U27537 (N_27537,N_27315,N_27007);
or U27538 (N_27538,N_27268,N_25799);
or U27539 (N_27539,N_25824,N_25754);
and U27540 (N_27540,N_26140,N_26566);
or U27541 (N_27541,N_26277,N_25060);
nand U27542 (N_27542,N_27100,N_26141);
and U27543 (N_27543,N_26964,N_25874);
xor U27544 (N_27544,N_26858,N_26004);
xor U27545 (N_27545,N_27204,N_26303);
nand U27546 (N_27546,N_26682,N_26129);
xor U27547 (N_27547,N_25202,N_25107);
nor U27548 (N_27548,N_25231,N_26672);
nand U27549 (N_27549,N_27206,N_26745);
nor U27550 (N_27550,N_27491,N_27401);
and U27551 (N_27551,N_26528,N_27116);
and U27552 (N_27552,N_26544,N_26323);
xnor U27553 (N_27553,N_25076,N_25437);
or U27554 (N_27554,N_25480,N_27396);
or U27555 (N_27555,N_26762,N_25000);
nor U27556 (N_27556,N_26316,N_25808);
nand U27557 (N_27557,N_27189,N_26982);
or U27558 (N_27558,N_26231,N_26574);
xor U27559 (N_27559,N_26287,N_26027);
nor U27560 (N_27560,N_26909,N_25609);
or U27561 (N_27561,N_26872,N_25708);
or U27562 (N_27562,N_26483,N_27203);
or U27563 (N_27563,N_26530,N_26186);
nand U27564 (N_27564,N_25127,N_26409);
nand U27565 (N_27565,N_26616,N_25881);
nand U27566 (N_27566,N_26191,N_27261);
xor U27567 (N_27567,N_25298,N_25380);
nor U27568 (N_27568,N_25266,N_27480);
nor U27569 (N_27569,N_26591,N_26996);
and U27570 (N_27570,N_26773,N_25510);
nor U27571 (N_27571,N_25080,N_25674);
or U27572 (N_27572,N_26061,N_26601);
nor U27573 (N_27573,N_26881,N_26758);
xor U27574 (N_27574,N_27356,N_26487);
or U27575 (N_27575,N_25650,N_27037);
xor U27576 (N_27576,N_26042,N_26243);
and U27577 (N_27577,N_25645,N_27106);
nand U27578 (N_27578,N_26580,N_26377);
and U27579 (N_27579,N_27321,N_25018);
nor U27580 (N_27580,N_27458,N_25253);
nor U27581 (N_27581,N_27193,N_26337);
xnor U27582 (N_27582,N_25557,N_25230);
nor U27583 (N_27583,N_26602,N_27280);
nand U27584 (N_27584,N_27058,N_25325);
or U27585 (N_27585,N_25252,N_25839);
or U27586 (N_27586,N_26922,N_26609);
and U27587 (N_27587,N_27045,N_26265);
nand U27588 (N_27588,N_25104,N_26458);
and U27589 (N_27589,N_25381,N_25337);
and U27590 (N_27590,N_27466,N_25320);
and U27591 (N_27591,N_26146,N_25710);
nor U27592 (N_27592,N_27051,N_25878);
or U27593 (N_27593,N_26012,N_25239);
nor U27594 (N_27594,N_26148,N_25830);
and U27595 (N_27595,N_26234,N_25921);
xor U27596 (N_27596,N_26671,N_27409);
and U27597 (N_27597,N_26080,N_25474);
nor U27598 (N_27598,N_26262,N_27242);
nor U27599 (N_27599,N_25341,N_26485);
and U27600 (N_27600,N_25917,N_27085);
nor U27601 (N_27601,N_27436,N_25625);
or U27602 (N_27602,N_26005,N_25091);
and U27603 (N_27603,N_25677,N_27194);
xor U27604 (N_27604,N_26576,N_25940);
or U27605 (N_27605,N_26403,N_27416);
xnor U27606 (N_27606,N_26070,N_25442);
xor U27607 (N_27607,N_26166,N_25098);
nor U27608 (N_27608,N_26361,N_27446);
nor U27609 (N_27609,N_25670,N_27265);
nor U27610 (N_27610,N_26217,N_26880);
nand U27611 (N_27611,N_26763,N_26138);
xor U27612 (N_27612,N_25583,N_26687);
nor U27613 (N_27613,N_27197,N_26479);
nor U27614 (N_27614,N_25351,N_27190);
nor U27615 (N_27615,N_26803,N_26807);
nor U27616 (N_27616,N_27053,N_26368);
or U27617 (N_27617,N_26087,N_26689);
nor U27618 (N_27618,N_25276,N_26235);
nand U27619 (N_27619,N_26205,N_25365);
nand U27620 (N_27620,N_26966,N_26662);
and U27621 (N_27621,N_26674,N_25847);
nand U27622 (N_27622,N_27047,N_26617);
xnor U27623 (N_27623,N_27434,N_27428);
and U27624 (N_27624,N_26536,N_25511);
xor U27625 (N_27625,N_26753,N_26282);
or U27626 (N_27626,N_25033,N_26976);
nor U27627 (N_27627,N_25880,N_25742);
and U27628 (N_27628,N_26144,N_26113);
nor U27629 (N_27629,N_25475,N_26865);
nand U27630 (N_27630,N_25129,N_26371);
or U27631 (N_27631,N_26471,N_27325);
nand U27632 (N_27632,N_25218,N_27167);
and U27633 (N_27633,N_26607,N_25775);
or U27634 (N_27634,N_25321,N_26153);
or U27635 (N_27635,N_26133,N_27447);
nor U27636 (N_27636,N_26009,N_27181);
or U27637 (N_27637,N_27288,N_25621);
and U27638 (N_27638,N_25532,N_25013);
nand U27639 (N_27639,N_26990,N_27452);
and U27640 (N_27640,N_25610,N_26218);
xnor U27641 (N_27641,N_26278,N_27032);
and U27642 (N_27642,N_26295,N_25911);
or U27643 (N_27643,N_25637,N_25812);
or U27644 (N_27644,N_26346,N_26119);
nand U27645 (N_27645,N_25017,N_27122);
xnor U27646 (N_27646,N_26221,N_25162);
or U27647 (N_27647,N_27298,N_26721);
xnor U27648 (N_27648,N_25001,N_26508);
and U27649 (N_27649,N_27294,N_27324);
nor U27650 (N_27650,N_27459,N_27077);
nand U27651 (N_27651,N_26577,N_25778);
nand U27652 (N_27652,N_27208,N_26389);
xor U27653 (N_27653,N_26756,N_27161);
nand U27654 (N_27654,N_26761,N_25420);
and U27655 (N_27655,N_26385,N_25560);
nor U27656 (N_27656,N_25906,N_26885);
nand U27657 (N_27657,N_26860,N_26311);
nand U27658 (N_27658,N_25310,N_26811);
xnor U27659 (N_27659,N_27140,N_27198);
xor U27660 (N_27660,N_25372,N_25472);
or U27661 (N_27661,N_26586,N_26684);
xor U27662 (N_27662,N_27254,N_26501);
nand U27663 (N_27663,N_27043,N_25408);
xor U27664 (N_27664,N_25722,N_27087);
or U27665 (N_27665,N_25977,N_27152);
xor U27666 (N_27666,N_26043,N_27367);
xnor U27667 (N_27667,N_26683,N_26703);
xnor U27668 (N_27668,N_25173,N_26456);
and U27669 (N_27669,N_26810,N_26380);
xor U27670 (N_27670,N_27166,N_25081);
nor U27671 (N_27671,N_25758,N_26018);
nor U27672 (N_27672,N_26582,N_26540);
xor U27673 (N_27673,N_26961,N_25980);
or U27674 (N_27674,N_25415,N_25692);
nor U27675 (N_27675,N_26420,N_25592);
xor U27676 (N_27676,N_26161,N_25125);
and U27677 (N_27677,N_27253,N_27155);
or U27678 (N_27678,N_25431,N_26825);
xnor U27679 (N_27679,N_26852,N_26719);
or U27680 (N_27680,N_25015,N_26959);
and U27681 (N_27681,N_25750,N_26354);
nor U27682 (N_27682,N_27091,N_25897);
xnor U27683 (N_27683,N_26275,N_27052);
nor U27684 (N_27684,N_26804,N_26621);
nand U27685 (N_27685,N_26686,N_25434);
nand U27686 (N_27686,N_26291,N_27080);
and U27687 (N_27687,N_27448,N_27498);
nand U27688 (N_27688,N_25130,N_25678);
nor U27689 (N_27689,N_27031,N_25100);
xnor U27690 (N_27690,N_26294,N_26759);
and U27691 (N_27691,N_25082,N_27148);
or U27692 (N_27692,N_27259,N_26192);
nor U27693 (N_27693,N_27171,N_25279);
nand U27694 (N_27694,N_26725,N_25261);
nand U27695 (N_27695,N_25003,N_27277);
xnor U27696 (N_27696,N_26707,N_26980);
nand U27697 (N_27697,N_27114,N_26222);
or U27698 (N_27698,N_25248,N_27250);
nand U27699 (N_27699,N_25049,N_25546);
nor U27700 (N_27700,N_25355,N_26279);
or U27701 (N_27701,N_26023,N_25025);
or U27702 (N_27702,N_25823,N_26359);
and U27703 (N_27703,N_26417,N_26747);
nor U27704 (N_27704,N_25155,N_25986);
or U27705 (N_27705,N_27432,N_25293);
nand U27706 (N_27706,N_25660,N_26962);
or U27707 (N_27707,N_26655,N_26488);
xnor U27708 (N_27708,N_25953,N_25760);
or U27709 (N_27709,N_25469,N_26421);
and U27710 (N_27710,N_26636,N_25443);
or U27711 (N_27711,N_25726,N_26125);
or U27712 (N_27712,N_26679,N_27453);
nand U27713 (N_27713,N_26335,N_26283);
nand U27714 (N_27714,N_27378,N_27439);
nand U27715 (N_27715,N_26912,N_25174);
nor U27716 (N_27716,N_26644,N_25647);
nand U27717 (N_27717,N_26246,N_25707);
nand U27718 (N_27718,N_25181,N_26928);
xnor U27719 (N_27719,N_26227,N_26948);
xnor U27720 (N_27720,N_27297,N_27327);
nor U27721 (N_27721,N_27243,N_27186);
and U27722 (N_27722,N_26363,N_26604);
or U27723 (N_27723,N_25142,N_27231);
nand U27724 (N_27724,N_25446,N_27317);
or U27725 (N_27725,N_27038,N_25969);
xor U27726 (N_27726,N_27490,N_25619);
and U27727 (N_27727,N_25387,N_25074);
nand U27728 (N_27728,N_25785,N_25236);
nand U27729 (N_27729,N_25496,N_25576);
or U27730 (N_27730,N_25894,N_27121);
or U27731 (N_27731,N_26696,N_26787);
nand U27732 (N_27732,N_25028,N_25551);
nand U27733 (N_27733,N_27082,N_25456);
and U27734 (N_27734,N_25109,N_27060);
and U27735 (N_27735,N_25587,N_25809);
and U27736 (N_27736,N_25640,N_26194);
nand U27737 (N_27737,N_26358,N_27408);
nand U27738 (N_27738,N_25507,N_26727);
and U27739 (N_27739,N_26779,N_26252);
xnor U27740 (N_27740,N_26668,N_25085);
and U27741 (N_27741,N_26520,N_25055);
nand U27742 (N_27742,N_25864,N_26370);
nand U27743 (N_27743,N_26986,N_25283);
and U27744 (N_27744,N_26466,N_26190);
or U27745 (N_27745,N_26270,N_26890);
and U27746 (N_27746,N_25762,N_25791);
nor U27747 (N_27747,N_26338,N_27272);
and U27748 (N_27748,N_25994,N_27101);
xnor U27749 (N_27749,N_25304,N_25334);
nand U27750 (N_27750,N_25251,N_25704);
xor U27751 (N_27751,N_26984,N_25756);
xnor U27752 (N_27752,N_26706,N_26008);
and U27753 (N_27753,N_25187,N_25468);
and U27754 (N_27754,N_26264,N_26647);
or U27755 (N_27755,N_26569,N_25976);
nor U27756 (N_27756,N_25077,N_25342);
or U27757 (N_27757,N_26006,N_25838);
and U27758 (N_27758,N_26101,N_26063);
nand U27759 (N_27759,N_26808,N_26648);
or U27760 (N_27760,N_25141,N_25548);
nand U27761 (N_27761,N_26209,N_25935);
and U27762 (N_27762,N_25851,N_26053);
or U27763 (N_27763,N_26500,N_26341);
nor U27764 (N_27764,N_27341,N_26603);
and U27765 (N_27765,N_26940,N_25852);
or U27766 (N_27766,N_25582,N_27074);
nand U27767 (N_27767,N_25300,N_25689);
xnor U27768 (N_27768,N_25748,N_25117);
xor U27769 (N_27769,N_25326,N_27102);
or U27770 (N_27770,N_25634,N_25822);
and U27771 (N_27771,N_26641,N_25745);
and U27772 (N_27772,N_26065,N_25781);
and U27773 (N_27773,N_27178,N_25233);
nor U27774 (N_27774,N_27454,N_27390);
xnor U27775 (N_27775,N_25752,N_25247);
xnor U27776 (N_27776,N_27316,N_25598);
nand U27777 (N_27777,N_27111,N_25163);
nor U27778 (N_27778,N_25414,N_26178);
nand U27779 (N_27779,N_27456,N_26935);
or U27780 (N_27780,N_26093,N_26669);
and U27781 (N_27781,N_25491,N_25256);
nor U27782 (N_27782,N_25140,N_27266);
nor U27783 (N_27783,N_25811,N_27263);
nor U27784 (N_27784,N_25223,N_25899);
and U27785 (N_27785,N_25875,N_26304);
nor U27786 (N_27786,N_25292,N_25856);
and U27787 (N_27787,N_26273,N_26260);
nand U27788 (N_27788,N_25157,N_26952);
xor U27789 (N_27789,N_26039,N_26728);
and U27790 (N_27790,N_27041,N_26765);
or U27791 (N_27791,N_25702,N_25370);
xnor U27792 (N_27792,N_27219,N_26364);
xnor U27793 (N_27793,N_25034,N_25144);
or U27794 (N_27794,N_26493,N_25108);
nand U27795 (N_27795,N_25889,N_27025);
nand U27796 (N_27796,N_26742,N_27068);
and U27797 (N_27797,N_25086,N_27461);
xnor U27798 (N_27798,N_25620,N_25193);
nor U27799 (N_27799,N_25730,N_25542);
xnor U27800 (N_27800,N_26318,N_26159);
nor U27801 (N_27801,N_26637,N_26357);
or U27802 (N_27802,N_26086,N_26664);
xnor U27803 (N_27803,N_26916,N_25923);
nand U27804 (N_27804,N_26438,N_26846);
and U27805 (N_27805,N_26289,N_25361);
or U27806 (N_27806,N_27300,N_26778);
nand U27807 (N_27807,N_25254,N_25078);
and U27808 (N_27808,N_26542,N_25888);
nor U27809 (N_27809,N_25749,N_26734);
nand U27810 (N_27810,N_25030,N_26660);
nor U27811 (N_27811,N_25596,N_26347);
nor U27812 (N_27812,N_27094,N_26333);
nand U27813 (N_27813,N_25366,N_27365);
and U27814 (N_27814,N_27017,N_25501);
xnor U27815 (N_27815,N_25925,N_26945);
and U27816 (N_27816,N_25633,N_25736);
nor U27817 (N_27817,N_26381,N_25920);
nand U27818 (N_27818,N_27175,N_25201);
and U27819 (N_27819,N_26533,N_25432);
nor U27820 (N_27820,N_26897,N_25398);
nand U27821 (N_27821,N_27162,N_25166);
and U27822 (N_27822,N_26010,N_25769);
or U27823 (N_27823,N_25763,N_26077);
or U27824 (N_27824,N_26415,N_25840);
nor U27825 (N_27825,N_25413,N_27176);
or U27826 (N_27826,N_25336,N_27495);
nand U27827 (N_27827,N_25330,N_26785);
xor U27828 (N_27828,N_25221,N_25084);
nor U27829 (N_27829,N_25079,N_25800);
and U27830 (N_27830,N_26892,N_25394);
and U27831 (N_27831,N_25250,N_26312);
xnor U27832 (N_27832,N_25473,N_25814);
xor U27833 (N_27833,N_26470,N_25612);
and U27834 (N_27834,N_26794,N_26550);
xnor U27835 (N_27835,N_25558,N_26896);
nand U27836 (N_27836,N_25198,N_26649);
and U27837 (N_27837,N_26901,N_25908);
nand U27838 (N_27838,N_25712,N_27361);
nor U27839 (N_27839,N_25418,N_26177);
or U27840 (N_27840,N_25784,N_26048);
and U27841 (N_27841,N_26579,N_26407);
xor U27842 (N_27842,N_25553,N_25407);
xor U27843 (N_27843,N_25919,N_25455);
or U27844 (N_27844,N_25416,N_25611);
nor U27845 (N_27845,N_25913,N_26482);
and U27846 (N_27846,N_25618,N_26766);
nor U27847 (N_27847,N_25943,N_27240);
or U27848 (N_27848,N_26934,N_25701);
or U27849 (N_27849,N_26981,N_27230);
nand U27850 (N_27850,N_25570,N_27120);
xor U27851 (N_27851,N_25178,N_26799);
xor U27852 (N_27852,N_25516,N_25624);
or U27853 (N_27853,N_25389,N_25541);
nor U27854 (N_27854,N_27147,N_27020);
nor U27855 (N_27855,N_25268,N_27286);
and U27856 (N_27856,N_25119,N_27233);
nand U27857 (N_27857,N_25843,N_25374);
nor U27858 (N_27858,N_26749,N_26401);
xor U27859 (N_27859,N_26849,N_26911);
nand U27860 (N_27860,N_25832,N_25514);
nor U27861 (N_27861,N_25787,N_26240);
and U27862 (N_27862,N_25347,N_25697);
xor U27863 (N_27863,N_25961,N_27287);
and U27864 (N_27864,N_25631,N_27044);
nor U27865 (N_27865,N_26998,N_26317);
nand U27866 (N_27866,N_26864,N_26397);
or U27867 (N_27867,N_25483,N_25687);
nor U27868 (N_27868,N_27137,N_26132);
or U27869 (N_27869,N_25410,N_25821);
nand U27870 (N_27870,N_26848,N_27146);
nand U27871 (N_27871,N_26828,N_25275);
or U27872 (N_27872,N_26238,N_26941);
or U27873 (N_27873,N_26134,N_25605);
and U27874 (N_27874,N_26772,N_25213);
nand U27875 (N_27875,N_26947,N_27118);
nor U27876 (N_27876,N_26507,N_26248);
and U27877 (N_27877,N_25484,N_27196);
and U27878 (N_27878,N_26836,N_27353);
and U27879 (N_27879,N_27403,N_25694);
xor U27880 (N_27880,N_25007,N_26541);
xor U27881 (N_27881,N_25520,N_27063);
xnor U27882 (N_27882,N_27030,N_26534);
or U27883 (N_27883,N_25519,N_27220);
nor U27884 (N_27884,N_26791,N_26047);
nor U27885 (N_27885,N_25972,N_25740);
xnor U27886 (N_27886,N_27050,N_25345);
or U27887 (N_27887,N_26244,N_25022);
and U27888 (N_27888,N_25837,N_25693);
or U27889 (N_27889,N_27108,N_26960);
and U27890 (N_27890,N_26328,N_25797);
nand U27891 (N_27891,N_27226,N_26418);
and U27892 (N_27892,N_27083,N_25617);
or U27893 (N_27893,N_25757,N_25448);
or U27894 (N_27894,N_26054,N_26627);
nor U27895 (N_27895,N_25792,N_25167);
or U27896 (N_27896,N_25360,N_26233);
xnor U27897 (N_27897,N_25657,N_25695);
nand U27898 (N_27898,N_25984,N_26147);
and U27899 (N_27899,N_26123,N_25973);
and U27900 (N_27900,N_27389,N_25177);
or U27901 (N_27901,N_27229,N_26379);
nand U27902 (N_27902,N_26863,N_26526);
or U27903 (N_27903,N_26963,N_25877);
nand U27904 (N_27904,N_26437,N_25280);
nand U27905 (N_27905,N_26505,N_25403);
or U27906 (N_27906,N_27089,N_26565);
nand U27907 (N_27907,N_25220,N_26886);
or U27908 (N_27908,N_26882,N_25998);
nand U27909 (N_27909,N_26531,N_26075);
nand U27910 (N_27910,N_25948,N_26771);
xnor U27911 (N_27911,N_27323,N_27497);
or U27912 (N_27912,N_26176,N_25132);
nand U27913 (N_27913,N_27257,N_25296);
and U27914 (N_27914,N_25635,N_26658);
xor U27915 (N_27915,N_26297,N_26904);
nor U27916 (N_27916,N_27392,N_26549);
xnor U27917 (N_27917,N_26416,N_27333);
or U27918 (N_27918,N_25136,N_27252);
nor U27919 (N_27919,N_25688,N_25751);
nor U27920 (N_27920,N_26411,N_25421);
and U27921 (N_27921,N_26600,N_25259);
or U27922 (N_27922,N_25008,N_25767);
or U27923 (N_27923,N_25146,N_26143);
or U27924 (N_27924,N_26163,N_27465);
nand U27925 (N_27925,N_26921,N_25666);
and U27926 (N_27926,N_25776,N_26453);
nor U27927 (N_27927,N_26028,N_26900);
xor U27928 (N_27928,N_25463,N_26097);
or U27929 (N_27929,N_25574,N_25842);
and U27930 (N_27930,N_26106,N_25430);
xnor U27931 (N_27931,N_27125,N_25244);
nand U27932 (N_27932,N_25409,N_25158);
and U27933 (N_27933,N_27345,N_26268);
and U27934 (N_27934,N_25467,N_26592);
nand U27935 (N_27935,N_27142,N_26782);
nor U27936 (N_27936,N_27014,N_25440);
or U27937 (N_27937,N_27098,N_26019);
nor U27938 (N_27938,N_27010,N_25428);
nand U27939 (N_27939,N_25552,N_26983);
or U27940 (N_27940,N_25376,N_25928);
and U27941 (N_27941,N_26013,N_25048);
nor U27942 (N_27942,N_25105,N_25535);
xor U27943 (N_27943,N_26350,N_25445);
or U27944 (N_27944,N_25951,N_26216);
and U27945 (N_27945,N_25329,N_27064);
and U27946 (N_27946,N_26472,N_25589);
nand U27947 (N_27947,N_27475,N_26556);
and U27948 (N_27948,N_26735,N_25094);
or U27949 (N_27949,N_26700,N_27411);
nand U27950 (N_27950,N_25934,N_25278);
nand U27951 (N_27951,N_25490,N_27133);
xnor U27952 (N_27952,N_26029,N_25183);
or U27953 (N_27953,N_26740,N_26340);
nor U27954 (N_27954,N_25012,N_26623);
nand U27955 (N_27955,N_26924,N_25281);
nand U27956 (N_27956,N_27394,N_26625);
nand U27957 (N_27957,N_25870,N_26838);
nand U27958 (N_27958,N_25664,N_26851);
and U27959 (N_27959,N_26694,N_27296);
and U27960 (N_27960,N_25717,N_26365);
xnor U27961 (N_27961,N_26189,N_26902);
or U27962 (N_27962,N_25713,N_25853);
and U27963 (N_27963,N_26820,N_25826);
or U27964 (N_27964,N_26926,N_26732);
or U27965 (N_27965,N_26412,N_26382);
nand U27966 (N_27966,N_27097,N_26561);
nand U27967 (N_27967,N_26840,N_26770);
or U27968 (N_27968,N_26914,N_25313);
and U27969 (N_27969,N_26305,N_25289);
and U27970 (N_27970,N_26906,N_27160);
xor U27971 (N_27971,N_26847,N_26789);
nor U27972 (N_27972,N_26572,N_27026);
and U27973 (N_27973,N_25195,N_25063);
and U27974 (N_27974,N_26459,N_25989);
nand U27975 (N_27975,N_25367,N_25106);
nor U27976 (N_27976,N_26539,N_26717);
and U27977 (N_27977,N_25720,N_26888);
and U27978 (N_27978,N_25854,N_26041);
nor U27979 (N_27979,N_25056,N_25126);
xor U27980 (N_27980,N_25404,N_27217);
nor U27981 (N_27981,N_26513,N_25914);
nor U27982 (N_27982,N_25690,N_25773);
nor U27983 (N_27983,N_27444,N_27228);
nor U27984 (N_27984,N_25993,N_25987);
and U27985 (N_27985,N_26588,N_25069);
nand U27986 (N_27986,N_27164,N_26263);
or U27987 (N_27987,N_26130,N_26519);
and U27988 (N_27988,N_26236,N_27374);
and U27989 (N_27989,N_27467,N_27366);
or U27990 (N_27990,N_25663,N_25046);
nand U27991 (N_27991,N_26868,N_26843);
or U27992 (N_27992,N_25947,N_26590);
nand U27993 (N_27993,N_26136,N_26818);
and U27994 (N_27994,N_26552,N_25176);
nor U27995 (N_27995,N_25902,N_25892);
and U27996 (N_27996,N_25302,N_25867);
nor U27997 (N_27997,N_25863,N_26336);
xnor U27998 (N_27998,N_25721,N_27419);
or U27999 (N_27999,N_26419,N_25171);
nor U28000 (N_28000,N_26056,N_26331);
xor U28001 (N_28001,N_27372,N_25186);
xor U28002 (N_28002,N_25580,N_25658);
nand U28003 (N_28003,N_26214,N_26105);
and U28004 (N_28004,N_26334,N_26068);
or U28005 (N_28005,N_25924,N_25898);
nor U28006 (N_28006,N_27309,N_26809);
and U28007 (N_28007,N_25343,N_27004);
nand U28008 (N_28008,N_26111,N_25453);
nor U28009 (N_28009,N_26388,N_26284);
or U28010 (N_28010,N_27469,N_27195);
nor U28011 (N_28011,N_26593,N_25331);
and U28012 (N_28012,N_25727,N_26757);
and U28013 (N_28013,N_25489,N_26833);
and U28014 (N_28014,N_25032,N_25447);
xor U28015 (N_28015,N_25561,N_26856);
xor U28016 (N_28016,N_26455,N_27090);
nor U28017 (N_28017,N_27391,N_26713);
or U28018 (N_28018,N_26116,N_26139);
nor U28019 (N_28019,N_27199,N_26271);
or U28020 (N_28020,N_27470,N_25096);
xor U28021 (N_28021,N_26400,N_25211);
nor U28022 (N_28022,N_25955,N_26790);
nor U28023 (N_28023,N_26760,N_26180);
nand U28024 (N_28024,N_26399,N_26308);
and U28025 (N_28025,N_26575,N_27313);
nand U28026 (N_28026,N_25765,N_27003);
or U28027 (N_28027,N_27338,N_25788);
or U28028 (N_28028,N_27241,N_26510);
nand U28029 (N_28029,N_27437,N_26614);
xor U28030 (N_28030,N_27273,N_25087);
or U28031 (N_28031,N_27154,N_25209);
xnor U28032 (N_28032,N_25643,N_26731);
or U28033 (N_28033,N_25073,N_27222);
xnor U28034 (N_28034,N_26730,N_26560);
nand U28035 (N_28035,N_26884,N_26237);
nor U28036 (N_28036,N_26210,N_25499);
nand U28037 (N_28037,N_26454,N_26801);
or U28038 (N_28038,N_26930,N_26187);
or U28039 (N_28039,N_26184,N_26690);
xnor U28040 (N_28040,N_25779,N_27258);
and U28041 (N_28041,N_27019,N_25041);
xnor U28042 (N_28042,N_27248,N_26973);
or U28043 (N_28043,N_25139,N_26769);
and U28044 (N_28044,N_25191,N_26465);
xnor U28045 (N_28045,N_27283,N_25005);
nor U28046 (N_28046,N_26557,N_27385);
nand U28047 (N_28047,N_25378,N_25422);
nand U28048 (N_28048,N_27328,N_27429);
xor U28049 (N_28049,N_26494,N_26876);
and U28050 (N_28050,N_27386,N_26942);
nor U28051 (N_28051,N_25185,N_26293);
nor U28052 (N_28052,N_25556,N_25306);
or U28053 (N_28053,N_26639,N_27292);
and U28054 (N_28054,N_26819,N_26285);
or U28055 (N_28055,N_26518,N_27499);
nor U28056 (N_28056,N_27221,N_27039);
xnor U28057 (N_28057,N_25855,N_25044);
and U28058 (N_28058,N_27468,N_26319);
or U28059 (N_28059,N_26788,N_27293);
nand U28060 (N_28060,N_26943,N_26845);
or U28061 (N_28061,N_25124,N_26188);
nand U28062 (N_28062,N_26172,N_27234);
or U28063 (N_28063,N_25794,N_26448);
or U28064 (N_28064,N_26985,N_26780);
nand U28065 (N_28065,N_25850,N_25246);
or U28066 (N_28066,N_25452,N_26720);
and U28067 (N_28067,N_25500,N_26154);
or U28068 (N_28068,N_27086,N_26229);
nor U28069 (N_28069,N_26768,N_25255);
or U28070 (N_28070,N_26201,N_26444);
and U28071 (N_28071,N_26302,N_27346);
or U28072 (N_28072,N_26670,N_26392);
and U28073 (N_28073,N_25734,N_26480);
nand U28074 (N_28074,N_25804,N_25053);
nand U28075 (N_28075,N_25390,N_25819);
and U28076 (N_28076,N_25010,N_27081);
and U28077 (N_28077,N_25212,N_27119);
or U28078 (N_28078,N_25723,N_25057);
xor U28079 (N_28079,N_26256,N_26537);
and U28080 (N_28080,N_26290,N_25882);
xor U28081 (N_28081,N_27332,N_25893);
nand U28082 (N_28082,N_26391,N_26821);
nor U28083 (N_28083,N_25135,N_25009);
nand U28084 (N_28084,N_25918,N_26230);
nand U28085 (N_28085,N_25790,N_26968);
nor U28086 (N_28086,N_25287,N_26157);
xor U28087 (N_28087,N_27473,N_25667);
nor U28088 (N_28088,N_25435,N_25970);
and U28089 (N_28089,N_25227,N_25401);
nand U28090 (N_28090,N_25579,N_25297);
and U28091 (N_28091,N_26502,N_25528);
or U28092 (N_28092,N_27489,N_27040);
nor U28093 (N_28093,N_26432,N_26891);
or U28094 (N_28094,N_25833,N_25494);
and U28095 (N_28095,N_25172,N_26927);
or U28096 (N_28096,N_26826,N_25358);
nor U28097 (N_28097,N_27131,N_25175);
xor U28098 (N_28098,N_26150,N_25595);
nand U28099 (N_28099,N_27245,N_26055);
xnor U28100 (N_28100,N_26971,N_26701);
nor U28101 (N_28101,N_25131,N_25493);
or U28102 (N_28102,N_27130,N_25997);
and U28103 (N_28103,N_26211,N_25806);
or U28104 (N_28104,N_25210,N_26498);
nor U28105 (N_28105,N_26345,N_26546);
nand U28106 (N_28106,N_26193,N_26598);
xnor U28107 (N_28107,N_27359,N_26514);
nand U28108 (N_28108,N_25782,N_26182);
nor U28109 (N_28109,N_26814,N_27308);
xnor U28110 (N_28110,N_25328,N_26425);
nor U28111 (N_28111,N_26402,N_26095);
nand U28112 (N_28112,N_26414,N_25866);
xnor U28113 (N_28113,N_26975,N_25312);
or U28114 (N_28114,N_27278,N_25719);
or U28115 (N_28115,N_27153,N_26484);
or U28116 (N_28116,N_25903,N_25636);
xor U28117 (N_28117,N_26521,N_25219);
nand U28118 (N_28118,N_26375,N_27312);
nor U28119 (N_28119,N_25269,N_26475);
nand U28120 (N_28120,N_25027,N_26067);
nand U28121 (N_28121,N_26044,N_25766);
xnor U28122 (N_28122,N_26326,N_26812);
nand U28123 (N_28123,N_27255,N_25952);
nand U28124 (N_28124,N_27141,N_26267);
xnor U28125 (N_28125,N_26511,N_26677);
nor U28126 (N_28126,N_26387,N_27169);
or U28127 (N_28127,N_25502,N_26527);
nor U28128 (N_28128,N_25681,N_25333);
nor U28129 (N_28129,N_27249,N_26492);
and U28130 (N_28130,N_25462,N_26126);
nand U28131 (N_28131,N_26585,N_25190);
xnor U28132 (N_28132,N_25368,N_27352);
xor U28133 (N_28133,N_25340,N_26805);
nand U28134 (N_28134,N_25152,N_26241);
xor U28135 (N_28135,N_27318,N_25216);
or U28136 (N_28136,N_26525,N_26877);
nor U28137 (N_28137,N_27056,N_27096);
nand U28138 (N_28138,N_27009,N_25097);
nand U28139 (N_28139,N_26581,N_25651);
or U28140 (N_28140,N_25242,N_27299);
or U28141 (N_28141,N_26128,N_25050);
or U28142 (N_28142,N_26853,N_25203);
or U28143 (N_28143,N_27440,N_27151);
or U28144 (N_28144,N_25529,N_26046);
or U28145 (N_28145,N_25741,N_26169);
or U28146 (N_28146,N_26183,N_25147);
nor U28147 (N_28147,N_26887,N_25858);
nor U28148 (N_28148,N_25682,N_25120);
nand U28149 (N_28149,N_25938,N_27450);
nand U28150 (N_28150,N_27015,N_25876);
nand U28151 (N_28151,N_25783,N_26215);
nor U28152 (N_28152,N_27187,N_25725);
nand U28153 (N_28153,N_26052,N_26993);
or U28154 (N_28154,N_26495,N_25523);
or U28155 (N_28155,N_26504,N_27424);
nand U28156 (N_28156,N_25427,N_26149);
nand U28157 (N_28157,N_27023,N_25698);
nor U28158 (N_28158,N_26562,N_27285);
or U28159 (N_28159,N_25391,N_26997);
or U28160 (N_28160,N_25425,N_25981);
nor U28161 (N_28161,N_27011,N_25040);
or U28162 (N_28162,N_25272,N_25006);
and U28163 (N_28163,N_27127,N_25768);
nand U28164 (N_28164,N_27270,N_25047);
and U28165 (N_28165,N_26185,N_27393);
nand U28166 (N_28166,N_26869,N_27284);
xnor U28167 (N_28167,N_26439,N_27322);
and U28168 (N_28168,N_27059,N_25123);
nand U28169 (N_28169,N_27383,N_26726);
nand U28170 (N_28170,N_25991,N_26729);
xor U28171 (N_28171,N_25153,N_25215);
nand U28172 (N_28172,N_25311,N_25377);
and U28173 (N_28173,N_26657,N_27379);
and U28174 (N_28174,N_26274,N_25669);
nand U28175 (N_28175,N_25083,N_25659);
and U28176 (N_28176,N_25517,N_25121);
and U28177 (N_28177,N_25379,N_25458);
or U28178 (N_28178,N_25739,N_26624);
nor U28179 (N_28179,N_26933,N_25861);
xnor U28180 (N_28180,N_26978,N_26532);
or U28181 (N_28181,N_25533,N_26072);
and U28182 (N_28182,N_25630,N_25944);
nor U28183 (N_28183,N_26793,N_25396);
or U28184 (N_28184,N_27360,N_26710);
xor U28185 (N_28185,N_25249,N_26118);
and U28186 (N_28186,N_26491,N_25257);
nor U28187 (N_28187,N_26045,N_26659);
nand U28188 (N_28188,N_25718,N_26478);
xnor U28189 (N_28189,N_25732,N_26373);
nor U28190 (N_28190,N_26867,N_26889);
nand U28191 (N_28191,N_26057,N_25868);
xnor U28192 (N_28192,N_25545,N_25460);
or U28193 (N_28193,N_26259,N_26638);
nand U28194 (N_28194,N_25845,N_26158);
xor U28195 (N_28195,N_26195,N_25978);
and U28196 (N_28196,N_26424,N_27289);
or U28197 (N_28197,N_26162,N_26098);
nand U28198 (N_28198,N_26878,N_26893);
and U28199 (N_28199,N_25402,N_25192);
nand U28200 (N_28200,N_26074,N_25503);
or U28201 (N_28201,N_26002,N_27170);
or U28202 (N_28202,N_26925,N_25498);
nand U28203 (N_28203,N_26693,N_26175);
nor U28204 (N_28204,N_26025,N_25024);
nand U28205 (N_28205,N_27451,N_26548);
nor U28206 (N_28206,N_27431,N_26094);
and U28207 (N_28207,N_26907,N_26797);
or U28208 (N_28208,N_26344,N_27049);
or U28209 (N_28209,N_27172,N_25956);
and U28210 (N_28210,N_25488,N_26396);
nor U28211 (N_28211,N_26538,N_26619);
or U28212 (N_28212,N_26443,N_26917);
and U28213 (N_28213,N_26835,N_26436);
nor U28214 (N_28214,N_26654,N_26736);
and U28215 (N_28215,N_26145,N_26451);
xor U28216 (N_28216,N_25093,N_27387);
and U28217 (N_28217,N_26001,N_25196);
and U28218 (N_28218,N_26866,N_25457);
nand U28219 (N_28219,N_25731,N_26932);
nand U28220 (N_28220,N_25622,N_26676);
and U28221 (N_28221,N_26875,N_27342);
nand U28222 (N_28222,N_25386,N_25011);
nor U28223 (N_28223,N_25150,N_25477);
and U28224 (N_28224,N_25309,N_26712);
xnor U28225 (N_28225,N_26249,N_26972);
nand U28226 (N_28226,N_27061,N_27066);
nand U28227 (N_28227,N_26281,N_25577);
nand U28228 (N_28228,N_25308,N_25831);
and U28229 (N_28229,N_26802,N_27314);
and U28230 (N_28230,N_25429,N_25629);
or U28231 (N_28231,N_25512,N_25646);
and U28232 (N_28232,N_26431,N_25222);
and U28233 (N_28233,N_26355,N_25777);
and U28234 (N_28234,N_27483,N_25243);
and U28235 (N_28235,N_25240,N_26688);
nor U28236 (N_28236,N_27382,N_26322);
nor U28237 (N_28237,N_27276,N_26251);
nor U28238 (N_28238,N_25090,N_27421);
nand U28239 (N_28239,N_26476,N_27442);
and U28240 (N_28240,N_26332,N_25550);
or U28241 (N_28241,N_25886,N_25971);
nand U28242 (N_28242,N_26953,N_26738);
or U28243 (N_28243,N_26564,N_26245);
nor U28244 (N_28244,N_26035,N_25052);
nand U28245 (N_28245,N_25648,N_25590);
or U28246 (N_28246,N_26079,N_26632);
or U28247 (N_28247,N_26254,N_25802);
xnor U28248 (N_28248,N_25459,N_26977);
xor U28249 (N_28249,N_26958,N_26698);
xnor U28250 (N_28250,N_27134,N_27210);
nand U28251 (N_28251,N_26324,N_27486);
or U28252 (N_28252,N_25439,N_26784);
nand U28253 (N_28253,N_25891,N_27158);
nand U28254 (N_28254,N_25930,N_25128);
and U28255 (N_28255,N_26666,N_27013);
xnor U28256 (N_28256,N_25037,N_25031);
xnor U28257 (N_28257,N_26353,N_27128);
nand U28258 (N_28258,N_26578,N_27192);
or U28259 (N_28259,N_26122,N_25224);
or U28260 (N_28260,N_25316,N_25319);
xor U28261 (N_28261,N_26255,N_25628);
nor U28262 (N_28262,N_26918,N_26257);
nand U28263 (N_28263,N_26342,N_27355);
nand U28264 (N_28264,N_26461,N_25879);
xnor U28265 (N_28265,N_27029,N_25264);
or U28266 (N_28266,N_27329,N_25092);
and U28267 (N_28267,N_26667,N_25004);
or U28268 (N_28268,N_27006,N_27054);
and U28269 (N_28269,N_26571,N_26716);
nand U28270 (N_28270,N_25887,N_26737);
or U28271 (N_28271,N_25241,N_26081);
and U28272 (N_28272,N_25795,N_25441);
and U28273 (N_28273,N_25703,N_27494);
and U28274 (N_28274,N_25197,N_27271);
nand U28275 (N_28275,N_26599,N_26800);
xnor U28276 (N_28276,N_25607,N_26490);
nand U28277 (N_28277,N_25526,N_25798);
nor U28278 (N_28278,N_25314,N_26367);
or U28279 (N_28279,N_26499,N_25271);
xor U28280 (N_28280,N_26506,N_26946);
nand U28281 (N_28281,N_27109,N_26089);
xor U28282 (N_28282,N_27224,N_26543);
or U28283 (N_28283,N_27095,N_26301);
xnor U28284 (N_28284,N_27354,N_26774);
nor U28285 (N_28285,N_26776,N_26939);
xnor U28286 (N_28286,N_25912,N_26300);
xnor U28287 (N_28287,N_27034,N_26630);
or U28288 (N_28288,N_25290,N_25170);
nor U28289 (N_28289,N_25568,N_25112);
nand U28290 (N_28290,N_26007,N_25884);
nor U28291 (N_28291,N_26724,N_25522);
or U28292 (N_28292,N_26173,N_27371);
or U28293 (N_28293,N_25549,N_26206);
nand U28294 (N_28294,N_27422,N_25262);
nand U28295 (N_28295,N_25564,N_26970);
and U28296 (N_28296,N_27326,N_25743);
xor U28297 (N_28297,N_25613,N_25035);
and U28298 (N_28298,N_26224,N_27381);
or U28299 (N_28299,N_26610,N_25338);
nor U28300 (N_28300,N_25827,N_25764);
and U28301 (N_28301,N_25054,N_26486);
nor U28302 (N_28302,N_25916,N_26299);
nor U28303 (N_28303,N_25299,N_25895);
or U28304 (N_28304,N_25915,N_26920);
xnor U28305 (N_28305,N_26767,N_25267);
nor U28306 (N_28306,N_27413,N_26606);
or U28307 (N_28307,N_25563,N_27110);
nor U28308 (N_28308,N_25068,N_27339);
nor U28309 (N_28309,N_25539,N_27107);
and U28310 (N_28310,N_25890,N_26393);
or U28311 (N_28311,N_26751,N_27202);
and U28312 (N_28312,N_26076,N_25639);
nand U28313 (N_28313,N_25836,N_27336);
xor U28314 (N_28314,N_26196,N_25995);
nor U28315 (N_28315,N_25780,N_26680);
nand U28316 (N_28316,N_25134,N_25638);
or U28317 (N_28317,N_25384,N_26515);
xor U28318 (N_28318,N_26862,N_26830);
nand U28319 (N_28319,N_26329,N_27227);
and U28320 (N_28320,N_25369,N_25352);
and U28321 (N_28321,N_26121,N_27343);
xor U28322 (N_28322,N_27079,N_25530);
and U28323 (N_28323,N_25841,N_26991);
nor U28324 (N_28324,N_25654,N_25835);
nand U28325 (N_28325,N_26383,N_25066);
and U28326 (N_28326,N_25156,N_26446);
xor U28327 (N_28327,N_26489,N_26306);
nor U28328 (N_28328,N_26640,N_25232);
or U28329 (N_28329,N_26117,N_27123);
or U28330 (N_28330,N_26022,N_25479);
or U28331 (N_28331,N_26406,N_26832);
and U28332 (N_28332,N_26910,N_27145);
xnor U28333 (N_28333,N_26225,N_25616);
nor U28334 (N_28334,N_27430,N_25089);
nand U28335 (N_28335,N_25169,N_26374);
nand U28336 (N_28336,N_25801,N_26563);
xor U28337 (N_28337,N_26813,N_27380);
and U28338 (N_28338,N_27062,N_27427);
and U28339 (N_28339,N_27397,N_25235);
or U28340 (N_28340,N_25449,N_26253);
xor U28341 (N_28341,N_26426,N_25929);
nand U28342 (N_28342,N_25497,N_26708);
and U28343 (N_28343,N_26589,N_27092);
or U28344 (N_28344,N_27163,N_25072);
xnor U28345 (N_28345,N_26873,N_27415);
or U28346 (N_28346,N_26049,N_27274);
nand U28347 (N_28347,N_25602,N_25182);
xnor U28348 (N_28348,N_27027,N_26219);
and U28349 (N_28349,N_27012,N_25983);
and U28350 (N_28350,N_25676,N_25444);
xor U28351 (N_28351,N_26091,N_26360);
nand U28352 (N_28352,N_25039,N_26449);
nand U28353 (N_28353,N_25180,N_25451);
nand U28354 (N_28354,N_27165,N_26423);
and U28355 (N_28355,N_25204,N_25353);
xnor U28356 (N_28356,N_25623,N_26120);
xnor U28357 (N_28357,N_26844,N_26124);
nor U28358 (N_28358,N_25554,N_26777);
nand U28359 (N_28359,N_25988,N_26894);
xor U28360 (N_28360,N_25655,N_27042);
or U28361 (N_28361,N_25019,N_25088);
and U28362 (N_28362,N_25813,N_26441);
nor U28363 (N_28363,N_26559,N_25388);
xnor U28364 (N_28364,N_25600,N_25014);
nand U28365 (N_28365,N_27407,N_25485);
xnor U28366 (N_28366,N_26595,N_25649);
nand U28367 (N_28367,N_26979,N_26384);
nor U28368 (N_28368,N_25258,N_26645);
xnor U28369 (N_28369,N_25318,N_27185);
xor U28370 (N_28370,N_26786,N_25537);
nand U28371 (N_28371,N_27157,N_25653);
or U28372 (N_28372,N_27214,N_27236);
nor U28373 (N_28373,N_26796,N_26999);
nand U28374 (N_28374,N_26474,N_25706);
and U28375 (N_28375,N_25114,N_26628);
xnor U28376 (N_28376,N_26000,N_27216);
and U28377 (N_28377,N_25926,N_25138);
or U28378 (N_28378,N_25419,N_25161);
nand U28379 (N_28379,N_25817,N_27028);
xor U28380 (N_28380,N_26477,N_27405);
or U28381 (N_28381,N_25423,N_26573);
nand U28382 (N_28382,N_25525,N_25122);
and U28383 (N_28383,N_25199,N_26781);
xor U28384 (N_28384,N_25584,N_25059);
nand U28385 (N_28385,N_25818,N_27375);
or U28386 (N_28386,N_25466,N_25996);
and U28387 (N_28387,N_25346,N_26895);
nand U28388 (N_28388,N_26261,N_25680);
nor U28389 (N_28389,N_25277,N_26339);
or U28390 (N_28390,N_26622,N_26199);
nor U28391 (N_28391,N_26596,N_27132);
or U28392 (N_28392,N_26469,N_26535);
nand U28393 (N_28393,N_26587,N_25922);
and U28394 (N_28394,N_27205,N_26151);
nor U28395 (N_28395,N_27150,N_25067);
xnor U28396 (N_28396,N_25487,N_25392);
nor U28397 (N_28397,N_27067,N_27420);
and U28398 (N_28398,N_27239,N_26352);
nand U28399 (N_28399,N_27304,N_27474);
and U28400 (N_28400,N_25770,N_26325);
and U28401 (N_28401,N_26764,N_26362);
and U28402 (N_28402,N_26723,N_25644);
or U28403 (N_28403,N_25286,N_27496);
and U28404 (N_28404,N_26629,N_27384);
nor U28405 (N_28405,N_26378,N_27093);
nor U28406 (N_28406,N_25848,N_25885);
xnor U28407 (N_28407,N_25946,N_25294);
or U28408 (N_28408,N_26171,N_27462);
or U28409 (N_28409,N_26850,N_26408);
and U28410 (N_28410,N_25711,N_27018);
nand U28411 (N_28411,N_26697,N_25454);
xor U28412 (N_28412,N_25021,N_25957);
or U28413 (N_28413,N_26078,N_26750);
and U28414 (N_28414,N_26404,N_26085);
and U28415 (N_28415,N_27008,N_26855);
xor U28416 (N_28416,N_27184,N_25411);
and U28417 (N_28417,N_26131,N_26100);
nor U28418 (N_28418,N_26692,N_26936);
xnor U28419 (N_28419,N_26174,N_26691);
xnor U28420 (N_28420,N_25939,N_26197);
nand U28421 (N_28421,N_26307,N_25023);
xor U28422 (N_28422,N_25982,N_27485);
nor U28423 (N_28423,N_25543,N_27275);
nor U28424 (N_28424,N_25234,N_27103);
nor U28425 (N_28425,N_25964,N_25820);
nor U28426 (N_28426,N_25575,N_25656);
xnor U28427 (N_28427,N_26618,N_26090);
nand U28428 (N_28428,N_27410,N_27260);
or U28429 (N_28429,N_26841,N_26434);
xor U28430 (N_28430,N_26024,N_25274);
xnor U28431 (N_28431,N_25531,N_26313);
xor U28432 (N_28432,N_26994,N_27488);
nand U28433 (N_28433,N_25375,N_26714);
and U28434 (N_28434,N_25417,N_26815);
nand U28435 (N_28435,N_26675,N_26330);
nand U28436 (N_28436,N_26806,N_27433);
and U28437 (N_28437,N_25344,N_25907);
nor U28438 (N_28438,N_27426,N_26109);
nand U28439 (N_28439,N_25979,N_25793);
and U28440 (N_28440,N_26898,N_25164);
or U28441 (N_28441,N_25509,N_26711);
xnor U28442 (N_28442,N_27247,N_27348);
xnor U28443 (N_28443,N_26989,N_27492);
or U28444 (N_28444,N_26903,N_27207);
or U28445 (N_28445,N_26102,N_26272);
nand U28446 (N_28446,N_27084,N_26752);
or U28447 (N_28447,N_26321,N_25714);
and U28448 (N_28448,N_26643,N_27188);
xnor U28449 (N_28449,N_26170,N_25672);
xor U28450 (N_28450,N_26481,N_25959);
or U28451 (N_28451,N_27455,N_25238);
or U28452 (N_28452,N_25753,N_26462);
or U28453 (N_28453,N_27311,N_25260);
or U28454 (N_28454,N_26059,N_26356);
or U28455 (N_28455,N_26913,N_25755);
nand U28456 (N_28456,N_25518,N_25606);
xnor U28457 (N_28457,N_26114,N_26584);
and U28458 (N_28458,N_25599,N_25642);
nand U28459 (N_28459,N_25062,N_25486);
nor U28460 (N_28460,N_25115,N_25747);
and U28461 (N_28461,N_25873,N_26092);
and U28462 (N_28462,N_27464,N_26899);
or U28463 (N_28463,N_26915,N_25527);
nand U28464 (N_28464,N_27388,N_26422);
nor U28465 (N_28465,N_25505,N_25661);
and U28466 (N_28466,N_26348,N_26651);
or U28467 (N_28467,N_25869,N_25051);
or U28468 (N_28468,N_25159,N_25699);
nand U28469 (N_28469,N_27423,N_26685);
nand U28470 (N_28470,N_25562,N_26082);
and U28471 (N_28471,N_27138,N_25871);
xor U28472 (N_28472,N_25226,N_26568);
xor U28473 (N_28473,N_26613,N_25506);
and U28474 (N_28474,N_25685,N_26433);
nand U28475 (N_28475,N_26410,N_27478);
and U28476 (N_28476,N_25515,N_25673);
xor U28477 (N_28477,N_25571,N_25263);
and U28478 (N_28478,N_27156,N_25165);
nor U28479 (N_28479,N_25534,N_25481);
and U28480 (N_28480,N_25436,N_26699);
or U28481 (N_28481,N_26247,N_27144);
xor U28482 (N_28482,N_27113,N_26213);
xnor U28483 (N_28483,N_25759,N_25807);
nand U28484 (N_28484,N_25433,N_26276);
nor U28485 (N_28485,N_25350,N_25118);
and U28486 (N_28486,N_25504,N_27358);
or U28487 (N_28487,N_25284,N_26702);
or U28488 (N_28488,N_25865,N_26464);
or U28489 (N_28489,N_25559,N_25683);
xor U28490 (N_28490,N_26754,N_25632);
or U28491 (N_28491,N_25536,N_25771);
nor U28492 (N_28492,N_27115,N_26652);
and U28493 (N_28493,N_27307,N_25569);
nand U28494 (N_28494,N_26430,N_25857);
nor U28495 (N_28495,N_25508,N_26570);
nor U28496 (N_28496,N_27279,N_25295);
nor U28497 (N_28497,N_26992,N_27457);
xnor U28498 (N_28498,N_27414,N_26615);
and U28499 (N_28499,N_27168,N_27400);
or U28500 (N_28500,N_25285,N_25603);
and U28501 (N_28501,N_25399,N_26314);
and U28502 (N_28502,N_25684,N_27211);
nand U28503 (N_28503,N_27377,N_26937);
nand U28504 (N_28504,N_25941,N_27460);
xnor U28505 (N_28505,N_25860,N_26605);
nor U28506 (N_28506,N_26429,N_26069);
or U28507 (N_28507,N_25154,N_26220);
and U28508 (N_28508,N_25042,N_25990);
nand U28509 (N_28509,N_26207,N_26608);
nand U28510 (N_28510,N_26551,N_27149);
and U28511 (N_28511,N_26931,N_26286);
and U28512 (N_28512,N_26228,N_27112);
xor U28513 (N_28513,N_27135,N_25382);
nor U28514 (N_28514,N_25291,N_26517);
xor U28515 (N_28515,N_25470,N_26905);
nand U28516 (N_28516,N_26112,N_26181);
nand U28517 (N_28517,N_26107,N_25206);
nand U28518 (N_28518,N_25137,N_27363);
nor U28519 (N_28519,N_26298,N_26062);
or U28520 (N_28520,N_25963,N_27173);
or U28521 (N_28521,N_26440,N_25356);
or U28522 (N_28522,N_25373,N_26529);
or U28523 (N_28523,N_25724,N_25099);
and U28524 (N_28524,N_25909,N_27310);
nor U28525 (N_28525,N_25716,N_25179);
and U28526 (N_28526,N_25958,N_26269);
xnor U28527 (N_28527,N_25133,N_26715);
or U28528 (N_28528,N_26405,N_27449);
nor U28529 (N_28529,N_25700,N_26467);
nor U28530 (N_28530,N_26956,N_26650);
or U28531 (N_28531,N_25950,N_27331);
and U28532 (N_28532,N_26823,N_26950);
or U28533 (N_28533,N_25461,N_26923);
and U28534 (N_28534,N_26558,N_25339);
or U28535 (N_28535,N_25931,N_25586);
or U28536 (N_28536,N_27177,N_26160);
xor U28537 (N_28537,N_26017,N_27071);
nor U28538 (N_28538,N_27340,N_25113);
and U28539 (N_28539,N_25273,N_26003);
and U28540 (N_28540,N_25354,N_26620);
nor U28541 (N_28541,N_25999,N_26011);
and U28542 (N_28542,N_26824,N_27218);
nand U28543 (N_28543,N_27251,N_25016);
xor U28544 (N_28544,N_26058,N_27493);
nand U28545 (N_28545,N_25846,N_26827);
and U28546 (N_28546,N_27435,N_26051);
or U28547 (N_28547,N_25482,N_26266);
or U28548 (N_28548,N_27174,N_25359);
xor U28549 (N_28549,N_25744,N_27344);
nor U28550 (N_28550,N_26239,N_25143);
xnor U28551 (N_28551,N_25070,N_25002);
and U28552 (N_28552,N_25524,N_26497);
or U28553 (N_28553,N_25207,N_26611);
nand U28554 (N_28554,N_26450,N_26060);
xnor U28555 (N_28555,N_25668,N_25581);
nor U28556 (N_28556,N_26033,N_25265);
nor U28557 (N_28557,N_25796,N_25933);
nor U28558 (N_28558,N_25228,N_26954);
and U28559 (N_28559,N_26957,N_27301);
and U28560 (N_28560,N_27179,N_26250);
xnor U28561 (N_28561,N_26522,N_25225);
and U28562 (N_28562,N_25992,N_26854);
and U28563 (N_28563,N_25065,N_25521);
nand U28564 (N_28564,N_26167,N_25043);
or U28565 (N_28565,N_25111,N_25927);
and U28566 (N_28566,N_26026,N_25905);
and U28567 (N_28567,N_26634,N_26503);
nor U28568 (N_28568,N_25029,N_26034);
and U28569 (N_28569,N_27373,N_26212);
xnor U28570 (N_28570,N_25245,N_25772);
nand U28571 (N_28571,N_26223,N_26661);
and U28572 (N_28572,N_25301,N_27159);
xor U28573 (N_28573,N_25862,N_26705);
nand U28574 (N_28574,N_25188,N_25735);
nand U28575 (N_28575,N_27078,N_27264);
and U28576 (N_28576,N_25904,N_27404);
xnor U28577 (N_28577,N_25061,N_25400);
nand U28578 (N_28578,N_25728,N_27246);
and U28579 (N_28579,N_26524,N_26626);
or U28580 (N_28580,N_25323,N_25101);
and U28581 (N_28581,N_25363,N_25615);
and U28582 (N_28582,N_25567,N_27136);
and U28583 (N_28583,N_27441,N_26366);
xor U28584 (N_28584,N_26743,N_26064);
or U28585 (N_28585,N_25937,N_26646);
or U28586 (N_28586,N_26208,N_25349);
nand U28587 (N_28587,N_26783,N_26135);
or U28588 (N_28588,N_25594,N_26310);
and U28589 (N_28589,N_27005,N_26395);
or U28590 (N_28590,N_27191,N_26974);
nand U28591 (N_28591,N_25317,N_26944);
xnor U28592 (N_28592,N_26428,N_27481);
or U28593 (N_28593,N_26673,N_26516);
xnor U28594 (N_28594,N_26512,N_26104);
nand U28595 (N_28595,N_25036,N_26744);
and U28596 (N_28596,N_27334,N_25844);
xnor U28597 (N_28597,N_27281,N_26309);
xnor U28598 (N_28598,N_25849,N_25675);
xnor U28599 (N_28599,N_27347,N_25229);
nand U28600 (N_28600,N_26816,N_27201);
or U28601 (N_28601,N_25102,N_27305);
xor U28602 (N_28602,N_26457,N_26327);
or U28603 (N_28603,N_26969,N_26021);
or U28604 (N_28604,N_26831,N_26038);
nand U28605 (N_28605,N_25194,N_27291);
xor U28606 (N_28606,N_27412,N_27443);
or U28607 (N_28607,N_25383,N_26390);
nand U28608 (N_28608,N_25145,N_27463);
nand U28609 (N_28609,N_27180,N_25662);
nor U28610 (N_28610,N_26665,N_25095);
nand U28611 (N_28611,N_27232,N_25686);
nand U28612 (N_28612,N_26496,N_25116);
nor U28613 (N_28613,N_27362,N_26554);
nor U28614 (N_28614,N_27225,N_26837);
and U28615 (N_28615,N_25962,N_27349);
and U28616 (N_28616,N_27139,N_27479);
nand U28617 (N_28617,N_25208,N_25665);
and U28618 (N_28618,N_27070,N_25729);
or U28619 (N_28619,N_27295,N_25954);
nor U28620 (N_28620,N_25405,N_25064);
and U28621 (N_28621,N_25604,N_25513);
or U28622 (N_28622,N_26127,N_25438);
or U28623 (N_28623,N_25315,N_26445);
or U28624 (N_28624,N_26110,N_26857);
and U28625 (N_28625,N_27124,N_25168);
nand U28626 (N_28626,N_26036,N_27046);
or U28627 (N_28627,N_26829,N_26798);
and U28628 (N_28628,N_25932,N_27099);
nor U28629 (N_28629,N_25148,N_27267);
and U28630 (N_28630,N_26108,N_25738);
nand U28631 (N_28631,N_25357,N_25883);
xor U28632 (N_28632,N_27482,N_26376);
and U28633 (N_28633,N_27303,N_25626);
xor U28634 (N_28634,N_26553,N_26473);
or U28635 (N_28635,N_26987,N_25789);
and U28636 (N_28636,N_27337,N_27065);
nor U28637 (N_28637,N_25671,N_27335);
nand U28638 (N_28638,N_26015,N_26242);
xor U28639 (N_28639,N_26292,N_26748);
or U28640 (N_28640,N_26288,N_26681);
and U28641 (N_28641,N_27002,N_26050);
nand U28642 (N_28642,N_25495,N_27351);
nor U28643 (N_28643,N_25184,N_26919);
nand U28644 (N_28644,N_27183,N_25307);
nand U28645 (N_28645,N_27402,N_25151);
nand U28646 (N_28646,N_27445,N_27073);
xnor U28647 (N_28647,N_26164,N_25364);
or U28648 (N_28648,N_26203,N_25348);
or U28649 (N_28649,N_25189,N_26115);
and U28650 (N_28650,N_26929,N_25816);
nand U28651 (N_28651,N_25705,N_25464);
and U28652 (N_28652,N_25555,N_26859);
or U28653 (N_28653,N_25478,N_26612);
nand U28654 (N_28654,N_26258,N_25936);
nor U28655 (N_28655,N_26014,N_27306);
nand U28656 (N_28656,N_26315,N_26073);
xor U28657 (N_28657,N_26103,N_27213);
xor U28658 (N_28658,N_27000,N_26741);
and U28659 (N_28659,N_25424,N_26083);
or U28660 (N_28660,N_26016,N_27223);
nand U28661 (N_28661,N_27418,N_25058);
nand U28662 (N_28662,N_25968,N_26142);
and U28663 (N_28663,N_27117,N_27212);
and U28664 (N_28664,N_25288,N_26817);
or U28665 (N_28665,N_25652,N_26722);
and U28666 (N_28666,N_25974,N_27209);
nand U28667 (N_28667,N_27484,N_26372);
nand U28668 (N_28668,N_26755,N_25476);
or U28669 (N_28669,N_26369,N_25585);
nand U28670 (N_28670,N_25026,N_26200);
or U28671 (N_28671,N_27104,N_27048);
nor U28672 (N_28672,N_25385,N_25737);
nand U28673 (N_28673,N_27369,N_26795);
nand U28674 (N_28674,N_26955,N_25761);
nand U28675 (N_28675,N_27237,N_25975);
and U28676 (N_28676,N_26031,N_26908);
xnor U28677 (N_28677,N_26460,N_26156);
xnor U28678 (N_28678,N_25322,N_27370);
and U28679 (N_28679,N_25910,N_26874);
nand U28680 (N_28680,N_26583,N_26704);
nor U28681 (N_28681,N_27022,N_26463);
xnor U28682 (N_28682,N_25038,N_27001);
nand U28683 (N_28683,N_27055,N_26633);
or U28684 (N_28684,N_25465,N_27425);
or U28685 (N_28685,N_25020,N_27126);
nand U28686 (N_28686,N_26202,N_25544);
xnor U28687 (N_28687,N_26567,N_25412);
and U28688 (N_28688,N_25303,N_26343);
nor U28689 (N_28689,N_25985,N_25578);
and U28690 (N_28690,N_25110,N_26594);
nor U28691 (N_28691,N_25901,N_25715);
xor U28692 (N_28692,N_26545,N_25829);
and U28693 (N_28693,N_26597,N_27417);
and U28694 (N_28694,N_26631,N_25149);
or U28695 (N_28695,N_27368,N_25900);
xor U28696 (N_28696,N_27406,N_25601);
or U28697 (N_28697,N_25825,N_26555);
nand U28698 (N_28698,N_25200,N_27072);
or U28699 (N_28699,N_27021,N_27319);
xor U28700 (N_28700,N_27143,N_27350);
or U28701 (N_28701,N_25565,N_25573);
and U28702 (N_28702,N_25393,N_26733);
nand U28703 (N_28703,N_26509,N_25774);
nand U28704 (N_28704,N_25332,N_26198);
xnor U28705 (N_28705,N_27476,N_27269);
nor U28706 (N_28706,N_26642,N_26066);
nand U28707 (N_28707,N_26775,N_26084);
nor U28708 (N_28708,N_25803,N_26678);
xnor U28709 (N_28709,N_25471,N_27088);
and U28710 (N_28710,N_26349,N_25896);
xor U28711 (N_28711,N_25572,N_26398);
xnor U28712 (N_28712,N_26839,N_26452);
and U28713 (N_28713,N_25426,N_26879);
or U28714 (N_28714,N_26656,N_25942);
or U28715 (N_28715,N_26792,N_27438);
xor U28716 (N_28716,N_26088,N_25597);
nor U28717 (N_28717,N_25327,N_25945);
xnor U28718 (N_28718,N_26427,N_26695);
nor U28719 (N_28719,N_25205,N_27376);
xnor U28720 (N_28720,N_25679,N_27076);
and U28721 (N_28721,N_26155,N_27477);
nand U28722 (N_28722,N_26938,N_26709);
nand U28723 (N_28723,N_26739,N_26435);
or U28724 (N_28724,N_27262,N_27024);
xnor U28725 (N_28725,N_26099,N_25450);
or U28726 (N_28726,N_26413,N_25810);
or U28727 (N_28727,N_26232,N_26020);
and U28728 (N_28728,N_25967,N_27399);
nand U28729 (N_28729,N_26988,N_25872);
and U28730 (N_28730,N_25591,N_27364);
nand U28731 (N_28731,N_27357,N_27487);
and U28732 (N_28732,N_25733,N_26951);
and U28733 (N_28733,N_25834,N_25815);
and U28734 (N_28734,N_25492,N_25966);
xor U28735 (N_28735,N_25709,N_27235);
nand U28736 (N_28736,N_25691,N_25965);
nand U28737 (N_28737,N_26995,N_27395);
or U28738 (N_28738,N_26861,N_27033);
or U28739 (N_28739,N_25270,N_26870);
nor U28740 (N_28740,N_26718,N_27330);
nand U28741 (N_28741,N_26447,N_25362);
nor U28742 (N_28742,N_27069,N_25859);
nand U28743 (N_28743,N_25614,N_26032);
xor U28744 (N_28744,N_26096,N_25214);
nand U28745 (N_28745,N_26296,N_27016);
nor U28746 (N_28746,N_25406,N_26949);
or U28747 (N_28747,N_25566,N_26468);
xor U28748 (N_28748,N_26071,N_27290);
or U28749 (N_28749,N_26179,N_26663);
xor U28750 (N_28750,N_27153,N_27032);
or U28751 (N_28751,N_26132,N_26416);
nor U28752 (N_28752,N_27240,N_25001);
nand U28753 (N_28753,N_26092,N_26166);
nor U28754 (N_28754,N_27091,N_26477);
xnor U28755 (N_28755,N_26323,N_25816);
or U28756 (N_28756,N_25665,N_27021);
xor U28757 (N_28757,N_25140,N_26031);
xor U28758 (N_28758,N_26054,N_26601);
nand U28759 (N_28759,N_25140,N_25476);
nor U28760 (N_28760,N_26273,N_25951);
nor U28761 (N_28761,N_26821,N_25457);
nor U28762 (N_28762,N_26662,N_26444);
or U28763 (N_28763,N_25631,N_27437);
nor U28764 (N_28764,N_25618,N_25698);
xor U28765 (N_28765,N_25435,N_26143);
and U28766 (N_28766,N_25495,N_27170);
or U28767 (N_28767,N_26601,N_25651);
nand U28768 (N_28768,N_26910,N_25917);
or U28769 (N_28769,N_25135,N_27097);
nor U28770 (N_28770,N_25268,N_25052);
or U28771 (N_28771,N_27498,N_27240);
and U28772 (N_28772,N_25055,N_25775);
or U28773 (N_28773,N_25887,N_26252);
nor U28774 (N_28774,N_25409,N_25322);
nor U28775 (N_28775,N_26516,N_26475);
or U28776 (N_28776,N_25085,N_27360);
nand U28777 (N_28777,N_26509,N_25158);
or U28778 (N_28778,N_26206,N_26175);
or U28779 (N_28779,N_26460,N_26385);
and U28780 (N_28780,N_26913,N_25512);
or U28781 (N_28781,N_26554,N_25592);
and U28782 (N_28782,N_25319,N_26140);
nand U28783 (N_28783,N_26262,N_25583);
and U28784 (N_28784,N_27426,N_26735);
or U28785 (N_28785,N_27341,N_26298);
or U28786 (N_28786,N_26535,N_27001);
nor U28787 (N_28787,N_25194,N_26592);
nand U28788 (N_28788,N_25687,N_26094);
and U28789 (N_28789,N_27187,N_25565);
xor U28790 (N_28790,N_27323,N_26845);
xor U28791 (N_28791,N_27186,N_26852);
and U28792 (N_28792,N_25160,N_25699);
and U28793 (N_28793,N_25442,N_26403);
nor U28794 (N_28794,N_25224,N_27145);
nand U28795 (N_28795,N_27239,N_26672);
xnor U28796 (N_28796,N_25848,N_25843);
xnor U28797 (N_28797,N_25919,N_27109);
or U28798 (N_28798,N_26949,N_25871);
or U28799 (N_28799,N_26780,N_26808);
and U28800 (N_28800,N_25840,N_25836);
xor U28801 (N_28801,N_27322,N_25758);
or U28802 (N_28802,N_25268,N_25853);
nand U28803 (N_28803,N_25339,N_27028);
nand U28804 (N_28804,N_25418,N_27179);
nand U28805 (N_28805,N_25368,N_26312);
and U28806 (N_28806,N_27037,N_25315);
or U28807 (N_28807,N_25720,N_27228);
xnor U28808 (N_28808,N_26259,N_26708);
and U28809 (N_28809,N_25688,N_26650);
and U28810 (N_28810,N_25645,N_26068);
or U28811 (N_28811,N_27078,N_25473);
nor U28812 (N_28812,N_25525,N_27365);
nor U28813 (N_28813,N_27364,N_26725);
and U28814 (N_28814,N_26647,N_26709);
and U28815 (N_28815,N_27169,N_25123);
or U28816 (N_28816,N_26996,N_25124);
nor U28817 (N_28817,N_25766,N_25452);
xor U28818 (N_28818,N_26405,N_26973);
nor U28819 (N_28819,N_27390,N_27053);
xnor U28820 (N_28820,N_25721,N_27245);
nor U28821 (N_28821,N_26058,N_25638);
or U28822 (N_28822,N_25703,N_25456);
or U28823 (N_28823,N_26260,N_25785);
nand U28824 (N_28824,N_26382,N_25924);
and U28825 (N_28825,N_25758,N_26244);
nor U28826 (N_28826,N_27329,N_26328);
xor U28827 (N_28827,N_26313,N_27277);
or U28828 (N_28828,N_26968,N_27065);
and U28829 (N_28829,N_26095,N_26759);
nand U28830 (N_28830,N_26195,N_25368);
and U28831 (N_28831,N_25065,N_25258);
and U28832 (N_28832,N_25865,N_26055);
nand U28833 (N_28833,N_27189,N_25548);
nand U28834 (N_28834,N_27001,N_26048);
xor U28835 (N_28835,N_27408,N_26053);
nor U28836 (N_28836,N_26246,N_25200);
nor U28837 (N_28837,N_25777,N_25770);
nor U28838 (N_28838,N_27456,N_26167);
and U28839 (N_28839,N_25030,N_25142);
or U28840 (N_28840,N_25829,N_27274);
or U28841 (N_28841,N_25135,N_27166);
nor U28842 (N_28842,N_25846,N_25447);
nor U28843 (N_28843,N_26693,N_25846);
and U28844 (N_28844,N_26376,N_25937);
nand U28845 (N_28845,N_26094,N_25585);
xnor U28846 (N_28846,N_25068,N_25657);
and U28847 (N_28847,N_26949,N_26722);
nor U28848 (N_28848,N_26525,N_27110);
xnor U28849 (N_28849,N_25855,N_26621);
nand U28850 (N_28850,N_26918,N_26026);
xor U28851 (N_28851,N_26895,N_26608);
nor U28852 (N_28852,N_25650,N_25903);
or U28853 (N_28853,N_25658,N_25867);
nor U28854 (N_28854,N_26062,N_26033);
nor U28855 (N_28855,N_25448,N_25606);
nor U28856 (N_28856,N_25877,N_26011);
and U28857 (N_28857,N_25421,N_25537);
xnor U28858 (N_28858,N_26395,N_26905);
nand U28859 (N_28859,N_26612,N_25659);
nor U28860 (N_28860,N_25563,N_25677);
and U28861 (N_28861,N_27269,N_26985);
nor U28862 (N_28862,N_26594,N_25423);
xor U28863 (N_28863,N_25926,N_25391);
nor U28864 (N_28864,N_25002,N_25518);
nor U28865 (N_28865,N_25373,N_25338);
or U28866 (N_28866,N_27214,N_25781);
and U28867 (N_28867,N_27104,N_26967);
nand U28868 (N_28868,N_26837,N_26492);
xnor U28869 (N_28869,N_27460,N_25663);
nand U28870 (N_28870,N_26945,N_26300);
or U28871 (N_28871,N_25701,N_26964);
or U28872 (N_28872,N_25914,N_25732);
nor U28873 (N_28873,N_26706,N_27074);
or U28874 (N_28874,N_25961,N_25863);
nor U28875 (N_28875,N_25849,N_26024);
or U28876 (N_28876,N_27283,N_26435);
nor U28877 (N_28877,N_25753,N_27280);
nor U28878 (N_28878,N_26530,N_25989);
nand U28879 (N_28879,N_26773,N_26709);
nor U28880 (N_28880,N_25152,N_26332);
nor U28881 (N_28881,N_25376,N_27134);
or U28882 (N_28882,N_25093,N_26788);
and U28883 (N_28883,N_25421,N_26271);
nand U28884 (N_28884,N_26784,N_26386);
nor U28885 (N_28885,N_25229,N_27213);
nor U28886 (N_28886,N_27197,N_26269);
and U28887 (N_28887,N_25853,N_26066);
and U28888 (N_28888,N_25399,N_25959);
nor U28889 (N_28889,N_25163,N_25645);
or U28890 (N_28890,N_26428,N_27286);
or U28891 (N_28891,N_25743,N_26687);
nor U28892 (N_28892,N_25661,N_25909);
or U28893 (N_28893,N_26062,N_27080);
and U28894 (N_28894,N_25134,N_25240);
xor U28895 (N_28895,N_26766,N_25914);
nor U28896 (N_28896,N_25075,N_25882);
and U28897 (N_28897,N_25445,N_26527);
and U28898 (N_28898,N_26955,N_25585);
xnor U28899 (N_28899,N_25945,N_25072);
or U28900 (N_28900,N_25728,N_26310);
xor U28901 (N_28901,N_26742,N_25769);
nor U28902 (N_28902,N_25264,N_26220);
or U28903 (N_28903,N_27358,N_25537);
nor U28904 (N_28904,N_25018,N_25379);
or U28905 (N_28905,N_27401,N_26751);
or U28906 (N_28906,N_26502,N_25697);
nor U28907 (N_28907,N_25602,N_25682);
xnor U28908 (N_28908,N_26189,N_25626);
or U28909 (N_28909,N_25177,N_25848);
nor U28910 (N_28910,N_26267,N_26890);
nor U28911 (N_28911,N_26770,N_26991);
nand U28912 (N_28912,N_25154,N_25520);
nor U28913 (N_28913,N_25524,N_26156);
and U28914 (N_28914,N_27052,N_27006);
and U28915 (N_28915,N_25939,N_25203);
nand U28916 (N_28916,N_26384,N_25870);
nand U28917 (N_28917,N_25964,N_26959);
nand U28918 (N_28918,N_25991,N_26109);
xor U28919 (N_28919,N_25869,N_27038);
and U28920 (N_28920,N_27324,N_27197);
nor U28921 (N_28921,N_26430,N_25391);
and U28922 (N_28922,N_26195,N_25155);
and U28923 (N_28923,N_26870,N_27469);
or U28924 (N_28924,N_27257,N_25277);
and U28925 (N_28925,N_26209,N_27250);
nor U28926 (N_28926,N_27495,N_26666);
xor U28927 (N_28927,N_26925,N_27299);
and U28928 (N_28928,N_26046,N_25917);
nor U28929 (N_28929,N_26086,N_25696);
or U28930 (N_28930,N_26580,N_25557);
xnor U28931 (N_28931,N_27328,N_27465);
nand U28932 (N_28932,N_26164,N_27137);
and U28933 (N_28933,N_25763,N_27320);
and U28934 (N_28934,N_27027,N_25179);
nand U28935 (N_28935,N_26593,N_26188);
nor U28936 (N_28936,N_27321,N_26415);
xor U28937 (N_28937,N_26349,N_25703);
or U28938 (N_28938,N_27340,N_25871);
and U28939 (N_28939,N_27204,N_26214);
nor U28940 (N_28940,N_26166,N_26443);
and U28941 (N_28941,N_25417,N_25376);
or U28942 (N_28942,N_26696,N_25358);
xnor U28943 (N_28943,N_26129,N_25544);
nand U28944 (N_28944,N_25642,N_26730);
xor U28945 (N_28945,N_25782,N_26922);
nor U28946 (N_28946,N_25696,N_25474);
and U28947 (N_28947,N_27053,N_25656);
or U28948 (N_28948,N_25175,N_26893);
nor U28949 (N_28949,N_26360,N_25090);
or U28950 (N_28950,N_25363,N_26005);
and U28951 (N_28951,N_26510,N_27139);
nor U28952 (N_28952,N_27330,N_26567);
nand U28953 (N_28953,N_25189,N_25036);
nand U28954 (N_28954,N_25727,N_27084);
nand U28955 (N_28955,N_25990,N_27447);
xnor U28956 (N_28956,N_27111,N_27015);
nand U28957 (N_28957,N_26761,N_25974);
nand U28958 (N_28958,N_26946,N_25161);
xor U28959 (N_28959,N_27141,N_25924);
or U28960 (N_28960,N_25474,N_26244);
nor U28961 (N_28961,N_26516,N_26170);
xnor U28962 (N_28962,N_25343,N_27130);
or U28963 (N_28963,N_27159,N_25898);
nor U28964 (N_28964,N_26133,N_26251);
xnor U28965 (N_28965,N_27341,N_26079);
nor U28966 (N_28966,N_26707,N_26577);
and U28967 (N_28967,N_25323,N_25488);
nand U28968 (N_28968,N_25772,N_26230);
or U28969 (N_28969,N_27062,N_27367);
xnor U28970 (N_28970,N_27291,N_26889);
and U28971 (N_28971,N_26275,N_26708);
nand U28972 (N_28972,N_26923,N_26542);
nor U28973 (N_28973,N_26023,N_25001);
nand U28974 (N_28974,N_26335,N_26714);
and U28975 (N_28975,N_25459,N_26701);
nor U28976 (N_28976,N_25716,N_27495);
or U28977 (N_28977,N_25598,N_26257);
or U28978 (N_28978,N_26145,N_25627);
nand U28979 (N_28979,N_26586,N_25260);
and U28980 (N_28980,N_27273,N_26769);
nor U28981 (N_28981,N_25396,N_25416);
or U28982 (N_28982,N_25891,N_25376);
and U28983 (N_28983,N_26283,N_27110);
xnor U28984 (N_28984,N_25622,N_25784);
nor U28985 (N_28985,N_26166,N_25649);
nor U28986 (N_28986,N_27417,N_27132);
nand U28987 (N_28987,N_27325,N_25673);
nor U28988 (N_28988,N_25891,N_26118);
and U28989 (N_28989,N_25359,N_26132);
and U28990 (N_28990,N_26780,N_26710);
nor U28991 (N_28991,N_26841,N_25939);
or U28992 (N_28992,N_25222,N_26628);
xor U28993 (N_28993,N_26785,N_26772);
nor U28994 (N_28994,N_26883,N_27209);
nand U28995 (N_28995,N_25109,N_26607);
or U28996 (N_28996,N_25541,N_27301);
and U28997 (N_28997,N_25971,N_25654);
or U28998 (N_28998,N_27121,N_26746);
and U28999 (N_28999,N_27302,N_27323);
xnor U29000 (N_29000,N_26493,N_25215);
and U29001 (N_29001,N_26566,N_26020);
and U29002 (N_29002,N_25395,N_26403);
nor U29003 (N_29003,N_26314,N_25618);
nand U29004 (N_29004,N_26456,N_25024);
and U29005 (N_29005,N_27001,N_26460);
nor U29006 (N_29006,N_25482,N_27315);
and U29007 (N_29007,N_25773,N_26094);
or U29008 (N_29008,N_25350,N_25112);
or U29009 (N_29009,N_26486,N_25794);
xor U29010 (N_29010,N_26005,N_27300);
or U29011 (N_29011,N_26141,N_25540);
or U29012 (N_29012,N_25133,N_25303);
xnor U29013 (N_29013,N_26439,N_27215);
nand U29014 (N_29014,N_26295,N_25348);
xnor U29015 (N_29015,N_26290,N_25294);
or U29016 (N_29016,N_25037,N_26691);
or U29017 (N_29017,N_26676,N_25521);
nor U29018 (N_29018,N_25693,N_26368);
and U29019 (N_29019,N_26445,N_27426);
nand U29020 (N_29020,N_25986,N_26467);
nor U29021 (N_29021,N_26272,N_26018);
or U29022 (N_29022,N_25008,N_25476);
nor U29023 (N_29023,N_26606,N_26079);
nand U29024 (N_29024,N_27115,N_26025);
xnor U29025 (N_29025,N_27181,N_25599);
or U29026 (N_29026,N_26874,N_26651);
nand U29027 (N_29027,N_26144,N_25724);
and U29028 (N_29028,N_25727,N_25800);
nand U29029 (N_29029,N_25858,N_26161);
or U29030 (N_29030,N_25201,N_26943);
and U29031 (N_29031,N_25939,N_26714);
nand U29032 (N_29032,N_25405,N_26857);
nor U29033 (N_29033,N_26457,N_26155);
nor U29034 (N_29034,N_27208,N_27150);
xnor U29035 (N_29035,N_26721,N_27140);
or U29036 (N_29036,N_26525,N_27017);
nor U29037 (N_29037,N_25523,N_27192);
nor U29038 (N_29038,N_25990,N_27464);
and U29039 (N_29039,N_26544,N_27243);
nor U29040 (N_29040,N_26075,N_25968);
and U29041 (N_29041,N_27020,N_26321);
and U29042 (N_29042,N_25512,N_25683);
nand U29043 (N_29043,N_26929,N_26582);
xor U29044 (N_29044,N_26760,N_27037);
nand U29045 (N_29045,N_26985,N_26787);
and U29046 (N_29046,N_26160,N_25697);
or U29047 (N_29047,N_26811,N_25815);
nor U29048 (N_29048,N_25122,N_27141);
or U29049 (N_29049,N_27055,N_25425);
and U29050 (N_29050,N_25426,N_27475);
xor U29051 (N_29051,N_27089,N_26415);
and U29052 (N_29052,N_25317,N_26142);
and U29053 (N_29053,N_25637,N_25377);
xor U29054 (N_29054,N_26916,N_25090);
or U29055 (N_29055,N_26684,N_26837);
nand U29056 (N_29056,N_26866,N_26194);
xor U29057 (N_29057,N_25065,N_26438);
or U29058 (N_29058,N_27084,N_25072);
and U29059 (N_29059,N_27055,N_25940);
or U29060 (N_29060,N_26551,N_25037);
nor U29061 (N_29061,N_26606,N_27154);
nand U29062 (N_29062,N_25467,N_25425);
nor U29063 (N_29063,N_27356,N_26434);
nand U29064 (N_29064,N_27281,N_26467);
nor U29065 (N_29065,N_26688,N_26306);
or U29066 (N_29066,N_27001,N_25029);
nor U29067 (N_29067,N_25922,N_26611);
nor U29068 (N_29068,N_25222,N_26949);
nand U29069 (N_29069,N_26648,N_26732);
nand U29070 (N_29070,N_25289,N_26931);
nor U29071 (N_29071,N_25406,N_25512);
and U29072 (N_29072,N_26728,N_25654);
nand U29073 (N_29073,N_25540,N_26855);
nand U29074 (N_29074,N_26838,N_26869);
xor U29075 (N_29075,N_27062,N_27449);
xnor U29076 (N_29076,N_25099,N_26988);
and U29077 (N_29077,N_25464,N_26707);
nor U29078 (N_29078,N_27311,N_26909);
xnor U29079 (N_29079,N_26577,N_25562);
nand U29080 (N_29080,N_25432,N_27416);
and U29081 (N_29081,N_25694,N_27209);
or U29082 (N_29082,N_27391,N_25918);
xor U29083 (N_29083,N_25233,N_25684);
or U29084 (N_29084,N_26158,N_26876);
or U29085 (N_29085,N_26507,N_25677);
or U29086 (N_29086,N_27093,N_27253);
and U29087 (N_29087,N_25925,N_25218);
xor U29088 (N_29088,N_25676,N_26643);
nand U29089 (N_29089,N_27165,N_27217);
nor U29090 (N_29090,N_25683,N_25794);
nand U29091 (N_29091,N_26218,N_25920);
nand U29092 (N_29092,N_26671,N_25169);
nor U29093 (N_29093,N_26322,N_25352);
and U29094 (N_29094,N_26021,N_25234);
nand U29095 (N_29095,N_25383,N_25556);
nand U29096 (N_29096,N_26013,N_26231);
nand U29097 (N_29097,N_26262,N_25511);
and U29098 (N_29098,N_27114,N_25517);
nand U29099 (N_29099,N_26545,N_25073);
and U29100 (N_29100,N_27105,N_25118);
nand U29101 (N_29101,N_25783,N_25308);
nand U29102 (N_29102,N_25969,N_25837);
nor U29103 (N_29103,N_26413,N_26101);
and U29104 (N_29104,N_26107,N_25577);
and U29105 (N_29105,N_25023,N_26036);
nand U29106 (N_29106,N_27171,N_25761);
nor U29107 (N_29107,N_26666,N_25952);
and U29108 (N_29108,N_27156,N_26009);
xnor U29109 (N_29109,N_26337,N_26303);
and U29110 (N_29110,N_27293,N_25690);
or U29111 (N_29111,N_27174,N_25327);
nand U29112 (N_29112,N_25450,N_26909);
and U29113 (N_29113,N_26702,N_26413);
and U29114 (N_29114,N_25164,N_25491);
nor U29115 (N_29115,N_25869,N_25293);
nor U29116 (N_29116,N_27492,N_25802);
and U29117 (N_29117,N_27093,N_26438);
nand U29118 (N_29118,N_25599,N_26490);
nand U29119 (N_29119,N_26391,N_27462);
or U29120 (N_29120,N_25214,N_26453);
nand U29121 (N_29121,N_25147,N_26063);
and U29122 (N_29122,N_27460,N_27492);
nor U29123 (N_29123,N_26755,N_26055);
nor U29124 (N_29124,N_26029,N_27077);
xnor U29125 (N_29125,N_25456,N_25423);
nor U29126 (N_29126,N_26640,N_25116);
and U29127 (N_29127,N_25304,N_26592);
nor U29128 (N_29128,N_26531,N_27272);
xor U29129 (N_29129,N_26332,N_25883);
or U29130 (N_29130,N_27001,N_25662);
nand U29131 (N_29131,N_27221,N_25730);
xor U29132 (N_29132,N_26611,N_25589);
nor U29133 (N_29133,N_25514,N_26991);
nor U29134 (N_29134,N_27361,N_26422);
and U29135 (N_29135,N_25854,N_25367);
or U29136 (N_29136,N_26823,N_25182);
xor U29137 (N_29137,N_27135,N_27179);
and U29138 (N_29138,N_26092,N_26136);
xnor U29139 (N_29139,N_26925,N_27090);
nor U29140 (N_29140,N_25835,N_25449);
nor U29141 (N_29141,N_27271,N_25061);
or U29142 (N_29142,N_26989,N_26327);
nand U29143 (N_29143,N_26214,N_25538);
or U29144 (N_29144,N_25371,N_27229);
nor U29145 (N_29145,N_25194,N_25124);
nor U29146 (N_29146,N_26860,N_26447);
and U29147 (N_29147,N_26160,N_25484);
nor U29148 (N_29148,N_26676,N_27368);
nand U29149 (N_29149,N_25852,N_25090);
xor U29150 (N_29150,N_26836,N_25542);
and U29151 (N_29151,N_26963,N_25424);
nor U29152 (N_29152,N_27336,N_26835);
and U29153 (N_29153,N_25912,N_27142);
or U29154 (N_29154,N_25876,N_27375);
and U29155 (N_29155,N_26024,N_26858);
nor U29156 (N_29156,N_27341,N_25152);
nand U29157 (N_29157,N_27148,N_27453);
xor U29158 (N_29158,N_25616,N_27079);
nand U29159 (N_29159,N_26844,N_26298);
or U29160 (N_29160,N_25341,N_26603);
xor U29161 (N_29161,N_25835,N_26593);
xor U29162 (N_29162,N_25672,N_25890);
xnor U29163 (N_29163,N_25789,N_25638);
xor U29164 (N_29164,N_25506,N_26384);
nand U29165 (N_29165,N_26629,N_27122);
or U29166 (N_29166,N_25315,N_26706);
xor U29167 (N_29167,N_25514,N_25874);
nand U29168 (N_29168,N_25395,N_26941);
nand U29169 (N_29169,N_27270,N_25330);
and U29170 (N_29170,N_27044,N_26280);
xnor U29171 (N_29171,N_27376,N_26426);
and U29172 (N_29172,N_26932,N_27431);
xor U29173 (N_29173,N_27025,N_26936);
nor U29174 (N_29174,N_27373,N_25619);
and U29175 (N_29175,N_27097,N_26929);
nor U29176 (N_29176,N_25861,N_26902);
nand U29177 (N_29177,N_27424,N_26996);
nand U29178 (N_29178,N_26794,N_25471);
nand U29179 (N_29179,N_26219,N_25501);
nor U29180 (N_29180,N_26506,N_25521);
xnor U29181 (N_29181,N_25383,N_25815);
nor U29182 (N_29182,N_27358,N_25749);
nor U29183 (N_29183,N_25466,N_27094);
or U29184 (N_29184,N_26710,N_26198);
and U29185 (N_29185,N_27342,N_27276);
nand U29186 (N_29186,N_25976,N_25265);
and U29187 (N_29187,N_27315,N_27418);
xnor U29188 (N_29188,N_26546,N_25733);
or U29189 (N_29189,N_25697,N_27351);
or U29190 (N_29190,N_25975,N_26105);
nand U29191 (N_29191,N_25872,N_25156);
nor U29192 (N_29192,N_25833,N_25938);
or U29193 (N_29193,N_25319,N_26088);
xor U29194 (N_29194,N_26226,N_26731);
or U29195 (N_29195,N_27048,N_26219);
or U29196 (N_29196,N_27260,N_25171);
and U29197 (N_29197,N_27132,N_25940);
and U29198 (N_29198,N_27398,N_25376);
or U29199 (N_29199,N_27349,N_27147);
nand U29200 (N_29200,N_25117,N_25532);
xor U29201 (N_29201,N_26308,N_26047);
or U29202 (N_29202,N_25817,N_26520);
xor U29203 (N_29203,N_26835,N_25120);
nor U29204 (N_29204,N_26278,N_26109);
nor U29205 (N_29205,N_26958,N_25387);
or U29206 (N_29206,N_27248,N_26110);
nand U29207 (N_29207,N_26971,N_26667);
and U29208 (N_29208,N_26344,N_25058);
or U29209 (N_29209,N_25839,N_25744);
xor U29210 (N_29210,N_25114,N_26812);
or U29211 (N_29211,N_26511,N_25148);
nor U29212 (N_29212,N_26968,N_25212);
and U29213 (N_29213,N_25189,N_25263);
or U29214 (N_29214,N_25851,N_26180);
and U29215 (N_29215,N_26529,N_26760);
and U29216 (N_29216,N_26605,N_26241);
nor U29217 (N_29217,N_25984,N_27263);
nand U29218 (N_29218,N_25129,N_25603);
nor U29219 (N_29219,N_25720,N_26657);
and U29220 (N_29220,N_25120,N_26623);
nor U29221 (N_29221,N_26325,N_26223);
and U29222 (N_29222,N_27138,N_27330);
and U29223 (N_29223,N_26047,N_25836);
or U29224 (N_29224,N_27453,N_26837);
nor U29225 (N_29225,N_27475,N_25495);
nand U29226 (N_29226,N_27388,N_26091);
nor U29227 (N_29227,N_25097,N_25416);
and U29228 (N_29228,N_26811,N_25190);
and U29229 (N_29229,N_26330,N_26138);
and U29230 (N_29230,N_26361,N_27130);
or U29231 (N_29231,N_25579,N_25228);
xor U29232 (N_29232,N_26017,N_25660);
and U29233 (N_29233,N_27323,N_26731);
xor U29234 (N_29234,N_26761,N_26944);
nand U29235 (N_29235,N_26135,N_26839);
nand U29236 (N_29236,N_26446,N_26391);
and U29237 (N_29237,N_25219,N_25277);
nor U29238 (N_29238,N_27250,N_26890);
and U29239 (N_29239,N_26297,N_25562);
nand U29240 (N_29240,N_27317,N_27176);
and U29241 (N_29241,N_27085,N_27373);
and U29242 (N_29242,N_25675,N_25124);
or U29243 (N_29243,N_25971,N_25074);
nor U29244 (N_29244,N_25999,N_27045);
or U29245 (N_29245,N_26441,N_27142);
and U29246 (N_29246,N_25683,N_27456);
or U29247 (N_29247,N_26325,N_26004);
nand U29248 (N_29248,N_27309,N_25559);
nor U29249 (N_29249,N_26967,N_26359);
and U29250 (N_29250,N_25928,N_26365);
xor U29251 (N_29251,N_26211,N_25453);
nor U29252 (N_29252,N_26850,N_25597);
nor U29253 (N_29253,N_27385,N_25414);
nand U29254 (N_29254,N_25167,N_27211);
nor U29255 (N_29255,N_25172,N_27396);
xnor U29256 (N_29256,N_27126,N_26428);
and U29257 (N_29257,N_25079,N_25967);
and U29258 (N_29258,N_26088,N_27148);
or U29259 (N_29259,N_26570,N_25482);
and U29260 (N_29260,N_27240,N_27496);
and U29261 (N_29261,N_26582,N_26457);
and U29262 (N_29262,N_26079,N_27438);
and U29263 (N_29263,N_25343,N_25822);
nand U29264 (N_29264,N_26786,N_25785);
or U29265 (N_29265,N_26265,N_26319);
and U29266 (N_29266,N_25077,N_25055);
or U29267 (N_29267,N_27176,N_25138);
and U29268 (N_29268,N_25639,N_25996);
and U29269 (N_29269,N_27080,N_25573);
and U29270 (N_29270,N_25501,N_25972);
nor U29271 (N_29271,N_25428,N_26242);
nor U29272 (N_29272,N_26224,N_25325);
nor U29273 (N_29273,N_26300,N_25440);
xor U29274 (N_29274,N_26973,N_26303);
nor U29275 (N_29275,N_26760,N_26331);
nand U29276 (N_29276,N_27460,N_25286);
nor U29277 (N_29277,N_26743,N_25662);
nand U29278 (N_29278,N_26206,N_25548);
xor U29279 (N_29279,N_25889,N_25796);
or U29280 (N_29280,N_25576,N_25480);
and U29281 (N_29281,N_25472,N_26768);
or U29282 (N_29282,N_25405,N_26299);
xor U29283 (N_29283,N_25328,N_26717);
nor U29284 (N_29284,N_25542,N_27023);
and U29285 (N_29285,N_25201,N_26383);
or U29286 (N_29286,N_25397,N_25362);
nor U29287 (N_29287,N_25415,N_27248);
nand U29288 (N_29288,N_27335,N_26033);
xor U29289 (N_29289,N_25652,N_25618);
and U29290 (N_29290,N_26699,N_27182);
nor U29291 (N_29291,N_25929,N_27494);
or U29292 (N_29292,N_25627,N_27209);
nor U29293 (N_29293,N_26017,N_25823);
nand U29294 (N_29294,N_26793,N_26070);
and U29295 (N_29295,N_25457,N_25890);
nand U29296 (N_29296,N_26334,N_26221);
or U29297 (N_29297,N_26142,N_26826);
nand U29298 (N_29298,N_25602,N_25648);
or U29299 (N_29299,N_25762,N_26975);
xnor U29300 (N_29300,N_27233,N_26497);
and U29301 (N_29301,N_27188,N_25035);
xnor U29302 (N_29302,N_27484,N_26522);
xor U29303 (N_29303,N_26952,N_25589);
or U29304 (N_29304,N_25908,N_26736);
nor U29305 (N_29305,N_25114,N_26605);
nand U29306 (N_29306,N_27284,N_26649);
nor U29307 (N_29307,N_25774,N_27267);
or U29308 (N_29308,N_27276,N_27435);
nor U29309 (N_29309,N_26050,N_26181);
nand U29310 (N_29310,N_26217,N_26620);
nand U29311 (N_29311,N_26911,N_27074);
xnor U29312 (N_29312,N_25970,N_27076);
nand U29313 (N_29313,N_26642,N_25951);
nor U29314 (N_29314,N_26850,N_26917);
or U29315 (N_29315,N_25210,N_27066);
xor U29316 (N_29316,N_26716,N_25098);
nand U29317 (N_29317,N_27054,N_26091);
or U29318 (N_29318,N_25625,N_26273);
nand U29319 (N_29319,N_25247,N_26091);
nand U29320 (N_29320,N_25610,N_25311);
and U29321 (N_29321,N_25666,N_26123);
or U29322 (N_29322,N_26438,N_25023);
nor U29323 (N_29323,N_25778,N_25199);
nand U29324 (N_29324,N_25654,N_27206);
nand U29325 (N_29325,N_25886,N_26440);
xor U29326 (N_29326,N_25896,N_25826);
and U29327 (N_29327,N_25188,N_25161);
nor U29328 (N_29328,N_26299,N_25350);
nand U29329 (N_29329,N_27109,N_27195);
nand U29330 (N_29330,N_26385,N_26775);
and U29331 (N_29331,N_27291,N_25731);
nor U29332 (N_29332,N_27301,N_25564);
nand U29333 (N_29333,N_25139,N_25060);
or U29334 (N_29334,N_27428,N_27388);
or U29335 (N_29335,N_26898,N_25594);
nand U29336 (N_29336,N_26265,N_26321);
xor U29337 (N_29337,N_25783,N_26514);
nand U29338 (N_29338,N_25813,N_26403);
xnor U29339 (N_29339,N_25893,N_25566);
nand U29340 (N_29340,N_27105,N_25856);
and U29341 (N_29341,N_25292,N_25175);
nand U29342 (N_29342,N_25299,N_26357);
xnor U29343 (N_29343,N_26309,N_25715);
xnor U29344 (N_29344,N_26944,N_26760);
nand U29345 (N_29345,N_26430,N_26767);
nor U29346 (N_29346,N_25789,N_26753);
nand U29347 (N_29347,N_25792,N_26117);
and U29348 (N_29348,N_26669,N_27001);
xnor U29349 (N_29349,N_25475,N_26999);
xnor U29350 (N_29350,N_25327,N_26199);
nand U29351 (N_29351,N_26784,N_25528);
or U29352 (N_29352,N_26252,N_27128);
and U29353 (N_29353,N_25383,N_27417);
or U29354 (N_29354,N_25106,N_27265);
nand U29355 (N_29355,N_27067,N_26994);
nor U29356 (N_29356,N_27018,N_26818);
nor U29357 (N_29357,N_26517,N_25575);
nor U29358 (N_29358,N_25264,N_26476);
xor U29359 (N_29359,N_25080,N_27454);
xnor U29360 (N_29360,N_26532,N_26210);
and U29361 (N_29361,N_27260,N_26676);
and U29362 (N_29362,N_27106,N_25087);
and U29363 (N_29363,N_25884,N_25776);
xnor U29364 (N_29364,N_25374,N_27191);
or U29365 (N_29365,N_25020,N_26985);
nand U29366 (N_29366,N_25485,N_25103);
nand U29367 (N_29367,N_27482,N_27120);
and U29368 (N_29368,N_25274,N_25433);
nand U29369 (N_29369,N_26827,N_25959);
or U29370 (N_29370,N_26306,N_27063);
or U29371 (N_29371,N_26849,N_26736);
or U29372 (N_29372,N_25267,N_26950);
or U29373 (N_29373,N_27181,N_25694);
nor U29374 (N_29374,N_25056,N_26314);
xnor U29375 (N_29375,N_26330,N_26693);
and U29376 (N_29376,N_27138,N_27333);
nand U29377 (N_29377,N_26541,N_27050);
nor U29378 (N_29378,N_26311,N_25857);
nor U29379 (N_29379,N_27000,N_25524);
xor U29380 (N_29380,N_25553,N_26517);
or U29381 (N_29381,N_27412,N_27200);
xnor U29382 (N_29382,N_25104,N_25231);
or U29383 (N_29383,N_26924,N_26305);
xor U29384 (N_29384,N_27405,N_27062);
or U29385 (N_29385,N_25779,N_26064);
or U29386 (N_29386,N_26177,N_26129);
nor U29387 (N_29387,N_27273,N_25291);
or U29388 (N_29388,N_26346,N_25812);
or U29389 (N_29389,N_25184,N_26687);
or U29390 (N_29390,N_26496,N_25615);
and U29391 (N_29391,N_25131,N_26042);
nand U29392 (N_29392,N_26183,N_26877);
xor U29393 (N_29393,N_26325,N_26837);
nor U29394 (N_29394,N_26167,N_26771);
xor U29395 (N_29395,N_27175,N_26408);
and U29396 (N_29396,N_27454,N_26234);
nor U29397 (N_29397,N_26358,N_25254);
and U29398 (N_29398,N_26479,N_25214);
and U29399 (N_29399,N_25235,N_27302);
nand U29400 (N_29400,N_25523,N_25062);
nor U29401 (N_29401,N_27230,N_27311);
and U29402 (N_29402,N_25144,N_25408);
nand U29403 (N_29403,N_27411,N_26232);
xor U29404 (N_29404,N_25068,N_26106);
nor U29405 (N_29405,N_25534,N_27446);
xnor U29406 (N_29406,N_25363,N_25595);
and U29407 (N_29407,N_25474,N_25419);
xnor U29408 (N_29408,N_25290,N_25414);
or U29409 (N_29409,N_27200,N_25477);
or U29410 (N_29410,N_25458,N_27336);
and U29411 (N_29411,N_27234,N_26430);
nand U29412 (N_29412,N_27039,N_27004);
or U29413 (N_29413,N_26557,N_26493);
xnor U29414 (N_29414,N_26244,N_27118);
or U29415 (N_29415,N_26566,N_26843);
nand U29416 (N_29416,N_25397,N_27147);
and U29417 (N_29417,N_27440,N_26366);
or U29418 (N_29418,N_26466,N_25990);
or U29419 (N_29419,N_26283,N_26257);
and U29420 (N_29420,N_26157,N_27043);
xor U29421 (N_29421,N_25154,N_25287);
and U29422 (N_29422,N_26424,N_26630);
xnor U29423 (N_29423,N_26763,N_26894);
nand U29424 (N_29424,N_25319,N_26363);
and U29425 (N_29425,N_27365,N_25438);
xnor U29426 (N_29426,N_25991,N_25958);
and U29427 (N_29427,N_26069,N_25984);
xor U29428 (N_29428,N_26106,N_25723);
nor U29429 (N_29429,N_25588,N_27087);
or U29430 (N_29430,N_27071,N_26670);
or U29431 (N_29431,N_26166,N_25875);
xor U29432 (N_29432,N_26323,N_26024);
and U29433 (N_29433,N_26221,N_27391);
xor U29434 (N_29434,N_26546,N_27199);
xor U29435 (N_29435,N_25104,N_26952);
nand U29436 (N_29436,N_25728,N_25655);
or U29437 (N_29437,N_25802,N_26081);
or U29438 (N_29438,N_26945,N_26620);
nor U29439 (N_29439,N_25518,N_25533);
and U29440 (N_29440,N_26248,N_27153);
nand U29441 (N_29441,N_27027,N_26099);
xnor U29442 (N_29442,N_25631,N_25466);
nor U29443 (N_29443,N_25831,N_26728);
and U29444 (N_29444,N_25965,N_25150);
nor U29445 (N_29445,N_26247,N_25098);
xnor U29446 (N_29446,N_25113,N_27260);
xnor U29447 (N_29447,N_27411,N_26121);
nand U29448 (N_29448,N_25201,N_25403);
xnor U29449 (N_29449,N_25603,N_25878);
nor U29450 (N_29450,N_27391,N_25434);
and U29451 (N_29451,N_26927,N_27080);
nor U29452 (N_29452,N_27037,N_25154);
or U29453 (N_29453,N_27120,N_27255);
nand U29454 (N_29454,N_27442,N_26235);
or U29455 (N_29455,N_26240,N_26957);
or U29456 (N_29456,N_25036,N_27391);
or U29457 (N_29457,N_26194,N_26682);
and U29458 (N_29458,N_25164,N_26822);
nor U29459 (N_29459,N_26398,N_26827);
nor U29460 (N_29460,N_27409,N_26135);
or U29461 (N_29461,N_25082,N_25607);
and U29462 (N_29462,N_26587,N_27249);
or U29463 (N_29463,N_27229,N_25440);
and U29464 (N_29464,N_25277,N_26908);
and U29465 (N_29465,N_26655,N_27357);
nand U29466 (N_29466,N_26060,N_25186);
nand U29467 (N_29467,N_27184,N_26881);
and U29468 (N_29468,N_26231,N_26776);
nand U29469 (N_29469,N_26692,N_25643);
xor U29470 (N_29470,N_26068,N_26748);
nand U29471 (N_29471,N_26329,N_27061);
nand U29472 (N_29472,N_26094,N_26352);
nand U29473 (N_29473,N_25167,N_27303);
and U29474 (N_29474,N_26645,N_26709);
or U29475 (N_29475,N_26718,N_25010);
or U29476 (N_29476,N_26020,N_25684);
or U29477 (N_29477,N_26455,N_26860);
or U29478 (N_29478,N_26868,N_27036);
nand U29479 (N_29479,N_27464,N_25517);
and U29480 (N_29480,N_27083,N_25804);
nand U29481 (N_29481,N_27307,N_26515);
nor U29482 (N_29482,N_25806,N_27264);
and U29483 (N_29483,N_25020,N_25050);
and U29484 (N_29484,N_25725,N_25925);
or U29485 (N_29485,N_27109,N_27203);
nand U29486 (N_29486,N_25227,N_27264);
nor U29487 (N_29487,N_25391,N_26788);
nand U29488 (N_29488,N_25418,N_25527);
xnor U29489 (N_29489,N_26183,N_26262);
nand U29490 (N_29490,N_25588,N_25188);
nor U29491 (N_29491,N_26088,N_27115);
nor U29492 (N_29492,N_25514,N_26487);
nor U29493 (N_29493,N_25096,N_26383);
and U29494 (N_29494,N_25169,N_25204);
xor U29495 (N_29495,N_27466,N_27103);
xor U29496 (N_29496,N_26748,N_27402);
and U29497 (N_29497,N_27357,N_26210);
nor U29498 (N_29498,N_26806,N_26617);
and U29499 (N_29499,N_25635,N_27327);
nor U29500 (N_29500,N_27388,N_27367);
xnor U29501 (N_29501,N_25799,N_27367);
or U29502 (N_29502,N_25146,N_26323);
and U29503 (N_29503,N_25795,N_25789);
xnor U29504 (N_29504,N_26327,N_26659);
nand U29505 (N_29505,N_25762,N_27393);
xor U29506 (N_29506,N_26256,N_27109);
nor U29507 (N_29507,N_26109,N_27335);
nor U29508 (N_29508,N_27178,N_26167);
xnor U29509 (N_29509,N_26869,N_27411);
xnor U29510 (N_29510,N_27129,N_25833);
xor U29511 (N_29511,N_27064,N_27428);
or U29512 (N_29512,N_26595,N_26063);
nand U29513 (N_29513,N_26979,N_25123);
xnor U29514 (N_29514,N_27262,N_26210);
nand U29515 (N_29515,N_25445,N_27380);
and U29516 (N_29516,N_25256,N_26363);
nor U29517 (N_29517,N_26905,N_26741);
xor U29518 (N_29518,N_25146,N_27415);
xor U29519 (N_29519,N_27367,N_25984);
or U29520 (N_29520,N_25424,N_27061);
nor U29521 (N_29521,N_26807,N_25524);
xnor U29522 (N_29522,N_27202,N_25487);
nor U29523 (N_29523,N_25572,N_26125);
nor U29524 (N_29524,N_26851,N_25290);
nor U29525 (N_29525,N_25700,N_26552);
and U29526 (N_29526,N_25260,N_25262);
nand U29527 (N_29527,N_25451,N_27374);
and U29528 (N_29528,N_26518,N_25002);
xnor U29529 (N_29529,N_25008,N_26742);
and U29530 (N_29530,N_26237,N_26552);
xnor U29531 (N_29531,N_25484,N_26065);
nand U29532 (N_29532,N_27122,N_26059);
nand U29533 (N_29533,N_26067,N_25813);
and U29534 (N_29534,N_26171,N_25488);
and U29535 (N_29535,N_25336,N_25769);
nand U29536 (N_29536,N_26316,N_25032);
nor U29537 (N_29537,N_27233,N_25532);
xor U29538 (N_29538,N_26745,N_26038);
xnor U29539 (N_29539,N_26474,N_26387);
xor U29540 (N_29540,N_27062,N_25018);
xnor U29541 (N_29541,N_27167,N_26911);
nand U29542 (N_29542,N_27335,N_27087);
or U29543 (N_29543,N_25841,N_26885);
or U29544 (N_29544,N_26831,N_27159);
xor U29545 (N_29545,N_25785,N_27492);
and U29546 (N_29546,N_27000,N_27181);
nand U29547 (N_29547,N_26602,N_25625);
nand U29548 (N_29548,N_26790,N_26665);
nand U29549 (N_29549,N_25176,N_25310);
nand U29550 (N_29550,N_25054,N_26729);
nor U29551 (N_29551,N_26700,N_25239);
xor U29552 (N_29552,N_27273,N_25481);
nand U29553 (N_29553,N_27161,N_25532);
nor U29554 (N_29554,N_26002,N_25335);
nor U29555 (N_29555,N_26517,N_26950);
nand U29556 (N_29556,N_25323,N_26075);
or U29557 (N_29557,N_27307,N_27103);
or U29558 (N_29558,N_26046,N_27160);
xor U29559 (N_29559,N_26877,N_25714);
xnor U29560 (N_29560,N_25645,N_25842);
nor U29561 (N_29561,N_26068,N_27196);
or U29562 (N_29562,N_25879,N_26316);
nand U29563 (N_29563,N_26013,N_25724);
or U29564 (N_29564,N_26958,N_25137);
and U29565 (N_29565,N_26392,N_27024);
or U29566 (N_29566,N_25943,N_25579);
or U29567 (N_29567,N_26435,N_26887);
or U29568 (N_29568,N_25300,N_26585);
and U29569 (N_29569,N_26048,N_25391);
and U29570 (N_29570,N_26697,N_25395);
or U29571 (N_29571,N_27294,N_27362);
nor U29572 (N_29572,N_27332,N_25090);
and U29573 (N_29573,N_25986,N_26535);
and U29574 (N_29574,N_26732,N_26442);
or U29575 (N_29575,N_26680,N_25823);
and U29576 (N_29576,N_26696,N_27317);
or U29577 (N_29577,N_25171,N_26062);
and U29578 (N_29578,N_25345,N_25300);
xor U29579 (N_29579,N_25871,N_26766);
xnor U29580 (N_29580,N_26259,N_26384);
or U29581 (N_29581,N_25207,N_26128);
xor U29582 (N_29582,N_26937,N_25452);
and U29583 (N_29583,N_26297,N_26974);
and U29584 (N_29584,N_25046,N_26358);
nor U29585 (N_29585,N_26783,N_27156);
nor U29586 (N_29586,N_25222,N_25551);
and U29587 (N_29587,N_25817,N_27144);
nor U29588 (N_29588,N_26740,N_25673);
or U29589 (N_29589,N_26248,N_25857);
xor U29590 (N_29590,N_26824,N_26378);
nand U29591 (N_29591,N_27166,N_26661);
or U29592 (N_29592,N_26583,N_25232);
nand U29593 (N_29593,N_26117,N_26107);
xnor U29594 (N_29594,N_26012,N_27004);
nand U29595 (N_29595,N_25433,N_26274);
or U29596 (N_29596,N_25400,N_26269);
xor U29597 (N_29597,N_25209,N_25893);
xnor U29598 (N_29598,N_25964,N_26262);
or U29599 (N_29599,N_26664,N_25671);
nor U29600 (N_29600,N_25922,N_25083);
or U29601 (N_29601,N_25918,N_27377);
nand U29602 (N_29602,N_25538,N_26674);
xor U29603 (N_29603,N_27337,N_26619);
nor U29604 (N_29604,N_26625,N_26120);
nand U29605 (N_29605,N_26892,N_27380);
nand U29606 (N_29606,N_26194,N_25236);
xnor U29607 (N_29607,N_27204,N_26276);
and U29608 (N_29608,N_25487,N_27087);
xnor U29609 (N_29609,N_25568,N_26890);
xnor U29610 (N_29610,N_25794,N_27497);
and U29611 (N_29611,N_25212,N_25023);
and U29612 (N_29612,N_25391,N_26927);
and U29613 (N_29613,N_27339,N_25616);
xor U29614 (N_29614,N_25098,N_25564);
or U29615 (N_29615,N_26547,N_25285);
nand U29616 (N_29616,N_25418,N_25723);
nand U29617 (N_29617,N_25875,N_26384);
or U29618 (N_29618,N_26194,N_27321);
or U29619 (N_29619,N_25706,N_26449);
or U29620 (N_29620,N_26962,N_25261);
xor U29621 (N_29621,N_26402,N_27012);
nand U29622 (N_29622,N_26651,N_27009);
nor U29623 (N_29623,N_26638,N_25319);
xor U29624 (N_29624,N_25632,N_25070);
and U29625 (N_29625,N_25500,N_25775);
xor U29626 (N_29626,N_25082,N_27362);
or U29627 (N_29627,N_26880,N_26964);
nor U29628 (N_29628,N_25887,N_25769);
or U29629 (N_29629,N_26938,N_25806);
and U29630 (N_29630,N_25457,N_27416);
nand U29631 (N_29631,N_26101,N_26483);
xnor U29632 (N_29632,N_25410,N_26725);
nor U29633 (N_29633,N_27441,N_25805);
or U29634 (N_29634,N_25495,N_26880);
or U29635 (N_29635,N_25347,N_26555);
nand U29636 (N_29636,N_25606,N_26197);
nor U29637 (N_29637,N_27336,N_25322);
nand U29638 (N_29638,N_26494,N_25911);
nand U29639 (N_29639,N_26096,N_25961);
xor U29640 (N_29640,N_26046,N_27437);
nor U29641 (N_29641,N_25049,N_26886);
nand U29642 (N_29642,N_25170,N_25440);
nor U29643 (N_29643,N_25964,N_25892);
and U29644 (N_29644,N_25730,N_25977);
or U29645 (N_29645,N_27468,N_25382);
nand U29646 (N_29646,N_26168,N_27203);
nor U29647 (N_29647,N_26033,N_25307);
or U29648 (N_29648,N_25618,N_25670);
and U29649 (N_29649,N_25704,N_27335);
and U29650 (N_29650,N_25928,N_26001);
and U29651 (N_29651,N_26058,N_25654);
and U29652 (N_29652,N_26395,N_26337);
xnor U29653 (N_29653,N_25825,N_25563);
and U29654 (N_29654,N_26190,N_25793);
or U29655 (N_29655,N_26695,N_27100);
or U29656 (N_29656,N_25011,N_26790);
nand U29657 (N_29657,N_27089,N_26303);
or U29658 (N_29658,N_26529,N_27411);
and U29659 (N_29659,N_25758,N_26100);
or U29660 (N_29660,N_25837,N_25869);
nor U29661 (N_29661,N_25917,N_26017);
nand U29662 (N_29662,N_26198,N_26358);
or U29663 (N_29663,N_25565,N_25907);
xor U29664 (N_29664,N_27016,N_25716);
nand U29665 (N_29665,N_25880,N_25060);
nand U29666 (N_29666,N_25191,N_27405);
or U29667 (N_29667,N_27004,N_25999);
nor U29668 (N_29668,N_26420,N_26317);
xnor U29669 (N_29669,N_27365,N_26780);
or U29670 (N_29670,N_25437,N_26238);
nor U29671 (N_29671,N_25768,N_25106);
nor U29672 (N_29672,N_25323,N_26485);
and U29673 (N_29673,N_25903,N_27253);
nor U29674 (N_29674,N_25406,N_27369);
xor U29675 (N_29675,N_25202,N_25888);
and U29676 (N_29676,N_26096,N_26113);
or U29677 (N_29677,N_25112,N_25224);
nand U29678 (N_29678,N_27170,N_25677);
nand U29679 (N_29679,N_27051,N_27458);
nand U29680 (N_29680,N_25156,N_27353);
and U29681 (N_29681,N_25164,N_26436);
xor U29682 (N_29682,N_27306,N_26944);
and U29683 (N_29683,N_27480,N_26979);
xor U29684 (N_29684,N_27015,N_26968);
nand U29685 (N_29685,N_27406,N_26788);
xor U29686 (N_29686,N_27409,N_27256);
nor U29687 (N_29687,N_26614,N_26964);
nand U29688 (N_29688,N_25510,N_26793);
nor U29689 (N_29689,N_27001,N_25571);
xor U29690 (N_29690,N_26187,N_25602);
and U29691 (N_29691,N_26098,N_25340);
xor U29692 (N_29692,N_26965,N_27013);
nand U29693 (N_29693,N_26867,N_25312);
xnor U29694 (N_29694,N_27449,N_27464);
xnor U29695 (N_29695,N_27474,N_25629);
xnor U29696 (N_29696,N_27105,N_26532);
and U29697 (N_29697,N_25441,N_25973);
xnor U29698 (N_29698,N_26961,N_26515);
nand U29699 (N_29699,N_26817,N_26846);
and U29700 (N_29700,N_27467,N_25347);
nand U29701 (N_29701,N_26762,N_25188);
xor U29702 (N_29702,N_27008,N_25433);
and U29703 (N_29703,N_25167,N_27457);
nand U29704 (N_29704,N_25569,N_25654);
nor U29705 (N_29705,N_26338,N_25032);
xor U29706 (N_29706,N_25429,N_26667);
and U29707 (N_29707,N_26528,N_25170);
or U29708 (N_29708,N_26046,N_27169);
and U29709 (N_29709,N_26356,N_27073);
and U29710 (N_29710,N_26424,N_25179);
or U29711 (N_29711,N_25314,N_27476);
xor U29712 (N_29712,N_27207,N_26248);
xor U29713 (N_29713,N_25878,N_26564);
xor U29714 (N_29714,N_27452,N_26706);
xnor U29715 (N_29715,N_26510,N_25901);
nand U29716 (N_29716,N_26392,N_25387);
xnor U29717 (N_29717,N_25276,N_26179);
nor U29718 (N_29718,N_26341,N_26919);
or U29719 (N_29719,N_26449,N_25565);
and U29720 (N_29720,N_26628,N_26868);
xor U29721 (N_29721,N_26930,N_25595);
nand U29722 (N_29722,N_27401,N_27400);
nand U29723 (N_29723,N_26708,N_26240);
nor U29724 (N_29724,N_27460,N_26125);
nand U29725 (N_29725,N_27198,N_25824);
xor U29726 (N_29726,N_25325,N_25263);
or U29727 (N_29727,N_26222,N_25791);
or U29728 (N_29728,N_27453,N_26239);
and U29729 (N_29729,N_25955,N_26202);
or U29730 (N_29730,N_26084,N_26874);
and U29731 (N_29731,N_26650,N_27044);
or U29732 (N_29732,N_27413,N_27070);
and U29733 (N_29733,N_25177,N_25522);
and U29734 (N_29734,N_26631,N_27285);
or U29735 (N_29735,N_26896,N_25004);
nor U29736 (N_29736,N_26936,N_26974);
or U29737 (N_29737,N_25696,N_26299);
and U29738 (N_29738,N_26106,N_25055);
or U29739 (N_29739,N_26959,N_27176);
or U29740 (N_29740,N_26917,N_25815);
nor U29741 (N_29741,N_26380,N_26336);
nor U29742 (N_29742,N_27306,N_25692);
nand U29743 (N_29743,N_25094,N_25291);
or U29744 (N_29744,N_25799,N_26958);
and U29745 (N_29745,N_25289,N_27004);
nand U29746 (N_29746,N_26760,N_27309);
nand U29747 (N_29747,N_27186,N_25131);
or U29748 (N_29748,N_26634,N_25183);
or U29749 (N_29749,N_26266,N_25993);
or U29750 (N_29750,N_26138,N_27285);
nand U29751 (N_29751,N_27088,N_26644);
and U29752 (N_29752,N_25320,N_27137);
and U29753 (N_29753,N_25602,N_26831);
nor U29754 (N_29754,N_25583,N_27116);
nor U29755 (N_29755,N_25433,N_25543);
nor U29756 (N_29756,N_25832,N_26361);
nand U29757 (N_29757,N_25253,N_27297);
and U29758 (N_29758,N_26410,N_25219);
and U29759 (N_29759,N_25760,N_25801);
xnor U29760 (N_29760,N_26790,N_25199);
nor U29761 (N_29761,N_26483,N_25703);
nor U29762 (N_29762,N_27373,N_26466);
nand U29763 (N_29763,N_26229,N_25870);
nor U29764 (N_29764,N_27496,N_26310);
nor U29765 (N_29765,N_26093,N_25226);
xnor U29766 (N_29766,N_25812,N_25046);
or U29767 (N_29767,N_26809,N_25450);
or U29768 (N_29768,N_25350,N_26114);
xor U29769 (N_29769,N_27078,N_25405);
and U29770 (N_29770,N_25991,N_25847);
or U29771 (N_29771,N_25592,N_25880);
nand U29772 (N_29772,N_25571,N_25232);
nor U29773 (N_29773,N_26561,N_27402);
nand U29774 (N_29774,N_26799,N_25145);
or U29775 (N_29775,N_27170,N_26888);
and U29776 (N_29776,N_25351,N_27289);
xor U29777 (N_29777,N_25337,N_26900);
nor U29778 (N_29778,N_26888,N_27349);
or U29779 (N_29779,N_25573,N_25216);
xor U29780 (N_29780,N_25016,N_25378);
or U29781 (N_29781,N_27235,N_26073);
and U29782 (N_29782,N_26633,N_25996);
xnor U29783 (N_29783,N_25063,N_25393);
and U29784 (N_29784,N_26686,N_27451);
and U29785 (N_29785,N_26574,N_26047);
and U29786 (N_29786,N_25085,N_25262);
nand U29787 (N_29787,N_26632,N_26793);
xnor U29788 (N_29788,N_25659,N_25021);
or U29789 (N_29789,N_25662,N_25688);
nand U29790 (N_29790,N_25908,N_26299);
nand U29791 (N_29791,N_25274,N_25502);
nor U29792 (N_29792,N_26953,N_26501);
and U29793 (N_29793,N_27045,N_26614);
or U29794 (N_29794,N_25247,N_26117);
and U29795 (N_29795,N_27251,N_25804);
xor U29796 (N_29796,N_25244,N_27256);
xor U29797 (N_29797,N_25847,N_25506);
nand U29798 (N_29798,N_27422,N_25630);
nand U29799 (N_29799,N_26352,N_27374);
and U29800 (N_29800,N_26134,N_26479);
nor U29801 (N_29801,N_25273,N_25430);
nor U29802 (N_29802,N_25073,N_27013);
nor U29803 (N_29803,N_25631,N_25764);
or U29804 (N_29804,N_25264,N_26520);
or U29805 (N_29805,N_25236,N_25782);
xor U29806 (N_29806,N_26284,N_25723);
and U29807 (N_29807,N_25166,N_25107);
nor U29808 (N_29808,N_27370,N_26441);
xnor U29809 (N_29809,N_27391,N_25012);
xnor U29810 (N_29810,N_25322,N_27199);
nand U29811 (N_29811,N_25664,N_26396);
xnor U29812 (N_29812,N_26718,N_26843);
xnor U29813 (N_29813,N_25283,N_26030);
xor U29814 (N_29814,N_26742,N_25807);
and U29815 (N_29815,N_25161,N_27420);
and U29816 (N_29816,N_25458,N_27371);
or U29817 (N_29817,N_27155,N_26001);
nand U29818 (N_29818,N_26761,N_27465);
or U29819 (N_29819,N_26641,N_25085);
xnor U29820 (N_29820,N_26794,N_26991);
nand U29821 (N_29821,N_25248,N_25157);
and U29822 (N_29822,N_25165,N_25713);
or U29823 (N_29823,N_25651,N_27225);
nand U29824 (N_29824,N_25238,N_26481);
xor U29825 (N_29825,N_25745,N_25928);
xnor U29826 (N_29826,N_26922,N_26938);
and U29827 (N_29827,N_25975,N_27490);
nand U29828 (N_29828,N_26042,N_27469);
and U29829 (N_29829,N_27125,N_27429);
nand U29830 (N_29830,N_26782,N_25317);
nand U29831 (N_29831,N_27296,N_25418);
or U29832 (N_29832,N_26298,N_26919);
nand U29833 (N_29833,N_27054,N_26539);
and U29834 (N_29834,N_27195,N_26444);
xnor U29835 (N_29835,N_27263,N_26196);
xor U29836 (N_29836,N_27288,N_27301);
and U29837 (N_29837,N_26102,N_26948);
or U29838 (N_29838,N_27111,N_27304);
nand U29839 (N_29839,N_25216,N_27468);
nand U29840 (N_29840,N_25874,N_25357);
nand U29841 (N_29841,N_27086,N_27197);
nand U29842 (N_29842,N_25952,N_25892);
nand U29843 (N_29843,N_27432,N_25309);
nor U29844 (N_29844,N_25102,N_27272);
nor U29845 (N_29845,N_25536,N_27440);
and U29846 (N_29846,N_27150,N_25347);
nand U29847 (N_29847,N_26694,N_25464);
and U29848 (N_29848,N_25481,N_26654);
nand U29849 (N_29849,N_26268,N_27414);
nor U29850 (N_29850,N_26238,N_26518);
and U29851 (N_29851,N_27407,N_25126);
nor U29852 (N_29852,N_25319,N_26258);
nand U29853 (N_29853,N_26312,N_25406);
nand U29854 (N_29854,N_26227,N_25574);
or U29855 (N_29855,N_25617,N_25197);
nand U29856 (N_29856,N_26389,N_27299);
or U29857 (N_29857,N_25922,N_25361);
nand U29858 (N_29858,N_25500,N_26925);
nor U29859 (N_29859,N_25034,N_25106);
xnor U29860 (N_29860,N_27031,N_26161);
nor U29861 (N_29861,N_25743,N_25778);
or U29862 (N_29862,N_26855,N_25139);
nor U29863 (N_29863,N_27029,N_26910);
or U29864 (N_29864,N_26413,N_25022);
or U29865 (N_29865,N_25490,N_26377);
xnor U29866 (N_29866,N_26503,N_26862);
xor U29867 (N_29867,N_25427,N_26114);
nor U29868 (N_29868,N_25209,N_26274);
or U29869 (N_29869,N_25153,N_27238);
and U29870 (N_29870,N_25661,N_26778);
or U29871 (N_29871,N_25612,N_25713);
nor U29872 (N_29872,N_25639,N_27030);
nand U29873 (N_29873,N_25543,N_26563);
and U29874 (N_29874,N_25848,N_26169);
xnor U29875 (N_29875,N_26966,N_25528);
xor U29876 (N_29876,N_26178,N_25644);
and U29877 (N_29877,N_25146,N_26717);
nand U29878 (N_29878,N_26343,N_25407);
xnor U29879 (N_29879,N_27234,N_26236);
xnor U29880 (N_29880,N_26792,N_26169);
nand U29881 (N_29881,N_25071,N_25887);
nor U29882 (N_29882,N_25176,N_26888);
xnor U29883 (N_29883,N_27120,N_26430);
xnor U29884 (N_29884,N_26022,N_25556);
and U29885 (N_29885,N_25792,N_27456);
and U29886 (N_29886,N_27473,N_25163);
xor U29887 (N_29887,N_25895,N_26152);
nor U29888 (N_29888,N_27276,N_26511);
nand U29889 (N_29889,N_26774,N_25450);
nor U29890 (N_29890,N_25414,N_25430);
xor U29891 (N_29891,N_26507,N_25650);
nand U29892 (N_29892,N_27183,N_26710);
or U29893 (N_29893,N_25167,N_25564);
or U29894 (N_29894,N_27328,N_26878);
nand U29895 (N_29895,N_25276,N_27327);
nand U29896 (N_29896,N_25363,N_27468);
nand U29897 (N_29897,N_25453,N_26601);
xor U29898 (N_29898,N_26905,N_25674);
nand U29899 (N_29899,N_26628,N_27012);
and U29900 (N_29900,N_26695,N_25592);
nor U29901 (N_29901,N_26741,N_27454);
or U29902 (N_29902,N_25179,N_26223);
xnor U29903 (N_29903,N_25534,N_26442);
xnor U29904 (N_29904,N_25117,N_26465);
or U29905 (N_29905,N_26720,N_26014);
nor U29906 (N_29906,N_26883,N_25817);
xnor U29907 (N_29907,N_26096,N_27185);
and U29908 (N_29908,N_27426,N_26299);
nand U29909 (N_29909,N_26580,N_26277);
and U29910 (N_29910,N_27019,N_25246);
nand U29911 (N_29911,N_27020,N_25678);
xor U29912 (N_29912,N_25763,N_26398);
xnor U29913 (N_29913,N_26818,N_26055);
and U29914 (N_29914,N_25114,N_25038);
and U29915 (N_29915,N_25194,N_26831);
or U29916 (N_29916,N_26254,N_26377);
nor U29917 (N_29917,N_25411,N_27300);
xnor U29918 (N_29918,N_25789,N_27183);
xnor U29919 (N_29919,N_27204,N_25679);
nor U29920 (N_29920,N_25014,N_26882);
nand U29921 (N_29921,N_26255,N_26893);
nand U29922 (N_29922,N_25162,N_27197);
nand U29923 (N_29923,N_25716,N_26719);
nor U29924 (N_29924,N_26408,N_25493);
xnor U29925 (N_29925,N_25475,N_26238);
and U29926 (N_29926,N_25563,N_26725);
or U29927 (N_29927,N_26724,N_25055);
nor U29928 (N_29928,N_25720,N_25779);
nor U29929 (N_29929,N_25370,N_25634);
nand U29930 (N_29930,N_25539,N_25001);
or U29931 (N_29931,N_25667,N_25017);
nor U29932 (N_29932,N_27481,N_27052);
or U29933 (N_29933,N_25480,N_26972);
or U29934 (N_29934,N_25387,N_26506);
or U29935 (N_29935,N_27405,N_26261);
or U29936 (N_29936,N_25505,N_25951);
and U29937 (N_29937,N_26601,N_26948);
nand U29938 (N_29938,N_26384,N_27217);
and U29939 (N_29939,N_25484,N_26325);
or U29940 (N_29940,N_25406,N_25529);
xor U29941 (N_29941,N_25820,N_26316);
xor U29942 (N_29942,N_26886,N_27242);
xnor U29943 (N_29943,N_26025,N_26587);
nand U29944 (N_29944,N_27129,N_25903);
xor U29945 (N_29945,N_25899,N_26952);
nor U29946 (N_29946,N_26500,N_25477);
and U29947 (N_29947,N_25623,N_26916);
nand U29948 (N_29948,N_26259,N_25360);
and U29949 (N_29949,N_27216,N_27069);
nand U29950 (N_29950,N_26004,N_26394);
xor U29951 (N_29951,N_26972,N_25288);
nand U29952 (N_29952,N_25509,N_25867);
nand U29953 (N_29953,N_25762,N_25587);
or U29954 (N_29954,N_25275,N_26710);
or U29955 (N_29955,N_26466,N_25708);
xor U29956 (N_29956,N_27317,N_25870);
nor U29957 (N_29957,N_27185,N_26476);
and U29958 (N_29958,N_25635,N_26162);
or U29959 (N_29959,N_25023,N_25707);
xnor U29960 (N_29960,N_27136,N_26701);
nand U29961 (N_29961,N_25365,N_27202);
or U29962 (N_29962,N_26850,N_25604);
xor U29963 (N_29963,N_25875,N_25996);
or U29964 (N_29964,N_25302,N_25466);
nor U29965 (N_29965,N_25066,N_26705);
or U29966 (N_29966,N_26328,N_25950);
nor U29967 (N_29967,N_26697,N_26400);
or U29968 (N_29968,N_27159,N_25468);
nor U29969 (N_29969,N_25158,N_25913);
and U29970 (N_29970,N_27384,N_26519);
xnor U29971 (N_29971,N_26613,N_25243);
nand U29972 (N_29972,N_26564,N_26020);
nand U29973 (N_29973,N_26081,N_26738);
nand U29974 (N_29974,N_25610,N_25772);
and U29975 (N_29975,N_27437,N_26780);
nor U29976 (N_29976,N_26177,N_26890);
or U29977 (N_29977,N_25498,N_25790);
and U29978 (N_29978,N_25122,N_26590);
xnor U29979 (N_29979,N_26521,N_26269);
nor U29980 (N_29980,N_27221,N_27084);
nor U29981 (N_29981,N_26774,N_26348);
xnor U29982 (N_29982,N_25289,N_26734);
nor U29983 (N_29983,N_25756,N_25538);
and U29984 (N_29984,N_26427,N_27352);
and U29985 (N_29985,N_26223,N_25645);
or U29986 (N_29986,N_25133,N_26630);
and U29987 (N_29987,N_25373,N_25284);
or U29988 (N_29988,N_27231,N_26498);
nor U29989 (N_29989,N_25344,N_26852);
nor U29990 (N_29990,N_26916,N_26874);
xnor U29991 (N_29991,N_25695,N_26535);
xnor U29992 (N_29992,N_27106,N_25557);
nand U29993 (N_29993,N_27140,N_25862);
or U29994 (N_29994,N_25836,N_25179);
xor U29995 (N_29995,N_25997,N_26004);
or U29996 (N_29996,N_26882,N_26287);
and U29997 (N_29997,N_26598,N_26280);
or U29998 (N_29998,N_27498,N_26229);
nand U29999 (N_29999,N_26482,N_25028);
and U30000 (N_30000,N_28685,N_28303);
or U30001 (N_30001,N_29218,N_27708);
xnor U30002 (N_30002,N_29199,N_29651);
nor U30003 (N_30003,N_28390,N_28910);
or U30004 (N_30004,N_29934,N_28863);
or U30005 (N_30005,N_29588,N_28294);
and U30006 (N_30006,N_28393,N_27951);
or U30007 (N_30007,N_27666,N_28669);
xor U30008 (N_30008,N_29424,N_28712);
nand U30009 (N_30009,N_29669,N_28679);
and U30010 (N_30010,N_28804,N_28717);
and U30011 (N_30011,N_27880,N_29341);
or U30012 (N_30012,N_28167,N_27603);
nor U30013 (N_30013,N_28774,N_28029);
or U30014 (N_30014,N_28553,N_28620);
and U30015 (N_30015,N_28784,N_29886);
nor U30016 (N_30016,N_28858,N_28698);
and U30017 (N_30017,N_28762,N_28495);
xor U30018 (N_30018,N_29155,N_27914);
and U30019 (N_30019,N_28246,N_29332);
nand U30020 (N_30020,N_28596,N_28231);
or U30021 (N_30021,N_29164,N_29791);
nand U30022 (N_30022,N_28782,N_28444);
nand U30023 (N_30023,N_29027,N_29132);
nand U30024 (N_30024,N_28342,N_28375);
or U30025 (N_30025,N_28697,N_29339);
nor U30026 (N_30026,N_27521,N_29510);
nor U30027 (N_30027,N_28832,N_29709);
xor U30028 (N_30028,N_29862,N_29197);
nor U30029 (N_30029,N_29222,N_29097);
and U30030 (N_30030,N_28986,N_28194);
nand U30031 (N_30031,N_29698,N_28592);
nand U30032 (N_30032,N_28451,N_28569);
or U30033 (N_30033,N_29327,N_27778);
or U30034 (N_30034,N_27531,N_28790);
or U30035 (N_30035,N_28502,N_28023);
nor U30036 (N_30036,N_27511,N_29973);
nor U30037 (N_30037,N_28976,N_29177);
and U30038 (N_30038,N_29106,N_28438);
nor U30039 (N_30039,N_28630,N_29090);
or U30040 (N_30040,N_29035,N_28766);
xnor U30041 (N_30041,N_28270,N_28966);
nand U30042 (N_30042,N_28183,N_27660);
and U30043 (N_30043,N_28346,N_29885);
and U30044 (N_30044,N_28394,N_27824);
or U30045 (N_30045,N_28551,N_29751);
or U30046 (N_30046,N_29874,N_29501);
nor U30047 (N_30047,N_27990,N_29154);
nor U30048 (N_30048,N_28733,N_29546);
and U30049 (N_30049,N_29084,N_29869);
nand U30050 (N_30050,N_29320,N_29729);
nand U30051 (N_30051,N_29270,N_29919);
and U30052 (N_30052,N_29716,N_29948);
nand U30053 (N_30053,N_28958,N_28961);
xor U30054 (N_30054,N_28111,N_29153);
xor U30055 (N_30055,N_29717,N_28508);
and U30056 (N_30056,N_29061,N_29721);
nor U30057 (N_30057,N_28900,N_29640);
nand U30058 (N_30058,N_29771,N_28771);
and U30059 (N_30059,N_29151,N_29792);
xnor U30060 (N_30060,N_29010,N_29219);
or U30061 (N_30061,N_28476,N_29932);
nor U30062 (N_30062,N_29003,N_28157);
nor U30063 (N_30063,N_27535,N_28973);
nor U30064 (N_30064,N_29605,N_29582);
and U30065 (N_30065,N_28283,N_28469);
and U30066 (N_30066,N_28038,N_28730);
nor U30067 (N_30067,N_27758,N_29690);
nand U30068 (N_30068,N_29921,N_29295);
xor U30069 (N_30069,N_29333,N_28302);
xor U30070 (N_30070,N_29268,N_29530);
nand U30071 (N_30071,N_28586,N_28646);
nor U30072 (N_30072,N_29607,N_29784);
or U30073 (N_30073,N_29685,N_29355);
or U30074 (N_30074,N_29023,N_29451);
nand U30075 (N_30075,N_28185,N_27950);
nor U30076 (N_30076,N_29054,N_28627);
and U30077 (N_30077,N_28033,N_29654);
or U30078 (N_30078,N_29529,N_28887);
xnor U30079 (N_30079,N_28664,N_29827);
and U30080 (N_30080,N_27887,N_29009);
nor U30081 (N_30081,N_29042,N_29947);
or U30082 (N_30082,N_28844,N_28396);
and U30083 (N_30083,N_28625,N_27957);
nor U30084 (N_30084,N_29311,N_28843);
nor U30085 (N_30085,N_29748,N_28888);
xnor U30086 (N_30086,N_27934,N_29787);
nand U30087 (N_30087,N_28097,N_27811);
xor U30088 (N_30088,N_28120,N_28427);
nand U30089 (N_30089,N_28192,N_28942);
xnor U30090 (N_30090,N_27828,N_28074);
nor U30091 (N_30091,N_29229,N_29838);
or U30092 (N_30092,N_29481,N_28372);
nand U30093 (N_30093,N_29941,N_28387);
xnor U30094 (N_30094,N_29062,N_28607);
nand U30095 (N_30095,N_29294,N_29898);
nor U30096 (N_30096,N_27840,N_29692);
nor U30097 (N_30097,N_28518,N_28603);
nor U30098 (N_30098,N_27772,N_28773);
nor U30099 (N_30099,N_28959,N_27919);
nor U30100 (N_30100,N_29920,N_28795);
and U30101 (N_30101,N_29292,N_29200);
nor U30102 (N_30102,N_29979,N_28359);
nor U30103 (N_30103,N_28447,N_28078);
and U30104 (N_30104,N_29052,N_27541);
and U30105 (N_30105,N_28741,N_29191);
or U30106 (N_30106,N_27800,N_27876);
and U30107 (N_30107,N_27564,N_29967);
nand U30108 (N_30108,N_27598,N_29499);
nand U30109 (N_30109,N_28886,N_28904);
and U30110 (N_30110,N_28535,N_27810);
nand U30111 (N_30111,N_28936,N_27547);
nand U30112 (N_30112,N_27799,N_28054);
and U30113 (N_30113,N_28533,N_29823);
and U30114 (N_30114,N_28373,N_28732);
nand U30115 (N_30115,N_29150,N_29893);
or U30116 (N_30116,N_29524,N_29812);
nand U30117 (N_30117,N_29756,N_29083);
nor U30118 (N_30118,N_28457,N_29868);
or U30119 (N_30119,N_28780,N_28017);
and U30120 (N_30120,N_29627,N_29395);
and U30121 (N_30121,N_27915,N_28590);
xnor U30122 (N_30122,N_28031,N_29015);
xor U30123 (N_30123,N_29835,N_27871);
and U30124 (N_30124,N_29033,N_27529);
and U30125 (N_30125,N_29282,N_29336);
nand U30126 (N_30126,N_29039,N_29321);
or U30127 (N_30127,N_29840,N_27899);
and U30128 (N_30128,N_29082,N_28446);
or U30129 (N_30129,N_29537,N_28005);
nand U30130 (N_30130,N_28001,N_29381);
or U30131 (N_30131,N_28172,N_28995);
or U30132 (N_30132,N_28550,N_29492);
nor U30133 (N_30133,N_28713,N_29673);
and U30134 (N_30134,N_29970,N_29094);
and U30135 (N_30135,N_29727,N_29689);
and U30136 (N_30136,N_28785,N_28814);
nor U30137 (N_30137,N_28140,N_28536);
or U30138 (N_30138,N_27684,N_27570);
and U30139 (N_30139,N_28460,N_27993);
and U30140 (N_30140,N_29017,N_28361);
and U30141 (N_30141,N_27581,N_27754);
xnor U30142 (N_30142,N_28520,N_29450);
and U30143 (N_30143,N_29620,N_29731);
xnor U30144 (N_30144,N_28775,N_28134);
nand U30145 (N_30145,N_29517,N_28663);
nor U30146 (N_30146,N_28441,N_29079);
or U30147 (N_30147,N_28268,N_29794);
and U30148 (N_30148,N_27734,N_29684);
xnor U30149 (N_30149,N_29750,N_28133);
xor U30150 (N_30150,N_27788,N_28840);
nor U30151 (N_30151,N_29484,N_28874);
or U30152 (N_30152,N_28316,N_27943);
nand U30153 (N_30153,N_27738,N_28211);
or U30154 (N_30154,N_28847,N_27677);
nand U30155 (N_30155,N_28295,N_29190);
nor U30156 (N_30156,N_29906,N_29954);
nor U30157 (N_30157,N_29531,N_29486);
xor U30158 (N_30158,N_29045,N_29390);
nor U30159 (N_30159,N_27673,N_27700);
nor U30160 (N_30160,N_29589,N_27662);
and U30161 (N_30161,N_29819,N_29148);
nand U30162 (N_30162,N_29647,N_28560);
nand U30163 (N_30163,N_27869,N_27675);
or U30164 (N_30164,N_29785,N_28030);
nand U30165 (N_30165,N_28352,N_27544);
or U30166 (N_30166,N_29859,N_28252);
and U30167 (N_30167,N_28816,N_29186);
nor U30168 (N_30168,N_28368,N_29158);
nand U30169 (N_30169,N_28424,N_29918);
nand U30170 (N_30170,N_29245,N_28251);
and U30171 (N_30171,N_28941,N_28952);
nand U30172 (N_30172,N_28265,N_28682);
and U30173 (N_30173,N_28481,N_28350);
nor U30174 (N_30174,N_29686,N_28062);
nor U30175 (N_30175,N_28839,N_29714);
and U30176 (N_30176,N_27966,N_29317);
xnor U30177 (N_30177,N_29236,N_29584);
or U30178 (N_30178,N_29060,N_28641);
xor U30179 (N_30179,N_27906,N_28921);
and U30180 (N_30180,N_28275,N_27510);
nand U30181 (N_30181,N_29183,N_29497);
xor U30182 (N_30182,N_28081,N_28637);
or U30183 (N_30183,N_27515,N_29765);
nor U30184 (N_30184,N_29801,N_29570);
xnor U30185 (N_30185,N_27932,N_27792);
nor U30186 (N_30186,N_29305,N_27605);
xnor U30187 (N_30187,N_28391,N_27972);
and U30188 (N_30188,N_28738,N_28435);
xnor U30189 (N_30189,N_29961,N_29826);
xnor U30190 (N_30190,N_28497,N_27536);
nand U30191 (N_30191,N_28875,N_29952);
or U30192 (N_30192,N_28528,N_27837);
nand U30193 (N_30193,N_27711,N_29007);
nor U30194 (N_30194,N_29867,N_29900);
nand U30195 (N_30195,N_27577,N_28517);
and U30196 (N_30196,N_29697,N_27834);
or U30197 (N_30197,N_29758,N_28201);
or U30198 (N_30198,N_28594,N_29048);
xnor U30199 (N_30199,N_29828,N_29703);
and U30200 (N_30200,N_28199,N_29202);
xnor U30201 (N_30201,N_27981,N_27558);
nor U30202 (N_30202,N_28515,N_29005);
nand U30203 (N_30203,N_27879,N_28675);
nor U30204 (N_30204,N_27682,N_29230);
nand U30205 (N_30205,N_29943,N_27822);
nor U30206 (N_30206,N_28753,N_29092);
nand U30207 (N_30207,N_28512,N_29457);
xnor U30208 (N_30208,N_27670,N_29897);
nor U30209 (N_30209,N_28004,N_28020);
or U30210 (N_30210,N_29024,N_27881);
nand U30211 (N_30211,N_28636,N_29085);
xor U30212 (N_30212,N_28107,N_28112);
or U30213 (N_30213,N_29944,N_29553);
nand U30214 (N_30214,N_29960,N_29880);
nand U30215 (N_30215,N_29656,N_29460);
xor U30216 (N_30216,N_29632,N_28127);
and U30217 (N_30217,N_28543,N_28108);
and U30218 (N_30218,N_28170,N_29798);
or U30219 (N_30219,N_29019,N_28947);
and U30220 (N_30220,N_29873,N_29340);
or U30221 (N_30221,N_27593,N_28657);
xnor U30222 (N_30222,N_29187,N_29345);
and U30223 (N_30223,N_29400,N_27953);
nand U30224 (N_30224,N_29300,N_28604);
nand U30225 (N_30225,N_29490,N_28818);
xor U30226 (N_30226,N_29662,N_29608);
nand U30227 (N_30227,N_29876,N_28046);
xor U30228 (N_30228,N_29149,N_29385);
xnor U30229 (N_30229,N_29398,N_28779);
and U30230 (N_30230,N_29845,N_27999);
xnor U30231 (N_30231,N_28949,N_28349);
and U30232 (N_30232,N_28667,N_29806);
nor U30233 (N_30233,N_29763,N_27744);
and U30234 (N_30234,N_27980,N_29969);
nor U30235 (N_30235,N_29797,N_28969);
or U30236 (N_30236,N_27528,N_29382);
and U30237 (N_30237,N_27769,N_29215);
and U30238 (N_30238,N_27729,N_27585);
xor U30239 (N_30239,N_28466,N_29870);
xor U30240 (N_30240,N_27557,N_27912);
or U30241 (N_30241,N_27829,N_28545);
and U30242 (N_30242,N_28115,N_28129);
nor U30243 (N_30243,N_29810,N_29515);
xor U30244 (N_30244,N_27893,N_29166);
or U30245 (N_30245,N_29234,N_29986);
nand U30246 (N_30246,N_29313,N_29682);
nand U30247 (N_30247,N_29691,N_28661);
and U30248 (N_30248,N_28420,N_28212);
and U30249 (N_30249,N_28742,N_29380);
xnor U30250 (N_30250,N_29718,N_27783);
and U30251 (N_30251,N_29958,N_29988);
and U30252 (N_30252,N_28516,N_29905);
and U30253 (N_30253,N_29491,N_27731);
nor U30254 (N_30254,N_29281,N_29246);
nor U30255 (N_30255,N_28018,N_29427);
nor U30256 (N_30256,N_28452,N_28026);
nand U30257 (N_30257,N_29091,N_28002);
xor U30258 (N_30258,N_29115,N_28015);
or U30259 (N_30259,N_28873,N_28383);
and U30260 (N_30260,N_28866,N_29034);
nand U30261 (N_30261,N_28056,N_27562);
or U30262 (N_30262,N_29306,N_28221);
xnor U30263 (N_30263,N_27742,N_28422);
and U30264 (N_30264,N_28997,N_27533);
nand U30265 (N_30265,N_27693,N_28255);
or U30266 (N_30266,N_28826,N_28812);
and U30267 (N_30267,N_29285,N_27833);
or U30268 (N_30268,N_29800,N_29001);
nand U30269 (N_30269,N_28808,N_27813);
nand U30270 (N_30270,N_28357,N_28204);
and U30271 (N_30271,N_29393,N_29705);
nand U30272 (N_30272,N_29417,N_28378);
nor U30273 (N_30273,N_28721,N_28800);
xor U30274 (N_30274,N_29263,N_29216);
nor U30275 (N_30275,N_28531,N_27672);
xor U30276 (N_30276,N_27534,N_28392);
nor U30277 (N_30277,N_27955,N_28198);
and U30278 (N_30278,N_29680,N_29272);
xor U30279 (N_30279,N_28960,N_28648);
or U30280 (N_30280,N_29111,N_28370);
nand U30281 (N_30281,N_29414,N_29770);
nor U30282 (N_30282,N_27940,N_29470);
xnor U30283 (N_30283,N_28925,N_27601);
xor U30284 (N_30284,N_28867,N_28504);
nor U30285 (N_30285,N_28834,N_29804);
xor U30286 (N_30286,N_28035,N_29167);
and U30287 (N_30287,N_27992,N_28000);
nand U30288 (N_30288,N_27860,N_28178);
nand U30289 (N_30289,N_29799,N_29103);
and U30290 (N_30290,N_28609,N_29520);
or U30291 (N_30291,N_28567,N_29937);
and U30292 (N_30292,N_29707,N_29518);
or U30293 (N_30293,N_27795,N_29221);
or U30294 (N_30294,N_29639,N_28311);
or U30295 (N_30295,N_28967,N_28868);
or U30296 (N_30296,N_28527,N_29715);
nor U30297 (N_30297,N_29182,N_29983);
or U30298 (N_30298,N_27948,N_29883);
and U30299 (N_30299,N_29675,N_29775);
xor U30300 (N_30300,N_27973,N_29243);
or U30301 (N_30301,N_29645,N_29681);
nor U30302 (N_30302,N_28439,N_29976);
nand U30303 (N_30303,N_27559,N_28174);
or U30304 (N_30304,N_29593,N_28987);
and U30305 (N_30305,N_28701,N_29927);
or U30306 (N_30306,N_28499,N_27513);
nor U30307 (N_30307,N_29899,N_29946);
and U30308 (N_30308,N_27835,N_27851);
nor U30309 (N_30309,N_29047,N_29556);
nand U30310 (N_30310,N_28981,N_28171);
xor U30311 (N_30311,N_28723,N_28436);
nor U30312 (N_30312,N_29829,N_27884);
nor U30313 (N_30313,N_28579,N_28837);
xnor U30314 (N_30314,N_28506,N_28964);
xnor U30315 (N_30315,N_28990,N_28253);
xor U30316 (N_30316,N_28631,N_27669);
nor U30317 (N_30317,N_27604,N_28468);
nor U30318 (N_30318,N_28786,N_27985);
xnor U30319 (N_30319,N_29957,N_29852);
nor U30320 (N_30320,N_27571,N_29494);
nand U30321 (N_30321,N_28909,N_27781);
and U30322 (N_30322,N_28092,N_29722);
and U30323 (N_30323,N_28623,N_28621);
xnor U30324 (N_30324,N_29642,N_28864);
or U30325 (N_30325,N_28314,N_27929);
and U30326 (N_30326,N_28297,N_28122);
nor U30327 (N_30327,N_28937,N_29472);
nand U30328 (N_30328,N_28678,N_27964);
xor U30329 (N_30329,N_27956,N_29790);
nand U30330 (N_30330,N_29614,N_27615);
and U30331 (N_30331,N_29374,N_29296);
and U30332 (N_30332,N_28582,N_29248);
nor U30333 (N_30333,N_29950,N_27576);
xor U30334 (N_30334,N_29901,N_29863);
and U30335 (N_30335,N_28069,N_28856);
xnor U30336 (N_30336,N_29617,N_28872);
nand U30337 (N_30337,N_27905,N_29028);
or U30338 (N_30338,N_28155,N_28066);
nand U30339 (N_30339,N_29534,N_27629);
xor U30340 (N_30340,N_27875,N_28794);
xor U30341 (N_30341,N_29399,N_28606);
xor U30342 (N_30342,N_28068,N_28570);
xnor U30343 (N_30343,N_29657,N_29217);
and U30344 (N_30344,N_29601,N_27983);
and U30345 (N_30345,N_27674,N_29309);
and U30346 (N_30346,N_29433,N_27760);
or U30347 (N_30347,N_27686,N_29541);
and U30348 (N_30348,N_27640,N_28432);
nor U30349 (N_30349,N_28400,N_29014);
and U30350 (N_30350,N_28768,N_28058);
or U30351 (N_30351,N_27969,N_28827);
and U30352 (N_30352,N_29987,N_27736);
or U30353 (N_30353,N_28259,N_27987);
nor U30354 (N_30354,N_27988,N_29755);
xnor U30355 (N_30355,N_28789,N_29206);
nand U30356 (N_30356,N_28974,N_28511);
nor U30357 (N_30357,N_29360,N_29644);
nor U30358 (N_30358,N_29471,N_28256);
nor U30359 (N_30359,N_28923,N_28666);
nor U30360 (N_30360,N_27602,N_27959);
xor U30361 (N_30361,N_28707,N_27546);
and U30362 (N_30362,N_29358,N_28492);
nor U30363 (N_30363,N_29887,N_28809);
nand U30364 (N_30364,N_28100,N_29324);
and U30365 (N_30365,N_27804,N_27763);
xnor U30366 (N_30366,N_28770,N_29310);
and U30367 (N_30367,N_29051,N_28980);
nand U30368 (N_30368,N_29384,N_28010);
or U30369 (N_30369,N_29116,N_29031);
or U30370 (N_30370,N_29891,N_28117);
nor U30371 (N_30371,N_28474,N_27607);
nor U30372 (N_30372,N_27637,N_28239);
and U30373 (N_30373,N_28578,N_29574);
and U30374 (N_30374,N_29018,N_29426);
nor U30375 (N_30375,N_27895,N_27962);
xor U30376 (N_30376,N_29581,N_28224);
nor U30377 (N_30377,N_28658,N_28250);
xnor U30378 (N_30378,N_28719,N_27505);
and U30379 (N_30379,N_28276,N_28477);
or U30380 (N_30380,N_29179,N_29477);
nor U30381 (N_30381,N_27500,N_29674);
and U30382 (N_30382,N_28273,N_28860);
xnor U30383 (N_30383,N_27916,N_28815);
nand U30384 (N_30384,N_28805,N_29578);
and U30385 (N_30385,N_29625,N_27963);
xnor U30386 (N_30386,N_28347,N_29098);
xor U30387 (N_30387,N_28105,N_28077);
and U30388 (N_30388,N_29423,N_28534);
or U30389 (N_30389,N_28931,N_29889);
xor U30390 (N_30390,N_28589,N_28095);
xor U30391 (N_30391,N_28668,N_28954);
nand U30392 (N_30392,N_29361,N_28616);
xor U30393 (N_30393,N_27856,N_29169);
nor U30394 (N_30394,N_29908,N_27801);
or U30395 (N_30395,N_27995,N_29378);
and U30396 (N_30396,N_27648,N_27768);
and U30397 (N_30397,N_29249,N_29815);
xor U30398 (N_30398,N_29805,N_29220);
nor U30399 (N_30399,N_29498,N_29156);
nor U30400 (N_30400,N_28982,N_28047);
nand U30401 (N_30401,N_29878,N_28067);
xnor U30402 (N_30402,N_27970,N_29650);
nor U30403 (N_30403,N_27654,N_27589);
xor U30404 (N_30404,N_28992,N_28085);
xnor U30405 (N_30405,N_28680,N_28890);
and U30406 (N_30406,N_28043,N_27540);
xnor U30407 (N_30407,N_29628,N_28912);
or U30408 (N_30408,N_29247,N_27718);
or U30409 (N_30409,N_27945,N_29576);
nor U30410 (N_30410,N_27762,N_29344);
or U30411 (N_30411,N_29388,N_29701);
nand U30412 (N_30412,N_29571,N_28341);
or U30413 (N_30413,N_27892,N_28524);
and U30414 (N_30414,N_28191,N_27658);
nand U30415 (N_30415,N_29401,N_29185);
or U30416 (N_30416,N_27647,N_28684);
and U30417 (N_30417,N_28164,N_29549);
or U30418 (N_30418,N_28162,N_28089);
and U30419 (N_30419,N_29602,N_28521);
nor U30420 (N_30420,N_27657,N_29495);
xor U30421 (N_30421,N_27703,N_29736);
or U30422 (N_30422,N_29203,N_28583);
nand U30423 (N_30423,N_27991,N_28822);
or U30424 (N_30424,N_28381,N_28453);
nand U30425 (N_30425,N_29538,N_29746);
or U30426 (N_30426,N_29449,N_28626);
and U30427 (N_30427,N_29274,N_29851);
nand U30428 (N_30428,N_28345,N_29174);
nor U30429 (N_30429,N_28414,N_28993);
xor U30430 (N_30430,N_27918,N_28286);
or U30431 (N_30431,N_29866,N_28687);
nor U30432 (N_30432,N_28425,N_29997);
nand U30433 (N_30433,N_27507,N_29540);
nand U30434 (N_30434,N_29466,N_29843);
xnor U30435 (N_30435,N_28801,N_28406);
xnor U30436 (N_30436,N_29567,N_28752);
or U30437 (N_30437,N_29262,N_27808);
and U30438 (N_30438,N_27650,N_29102);
xor U30439 (N_30439,N_27638,N_29440);
nor U30440 (N_30440,N_28725,N_29591);
xor U30441 (N_30441,N_28737,N_28202);
nor U30442 (N_30442,N_27831,N_29404);
nand U30443 (N_30443,N_27526,N_29809);
or U30444 (N_30444,N_27847,N_29741);
nand U30445 (N_30445,N_29532,N_27538);
or U30446 (N_30446,N_28149,N_29368);
and U30447 (N_30447,N_29949,N_29637);
nand U30448 (N_30448,N_27770,N_29613);
nor U30449 (N_30449,N_28735,N_29483);
and U30450 (N_30450,N_29778,N_27809);
nor U30451 (N_30451,N_28576,N_28187);
and U30452 (N_30452,N_27921,N_27941);
nand U30453 (N_30453,N_29121,N_28799);
xnor U30454 (N_30454,N_29788,N_29560);
nand U30455 (N_30455,N_28756,N_27679);
xnor U30456 (N_30456,N_29485,N_29269);
xor U30457 (N_30457,N_27774,N_29459);
xnor U30458 (N_30458,N_29688,N_29419);
nand U30459 (N_30459,N_27787,N_27883);
nor U30460 (N_30460,N_29043,N_28615);
nor U30461 (N_30461,N_27873,N_28369);
nor U30462 (N_30462,N_28291,N_29022);
and U30463 (N_30463,N_27803,N_27572);
nand U30464 (N_30464,N_29383,N_29142);
nor U30465 (N_30465,N_27539,N_29415);
and U30466 (N_30466,N_28984,N_29562);
nand U30467 (N_30467,N_29635,N_28242);
nor U30468 (N_30468,N_28880,N_28728);
and U30469 (N_30469,N_29670,N_28597);
xor U30470 (N_30470,N_27683,N_27690);
nor U30471 (N_30471,N_29139,N_28977);
nor U30472 (N_30472,N_28704,N_28983);
nand U30473 (N_30473,N_27639,N_29535);
nor U30474 (N_30474,N_27939,N_28632);
or U30475 (N_30475,N_29067,N_28364);
nand U30476 (N_30476,N_28036,N_29448);
and U30477 (N_30477,N_28628,N_29016);
nand U30478 (N_30478,N_27930,N_29533);
and U30479 (N_30479,N_28945,N_29038);
xor U30480 (N_30480,N_27642,N_28267);
or U30481 (N_30481,N_28859,N_29816);
nand U30482 (N_30482,N_28177,N_29453);
and U30483 (N_30483,N_29025,N_29157);
or U30484 (N_30484,N_27551,N_27689);
nor U30485 (N_30485,N_29712,N_28153);
nor U30486 (N_30486,N_28146,N_28587);
or U30487 (N_30487,N_29693,N_29523);
or U30488 (N_30488,N_28736,N_28978);
and U30489 (N_30489,N_28417,N_29231);
or U30490 (N_30490,N_28009,N_27550);
nand U30491 (N_30491,N_28467,N_28410);
or U30492 (N_30492,N_28322,N_28113);
and U30493 (N_30493,N_27798,N_27761);
and U30494 (N_30494,N_27877,N_29505);
nand U30495 (N_30495,N_29265,N_29273);
or U30496 (N_30496,N_29180,N_28841);
nor U30497 (N_30497,N_29211,N_29053);
nand U30498 (N_30498,N_29487,N_27900);
nor U30499 (N_30499,N_28710,N_29322);
xnor U30500 (N_30500,N_28395,N_29879);
nor U30501 (N_30501,N_29547,N_29235);
nor U30502 (N_30502,N_28374,N_29996);
nand U30503 (N_30503,N_28878,N_28338);
nand U30504 (N_30504,N_28633,N_29212);
nand U30505 (N_30505,N_29369,N_29343);
xnor U30506 (N_30506,N_28091,N_29604);
or U30507 (N_30507,N_28884,N_29832);
or U30508 (N_30508,N_28064,N_27909);
nand U30509 (N_30509,N_27764,N_27709);
nand U30510 (N_30510,N_29239,N_27782);
and U30511 (N_30511,N_28473,N_28988);
or U30512 (N_30512,N_28883,N_28028);
xnor U30513 (N_30513,N_28102,N_29990);
nor U30514 (N_30514,N_28509,N_27961);
nand U30515 (N_30515,N_29679,N_29521);
nand U30516 (N_30516,N_29720,N_28561);
nand U30517 (N_30517,N_28998,N_27989);
or U30518 (N_30518,N_28116,N_28434);
xor U30519 (N_30519,N_27671,N_28057);
nor U30520 (N_30520,N_27617,N_29410);
nand U30521 (N_30521,N_29474,N_29008);
nand U30522 (N_30522,N_28693,N_27854);
nand U30523 (N_30523,N_29392,N_29351);
or U30524 (N_30524,N_29783,N_29732);
nand U30525 (N_30525,N_27848,N_27676);
nor U30526 (N_30526,N_28299,N_28911);
or U30527 (N_30527,N_27859,N_27780);
nand U30528 (N_30528,N_28104,N_27777);
nand U30529 (N_30529,N_28836,N_27942);
and U30530 (N_30530,N_29432,N_29334);
or U30531 (N_30531,N_29096,N_28235);
nor U30532 (N_30532,N_27661,N_29730);
or U30533 (N_30533,N_29473,N_29551);
nor U30534 (N_30534,N_27832,N_28193);
xnor U30535 (N_30535,N_27815,N_28505);
nand U30536 (N_30536,N_27865,N_27858);
or U30537 (N_30537,N_27979,N_29726);
and U30538 (N_30538,N_29877,N_29633);
and U30539 (N_30539,N_29909,N_27894);
or U30540 (N_30540,N_27960,N_29413);
and U30541 (N_30541,N_28013,N_28924);
nor U30542 (N_30542,N_28156,N_28761);
xnor U30543 (N_30543,N_29093,N_29468);
nand U30544 (N_30544,N_27842,N_27624);
xnor U30545 (N_30545,N_27868,N_28940);
nor U30546 (N_30546,N_29989,N_28330);
xor U30547 (N_30547,N_29335,N_29205);
nor U30548 (N_30548,N_28871,N_29134);
xor U30549 (N_30549,N_29371,N_28082);
and U30550 (N_30550,N_29080,N_29125);
and U30551 (N_30551,N_29516,N_28879);
xor U30552 (N_30552,N_28650,N_27907);
nand U30553 (N_30553,N_28471,N_29938);
and U30554 (N_30554,N_29548,N_29740);
xnor U30555 (N_30555,N_28622,N_29437);
and U30556 (N_30556,N_28647,N_29331);
nor U30557 (N_30557,N_29575,N_29699);
and U30558 (N_30558,N_28042,N_29762);
or U30559 (N_30559,N_28584,N_28094);
or U30560 (N_30560,N_28173,N_28109);
xor U30561 (N_30561,N_29861,N_28429);
or U30562 (N_30562,N_27611,N_28334);
nor U30563 (N_30563,N_29464,N_28247);
or U30564 (N_30564,N_28228,N_28483);
nand U30565 (N_30565,N_28470,N_27628);
nor U30566 (N_30566,N_27751,N_27935);
or U30567 (N_30567,N_29713,N_28908);
and U30568 (N_30568,N_28580,N_29882);
nor U30569 (N_30569,N_28585,N_28963);
nand U30570 (N_30570,N_29733,N_29438);
nand U30571 (N_30571,N_29099,N_29475);
or U30572 (N_30572,N_29290,N_29389);
or U30573 (N_30573,N_27619,N_29255);
and U30574 (N_30574,N_29789,N_28554);
and U30575 (N_30575,N_27794,N_29708);
or U30576 (N_30576,N_28449,N_28306);
or U30577 (N_30577,N_27687,N_28611);
xor U30578 (N_30578,N_28006,N_29624);
nand U30579 (N_30579,N_27779,N_29597);
and U30580 (N_30580,N_28853,N_29021);
nor U30581 (N_30581,N_29696,N_28591);
and U30582 (N_30582,N_27791,N_29461);
or U30583 (N_30583,N_28220,N_29297);
nor U30584 (N_30584,N_27728,N_28662);
xnor U30585 (N_30585,N_29545,N_27635);
and U30586 (N_30586,N_28544,N_29455);
nand U30587 (N_30587,N_28731,N_29223);
nand U30588 (N_30588,N_28331,N_28744);
xor U30589 (N_30589,N_29244,N_27927);
or U30590 (N_30590,N_29133,N_29700);
nor U30591 (N_30591,N_29592,N_28141);
nand U30592 (N_30592,N_29159,N_28365);
xnor U30593 (N_30593,N_29586,N_28493);
nand U30594 (N_30594,N_27652,N_28323);
nand U30595 (N_30595,N_28180,N_28749);
nand U30596 (N_30596,N_28229,N_27733);
nor U30597 (N_30597,N_27775,N_28614);
nor U30598 (N_30598,N_28227,N_27819);
and U30599 (N_30599,N_28355,N_28261);
nand U30600 (N_30600,N_29163,N_27853);
nor U30601 (N_30601,N_27506,N_29621);
and U30602 (N_30602,N_27574,N_28135);
nand U30603 (N_30603,N_29172,N_28456);
and U30604 (N_30604,N_27706,N_27784);
nand U30605 (N_30605,N_29834,N_28161);
xnor U30606 (N_30606,N_29436,N_28613);
xor U30607 (N_30607,N_28796,N_27846);
nand U30608 (N_30608,N_28053,N_28217);
nor U30609 (N_30609,N_27741,N_28727);
xor U30610 (N_30610,N_29489,N_28817);
and U30611 (N_30611,N_28325,N_28049);
nor U30612 (N_30612,N_28807,N_29926);
nand U30613 (N_30613,N_28237,N_29841);
xor U30614 (N_30614,N_28672,N_28915);
and U30615 (N_30615,N_29041,N_28739);
xnor U30616 (N_30616,N_28927,N_29702);
xor U30617 (N_30617,N_27664,N_28708);
nand U30618 (N_30618,N_28895,N_28711);
xor U30619 (N_30619,N_28126,N_28139);
nand U30620 (N_30620,N_29888,N_28559);
xnor U30621 (N_30621,N_27917,N_28249);
nor U30622 (N_30622,N_27724,N_29507);
nor U30623 (N_30623,N_28696,N_27656);
nor U30624 (N_30624,N_28271,N_28500);
xor U30625 (N_30625,N_29020,N_28025);
or U30626 (N_30626,N_29232,N_29479);
and U30627 (N_30627,N_28781,N_29522);
and U30628 (N_30628,N_27659,N_28478);
nor U30629 (N_30629,N_28354,N_28213);
or U30630 (N_30630,N_28918,N_28019);
and U30631 (N_30631,N_28933,N_28443);
xor U30632 (N_30632,N_27857,N_29407);
nor U30633 (N_30633,N_28491,N_27591);
xnor U30634 (N_30634,N_29303,N_28210);
xor U30635 (N_30635,N_27502,N_28546);
or U30636 (N_30636,N_28957,N_28702);
xnor U30637 (N_30637,N_29373,N_27599);
and U30638 (N_30638,N_28463,N_27790);
or U30639 (N_30639,N_29059,N_29890);
nor U30640 (N_30640,N_28519,N_28296);
and U30641 (N_30641,N_28722,N_28548);
xnor U30642 (N_30642,N_29002,N_27924);
nor U30643 (N_30643,N_28479,N_29971);
xor U30644 (N_30644,N_29768,N_29653);
and U30645 (N_30645,N_27925,N_27923);
and U30646 (N_30646,N_28514,N_27785);
nand U30647 (N_30647,N_27882,N_28226);
and U30648 (N_30648,N_27606,N_29634);
nand U30649 (N_30649,N_28999,N_29744);
nand U30650 (N_30650,N_29661,N_28670);
and U30651 (N_30651,N_28542,N_29603);
or U30652 (N_30652,N_28450,N_27644);
nand U30653 (N_30653,N_28280,N_28200);
and U30654 (N_30654,N_27773,N_29075);
nand U30655 (N_30655,N_29469,N_28152);
nor U30656 (N_30656,N_28462,N_28892);
and U30657 (N_30657,N_28938,N_28219);
nor U30658 (N_30658,N_28747,N_27516);
xnor U30659 (N_30659,N_28052,N_29956);
and U30660 (N_30660,N_29536,N_28384);
or U30661 (N_30661,N_29101,N_29710);
nand U30662 (N_30662,N_29353,N_28539);
or U30663 (N_30663,N_29118,N_28709);
and U30664 (N_30664,N_28595,N_28040);
and U30665 (N_30665,N_28233,N_29526);
nand U30666 (N_30666,N_28760,N_28371);
nand U30667 (N_30667,N_29892,N_28379);
and U30668 (N_30668,N_27634,N_29108);
and U30669 (N_30669,N_27910,N_28179);
and U30670 (N_30670,N_28996,N_28944);
or U30671 (N_30671,N_29824,N_29396);
and U30672 (N_30672,N_29251,N_29254);
xor U30673 (N_30673,N_28158,N_29168);
nand U30674 (N_30674,N_29291,N_27821);
nand U30675 (N_30675,N_28652,N_29352);
nand U30676 (N_30676,N_28309,N_29319);
xnor U30677 (N_30677,N_27542,N_29519);
xnor U30678 (N_30678,N_28339,N_27549);
and U30679 (N_30679,N_28862,N_28985);
nand U30680 (N_30680,N_29853,N_28114);
and U30681 (N_30681,N_27863,N_28101);
nand U30682 (N_30682,N_27977,N_28412);
nand U30683 (N_30683,N_28336,N_28022);
nor U30684 (N_30684,N_28897,N_29995);
or U30685 (N_30685,N_27717,N_27530);
xor U30686 (N_30686,N_29482,N_27984);
or U30687 (N_30687,N_29564,N_27861);
or U30688 (N_30688,N_27627,N_27997);
and U30689 (N_30689,N_29114,N_29807);
xor U30690 (N_30690,N_29377,N_28605);
nor U30691 (N_30691,N_28189,N_27527);
nor U30692 (N_30692,N_27609,N_29391);
or U30693 (N_30693,N_29858,N_27563);
and U30694 (N_30694,N_28160,N_27730);
xor U30695 (N_30695,N_27749,N_28398);
xor U30696 (N_30696,N_27816,N_28304);
nand U30697 (N_30697,N_29257,N_29095);
nor U30698 (N_30698,N_27740,N_27771);
or U30699 (N_30699,N_28209,N_28310);
and U30700 (N_30700,N_29953,N_27600);
xor U30701 (N_30701,N_28490,N_28939);
nor U30702 (N_30702,N_28222,N_29616);
nor U30703 (N_30703,N_28651,N_29663);
nand U30704 (N_30704,N_27874,N_28367);
nand U30705 (N_30705,N_28644,N_28003);
xnor U30706 (N_30706,N_27975,N_28891);
or U30707 (N_30707,N_28260,N_27714);
and U30708 (N_30708,N_27805,N_28638);
and U30709 (N_30709,N_29942,N_28772);
nor U30710 (N_30710,N_28759,N_28136);
nor U30711 (N_30711,N_29648,N_28537);
or U30712 (N_30712,N_27838,N_29924);
nor U30713 (N_30713,N_29214,N_29316);
nor U30714 (N_30714,N_28917,N_29195);
or U30715 (N_30715,N_28070,N_28041);
xnor U30716 (N_30716,N_29283,N_29871);
and U30717 (N_30717,N_29176,N_28810);
xor U30718 (N_30718,N_29754,N_29933);
and U30719 (N_30719,N_29452,N_29817);
nand U30720 (N_30720,N_28351,N_28197);
and U30721 (N_30721,N_28175,N_29902);
and U30722 (N_30722,N_29078,N_28549);
nor U30723 (N_30723,N_29856,N_28324);
xnor U30724 (N_30724,N_28337,N_29359);
nor U30725 (N_30725,N_28571,N_28573);
and U30726 (N_30726,N_29488,N_28758);
nand U30727 (N_30727,N_29678,N_27612);
nand U30728 (N_30728,N_28547,N_28556);
or U30729 (N_30729,N_28566,N_29683);
nor U30730 (N_30730,N_28181,N_28743);
nand U30731 (N_30731,N_29318,N_29929);
or U30732 (N_30732,N_28979,N_29550);
xnor U30733 (N_30733,N_28919,N_27836);
nor U30734 (N_30734,N_28051,N_29350);
nor U30735 (N_30735,N_27789,N_29577);
and U30736 (N_30736,N_28382,N_29068);
nor U30737 (N_30737,N_28190,N_28437);
nor U30738 (N_30738,N_28465,N_28388);
nand U30739 (N_30739,N_27936,N_28558);
and U30740 (N_30740,N_28360,N_29162);
xnor U30741 (N_30741,N_29443,N_28842);
and U30742 (N_30742,N_28344,N_28014);
xnor U30743 (N_30743,N_29087,N_29641);
or U30744 (N_30744,N_29981,N_28928);
xnor U30745 (N_30745,N_28541,N_27586);
and U30746 (N_30746,N_28482,N_27726);
or U30747 (N_30747,N_27890,N_29839);
nand U30748 (N_30748,N_27755,N_28734);
and U30749 (N_30749,N_27501,N_27626);
nor U30750 (N_30750,N_28196,N_29963);
nand U30751 (N_30751,N_28034,N_29192);
nand U30752 (N_30752,N_29013,N_29552);
and U30753 (N_30753,N_28485,N_29672);
or U30754 (N_30754,N_27720,N_29743);
xor U30755 (N_30755,N_29594,N_29998);
or U30756 (N_30756,N_28865,N_28602);
nor U30757 (N_30757,N_28225,N_29004);
and U30758 (N_30758,N_29780,N_27552);
nor U30759 (N_30759,N_27610,N_27705);
or U30760 (N_30760,N_28905,N_28562);
or U30761 (N_30761,N_27996,N_27694);
or U30762 (N_30762,N_29814,N_29706);
and U30763 (N_30763,N_29425,N_29506);
and U30764 (N_30764,N_28948,N_27616);
xor U30765 (N_30765,N_29757,N_28048);
nor U30766 (N_30766,N_27503,N_28778);
nand U30767 (N_30767,N_29904,N_29420);
nor U30768 (N_30768,N_28575,N_29403);
nor U30769 (N_30769,N_29619,N_29609);
xor U30770 (N_30770,N_27696,N_28557);
xnor U30771 (N_30771,N_29781,N_28695);
xnor U30772 (N_30772,N_28169,N_28032);
xnor U30773 (N_30773,N_28935,N_28285);
and U30774 (N_30774,N_28729,N_29509);
or U30775 (N_30775,N_28098,N_29204);
or U30776 (N_30776,N_28532,N_29356);
nor U30777 (N_30777,N_28686,N_29910);
nor U30778 (N_30778,N_28660,N_28278);
and U30779 (N_30779,N_28823,N_27839);
nand U30780 (N_30780,N_29940,N_29749);
or U30781 (N_30781,N_28272,N_28289);
nor U30782 (N_30782,N_28968,N_28577);
nand U30783 (N_30783,N_28946,N_29962);
xor U30784 (N_30784,N_28838,N_29145);
nor U30785 (N_30785,N_29769,N_29583);
and U30786 (N_30786,N_29171,N_28764);
xnor U30787 (N_30787,N_28835,N_28423);
nor U30788 (N_30788,N_27757,N_28335);
and U30789 (N_30789,N_27812,N_29135);
nand U30790 (N_30790,N_28824,N_27888);
xor U30791 (N_30791,N_28206,N_29512);
xnor U30792 (N_30792,N_29630,N_27543);
and U30793 (N_30793,N_28943,N_28994);
or U30794 (N_30794,N_29568,N_27633);
nor U30795 (N_30795,N_29074,N_28218);
and U30796 (N_30796,N_29467,N_29070);
and U30797 (N_30797,N_29366,N_27807);
and U30798 (N_30798,N_27566,N_27707);
nand U30799 (N_30799,N_28458,N_28813);
or U30800 (N_30800,N_28060,N_29854);
and U30801 (N_30801,N_29966,N_29811);
and U30802 (N_30802,N_28154,N_28366);
nand U30803 (N_30803,N_28618,N_28718);
and U30804 (N_30804,N_29922,N_29855);
nand U30805 (N_30805,N_29513,N_27561);
nor U30806 (N_30806,N_29825,N_28525);
nor U30807 (N_30807,N_28953,N_27595);
xor U30808 (N_30808,N_28288,N_28319);
and U30809 (N_30809,N_29429,N_28881);
or U30810 (N_30810,N_29964,N_28498);
nor U30811 (N_30811,N_28008,N_29496);
xor U30812 (N_30812,N_27710,N_27965);
or U30813 (N_30813,N_28281,N_27665);
or U30814 (N_30814,N_29955,N_28232);
and U30815 (N_30815,N_27796,N_29271);
or U30816 (N_30816,N_28962,N_29446);
nand U30817 (N_30817,N_28176,N_27645);
nor U30818 (N_30818,N_27587,N_27596);
nand U30819 (N_30819,N_28405,N_28692);
nor U30820 (N_30820,N_29250,N_28746);
and U30821 (N_30821,N_28459,N_29782);
nor U30822 (N_30822,N_28145,N_28386);
and U30823 (N_30823,N_28700,N_28184);
nor U30824 (N_30824,N_28418,N_27568);
nor U30825 (N_30825,N_28182,N_28480);
and U30826 (N_30826,N_29747,N_28142);
nor U30827 (N_30827,N_29566,N_28861);
or U30828 (N_30828,N_29561,N_28248);
and U30829 (N_30829,N_28750,N_29822);
and U30830 (N_30830,N_29012,N_27509);
nand U30831 (N_30831,N_29599,N_29405);
or U30832 (N_30832,N_28494,N_29636);
nand U30833 (N_30833,N_29124,N_28849);
and U30834 (N_30834,N_29055,N_28326);
or U30835 (N_30835,N_29842,N_28243);
xnor U30836 (N_30836,N_27630,N_27986);
and U30837 (N_30837,N_29259,N_27841);
xor U30838 (N_30838,N_27667,N_29402);
and U30839 (N_30839,N_29409,N_29821);
xnor U30840 (N_30840,N_28629,N_29226);
nor U30841 (N_30841,N_28568,N_28610);
nor U30842 (N_30842,N_28971,N_29240);
or U30843 (N_30843,N_29127,N_27578);
nand U30844 (N_30844,N_29569,N_28244);
xnor U30845 (N_30845,N_27555,N_28072);
or U30846 (N_30846,N_28110,N_29764);
nor U30847 (N_30847,N_29864,N_27702);
nand U30848 (N_30848,N_28096,N_28472);
and U30849 (N_30849,N_28673,N_27750);
xnor U30850 (N_30850,N_28674,N_29965);
or U30851 (N_30851,N_28088,N_28932);
nor U30852 (N_30852,N_28788,N_29652);
or U30853 (N_30853,N_29069,N_28084);
or U30854 (N_30854,N_28307,N_28572);
nor U30855 (N_30855,N_27922,N_29130);
or U30856 (N_30856,N_27588,N_29113);
or U30857 (N_30857,N_29040,N_28266);
and U30858 (N_30858,N_28600,N_29884);
xor U30859 (N_30859,N_29073,N_27520);
nand U30860 (N_30860,N_29915,N_29144);
or U30861 (N_30861,N_29724,N_27793);
nor U30862 (N_30862,N_29930,N_27938);
and U30863 (N_30863,N_29895,N_28783);
or U30864 (N_30864,N_29974,N_29088);
or U30865 (N_30865,N_29178,N_29836);
xor U30866 (N_30866,N_28421,N_28234);
nor U30867 (N_30867,N_29931,N_29734);
nand U30868 (N_30868,N_29543,N_27937);
and U30869 (N_30869,N_29428,N_28131);
or U30870 (N_30870,N_29623,N_27631);
nor U30871 (N_30871,N_27817,N_29458);
nand U30872 (N_30872,N_28507,N_29928);
xnor U30873 (N_30873,N_29923,N_28598);
or U30874 (N_30874,N_28599,N_27753);
nand U30875 (N_30875,N_29147,N_28563);
nor U30876 (N_30876,N_28340,N_28123);
nor U30877 (N_30877,N_29107,N_27525);
nand U30878 (N_30878,N_29264,N_29201);
or U30879 (N_30879,N_29837,N_28413);
xnor U30880 (N_30880,N_29985,N_28287);
or U30881 (N_30881,N_28681,N_28059);
nand U30882 (N_30882,N_28777,N_27567);
and U30883 (N_30883,N_28564,N_27866);
nand U30884 (N_30884,N_29925,N_29911);
nand U30885 (N_30885,N_27721,N_28430);
nand U30886 (N_30886,N_28151,N_28903);
and U30887 (N_30887,N_28751,N_29525);
or U30888 (N_30888,N_27830,N_28230);
and U30889 (N_30889,N_29978,N_28645);
or U30890 (N_30890,N_29299,N_28588);
xnor U30891 (N_30891,N_29735,N_28241);
or U30892 (N_30892,N_29329,N_28027);
nor U30893 (N_30893,N_28130,N_27620);
or U30894 (N_30894,N_28207,N_29659);
nor U30895 (N_30895,N_28044,N_27594);
nor U30896 (N_30896,N_27974,N_28501);
nand U30897 (N_30897,N_27537,N_29129);
xor U30898 (N_30898,N_28454,N_27766);
nor U30899 (N_30899,N_28755,N_28806);
or U30900 (N_30900,N_29454,N_27867);
or U30901 (N_30901,N_29480,N_28828);
nand U30902 (N_30902,N_27523,N_29646);
or U30903 (N_30903,N_28343,N_28522);
nor U30904 (N_30904,N_29872,N_29314);
and U30905 (N_30905,N_28138,N_28975);
xnor U30906 (N_30906,N_27814,N_28461);
and U30907 (N_30907,N_29704,N_28885);
or U30908 (N_30908,N_28061,N_28312);
xor U30909 (N_30909,N_28820,N_28540);
or U30910 (N_30910,N_29237,N_28411);
xor U30911 (N_30911,N_28757,N_27855);
xnor U30912 (N_30912,N_28318,N_28292);
or U30913 (N_30913,N_27681,N_28705);
nor U30914 (N_30914,N_27712,N_27933);
xnor U30915 (N_30915,N_27582,N_28076);
nor U30916 (N_30916,N_29558,N_28313);
or U30917 (N_30917,N_29618,N_28920);
or U30918 (N_30918,N_27897,N_27699);
nor U30919 (N_30919,N_29100,N_28510);
xnor U30920 (N_30920,N_29664,N_29728);
or U30921 (N_30921,N_29579,N_29276);
and U30922 (N_30922,N_29143,N_28950);
and U30923 (N_30923,N_29462,N_29666);
nor U30924 (N_30924,N_29968,N_29208);
nand U30925 (N_30925,N_28332,N_28099);
nor U30926 (N_30926,N_28484,N_28870);
nor U30927 (N_30927,N_29298,N_27765);
and U30928 (N_30928,N_29846,N_27522);
or U30929 (N_30929,N_29165,N_28802);
or U30930 (N_30930,N_29612,N_28063);
nand U30931 (N_30931,N_28639,N_29326);
xor U30932 (N_30932,N_29773,N_29252);
nor U30933 (N_30933,N_29181,N_28855);
nand U30934 (N_30934,N_29742,N_29917);
nor U30935 (N_30935,N_29585,N_29914);
xnor U30936 (N_30936,N_29253,N_29590);
and U30937 (N_30937,N_29348,N_29049);
nor U30938 (N_30938,N_27646,N_28433);
xnor U30939 (N_30939,N_27655,N_28825);
or U30940 (N_30940,N_28724,N_28612);
xnor U30941 (N_30941,N_29774,N_28489);
xor U30942 (N_30942,N_29224,N_29994);
nand U30943 (N_30943,N_27723,N_29026);
xnor U30944 (N_30944,N_28254,N_28811);
nor U30945 (N_30945,N_28754,N_29227);
xor U30946 (N_30946,N_29439,N_29980);
or U30947 (N_30947,N_27621,N_27928);
or U30948 (N_30948,N_27737,N_29850);
and U30949 (N_30949,N_28083,N_29745);
nand U30950 (N_30950,N_29293,N_28965);
or U30951 (N_30951,N_29308,N_28676);
nor U30952 (N_30952,N_29109,N_27759);
nand U30953 (N_30953,N_28408,N_29528);
nor U30954 (N_30954,N_27994,N_28486);
and U30955 (N_30955,N_29694,N_28513);
nor U30956 (N_30956,N_27958,N_28277);
nor U30957 (N_30957,N_27797,N_28103);
and U30958 (N_30958,N_29761,N_28416);
nand U30959 (N_30959,N_27608,N_27532);
nor U30960 (N_30960,N_28635,N_28415);
xnor U30961 (N_30961,N_28740,N_29982);
xnor U30962 (N_30962,N_29029,N_28039);
or U30963 (N_30963,N_28125,N_28748);
and U30964 (N_30964,N_27826,N_27886);
and U30965 (N_30965,N_29160,N_29444);
xor U30966 (N_30966,N_27653,N_29881);
nand U30967 (N_30967,N_28797,N_28329);
and U30968 (N_30968,N_28930,N_28320);
and U30969 (N_30969,N_28529,N_28845);
xor U30970 (N_30970,N_27825,N_28819);
nor U30971 (N_30971,N_29959,N_29406);
nand U30972 (N_30972,N_28956,N_29112);
nand U30973 (N_30973,N_29076,N_28907);
or U30974 (N_30974,N_28765,N_29643);
nand U30975 (N_30975,N_27649,N_27776);
nor U30976 (N_30976,N_29367,N_29184);
or U30977 (N_30977,N_28487,N_28991);
and U30978 (N_30978,N_29975,N_29767);
or U30979 (N_30979,N_29992,N_28195);
and U30980 (N_30980,N_28118,N_27767);
or U30981 (N_30981,N_28475,N_29626);
and U30982 (N_30982,N_29301,N_28850);
and U30983 (N_30983,N_27668,N_29064);
or U30984 (N_30984,N_28617,N_29188);
nor U30985 (N_30985,N_29435,N_28240);
xor U30986 (N_30986,N_29056,N_28689);
nor U30987 (N_30987,N_27739,N_27976);
nor U30988 (N_30988,N_29779,N_29347);
and U30989 (N_30989,N_28353,N_28846);
nand U30990 (N_30990,N_28147,N_28358);
or U30991 (N_30991,N_29655,N_29638);
nor U30992 (N_30992,N_29119,N_28726);
xor U30993 (N_30993,N_29665,N_29668);
xnor U30994 (N_30994,N_29936,N_27713);
or U30995 (N_30995,N_28389,N_29631);
or U30996 (N_30996,N_28090,N_28634);
xnor U30997 (N_30997,N_29580,N_27698);
and U30998 (N_30998,N_29833,N_27920);
and U30999 (N_30999,N_27704,N_28258);
or U31000 (N_31000,N_27732,N_29131);
and U31001 (N_31001,N_29412,N_28989);
and U31002 (N_31002,N_28093,N_29242);
xor U31003 (N_31003,N_28821,N_29330);
xnor U31004 (N_31004,N_28857,N_29196);
and U31005 (N_31005,N_27889,N_27845);
nand U31006 (N_31006,N_27643,N_28526);
nand U31007 (N_31007,N_29338,N_29376);
or U31008 (N_31008,N_27944,N_27613);
nand U31009 (N_31009,N_28399,N_28144);
or U31010 (N_31010,N_29514,N_28745);
nand U31011 (N_31011,N_27947,N_28403);
xnor U31012 (N_31012,N_28426,N_28916);
or U31013 (N_31013,N_27870,N_28401);
and U31014 (N_31014,N_29136,N_29120);
nand U31015 (N_31015,N_27823,N_28714);
xnor U31016 (N_31016,N_29277,N_28440);
nand U31017 (N_31017,N_29011,N_29421);
nor U31018 (N_31018,N_28688,N_29434);
nand U31019 (N_31019,N_27623,N_27722);
nand U31020 (N_31020,N_28050,N_29629);
xnor U31021 (N_31021,N_29213,N_28137);
nor U31022 (N_31022,N_29831,N_28205);
nor U31023 (N_31023,N_28703,N_29422);
nand U31024 (N_31024,N_29260,N_28402);
xor U31025 (N_31025,N_28071,N_27908);
or U31026 (N_31026,N_27850,N_28530);
nand U31027 (N_31027,N_29044,N_29349);
and U31028 (N_31028,N_28555,N_29411);
xnor U31029 (N_31029,N_29057,N_29511);
xor U31030 (N_31030,N_27688,N_29146);
or U31031 (N_31031,N_28793,N_27896);
nor U31032 (N_31032,N_27949,N_28665);
nor U31033 (N_31033,N_28284,N_28706);
nor U31034 (N_31034,N_28315,N_29307);
or U31035 (N_31035,N_29110,N_29993);
nor U31036 (N_31036,N_29848,N_29615);
xnor U31037 (N_31037,N_28148,N_27641);
nand U31038 (N_31038,N_28893,N_29289);
xnor U31039 (N_31039,N_27625,N_27583);
or U31040 (N_31040,N_29587,N_29795);
xor U31041 (N_31041,N_29573,N_28203);
xnor U31042 (N_31042,N_29991,N_29555);
nor U31043 (N_31043,N_28168,N_29225);
nand U31044 (N_31044,N_29739,N_28007);
and U31045 (N_31045,N_28124,N_27519);
or U31046 (N_31046,N_29387,N_28262);
nand U31047 (N_31047,N_27560,N_27931);
nor U31048 (N_31048,N_28642,N_29606);
or U31049 (N_31049,N_28328,N_28119);
or U31050 (N_31050,N_29695,N_28715);
nand U31051 (N_31051,N_29711,N_28377);
and U31052 (N_31052,N_29065,N_28397);
and U31053 (N_31053,N_28565,N_29152);
nand U31054 (N_31054,N_29328,N_28955);
or U31055 (N_31055,N_28293,N_29288);
xnor U31056 (N_31056,N_29865,N_28464);
and U31057 (N_31057,N_28065,N_28503);
and U31058 (N_31058,N_28428,N_29279);
nor U31059 (N_31059,N_29803,N_28263);
nand U31060 (N_31060,N_29086,N_29671);
nor U31061 (N_31061,N_29037,N_28024);
nor U31062 (N_31062,N_28016,N_27580);
xor U31063 (N_31063,N_28298,N_28649);
nand U31064 (N_31064,N_29723,N_28654);
xnor U31065 (N_31065,N_29058,N_29280);
xnor U31066 (N_31066,N_28216,N_28523);
nand U31067 (N_31067,N_29379,N_29667);
or U31068 (N_31068,N_29228,N_27820);
nor U31069 (N_31069,N_28869,N_29442);
nand U31070 (N_31070,N_28803,N_28238);
nor U31071 (N_31071,N_29189,N_28300);
xnor U31072 (N_31072,N_29951,N_29984);
or U31073 (N_31073,N_28852,N_29972);
nor U31074 (N_31074,N_28934,N_28763);
xnor U31075 (N_31075,N_29857,N_27618);
nor U31076 (N_31076,N_29611,N_28321);
nand U31077 (N_31077,N_29372,N_28080);
or U31078 (N_31078,N_29875,N_29267);
and U31079 (N_31079,N_27747,N_28445);
xor U31080 (N_31080,N_29813,N_28012);
or U31081 (N_31081,N_28404,N_27852);
or U31082 (N_31082,N_27786,N_27911);
xor U31083 (N_31083,N_29365,N_29122);
and U31084 (N_31084,N_28186,N_27504);
or U31085 (N_31085,N_27716,N_28901);
nand U31086 (N_31086,N_29658,N_27663);
nor U31087 (N_31087,N_29818,N_28831);
nand U31088 (N_31088,N_29364,N_27748);
and U31089 (N_31089,N_29830,N_29896);
and U31090 (N_31090,N_27818,N_29323);
nor U31091 (N_31091,N_29193,N_27678);
or U31092 (N_31092,N_27864,N_29194);
nor U31093 (N_31093,N_28407,N_29478);
nand U31094 (N_31094,N_29598,N_28914);
or U31095 (N_31095,N_28128,N_28257);
and U31096 (N_31096,N_29430,N_28165);
xnor U31097 (N_31097,N_27597,N_29030);
and U31098 (N_31098,N_27967,N_28223);
nand U31099 (N_31099,N_29939,N_28236);
nand U31100 (N_31100,N_28913,N_27806);
nand U31101 (N_31101,N_28538,N_27898);
and U31102 (N_31102,N_29325,N_28055);
nand U31103 (N_31103,N_28317,N_27849);
nand U31104 (N_31104,N_29793,N_28854);
and U31105 (N_31105,N_28327,N_29493);
and U31106 (N_31106,N_29610,N_29760);
nor U31107 (N_31107,N_27902,N_28601);
or U31108 (N_31108,N_28073,N_29104);
nand U31109 (N_31109,N_28348,N_29539);
nand U31110 (N_31110,N_29563,N_29238);
or U31111 (N_31111,N_29557,N_29394);
nand U31112 (N_31112,N_29456,N_27878);
nand U31113 (N_31113,N_27514,N_27954);
or U31114 (N_31114,N_27746,N_29752);
and U31115 (N_31115,N_29912,N_29508);
and U31116 (N_31116,N_28581,N_28269);
xor U31117 (N_31117,N_27735,N_29463);
or U31118 (N_31118,N_29622,N_29312);
nor U31119 (N_31119,N_27998,N_29844);
nand U31120 (N_31120,N_28376,N_27978);
nand U31121 (N_31121,N_28683,N_28769);
nor U31122 (N_31122,N_29386,N_28691);
xor U31123 (N_31123,N_29046,N_28690);
nor U31124 (N_31124,N_28882,N_29089);
xnor U31125 (N_31125,N_28333,N_29820);
xnor U31126 (N_31126,N_27971,N_27946);
or U31127 (N_31127,N_27872,N_29408);
nand U31128 (N_31128,N_27592,N_28552);
nor U31129 (N_31129,N_29066,N_27517);
or U31130 (N_31130,N_29527,N_29138);
and U31131 (N_31131,N_28106,N_27524);
or U31132 (N_31132,N_27508,N_28380);
or U31133 (N_31133,N_29342,N_29117);
nor U31134 (N_31134,N_28021,N_28011);
nor U31135 (N_31135,N_28922,N_29572);
xnor U31136 (N_31136,N_29209,N_28624);
nand U31137 (N_31137,N_29304,N_29207);
nand U31138 (N_31138,N_29753,N_28889);
and U31139 (N_31139,N_29687,N_28640);
nand U31140 (N_31140,N_29278,N_29286);
nor U31141 (N_31141,N_27695,N_29284);
nand U31142 (N_31142,N_29596,N_29105);
nor U31143 (N_31143,N_28496,N_29256);
nor U31144 (N_31144,N_29476,N_28150);
or U31145 (N_31145,N_28767,N_27885);
and U31146 (N_31146,N_28902,N_29565);
nand U31147 (N_31147,N_27697,N_29036);
or U31148 (N_31148,N_29071,N_29032);
xnor U31149 (N_31149,N_28488,N_28264);
nand U31150 (N_31150,N_28274,N_29137);
and U31151 (N_31151,N_29660,N_28385);
and U31152 (N_31152,N_29504,N_27743);
or U31153 (N_31153,N_28245,N_29916);
nand U31154 (N_31154,N_29261,N_27573);
nor U31155 (N_31155,N_29777,N_28791);
xor U31156 (N_31156,N_28656,N_27843);
nand U31157 (N_31157,N_29198,N_29173);
or U31158 (N_31158,N_29894,N_29081);
and U31159 (N_31159,N_27691,N_28787);
nand U31160 (N_31160,N_29416,N_28833);
nand U31161 (N_31161,N_29397,N_28643);
xor U31162 (N_31162,N_29977,N_29808);
and U31163 (N_31163,N_27901,N_28894);
xor U31164 (N_31164,N_29006,N_27968);
nor U31165 (N_31165,N_28877,N_28143);
nor U31166 (N_31166,N_28356,N_29357);
xnor U31167 (N_31167,N_29445,N_29554);
and U31168 (N_31168,N_28282,N_28301);
or U31169 (N_31169,N_27692,N_29649);
or U31170 (N_31170,N_28208,N_27651);
xor U31171 (N_31171,N_29072,N_29465);
and U31172 (N_31172,N_28159,N_28851);
nor U31173 (N_31173,N_27727,N_28776);
xor U31174 (N_31174,N_29050,N_28593);
nand U31175 (N_31175,N_27844,N_27903);
nor U31176 (N_31176,N_29123,N_28716);
and U31177 (N_31177,N_29776,N_29737);
nor U31178 (N_31178,N_28166,N_27553);
and U31179 (N_31179,N_28442,N_29847);
or U31180 (N_31180,N_29126,N_27579);
xor U31181 (N_31181,N_27982,N_27556);
and U31182 (N_31182,N_27752,N_28121);
nor U31183 (N_31183,N_27719,N_28279);
nand U31184 (N_31184,N_29766,N_28898);
or U31185 (N_31185,N_28792,N_29503);
and U31186 (N_31186,N_28830,N_27685);
xnor U31187 (N_31187,N_29500,N_29719);
nor U31188 (N_31188,N_28720,N_28087);
and U31189 (N_31189,N_29241,N_27725);
nand U31190 (N_31190,N_28045,N_27565);
and U31191 (N_31191,N_28362,N_27590);
nand U31192 (N_31192,N_29738,N_27636);
xnor U31193 (N_31193,N_29063,N_29677);
or U31194 (N_31194,N_27913,N_28163);
nor U31195 (N_31195,N_28214,N_29140);
nor U31196 (N_31196,N_28305,N_27891);
xnor U31197 (N_31197,N_28899,N_28409);
nand U31198 (N_31198,N_28829,N_29935);
or U31199 (N_31199,N_29141,N_28448);
and U31200 (N_31200,N_29266,N_27622);
nor U31201 (N_31201,N_29077,N_29128);
xnor U31202 (N_31202,N_28671,N_29275);
or U31203 (N_31203,N_29233,N_27802);
nor U31204 (N_31204,N_28608,N_27904);
or U31205 (N_31205,N_29913,N_27584);
nor U31206 (N_31206,N_29849,N_28659);
and U31207 (N_31207,N_29945,N_29559);
and U31208 (N_31208,N_29447,N_29860);
nand U31209 (N_31209,N_29772,N_29362);
nor U31210 (N_31210,N_28972,N_27569);
nor U31211 (N_31211,N_29441,N_29600);
or U31212 (N_31212,N_27701,N_29595);
or U31213 (N_31213,N_27614,N_28363);
nor U31214 (N_31214,N_28694,N_28574);
nand U31215 (N_31215,N_29375,N_29544);
xor U31216 (N_31216,N_29725,N_29431);
or U31217 (N_31217,N_27632,N_28906);
xnor U31218 (N_31218,N_27548,N_28075);
nand U31219 (N_31219,N_28037,N_27512);
nand U31220 (N_31220,N_27926,N_29302);
xnor U31221 (N_31221,N_28188,N_29161);
and U31222 (N_31222,N_28929,N_28431);
xor U31223 (N_31223,N_29802,N_28308);
nor U31224 (N_31224,N_28896,N_29363);
or U31225 (N_31225,N_28848,N_27680);
and U31226 (N_31226,N_28951,N_29170);
and U31227 (N_31227,N_29786,N_27545);
or U31228 (N_31228,N_29502,N_28290);
nor U31229 (N_31229,N_28419,N_29346);
xor U31230 (N_31230,N_27745,N_29175);
or U31231 (N_31231,N_29370,N_27756);
xnor U31232 (N_31232,N_28655,N_28455);
xnor U31233 (N_31233,N_29337,N_27862);
or U31234 (N_31234,N_27715,N_27554);
nor U31235 (N_31235,N_29354,N_29210);
nor U31236 (N_31236,N_29418,N_29542);
xnor U31237 (N_31237,N_27575,N_29287);
and U31238 (N_31238,N_29315,N_28132);
nand U31239 (N_31239,N_29903,N_28876);
and U31240 (N_31240,N_28926,N_29000);
and U31241 (N_31241,N_28653,N_29759);
nor U31242 (N_31242,N_29907,N_27827);
nor U31243 (N_31243,N_29258,N_28970);
xnor U31244 (N_31244,N_29796,N_28086);
xor U31245 (N_31245,N_28677,N_27952);
xnor U31246 (N_31246,N_28699,N_28079);
nor U31247 (N_31247,N_28619,N_28215);
nand U31248 (N_31248,N_29999,N_28798);
nand U31249 (N_31249,N_27518,N_29676);
and U31250 (N_31250,N_27843,N_29744);
or U31251 (N_31251,N_29809,N_28169);
or U31252 (N_31252,N_27915,N_29351);
xor U31253 (N_31253,N_28937,N_29217);
and U31254 (N_31254,N_27865,N_29831);
xnor U31255 (N_31255,N_27644,N_29047);
or U31256 (N_31256,N_28072,N_28494);
xor U31257 (N_31257,N_27670,N_29105);
nor U31258 (N_31258,N_29555,N_29465);
or U31259 (N_31259,N_28665,N_28443);
nand U31260 (N_31260,N_28005,N_29489);
and U31261 (N_31261,N_28858,N_29718);
or U31262 (N_31262,N_29198,N_27638);
or U31263 (N_31263,N_28621,N_27758);
xor U31264 (N_31264,N_29762,N_27773);
nand U31265 (N_31265,N_27730,N_29481);
or U31266 (N_31266,N_29761,N_29562);
or U31267 (N_31267,N_29500,N_28744);
or U31268 (N_31268,N_29895,N_29298);
and U31269 (N_31269,N_29168,N_28191);
nor U31270 (N_31270,N_29671,N_29233);
and U31271 (N_31271,N_29434,N_29363);
xnor U31272 (N_31272,N_27824,N_28042);
and U31273 (N_31273,N_27721,N_29148);
nand U31274 (N_31274,N_28047,N_28489);
and U31275 (N_31275,N_29886,N_27730);
nand U31276 (N_31276,N_27797,N_27961);
or U31277 (N_31277,N_28429,N_28232);
or U31278 (N_31278,N_28010,N_27637);
and U31279 (N_31279,N_27903,N_28864);
or U31280 (N_31280,N_29847,N_29921);
nor U31281 (N_31281,N_29667,N_28384);
nor U31282 (N_31282,N_27768,N_27737);
or U31283 (N_31283,N_29327,N_29631);
or U31284 (N_31284,N_29485,N_28188);
nor U31285 (N_31285,N_28989,N_28807);
xor U31286 (N_31286,N_27941,N_29836);
or U31287 (N_31287,N_27972,N_29363);
xor U31288 (N_31288,N_28261,N_29302);
nor U31289 (N_31289,N_27716,N_29502);
and U31290 (N_31290,N_29119,N_28218);
and U31291 (N_31291,N_29211,N_28359);
and U31292 (N_31292,N_28637,N_27980);
and U31293 (N_31293,N_29725,N_29210);
nand U31294 (N_31294,N_29971,N_28513);
and U31295 (N_31295,N_27846,N_29225);
nor U31296 (N_31296,N_29088,N_28507);
nor U31297 (N_31297,N_29247,N_29694);
nand U31298 (N_31298,N_27584,N_28551);
nor U31299 (N_31299,N_27501,N_29577);
nand U31300 (N_31300,N_29320,N_28682);
nand U31301 (N_31301,N_28020,N_29053);
xor U31302 (N_31302,N_27856,N_28831);
xor U31303 (N_31303,N_27989,N_29838);
and U31304 (N_31304,N_28139,N_28562);
xor U31305 (N_31305,N_27706,N_27979);
nor U31306 (N_31306,N_29313,N_29150);
or U31307 (N_31307,N_28679,N_29910);
and U31308 (N_31308,N_27708,N_28556);
or U31309 (N_31309,N_28058,N_29865);
or U31310 (N_31310,N_29267,N_28929);
nand U31311 (N_31311,N_29164,N_29081);
or U31312 (N_31312,N_28642,N_27942);
nand U31313 (N_31313,N_29203,N_29837);
and U31314 (N_31314,N_28268,N_28498);
or U31315 (N_31315,N_29425,N_29723);
or U31316 (N_31316,N_27713,N_28356);
xnor U31317 (N_31317,N_29628,N_28422);
or U31318 (N_31318,N_29586,N_29840);
xor U31319 (N_31319,N_28117,N_27867);
nand U31320 (N_31320,N_28522,N_28366);
xnor U31321 (N_31321,N_28352,N_29500);
xor U31322 (N_31322,N_29340,N_29988);
nor U31323 (N_31323,N_28104,N_28198);
and U31324 (N_31324,N_29628,N_28056);
and U31325 (N_31325,N_27584,N_29976);
and U31326 (N_31326,N_27858,N_29394);
xnor U31327 (N_31327,N_29488,N_29205);
nor U31328 (N_31328,N_27718,N_29424);
or U31329 (N_31329,N_28412,N_29328);
xor U31330 (N_31330,N_28732,N_29879);
or U31331 (N_31331,N_28976,N_29347);
nor U31332 (N_31332,N_28608,N_27696);
or U31333 (N_31333,N_28545,N_27940);
and U31334 (N_31334,N_29280,N_28330);
nor U31335 (N_31335,N_29248,N_29512);
nor U31336 (N_31336,N_28163,N_28843);
nor U31337 (N_31337,N_29172,N_28574);
nand U31338 (N_31338,N_29298,N_28585);
or U31339 (N_31339,N_29533,N_29057);
or U31340 (N_31340,N_29876,N_27824);
or U31341 (N_31341,N_28986,N_28671);
nor U31342 (N_31342,N_27813,N_27736);
xor U31343 (N_31343,N_27853,N_29774);
and U31344 (N_31344,N_29697,N_29830);
xor U31345 (N_31345,N_28677,N_27713);
xor U31346 (N_31346,N_29011,N_27566);
nand U31347 (N_31347,N_29188,N_28269);
and U31348 (N_31348,N_27919,N_27531);
and U31349 (N_31349,N_29067,N_27883);
or U31350 (N_31350,N_29279,N_29522);
nand U31351 (N_31351,N_28057,N_28882);
nor U31352 (N_31352,N_27605,N_27853);
and U31353 (N_31353,N_27846,N_29081);
or U31354 (N_31354,N_29057,N_29065);
xnor U31355 (N_31355,N_28237,N_27874);
and U31356 (N_31356,N_28233,N_28691);
and U31357 (N_31357,N_29876,N_28360);
xnor U31358 (N_31358,N_29096,N_28524);
and U31359 (N_31359,N_28562,N_28304);
and U31360 (N_31360,N_28602,N_27572);
nor U31361 (N_31361,N_29441,N_29498);
or U31362 (N_31362,N_27882,N_28096);
xor U31363 (N_31363,N_29837,N_28762);
nor U31364 (N_31364,N_28721,N_29948);
and U31365 (N_31365,N_29769,N_28643);
xor U31366 (N_31366,N_28183,N_28352);
xnor U31367 (N_31367,N_29288,N_28096);
nand U31368 (N_31368,N_29833,N_27667);
nor U31369 (N_31369,N_27891,N_27975);
nand U31370 (N_31370,N_29769,N_28915);
and U31371 (N_31371,N_28420,N_28636);
or U31372 (N_31372,N_28512,N_28676);
and U31373 (N_31373,N_29337,N_29585);
or U31374 (N_31374,N_28135,N_27567);
nand U31375 (N_31375,N_29648,N_27999);
nor U31376 (N_31376,N_28553,N_28980);
nor U31377 (N_31377,N_28600,N_28382);
or U31378 (N_31378,N_28899,N_28740);
and U31379 (N_31379,N_27594,N_29101);
xnor U31380 (N_31380,N_28197,N_27577);
nand U31381 (N_31381,N_29480,N_28545);
and U31382 (N_31382,N_28919,N_27922);
nand U31383 (N_31383,N_28828,N_29537);
and U31384 (N_31384,N_27502,N_28236);
and U31385 (N_31385,N_27699,N_29057);
nor U31386 (N_31386,N_28186,N_29302);
or U31387 (N_31387,N_29493,N_28143);
or U31388 (N_31388,N_29857,N_28018);
nor U31389 (N_31389,N_28083,N_29552);
nor U31390 (N_31390,N_28405,N_27764);
and U31391 (N_31391,N_27949,N_29626);
nand U31392 (N_31392,N_28452,N_28502);
and U31393 (N_31393,N_27532,N_27545);
xor U31394 (N_31394,N_27583,N_29190);
xnor U31395 (N_31395,N_29463,N_28277);
nor U31396 (N_31396,N_29467,N_29840);
xnor U31397 (N_31397,N_29419,N_27963);
xor U31398 (N_31398,N_29483,N_28143);
nand U31399 (N_31399,N_28006,N_28571);
nand U31400 (N_31400,N_28676,N_27678);
and U31401 (N_31401,N_29130,N_27813);
xor U31402 (N_31402,N_28565,N_29633);
nor U31403 (N_31403,N_28620,N_29187);
nor U31404 (N_31404,N_28176,N_27560);
xnor U31405 (N_31405,N_28153,N_28492);
nand U31406 (N_31406,N_27652,N_27970);
xor U31407 (N_31407,N_28666,N_28844);
or U31408 (N_31408,N_28946,N_27590);
nor U31409 (N_31409,N_28739,N_27786);
nor U31410 (N_31410,N_28332,N_27586);
and U31411 (N_31411,N_29396,N_28048);
nand U31412 (N_31412,N_28609,N_27784);
or U31413 (N_31413,N_28792,N_29633);
and U31414 (N_31414,N_28655,N_27854);
nor U31415 (N_31415,N_27871,N_29096);
or U31416 (N_31416,N_28632,N_27945);
xor U31417 (N_31417,N_29600,N_28797);
or U31418 (N_31418,N_28430,N_27774);
or U31419 (N_31419,N_29121,N_28064);
and U31420 (N_31420,N_27650,N_29692);
nor U31421 (N_31421,N_28492,N_27846);
or U31422 (N_31422,N_27502,N_28356);
xor U31423 (N_31423,N_28444,N_27869);
and U31424 (N_31424,N_29865,N_28075);
nor U31425 (N_31425,N_29543,N_28034);
xor U31426 (N_31426,N_29323,N_28641);
nor U31427 (N_31427,N_28276,N_29128);
xor U31428 (N_31428,N_28916,N_27503);
nand U31429 (N_31429,N_29851,N_28828);
and U31430 (N_31430,N_28040,N_28971);
and U31431 (N_31431,N_28559,N_29855);
nor U31432 (N_31432,N_27620,N_29648);
and U31433 (N_31433,N_29845,N_29040);
and U31434 (N_31434,N_29439,N_28015);
and U31435 (N_31435,N_29296,N_27560);
and U31436 (N_31436,N_28120,N_29178);
xor U31437 (N_31437,N_29015,N_29955);
xnor U31438 (N_31438,N_29846,N_29173);
and U31439 (N_31439,N_27703,N_29029);
nor U31440 (N_31440,N_29288,N_29211);
or U31441 (N_31441,N_27794,N_29297);
xnor U31442 (N_31442,N_28595,N_28525);
nor U31443 (N_31443,N_29324,N_29428);
nand U31444 (N_31444,N_28875,N_28314);
or U31445 (N_31445,N_27647,N_29380);
or U31446 (N_31446,N_29062,N_29308);
nand U31447 (N_31447,N_28130,N_29891);
xnor U31448 (N_31448,N_28916,N_27756);
xnor U31449 (N_31449,N_27783,N_29828);
xnor U31450 (N_31450,N_28261,N_29690);
xnor U31451 (N_31451,N_29684,N_28405);
nand U31452 (N_31452,N_28486,N_28838);
xnor U31453 (N_31453,N_28101,N_28493);
or U31454 (N_31454,N_28277,N_29356);
and U31455 (N_31455,N_28118,N_28979);
nor U31456 (N_31456,N_27629,N_29934);
nand U31457 (N_31457,N_29283,N_29982);
or U31458 (N_31458,N_29347,N_29698);
nor U31459 (N_31459,N_28193,N_29809);
and U31460 (N_31460,N_27987,N_29318);
xnor U31461 (N_31461,N_29948,N_29509);
xnor U31462 (N_31462,N_28926,N_28184);
or U31463 (N_31463,N_29018,N_27552);
nor U31464 (N_31464,N_28075,N_27731);
or U31465 (N_31465,N_28671,N_29166);
xor U31466 (N_31466,N_29117,N_28947);
or U31467 (N_31467,N_27962,N_28846);
or U31468 (N_31468,N_28443,N_28677);
or U31469 (N_31469,N_29465,N_29616);
or U31470 (N_31470,N_28174,N_29398);
or U31471 (N_31471,N_29372,N_28432);
nand U31472 (N_31472,N_29652,N_29952);
or U31473 (N_31473,N_29651,N_29615);
nand U31474 (N_31474,N_29086,N_29867);
nor U31475 (N_31475,N_27641,N_28412);
or U31476 (N_31476,N_28105,N_29779);
xnor U31477 (N_31477,N_29588,N_29539);
or U31478 (N_31478,N_29332,N_29294);
nor U31479 (N_31479,N_28324,N_27822);
or U31480 (N_31480,N_29409,N_29289);
xor U31481 (N_31481,N_28259,N_29977);
and U31482 (N_31482,N_28586,N_28854);
or U31483 (N_31483,N_29755,N_28757);
xnor U31484 (N_31484,N_27749,N_28307);
and U31485 (N_31485,N_27838,N_28909);
nand U31486 (N_31486,N_29043,N_29255);
or U31487 (N_31487,N_27850,N_29415);
and U31488 (N_31488,N_29299,N_29127);
nor U31489 (N_31489,N_28284,N_29873);
or U31490 (N_31490,N_28582,N_28745);
xnor U31491 (N_31491,N_28433,N_29080);
and U31492 (N_31492,N_28305,N_28103);
nand U31493 (N_31493,N_29529,N_28242);
and U31494 (N_31494,N_28094,N_27911);
xor U31495 (N_31495,N_29031,N_29610);
xnor U31496 (N_31496,N_28984,N_28494);
or U31497 (N_31497,N_27822,N_29335);
nor U31498 (N_31498,N_29590,N_29166);
and U31499 (N_31499,N_27831,N_28630);
xor U31500 (N_31500,N_29152,N_29139);
or U31501 (N_31501,N_28554,N_27684);
and U31502 (N_31502,N_29416,N_28687);
or U31503 (N_31503,N_29540,N_29421);
nor U31504 (N_31504,N_28470,N_27707);
or U31505 (N_31505,N_28188,N_29583);
nand U31506 (N_31506,N_27727,N_27704);
nor U31507 (N_31507,N_29656,N_29149);
xor U31508 (N_31508,N_29422,N_29219);
xor U31509 (N_31509,N_27967,N_27795);
nand U31510 (N_31510,N_29135,N_28497);
nand U31511 (N_31511,N_28518,N_28609);
nor U31512 (N_31512,N_28509,N_28726);
and U31513 (N_31513,N_29727,N_28859);
nor U31514 (N_31514,N_27770,N_28486);
and U31515 (N_31515,N_27902,N_28906);
nor U31516 (N_31516,N_28416,N_28656);
xnor U31517 (N_31517,N_29314,N_29249);
nor U31518 (N_31518,N_29094,N_28009);
xnor U31519 (N_31519,N_28483,N_28400);
or U31520 (N_31520,N_29438,N_29439);
xnor U31521 (N_31521,N_28820,N_29847);
nor U31522 (N_31522,N_29980,N_29681);
xor U31523 (N_31523,N_29463,N_27939);
and U31524 (N_31524,N_29954,N_29645);
xnor U31525 (N_31525,N_29785,N_29589);
and U31526 (N_31526,N_29469,N_28759);
or U31527 (N_31527,N_28438,N_29874);
and U31528 (N_31528,N_28741,N_29591);
and U31529 (N_31529,N_28280,N_28893);
or U31530 (N_31530,N_28804,N_27820);
nand U31531 (N_31531,N_29649,N_29552);
nand U31532 (N_31532,N_29144,N_28251);
xor U31533 (N_31533,N_27505,N_27907);
nand U31534 (N_31534,N_29646,N_28051);
nand U31535 (N_31535,N_28646,N_28378);
xnor U31536 (N_31536,N_27926,N_28051);
or U31537 (N_31537,N_28376,N_29097);
xnor U31538 (N_31538,N_28300,N_28614);
and U31539 (N_31539,N_29313,N_28920);
xnor U31540 (N_31540,N_28691,N_29914);
xor U31541 (N_31541,N_28428,N_27835);
xor U31542 (N_31542,N_27948,N_27824);
nand U31543 (N_31543,N_28115,N_28612);
nor U31544 (N_31544,N_28281,N_29684);
nand U31545 (N_31545,N_28534,N_29594);
xnor U31546 (N_31546,N_27598,N_28299);
nand U31547 (N_31547,N_28291,N_28317);
or U31548 (N_31548,N_28520,N_28823);
or U31549 (N_31549,N_27880,N_27949);
nor U31550 (N_31550,N_28421,N_27904);
nand U31551 (N_31551,N_28967,N_29124);
nor U31552 (N_31552,N_28512,N_28491);
or U31553 (N_31553,N_29048,N_29784);
xor U31554 (N_31554,N_29647,N_28161);
xor U31555 (N_31555,N_29940,N_28232);
and U31556 (N_31556,N_29016,N_28727);
nor U31557 (N_31557,N_28642,N_29609);
xnor U31558 (N_31558,N_29550,N_29588);
xnor U31559 (N_31559,N_28563,N_28807);
nand U31560 (N_31560,N_28536,N_29622);
nor U31561 (N_31561,N_28341,N_27951);
xor U31562 (N_31562,N_29130,N_28015);
nand U31563 (N_31563,N_29485,N_28649);
and U31564 (N_31564,N_27966,N_28569);
xnor U31565 (N_31565,N_27728,N_28461);
or U31566 (N_31566,N_28766,N_29616);
xnor U31567 (N_31567,N_28475,N_29623);
nor U31568 (N_31568,N_28812,N_28421);
or U31569 (N_31569,N_29423,N_28817);
nor U31570 (N_31570,N_27546,N_28879);
xnor U31571 (N_31571,N_29826,N_29554);
nand U31572 (N_31572,N_29580,N_29408);
xor U31573 (N_31573,N_29590,N_28997);
nand U31574 (N_31574,N_29837,N_28708);
or U31575 (N_31575,N_29345,N_27973);
nor U31576 (N_31576,N_27964,N_28297);
and U31577 (N_31577,N_27802,N_28298);
nor U31578 (N_31578,N_29007,N_28834);
or U31579 (N_31579,N_27710,N_29589);
and U31580 (N_31580,N_28927,N_28897);
xor U31581 (N_31581,N_28904,N_27624);
nand U31582 (N_31582,N_28611,N_29777);
or U31583 (N_31583,N_29294,N_27513);
xor U31584 (N_31584,N_29036,N_27998);
or U31585 (N_31585,N_28003,N_28168);
or U31586 (N_31586,N_29088,N_28457);
nor U31587 (N_31587,N_28500,N_28585);
nor U31588 (N_31588,N_28363,N_29164);
and U31589 (N_31589,N_29918,N_29546);
xnor U31590 (N_31590,N_27797,N_27832);
nand U31591 (N_31591,N_28812,N_27600);
or U31592 (N_31592,N_28175,N_28413);
nand U31593 (N_31593,N_28622,N_28798);
nand U31594 (N_31594,N_27965,N_28920);
and U31595 (N_31595,N_27673,N_29657);
or U31596 (N_31596,N_29963,N_28507);
xor U31597 (N_31597,N_29740,N_27992);
and U31598 (N_31598,N_28673,N_28366);
nand U31599 (N_31599,N_27520,N_28321);
xor U31600 (N_31600,N_29708,N_29934);
nor U31601 (N_31601,N_27694,N_28840);
or U31602 (N_31602,N_28748,N_27714);
xor U31603 (N_31603,N_28094,N_28819);
nand U31604 (N_31604,N_29562,N_28226);
nor U31605 (N_31605,N_29749,N_29913);
and U31606 (N_31606,N_29718,N_28654);
xnor U31607 (N_31607,N_29789,N_27830);
nand U31608 (N_31608,N_29421,N_28803);
xor U31609 (N_31609,N_28270,N_28597);
and U31610 (N_31610,N_27697,N_28438);
xnor U31611 (N_31611,N_28797,N_28753);
nand U31612 (N_31612,N_27544,N_29666);
and U31613 (N_31613,N_28812,N_27934);
or U31614 (N_31614,N_29999,N_29101);
or U31615 (N_31615,N_28177,N_29754);
nand U31616 (N_31616,N_29436,N_29887);
and U31617 (N_31617,N_28347,N_28158);
nor U31618 (N_31618,N_27521,N_28799);
xor U31619 (N_31619,N_28811,N_29559);
or U31620 (N_31620,N_27502,N_28960);
xor U31621 (N_31621,N_28258,N_28731);
nor U31622 (N_31622,N_29188,N_29369);
and U31623 (N_31623,N_28585,N_28543);
or U31624 (N_31624,N_29296,N_29324);
nand U31625 (N_31625,N_28528,N_28714);
nand U31626 (N_31626,N_28088,N_28141);
and U31627 (N_31627,N_28319,N_29663);
nand U31628 (N_31628,N_28988,N_29690);
xor U31629 (N_31629,N_29275,N_28213);
nor U31630 (N_31630,N_28780,N_28652);
nor U31631 (N_31631,N_29486,N_27560);
and U31632 (N_31632,N_28305,N_29156);
nor U31633 (N_31633,N_27765,N_29224);
nand U31634 (N_31634,N_29042,N_27664);
nand U31635 (N_31635,N_29963,N_29898);
nand U31636 (N_31636,N_29784,N_28298);
nor U31637 (N_31637,N_27948,N_27979);
and U31638 (N_31638,N_28382,N_28320);
nand U31639 (N_31639,N_29809,N_29888);
nor U31640 (N_31640,N_29614,N_29430);
and U31641 (N_31641,N_28333,N_29452);
nand U31642 (N_31642,N_29320,N_27746);
or U31643 (N_31643,N_28936,N_29785);
and U31644 (N_31644,N_29807,N_27571);
xor U31645 (N_31645,N_29320,N_29476);
and U31646 (N_31646,N_29367,N_29168);
nand U31647 (N_31647,N_29393,N_27628);
xnor U31648 (N_31648,N_29351,N_29154);
and U31649 (N_31649,N_27862,N_29131);
nand U31650 (N_31650,N_29705,N_27939);
nand U31651 (N_31651,N_28170,N_28074);
xor U31652 (N_31652,N_28150,N_27727);
nor U31653 (N_31653,N_28376,N_28527);
or U31654 (N_31654,N_28901,N_27715);
and U31655 (N_31655,N_27669,N_28882);
nor U31656 (N_31656,N_28231,N_27940);
nor U31657 (N_31657,N_29838,N_29104);
and U31658 (N_31658,N_28951,N_29779);
or U31659 (N_31659,N_28873,N_29389);
nor U31660 (N_31660,N_27682,N_28043);
nor U31661 (N_31661,N_29678,N_27987);
nor U31662 (N_31662,N_27500,N_29511);
and U31663 (N_31663,N_27774,N_29958);
xor U31664 (N_31664,N_27662,N_27859);
xnor U31665 (N_31665,N_29417,N_29226);
nand U31666 (N_31666,N_27635,N_27787);
xor U31667 (N_31667,N_28183,N_27517);
nand U31668 (N_31668,N_29442,N_28525);
nor U31669 (N_31669,N_28381,N_28962);
nor U31670 (N_31670,N_29881,N_29660);
and U31671 (N_31671,N_29539,N_27796);
nor U31672 (N_31672,N_29152,N_28756);
or U31673 (N_31673,N_28188,N_28107);
nand U31674 (N_31674,N_28554,N_29233);
nand U31675 (N_31675,N_27916,N_29321);
or U31676 (N_31676,N_29427,N_29836);
or U31677 (N_31677,N_28492,N_28238);
nand U31678 (N_31678,N_29478,N_28983);
or U31679 (N_31679,N_28345,N_28568);
or U31680 (N_31680,N_27999,N_28872);
nor U31681 (N_31681,N_28548,N_28224);
xor U31682 (N_31682,N_29334,N_27895);
and U31683 (N_31683,N_27506,N_29064);
and U31684 (N_31684,N_27738,N_29049);
or U31685 (N_31685,N_29865,N_27514);
nand U31686 (N_31686,N_29736,N_28982);
and U31687 (N_31687,N_29058,N_28336);
nand U31688 (N_31688,N_27535,N_28526);
and U31689 (N_31689,N_27797,N_27909);
nand U31690 (N_31690,N_28079,N_28494);
and U31691 (N_31691,N_27540,N_29814);
nand U31692 (N_31692,N_29189,N_29537);
and U31693 (N_31693,N_28019,N_27953);
or U31694 (N_31694,N_27707,N_28120);
and U31695 (N_31695,N_29934,N_28618);
nor U31696 (N_31696,N_28045,N_27699);
xor U31697 (N_31697,N_29430,N_29636);
and U31698 (N_31698,N_27672,N_29887);
and U31699 (N_31699,N_28197,N_29901);
or U31700 (N_31700,N_29969,N_28337);
or U31701 (N_31701,N_28919,N_29810);
xor U31702 (N_31702,N_28916,N_29409);
xnor U31703 (N_31703,N_28831,N_28318);
and U31704 (N_31704,N_29381,N_28599);
nor U31705 (N_31705,N_28805,N_29892);
xor U31706 (N_31706,N_28876,N_27509);
xnor U31707 (N_31707,N_28869,N_27777);
nand U31708 (N_31708,N_28360,N_27920);
nand U31709 (N_31709,N_27649,N_28910);
or U31710 (N_31710,N_27512,N_27542);
nand U31711 (N_31711,N_29958,N_28802);
nor U31712 (N_31712,N_29203,N_28572);
and U31713 (N_31713,N_28033,N_27531);
nand U31714 (N_31714,N_28891,N_28394);
or U31715 (N_31715,N_29115,N_29037);
xnor U31716 (N_31716,N_29713,N_28651);
and U31717 (N_31717,N_28456,N_28213);
or U31718 (N_31718,N_28838,N_29422);
or U31719 (N_31719,N_27654,N_29989);
nor U31720 (N_31720,N_28164,N_28775);
and U31721 (N_31721,N_28933,N_29817);
nor U31722 (N_31722,N_28210,N_29335);
and U31723 (N_31723,N_28899,N_28727);
nor U31724 (N_31724,N_28629,N_29482);
or U31725 (N_31725,N_28800,N_29988);
nor U31726 (N_31726,N_29065,N_29145);
nor U31727 (N_31727,N_29824,N_28034);
xor U31728 (N_31728,N_28363,N_28772);
or U31729 (N_31729,N_28793,N_28642);
or U31730 (N_31730,N_28823,N_29603);
and U31731 (N_31731,N_29575,N_29762);
xnor U31732 (N_31732,N_27516,N_29094);
nand U31733 (N_31733,N_28525,N_29891);
and U31734 (N_31734,N_29811,N_29703);
xnor U31735 (N_31735,N_29187,N_29191);
nor U31736 (N_31736,N_28511,N_28526);
xor U31737 (N_31737,N_29047,N_29607);
or U31738 (N_31738,N_28937,N_27684);
or U31739 (N_31739,N_28301,N_27539);
nor U31740 (N_31740,N_28456,N_29390);
and U31741 (N_31741,N_28680,N_29493);
or U31742 (N_31742,N_27882,N_29848);
xor U31743 (N_31743,N_28550,N_29471);
xnor U31744 (N_31744,N_29195,N_28951);
or U31745 (N_31745,N_28123,N_27733);
xor U31746 (N_31746,N_29985,N_28060);
nor U31747 (N_31747,N_28225,N_28649);
nor U31748 (N_31748,N_27725,N_28352);
or U31749 (N_31749,N_29725,N_28994);
xnor U31750 (N_31750,N_29160,N_27590);
and U31751 (N_31751,N_27857,N_28969);
and U31752 (N_31752,N_28393,N_28377);
xnor U31753 (N_31753,N_29758,N_28117);
nand U31754 (N_31754,N_29293,N_27977);
nor U31755 (N_31755,N_28037,N_29779);
nand U31756 (N_31756,N_27919,N_28248);
xnor U31757 (N_31757,N_28364,N_29585);
and U31758 (N_31758,N_28016,N_29073);
xnor U31759 (N_31759,N_29544,N_29589);
or U31760 (N_31760,N_27596,N_29267);
xor U31761 (N_31761,N_29876,N_29996);
xor U31762 (N_31762,N_28360,N_29360);
xnor U31763 (N_31763,N_29964,N_29363);
and U31764 (N_31764,N_28332,N_28509);
and U31765 (N_31765,N_29832,N_27596);
nand U31766 (N_31766,N_27618,N_28803);
xnor U31767 (N_31767,N_28390,N_27599);
and U31768 (N_31768,N_29668,N_29309);
nand U31769 (N_31769,N_28656,N_29064);
xnor U31770 (N_31770,N_28977,N_28109);
and U31771 (N_31771,N_29269,N_29780);
or U31772 (N_31772,N_28067,N_28484);
nor U31773 (N_31773,N_29900,N_27544);
nand U31774 (N_31774,N_29633,N_29227);
or U31775 (N_31775,N_27566,N_27685);
xnor U31776 (N_31776,N_29832,N_28388);
nand U31777 (N_31777,N_29246,N_29205);
nand U31778 (N_31778,N_28929,N_28954);
nor U31779 (N_31779,N_29536,N_28646);
or U31780 (N_31780,N_29276,N_29841);
or U31781 (N_31781,N_29634,N_28020);
or U31782 (N_31782,N_27700,N_28460);
xnor U31783 (N_31783,N_28891,N_28642);
and U31784 (N_31784,N_28489,N_29452);
and U31785 (N_31785,N_27895,N_28489);
nand U31786 (N_31786,N_29390,N_28033);
or U31787 (N_31787,N_28902,N_27564);
and U31788 (N_31788,N_27537,N_29073);
and U31789 (N_31789,N_29986,N_29606);
and U31790 (N_31790,N_27502,N_29012);
xor U31791 (N_31791,N_29979,N_27929);
nor U31792 (N_31792,N_28186,N_29791);
or U31793 (N_31793,N_28714,N_27815);
and U31794 (N_31794,N_28448,N_29711);
xor U31795 (N_31795,N_27513,N_28815);
nor U31796 (N_31796,N_28814,N_29124);
xnor U31797 (N_31797,N_28678,N_28030);
xnor U31798 (N_31798,N_29415,N_29802);
or U31799 (N_31799,N_29421,N_28660);
and U31800 (N_31800,N_28415,N_29393);
or U31801 (N_31801,N_27900,N_29659);
xor U31802 (N_31802,N_28635,N_29700);
xor U31803 (N_31803,N_28744,N_29614);
nand U31804 (N_31804,N_28089,N_28982);
or U31805 (N_31805,N_28158,N_28751);
xnor U31806 (N_31806,N_28139,N_28827);
nor U31807 (N_31807,N_29330,N_29668);
and U31808 (N_31808,N_28254,N_28471);
xor U31809 (N_31809,N_29798,N_29286);
nand U31810 (N_31810,N_29682,N_28106);
and U31811 (N_31811,N_27764,N_27942);
or U31812 (N_31812,N_29651,N_28217);
and U31813 (N_31813,N_28313,N_28340);
xnor U31814 (N_31814,N_28204,N_28533);
and U31815 (N_31815,N_29773,N_29917);
nand U31816 (N_31816,N_29099,N_29831);
or U31817 (N_31817,N_29470,N_29866);
or U31818 (N_31818,N_27705,N_29437);
and U31819 (N_31819,N_27526,N_28103);
nor U31820 (N_31820,N_27580,N_29746);
or U31821 (N_31821,N_29065,N_27582);
xnor U31822 (N_31822,N_28451,N_27576);
nand U31823 (N_31823,N_28885,N_28408);
xor U31824 (N_31824,N_27987,N_28881);
and U31825 (N_31825,N_27667,N_28559);
xor U31826 (N_31826,N_28074,N_27875);
and U31827 (N_31827,N_29959,N_28783);
nor U31828 (N_31828,N_29897,N_28658);
xnor U31829 (N_31829,N_29446,N_28969);
or U31830 (N_31830,N_27685,N_28845);
or U31831 (N_31831,N_28894,N_29597);
xnor U31832 (N_31832,N_28787,N_28105);
and U31833 (N_31833,N_29687,N_29276);
and U31834 (N_31834,N_29360,N_27977);
xor U31835 (N_31835,N_28374,N_29274);
xor U31836 (N_31836,N_28691,N_28343);
xnor U31837 (N_31837,N_28740,N_28849);
xor U31838 (N_31838,N_27813,N_29176);
nor U31839 (N_31839,N_29955,N_27970);
or U31840 (N_31840,N_28215,N_28004);
xor U31841 (N_31841,N_28967,N_27628);
nor U31842 (N_31842,N_29410,N_28879);
nand U31843 (N_31843,N_29190,N_28347);
nand U31844 (N_31844,N_28057,N_29738);
or U31845 (N_31845,N_28638,N_27831);
and U31846 (N_31846,N_28769,N_28964);
nor U31847 (N_31847,N_29454,N_29674);
or U31848 (N_31848,N_27646,N_27853);
or U31849 (N_31849,N_28346,N_28391);
and U31850 (N_31850,N_27905,N_29394);
and U31851 (N_31851,N_29064,N_29044);
and U31852 (N_31852,N_29944,N_29086);
xnor U31853 (N_31853,N_29440,N_29757);
and U31854 (N_31854,N_29315,N_29256);
nand U31855 (N_31855,N_29811,N_29786);
xor U31856 (N_31856,N_28076,N_29517);
and U31857 (N_31857,N_29043,N_29069);
nand U31858 (N_31858,N_28345,N_28110);
and U31859 (N_31859,N_29758,N_29129);
nor U31860 (N_31860,N_28462,N_29870);
and U31861 (N_31861,N_29470,N_28372);
nand U31862 (N_31862,N_29129,N_27844);
nor U31863 (N_31863,N_28847,N_29673);
xnor U31864 (N_31864,N_28683,N_29540);
or U31865 (N_31865,N_28900,N_29700);
xnor U31866 (N_31866,N_28894,N_29222);
nor U31867 (N_31867,N_29954,N_27977);
xnor U31868 (N_31868,N_27984,N_29991);
nor U31869 (N_31869,N_28026,N_27754);
nor U31870 (N_31870,N_28852,N_29501);
and U31871 (N_31871,N_28811,N_27785);
nand U31872 (N_31872,N_29426,N_27752);
nand U31873 (N_31873,N_28043,N_29347);
nor U31874 (N_31874,N_29348,N_29297);
nor U31875 (N_31875,N_28855,N_29295);
nor U31876 (N_31876,N_29617,N_29826);
xor U31877 (N_31877,N_29390,N_29844);
and U31878 (N_31878,N_27850,N_29901);
nor U31879 (N_31879,N_28408,N_27538);
and U31880 (N_31880,N_28889,N_29625);
nand U31881 (N_31881,N_29136,N_29899);
xor U31882 (N_31882,N_29067,N_29342);
xor U31883 (N_31883,N_29534,N_28855);
and U31884 (N_31884,N_29335,N_29183);
nor U31885 (N_31885,N_28347,N_29962);
or U31886 (N_31886,N_29429,N_29746);
nor U31887 (N_31887,N_27913,N_29538);
nor U31888 (N_31888,N_28206,N_28813);
or U31889 (N_31889,N_29480,N_28747);
or U31890 (N_31890,N_28707,N_28979);
nor U31891 (N_31891,N_27926,N_29110);
xnor U31892 (N_31892,N_28055,N_28254);
xor U31893 (N_31893,N_27686,N_28331);
and U31894 (N_31894,N_29452,N_29496);
xnor U31895 (N_31895,N_28339,N_29865);
nand U31896 (N_31896,N_28786,N_29957);
nand U31897 (N_31897,N_29875,N_28825);
nor U31898 (N_31898,N_28358,N_28573);
or U31899 (N_31899,N_27972,N_29997);
or U31900 (N_31900,N_29764,N_29131);
xnor U31901 (N_31901,N_27974,N_29474);
or U31902 (N_31902,N_28536,N_29586);
xor U31903 (N_31903,N_28883,N_28634);
and U31904 (N_31904,N_27532,N_29007);
nor U31905 (N_31905,N_28577,N_29088);
xnor U31906 (N_31906,N_29597,N_28039);
and U31907 (N_31907,N_29394,N_29133);
or U31908 (N_31908,N_28930,N_29244);
nand U31909 (N_31909,N_29452,N_29823);
and U31910 (N_31910,N_29855,N_29755);
or U31911 (N_31911,N_29746,N_29709);
or U31912 (N_31912,N_29399,N_29617);
or U31913 (N_31913,N_29705,N_29105);
nand U31914 (N_31914,N_27950,N_29171);
nor U31915 (N_31915,N_29789,N_28694);
xor U31916 (N_31916,N_28244,N_28001);
nor U31917 (N_31917,N_28111,N_27961);
or U31918 (N_31918,N_29572,N_29671);
and U31919 (N_31919,N_29589,N_28793);
or U31920 (N_31920,N_29050,N_28615);
nor U31921 (N_31921,N_28764,N_28721);
xnor U31922 (N_31922,N_29284,N_29112);
or U31923 (N_31923,N_27558,N_29420);
or U31924 (N_31924,N_29405,N_28867);
nand U31925 (N_31925,N_28983,N_29530);
and U31926 (N_31926,N_28824,N_28633);
nor U31927 (N_31927,N_29557,N_29538);
nor U31928 (N_31928,N_29753,N_28460);
nor U31929 (N_31929,N_27868,N_28922);
and U31930 (N_31930,N_28442,N_28028);
or U31931 (N_31931,N_29689,N_27649);
nor U31932 (N_31932,N_28552,N_28003);
and U31933 (N_31933,N_28752,N_29367);
and U31934 (N_31934,N_29535,N_27538);
and U31935 (N_31935,N_28263,N_29703);
or U31936 (N_31936,N_29539,N_28002);
nor U31937 (N_31937,N_27551,N_28649);
nor U31938 (N_31938,N_28775,N_29052);
and U31939 (N_31939,N_29935,N_27679);
xnor U31940 (N_31940,N_29393,N_29339);
and U31941 (N_31941,N_29297,N_28890);
xor U31942 (N_31942,N_27602,N_28212);
or U31943 (N_31943,N_29585,N_27766);
or U31944 (N_31944,N_27707,N_29916);
nor U31945 (N_31945,N_28512,N_28250);
or U31946 (N_31946,N_27861,N_28572);
nand U31947 (N_31947,N_28603,N_29790);
or U31948 (N_31948,N_29074,N_29145);
nor U31949 (N_31949,N_28269,N_29534);
or U31950 (N_31950,N_28954,N_29697);
and U31951 (N_31951,N_28555,N_28143);
and U31952 (N_31952,N_29575,N_29200);
nor U31953 (N_31953,N_28605,N_27546);
nor U31954 (N_31954,N_28673,N_28544);
or U31955 (N_31955,N_28249,N_29946);
or U31956 (N_31956,N_27566,N_28659);
xnor U31957 (N_31957,N_27571,N_29117);
or U31958 (N_31958,N_29624,N_29935);
and U31959 (N_31959,N_29763,N_29558);
nor U31960 (N_31960,N_29723,N_27957);
xor U31961 (N_31961,N_27632,N_29826);
and U31962 (N_31962,N_28059,N_29845);
nand U31963 (N_31963,N_29340,N_29593);
xnor U31964 (N_31964,N_29065,N_28496);
nand U31965 (N_31965,N_29042,N_27573);
nor U31966 (N_31966,N_28944,N_29320);
and U31967 (N_31967,N_29901,N_29366);
or U31968 (N_31968,N_28427,N_29494);
and U31969 (N_31969,N_28736,N_29975);
xnor U31970 (N_31970,N_28031,N_29182);
or U31971 (N_31971,N_28258,N_28680);
xor U31972 (N_31972,N_29722,N_28646);
xor U31973 (N_31973,N_29726,N_29446);
nor U31974 (N_31974,N_29614,N_29260);
xor U31975 (N_31975,N_29661,N_27851);
nor U31976 (N_31976,N_29435,N_28686);
xnor U31977 (N_31977,N_29236,N_28306);
nand U31978 (N_31978,N_29722,N_27718);
and U31979 (N_31979,N_29795,N_28322);
nor U31980 (N_31980,N_29033,N_27722);
nand U31981 (N_31981,N_28262,N_28050);
and U31982 (N_31982,N_29755,N_29878);
and U31983 (N_31983,N_28266,N_28739);
nor U31984 (N_31984,N_28057,N_27938);
nor U31985 (N_31985,N_27712,N_27522);
nand U31986 (N_31986,N_28762,N_27812);
nor U31987 (N_31987,N_27881,N_28872);
nand U31988 (N_31988,N_29170,N_28693);
xnor U31989 (N_31989,N_27634,N_28120);
xnor U31990 (N_31990,N_28588,N_29513);
xnor U31991 (N_31991,N_28471,N_28238);
and U31992 (N_31992,N_27825,N_28276);
nand U31993 (N_31993,N_29670,N_29096);
or U31994 (N_31994,N_27762,N_29530);
nor U31995 (N_31995,N_27737,N_28941);
xor U31996 (N_31996,N_29912,N_29436);
or U31997 (N_31997,N_29723,N_28655);
nand U31998 (N_31998,N_27952,N_29754);
or U31999 (N_31999,N_28411,N_28127);
nand U32000 (N_32000,N_28202,N_28017);
and U32001 (N_32001,N_28169,N_29691);
xor U32002 (N_32002,N_28002,N_27822);
and U32003 (N_32003,N_27607,N_29205);
xnor U32004 (N_32004,N_28479,N_28913);
nor U32005 (N_32005,N_28625,N_27722);
xor U32006 (N_32006,N_29028,N_29663);
and U32007 (N_32007,N_29263,N_28580);
nor U32008 (N_32008,N_28712,N_27969);
or U32009 (N_32009,N_28205,N_29555);
nand U32010 (N_32010,N_28072,N_28496);
nor U32011 (N_32011,N_28037,N_29255);
or U32012 (N_32012,N_29647,N_28722);
nand U32013 (N_32013,N_29910,N_27679);
nor U32014 (N_32014,N_29286,N_28258);
xnor U32015 (N_32015,N_28194,N_28257);
or U32016 (N_32016,N_28206,N_29801);
or U32017 (N_32017,N_27922,N_29013);
or U32018 (N_32018,N_27552,N_28688);
and U32019 (N_32019,N_27809,N_29420);
nor U32020 (N_32020,N_29796,N_28862);
and U32021 (N_32021,N_27794,N_27559);
nand U32022 (N_32022,N_28324,N_29543);
xnor U32023 (N_32023,N_29763,N_28485);
and U32024 (N_32024,N_29736,N_29841);
xnor U32025 (N_32025,N_28357,N_29512);
nand U32026 (N_32026,N_29090,N_29622);
and U32027 (N_32027,N_27832,N_29975);
and U32028 (N_32028,N_29801,N_29504);
and U32029 (N_32029,N_28375,N_28540);
and U32030 (N_32030,N_27725,N_27588);
and U32031 (N_32031,N_29879,N_29586);
nand U32032 (N_32032,N_29766,N_28381);
nor U32033 (N_32033,N_29970,N_28864);
nand U32034 (N_32034,N_29703,N_29087);
and U32035 (N_32035,N_28314,N_28534);
nor U32036 (N_32036,N_29790,N_27759);
xor U32037 (N_32037,N_27598,N_28389);
and U32038 (N_32038,N_29210,N_27526);
and U32039 (N_32039,N_27914,N_28068);
nand U32040 (N_32040,N_29499,N_27801);
nand U32041 (N_32041,N_28628,N_28059);
and U32042 (N_32042,N_28954,N_29726);
and U32043 (N_32043,N_29048,N_29662);
nor U32044 (N_32044,N_27781,N_27667);
nand U32045 (N_32045,N_28778,N_28249);
nand U32046 (N_32046,N_28418,N_27832);
or U32047 (N_32047,N_29967,N_29407);
nor U32048 (N_32048,N_28271,N_28840);
nand U32049 (N_32049,N_28836,N_29884);
nor U32050 (N_32050,N_29050,N_29442);
xnor U32051 (N_32051,N_28985,N_29759);
xor U32052 (N_32052,N_29910,N_29279);
or U32053 (N_32053,N_27513,N_27795);
and U32054 (N_32054,N_28960,N_28635);
nor U32055 (N_32055,N_27783,N_29360);
and U32056 (N_32056,N_29425,N_29719);
or U32057 (N_32057,N_27639,N_28735);
nand U32058 (N_32058,N_28317,N_27861);
and U32059 (N_32059,N_27614,N_27992);
nor U32060 (N_32060,N_29971,N_28076);
nor U32061 (N_32061,N_28365,N_28480);
nor U32062 (N_32062,N_28811,N_29172);
xor U32063 (N_32063,N_29815,N_28937);
or U32064 (N_32064,N_28396,N_28029);
nand U32065 (N_32065,N_29489,N_28556);
or U32066 (N_32066,N_28602,N_29232);
nand U32067 (N_32067,N_28710,N_28513);
nand U32068 (N_32068,N_29739,N_28109);
or U32069 (N_32069,N_29740,N_27984);
and U32070 (N_32070,N_29254,N_29859);
nor U32071 (N_32071,N_28495,N_29454);
or U32072 (N_32072,N_27762,N_29130);
nor U32073 (N_32073,N_28772,N_28277);
xor U32074 (N_32074,N_29794,N_28765);
and U32075 (N_32075,N_28111,N_28698);
nand U32076 (N_32076,N_28802,N_28368);
and U32077 (N_32077,N_28800,N_27908);
and U32078 (N_32078,N_29330,N_29891);
nor U32079 (N_32079,N_29769,N_29241);
nor U32080 (N_32080,N_28792,N_29091);
nand U32081 (N_32081,N_29318,N_28901);
nor U32082 (N_32082,N_28222,N_29680);
and U32083 (N_32083,N_28155,N_27557);
and U32084 (N_32084,N_28675,N_28733);
and U32085 (N_32085,N_28157,N_28449);
xor U32086 (N_32086,N_29761,N_27749);
and U32087 (N_32087,N_29550,N_28083);
or U32088 (N_32088,N_28477,N_29437);
xor U32089 (N_32089,N_29901,N_29355);
or U32090 (N_32090,N_28307,N_28512);
nor U32091 (N_32091,N_29498,N_27786);
nand U32092 (N_32092,N_27642,N_27911);
or U32093 (N_32093,N_29759,N_29341);
and U32094 (N_32094,N_28347,N_28027);
or U32095 (N_32095,N_28227,N_28486);
nand U32096 (N_32096,N_28774,N_27580);
nor U32097 (N_32097,N_28929,N_28670);
nor U32098 (N_32098,N_27960,N_29821);
and U32099 (N_32099,N_28790,N_28809);
and U32100 (N_32100,N_29558,N_28325);
nor U32101 (N_32101,N_28896,N_28361);
or U32102 (N_32102,N_29611,N_28051);
xnor U32103 (N_32103,N_28239,N_27613);
nor U32104 (N_32104,N_28705,N_28569);
or U32105 (N_32105,N_28622,N_29305);
and U32106 (N_32106,N_29337,N_27964);
nand U32107 (N_32107,N_29791,N_28904);
nand U32108 (N_32108,N_29994,N_27780);
xnor U32109 (N_32109,N_28009,N_29025);
or U32110 (N_32110,N_29688,N_28495);
xor U32111 (N_32111,N_27717,N_28553);
nor U32112 (N_32112,N_29530,N_27544);
xnor U32113 (N_32113,N_29228,N_28780);
or U32114 (N_32114,N_29144,N_29463);
nand U32115 (N_32115,N_28165,N_28936);
or U32116 (N_32116,N_29503,N_27519);
nand U32117 (N_32117,N_27697,N_29164);
nor U32118 (N_32118,N_29290,N_28435);
or U32119 (N_32119,N_27648,N_29604);
and U32120 (N_32120,N_27847,N_29485);
nand U32121 (N_32121,N_27984,N_29806);
xor U32122 (N_32122,N_28101,N_29396);
or U32123 (N_32123,N_28292,N_29760);
nor U32124 (N_32124,N_27991,N_28049);
and U32125 (N_32125,N_28063,N_28169);
nor U32126 (N_32126,N_27625,N_29883);
nand U32127 (N_32127,N_29132,N_29792);
or U32128 (N_32128,N_28888,N_28831);
and U32129 (N_32129,N_29777,N_29956);
or U32130 (N_32130,N_27540,N_29038);
nand U32131 (N_32131,N_27835,N_28230);
nor U32132 (N_32132,N_29520,N_29246);
xor U32133 (N_32133,N_28484,N_28040);
or U32134 (N_32134,N_27969,N_27581);
and U32135 (N_32135,N_27856,N_29675);
nand U32136 (N_32136,N_29822,N_29240);
nor U32137 (N_32137,N_29756,N_29815);
and U32138 (N_32138,N_29005,N_27729);
and U32139 (N_32139,N_29884,N_28037);
nor U32140 (N_32140,N_28375,N_28137);
and U32141 (N_32141,N_27697,N_29393);
xor U32142 (N_32142,N_27884,N_28586);
or U32143 (N_32143,N_27660,N_28610);
xnor U32144 (N_32144,N_28022,N_28639);
nand U32145 (N_32145,N_29770,N_29317);
and U32146 (N_32146,N_28484,N_29727);
nor U32147 (N_32147,N_29596,N_28361);
nand U32148 (N_32148,N_28339,N_28160);
nand U32149 (N_32149,N_27926,N_29759);
nand U32150 (N_32150,N_27957,N_28189);
nand U32151 (N_32151,N_29929,N_27953);
and U32152 (N_32152,N_29695,N_29444);
or U32153 (N_32153,N_28351,N_28265);
nor U32154 (N_32154,N_28955,N_28982);
or U32155 (N_32155,N_29970,N_29565);
and U32156 (N_32156,N_27857,N_29722);
nor U32157 (N_32157,N_28273,N_29047);
or U32158 (N_32158,N_29093,N_27591);
nand U32159 (N_32159,N_29271,N_27542);
nand U32160 (N_32160,N_28921,N_27564);
or U32161 (N_32161,N_29676,N_29929);
nand U32162 (N_32162,N_27837,N_27984);
or U32163 (N_32163,N_29667,N_28244);
nor U32164 (N_32164,N_29507,N_29370);
and U32165 (N_32165,N_28676,N_28942);
nor U32166 (N_32166,N_29667,N_29560);
and U32167 (N_32167,N_28066,N_29071);
or U32168 (N_32168,N_27677,N_29542);
nor U32169 (N_32169,N_29959,N_28957);
or U32170 (N_32170,N_28376,N_29257);
and U32171 (N_32171,N_28640,N_29894);
nand U32172 (N_32172,N_29683,N_28194);
or U32173 (N_32173,N_27544,N_27503);
or U32174 (N_32174,N_27659,N_28568);
nand U32175 (N_32175,N_27999,N_28854);
xnor U32176 (N_32176,N_28679,N_28058);
or U32177 (N_32177,N_29740,N_28092);
and U32178 (N_32178,N_29154,N_29655);
nor U32179 (N_32179,N_29271,N_27840);
xor U32180 (N_32180,N_28715,N_29473);
and U32181 (N_32181,N_27645,N_28740);
nand U32182 (N_32182,N_28633,N_28645);
and U32183 (N_32183,N_27543,N_28102);
xnor U32184 (N_32184,N_29849,N_28626);
or U32185 (N_32185,N_29112,N_29697);
or U32186 (N_32186,N_28076,N_29415);
nor U32187 (N_32187,N_28128,N_27783);
and U32188 (N_32188,N_29537,N_28084);
and U32189 (N_32189,N_27768,N_29375);
and U32190 (N_32190,N_27537,N_28157);
nor U32191 (N_32191,N_29568,N_28303);
xnor U32192 (N_32192,N_29128,N_28827);
or U32193 (N_32193,N_28526,N_29461);
xor U32194 (N_32194,N_28014,N_28052);
nand U32195 (N_32195,N_29268,N_28644);
nand U32196 (N_32196,N_29401,N_29682);
nor U32197 (N_32197,N_29867,N_28255);
xor U32198 (N_32198,N_28672,N_29122);
xnor U32199 (N_32199,N_28512,N_27623);
xor U32200 (N_32200,N_28766,N_29324);
nor U32201 (N_32201,N_28964,N_29260);
nor U32202 (N_32202,N_27677,N_28899);
nor U32203 (N_32203,N_28381,N_28963);
and U32204 (N_32204,N_28527,N_27999);
and U32205 (N_32205,N_29448,N_27655);
nand U32206 (N_32206,N_28185,N_29556);
and U32207 (N_32207,N_28866,N_29321);
xor U32208 (N_32208,N_28901,N_28395);
nand U32209 (N_32209,N_28285,N_27611);
and U32210 (N_32210,N_27938,N_29237);
nand U32211 (N_32211,N_29791,N_29362);
and U32212 (N_32212,N_29642,N_29982);
and U32213 (N_32213,N_29602,N_29437);
or U32214 (N_32214,N_28613,N_27521);
and U32215 (N_32215,N_29750,N_29801);
nor U32216 (N_32216,N_28409,N_28489);
nor U32217 (N_32217,N_29719,N_28120);
or U32218 (N_32218,N_29026,N_29340);
nand U32219 (N_32219,N_28979,N_27862);
or U32220 (N_32220,N_29820,N_28423);
xnor U32221 (N_32221,N_29300,N_28965);
xnor U32222 (N_32222,N_27882,N_27792);
nand U32223 (N_32223,N_29723,N_27578);
nand U32224 (N_32224,N_27973,N_27974);
nand U32225 (N_32225,N_27614,N_28305);
or U32226 (N_32226,N_28195,N_28514);
nor U32227 (N_32227,N_29798,N_29360);
nand U32228 (N_32228,N_28568,N_28343);
xor U32229 (N_32229,N_29511,N_27594);
or U32230 (N_32230,N_28267,N_29471);
and U32231 (N_32231,N_27948,N_28308);
or U32232 (N_32232,N_29694,N_27653);
and U32233 (N_32233,N_29900,N_28800);
nor U32234 (N_32234,N_29567,N_29592);
nor U32235 (N_32235,N_27968,N_29320);
and U32236 (N_32236,N_29442,N_27619);
or U32237 (N_32237,N_29693,N_29055);
xor U32238 (N_32238,N_29635,N_29929);
or U32239 (N_32239,N_29394,N_28265);
or U32240 (N_32240,N_29849,N_27810);
nand U32241 (N_32241,N_28117,N_27610);
or U32242 (N_32242,N_28734,N_28869);
nand U32243 (N_32243,N_28236,N_29148);
nor U32244 (N_32244,N_29847,N_29079);
xnor U32245 (N_32245,N_27625,N_28567);
or U32246 (N_32246,N_27660,N_28754);
nand U32247 (N_32247,N_29584,N_29414);
xnor U32248 (N_32248,N_28500,N_29630);
nand U32249 (N_32249,N_27544,N_29360);
xor U32250 (N_32250,N_29597,N_29607);
xnor U32251 (N_32251,N_27552,N_27593);
nor U32252 (N_32252,N_28607,N_29833);
and U32253 (N_32253,N_27584,N_27621);
and U32254 (N_32254,N_29067,N_28697);
xnor U32255 (N_32255,N_29285,N_28372);
nor U32256 (N_32256,N_29734,N_29808);
nand U32257 (N_32257,N_29620,N_28969);
or U32258 (N_32258,N_29984,N_28965);
xnor U32259 (N_32259,N_29251,N_29476);
and U32260 (N_32260,N_29685,N_29775);
and U32261 (N_32261,N_29511,N_29173);
xor U32262 (N_32262,N_27650,N_29525);
nor U32263 (N_32263,N_29345,N_27998);
xnor U32264 (N_32264,N_29026,N_29363);
nor U32265 (N_32265,N_28916,N_29019);
or U32266 (N_32266,N_27926,N_29189);
xnor U32267 (N_32267,N_27782,N_28882);
xor U32268 (N_32268,N_29160,N_29643);
nand U32269 (N_32269,N_29721,N_28139);
nor U32270 (N_32270,N_28995,N_28229);
xor U32271 (N_32271,N_28681,N_28927);
xor U32272 (N_32272,N_28573,N_29335);
and U32273 (N_32273,N_29158,N_29555);
nor U32274 (N_32274,N_28653,N_27512);
xnor U32275 (N_32275,N_27580,N_27848);
xnor U32276 (N_32276,N_29066,N_29908);
or U32277 (N_32277,N_28126,N_28079);
nor U32278 (N_32278,N_29787,N_28684);
or U32279 (N_32279,N_27529,N_28105);
nand U32280 (N_32280,N_29611,N_28232);
xor U32281 (N_32281,N_27866,N_27580);
nand U32282 (N_32282,N_28418,N_28433);
nand U32283 (N_32283,N_29191,N_28667);
nor U32284 (N_32284,N_29055,N_27784);
or U32285 (N_32285,N_29788,N_27551);
xor U32286 (N_32286,N_28796,N_28772);
nand U32287 (N_32287,N_28205,N_28461);
nor U32288 (N_32288,N_29493,N_28581);
nand U32289 (N_32289,N_29485,N_28522);
nor U32290 (N_32290,N_27849,N_29056);
nand U32291 (N_32291,N_28639,N_28717);
xnor U32292 (N_32292,N_29323,N_27803);
nand U32293 (N_32293,N_29756,N_27537);
and U32294 (N_32294,N_28661,N_29337);
nor U32295 (N_32295,N_29899,N_28066);
or U32296 (N_32296,N_28097,N_29893);
or U32297 (N_32297,N_29757,N_28390);
or U32298 (N_32298,N_28179,N_29169);
or U32299 (N_32299,N_29711,N_27661);
or U32300 (N_32300,N_27860,N_29584);
nand U32301 (N_32301,N_29783,N_28980);
nor U32302 (N_32302,N_28917,N_28592);
nand U32303 (N_32303,N_29786,N_28033);
nand U32304 (N_32304,N_28911,N_29803);
nand U32305 (N_32305,N_28449,N_28729);
or U32306 (N_32306,N_28126,N_28584);
nor U32307 (N_32307,N_27814,N_27980);
and U32308 (N_32308,N_27906,N_28192);
or U32309 (N_32309,N_29336,N_29495);
nand U32310 (N_32310,N_28403,N_28574);
nor U32311 (N_32311,N_28380,N_28069);
nand U32312 (N_32312,N_29069,N_28403);
nor U32313 (N_32313,N_28536,N_27818);
xnor U32314 (N_32314,N_27641,N_29166);
xnor U32315 (N_32315,N_29316,N_28701);
nand U32316 (N_32316,N_28289,N_29384);
nand U32317 (N_32317,N_29521,N_29922);
nor U32318 (N_32318,N_28420,N_29716);
xnor U32319 (N_32319,N_28389,N_28721);
nor U32320 (N_32320,N_29825,N_28389);
nand U32321 (N_32321,N_27845,N_28279);
or U32322 (N_32322,N_28653,N_27875);
xor U32323 (N_32323,N_29367,N_29501);
or U32324 (N_32324,N_28331,N_29790);
xnor U32325 (N_32325,N_29910,N_29021);
nand U32326 (N_32326,N_27955,N_28026);
nand U32327 (N_32327,N_28829,N_28297);
and U32328 (N_32328,N_29420,N_29871);
or U32329 (N_32329,N_29004,N_28637);
nor U32330 (N_32330,N_29388,N_29159);
and U32331 (N_32331,N_28690,N_27859);
xnor U32332 (N_32332,N_28057,N_28704);
or U32333 (N_32333,N_27630,N_29627);
xor U32334 (N_32334,N_29557,N_28843);
or U32335 (N_32335,N_28951,N_29623);
xor U32336 (N_32336,N_28715,N_29648);
nand U32337 (N_32337,N_28007,N_28184);
nor U32338 (N_32338,N_29579,N_29952);
and U32339 (N_32339,N_29224,N_28005);
xnor U32340 (N_32340,N_29985,N_28591);
and U32341 (N_32341,N_29482,N_27503);
nand U32342 (N_32342,N_29058,N_29100);
and U32343 (N_32343,N_28616,N_29980);
or U32344 (N_32344,N_29252,N_28228);
nand U32345 (N_32345,N_29537,N_27820);
nor U32346 (N_32346,N_29457,N_29887);
or U32347 (N_32347,N_27618,N_28012);
nand U32348 (N_32348,N_29197,N_29038);
nand U32349 (N_32349,N_27724,N_28235);
and U32350 (N_32350,N_29641,N_29974);
xnor U32351 (N_32351,N_27740,N_28916);
or U32352 (N_32352,N_29813,N_29459);
nor U32353 (N_32353,N_28505,N_29126);
xor U32354 (N_32354,N_29232,N_29195);
and U32355 (N_32355,N_28949,N_29764);
xnor U32356 (N_32356,N_28926,N_28616);
nand U32357 (N_32357,N_29277,N_28538);
and U32358 (N_32358,N_28295,N_28877);
nand U32359 (N_32359,N_29105,N_27734);
or U32360 (N_32360,N_27603,N_28126);
and U32361 (N_32361,N_28422,N_28162);
nor U32362 (N_32362,N_27694,N_29774);
nand U32363 (N_32363,N_29942,N_28647);
and U32364 (N_32364,N_29970,N_29478);
or U32365 (N_32365,N_28809,N_28770);
xor U32366 (N_32366,N_29319,N_28525);
nor U32367 (N_32367,N_29869,N_27960);
and U32368 (N_32368,N_28830,N_29632);
or U32369 (N_32369,N_29630,N_29890);
and U32370 (N_32370,N_29557,N_28407);
or U32371 (N_32371,N_29880,N_29939);
nand U32372 (N_32372,N_28898,N_28725);
xnor U32373 (N_32373,N_29742,N_28724);
nand U32374 (N_32374,N_29636,N_27589);
and U32375 (N_32375,N_29278,N_27761);
nand U32376 (N_32376,N_29407,N_29530);
nand U32377 (N_32377,N_27667,N_29666);
nor U32378 (N_32378,N_27719,N_27762);
xor U32379 (N_32379,N_28444,N_29723);
nor U32380 (N_32380,N_29978,N_28753);
and U32381 (N_32381,N_27764,N_27792);
xnor U32382 (N_32382,N_28029,N_29887);
or U32383 (N_32383,N_29375,N_27669);
xnor U32384 (N_32384,N_29322,N_29928);
xor U32385 (N_32385,N_28814,N_27849);
nor U32386 (N_32386,N_27760,N_27893);
and U32387 (N_32387,N_27933,N_28760);
xor U32388 (N_32388,N_29189,N_28245);
nand U32389 (N_32389,N_28875,N_27545);
xor U32390 (N_32390,N_29484,N_28732);
or U32391 (N_32391,N_27586,N_29295);
and U32392 (N_32392,N_28347,N_29966);
xor U32393 (N_32393,N_27934,N_29590);
xor U32394 (N_32394,N_29142,N_28009);
and U32395 (N_32395,N_29332,N_29126);
xnor U32396 (N_32396,N_27813,N_29965);
and U32397 (N_32397,N_28571,N_29335);
and U32398 (N_32398,N_29538,N_28098);
nor U32399 (N_32399,N_29803,N_29856);
or U32400 (N_32400,N_27705,N_28215);
and U32401 (N_32401,N_27967,N_29043);
and U32402 (N_32402,N_29945,N_29873);
nor U32403 (N_32403,N_28754,N_28497);
and U32404 (N_32404,N_27866,N_28018);
xnor U32405 (N_32405,N_29902,N_28608);
xor U32406 (N_32406,N_28568,N_28862);
nand U32407 (N_32407,N_27767,N_29218);
xor U32408 (N_32408,N_28444,N_28341);
nor U32409 (N_32409,N_28298,N_27684);
or U32410 (N_32410,N_28672,N_29912);
and U32411 (N_32411,N_28620,N_28379);
xnor U32412 (N_32412,N_27525,N_28768);
nor U32413 (N_32413,N_29196,N_29833);
nand U32414 (N_32414,N_29574,N_29632);
xor U32415 (N_32415,N_29660,N_29946);
nor U32416 (N_32416,N_28900,N_28341);
xor U32417 (N_32417,N_28492,N_29274);
xnor U32418 (N_32418,N_28762,N_28223);
or U32419 (N_32419,N_29301,N_27504);
xnor U32420 (N_32420,N_29422,N_29525);
nand U32421 (N_32421,N_29313,N_29801);
nor U32422 (N_32422,N_28054,N_29610);
xnor U32423 (N_32423,N_28241,N_28875);
and U32424 (N_32424,N_28700,N_28577);
nand U32425 (N_32425,N_29260,N_29500);
nor U32426 (N_32426,N_28304,N_28021);
xor U32427 (N_32427,N_27663,N_28286);
nor U32428 (N_32428,N_29513,N_27663);
or U32429 (N_32429,N_28242,N_28461);
or U32430 (N_32430,N_28989,N_29669);
xor U32431 (N_32431,N_29879,N_29259);
and U32432 (N_32432,N_28134,N_29936);
or U32433 (N_32433,N_29822,N_29812);
nand U32434 (N_32434,N_28307,N_28302);
or U32435 (N_32435,N_29895,N_29497);
xnor U32436 (N_32436,N_29029,N_27941);
or U32437 (N_32437,N_29854,N_29518);
and U32438 (N_32438,N_27713,N_28996);
nor U32439 (N_32439,N_27526,N_27949);
or U32440 (N_32440,N_27895,N_29852);
or U32441 (N_32441,N_27971,N_28186);
or U32442 (N_32442,N_28443,N_27749);
or U32443 (N_32443,N_27651,N_28515);
and U32444 (N_32444,N_28748,N_28606);
nor U32445 (N_32445,N_27698,N_29530);
or U32446 (N_32446,N_29933,N_28504);
or U32447 (N_32447,N_27975,N_28179);
nor U32448 (N_32448,N_28187,N_28627);
nor U32449 (N_32449,N_29360,N_28584);
or U32450 (N_32450,N_27585,N_28176);
or U32451 (N_32451,N_29930,N_29636);
nand U32452 (N_32452,N_28438,N_29393);
or U32453 (N_32453,N_27799,N_28763);
nor U32454 (N_32454,N_28204,N_27561);
nand U32455 (N_32455,N_29669,N_29090);
xnor U32456 (N_32456,N_28545,N_29417);
xnor U32457 (N_32457,N_27750,N_28573);
nor U32458 (N_32458,N_29268,N_28766);
or U32459 (N_32459,N_28175,N_29240);
and U32460 (N_32460,N_29672,N_28559);
xnor U32461 (N_32461,N_29361,N_29376);
nand U32462 (N_32462,N_27634,N_29059);
nor U32463 (N_32463,N_27710,N_29118);
nor U32464 (N_32464,N_28871,N_29882);
or U32465 (N_32465,N_27610,N_27793);
or U32466 (N_32466,N_27716,N_29647);
xnor U32467 (N_32467,N_28460,N_27614);
and U32468 (N_32468,N_28488,N_27695);
nor U32469 (N_32469,N_28695,N_28685);
nor U32470 (N_32470,N_28952,N_28208);
or U32471 (N_32471,N_29998,N_28548);
nor U32472 (N_32472,N_29570,N_28719);
nand U32473 (N_32473,N_29282,N_29705);
nand U32474 (N_32474,N_29567,N_29163);
and U32475 (N_32475,N_28210,N_27900);
and U32476 (N_32476,N_28677,N_27755);
xor U32477 (N_32477,N_29193,N_29758);
and U32478 (N_32478,N_29251,N_29852);
xnor U32479 (N_32479,N_29954,N_29008);
and U32480 (N_32480,N_29361,N_27985);
or U32481 (N_32481,N_29747,N_29596);
or U32482 (N_32482,N_28812,N_29716);
nand U32483 (N_32483,N_29683,N_29120);
nand U32484 (N_32484,N_28873,N_28221);
xnor U32485 (N_32485,N_28576,N_28625);
nand U32486 (N_32486,N_28488,N_28010);
nor U32487 (N_32487,N_29039,N_28058);
nand U32488 (N_32488,N_29156,N_27648);
xnor U32489 (N_32489,N_28248,N_29053);
xor U32490 (N_32490,N_29028,N_27614);
xnor U32491 (N_32491,N_28274,N_28985);
and U32492 (N_32492,N_28303,N_29025);
and U32493 (N_32493,N_27828,N_29973);
or U32494 (N_32494,N_27924,N_29656);
and U32495 (N_32495,N_28566,N_29231);
and U32496 (N_32496,N_28231,N_28669);
xor U32497 (N_32497,N_29121,N_27789);
and U32498 (N_32498,N_28551,N_29365);
and U32499 (N_32499,N_28475,N_29842);
nor U32500 (N_32500,N_31808,N_30930);
nand U32501 (N_32501,N_30647,N_31157);
and U32502 (N_32502,N_30623,N_32438);
nor U32503 (N_32503,N_30192,N_31256);
nor U32504 (N_32504,N_30935,N_30860);
xor U32505 (N_32505,N_32091,N_31998);
nor U32506 (N_32506,N_30887,N_30363);
nor U32507 (N_32507,N_30581,N_32492);
nand U32508 (N_32508,N_31300,N_31355);
nor U32509 (N_32509,N_31342,N_31446);
nand U32510 (N_32510,N_30524,N_30520);
and U32511 (N_32511,N_30678,N_31559);
xnor U32512 (N_32512,N_31877,N_30196);
nand U32513 (N_32513,N_32055,N_32078);
nand U32514 (N_32514,N_31409,N_30869);
and U32515 (N_32515,N_31085,N_32083);
nand U32516 (N_32516,N_30364,N_31201);
and U32517 (N_32517,N_30531,N_30644);
nor U32518 (N_32518,N_31687,N_30304);
nor U32519 (N_32519,N_31140,N_31326);
or U32520 (N_32520,N_31681,N_31434);
nor U32521 (N_32521,N_30573,N_31141);
and U32522 (N_32522,N_30455,N_30692);
and U32523 (N_32523,N_31927,N_30037);
nor U32524 (N_32524,N_31031,N_32307);
or U32525 (N_32525,N_32139,N_31814);
xnor U32526 (N_32526,N_31054,N_30579);
or U32527 (N_32527,N_31796,N_31734);
nand U32528 (N_32528,N_31873,N_30297);
nor U32529 (N_32529,N_32272,N_31209);
or U32530 (N_32530,N_30981,N_30092);
or U32531 (N_32531,N_31632,N_31875);
nand U32532 (N_32532,N_30208,N_31255);
nand U32533 (N_32533,N_30239,N_30976);
xor U32534 (N_32534,N_32169,N_31723);
and U32535 (N_32535,N_31106,N_30228);
or U32536 (N_32536,N_30096,N_32453);
nor U32537 (N_32537,N_32440,N_31672);
and U32538 (N_32538,N_31414,N_31533);
nand U32539 (N_32539,N_31668,N_32403);
xnor U32540 (N_32540,N_30314,N_31306);
xnor U32541 (N_32541,N_31768,N_32327);
and U32542 (N_32542,N_31464,N_30937);
nor U32543 (N_32543,N_30979,N_32496);
or U32544 (N_32544,N_32431,N_30511);
and U32545 (N_32545,N_32491,N_32464);
nor U32546 (N_32546,N_31882,N_30370);
xor U32547 (N_32547,N_31562,N_32424);
nand U32548 (N_32548,N_30767,N_32472);
nand U32549 (N_32549,N_30257,N_32216);
and U32550 (N_32550,N_32398,N_30823);
nand U32551 (N_32551,N_30419,N_31199);
xor U32552 (N_32552,N_30048,N_30266);
xor U32553 (N_32553,N_31754,N_30832);
and U32554 (N_32554,N_32456,N_31457);
nand U32555 (N_32555,N_31631,N_31805);
nor U32556 (N_32556,N_30540,N_30568);
or U32557 (N_32557,N_31893,N_31978);
and U32558 (N_32558,N_30260,N_31293);
or U32559 (N_32559,N_32392,N_30378);
and U32560 (N_32560,N_30781,N_32136);
and U32561 (N_32561,N_32474,N_32363);
xor U32562 (N_32562,N_30900,N_30888);
nor U32563 (N_32563,N_31186,N_31586);
xor U32564 (N_32564,N_31712,N_30576);
xor U32565 (N_32565,N_30843,N_30152);
and U32566 (N_32566,N_32231,N_30677);
or U32567 (N_32567,N_30151,N_30845);
or U32568 (N_32568,N_32079,N_30502);
or U32569 (N_32569,N_32206,N_31462);
and U32570 (N_32570,N_31541,N_30599);
and U32571 (N_32571,N_31968,N_31705);
nor U32572 (N_32572,N_31155,N_30594);
and U32573 (N_32573,N_30912,N_30470);
and U32574 (N_32574,N_31384,N_31400);
nand U32575 (N_32575,N_31390,N_30063);
and U32576 (N_32576,N_30654,N_31799);
nor U32577 (N_32577,N_30789,N_30414);
nor U32578 (N_32578,N_32160,N_31469);
or U32579 (N_32579,N_30244,N_30880);
nand U32580 (N_32580,N_30727,N_30309);
xnor U32581 (N_32581,N_32113,N_30839);
or U32582 (N_32582,N_31424,N_30634);
nor U32583 (N_32583,N_30911,N_31718);
xnor U32584 (N_32584,N_32332,N_30676);
and U32585 (N_32585,N_31596,N_30876);
xnor U32586 (N_32586,N_32429,N_32427);
and U32587 (N_32587,N_30629,N_31688);
nand U32588 (N_32588,N_31766,N_31884);
nor U32589 (N_32589,N_31092,N_32285);
nand U32590 (N_32590,N_30826,N_32248);
nand U32591 (N_32591,N_30423,N_31996);
nor U32592 (N_32592,N_30174,N_31821);
xnor U32593 (N_32593,N_31251,N_32064);
nand U32594 (N_32594,N_30235,N_31812);
nand U32595 (N_32595,N_31589,N_30401);
nor U32596 (N_32596,N_32466,N_31895);
and U32597 (N_32597,N_30464,N_31704);
nand U32598 (N_32598,N_30936,N_30746);
or U32599 (N_32599,N_30420,N_30012);
nand U32600 (N_32600,N_31425,N_30903);
nor U32601 (N_32601,N_31932,N_31080);
or U32602 (N_32602,N_30136,N_32020);
nor U32603 (N_32603,N_30042,N_30904);
nor U32604 (N_32604,N_30881,N_31018);
xor U32605 (N_32605,N_31608,N_31544);
xor U32606 (N_32606,N_31685,N_31381);
and U32607 (N_32607,N_30486,N_32195);
nor U32608 (N_32608,N_32479,N_31297);
nand U32609 (N_32609,N_30929,N_32435);
xnor U32610 (N_32610,N_31122,N_32243);
xor U32611 (N_32611,N_30120,N_32372);
and U32612 (N_32612,N_30480,N_30171);
or U32613 (N_32613,N_31200,N_31530);
nor U32614 (N_32614,N_30569,N_31207);
or U32615 (N_32615,N_31732,N_31599);
nand U32616 (N_32616,N_30340,N_31843);
xnor U32617 (N_32617,N_31967,N_30906);
or U32618 (N_32618,N_31517,N_31745);
nand U32619 (N_32619,N_31477,N_31327);
nand U32620 (N_32620,N_30245,N_30289);
xnor U32621 (N_32621,N_30834,N_32349);
and U32622 (N_32622,N_30805,N_30765);
and U32623 (N_32623,N_31747,N_30915);
xnor U32624 (N_32624,N_30108,N_31412);
nor U32625 (N_32625,N_31973,N_32146);
and U32626 (N_32626,N_31602,N_31289);
nor U32627 (N_32627,N_32408,N_31815);
xnor U32628 (N_32628,N_31992,N_31146);
and U32629 (N_32629,N_30205,N_30794);
or U32630 (N_32630,N_31793,N_30555);
xor U32631 (N_32631,N_32331,N_30791);
xor U32632 (N_32632,N_30089,N_31062);
or U32633 (N_32633,N_30327,N_32066);
or U32634 (N_32634,N_32425,N_32144);
xor U32635 (N_32635,N_31673,N_31635);
and U32636 (N_32636,N_31795,N_31729);
nor U32637 (N_32637,N_30849,N_30750);
or U32638 (N_32638,N_30782,N_32121);
and U32639 (N_32639,N_31613,N_32324);
nor U32640 (N_32640,N_31550,N_31662);
nor U32641 (N_32641,N_30748,N_31553);
xnor U32642 (N_32642,N_31466,N_30992);
nand U32643 (N_32643,N_32196,N_31733);
xor U32644 (N_32644,N_30532,N_32090);
xor U32645 (N_32645,N_30119,N_30864);
and U32646 (N_32646,N_30813,N_31402);
or U32647 (N_32647,N_30559,N_32375);
and U32648 (N_32648,N_30662,N_31442);
nand U32649 (N_32649,N_31284,N_31831);
and U32650 (N_32650,N_31489,N_31413);
nand U32651 (N_32651,N_31842,N_31339);
or U32652 (N_32652,N_30291,N_31811);
xor U32653 (N_32653,N_32274,N_30492);
xnor U32654 (N_32654,N_30332,N_32057);
or U32655 (N_32655,N_31593,N_31880);
or U32656 (N_32656,N_31696,N_32114);
or U32657 (N_32657,N_31387,N_30969);
nor U32658 (N_32658,N_32426,N_31878);
nand U32659 (N_32659,N_32180,N_30347);
and U32660 (N_32660,N_31791,N_31790);
xor U32661 (N_32661,N_30035,N_31922);
nor U32662 (N_32662,N_30770,N_31154);
nand U32663 (N_32663,N_32380,N_30557);
nor U32664 (N_32664,N_30875,N_32316);
nor U32665 (N_32665,N_30683,N_31272);
or U32666 (N_32666,N_30563,N_31810);
xor U32667 (N_32667,N_30796,N_30998);
nor U32668 (N_32668,N_30752,N_31153);
nor U32669 (N_32669,N_30001,N_32152);
nor U32670 (N_32670,N_31214,N_31436);
or U32671 (N_32671,N_31134,N_30085);
nand U32672 (N_32672,N_31962,N_31282);
and U32673 (N_32673,N_31262,N_31483);
nand U32674 (N_32674,N_30409,N_32137);
and U32675 (N_32675,N_30682,N_30575);
or U32676 (N_32676,N_31012,N_31742);
xor U32677 (N_32677,N_32032,N_31983);
and U32678 (N_32678,N_32489,N_32107);
nand U32679 (N_32679,N_30605,N_31296);
xor U32680 (N_32680,N_32232,N_31775);
nor U32681 (N_32681,N_31249,N_31163);
xor U32682 (N_32682,N_32060,N_31763);
nor U32683 (N_32683,N_30919,N_31735);
xor U32684 (N_32684,N_30204,N_30072);
xnor U32685 (N_32685,N_30467,N_31902);
and U32686 (N_32686,N_31897,N_30278);
or U32687 (N_32687,N_31234,N_31335);
and U32688 (N_32688,N_30893,N_31051);
xor U32689 (N_32689,N_31676,N_30952);
nor U32690 (N_32690,N_32458,N_31785);
xnor U32691 (N_32691,N_30039,N_30809);
or U32692 (N_32692,N_31159,N_31659);
or U32693 (N_32693,N_31714,N_32125);
nor U32694 (N_32694,N_32183,N_31855);
and U32695 (N_32695,N_32279,N_30527);
and U32696 (N_32696,N_31020,N_30169);
nand U32697 (N_32697,N_30537,N_30167);
nor U32698 (N_32698,N_31711,N_31839);
nand U32699 (N_32699,N_31925,N_30997);
nand U32700 (N_32700,N_30804,N_31292);
xor U32701 (N_32701,N_31769,N_31247);
and U32702 (N_32702,N_31373,N_30261);
and U32703 (N_32703,N_31611,N_31514);
and U32704 (N_32704,N_30317,N_32014);
nor U32705 (N_32705,N_30276,N_31910);
or U32706 (N_32706,N_30300,N_31677);
nor U32707 (N_32707,N_31242,N_30392);
and U32708 (N_32708,N_32447,N_31231);
or U32709 (N_32709,N_32321,N_32271);
or U32710 (N_32710,N_32277,N_30456);
nor U32711 (N_32711,N_32038,N_30847);
and U32712 (N_32712,N_32494,N_31478);
nor U32713 (N_32713,N_31379,N_31304);
nand U32714 (N_32714,N_30764,N_31573);
nand U32715 (N_32715,N_30482,N_31912);
or U32716 (N_32716,N_31032,N_31107);
xor U32717 (N_32717,N_31235,N_31951);
nand U32718 (N_32718,N_30259,N_32289);
and U32719 (N_32719,N_31254,N_31885);
nor U32720 (N_32720,N_31828,N_31082);
and U32721 (N_32721,N_31090,N_32048);
and U32722 (N_32722,N_31052,N_32360);
or U32723 (N_32723,N_30144,N_30716);
or U32724 (N_32724,N_31376,N_30908);
nand U32725 (N_32725,N_30509,N_31377);
nand U32726 (N_32726,N_32188,N_31465);
nand U32727 (N_32727,N_31104,N_30610);
nor U32728 (N_32728,N_30074,N_32340);
nor U32729 (N_32729,N_32390,N_30885);
xnor U32730 (N_32730,N_30595,N_30121);
xor U32731 (N_32731,N_31130,N_32190);
xor U32732 (N_32732,N_30666,N_31137);
nor U32733 (N_32733,N_31091,N_31535);
nor U32734 (N_32734,N_31460,N_32268);
xor U32735 (N_32735,N_31194,N_32320);
nand U32736 (N_32736,N_31337,N_30548);
nor U32737 (N_32737,N_32301,N_31813);
nand U32738 (N_32738,N_31127,N_32347);
nand U32739 (N_32739,N_30271,N_31846);
xnor U32740 (N_32740,N_31870,N_32251);
or U32741 (N_32741,N_32364,N_30268);
nor U32742 (N_32742,N_32077,N_31308);
nand U32743 (N_32743,N_32002,N_30381);
nand U32744 (N_32744,N_30129,N_31888);
xor U32745 (N_32745,N_31708,N_30941);
xor U32746 (N_32746,N_31307,N_30184);
xnor U32747 (N_32747,N_30863,N_30011);
and U32748 (N_32748,N_32123,N_31700);
and U32749 (N_32749,N_31522,N_31439);
and U32750 (N_32750,N_31277,N_31407);
or U32751 (N_32751,N_31906,N_30626);
and U32752 (N_32752,N_31829,N_31666);
nor U32753 (N_32753,N_30060,N_31603);
or U32754 (N_32754,N_31770,N_31389);
xor U32755 (N_32755,N_31626,N_31359);
or U32756 (N_32756,N_31473,N_30066);
nor U32757 (N_32757,N_30339,N_31179);
xnor U32758 (N_32758,N_32192,N_30925);
or U32759 (N_32759,N_32284,N_31240);
and U32760 (N_32760,N_30195,N_31375);
or U32761 (N_32761,N_31952,N_32345);
xor U32762 (N_32762,N_31505,N_30757);
or U32763 (N_32763,N_31679,N_32276);
nor U32764 (N_32764,N_32434,N_30909);
xnor U32765 (N_32765,N_30588,N_31601);
xnor U32766 (N_32766,N_32262,N_30833);
nor U32767 (N_32767,N_31901,N_31258);
xor U32768 (N_32768,N_31246,N_31279);
xnor U32769 (N_32769,N_30170,N_31622);
or U32770 (N_32770,N_31341,N_31364);
or U32771 (N_32771,N_32056,N_30681);
and U32772 (N_32772,N_30466,N_30080);
nor U32773 (N_32773,N_31642,N_30902);
xnor U32774 (N_32774,N_30735,N_30672);
or U32775 (N_32775,N_31315,N_32379);
nand U32776 (N_32776,N_30570,N_31614);
nand U32777 (N_32777,N_31241,N_30668);
and U32778 (N_32778,N_32267,N_30556);
or U32779 (N_32779,N_30358,N_31848);
nand U32780 (N_32780,N_31920,N_31328);
nor U32781 (N_32781,N_30730,N_32476);
nor U32782 (N_32782,N_30907,N_30384);
nor U32783 (N_32783,N_30091,N_30054);
nand U32784 (N_32784,N_30698,N_32407);
or U32785 (N_32785,N_30413,N_30516);
xor U32786 (N_32786,N_30792,N_30194);
nor U32787 (N_32787,N_30468,N_32328);
or U32788 (N_32788,N_30427,N_31017);
or U32789 (N_32789,N_32406,N_31545);
nor U32790 (N_32790,N_31369,N_31470);
xor U32791 (N_32791,N_30598,N_30739);
and U32792 (N_32792,N_32351,N_31064);
nand U32793 (N_32793,N_31050,N_32414);
xor U32794 (N_32794,N_30143,N_30868);
or U32795 (N_32795,N_30479,N_30236);
and U32796 (N_32796,N_30388,N_30172);
nor U32797 (N_32797,N_31405,N_31809);
nor U32798 (N_32798,N_30521,N_31817);
nand U32799 (N_32799,N_30015,N_31693);
or U32800 (N_32800,N_31010,N_30905);
and U32801 (N_32801,N_32215,N_30154);
nor U32802 (N_32802,N_31026,N_32235);
and U32803 (N_32803,N_30711,N_31926);
or U32804 (N_32804,N_30227,N_32105);
nor U32805 (N_32805,N_30652,N_31886);
or U32806 (N_32806,N_30950,N_30700);
and U32807 (N_32807,N_32281,N_31508);
and U32808 (N_32808,N_31836,N_31993);
nand U32809 (N_32809,N_32042,N_30865);
xnor U32810 (N_32810,N_32411,N_32388);
and U32811 (N_32811,N_31587,N_30801);
or U32812 (N_32812,N_31649,N_30251);
nor U32813 (N_32813,N_30994,N_30284);
or U32814 (N_32814,N_32145,N_31228);
xnor U32815 (N_32815,N_32443,N_31930);
nand U32816 (N_32816,N_30525,N_32186);
or U32817 (N_32817,N_30670,N_30397);
and U32818 (N_32818,N_30658,N_31792);
nor U32819 (N_32819,N_32256,N_32065);
xnor U32820 (N_32820,N_31382,N_30110);
or U32821 (N_32821,N_31372,N_30298);
nor U32822 (N_32822,N_31929,N_31556);
nand U32823 (N_32823,N_32369,N_31066);
nand U32824 (N_32824,N_30872,N_31536);
and U32825 (N_32825,N_31349,N_32040);
nand U32826 (N_32826,N_31911,N_31484);
nor U32827 (N_32827,N_30285,N_31969);
or U32828 (N_32828,N_30044,N_32087);
nand U32829 (N_32829,N_31285,N_30342);
xor U32830 (N_32830,N_30891,N_31816);
and U32831 (N_32831,N_32445,N_30879);
xnor U32832 (N_32832,N_31678,N_30924);
and U32833 (N_32833,N_32177,N_32166);
nand U32834 (N_32834,N_30368,N_32109);
nand U32835 (N_32835,N_30336,N_30371);
nand U32836 (N_32836,N_30009,N_32194);
or U32837 (N_32837,N_31741,N_30295);
nor U32838 (N_32838,N_30461,N_31049);
nand U32839 (N_32839,N_31954,N_32173);
xnor U32840 (N_32840,N_31955,N_31073);
or U32841 (N_32841,N_30441,N_31264);
nand U32842 (N_32842,N_31660,N_31220);
and U32843 (N_32843,N_31958,N_30761);
nand U32844 (N_32844,N_30506,N_30628);
nand U32845 (N_32845,N_31170,N_31851);
nor U32846 (N_32846,N_30258,N_31156);
nor U32847 (N_32847,N_31058,N_31534);
xor U32848 (N_32848,N_31502,N_32478);
nor U32849 (N_32849,N_30000,N_31298);
and U32850 (N_32850,N_30633,N_30232);
xnor U32851 (N_32851,N_30584,N_31761);
and U32852 (N_32852,N_30431,N_30667);
xor U32853 (N_32853,N_32158,N_31694);
or U32854 (N_32854,N_30953,N_31751);
and U32855 (N_32855,N_30661,N_31196);
nor U32856 (N_32856,N_32330,N_32312);
nand U32857 (N_32857,N_31459,N_30592);
nand U32858 (N_32858,N_32460,N_31498);
or U32859 (N_32859,N_30148,N_30665);
xor U32860 (N_32860,N_32462,N_32050);
and U32861 (N_32861,N_30100,N_32493);
xnor U32862 (N_32862,N_30591,N_30545);
or U32863 (N_32863,N_32204,N_31086);
xnor U32864 (N_32864,N_32227,N_30541);
nand U32865 (N_32865,N_30679,N_31725);
xnor U32866 (N_32866,N_30425,N_31715);
or U32867 (N_32867,N_32034,N_30737);
and U32868 (N_32868,N_30274,N_30505);
and U32869 (N_32869,N_30751,N_30487);
and U32870 (N_32870,N_31692,N_30828);
nand U32871 (N_32871,N_31128,N_30287);
nor U32872 (N_32872,N_30237,N_30624);
or U32873 (N_32873,N_32459,N_32314);
nor U32874 (N_32874,N_31362,N_30916);
and U32875 (N_32875,N_30411,N_31706);
and U32876 (N_32876,N_32412,N_30003);
nand U32877 (N_32877,N_31336,N_31480);
xor U32878 (N_32878,N_30533,N_32205);
nand U32879 (N_32879,N_32122,N_32488);
or U32880 (N_32880,N_32381,N_30835);
nand U32881 (N_32881,N_30215,N_30853);
xnor U32882 (N_32882,N_30951,N_31273);
and U32883 (N_32883,N_30694,N_30621);
or U32884 (N_32884,N_32170,N_30883);
and U32885 (N_32885,N_31744,N_31044);
and U32886 (N_32886,N_30355,N_31318);
xnor U32887 (N_32887,N_30117,N_30597);
and U32888 (N_32888,N_31585,N_31210);
nand U32889 (N_32889,N_30522,N_32242);
or U32890 (N_32890,N_31406,N_31762);
and U32891 (N_32891,N_30646,N_30252);
xor U32892 (N_32892,N_31604,N_31532);
xnor U32893 (N_32893,N_31310,N_31914);
nand U32894 (N_32894,N_30819,N_31617);
and U32895 (N_32895,N_30957,N_30326);
or U32896 (N_32896,N_31350,N_31640);
and U32897 (N_32897,N_32457,N_30097);
xor U32898 (N_32898,N_30377,N_32236);
or U32899 (N_32899,N_30412,N_30890);
nand U32900 (N_32900,N_30489,N_31616);
xnor U32901 (N_32901,N_31174,N_30292);
nand U32902 (N_32902,N_31096,N_30226);
and U32903 (N_32903,N_32322,N_31002);
xnor U32904 (N_32904,N_31689,N_32451);
nor U32905 (N_32905,N_31834,N_30973);
nand U32906 (N_32906,N_30281,N_31825);
nor U32907 (N_32907,N_30535,N_30216);
nor U32908 (N_32908,N_32337,N_30088);
nand U32909 (N_32909,N_32103,N_30926);
xor U32910 (N_32910,N_32278,N_31147);
nor U32911 (N_32911,N_30168,N_30510);
nand U32912 (N_32912,N_31495,N_31024);
or U32913 (N_32913,N_32413,N_30701);
and U32914 (N_32914,N_31995,N_32149);
nor U32915 (N_32915,N_31520,N_30762);
and U32916 (N_32916,N_31663,N_30434);
nand U32917 (N_32917,N_31084,N_32181);
and U32918 (N_32918,N_32023,N_31994);
or U32919 (N_32919,N_30897,N_32115);
xor U32920 (N_32920,N_30808,N_30083);
nor U32921 (N_32921,N_32348,N_31429);
or U32922 (N_32922,N_30240,N_32059);
or U32923 (N_32923,N_31109,N_32461);
xor U32924 (N_32924,N_30391,N_32467);
and U32925 (N_32925,N_30132,N_30210);
xor U32926 (N_32926,N_31612,N_31841);
and U32927 (N_32927,N_31760,N_30959);
or U32928 (N_32928,N_32172,N_31055);
and U32929 (N_32929,N_30852,N_30632);
nor U32930 (N_32930,N_30607,N_32303);
nor U32931 (N_32931,N_30433,N_31449);
nand U32932 (N_32932,N_30945,N_30577);
xnor U32933 (N_32933,N_32044,N_30145);
nor U32934 (N_32934,N_31664,N_30027);
nor U32935 (N_32935,N_31386,N_32350);
xor U32936 (N_32936,N_30002,N_30830);
nand U32937 (N_32937,N_32085,N_31868);
xor U32938 (N_32938,N_30558,N_31176);
nand U32939 (N_32939,N_32288,N_30488);
or U32940 (N_32940,N_30138,N_31312);
and U32941 (N_32941,N_31837,N_32399);
nand U32942 (N_32942,N_31583,N_32161);
xnor U32943 (N_32943,N_30709,N_31794);
nand U32944 (N_32944,N_32046,N_32419);
nand U32945 (N_32945,N_30810,N_31069);
and U32946 (N_32946,N_31396,N_31991);
or U32947 (N_32947,N_30723,N_32420);
nor U32948 (N_32948,N_30019,N_30798);
nand U32949 (N_32949,N_32253,N_31039);
and U32950 (N_32950,N_30648,N_30114);
and U32951 (N_32951,N_30986,N_30328);
nor U32952 (N_32952,N_32202,N_30301);
and U32953 (N_32953,N_31503,N_31866);
nand U32954 (N_32954,N_31288,N_31059);
xnor U32955 (N_32955,N_32179,N_31366);
xor U32956 (N_32956,N_31988,N_30014);
and U32957 (N_32957,N_31555,N_30552);
or U32958 (N_32958,N_31516,N_30504);
and U32959 (N_32959,N_30651,N_31531);
or U32960 (N_32960,N_32428,N_30566);
nand U32961 (N_32961,N_30346,N_31203);
nand U32962 (N_32962,N_32045,N_32036);
or U32963 (N_32963,N_31686,N_30203);
xor U32964 (N_32964,N_31270,N_30498);
nor U32965 (N_32965,N_30910,N_30724);
and U32966 (N_32966,N_30056,N_31680);
and U32967 (N_32967,N_31000,N_30574);
xor U32968 (N_32968,N_30061,N_30637);
and U32969 (N_32969,N_30878,N_31571);
or U32970 (N_32970,N_31110,N_32482);
nand U32971 (N_32971,N_31518,N_30721);
nor U32972 (N_32972,N_31226,N_30614);
xnor U32973 (N_32973,N_31456,N_30269);
and U32974 (N_32974,N_30107,N_31605);
and U32975 (N_32975,N_30547,N_30321);
and U32976 (N_32976,N_31195,N_30393);
xnor U32977 (N_32977,N_30838,N_31063);
or U32978 (N_32978,N_30696,N_32402);
and U32979 (N_32979,N_30688,N_31079);
nand U32980 (N_32980,N_30571,N_32218);
nor U32981 (N_32981,N_31504,N_32148);
nand U32982 (N_32982,N_31441,N_32336);
nor U32983 (N_32983,N_32027,N_31115);
or U32984 (N_32984,N_32257,N_30273);
xor U32985 (N_32985,N_31048,N_31303);
nand U32986 (N_32986,N_30198,N_30578);
or U32987 (N_32987,N_31942,N_32386);
nor U32988 (N_32988,N_30857,N_32473);
nand U32989 (N_32989,N_31144,N_31269);
nor U32990 (N_32990,N_30713,N_32401);
nor U32991 (N_32991,N_31351,N_32171);
or U32992 (N_32992,N_31568,N_30247);
and U32993 (N_32993,N_30918,N_31674);
and U32994 (N_32994,N_31779,N_31557);
or U32995 (N_32995,N_32199,N_30601);
or U32996 (N_32996,N_30113,N_31947);
nand U32997 (N_32997,N_30234,N_31083);
xnor U32998 (N_32998,N_31691,N_30766);
and U32999 (N_32999,N_30534,N_31636);
and U33000 (N_33000,N_30279,N_31899);
xor U33001 (N_33001,N_31365,N_31987);
nor U33002 (N_33002,N_30786,N_32224);
xnor U33003 (N_33003,N_31900,N_32287);
and U33004 (N_33004,N_32082,N_31784);
nand U33005 (N_33005,N_30821,N_30740);
or U33006 (N_33006,N_30360,N_32047);
nand U33007 (N_33007,N_32230,N_30586);
nand U33008 (N_33008,N_31184,N_31801);
nor U33009 (N_33009,N_31776,N_30150);
nand U33010 (N_33010,N_32200,N_31871);
xor U33011 (N_33011,N_30407,N_30977);
nor U33012 (N_33012,N_31782,N_31509);
xor U33013 (N_33013,N_30882,N_32396);
xnor U33014 (N_33014,N_32254,N_30109);
and U33015 (N_33015,N_31126,N_30710);
xor U33016 (N_33016,N_32151,N_31510);
nand U33017 (N_33017,N_31324,N_30090);
nand U33018 (N_33018,N_31116,N_31071);
xnor U33019 (N_33019,N_32081,N_31548);
or U33020 (N_33020,N_30350,N_31102);
nor U33021 (N_33021,N_30841,N_32100);
nor U33022 (N_33022,N_32415,N_31739);
nor U33023 (N_33023,N_31961,N_30288);
nor U33024 (N_33024,N_32093,N_31421);
nor U33025 (N_33025,N_31263,N_31078);
or U33026 (N_33026,N_31348,N_32086);
or U33027 (N_33027,N_32405,N_32339);
nand U33028 (N_33028,N_31035,N_30642);
or U33029 (N_33029,N_30779,N_30224);
and U33030 (N_33030,N_31832,N_30299);
or U33031 (N_33031,N_30069,N_32263);
or U33032 (N_33032,N_31697,N_30081);
nor U33033 (N_33033,N_32213,N_30084);
nor U33034 (N_33034,N_31178,N_31056);
or U33035 (N_33035,N_31094,N_31717);
xnor U33036 (N_33036,N_30697,N_30775);
xor U33037 (N_33037,N_32176,N_31447);
or U33038 (N_33038,N_30600,N_30310);
or U33039 (N_33039,N_32153,N_32247);
nor U33040 (N_33040,N_31780,N_30946);
and U33041 (N_33041,N_32361,N_32298);
xor U33042 (N_33042,N_30106,N_30337);
xor U33043 (N_33043,N_30387,N_30073);
nor U33044 (N_33044,N_31274,N_31112);
or U33045 (N_33045,N_32245,N_30348);
nand U33046 (N_33046,N_32132,N_30142);
or U33047 (N_33047,N_30485,N_30102);
nor U33048 (N_33048,N_32133,N_30410);
nand U33049 (N_33049,N_30783,N_31431);
nand U33050 (N_33050,N_31600,N_30331);
nor U33051 (N_33051,N_30917,N_30243);
nor U33052 (N_33052,N_31033,N_30565);
nor U33053 (N_33053,N_31892,N_30118);
nand U33054 (N_33054,N_31397,N_31476);
or U33055 (N_33055,N_30325,N_32201);
nor U33056 (N_33056,N_31638,N_30476);
nor U33057 (N_33057,N_31591,N_31171);
nor U33058 (N_33058,N_30450,N_30777);
nand U33059 (N_33059,N_30526,N_31850);
and U33060 (N_33060,N_31070,N_30983);
and U33061 (N_33061,N_31021,N_31399);
nor U33062 (N_33062,N_32317,N_31388);
nor U33063 (N_33063,N_30322,N_32442);
nand U33064 (N_33064,N_30311,N_30082);
nand U33065 (N_33065,N_31003,N_30160);
or U33066 (N_33066,N_31016,N_31551);
or U33067 (N_33067,N_32211,N_30589);
nor U33068 (N_33068,N_30923,N_32323);
nand U33069 (N_33069,N_30519,N_30616);
or U33070 (N_33070,N_31874,N_30884);
xor U33071 (N_33071,N_30754,N_31097);
nand U33072 (N_33072,N_31189,N_30277);
nor U33073 (N_33073,N_30333,N_30436);
or U33074 (N_33074,N_32117,N_30631);
or U33075 (N_33075,N_30189,N_30640);
nand U33076 (N_33076,N_32159,N_32450);
and U33077 (N_33077,N_31136,N_30617);
nand U33078 (N_33078,N_31481,N_32174);
xor U33079 (N_33079,N_31287,N_30999);
or U33080 (N_33080,N_32241,N_30312);
and U33081 (N_33081,N_31661,N_32229);
or U33082 (N_33082,N_30962,N_32355);
nor U33083 (N_33083,N_31634,N_31748);
or U33084 (N_33084,N_31103,N_32250);
or U33085 (N_33085,N_30124,N_30837);
or U33086 (N_33086,N_30454,N_30262);
and U33087 (N_33087,N_32189,N_32167);
nand U33088 (N_33088,N_30500,N_32147);
xor U33089 (N_33089,N_30901,N_32359);
and U33090 (N_33090,N_31230,N_32410);
and U33091 (N_33091,N_32225,N_30528);
or U33092 (N_33092,N_30725,N_30706);
or U33093 (N_33093,N_31863,N_32073);
nand U33094 (N_33094,N_32432,N_32469);
or U33095 (N_33095,N_31669,N_32378);
and U33096 (N_33096,N_31750,N_31423);
and U33097 (N_33097,N_32308,N_30302);
or U33098 (N_33098,N_31627,N_31781);
or U33099 (N_33099,N_32244,N_30316);
and U33100 (N_33100,N_32290,N_30459);
or U33101 (N_33101,N_31325,N_30372);
and U33102 (N_33102,N_32005,N_31019);
or U33103 (N_33103,N_32465,N_31597);
nand U33104 (N_33104,N_32313,N_31702);
or U33105 (N_33105,N_31047,N_31099);
or U33106 (N_33106,N_31212,N_30942);
or U33107 (N_33107,N_31528,N_30760);
or U33108 (N_33108,N_30715,N_30913);
xnor U33109 (N_33109,N_30769,N_30439);
nand U33110 (N_33110,N_30116,N_32017);
nand U33111 (N_33111,N_30474,N_30253);
xnor U33112 (N_33112,N_30099,N_30712);
nand U33113 (N_33113,N_31970,N_30442);
xnor U33114 (N_33114,N_31067,N_31463);
xor U33115 (N_33115,N_30432,N_31493);
nand U33116 (N_33116,N_30717,N_30030);
and U33117 (N_33117,N_30844,N_32140);
xor U33118 (N_33118,N_32452,N_30265);
xnor U33119 (N_33119,N_30395,N_30111);
and U33120 (N_33120,N_32395,N_32175);
and U33121 (N_33121,N_30306,N_30996);
or U33122 (N_33122,N_30703,N_31280);
nand U33123 (N_33123,N_31645,N_30836);
nand U33124 (N_33124,N_32041,N_30859);
or U33125 (N_33125,N_32184,N_30795);
xnor U33126 (N_33126,N_30553,N_30967);
nor U33127 (N_33127,N_31523,N_30460);
xnor U33128 (N_33128,N_30514,N_31213);
xnor U33129 (N_33129,N_31789,N_30799);
xor U33130 (N_33130,N_30481,N_31654);
nor U33131 (N_33131,N_32282,N_30156);
xor U33132 (N_33132,N_30307,N_31624);
nand U33133 (N_33133,N_30031,N_30686);
xor U33134 (N_33134,N_31707,N_32238);
nor U33135 (N_33135,N_30212,N_30745);
nand U33136 (N_33136,N_30660,N_30877);
xnor U33137 (N_33137,N_32422,N_31191);
and U33138 (N_33138,N_31629,N_32015);
nor U33139 (N_33139,N_32226,N_30975);
and U33140 (N_33140,N_31005,N_32185);
and U33141 (N_33141,N_31417,N_30286);
nand U33142 (N_33142,N_30771,N_30353);
nor U33143 (N_33143,N_31131,N_32304);
xnor U33144 (N_33144,N_31898,N_31344);
nand U33145 (N_33145,N_30440,N_31931);
nand U33146 (N_33146,N_32061,N_32119);
nand U33147 (N_33147,N_31824,N_30550);
nand U33148 (N_33148,N_32214,N_32371);
and U33149 (N_33149,N_30177,N_31598);
nor U33150 (N_33150,N_30889,N_31783);
nor U33151 (N_33151,N_31237,N_30583);
or U33152 (N_33152,N_32134,N_30033);
and U33153 (N_33153,N_30164,N_32273);
or U33154 (N_33154,N_30699,N_31823);
xor U33155 (N_33155,N_30990,N_31471);
and U33156 (N_33156,N_31552,N_31561);
nor U33157 (N_33157,N_30445,N_32449);
or U33158 (N_33158,N_30021,N_31857);
xnor U33159 (N_33159,N_30161,N_31265);
nand U33160 (N_33160,N_31180,N_30173);
nand U33161 (N_33161,N_30733,N_30140);
xor U33162 (N_33162,N_32283,N_30627);
or U33163 (N_33163,N_30155,N_30518);
nor U33164 (N_33164,N_30933,N_32129);
nand U33165 (N_33165,N_31488,N_31354);
or U33166 (N_33166,N_30680,N_32391);
or U33167 (N_33167,N_30815,N_30728);
and U33168 (N_33168,N_30267,N_31726);
xor U33169 (N_33169,N_30448,N_30484);
nor U33170 (N_33170,N_31574,N_31268);
xnor U33171 (N_33171,N_31455,N_30345);
or U33172 (N_33172,N_30246,N_30380);
or U33173 (N_33173,N_31957,N_32310);
nor U33174 (N_33174,N_30669,N_32338);
xor U33175 (N_33175,N_31081,N_30222);
nor U33176 (N_33176,N_30495,N_31965);
or U33177 (N_33177,N_30206,N_32068);
nand U33178 (N_33178,N_32097,N_31038);
xor U33179 (N_33179,N_30980,N_31068);
nor U33180 (N_33180,N_31383,N_30596);
nor U33181 (N_33181,N_31320,N_31401);
nor U33182 (N_33182,N_30949,N_30365);
xnor U33183 (N_33183,N_31361,N_30323);
or U33184 (N_33184,N_30283,N_32024);
nand U33185 (N_33185,N_30366,N_31135);
and U33186 (N_33186,N_30812,N_30593);
nor U33187 (N_33187,N_31858,N_32004);
xnor U33188 (N_33188,N_30705,N_30398);
xnor U33189 (N_33189,N_30147,N_31797);
xor U33190 (N_33190,N_30987,N_30225);
nand U33191 (N_33191,N_32028,N_32212);
nand U33192 (N_33192,N_32168,N_31853);
nand U33193 (N_33193,N_31515,N_30408);
or U33194 (N_33194,N_32069,N_31248);
or U33195 (N_33195,N_30126,N_31202);
nand U33196 (N_33196,N_30029,N_31916);
or U33197 (N_33197,N_30972,N_30984);
and U33198 (N_33198,N_30993,N_30604);
and U33199 (N_33199,N_31822,N_31773);
nand U33200 (N_33200,N_30068,N_32062);
nor U33201 (N_33201,N_31655,N_31295);
xor U33202 (N_33202,N_31166,N_30004);
or U33203 (N_33203,N_31291,N_30221);
nand U33204 (N_33204,N_30790,N_32088);
nor U33205 (N_33205,N_30463,N_31187);
or U33206 (N_33206,N_30280,N_30970);
nand U33207 (N_33207,N_31519,N_31290);
nand U33208 (N_33208,N_31225,N_30931);
nand U33209 (N_33209,N_30708,N_32437);
xor U33210 (N_33210,N_31087,N_30856);
or U33211 (N_33211,N_31343,N_30361);
nand U33212 (N_33212,N_30512,N_32111);
nand U33213 (N_33213,N_31474,N_30862);
nand U33214 (N_33214,N_30655,N_31521);
and U33215 (N_33215,N_30820,N_31615);
and U33216 (N_33216,N_31798,N_30026);
and U33217 (N_33217,N_32280,N_31197);
nor U33218 (N_33218,N_31525,N_30146);
or U33219 (N_33219,N_30536,N_31963);
xnor U33220 (N_33220,N_32156,N_32418);
xor U33221 (N_33221,N_30985,N_30747);
nor U33222 (N_33222,N_30207,N_30974);
nand U33223 (N_33223,N_32163,N_30417);
nor U33224 (N_33224,N_30421,N_31964);
xor U33225 (N_33225,N_30718,N_31844);
and U33226 (N_33226,N_31833,N_31740);
nand U33227 (N_33227,N_32498,N_31979);
and U33228 (N_33228,N_32016,N_31581);
nand U33229 (N_33229,N_30763,N_31646);
nor U33230 (N_33230,N_30734,N_31319);
or U33231 (N_33231,N_31639,N_32207);
nor U33232 (N_33232,N_30966,N_31524);
and U33233 (N_33233,N_31420,N_30202);
and U33234 (N_33234,N_30546,N_30065);
nand U33235 (N_33235,N_31499,N_32261);
and U33236 (N_33236,N_31252,N_31830);
or U33237 (N_33237,N_31864,N_31294);
nor U33238 (N_33238,N_30854,N_31028);
nor U33239 (N_33239,N_31630,N_30797);
nand U33240 (N_33240,N_30619,N_31223);
or U33241 (N_33241,N_30379,N_30047);
nor U33242 (N_33242,N_30773,N_31997);
nand U33243 (N_33243,N_32157,N_30714);
or U33244 (N_33244,N_31158,N_30422);
nand U33245 (N_33245,N_30007,N_31919);
xnor U33246 (N_33246,N_31305,N_30807);
xnor U33247 (N_33247,N_30720,N_30344);
nor U33248 (N_33248,N_30303,N_32233);
xor U33249 (N_33249,N_31856,N_32455);
nand U33250 (N_33250,N_31211,N_32219);
xor U33251 (N_33251,N_30443,N_31408);
and U33252 (N_33252,N_31786,N_30963);
and U33253 (N_33253,N_32297,N_30062);
and U33254 (N_33254,N_30811,N_30362);
nor U33255 (N_33255,N_31542,N_30645);
and U33256 (N_33256,N_32150,N_31378);
nand U33257 (N_33257,N_30656,N_30335);
or U33258 (N_33258,N_31314,N_30861);
nand U33259 (N_33259,N_32165,N_32485);
nand U33260 (N_33260,N_30620,N_30028);
or U33261 (N_33261,N_31358,N_32356);
nand U33262 (N_33262,N_30530,N_30806);
and U33263 (N_33263,N_31934,N_31360);
and U33264 (N_33264,N_31558,N_32477);
or U33265 (N_33265,N_30250,N_31577);
nand U33266 (N_33266,N_30390,N_32089);
xnor U33267 (N_33267,N_31398,N_31778);
xor U33268 (N_33268,N_31168,N_32300);
or U33269 (N_33269,N_31721,N_30191);
xnor U33270 (N_33270,N_31966,N_31299);
or U33271 (N_33271,N_31915,N_32051);
nor U33272 (N_33272,N_31415,N_32393);
or U33273 (N_33273,N_31445,N_30024);
nand U33274 (N_33274,N_31418,N_30991);
nor U33275 (N_33275,N_31309,N_30248);
xnor U33276 (N_33276,N_30612,N_31788);
and U33277 (N_33277,N_30451,N_31113);
nor U33278 (N_33278,N_32208,N_31283);
nand U33279 (N_33279,N_32258,N_31404);
xor U33280 (N_33280,N_30183,N_32334);
or U33281 (N_33281,N_32341,N_30824);
xor U33282 (N_33282,N_32108,N_30803);
xnor U33283 (N_33283,N_31564,N_30209);
nor U33284 (N_33284,N_31076,N_30939);
nand U33285 (N_33285,N_30149,N_30501);
nand U33286 (N_33286,N_30922,N_32448);
nor U33287 (N_33287,N_30964,N_31588);
or U33288 (N_33288,N_30756,N_31437);
and U33289 (N_33289,N_32011,N_30075);
or U33290 (N_33290,N_31152,N_31125);
and U33291 (N_33291,N_31347,N_30742);
xor U33292 (N_33292,N_30162,N_30971);
nand U33293 (N_33293,N_32423,N_30241);
or U33294 (N_33294,N_30130,N_30446);
xor U33295 (N_33295,N_32124,N_31435);
and U33296 (N_33296,N_30873,N_31746);
nand U33297 (N_33297,N_31894,N_31628);
xor U33298 (N_33298,N_32127,N_30503);
xnor U33299 (N_33299,N_31904,N_31363);
nor U33300 (N_33300,N_30139,N_30477);
and U33301 (N_33301,N_31037,N_31909);
and U33302 (N_33302,N_30473,N_32421);
and U33303 (N_33303,N_31749,N_31949);
and U33304 (N_33304,N_30095,N_31040);
or U33305 (N_33305,N_30270,N_31204);
xor U33306 (N_33306,N_30157,N_30018);
xor U33307 (N_33307,N_31710,N_31650);
xnor U33308 (N_33308,N_31185,N_30213);
nand U33309 (N_33309,N_32220,N_30472);
nand U33310 (N_33310,N_32385,N_30013);
or U33311 (N_33311,N_31777,N_32468);
or U33312 (N_33312,N_32164,N_30784);
and U33313 (N_33313,N_32487,N_32010);
xor U33314 (N_33314,N_30105,N_30214);
or U33315 (N_33315,N_31990,N_31913);
and U33316 (N_33316,N_31501,N_30726);
nand U33317 (N_33317,N_31448,N_31767);
nor U33318 (N_33318,N_30549,N_31606);
nor U33319 (N_33319,N_31245,N_30077);
xnor U33320 (N_33320,N_31940,N_32084);
or U33321 (N_33321,N_30389,N_31999);
nand U33322 (N_33322,N_30920,N_31034);
nor U33323 (N_33323,N_32029,N_31566);
and U33324 (N_33324,N_30785,N_30674);
or U33325 (N_33325,N_30772,N_30334);
xnor U33326 (N_33326,N_32352,N_30707);
nand U33327 (N_33327,N_30649,N_31346);
or U33328 (N_33328,N_31095,N_30671);
and U33329 (N_33329,N_30894,N_31117);
xnor U33330 (N_33330,N_31835,N_30606);
nor U33331 (N_33331,N_30094,N_32237);
xnor U33332 (N_33332,N_32362,N_32495);
and U33333 (N_33333,N_31006,N_31989);
or U33334 (N_33334,N_31215,N_30064);
and U33335 (N_33335,N_30137,N_31025);
and U33336 (N_33336,N_31267,N_30582);
xor U33337 (N_33337,N_32333,N_32198);
xor U33338 (N_33338,N_30639,N_32039);
nor U33339 (N_33339,N_31984,N_31787);
xnor U33340 (N_33340,N_31609,N_31675);
or U33341 (N_33341,N_30458,N_30217);
or U33342 (N_33342,N_30618,N_32116);
nand U33343 (N_33343,N_32354,N_30127);
and U33344 (N_33344,N_31921,N_32217);
or U33345 (N_33345,N_32102,N_32000);
xnor U33346 (N_33346,N_30050,N_30122);
nor U33347 (N_33347,N_31657,N_31867);
xnor U33348 (N_33348,N_31161,N_31392);
xor U33349 (N_33349,N_30038,N_30851);
or U33350 (N_33350,N_31699,N_30367);
nand U33351 (N_33351,N_30356,N_32439);
or U33352 (N_33352,N_30166,N_32306);
nand U33353 (N_33353,N_32475,N_30948);
xnor U33354 (N_33354,N_32329,N_31527);
nor U33355 (N_33355,N_30744,N_31500);
or U33356 (N_33356,N_30128,N_30469);
xor U33357 (N_33357,N_31590,N_30471);
nor U33358 (N_33358,N_32118,N_32021);
nand U33359 (N_33359,N_30995,N_31800);
xnor U33360 (N_33360,N_30230,N_30415);
nand U33361 (N_33361,N_31756,N_32131);
nor U33362 (N_33362,N_32033,N_30978);
nand U33363 (N_33363,N_31854,N_31009);
or U33364 (N_33364,N_31633,N_31022);
nor U33365 (N_33365,N_30135,N_31719);
and U33366 (N_33366,N_30641,N_30899);
nand U33367 (N_33367,N_30673,N_30057);
xor U33368 (N_33368,N_32318,N_31511);
xnor U33369 (N_33369,N_32299,N_30866);
nor U33370 (N_33370,N_32266,N_30223);
nand U33371 (N_33371,N_31001,N_31492);
nor U33372 (N_33372,N_30218,N_31494);
and U33373 (N_33373,N_32070,N_31944);
or U33374 (N_33374,N_30036,N_32293);
nor U33375 (N_33375,N_32389,N_32249);
and U33376 (N_33376,N_30653,N_30329);
and U33377 (N_33377,N_30827,N_31468);
xnor U33378 (N_33378,N_31887,N_31316);
or U33379 (N_33379,N_31043,N_31960);
xnor U33380 (N_33380,N_31238,N_32003);
or U33381 (N_33381,N_31946,N_30045);
or U33382 (N_33382,N_30517,N_32387);
nor U33383 (N_33383,N_30529,N_30523);
nor U33384 (N_33384,N_32191,N_32154);
xor U33385 (N_33385,N_31301,N_31948);
or U33386 (N_33386,N_30749,N_32483);
or U33387 (N_33387,N_30802,N_30846);
nor U33388 (N_33388,N_31579,N_32007);
and U33389 (N_33389,N_31621,N_30585);
xor U33390 (N_33390,N_30290,N_30732);
and U33391 (N_33391,N_32344,N_31956);
nor U33392 (N_33392,N_30182,N_31479);
and U33393 (N_33393,N_31623,N_31173);
nand U33394 (N_33394,N_30354,N_31271);
nand U33395 (N_33395,N_31329,N_32315);
nand U33396 (N_33396,N_31206,N_30622);
and U33397 (N_33397,N_31567,N_31497);
nand U33398 (N_33398,N_32481,N_31570);
nand U33399 (N_33399,N_30731,N_32187);
nand U33400 (N_33400,N_30141,N_31976);
and U33401 (N_33401,N_30437,N_31458);
and U33402 (N_33402,N_30041,N_32143);
nor U33403 (N_33403,N_30787,N_31029);
nand U33404 (N_33404,N_31667,N_31065);
and U33405 (N_33405,N_31757,N_31670);
nand U33406 (N_33406,N_31507,N_30496);
or U33407 (N_33407,N_30778,N_32228);
nor U33408 (N_33408,N_32383,N_30965);
and U33409 (N_33409,N_32067,N_31198);
xor U33410 (N_33410,N_30702,N_31653);
or U33411 (N_33411,N_30179,N_30774);
nor U33412 (N_33412,N_31190,N_30848);
nor U33413 (N_33413,N_30093,N_32096);
or U33414 (N_33414,N_30197,N_32013);
nor U33415 (N_33415,N_31937,N_30249);
xnor U33416 (N_33416,N_30822,N_31924);
or U33417 (N_33417,N_31443,N_32001);
or U33418 (N_33418,N_31371,N_31181);
nand U33419 (N_33419,N_30070,N_30055);
xnor U33420 (N_33420,N_31013,N_31731);
nand U33421 (N_33421,N_30609,N_30483);
nand U33422 (N_33422,N_32197,N_30211);
nand U33423 (N_33423,N_30176,N_30816);
xor U33424 (N_33424,N_30508,N_32006);
xor U33425 (N_33425,N_32074,N_31072);
and U33426 (N_33426,N_30693,N_30238);
or U33427 (N_33427,N_31860,N_30190);
xnor U33428 (N_33428,N_32365,N_31827);
xor U33429 (N_33429,N_32130,N_32309);
or U33430 (N_33430,N_31120,N_31427);
or U33431 (N_33431,N_31046,N_32259);
and U33432 (N_33432,N_31529,N_30374);
and U33433 (N_33433,N_30098,N_32377);
nor U33434 (N_33434,N_31982,N_30005);
xnor U33435 (N_33435,N_31089,N_30562);
nor U33436 (N_33436,N_31709,N_31101);
nand U33437 (N_33437,N_31008,N_31698);
nand U33438 (N_33438,N_31701,N_30308);
nor U33439 (N_33439,N_31876,N_31619);
nand U33440 (N_33440,N_30435,N_30493);
nand U33441 (N_33441,N_31730,N_30743);
or U33442 (N_33442,N_30741,N_30554);
xor U33443 (N_33443,N_30178,N_31410);
nand U33444 (N_33444,N_30032,N_30507);
nand U33445 (N_33445,N_32441,N_31053);
and U33446 (N_33446,N_31594,N_30800);
and U33447 (N_33447,N_31118,N_31133);
and U33448 (N_33448,N_30375,N_30611);
nor U33449 (N_33449,N_31208,N_30947);
nand U33450 (N_33450,N_30753,N_30023);
nand U33451 (N_33451,N_30403,N_31236);
or U33452 (N_33452,N_30043,N_30040);
nand U33453 (N_33453,N_31918,N_30960);
and U33454 (N_33454,N_32292,N_31023);
or U33455 (N_33455,N_31331,N_31943);
xor U33456 (N_33456,N_32384,N_31826);
nand U33457 (N_33457,N_31903,N_32240);
or U33458 (N_33458,N_31393,N_31737);
xor U33459 (N_33459,N_31385,N_31774);
xnor U33460 (N_33460,N_30625,N_30187);
nand U33461 (N_33461,N_31972,N_30180);
or U33462 (N_33462,N_31985,N_32374);
nand U33463 (N_33463,N_30755,N_31419);
nand U33464 (N_33464,N_30675,N_31641);
nand U33465 (N_33465,N_31266,N_31036);
nand U33466 (N_33466,N_30938,N_31703);
xor U33467 (N_33467,N_30687,N_31438);
nor U33468 (N_33468,N_32357,N_30349);
xor U33469 (N_33469,N_30025,N_31151);
and U33470 (N_33470,N_31260,N_31526);
xor U33471 (N_33471,N_32417,N_31620);
and U33472 (N_33472,N_30490,N_31060);
xnor U33473 (N_33473,N_31432,N_31980);
nand U33474 (N_33474,N_31818,N_31865);
xor U33475 (N_33475,N_30874,N_30793);
nor U33476 (N_33476,N_31847,N_31004);
nor U33477 (N_33477,N_30587,N_31467);
and U33478 (N_33478,N_31807,N_31736);
nand U33479 (N_33479,N_32264,N_31849);
xnor U33480 (N_33480,N_31695,N_31905);
nand U33481 (N_33481,N_31014,N_30053);
or U33482 (N_33482,N_30465,N_30602);
or U33483 (N_33483,N_32026,N_30016);
nand U33484 (N_33484,N_31352,N_31042);
xnor U33485 (N_33485,N_30318,N_30158);
or U33486 (N_33486,N_31644,N_31123);
and U33487 (N_33487,N_30351,N_32373);
nand U33488 (N_33488,N_31490,N_31945);
or U33489 (N_33489,N_31233,N_31119);
or U33490 (N_33490,N_30079,N_30357);
nor U33491 (N_33491,N_31205,N_30399);
xnor U33492 (N_33492,N_30341,N_31132);
and U33493 (N_33493,N_30231,N_32370);
or U33494 (N_33494,N_31950,N_30402);
and U33495 (N_33495,N_31175,N_30564);
and U33496 (N_33496,N_32054,N_30497);
and U33497 (N_33497,N_30636,N_30438);
nand U33498 (N_33498,N_30305,N_30561);
nor U33499 (N_33499,N_31537,N_31330);
nor U33500 (N_33500,N_32367,N_30125);
xnor U33501 (N_33501,N_31313,N_31491);
nand U33502 (N_33502,N_32358,N_31727);
xnor U33503 (N_33503,N_30272,N_31879);
nor U33504 (N_33504,N_30515,N_30051);
nand U33505 (N_33505,N_31311,N_30867);
xnor U33506 (N_33506,N_31416,N_32446);
nand U33507 (N_33507,N_31549,N_32342);
nand U33508 (N_33508,N_32221,N_32138);
xor U33509 (N_33509,N_32141,N_31239);
nand U33510 (N_33510,N_31138,N_30543);
and U33511 (N_33511,N_31333,N_30233);
and U33512 (N_33512,N_32099,N_30059);
nor U33513 (N_33513,N_31840,N_30982);
xor U33514 (N_33514,N_30932,N_30219);
nor U33515 (N_33515,N_31869,N_32075);
xor U33516 (N_33516,N_31370,N_31890);
and U33517 (N_33517,N_32499,N_30719);
or U33518 (N_33518,N_32222,N_30058);
or U33519 (N_33519,N_30201,N_30898);
nor U33520 (N_33520,N_30131,N_31889);
nand U33521 (N_33521,N_30338,N_30229);
nor U33522 (N_33522,N_32260,N_31648);
and U33523 (N_33523,N_30275,N_31941);
and U33524 (N_33524,N_30400,N_31077);
nor U33525 (N_33525,N_30386,N_31845);
xnor U33526 (N_33526,N_31908,N_30165);
or U33527 (N_33527,N_31164,N_32037);
nor U33528 (N_33528,N_31340,N_30163);
xnor U33529 (N_33529,N_30691,N_30940);
and U33530 (N_33530,N_30818,N_30544);
xnor U33531 (N_33531,N_30263,N_31753);
and U33532 (N_33532,N_31229,N_31572);
xnor U33533 (N_33533,N_31883,N_32416);
nand U33534 (N_33534,N_32376,N_32239);
nor U33535 (N_33535,N_31332,N_31222);
nand U33536 (N_33536,N_30689,N_31582);
nand U33537 (N_33537,N_31444,N_31936);
or U33538 (N_33538,N_30185,N_32072);
xnor U33539 (N_33539,N_32325,N_31357);
nand U33540 (N_33540,N_31041,N_30052);
nor U33541 (N_33541,N_32104,N_30426);
and U33542 (N_33542,N_31129,N_32246);
xnor U33543 (N_33543,N_32286,N_32343);
nor U33544 (N_33544,N_30017,N_32397);
nor U33545 (N_33545,N_32094,N_30199);
or U33546 (N_33546,N_30330,N_31224);
and U33547 (N_33547,N_32311,N_32252);
and U33548 (N_33548,N_30104,N_31074);
nand U33549 (N_33549,N_32294,N_30264);
and U33550 (N_33550,N_31618,N_31563);
and U33551 (N_33551,N_31453,N_31244);
nor U33552 (N_33552,N_32193,N_31935);
or U33553 (N_33553,N_31923,N_30320);
or U33554 (N_33554,N_32400,N_31512);
and U33555 (N_33555,N_31061,N_32463);
xor U33556 (N_33556,N_31971,N_31461);
nand U33557 (N_33557,N_31578,N_32035);
or U33558 (N_33558,N_31075,N_31160);
nor U33559 (N_33559,N_30175,N_31743);
nor U33560 (N_33560,N_31450,N_31953);
nor U33561 (N_33561,N_31148,N_31538);
or U33562 (N_33562,N_30315,N_30814);
xor U33563 (N_33563,N_32043,N_31554);
xnor U33564 (N_33564,N_30134,N_31565);
nand U33565 (N_33565,N_30369,N_30181);
xor U33566 (N_33566,N_30613,N_30590);
or U33567 (N_33567,N_32444,N_30650);
nor U33568 (N_33568,N_32326,N_30825);
or U33569 (N_33569,N_32346,N_32080);
nor U33570 (N_33570,N_32022,N_32110);
nand U33571 (N_33571,N_30580,N_30282);
or U33572 (N_33572,N_30831,N_31986);
xor U33573 (N_33573,N_31569,N_30664);
nor U33574 (N_33574,N_30087,N_31472);
nor U33575 (N_33575,N_31403,N_30457);
and U33576 (N_33576,N_30123,N_30567);
nor U33577 (N_33577,N_32436,N_32018);
or U33578 (N_33578,N_30638,N_30010);
xnor U33579 (N_33579,N_31891,N_31907);
and U33580 (N_33580,N_31543,N_31440);
and U33581 (N_33581,N_32335,N_30608);
and U33582 (N_33582,N_30768,N_31088);
or U33583 (N_33583,N_31658,N_31165);
xor U33584 (N_33584,N_32120,N_31802);
and U33585 (N_33585,N_31345,N_30049);
or U33586 (N_33586,N_30452,N_32071);
nand U33587 (N_33587,N_30758,N_30067);
xor U33588 (N_33588,N_32409,N_30928);
xor U33589 (N_33589,N_31539,N_30892);
xnor U33590 (N_33590,N_32178,N_32265);
and U33591 (N_33591,N_32135,N_31433);
nand U33592 (N_33592,N_30921,N_31015);
or U33593 (N_33593,N_31862,N_31232);
xnor U33594 (N_33594,N_31216,N_30255);
and U33595 (N_33595,N_31981,N_30046);
nand U33596 (N_33596,N_31217,N_32275);
nand U33597 (N_33597,N_31454,N_32454);
xor U33598 (N_33598,N_30663,N_31150);
nor U33599 (N_33599,N_30690,N_30538);
nand U33600 (N_33600,N_32296,N_31027);
nand U33601 (N_33601,N_30870,N_30643);
nand U33602 (N_33602,N_30008,N_30086);
xnor U33603 (N_33603,N_32203,N_32128);
or U33604 (N_33604,N_30956,N_32223);
and U33605 (N_33605,N_30840,N_30428);
xor U33606 (N_33606,N_31975,N_30254);
and U33607 (N_33607,N_31275,N_31451);
nand U33608 (N_33608,N_31513,N_31394);
nor U33609 (N_33609,N_30934,N_30376);
and U33610 (N_33610,N_30542,N_31391);
and U33611 (N_33611,N_31872,N_31243);
nand U33612 (N_33612,N_31100,N_31576);
and U33613 (N_33613,N_30988,N_31108);
nand U33614 (N_33614,N_31819,N_31183);
and U33615 (N_33615,N_32008,N_32430);
nand U33616 (N_33616,N_31188,N_31560);
xor U33617 (N_33617,N_31111,N_30071);
and U33618 (N_33618,N_32382,N_32126);
nand U33619 (N_33619,N_32490,N_30895);
or U33620 (N_33620,N_30684,N_30886);
nand U33621 (N_33621,N_30447,N_30491);
nand U33622 (N_33622,N_31755,N_30373);
nor U33623 (N_33623,N_31806,N_30444);
xor U33624 (N_33624,N_31682,N_30776);
nand U33625 (N_33625,N_32210,N_30133);
xnor U33626 (N_33626,N_30193,N_30159);
nor U33627 (N_33627,N_31540,N_31169);
nand U33628 (N_33628,N_30293,N_31716);
or U33629 (N_33629,N_32142,N_32291);
and U33630 (N_33630,N_32009,N_30759);
nor U33631 (N_33631,N_30453,N_30405);
or U33632 (N_33632,N_32305,N_30729);
nand U33633 (N_33633,N_32486,N_30494);
nor U33634 (N_33634,N_31651,N_30780);
nand U33635 (N_33635,N_31011,N_30242);
nor U33636 (N_33636,N_30462,N_32019);
or U33637 (N_33637,N_31422,N_31007);
and U33638 (N_33638,N_31764,N_30961);
and U33639 (N_33639,N_30022,N_30424);
or U33640 (N_33640,N_31317,N_31261);
nor U33641 (N_33641,N_30076,N_30256);
xnor U33642 (N_33642,N_30404,N_31105);
or U33643 (N_33643,N_30112,N_31143);
and U33644 (N_33644,N_31758,N_31356);
nand U33645 (N_33645,N_30020,N_31665);
nor U33646 (N_33646,N_31162,N_31192);
xor U33647 (N_33647,N_32269,N_31643);
xnor U33648 (N_33648,N_31652,N_30858);
nor U33649 (N_33649,N_31852,N_32366);
nor U33650 (N_33650,N_30603,N_30382);
nor U33651 (N_33651,N_30429,N_31647);
nor U33652 (N_33652,N_31820,N_30499);
or U33653 (N_33653,N_30659,N_30313);
nor U33654 (N_33654,N_32353,N_31475);
nor U33655 (N_33655,N_32112,N_31149);
nand U33656 (N_33656,N_30817,N_30855);
nand U33657 (N_33657,N_32394,N_31322);
nand U33658 (N_33658,N_30513,N_30220);
xnor U33659 (N_33659,N_30418,N_32295);
nor U33660 (N_33660,N_31804,N_31772);
or U33661 (N_33661,N_31030,N_31575);
or U33662 (N_33662,N_30685,N_32368);
nor U33663 (N_33663,N_30722,N_30539);
or U33664 (N_33664,N_31803,N_32484);
or U33665 (N_33665,N_30955,N_31145);
nor U33666 (N_33666,N_31428,N_32182);
xnor U33667 (N_33667,N_31580,N_30850);
and U33668 (N_33668,N_30115,N_30630);
nor U33669 (N_33669,N_31625,N_30478);
nand U33670 (N_33670,N_31281,N_30186);
nor U33671 (N_33671,N_31482,N_30842);
xor U33672 (N_33672,N_30103,N_30989);
and U33673 (N_33673,N_31121,N_31974);
or U33674 (N_33674,N_31859,N_30006);
nand U33675 (N_33675,N_30385,N_31182);
xnor U33676 (N_33676,N_32049,N_31610);
or U33677 (N_33677,N_31139,N_31276);
or U33678 (N_33678,N_31374,N_31765);
nor U33679 (N_33679,N_31367,N_32162);
nor U33680 (N_33680,N_32209,N_30551);
and U33681 (N_33681,N_32052,N_32031);
nor U33682 (N_33682,N_31452,N_31485);
or U33683 (N_33683,N_31656,N_31323);
xor U33684 (N_33684,N_30449,N_31690);
and U33685 (N_33685,N_32092,N_30927);
nand U33686 (N_33686,N_31257,N_31395);
nor U33687 (N_33687,N_30954,N_31752);
nand U33688 (N_33688,N_30829,N_31430);
nor U33689 (N_33689,N_31045,N_31607);
or U33690 (N_33690,N_30736,N_31683);
xnor U33691 (N_33691,N_30896,N_31218);
xnor U33692 (N_33692,N_32058,N_31933);
nand U33693 (N_33693,N_32404,N_31177);
xnor U33694 (N_33694,N_31253,N_31771);
or U33695 (N_33695,N_30343,N_30871);
nand U33696 (N_33696,N_30383,N_31221);
nand U33697 (N_33697,N_31368,N_31592);
xor U33698 (N_33698,N_31334,N_32470);
or U33699 (N_33699,N_31838,N_31338);
nor U33700 (N_33700,N_30394,N_30319);
or U33701 (N_33701,N_31724,N_30968);
xor U33702 (N_33702,N_31057,N_30788);
nand U33703 (N_33703,N_30657,N_30359);
nand U33704 (N_33704,N_31928,N_31759);
xor U33705 (N_33705,N_30296,N_31671);
nor U33706 (N_33706,N_31720,N_31547);
and U33707 (N_33707,N_30615,N_32471);
or U33708 (N_33708,N_31861,N_32095);
and U33709 (N_33709,N_31713,N_31167);
nor U33710 (N_33710,N_31426,N_31098);
xor U33711 (N_33711,N_30943,N_31219);
xnor U33712 (N_33712,N_32063,N_30695);
nand U33713 (N_33713,N_31487,N_30078);
nand U33714 (N_33714,N_32101,N_31917);
or U33715 (N_33715,N_31584,N_31114);
xor U33716 (N_33716,N_31938,N_32234);
nor U33717 (N_33717,N_30572,N_30635);
nand U33718 (N_33718,N_31896,N_32155);
or U33719 (N_33719,N_30200,N_32319);
or U33720 (N_33720,N_30352,N_32270);
or U33721 (N_33721,N_31881,N_31496);
nor U33722 (N_33722,N_31728,N_30430);
xor U33723 (N_33723,N_31302,N_31286);
xnor U33724 (N_33724,N_30406,N_30738);
and U33725 (N_33725,N_32025,N_31595);
nor U33726 (N_33726,N_31278,N_30914);
xnor U33727 (N_33727,N_32433,N_30324);
nand U33728 (N_33728,N_31250,N_31486);
nor U33729 (N_33729,N_32030,N_31321);
nand U33730 (N_33730,N_30944,N_32480);
or U33731 (N_33731,N_30475,N_31411);
nand U33732 (N_33732,N_31637,N_31722);
nand U33733 (N_33733,N_30396,N_31124);
nor U33734 (N_33734,N_31684,N_32106);
xnor U33735 (N_33735,N_32053,N_31172);
and U33736 (N_33736,N_31142,N_30416);
or U33737 (N_33737,N_31939,N_32497);
xnor U33738 (N_33738,N_32076,N_30294);
and U33739 (N_33739,N_32098,N_31353);
nand U33740 (N_33740,N_31738,N_30560);
nand U33741 (N_33741,N_31959,N_31093);
and U33742 (N_33742,N_31193,N_30034);
nand U33743 (N_33743,N_30704,N_30958);
and U33744 (N_33744,N_32255,N_31546);
xor U33745 (N_33745,N_30101,N_31259);
xor U33746 (N_33746,N_32302,N_31227);
nand U33747 (N_33747,N_32012,N_30153);
nor U33748 (N_33748,N_31380,N_30188);
nand U33749 (N_33749,N_31977,N_31506);
xor U33750 (N_33750,N_32148,N_30557);
nor U33751 (N_33751,N_30857,N_30955);
nand U33752 (N_33752,N_31839,N_30586);
nor U33753 (N_33753,N_30273,N_30705);
or U33754 (N_33754,N_32144,N_30170);
xor U33755 (N_33755,N_30580,N_31349);
nor U33756 (N_33756,N_31558,N_30033);
nand U33757 (N_33757,N_30828,N_31051);
xnor U33758 (N_33758,N_30188,N_30319);
or U33759 (N_33759,N_30976,N_30265);
nor U33760 (N_33760,N_31957,N_31011);
nor U33761 (N_33761,N_31199,N_32234);
and U33762 (N_33762,N_31469,N_30830);
nor U33763 (N_33763,N_30183,N_31384);
nand U33764 (N_33764,N_30735,N_32374);
and U33765 (N_33765,N_30064,N_31409);
xnor U33766 (N_33766,N_30228,N_32313);
nor U33767 (N_33767,N_31167,N_30005);
nand U33768 (N_33768,N_30631,N_30722);
nor U33769 (N_33769,N_32370,N_30160);
nand U33770 (N_33770,N_30191,N_30524);
and U33771 (N_33771,N_30091,N_31352);
nor U33772 (N_33772,N_32217,N_30132);
and U33773 (N_33773,N_30405,N_31098);
or U33774 (N_33774,N_32150,N_30066);
nand U33775 (N_33775,N_30547,N_32211);
or U33776 (N_33776,N_31317,N_31068);
nand U33777 (N_33777,N_31923,N_31698);
or U33778 (N_33778,N_32323,N_32445);
nor U33779 (N_33779,N_32263,N_31188);
xnor U33780 (N_33780,N_30999,N_30133);
xor U33781 (N_33781,N_32216,N_30544);
xor U33782 (N_33782,N_30147,N_30925);
nor U33783 (N_33783,N_30478,N_31542);
or U33784 (N_33784,N_31983,N_30907);
xnor U33785 (N_33785,N_30896,N_32281);
and U33786 (N_33786,N_30364,N_31974);
nand U33787 (N_33787,N_30495,N_30997);
nand U33788 (N_33788,N_30222,N_31219);
and U33789 (N_33789,N_32334,N_30285);
and U33790 (N_33790,N_30688,N_31033);
nor U33791 (N_33791,N_30345,N_30033);
xor U33792 (N_33792,N_31249,N_30115);
xnor U33793 (N_33793,N_32155,N_31318);
nor U33794 (N_33794,N_31203,N_31118);
nand U33795 (N_33795,N_32023,N_30945);
or U33796 (N_33796,N_31875,N_32131);
or U33797 (N_33797,N_30340,N_31633);
nand U33798 (N_33798,N_32167,N_31327);
nand U33799 (N_33799,N_30966,N_31786);
xnor U33800 (N_33800,N_31351,N_30795);
nor U33801 (N_33801,N_30432,N_30312);
nor U33802 (N_33802,N_32070,N_31245);
nor U33803 (N_33803,N_30925,N_31559);
xor U33804 (N_33804,N_31329,N_31361);
nor U33805 (N_33805,N_31645,N_31517);
nand U33806 (N_33806,N_31938,N_30153);
xnor U33807 (N_33807,N_30682,N_31841);
and U33808 (N_33808,N_31565,N_30219);
and U33809 (N_33809,N_32207,N_31629);
and U33810 (N_33810,N_31432,N_32303);
and U33811 (N_33811,N_31371,N_32066);
or U33812 (N_33812,N_32421,N_30674);
and U33813 (N_33813,N_31988,N_31954);
nor U33814 (N_33814,N_32145,N_31856);
or U33815 (N_33815,N_30398,N_31377);
or U33816 (N_33816,N_30360,N_30740);
nor U33817 (N_33817,N_32332,N_30284);
or U33818 (N_33818,N_30719,N_31326);
or U33819 (N_33819,N_31640,N_32364);
and U33820 (N_33820,N_30503,N_30267);
nand U33821 (N_33821,N_30684,N_31883);
nand U33822 (N_33822,N_30438,N_30465);
or U33823 (N_33823,N_30819,N_30584);
nor U33824 (N_33824,N_32480,N_30911);
and U33825 (N_33825,N_31908,N_31306);
nand U33826 (N_33826,N_31777,N_31086);
nor U33827 (N_33827,N_30424,N_30235);
and U33828 (N_33828,N_32477,N_31501);
nor U33829 (N_33829,N_31770,N_30151);
nand U33830 (N_33830,N_32437,N_32032);
and U33831 (N_33831,N_30506,N_31242);
and U33832 (N_33832,N_30627,N_31511);
xnor U33833 (N_33833,N_31111,N_30598);
or U33834 (N_33834,N_30077,N_31928);
and U33835 (N_33835,N_32268,N_30705);
nand U33836 (N_33836,N_32143,N_31812);
xor U33837 (N_33837,N_31824,N_31892);
nand U33838 (N_33838,N_30017,N_31385);
xor U33839 (N_33839,N_30674,N_31746);
and U33840 (N_33840,N_31136,N_30277);
nor U33841 (N_33841,N_30023,N_30241);
nor U33842 (N_33842,N_30790,N_31345);
or U33843 (N_33843,N_31787,N_30823);
nand U33844 (N_33844,N_30372,N_32096);
or U33845 (N_33845,N_31450,N_30868);
xor U33846 (N_33846,N_31477,N_31960);
nor U33847 (N_33847,N_31546,N_30243);
and U33848 (N_33848,N_31417,N_30837);
nand U33849 (N_33849,N_31570,N_31449);
nand U33850 (N_33850,N_30650,N_30747);
or U33851 (N_33851,N_30450,N_30624);
xnor U33852 (N_33852,N_30439,N_31403);
nor U33853 (N_33853,N_30039,N_31886);
nor U33854 (N_33854,N_30969,N_31265);
xnor U33855 (N_33855,N_32091,N_32169);
or U33856 (N_33856,N_30467,N_31376);
nand U33857 (N_33857,N_31251,N_31527);
or U33858 (N_33858,N_30474,N_32258);
nor U33859 (N_33859,N_31865,N_31698);
and U33860 (N_33860,N_31515,N_32396);
nand U33861 (N_33861,N_30198,N_30500);
nand U33862 (N_33862,N_30420,N_31230);
nor U33863 (N_33863,N_31822,N_32493);
nand U33864 (N_33864,N_31410,N_32253);
or U33865 (N_33865,N_31601,N_32208);
or U33866 (N_33866,N_32002,N_31126);
nand U33867 (N_33867,N_31324,N_31363);
or U33868 (N_33868,N_30025,N_30716);
nand U33869 (N_33869,N_30026,N_30225);
or U33870 (N_33870,N_30627,N_31997);
or U33871 (N_33871,N_31653,N_30096);
and U33872 (N_33872,N_32219,N_32413);
xor U33873 (N_33873,N_30769,N_31953);
and U33874 (N_33874,N_30658,N_31401);
nor U33875 (N_33875,N_30136,N_30250);
or U33876 (N_33876,N_30458,N_31973);
and U33877 (N_33877,N_31484,N_31801);
and U33878 (N_33878,N_30889,N_30846);
xnor U33879 (N_33879,N_30271,N_31596);
xnor U33880 (N_33880,N_31573,N_30393);
or U33881 (N_33881,N_30499,N_30787);
xnor U33882 (N_33882,N_32198,N_31908);
nand U33883 (N_33883,N_31560,N_32467);
xnor U33884 (N_33884,N_31896,N_32282);
or U33885 (N_33885,N_30618,N_30473);
or U33886 (N_33886,N_32414,N_30925);
xnor U33887 (N_33887,N_31561,N_30149);
xnor U33888 (N_33888,N_30494,N_32156);
xor U33889 (N_33889,N_30049,N_31259);
xor U33890 (N_33890,N_30027,N_32153);
xnor U33891 (N_33891,N_31780,N_32222);
nor U33892 (N_33892,N_31384,N_30087);
and U33893 (N_33893,N_30161,N_32160);
nand U33894 (N_33894,N_32239,N_31935);
and U33895 (N_33895,N_30126,N_30179);
xnor U33896 (N_33896,N_31513,N_30498);
and U33897 (N_33897,N_31921,N_31911);
xnor U33898 (N_33898,N_32244,N_31618);
nor U33899 (N_33899,N_31882,N_30137);
and U33900 (N_33900,N_30697,N_31530);
nand U33901 (N_33901,N_30493,N_30182);
or U33902 (N_33902,N_32312,N_31247);
nor U33903 (N_33903,N_30057,N_30035);
xnor U33904 (N_33904,N_30003,N_31762);
xnor U33905 (N_33905,N_31350,N_31263);
nand U33906 (N_33906,N_31473,N_30214);
or U33907 (N_33907,N_32329,N_31942);
xnor U33908 (N_33908,N_31320,N_30302);
or U33909 (N_33909,N_30359,N_32136);
nor U33910 (N_33910,N_32296,N_30394);
nor U33911 (N_33911,N_31617,N_32417);
or U33912 (N_33912,N_31913,N_31983);
and U33913 (N_33913,N_32495,N_32254);
or U33914 (N_33914,N_30828,N_31411);
nor U33915 (N_33915,N_30565,N_30274);
nor U33916 (N_33916,N_32030,N_32420);
or U33917 (N_33917,N_30530,N_31834);
or U33918 (N_33918,N_32107,N_31247);
xor U33919 (N_33919,N_31756,N_32125);
or U33920 (N_33920,N_30438,N_30865);
nand U33921 (N_33921,N_32331,N_30091);
nor U33922 (N_33922,N_30155,N_30658);
nor U33923 (N_33923,N_30072,N_30080);
xnor U33924 (N_33924,N_31825,N_32072);
or U33925 (N_33925,N_30245,N_31326);
nor U33926 (N_33926,N_31863,N_30411);
nand U33927 (N_33927,N_31347,N_32099);
or U33928 (N_33928,N_30893,N_30851);
and U33929 (N_33929,N_31006,N_30990);
xor U33930 (N_33930,N_32319,N_30140);
nor U33931 (N_33931,N_31214,N_32409);
or U33932 (N_33932,N_31900,N_30136);
and U33933 (N_33933,N_31605,N_31217);
nor U33934 (N_33934,N_32273,N_30569);
or U33935 (N_33935,N_30495,N_31719);
nor U33936 (N_33936,N_30088,N_31953);
nand U33937 (N_33937,N_31466,N_31718);
and U33938 (N_33938,N_30584,N_30938);
or U33939 (N_33939,N_31609,N_32461);
xnor U33940 (N_33940,N_30120,N_31970);
and U33941 (N_33941,N_32307,N_30527);
or U33942 (N_33942,N_30487,N_31981);
xor U33943 (N_33943,N_30001,N_31800);
nor U33944 (N_33944,N_30913,N_30030);
nor U33945 (N_33945,N_32012,N_32061);
nor U33946 (N_33946,N_30729,N_30612);
and U33947 (N_33947,N_31586,N_30997);
nor U33948 (N_33948,N_31861,N_31105);
or U33949 (N_33949,N_31118,N_31834);
nor U33950 (N_33950,N_30580,N_31567);
or U33951 (N_33951,N_30142,N_31275);
and U33952 (N_33952,N_30507,N_31632);
and U33953 (N_33953,N_30233,N_30430);
nor U33954 (N_33954,N_31045,N_31899);
nor U33955 (N_33955,N_32457,N_30680);
xnor U33956 (N_33956,N_31601,N_30032);
xnor U33957 (N_33957,N_32182,N_31457);
and U33958 (N_33958,N_31867,N_31152);
nor U33959 (N_33959,N_32061,N_30794);
nand U33960 (N_33960,N_30928,N_32023);
or U33961 (N_33961,N_31324,N_30005);
xnor U33962 (N_33962,N_31322,N_32230);
nor U33963 (N_33963,N_31600,N_31932);
or U33964 (N_33964,N_31147,N_30214);
and U33965 (N_33965,N_31819,N_30460);
and U33966 (N_33966,N_31346,N_31886);
nor U33967 (N_33967,N_31225,N_31485);
nor U33968 (N_33968,N_31216,N_31631);
nand U33969 (N_33969,N_30385,N_30891);
xor U33970 (N_33970,N_30540,N_31304);
nor U33971 (N_33971,N_30925,N_30079);
and U33972 (N_33972,N_32183,N_30843);
nor U33973 (N_33973,N_32067,N_32069);
and U33974 (N_33974,N_31956,N_32063);
and U33975 (N_33975,N_31198,N_31359);
xnor U33976 (N_33976,N_30425,N_31321);
or U33977 (N_33977,N_30801,N_31595);
nor U33978 (N_33978,N_30944,N_31995);
xnor U33979 (N_33979,N_31252,N_30432);
and U33980 (N_33980,N_32322,N_31967);
nor U33981 (N_33981,N_32225,N_31327);
nand U33982 (N_33982,N_32147,N_30855);
or U33983 (N_33983,N_32262,N_30197);
or U33984 (N_33984,N_30715,N_30269);
and U33985 (N_33985,N_30486,N_30316);
nor U33986 (N_33986,N_30665,N_30098);
nand U33987 (N_33987,N_30116,N_30368);
and U33988 (N_33988,N_30184,N_30911);
nand U33989 (N_33989,N_31400,N_32417);
or U33990 (N_33990,N_31047,N_30021);
nand U33991 (N_33991,N_31352,N_30024);
and U33992 (N_33992,N_31015,N_30547);
nor U33993 (N_33993,N_31530,N_31418);
or U33994 (N_33994,N_32060,N_30800);
and U33995 (N_33995,N_32467,N_31060);
or U33996 (N_33996,N_30642,N_31800);
nor U33997 (N_33997,N_32305,N_31770);
xor U33998 (N_33998,N_30466,N_31965);
nor U33999 (N_33999,N_31063,N_31938);
xor U34000 (N_34000,N_31362,N_30427);
xor U34001 (N_34001,N_32151,N_30881);
nand U34002 (N_34002,N_32084,N_32330);
xnor U34003 (N_34003,N_31326,N_31511);
nor U34004 (N_34004,N_31186,N_31079);
nand U34005 (N_34005,N_31384,N_30906);
or U34006 (N_34006,N_30669,N_31221);
nor U34007 (N_34007,N_30914,N_30240);
xnor U34008 (N_34008,N_32379,N_30575);
or U34009 (N_34009,N_31266,N_31076);
and U34010 (N_34010,N_31616,N_31088);
nand U34011 (N_34011,N_32158,N_31471);
nand U34012 (N_34012,N_32409,N_30599);
and U34013 (N_34013,N_31771,N_30435);
nand U34014 (N_34014,N_32456,N_31503);
or U34015 (N_34015,N_30734,N_31131);
nor U34016 (N_34016,N_31352,N_30661);
and U34017 (N_34017,N_31437,N_32090);
nand U34018 (N_34018,N_30345,N_32154);
nand U34019 (N_34019,N_31314,N_32127);
xor U34020 (N_34020,N_31654,N_30095);
nand U34021 (N_34021,N_31919,N_30894);
xnor U34022 (N_34022,N_30513,N_31694);
nand U34023 (N_34023,N_30807,N_30718);
xnor U34024 (N_34024,N_30531,N_31430);
and U34025 (N_34025,N_31468,N_31233);
xor U34026 (N_34026,N_30386,N_31110);
and U34027 (N_34027,N_30357,N_30350);
nor U34028 (N_34028,N_30726,N_30708);
nor U34029 (N_34029,N_32366,N_31274);
xnor U34030 (N_34030,N_32350,N_30212);
nand U34031 (N_34031,N_32000,N_31969);
xor U34032 (N_34032,N_31453,N_31974);
nor U34033 (N_34033,N_30976,N_32451);
xor U34034 (N_34034,N_31710,N_31661);
nor U34035 (N_34035,N_31759,N_32332);
xnor U34036 (N_34036,N_31404,N_31836);
xor U34037 (N_34037,N_30754,N_31775);
nor U34038 (N_34038,N_30957,N_31172);
xnor U34039 (N_34039,N_31531,N_30954);
xor U34040 (N_34040,N_32448,N_31274);
xnor U34041 (N_34041,N_30577,N_31000);
nand U34042 (N_34042,N_31504,N_30825);
and U34043 (N_34043,N_31712,N_32303);
xor U34044 (N_34044,N_30878,N_32353);
nor U34045 (N_34045,N_30766,N_31558);
or U34046 (N_34046,N_30623,N_31734);
xnor U34047 (N_34047,N_30002,N_31826);
xor U34048 (N_34048,N_30460,N_31079);
or U34049 (N_34049,N_32147,N_31933);
or U34050 (N_34050,N_30932,N_31650);
xor U34051 (N_34051,N_32124,N_31297);
and U34052 (N_34052,N_30601,N_31456);
or U34053 (N_34053,N_31685,N_30100);
xor U34054 (N_34054,N_31421,N_32205);
nand U34055 (N_34055,N_31971,N_32271);
nor U34056 (N_34056,N_31462,N_32454);
or U34057 (N_34057,N_31122,N_31564);
nor U34058 (N_34058,N_30956,N_30715);
xor U34059 (N_34059,N_31021,N_30880);
nand U34060 (N_34060,N_30210,N_30957);
nor U34061 (N_34061,N_31840,N_30322);
or U34062 (N_34062,N_32320,N_31067);
nand U34063 (N_34063,N_31372,N_31004);
nand U34064 (N_34064,N_31041,N_30982);
xnor U34065 (N_34065,N_32392,N_32154);
or U34066 (N_34066,N_30559,N_30455);
nand U34067 (N_34067,N_30091,N_30810);
or U34068 (N_34068,N_32183,N_31250);
nor U34069 (N_34069,N_30852,N_30982);
nand U34070 (N_34070,N_32122,N_30066);
nor U34071 (N_34071,N_30511,N_32200);
xnor U34072 (N_34072,N_31708,N_30185);
nand U34073 (N_34073,N_32015,N_32468);
nor U34074 (N_34074,N_31512,N_31474);
xor U34075 (N_34075,N_31865,N_31541);
xor U34076 (N_34076,N_30903,N_31505);
xor U34077 (N_34077,N_31746,N_30260);
nand U34078 (N_34078,N_32330,N_32059);
xor U34079 (N_34079,N_31973,N_30321);
nand U34080 (N_34080,N_31115,N_30977);
nor U34081 (N_34081,N_30887,N_31708);
nand U34082 (N_34082,N_30453,N_30214);
nand U34083 (N_34083,N_31023,N_31277);
xnor U34084 (N_34084,N_31757,N_30737);
and U34085 (N_34085,N_30520,N_30299);
nand U34086 (N_34086,N_31477,N_32057);
or U34087 (N_34087,N_30060,N_32371);
xor U34088 (N_34088,N_30800,N_30072);
nand U34089 (N_34089,N_32113,N_31451);
xor U34090 (N_34090,N_32251,N_31937);
xor U34091 (N_34091,N_32323,N_30558);
and U34092 (N_34092,N_32317,N_30573);
nand U34093 (N_34093,N_30049,N_31557);
nor U34094 (N_34094,N_32143,N_31402);
or U34095 (N_34095,N_32299,N_31811);
nor U34096 (N_34096,N_31725,N_30576);
nand U34097 (N_34097,N_31218,N_31478);
xor U34098 (N_34098,N_31627,N_30381);
nand U34099 (N_34099,N_30307,N_31172);
xnor U34100 (N_34100,N_31719,N_31772);
xor U34101 (N_34101,N_31078,N_32420);
nor U34102 (N_34102,N_30975,N_31222);
nor U34103 (N_34103,N_30626,N_31055);
nor U34104 (N_34104,N_31224,N_31083);
nor U34105 (N_34105,N_31933,N_31324);
or U34106 (N_34106,N_30282,N_31999);
and U34107 (N_34107,N_31789,N_30658);
xor U34108 (N_34108,N_30097,N_30491);
nand U34109 (N_34109,N_31609,N_30347);
nand U34110 (N_34110,N_31368,N_31527);
xnor U34111 (N_34111,N_32017,N_32127);
nor U34112 (N_34112,N_30496,N_31407);
and U34113 (N_34113,N_30750,N_30056);
xnor U34114 (N_34114,N_32292,N_31841);
or U34115 (N_34115,N_32247,N_31933);
or U34116 (N_34116,N_30283,N_30649);
and U34117 (N_34117,N_31268,N_30298);
nand U34118 (N_34118,N_31103,N_30313);
and U34119 (N_34119,N_31120,N_31704);
nand U34120 (N_34120,N_31508,N_31942);
and U34121 (N_34121,N_30506,N_31521);
nand U34122 (N_34122,N_30848,N_32107);
nor U34123 (N_34123,N_30786,N_32342);
and U34124 (N_34124,N_31848,N_32043);
and U34125 (N_34125,N_30193,N_30086);
xor U34126 (N_34126,N_31202,N_31795);
nor U34127 (N_34127,N_31315,N_30327);
xnor U34128 (N_34128,N_30714,N_30606);
nand U34129 (N_34129,N_32351,N_32359);
or U34130 (N_34130,N_31253,N_31190);
nand U34131 (N_34131,N_32367,N_31358);
and U34132 (N_34132,N_30094,N_32282);
or U34133 (N_34133,N_30186,N_32445);
nor U34134 (N_34134,N_30935,N_30302);
and U34135 (N_34135,N_32112,N_30565);
nand U34136 (N_34136,N_31179,N_31390);
nand U34137 (N_34137,N_31132,N_31528);
and U34138 (N_34138,N_30370,N_30327);
xor U34139 (N_34139,N_31781,N_30826);
and U34140 (N_34140,N_30012,N_31965);
nor U34141 (N_34141,N_30567,N_30430);
and U34142 (N_34142,N_31577,N_31135);
and U34143 (N_34143,N_30203,N_30727);
and U34144 (N_34144,N_30188,N_30728);
xor U34145 (N_34145,N_31588,N_30673);
or U34146 (N_34146,N_32264,N_31218);
xor U34147 (N_34147,N_30137,N_31878);
nor U34148 (N_34148,N_30802,N_30947);
nor U34149 (N_34149,N_30002,N_32170);
or U34150 (N_34150,N_31502,N_31762);
or U34151 (N_34151,N_30190,N_30202);
and U34152 (N_34152,N_30309,N_31313);
or U34153 (N_34153,N_32334,N_30498);
and U34154 (N_34154,N_30742,N_30837);
and U34155 (N_34155,N_30703,N_31770);
nand U34156 (N_34156,N_31845,N_31413);
nor U34157 (N_34157,N_31547,N_31456);
and U34158 (N_34158,N_30287,N_31227);
and U34159 (N_34159,N_31587,N_31562);
xnor U34160 (N_34160,N_30750,N_30824);
nor U34161 (N_34161,N_30609,N_30920);
or U34162 (N_34162,N_31730,N_30494);
nand U34163 (N_34163,N_31417,N_32147);
nor U34164 (N_34164,N_30780,N_31454);
nor U34165 (N_34165,N_31256,N_32428);
nor U34166 (N_34166,N_30431,N_30818);
or U34167 (N_34167,N_30652,N_31728);
nand U34168 (N_34168,N_30401,N_31961);
xnor U34169 (N_34169,N_31344,N_32039);
nand U34170 (N_34170,N_30725,N_31861);
and U34171 (N_34171,N_30818,N_31676);
nand U34172 (N_34172,N_32042,N_31109);
or U34173 (N_34173,N_30969,N_31243);
or U34174 (N_34174,N_32160,N_30985);
nand U34175 (N_34175,N_31313,N_31205);
and U34176 (N_34176,N_31460,N_30422);
and U34177 (N_34177,N_30567,N_32236);
nand U34178 (N_34178,N_30436,N_30806);
or U34179 (N_34179,N_30296,N_31371);
and U34180 (N_34180,N_32471,N_30868);
nand U34181 (N_34181,N_32361,N_31990);
nand U34182 (N_34182,N_32237,N_31657);
and U34183 (N_34183,N_31531,N_31076);
xor U34184 (N_34184,N_30788,N_31973);
or U34185 (N_34185,N_30228,N_31905);
and U34186 (N_34186,N_30894,N_31248);
xor U34187 (N_34187,N_32448,N_30662);
and U34188 (N_34188,N_31123,N_31605);
nand U34189 (N_34189,N_30901,N_31609);
nor U34190 (N_34190,N_30466,N_30213);
or U34191 (N_34191,N_30132,N_31898);
nand U34192 (N_34192,N_32211,N_31796);
or U34193 (N_34193,N_31505,N_32230);
or U34194 (N_34194,N_31073,N_30437);
nor U34195 (N_34195,N_32461,N_30031);
xor U34196 (N_34196,N_31087,N_31212);
and U34197 (N_34197,N_30854,N_31632);
nor U34198 (N_34198,N_31396,N_31321);
xnor U34199 (N_34199,N_30136,N_31042);
or U34200 (N_34200,N_30431,N_30944);
xnor U34201 (N_34201,N_31086,N_31008);
or U34202 (N_34202,N_32244,N_30993);
or U34203 (N_34203,N_30109,N_30634);
xor U34204 (N_34204,N_32157,N_32113);
or U34205 (N_34205,N_32189,N_31433);
nor U34206 (N_34206,N_30237,N_30038);
or U34207 (N_34207,N_30817,N_30073);
xnor U34208 (N_34208,N_32358,N_31649);
or U34209 (N_34209,N_30656,N_30271);
xnor U34210 (N_34210,N_31792,N_30694);
or U34211 (N_34211,N_30195,N_31190);
xor U34212 (N_34212,N_31164,N_32219);
xnor U34213 (N_34213,N_30812,N_30933);
xor U34214 (N_34214,N_32034,N_32223);
and U34215 (N_34215,N_30499,N_31963);
or U34216 (N_34216,N_30953,N_31406);
xor U34217 (N_34217,N_31012,N_30376);
nor U34218 (N_34218,N_30938,N_32146);
and U34219 (N_34219,N_30934,N_31230);
and U34220 (N_34220,N_30454,N_31591);
nor U34221 (N_34221,N_31021,N_32441);
xnor U34222 (N_34222,N_31756,N_32373);
nand U34223 (N_34223,N_30753,N_32365);
nand U34224 (N_34224,N_32147,N_31992);
and U34225 (N_34225,N_32348,N_31415);
xnor U34226 (N_34226,N_31726,N_31220);
or U34227 (N_34227,N_32277,N_31902);
or U34228 (N_34228,N_30603,N_31575);
nor U34229 (N_34229,N_32129,N_31299);
and U34230 (N_34230,N_31853,N_30730);
nor U34231 (N_34231,N_30537,N_32417);
nand U34232 (N_34232,N_30848,N_31963);
xor U34233 (N_34233,N_30573,N_30069);
and U34234 (N_34234,N_30392,N_31138);
nor U34235 (N_34235,N_31148,N_30451);
or U34236 (N_34236,N_32256,N_31003);
or U34237 (N_34237,N_32308,N_32377);
nand U34238 (N_34238,N_31979,N_31859);
or U34239 (N_34239,N_31704,N_31067);
xor U34240 (N_34240,N_31500,N_31835);
nand U34241 (N_34241,N_31235,N_31261);
nand U34242 (N_34242,N_30928,N_30051);
xor U34243 (N_34243,N_31032,N_32135);
xnor U34244 (N_34244,N_31395,N_30024);
and U34245 (N_34245,N_32452,N_30779);
nand U34246 (N_34246,N_32189,N_31267);
xor U34247 (N_34247,N_30632,N_30625);
xnor U34248 (N_34248,N_31145,N_31639);
or U34249 (N_34249,N_30226,N_31923);
or U34250 (N_34250,N_31698,N_31978);
and U34251 (N_34251,N_31347,N_30525);
xor U34252 (N_34252,N_31566,N_30935);
nor U34253 (N_34253,N_30078,N_31459);
nand U34254 (N_34254,N_32072,N_31216);
xor U34255 (N_34255,N_32316,N_30429);
xnor U34256 (N_34256,N_31273,N_31202);
nor U34257 (N_34257,N_30260,N_30144);
and U34258 (N_34258,N_31776,N_32136);
nor U34259 (N_34259,N_30841,N_31361);
nor U34260 (N_34260,N_31723,N_30422);
or U34261 (N_34261,N_31042,N_32119);
xnor U34262 (N_34262,N_31804,N_30025);
nor U34263 (N_34263,N_31896,N_31507);
nand U34264 (N_34264,N_30159,N_31123);
and U34265 (N_34265,N_31989,N_31005);
nand U34266 (N_34266,N_31399,N_31546);
xor U34267 (N_34267,N_31635,N_32221);
and U34268 (N_34268,N_31378,N_32472);
nor U34269 (N_34269,N_31170,N_31036);
nand U34270 (N_34270,N_30791,N_31718);
and U34271 (N_34271,N_31991,N_31021);
nor U34272 (N_34272,N_32282,N_31291);
nand U34273 (N_34273,N_31400,N_31662);
and U34274 (N_34274,N_30284,N_31629);
and U34275 (N_34275,N_31795,N_32205);
or U34276 (N_34276,N_31303,N_31286);
xnor U34277 (N_34277,N_30889,N_31701);
xnor U34278 (N_34278,N_30554,N_30123);
nor U34279 (N_34279,N_32396,N_31583);
nand U34280 (N_34280,N_31024,N_32403);
or U34281 (N_34281,N_32189,N_30766);
xnor U34282 (N_34282,N_31195,N_30476);
nand U34283 (N_34283,N_30304,N_31032);
nor U34284 (N_34284,N_30899,N_31926);
xor U34285 (N_34285,N_30604,N_32248);
nand U34286 (N_34286,N_32399,N_32212);
and U34287 (N_34287,N_30612,N_31541);
or U34288 (N_34288,N_30384,N_30818);
and U34289 (N_34289,N_31213,N_30175);
and U34290 (N_34290,N_30063,N_32408);
and U34291 (N_34291,N_31923,N_30314);
nand U34292 (N_34292,N_30371,N_32434);
nor U34293 (N_34293,N_30347,N_31003);
and U34294 (N_34294,N_31474,N_30860);
xor U34295 (N_34295,N_31506,N_30288);
nand U34296 (N_34296,N_32082,N_30472);
xnor U34297 (N_34297,N_31114,N_30812);
xnor U34298 (N_34298,N_30811,N_32167);
xor U34299 (N_34299,N_31033,N_31718);
xor U34300 (N_34300,N_30508,N_32180);
nand U34301 (N_34301,N_31784,N_31979);
nor U34302 (N_34302,N_30787,N_30210);
xnor U34303 (N_34303,N_30286,N_31756);
and U34304 (N_34304,N_32353,N_31867);
nand U34305 (N_34305,N_31703,N_30025);
and U34306 (N_34306,N_31387,N_31526);
xor U34307 (N_34307,N_31420,N_30859);
or U34308 (N_34308,N_31278,N_30321);
and U34309 (N_34309,N_30513,N_32321);
xnor U34310 (N_34310,N_30995,N_31698);
and U34311 (N_34311,N_30373,N_32321);
nor U34312 (N_34312,N_31945,N_32159);
and U34313 (N_34313,N_31689,N_32235);
and U34314 (N_34314,N_30763,N_30169);
nand U34315 (N_34315,N_32213,N_32245);
nand U34316 (N_34316,N_32137,N_31034);
and U34317 (N_34317,N_30719,N_30791);
nand U34318 (N_34318,N_30899,N_32450);
xor U34319 (N_34319,N_31101,N_31384);
xor U34320 (N_34320,N_30685,N_31824);
nor U34321 (N_34321,N_31708,N_31418);
and U34322 (N_34322,N_31896,N_32365);
xor U34323 (N_34323,N_30434,N_31056);
or U34324 (N_34324,N_31416,N_30801);
nor U34325 (N_34325,N_30320,N_30394);
or U34326 (N_34326,N_30894,N_30163);
or U34327 (N_34327,N_30959,N_31881);
xor U34328 (N_34328,N_30537,N_30840);
xor U34329 (N_34329,N_31893,N_31849);
or U34330 (N_34330,N_32140,N_31655);
xor U34331 (N_34331,N_32278,N_30392);
nor U34332 (N_34332,N_32120,N_32327);
nor U34333 (N_34333,N_31479,N_31030);
and U34334 (N_34334,N_31556,N_32405);
xnor U34335 (N_34335,N_32483,N_30344);
xor U34336 (N_34336,N_30002,N_31450);
or U34337 (N_34337,N_32118,N_31873);
or U34338 (N_34338,N_31544,N_31029);
xor U34339 (N_34339,N_31352,N_31424);
nand U34340 (N_34340,N_30985,N_31141);
nor U34341 (N_34341,N_31998,N_31484);
and U34342 (N_34342,N_30592,N_30962);
or U34343 (N_34343,N_30993,N_31457);
xor U34344 (N_34344,N_31975,N_30670);
and U34345 (N_34345,N_32483,N_32436);
or U34346 (N_34346,N_31299,N_32439);
nor U34347 (N_34347,N_30586,N_31937);
and U34348 (N_34348,N_31770,N_31332);
or U34349 (N_34349,N_31686,N_31443);
and U34350 (N_34350,N_30105,N_32307);
and U34351 (N_34351,N_30993,N_32449);
and U34352 (N_34352,N_30917,N_30246);
nor U34353 (N_34353,N_32176,N_31988);
nor U34354 (N_34354,N_32445,N_30818);
xnor U34355 (N_34355,N_31342,N_32111);
or U34356 (N_34356,N_30950,N_30871);
nand U34357 (N_34357,N_30738,N_30809);
and U34358 (N_34358,N_30702,N_31359);
xor U34359 (N_34359,N_31410,N_32248);
and U34360 (N_34360,N_30318,N_31925);
nand U34361 (N_34361,N_31703,N_31245);
or U34362 (N_34362,N_31257,N_31607);
nand U34363 (N_34363,N_30453,N_32390);
nor U34364 (N_34364,N_30514,N_30461);
nor U34365 (N_34365,N_32325,N_30881);
and U34366 (N_34366,N_31733,N_31181);
and U34367 (N_34367,N_30170,N_31184);
xnor U34368 (N_34368,N_31809,N_30830);
and U34369 (N_34369,N_30508,N_31451);
nand U34370 (N_34370,N_31630,N_32196);
nor U34371 (N_34371,N_30349,N_30449);
nor U34372 (N_34372,N_31512,N_31371);
xor U34373 (N_34373,N_32037,N_31701);
nor U34374 (N_34374,N_30778,N_31209);
or U34375 (N_34375,N_30232,N_30303);
xnor U34376 (N_34376,N_30060,N_30954);
or U34377 (N_34377,N_31661,N_31319);
nand U34378 (N_34378,N_31075,N_32493);
nand U34379 (N_34379,N_31299,N_31823);
xor U34380 (N_34380,N_31093,N_31350);
nor U34381 (N_34381,N_30834,N_32165);
nand U34382 (N_34382,N_31688,N_31406);
nor U34383 (N_34383,N_30668,N_30290);
nand U34384 (N_34384,N_31068,N_31579);
nor U34385 (N_34385,N_30441,N_30617);
nand U34386 (N_34386,N_30240,N_31850);
or U34387 (N_34387,N_31828,N_30213);
or U34388 (N_34388,N_30394,N_31768);
xor U34389 (N_34389,N_30500,N_30306);
nor U34390 (N_34390,N_31239,N_30794);
xor U34391 (N_34391,N_31076,N_30167);
or U34392 (N_34392,N_32117,N_30769);
nor U34393 (N_34393,N_31948,N_31107);
xor U34394 (N_34394,N_30254,N_30529);
nand U34395 (N_34395,N_31997,N_31761);
xor U34396 (N_34396,N_30018,N_32095);
nand U34397 (N_34397,N_32033,N_30092);
or U34398 (N_34398,N_30589,N_31324);
and U34399 (N_34399,N_30049,N_30466);
or U34400 (N_34400,N_31042,N_31190);
and U34401 (N_34401,N_30544,N_31712);
and U34402 (N_34402,N_31553,N_31006);
nor U34403 (N_34403,N_31639,N_32161);
xnor U34404 (N_34404,N_30349,N_30917);
or U34405 (N_34405,N_30050,N_31538);
and U34406 (N_34406,N_32045,N_32098);
xor U34407 (N_34407,N_32245,N_31067);
and U34408 (N_34408,N_31684,N_30056);
xor U34409 (N_34409,N_31492,N_31208);
and U34410 (N_34410,N_31490,N_30157);
or U34411 (N_34411,N_30206,N_31630);
or U34412 (N_34412,N_31051,N_30727);
or U34413 (N_34413,N_31338,N_30773);
nor U34414 (N_34414,N_31155,N_31134);
or U34415 (N_34415,N_30221,N_32447);
xnor U34416 (N_34416,N_30082,N_30329);
nand U34417 (N_34417,N_30593,N_31367);
xnor U34418 (N_34418,N_32401,N_30930);
or U34419 (N_34419,N_30952,N_31886);
and U34420 (N_34420,N_31307,N_30866);
or U34421 (N_34421,N_30437,N_31066);
xnor U34422 (N_34422,N_31195,N_32319);
xor U34423 (N_34423,N_31960,N_31151);
nand U34424 (N_34424,N_32142,N_32319);
and U34425 (N_34425,N_30808,N_30026);
or U34426 (N_34426,N_32336,N_32175);
nand U34427 (N_34427,N_30233,N_30853);
nor U34428 (N_34428,N_30875,N_30600);
and U34429 (N_34429,N_31513,N_31049);
or U34430 (N_34430,N_30727,N_31708);
xnor U34431 (N_34431,N_30743,N_31191);
and U34432 (N_34432,N_32449,N_32172);
nand U34433 (N_34433,N_31372,N_31497);
nand U34434 (N_34434,N_32187,N_31361);
nand U34435 (N_34435,N_31510,N_31908);
or U34436 (N_34436,N_31660,N_30259);
nand U34437 (N_34437,N_30793,N_31875);
xnor U34438 (N_34438,N_31762,N_32244);
xor U34439 (N_34439,N_31409,N_30480);
or U34440 (N_34440,N_31569,N_30310);
xor U34441 (N_34441,N_31285,N_32083);
nand U34442 (N_34442,N_30080,N_32159);
nand U34443 (N_34443,N_30941,N_30123);
or U34444 (N_34444,N_31724,N_30959);
and U34445 (N_34445,N_30322,N_30492);
or U34446 (N_34446,N_31210,N_30218);
xor U34447 (N_34447,N_31232,N_32488);
nor U34448 (N_34448,N_30817,N_32152);
nand U34449 (N_34449,N_30140,N_32207);
or U34450 (N_34450,N_31468,N_32080);
nand U34451 (N_34451,N_32492,N_31944);
and U34452 (N_34452,N_30798,N_30857);
xor U34453 (N_34453,N_31043,N_30727);
xnor U34454 (N_34454,N_32314,N_30111);
or U34455 (N_34455,N_31350,N_31374);
xor U34456 (N_34456,N_31195,N_30937);
xor U34457 (N_34457,N_30474,N_30305);
nor U34458 (N_34458,N_31449,N_31567);
or U34459 (N_34459,N_31863,N_31916);
nor U34460 (N_34460,N_31013,N_31737);
nor U34461 (N_34461,N_31079,N_31804);
xnor U34462 (N_34462,N_31196,N_30958);
or U34463 (N_34463,N_30646,N_30989);
nor U34464 (N_34464,N_30313,N_30780);
nand U34465 (N_34465,N_31659,N_30537);
xnor U34466 (N_34466,N_32219,N_31410);
or U34467 (N_34467,N_30252,N_31441);
nor U34468 (N_34468,N_31347,N_32278);
or U34469 (N_34469,N_30533,N_30357);
and U34470 (N_34470,N_32097,N_30458);
nand U34471 (N_34471,N_30070,N_31823);
nor U34472 (N_34472,N_31375,N_30503);
xnor U34473 (N_34473,N_32381,N_30822);
nand U34474 (N_34474,N_31129,N_30779);
or U34475 (N_34475,N_30517,N_31578);
nor U34476 (N_34476,N_30940,N_31846);
and U34477 (N_34477,N_30340,N_32116);
and U34478 (N_34478,N_32056,N_32167);
or U34479 (N_34479,N_30023,N_30422);
nor U34480 (N_34480,N_30236,N_30661);
nand U34481 (N_34481,N_31133,N_31286);
or U34482 (N_34482,N_31544,N_32446);
nor U34483 (N_34483,N_31692,N_30538);
nor U34484 (N_34484,N_32489,N_31866);
xor U34485 (N_34485,N_31515,N_30523);
and U34486 (N_34486,N_30840,N_30504);
or U34487 (N_34487,N_30699,N_31992);
nand U34488 (N_34488,N_31170,N_31265);
and U34489 (N_34489,N_30335,N_31288);
nand U34490 (N_34490,N_31791,N_30602);
or U34491 (N_34491,N_30414,N_30310);
or U34492 (N_34492,N_31225,N_31791);
and U34493 (N_34493,N_31847,N_32457);
or U34494 (N_34494,N_32200,N_31645);
xnor U34495 (N_34495,N_31406,N_31713);
nor U34496 (N_34496,N_32377,N_30834);
nand U34497 (N_34497,N_32071,N_30874);
xor U34498 (N_34498,N_31895,N_32299);
xor U34499 (N_34499,N_30721,N_31378);
or U34500 (N_34500,N_31760,N_30932);
or U34501 (N_34501,N_31504,N_31163);
xor U34502 (N_34502,N_32265,N_31306);
or U34503 (N_34503,N_31047,N_30930);
and U34504 (N_34504,N_30802,N_31288);
xor U34505 (N_34505,N_31514,N_31063);
nor U34506 (N_34506,N_30151,N_31165);
or U34507 (N_34507,N_31892,N_30809);
nor U34508 (N_34508,N_30109,N_30316);
and U34509 (N_34509,N_32232,N_30308);
and U34510 (N_34510,N_31179,N_32063);
or U34511 (N_34511,N_32313,N_31480);
and U34512 (N_34512,N_30731,N_30387);
nand U34513 (N_34513,N_30650,N_32339);
or U34514 (N_34514,N_30599,N_30755);
nor U34515 (N_34515,N_32460,N_31767);
and U34516 (N_34516,N_32292,N_32257);
nor U34517 (N_34517,N_31192,N_31535);
nor U34518 (N_34518,N_31339,N_31672);
nand U34519 (N_34519,N_31390,N_32048);
and U34520 (N_34520,N_32018,N_31035);
nand U34521 (N_34521,N_32160,N_32498);
or U34522 (N_34522,N_31610,N_30993);
and U34523 (N_34523,N_30910,N_30277);
nand U34524 (N_34524,N_32237,N_30347);
or U34525 (N_34525,N_31580,N_31127);
or U34526 (N_34526,N_30005,N_31232);
nand U34527 (N_34527,N_31613,N_32015);
and U34528 (N_34528,N_31660,N_30489);
nand U34529 (N_34529,N_31293,N_30189);
xor U34530 (N_34530,N_30725,N_31719);
nand U34531 (N_34531,N_31706,N_30746);
nand U34532 (N_34532,N_31783,N_31848);
or U34533 (N_34533,N_30924,N_30724);
nand U34534 (N_34534,N_31923,N_30338);
or U34535 (N_34535,N_30640,N_32490);
or U34536 (N_34536,N_30687,N_31764);
nor U34537 (N_34537,N_31977,N_32323);
nor U34538 (N_34538,N_30810,N_31272);
nand U34539 (N_34539,N_30234,N_30179);
and U34540 (N_34540,N_32054,N_31052);
nor U34541 (N_34541,N_30476,N_32375);
or U34542 (N_34542,N_31777,N_31899);
nand U34543 (N_34543,N_32029,N_31130);
and U34544 (N_34544,N_31189,N_30040);
xnor U34545 (N_34545,N_31059,N_32260);
and U34546 (N_34546,N_30760,N_31561);
and U34547 (N_34547,N_30614,N_30542);
nand U34548 (N_34548,N_30729,N_31119);
and U34549 (N_34549,N_30236,N_30546);
or U34550 (N_34550,N_32420,N_31164);
xnor U34551 (N_34551,N_31172,N_30472);
xor U34552 (N_34552,N_32056,N_30474);
xnor U34553 (N_34553,N_31574,N_31120);
nor U34554 (N_34554,N_30801,N_31282);
nand U34555 (N_34555,N_32064,N_31135);
and U34556 (N_34556,N_31515,N_31467);
nor U34557 (N_34557,N_31446,N_30122);
and U34558 (N_34558,N_31939,N_30380);
xnor U34559 (N_34559,N_30911,N_31969);
or U34560 (N_34560,N_31847,N_31492);
nor U34561 (N_34561,N_30945,N_32348);
and U34562 (N_34562,N_30786,N_31656);
or U34563 (N_34563,N_31356,N_31479);
nor U34564 (N_34564,N_30637,N_30132);
or U34565 (N_34565,N_31047,N_30795);
nand U34566 (N_34566,N_32151,N_30675);
and U34567 (N_34567,N_32466,N_31742);
xnor U34568 (N_34568,N_32189,N_30527);
nor U34569 (N_34569,N_32457,N_30225);
nor U34570 (N_34570,N_31365,N_30829);
or U34571 (N_34571,N_30455,N_32067);
xor U34572 (N_34572,N_30610,N_31614);
and U34573 (N_34573,N_31021,N_32077);
xnor U34574 (N_34574,N_31280,N_32053);
nand U34575 (N_34575,N_30062,N_32300);
nand U34576 (N_34576,N_30459,N_31259);
nand U34577 (N_34577,N_30235,N_32124);
xor U34578 (N_34578,N_31461,N_30219);
and U34579 (N_34579,N_31252,N_32253);
xor U34580 (N_34580,N_30483,N_32385);
or U34581 (N_34581,N_30765,N_30132);
xnor U34582 (N_34582,N_31391,N_31936);
nor U34583 (N_34583,N_30569,N_32425);
xnor U34584 (N_34584,N_32071,N_31455);
or U34585 (N_34585,N_30720,N_30275);
nor U34586 (N_34586,N_30633,N_31970);
or U34587 (N_34587,N_30259,N_30496);
nand U34588 (N_34588,N_30865,N_31680);
xnor U34589 (N_34589,N_32032,N_30397);
nor U34590 (N_34590,N_30600,N_30509);
or U34591 (N_34591,N_31696,N_32260);
nand U34592 (N_34592,N_32288,N_31117);
nand U34593 (N_34593,N_32064,N_31260);
nor U34594 (N_34594,N_32480,N_31271);
and U34595 (N_34595,N_30480,N_30177);
nor U34596 (N_34596,N_30961,N_32262);
and U34597 (N_34597,N_32112,N_31936);
xnor U34598 (N_34598,N_30323,N_30337);
or U34599 (N_34599,N_30297,N_31033);
xnor U34600 (N_34600,N_30161,N_32300);
or U34601 (N_34601,N_31119,N_31822);
nand U34602 (N_34602,N_32284,N_31212);
or U34603 (N_34603,N_30229,N_31137);
nand U34604 (N_34604,N_31397,N_32150);
nor U34605 (N_34605,N_32121,N_30555);
or U34606 (N_34606,N_30237,N_31031);
xnor U34607 (N_34607,N_32497,N_30096);
or U34608 (N_34608,N_31876,N_31031);
nor U34609 (N_34609,N_32101,N_31598);
or U34610 (N_34610,N_31426,N_31051);
or U34611 (N_34611,N_30062,N_32304);
nand U34612 (N_34612,N_32346,N_30710);
and U34613 (N_34613,N_32225,N_31663);
nand U34614 (N_34614,N_30034,N_30380);
or U34615 (N_34615,N_32341,N_30002);
and U34616 (N_34616,N_32479,N_30368);
and U34617 (N_34617,N_31313,N_30440);
nand U34618 (N_34618,N_31794,N_31360);
nand U34619 (N_34619,N_31007,N_30819);
nor U34620 (N_34620,N_31959,N_30219);
or U34621 (N_34621,N_30468,N_30158);
and U34622 (N_34622,N_30350,N_30108);
and U34623 (N_34623,N_31433,N_30012);
or U34624 (N_34624,N_32150,N_31715);
and U34625 (N_34625,N_32171,N_31495);
or U34626 (N_34626,N_30296,N_31527);
nor U34627 (N_34627,N_31311,N_30589);
xor U34628 (N_34628,N_32396,N_30981);
nand U34629 (N_34629,N_31135,N_30367);
or U34630 (N_34630,N_30817,N_32141);
nand U34631 (N_34631,N_30270,N_31669);
nand U34632 (N_34632,N_31537,N_30980);
or U34633 (N_34633,N_31686,N_30561);
nor U34634 (N_34634,N_32237,N_31079);
nand U34635 (N_34635,N_30489,N_32270);
xnor U34636 (N_34636,N_30293,N_30156);
or U34637 (N_34637,N_31462,N_32427);
nand U34638 (N_34638,N_31610,N_31788);
or U34639 (N_34639,N_31119,N_32124);
xnor U34640 (N_34640,N_32283,N_30149);
or U34641 (N_34641,N_31966,N_30207);
xor U34642 (N_34642,N_31885,N_30849);
nor U34643 (N_34643,N_30388,N_30355);
nor U34644 (N_34644,N_32023,N_30404);
xor U34645 (N_34645,N_31525,N_32266);
or U34646 (N_34646,N_30610,N_31417);
or U34647 (N_34647,N_31379,N_30035);
or U34648 (N_34648,N_31708,N_31792);
nor U34649 (N_34649,N_31544,N_31665);
nand U34650 (N_34650,N_32066,N_31409);
xnor U34651 (N_34651,N_31296,N_32017);
nor U34652 (N_34652,N_32269,N_31472);
xnor U34653 (N_34653,N_31844,N_30344);
nand U34654 (N_34654,N_32307,N_30577);
xor U34655 (N_34655,N_32025,N_30851);
nand U34656 (N_34656,N_30911,N_30101);
nand U34657 (N_34657,N_31534,N_30462);
or U34658 (N_34658,N_30241,N_30120);
nor U34659 (N_34659,N_31938,N_30595);
and U34660 (N_34660,N_30997,N_30668);
nor U34661 (N_34661,N_30904,N_31188);
or U34662 (N_34662,N_30093,N_30105);
or U34663 (N_34663,N_31642,N_31596);
xnor U34664 (N_34664,N_30847,N_30051);
and U34665 (N_34665,N_30278,N_31895);
nand U34666 (N_34666,N_30303,N_31269);
xor U34667 (N_34667,N_30565,N_30062);
xnor U34668 (N_34668,N_30783,N_31677);
xnor U34669 (N_34669,N_30143,N_32275);
or U34670 (N_34670,N_31106,N_31669);
and U34671 (N_34671,N_31923,N_30229);
xor U34672 (N_34672,N_30561,N_31964);
nand U34673 (N_34673,N_32178,N_32294);
xnor U34674 (N_34674,N_30513,N_32071);
or U34675 (N_34675,N_30059,N_32243);
nand U34676 (N_34676,N_30275,N_31062);
nor U34677 (N_34677,N_30661,N_30899);
nor U34678 (N_34678,N_30687,N_31676);
or U34679 (N_34679,N_31182,N_31568);
or U34680 (N_34680,N_31106,N_32396);
or U34681 (N_34681,N_31389,N_32347);
and U34682 (N_34682,N_30285,N_32460);
nand U34683 (N_34683,N_30497,N_31676);
and U34684 (N_34684,N_32169,N_32275);
nor U34685 (N_34685,N_30403,N_31040);
or U34686 (N_34686,N_31781,N_32423);
or U34687 (N_34687,N_31930,N_30876);
nor U34688 (N_34688,N_31322,N_30031);
nand U34689 (N_34689,N_31895,N_31961);
xnor U34690 (N_34690,N_30051,N_31086);
and U34691 (N_34691,N_30319,N_32331);
or U34692 (N_34692,N_30774,N_32326);
nor U34693 (N_34693,N_31067,N_30248);
or U34694 (N_34694,N_30073,N_32063);
nand U34695 (N_34695,N_32200,N_32424);
or U34696 (N_34696,N_30578,N_32388);
xor U34697 (N_34697,N_31549,N_31299);
nor U34698 (N_34698,N_31724,N_30338);
nor U34699 (N_34699,N_30134,N_31056);
nor U34700 (N_34700,N_31434,N_31777);
nand U34701 (N_34701,N_30311,N_31601);
or U34702 (N_34702,N_31836,N_30117);
and U34703 (N_34703,N_31029,N_31695);
or U34704 (N_34704,N_31223,N_30144);
nand U34705 (N_34705,N_31224,N_30289);
nand U34706 (N_34706,N_30912,N_31915);
nand U34707 (N_34707,N_32003,N_30449);
xor U34708 (N_34708,N_30327,N_30898);
or U34709 (N_34709,N_31176,N_31187);
xor U34710 (N_34710,N_30024,N_31184);
nor U34711 (N_34711,N_30620,N_31628);
xor U34712 (N_34712,N_32416,N_31084);
nor U34713 (N_34713,N_31781,N_30227);
nor U34714 (N_34714,N_31758,N_32110);
and U34715 (N_34715,N_30228,N_30836);
nor U34716 (N_34716,N_30568,N_31598);
xnor U34717 (N_34717,N_31976,N_30703);
or U34718 (N_34718,N_31236,N_31996);
nand U34719 (N_34719,N_30768,N_31543);
xnor U34720 (N_34720,N_31110,N_30472);
nor U34721 (N_34721,N_30372,N_32384);
and U34722 (N_34722,N_30273,N_32299);
and U34723 (N_34723,N_32239,N_31273);
and U34724 (N_34724,N_32223,N_31681);
or U34725 (N_34725,N_30720,N_30984);
xor U34726 (N_34726,N_32443,N_32217);
xor U34727 (N_34727,N_32094,N_31268);
or U34728 (N_34728,N_32133,N_30640);
or U34729 (N_34729,N_31194,N_30603);
or U34730 (N_34730,N_30730,N_30334);
and U34731 (N_34731,N_31844,N_31274);
and U34732 (N_34732,N_31233,N_30586);
nor U34733 (N_34733,N_32006,N_32173);
nor U34734 (N_34734,N_32099,N_30559);
xor U34735 (N_34735,N_31912,N_31099);
nor U34736 (N_34736,N_30506,N_31023);
xor U34737 (N_34737,N_30733,N_30966);
xnor U34738 (N_34738,N_30740,N_30008);
xnor U34739 (N_34739,N_30951,N_31657);
xor U34740 (N_34740,N_31866,N_31550);
xor U34741 (N_34741,N_31592,N_30974);
xor U34742 (N_34742,N_31438,N_30118);
and U34743 (N_34743,N_31024,N_31484);
nand U34744 (N_34744,N_32037,N_30545);
or U34745 (N_34745,N_32355,N_30628);
nand U34746 (N_34746,N_31986,N_31106);
and U34747 (N_34747,N_32477,N_31739);
nor U34748 (N_34748,N_31438,N_32021);
xnor U34749 (N_34749,N_31166,N_31469);
nor U34750 (N_34750,N_30972,N_31428);
nand U34751 (N_34751,N_32284,N_31923);
nand U34752 (N_34752,N_30394,N_31220);
nand U34753 (N_34753,N_31888,N_31367);
or U34754 (N_34754,N_30431,N_30919);
xnor U34755 (N_34755,N_30646,N_30948);
nand U34756 (N_34756,N_30391,N_30683);
and U34757 (N_34757,N_30426,N_31933);
nand U34758 (N_34758,N_30158,N_30532);
nand U34759 (N_34759,N_32136,N_31402);
nor U34760 (N_34760,N_31501,N_31583);
nand U34761 (N_34761,N_30473,N_30736);
xor U34762 (N_34762,N_31739,N_32343);
or U34763 (N_34763,N_32490,N_32405);
or U34764 (N_34764,N_31725,N_30386);
and U34765 (N_34765,N_30259,N_30173);
and U34766 (N_34766,N_31726,N_30355);
nand U34767 (N_34767,N_30106,N_32481);
nand U34768 (N_34768,N_32057,N_32462);
or U34769 (N_34769,N_31236,N_31826);
nor U34770 (N_34770,N_30336,N_31514);
nand U34771 (N_34771,N_30552,N_31315);
and U34772 (N_34772,N_30516,N_31471);
nor U34773 (N_34773,N_32194,N_31834);
xor U34774 (N_34774,N_31342,N_31543);
or U34775 (N_34775,N_31746,N_32182);
nor U34776 (N_34776,N_30504,N_30501);
nor U34777 (N_34777,N_31238,N_32135);
and U34778 (N_34778,N_30481,N_32180);
nand U34779 (N_34779,N_30260,N_30442);
xor U34780 (N_34780,N_30158,N_30181);
xor U34781 (N_34781,N_31002,N_31387);
nor U34782 (N_34782,N_30083,N_30427);
nand U34783 (N_34783,N_31584,N_30598);
xor U34784 (N_34784,N_31958,N_30066);
and U34785 (N_34785,N_30361,N_31625);
nand U34786 (N_34786,N_32229,N_31732);
nor U34787 (N_34787,N_31877,N_30841);
or U34788 (N_34788,N_30502,N_32276);
nor U34789 (N_34789,N_30676,N_31896);
or U34790 (N_34790,N_31767,N_30925);
nand U34791 (N_34791,N_30804,N_31705);
or U34792 (N_34792,N_31069,N_32495);
xnor U34793 (N_34793,N_31853,N_32002);
or U34794 (N_34794,N_30915,N_30295);
and U34795 (N_34795,N_31000,N_31649);
nor U34796 (N_34796,N_30987,N_32440);
or U34797 (N_34797,N_30817,N_30151);
nor U34798 (N_34798,N_30002,N_31348);
or U34799 (N_34799,N_30565,N_32008);
xor U34800 (N_34800,N_31805,N_31049);
or U34801 (N_34801,N_31196,N_31956);
and U34802 (N_34802,N_32288,N_31490);
nand U34803 (N_34803,N_31753,N_30776);
xor U34804 (N_34804,N_30930,N_30643);
nand U34805 (N_34805,N_30673,N_32063);
or U34806 (N_34806,N_30459,N_32096);
nor U34807 (N_34807,N_31197,N_31281);
nand U34808 (N_34808,N_31605,N_31105);
xor U34809 (N_34809,N_30659,N_30979);
nor U34810 (N_34810,N_32393,N_32438);
xor U34811 (N_34811,N_31105,N_31286);
nand U34812 (N_34812,N_30841,N_30934);
xor U34813 (N_34813,N_31986,N_30484);
and U34814 (N_34814,N_30182,N_32253);
or U34815 (N_34815,N_32185,N_30509);
nand U34816 (N_34816,N_30861,N_32075);
or U34817 (N_34817,N_31537,N_30263);
and U34818 (N_34818,N_31205,N_31672);
or U34819 (N_34819,N_30549,N_32290);
or U34820 (N_34820,N_31312,N_30686);
and U34821 (N_34821,N_31311,N_32194);
xor U34822 (N_34822,N_30101,N_31225);
or U34823 (N_34823,N_32178,N_31039);
nor U34824 (N_34824,N_30711,N_30026);
nand U34825 (N_34825,N_30014,N_32445);
nand U34826 (N_34826,N_30343,N_30292);
nand U34827 (N_34827,N_31631,N_31983);
xnor U34828 (N_34828,N_31756,N_30140);
nand U34829 (N_34829,N_31090,N_30876);
nand U34830 (N_34830,N_30463,N_31609);
or U34831 (N_34831,N_31442,N_31615);
xor U34832 (N_34832,N_30317,N_30571);
or U34833 (N_34833,N_32108,N_30209);
nor U34834 (N_34834,N_31885,N_31530);
or U34835 (N_34835,N_31436,N_31361);
nand U34836 (N_34836,N_30539,N_31134);
nand U34837 (N_34837,N_32363,N_31540);
nand U34838 (N_34838,N_31076,N_30315);
and U34839 (N_34839,N_31642,N_30285);
nor U34840 (N_34840,N_30834,N_30685);
and U34841 (N_34841,N_32143,N_32402);
and U34842 (N_34842,N_31142,N_31981);
or U34843 (N_34843,N_31377,N_31786);
xor U34844 (N_34844,N_31729,N_30259);
or U34845 (N_34845,N_31595,N_30163);
and U34846 (N_34846,N_30381,N_32205);
nor U34847 (N_34847,N_30509,N_31454);
nor U34848 (N_34848,N_30469,N_31150);
nand U34849 (N_34849,N_30021,N_30906);
nand U34850 (N_34850,N_30553,N_32314);
and U34851 (N_34851,N_32471,N_32426);
xor U34852 (N_34852,N_30735,N_32167);
nor U34853 (N_34853,N_30779,N_32004);
or U34854 (N_34854,N_30996,N_32085);
nor U34855 (N_34855,N_32157,N_30557);
xor U34856 (N_34856,N_32399,N_30282);
xnor U34857 (N_34857,N_31221,N_31723);
nand U34858 (N_34858,N_32172,N_30278);
and U34859 (N_34859,N_32319,N_31300);
xor U34860 (N_34860,N_31560,N_31290);
xnor U34861 (N_34861,N_30739,N_31222);
xor U34862 (N_34862,N_30085,N_31663);
xnor U34863 (N_34863,N_30478,N_31156);
nor U34864 (N_34864,N_30644,N_31561);
nor U34865 (N_34865,N_31343,N_31759);
nor U34866 (N_34866,N_30454,N_31585);
or U34867 (N_34867,N_30165,N_31053);
nand U34868 (N_34868,N_31998,N_31770);
or U34869 (N_34869,N_32253,N_30275);
or U34870 (N_34870,N_30248,N_30433);
or U34871 (N_34871,N_31737,N_32343);
or U34872 (N_34872,N_30105,N_30678);
and U34873 (N_34873,N_30497,N_30070);
and U34874 (N_34874,N_30960,N_31961);
or U34875 (N_34875,N_31241,N_32052);
nor U34876 (N_34876,N_31353,N_31402);
and U34877 (N_34877,N_32089,N_30424);
or U34878 (N_34878,N_30300,N_30284);
xor U34879 (N_34879,N_30174,N_30387);
or U34880 (N_34880,N_30678,N_30330);
or U34881 (N_34881,N_31817,N_31324);
nand U34882 (N_34882,N_32265,N_31218);
xnor U34883 (N_34883,N_31605,N_31941);
and U34884 (N_34884,N_30122,N_31817);
nand U34885 (N_34885,N_30984,N_31515);
nor U34886 (N_34886,N_31638,N_30803);
nand U34887 (N_34887,N_31566,N_31350);
or U34888 (N_34888,N_30670,N_31775);
nand U34889 (N_34889,N_32290,N_31142);
xor U34890 (N_34890,N_30443,N_30409);
nand U34891 (N_34891,N_31549,N_31183);
nor U34892 (N_34892,N_32028,N_32135);
nor U34893 (N_34893,N_32303,N_31488);
or U34894 (N_34894,N_30122,N_31867);
nand U34895 (N_34895,N_31102,N_31659);
nor U34896 (N_34896,N_30255,N_32245);
or U34897 (N_34897,N_32211,N_32432);
nor U34898 (N_34898,N_30036,N_32445);
and U34899 (N_34899,N_30596,N_31348);
nand U34900 (N_34900,N_32276,N_31207);
nand U34901 (N_34901,N_32284,N_31906);
xor U34902 (N_34902,N_31564,N_30627);
and U34903 (N_34903,N_30542,N_31161);
or U34904 (N_34904,N_31232,N_30221);
or U34905 (N_34905,N_30672,N_32247);
xnor U34906 (N_34906,N_31580,N_32097);
nor U34907 (N_34907,N_30868,N_31250);
and U34908 (N_34908,N_30890,N_30872);
nor U34909 (N_34909,N_32244,N_31229);
nor U34910 (N_34910,N_30093,N_32373);
xor U34911 (N_34911,N_32292,N_30369);
xor U34912 (N_34912,N_30984,N_30404);
or U34913 (N_34913,N_32339,N_32417);
and U34914 (N_34914,N_30327,N_32086);
nor U34915 (N_34915,N_30246,N_30568);
or U34916 (N_34916,N_30998,N_31540);
or U34917 (N_34917,N_31808,N_32436);
and U34918 (N_34918,N_30199,N_30879);
and U34919 (N_34919,N_31914,N_31203);
nand U34920 (N_34920,N_30328,N_31966);
or U34921 (N_34921,N_32184,N_31250);
nor U34922 (N_34922,N_31699,N_30345);
nor U34923 (N_34923,N_31902,N_31752);
xnor U34924 (N_34924,N_30524,N_31526);
xor U34925 (N_34925,N_31290,N_30750);
and U34926 (N_34926,N_30998,N_30064);
and U34927 (N_34927,N_32420,N_30424);
nor U34928 (N_34928,N_30447,N_31286);
and U34929 (N_34929,N_31308,N_30530);
or U34930 (N_34930,N_31355,N_30252);
xor U34931 (N_34931,N_31810,N_32249);
nand U34932 (N_34932,N_30407,N_30082);
nand U34933 (N_34933,N_31059,N_32330);
xnor U34934 (N_34934,N_32093,N_31407);
nor U34935 (N_34935,N_30717,N_32114);
nand U34936 (N_34936,N_30218,N_30743);
nor U34937 (N_34937,N_31582,N_30840);
nand U34938 (N_34938,N_31810,N_30799);
nor U34939 (N_34939,N_32270,N_30273);
xor U34940 (N_34940,N_31414,N_30860);
and U34941 (N_34941,N_30331,N_31962);
or U34942 (N_34942,N_30101,N_31410);
xor U34943 (N_34943,N_31741,N_32080);
nor U34944 (N_34944,N_30684,N_30235);
nand U34945 (N_34945,N_32455,N_30048);
nor U34946 (N_34946,N_30336,N_30619);
nor U34947 (N_34947,N_30337,N_31306);
and U34948 (N_34948,N_31123,N_31183);
or U34949 (N_34949,N_31770,N_30437);
nor U34950 (N_34950,N_32255,N_30509);
and U34951 (N_34951,N_30355,N_31532);
nand U34952 (N_34952,N_30392,N_31851);
xor U34953 (N_34953,N_30713,N_31221);
nand U34954 (N_34954,N_31511,N_31201);
nor U34955 (N_34955,N_31683,N_31110);
xnor U34956 (N_34956,N_32126,N_31807);
or U34957 (N_34957,N_31819,N_31221);
xor U34958 (N_34958,N_30832,N_31388);
nand U34959 (N_34959,N_30853,N_30729);
or U34960 (N_34960,N_31528,N_31081);
nand U34961 (N_34961,N_30956,N_32284);
or U34962 (N_34962,N_30601,N_30146);
nor U34963 (N_34963,N_30729,N_30638);
or U34964 (N_34964,N_31196,N_30715);
or U34965 (N_34965,N_30245,N_31981);
or U34966 (N_34966,N_31473,N_30589);
or U34967 (N_34967,N_30369,N_31579);
nand U34968 (N_34968,N_30214,N_31098);
or U34969 (N_34969,N_30462,N_30197);
or U34970 (N_34970,N_30683,N_30759);
and U34971 (N_34971,N_31733,N_31499);
xor U34972 (N_34972,N_30711,N_32114);
xor U34973 (N_34973,N_30779,N_31382);
nand U34974 (N_34974,N_31226,N_31079);
and U34975 (N_34975,N_30680,N_30907);
and U34976 (N_34976,N_30172,N_30805);
and U34977 (N_34977,N_31934,N_31954);
xnor U34978 (N_34978,N_31433,N_31166);
or U34979 (N_34979,N_30131,N_32282);
nand U34980 (N_34980,N_31033,N_31723);
nand U34981 (N_34981,N_31217,N_31835);
and U34982 (N_34982,N_31819,N_32410);
or U34983 (N_34983,N_30284,N_30122);
xor U34984 (N_34984,N_31264,N_31064);
xnor U34985 (N_34985,N_30209,N_30587);
nor U34986 (N_34986,N_30696,N_30691);
or U34987 (N_34987,N_30745,N_31057);
nor U34988 (N_34988,N_31946,N_30819);
nor U34989 (N_34989,N_30091,N_31271);
nor U34990 (N_34990,N_31774,N_32093);
or U34991 (N_34991,N_32090,N_30914);
and U34992 (N_34992,N_30653,N_32035);
nand U34993 (N_34993,N_31104,N_30919);
nor U34994 (N_34994,N_31283,N_31106);
xnor U34995 (N_34995,N_32403,N_30925);
nor U34996 (N_34996,N_31505,N_30071);
and U34997 (N_34997,N_30776,N_30112);
or U34998 (N_34998,N_31257,N_31702);
and U34999 (N_34999,N_30527,N_30788);
nor U35000 (N_35000,N_34051,N_33500);
nand U35001 (N_35001,N_32659,N_33651);
xor U35002 (N_35002,N_33449,N_34898);
nand U35003 (N_35003,N_33970,N_34009);
nor U35004 (N_35004,N_34304,N_34395);
nand U35005 (N_35005,N_33948,N_34241);
nand U35006 (N_35006,N_33698,N_34491);
and U35007 (N_35007,N_33736,N_32913);
and U35008 (N_35008,N_34360,N_33302);
and U35009 (N_35009,N_33501,N_34149);
nand U35010 (N_35010,N_33884,N_34642);
nand U35011 (N_35011,N_34772,N_34374);
xor U35012 (N_35012,N_33504,N_34493);
or U35013 (N_35013,N_34007,N_34072);
or U35014 (N_35014,N_34869,N_32661);
or U35015 (N_35015,N_33706,N_33831);
xnor U35016 (N_35016,N_34544,N_33576);
nand U35017 (N_35017,N_33080,N_33365);
nor U35018 (N_35018,N_33375,N_33180);
and U35019 (N_35019,N_32869,N_32666);
or U35020 (N_35020,N_34895,N_33479);
xor U35021 (N_35021,N_33011,N_34943);
or U35022 (N_35022,N_33029,N_34429);
nor U35023 (N_35023,N_33776,N_33895);
nor U35024 (N_35024,N_33155,N_33799);
and U35025 (N_35025,N_33523,N_34462);
nor U35026 (N_35026,N_32587,N_34680);
and U35027 (N_35027,N_34428,N_33014);
or U35028 (N_35028,N_33280,N_34319);
xor U35029 (N_35029,N_34981,N_34138);
xnor U35030 (N_35030,N_33463,N_33644);
nand U35031 (N_35031,N_33343,N_34970);
nor U35032 (N_35032,N_33245,N_33017);
nand U35033 (N_35033,N_34109,N_34351);
nand U35034 (N_35034,N_33168,N_33646);
or U35035 (N_35035,N_34802,N_33743);
nor U35036 (N_35036,N_34535,N_33596);
xnor U35037 (N_35037,N_32755,N_33927);
nor U35038 (N_35038,N_33385,N_33126);
nand U35039 (N_35039,N_33455,N_33432);
and U35040 (N_35040,N_33147,N_34592);
nor U35041 (N_35041,N_34847,N_32579);
xnor U35042 (N_35042,N_34426,N_34157);
nand U35043 (N_35043,N_33035,N_34466);
and U35044 (N_35044,N_33450,N_32675);
nor U35045 (N_35045,N_32532,N_33827);
xnor U35046 (N_35046,N_33969,N_33728);
nor U35047 (N_35047,N_34040,N_33765);
xnor U35048 (N_35048,N_34906,N_34407);
or U35049 (N_35049,N_34623,N_33384);
and U35050 (N_35050,N_33431,N_32912);
nand U35051 (N_35051,N_34356,N_33727);
nand U35052 (N_35052,N_34490,N_33874);
nand U35053 (N_35053,N_33466,N_34801);
or U35054 (N_35054,N_33770,N_33798);
nand U35055 (N_35055,N_33689,N_34763);
and U35056 (N_35056,N_34749,N_34222);
or U35057 (N_35057,N_33340,N_34261);
or U35058 (N_35058,N_32724,N_32989);
nor U35059 (N_35059,N_34787,N_32616);
nor U35060 (N_35060,N_33067,N_32549);
xor U35061 (N_35061,N_33772,N_33526);
nand U35062 (N_35062,N_32642,N_32542);
xnor U35063 (N_35063,N_32601,N_32538);
xnor U35064 (N_35064,N_34073,N_34103);
or U35065 (N_35065,N_34412,N_33634);
xnor U35066 (N_35066,N_34856,N_32737);
nor U35067 (N_35067,N_34722,N_34648);
nor U35068 (N_35068,N_34236,N_33332);
and U35069 (N_35069,N_32888,N_33069);
xor U35070 (N_35070,N_33790,N_34988);
nand U35071 (N_35071,N_34061,N_34067);
nor U35072 (N_35072,N_33879,N_34948);
xor U35073 (N_35073,N_34489,N_34525);
nor U35074 (N_35074,N_34724,N_34510);
nor U35075 (N_35075,N_33809,N_34273);
nand U35076 (N_35076,N_33774,N_33686);
nor U35077 (N_35077,N_32647,N_34287);
and U35078 (N_35078,N_34996,N_32882);
xor U35079 (N_35079,N_33252,N_32685);
and U35080 (N_35080,N_34438,N_33578);
and U35081 (N_35081,N_34101,N_33428);
or U35082 (N_35082,N_32861,N_34574);
nand U35083 (N_35083,N_33996,N_34968);
or U35084 (N_35084,N_34223,N_33172);
nor U35085 (N_35085,N_33543,N_32629);
xor U35086 (N_35086,N_34440,N_33341);
nand U35087 (N_35087,N_33232,N_34916);
nand U35088 (N_35088,N_33064,N_33581);
nand U35089 (N_35089,N_34068,N_32644);
or U35090 (N_35090,N_34899,N_34829);
nor U35091 (N_35091,N_32554,N_34288);
or U35092 (N_35092,N_32613,N_34914);
nor U35093 (N_35093,N_34667,N_34729);
and U35094 (N_35094,N_32658,N_34082);
and U35095 (N_35095,N_34536,N_34566);
nand U35096 (N_35096,N_32756,N_33617);
nor U35097 (N_35097,N_33200,N_33395);
and U35098 (N_35098,N_34352,N_34786);
nand U35099 (N_35099,N_33308,N_32621);
and U35100 (N_35100,N_32653,N_33603);
and U35101 (N_35101,N_34660,N_34366);
nor U35102 (N_35102,N_34714,N_32695);
nor U35103 (N_35103,N_34541,N_33256);
nand U35104 (N_35104,N_33366,N_34283);
nor U35105 (N_35105,N_34056,N_33307);
nand U35106 (N_35106,N_34766,N_32841);
or U35107 (N_35107,N_32997,N_32691);
nor U35108 (N_35108,N_32853,N_34629);
xnor U35109 (N_35109,N_33990,N_33908);
or U35110 (N_35110,N_33701,N_34759);
or U35111 (N_35111,N_33374,N_33606);
nor U35112 (N_35112,N_34591,N_34778);
nor U35113 (N_35113,N_33598,N_33751);
or U35114 (N_35114,N_33718,N_33278);
and U35115 (N_35115,N_34096,N_34839);
nand U35116 (N_35116,N_33199,N_32615);
and U35117 (N_35117,N_34765,N_33009);
nor U35118 (N_35118,N_32609,N_34270);
nor U35119 (N_35119,N_34628,N_34776);
and U35120 (N_35120,N_34310,N_33968);
xnor U35121 (N_35121,N_32707,N_34735);
nor U35122 (N_35122,N_34071,N_33730);
and U35123 (N_35123,N_34214,N_32610);
nor U35124 (N_35124,N_33789,N_32586);
or U35125 (N_35125,N_33091,N_32543);
and U35126 (N_35126,N_34523,N_33135);
or U35127 (N_35127,N_34646,N_33177);
nor U35128 (N_35128,N_34066,N_34882);
or U35129 (N_35129,N_33771,N_33847);
nand U35130 (N_35130,N_33213,N_33136);
or U35131 (N_35131,N_34728,N_32983);
nand U35132 (N_35132,N_32637,N_34922);
and U35133 (N_35133,N_34401,N_34368);
nor U35134 (N_35134,N_33773,N_34432);
nor U35135 (N_35135,N_34285,N_33465);
and U35136 (N_35136,N_33658,N_32598);
nor U35137 (N_35137,N_33854,N_33711);
xor U35138 (N_35138,N_33438,N_34550);
nand U35139 (N_35139,N_34422,N_33978);
or U35140 (N_35140,N_33269,N_34826);
or U35141 (N_35141,N_32725,N_33914);
xor U35142 (N_35142,N_34750,N_33058);
or U35143 (N_35143,N_32844,N_34427);
or U35144 (N_35144,N_32986,N_34833);
and U35145 (N_35145,N_32812,N_32561);
or U35146 (N_35146,N_34297,N_34183);
or U35147 (N_35147,N_32796,N_34411);
nand U35148 (N_35148,N_34569,N_32713);
xnor U35149 (N_35149,N_32995,N_33144);
nand U35150 (N_35150,N_33956,N_34681);
or U35151 (N_35151,N_33670,N_32806);
nand U35152 (N_35152,N_34028,N_33561);
xnor U35153 (N_35153,N_34150,N_34086);
nor U35154 (N_35154,N_32662,N_33247);
nor U35155 (N_35155,N_32577,N_32509);
and U35156 (N_35156,N_32596,N_33806);
nand U35157 (N_35157,N_33319,N_34805);
or U35158 (N_35158,N_32831,N_34713);
nor U35159 (N_35159,N_34572,N_34405);
or U35160 (N_35160,N_32846,N_32619);
xor U35161 (N_35161,N_33983,N_34980);
nand U35162 (N_35162,N_32952,N_34925);
nor U35163 (N_35163,N_34170,N_33794);
xor U35164 (N_35164,N_32593,N_34318);
and U35165 (N_35165,N_32594,N_33132);
and U35166 (N_35166,N_33497,N_33949);
or U35167 (N_35167,N_34142,N_34293);
or U35168 (N_35168,N_34791,N_33249);
xor U35169 (N_35169,N_33190,N_34307);
xor U35170 (N_35170,N_32851,N_34365);
and U35171 (N_35171,N_34348,N_34444);
and U35172 (N_35172,N_34737,N_33807);
and U35173 (N_35173,N_33092,N_34945);
or U35174 (N_35174,N_34121,N_33401);
or U35175 (N_35175,N_34404,N_33995);
nor U35176 (N_35176,N_33584,N_34420);
xnor U35177 (N_35177,N_34865,N_33755);
and U35178 (N_35178,N_33008,N_32575);
and U35179 (N_35179,N_34093,N_33894);
or U35180 (N_35180,N_33070,N_32710);
nor U35181 (N_35181,N_33369,N_34041);
and U35182 (N_35182,N_34091,N_34855);
or U35183 (N_35183,N_33242,N_32809);
xor U35184 (N_35184,N_33943,N_33205);
nor U35185 (N_35185,N_34083,N_34151);
or U35186 (N_35186,N_34389,N_32794);
xnor U35187 (N_35187,N_33417,N_34391);
or U35188 (N_35188,N_34141,N_34050);
or U35189 (N_35189,N_32860,N_33514);
and U35190 (N_35190,N_34036,N_32697);
xnor U35191 (N_35191,N_34232,N_34969);
nand U35192 (N_35192,N_33897,N_34809);
or U35193 (N_35193,N_33019,N_34956);
nor U35194 (N_35194,N_33437,N_34335);
and U35195 (N_35195,N_34709,N_34486);
xor U35196 (N_35196,N_33480,N_34345);
and U35197 (N_35197,N_34676,N_32501);
xor U35198 (N_35198,N_33625,N_33233);
nand U35199 (N_35199,N_33357,N_34530);
and U35200 (N_35200,N_34993,N_33442);
and U35201 (N_35201,N_34022,N_33925);
or U35202 (N_35202,N_34984,N_32772);
nor U35203 (N_35203,N_33193,N_32767);
xor U35204 (N_35204,N_34315,N_33866);
and U35205 (N_35205,N_34617,N_34613);
nor U35206 (N_35206,N_32673,N_34696);
xor U35207 (N_35207,N_33828,N_32514);
xnor U35208 (N_35208,N_33271,N_34218);
nor U35209 (N_35209,N_34099,N_34339);
and U35210 (N_35210,N_33660,N_33468);
or U35211 (N_35211,N_34529,N_33179);
nor U35212 (N_35212,N_34768,N_34894);
and U35213 (N_35213,N_32891,N_32699);
and U35214 (N_35214,N_34363,N_34974);
or U35215 (N_35215,N_33226,N_32742);
xnor U35216 (N_35216,N_34322,N_32605);
and U35217 (N_35217,N_33292,N_34215);
nand U35218 (N_35218,N_33074,N_33477);
or U35219 (N_35219,N_32789,N_33784);
nand U35220 (N_35220,N_32600,N_33492);
nor U35221 (N_35221,N_33682,N_34383);
nor U35222 (N_35222,N_33984,N_34501);
or U35223 (N_35223,N_33344,N_32604);
nand U35224 (N_35224,N_33093,N_33942);
or U35225 (N_35225,N_34048,N_34636);
xor U35226 (N_35226,N_33693,N_34020);
xor U35227 (N_35227,N_33918,N_34282);
or U35228 (N_35228,N_32540,N_34424);
and U35229 (N_35229,N_33766,N_32915);
or U35230 (N_35230,N_33397,N_34834);
nand U35231 (N_35231,N_34890,N_34299);
xor U35232 (N_35232,N_34399,N_33187);
xnor U35233 (N_35233,N_32592,N_33493);
nand U35234 (N_35234,N_34439,N_34519);
nor U35235 (N_35235,N_34732,N_34691);
nor U35236 (N_35236,N_32994,N_33039);
nand U35237 (N_35237,N_33522,N_33961);
or U35238 (N_35238,N_33184,N_34673);
and U35239 (N_35239,N_33315,N_34702);
xnor U35240 (N_35240,N_32674,N_34547);
xnor U35241 (N_35241,N_34131,N_34806);
or U35242 (N_35242,N_33778,N_34777);
and U35243 (N_35243,N_34761,N_34382);
or U35244 (N_35244,N_34447,N_32813);
and U35245 (N_35245,N_34989,N_33294);
xnor U35246 (N_35246,N_33456,N_33464);
and U35247 (N_35247,N_34252,N_33427);
xnor U35248 (N_35248,N_33178,N_34880);
and U35249 (N_35249,N_32611,N_34350);
or U35250 (N_35250,N_34184,N_34197);
nand U35251 (N_35251,N_32558,N_33508);
or U35252 (N_35252,N_34168,N_32907);
nand U35253 (N_35253,N_32832,N_32560);
xor U35254 (N_35254,N_34743,N_33348);
xnor U35255 (N_35255,N_34936,N_33785);
nand U35256 (N_35256,N_33065,N_32784);
nor U35257 (N_35257,N_34478,N_33745);
and U35258 (N_35258,N_34955,N_32749);
and U35259 (N_35259,N_32839,N_34002);
nor U35260 (N_35260,N_33157,N_33704);
nor U35261 (N_35261,N_32889,N_33273);
nand U35262 (N_35262,N_33947,N_33746);
and U35263 (N_35263,N_32706,N_34390);
or U35264 (N_35264,N_34094,N_32816);
and U35265 (N_35265,N_33295,N_34918);
nand U35266 (N_35266,N_34259,N_33687);
nor U35267 (N_35267,N_33933,N_33188);
nand U35268 (N_35268,N_34634,N_32909);
nand U35269 (N_35269,N_33118,N_32655);
xor U35270 (N_35270,N_34615,N_32643);
nand U35271 (N_35271,N_32871,N_34593);
xnor U35272 (N_35272,N_34790,N_32670);
nor U35273 (N_35273,N_33673,N_34556);
nor U35274 (N_35274,N_33243,N_34123);
and U35275 (N_35275,N_33692,N_34699);
xnor U35276 (N_35276,N_34563,N_34461);
nand U35277 (N_35277,N_34954,N_32879);
nand U35278 (N_35278,N_32566,N_33753);
nand U35279 (N_35279,N_34780,N_33000);
nor U35280 (N_35280,N_32897,N_34853);
xor U35281 (N_35281,N_33055,N_33031);
nor U35282 (N_35282,N_32735,N_34627);
or U35283 (N_35283,N_33140,N_32535);
nor U35284 (N_35284,N_34964,N_32572);
xor U35285 (N_35285,N_32720,N_34850);
and U35286 (N_35286,N_34748,N_33360);
xor U35287 (N_35287,N_34888,N_34129);
nor U35288 (N_35288,N_33872,N_33636);
and U35289 (N_35289,N_32625,N_34818);
nand U35290 (N_35290,N_34891,N_34637);
nand U35291 (N_35291,N_34507,N_33461);
and U35292 (N_35292,N_33980,N_32656);
or U35293 (N_35293,N_32555,N_33158);
and U35294 (N_35294,N_34385,N_34862);
and U35295 (N_35295,N_34973,N_32822);
or U35296 (N_35296,N_34276,N_32881);
or U35297 (N_35297,N_32530,N_32632);
or U35298 (N_35298,N_33429,N_33659);
nor U35299 (N_35299,N_32712,N_33703);
xor U35300 (N_35300,N_33439,N_33707);
nor U35301 (N_35301,N_34033,N_34364);
or U35302 (N_35302,N_34561,N_33123);
or U35303 (N_35303,N_33425,N_32526);
nor U35304 (N_35304,N_34941,N_33540);
nand U35305 (N_35305,N_33538,N_33505);
or U35306 (N_35306,N_34586,N_33353);
and U35307 (N_35307,N_32649,N_32719);
nor U35308 (N_35308,N_33619,N_32827);
xor U35309 (N_35309,N_33519,N_33839);
or U35310 (N_35310,N_34124,N_33214);
and U35311 (N_35311,N_32868,N_33222);
nand U35312 (N_35312,N_33648,N_33358);
nand U35313 (N_35313,N_33909,N_33930);
nand U35314 (N_35314,N_33877,N_34597);
nand U35315 (N_35315,N_34418,N_34088);
nand U35316 (N_35316,N_33272,N_33186);
and U35317 (N_35317,N_32534,N_33735);
and U35318 (N_35318,N_33038,N_34187);
and U35319 (N_35319,N_33856,N_32858);
xor U35320 (N_35320,N_33487,N_34957);
or U35321 (N_35321,N_34079,N_34582);
or U35322 (N_35322,N_33221,N_34843);
xor U35323 (N_35323,N_32867,N_33552);
xor U35324 (N_35324,N_32937,N_32834);
xnor U35325 (N_35325,N_33054,N_34603);
nand U35326 (N_35326,N_33414,N_33028);
and U35327 (N_35327,N_32957,N_33734);
nor U35328 (N_35328,N_34433,N_33533);
or U35329 (N_35329,N_34622,N_33881);
or U35330 (N_35330,N_32716,N_33892);
nor U35331 (N_35331,N_32896,N_32793);
or U35332 (N_35332,N_34267,N_33377);
nand U35333 (N_35333,N_33024,N_33104);
and U35334 (N_35334,N_34114,N_33667);
nand U35335 (N_35335,N_33623,N_32503);
nor U35336 (N_35336,N_33853,N_34610);
and U35337 (N_35337,N_33559,N_32739);
or U35338 (N_35338,N_33524,N_33915);
xor U35339 (N_35339,N_33868,N_33732);
or U35340 (N_35340,N_32588,N_32723);
nor U35341 (N_35341,N_34381,N_32802);
or U35342 (N_35342,N_32568,N_33657);
and U35343 (N_35343,N_33601,N_34278);
nand U35344 (N_35344,N_33400,N_32874);
xnor U35345 (N_35345,N_34375,N_32807);
and U35346 (N_35346,N_33708,N_33234);
nand U35347 (N_35347,N_32840,N_33800);
nor U35348 (N_35348,N_33850,N_33590);
nor U35349 (N_35349,N_33217,N_33393);
xnor U35350 (N_35350,N_34137,N_34357);
nand U35351 (N_35351,N_34775,N_33102);
nand U35352 (N_35352,N_34070,N_34528);
xor U35353 (N_35353,N_32582,N_33801);
xnor U35354 (N_35354,N_34122,N_34161);
xnor U35355 (N_35355,N_33237,N_33710);
xor U35356 (N_35356,N_32557,N_33321);
nor U35357 (N_35357,N_32602,N_33599);
and U35358 (N_35358,N_34298,N_33912);
nor U35359 (N_35359,N_33536,N_32968);
xor U35360 (N_35360,N_33904,N_32574);
nor U35361 (N_35361,N_34861,N_34851);
xnor U35362 (N_35362,N_33585,N_34867);
and U35363 (N_35363,N_32933,N_33920);
and U35364 (N_35364,N_33862,N_33629);
nor U35365 (N_35365,N_33460,N_34162);
nor U35366 (N_35366,N_33260,N_33923);
or U35367 (N_35367,N_34308,N_34542);
xnor U35368 (N_35368,N_34408,N_32500);
xnor U35369 (N_35369,N_32977,N_34744);
or U35370 (N_35370,N_34095,N_34499);
nor U35371 (N_35371,N_33027,N_33632);
xor U35372 (N_35372,N_34794,N_33022);
nand U35373 (N_35373,N_33971,N_32581);
and U35374 (N_35374,N_33472,N_34309);
xor U35375 (N_35375,N_34338,N_34224);
nor U35376 (N_35376,N_32519,N_33394);
xor U35377 (N_35377,N_33173,N_34125);
and U35378 (N_35378,N_33720,N_33363);
and U35379 (N_35379,N_33309,N_33499);
nor U35380 (N_35380,N_34576,N_32630);
or U35381 (N_35381,N_33901,N_32781);
nand U35382 (N_35382,N_32981,N_33210);
nand U35383 (N_35383,N_33435,N_33840);
and U35384 (N_35384,N_34192,N_33457);
and U35385 (N_35385,N_33891,N_34175);
xnor U35386 (N_35386,N_33001,N_33715);
and U35387 (N_35387,N_33724,N_34211);
nand U35388 (N_35388,N_34717,N_33317);
nand U35389 (N_35389,N_33835,N_34171);
nand U35390 (N_35390,N_33525,N_34746);
nand U35391 (N_35391,N_34396,N_32967);
or U35392 (N_35392,N_34872,N_34739);
and U35393 (N_35393,N_34479,N_33905);
nand U35394 (N_35394,N_33935,N_34024);
nand U35395 (N_35395,N_33287,N_33851);
and U35396 (N_35396,N_33580,N_33081);
xnor U35397 (N_35397,N_32898,N_34431);
nand U35398 (N_35398,N_32664,N_34392);
and U35399 (N_35399,N_34147,N_32761);
or U35400 (N_35400,N_32790,N_34182);
and U35401 (N_35401,N_33422,N_33462);
nand U35402 (N_35402,N_34231,N_33495);
xor U35403 (N_35403,N_33575,N_33227);
xor U35404 (N_35404,N_33577,N_32504);
and U35405 (N_35405,N_33645,N_32550);
and U35406 (N_35406,N_34130,N_34679);
and U35407 (N_35407,N_34081,N_32777);
nor U35408 (N_35408,N_34609,N_34303);
nor U35409 (N_35409,N_34376,N_34112);
or U35410 (N_35410,N_34860,N_32931);
and U35411 (N_35411,N_33822,N_33593);
and U35412 (N_35412,N_34706,N_33787);
nand U35413 (N_35413,N_32899,N_34233);
xor U35414 (N_35414,N_32750,N_33434);
or U35415 (N_35415,N_34032,N_32506);
nor U35416 (N_35416,N_34238,N_32734);
nand U35417 (N_35417,N_34783,N_32961);
or U35418 (N_35418,N_33663,N_34008);
and U35419 (N_35419,N_33758,N_34935);
nand U35420 (N_35420,N_33808,N_33383);
or U35421 (N_35421,N_34997,N_34027);
xnor U35422 (N_35422,N_34716,N_33826);
and U35423 (N_35423,N_33824,N_32752);
nor U35424 (N_35424,N_33007,N_33129);
and U35425 (N_35425,N_34452,N_34484);
and U35426 (N_35426,N_33446,N_34558);
nand U35427 (N_35427,N_33289,N_34849);
nor U35428 (N_35428,N_34191,N_33907);
nand U35429 (N_35429,N_32580,N_32786);
xor U35430 (N_35430,N_33324,N_33313);
xor U35431 (N_35431,N_33056,N_34858);
and U35432 (N_35432,N_32631,N_33231);
nor U35433 (N_35433,N_33113,N_33541);
nor U35434 (N_35434,N_32985,N_33328);
nor U35435 (N_35435,N_34471,N_33631);
xor U35436 (N_35436,N_34459,N_34864);
and U35437 (N_35437,N_34111,N_33690);
xnor U35438 (N_35438,N_33640,N_32792);
nor U35439 (N_35439,N_32892,N_34690);
nand U35440 (N_35440,N_33430,N_32953);
or U35441 (N_35441,N_32890,N_32799);
and U35442 (N_35442,N_33026,N_33744);
nand U35443 (N_35443,N_33731,N_33046);
and U35444 (N_35444,N_33875,N_34845);
nor U35445 (N_35445,N_34991,N_34193);
nor U35446 (N_35446,N_33396,N_34155);
nor U35447 (N_35447,N_34902,N_33684);
xor U35448 (N_35448,N_32911,N_33709);
and U35449 (N_35449,N_34979,N_32548);
and U35450 (N_35450,N_34503,N_33496);
nand U35451 (N_35451,N_33305,N_32971);
xnor U35452 (N_35452,N_32824,N_33752);
nand U35453 (N_35453,N_34107,N_34219);
and U35454 (N_35454,N_33254,N_34831);
xor U35455 (N_35455,N_32614,N_34403);
xor U35456 (N_35456,N_33739,N_34965);
and U35457 (N_35457,N_34552,N_34237);
or U35458 (N_35458,N_34506,N_34115);
or U35459 (N_35459,N_33964,N_32964);
or U35460 (N_35460,N_33564,N_34889);
or U35461 (N_35461,N_34460,N_34012);
xor U35462 (N_35462,N_33749,N_33270);
xor U35463 (N_35463,N_34631,N_34837);
and U35464 (N_35464,N_33981,N_34502);
and U35465 (N_35465,N_33005,N_34692);
or U35466 (N_35466,N_33532,N_32797);
nor U35467 (N_35467,N_34718,N_33291);
nor U35468 (N_35468,N_33040,N_33122);
nand U35469 (N_35469,N_33436,N_33481);
nand U35470 (N_35470,N_34240,N_34639);
xor U35471 (N_35471,N_34097,N_33661);
and U35472 (N_35472,N_34075,N_34999);
nand U35473 (N_35473,N_33286,N_33030);
nor U35474 (N_35474,N_34417,N_34788);
nand U35475 (N_35475,N_34291,N_33671);
or U35476 (N_35476,N_32516,N_32754);
and U35477 (N_35477,N_33403,N_33106);
xnor U35478 (N_35478,N_34693,N_33349);
nand U35479 (N_35479,N_33676,N_33662);
nand U35480 (N_35480,N_34146,N_33236);
nand U35481 (N_35481,N_32800,N_34540);
or U35482 (N_35482,N_33379,N_33795);
or U35483 (N_35483,N_34225,N_34173);
nand U35484 (N_35484,N_33721,N_34456);
nand U35485 (N_35485,N_33111,N_32870);
nand U35486 (N_35486,N_34442,N_33890);
nand U35487 (N_35487,N_32830,N_34004);
or U35488 (N_35488,N_34458,N_33107);
xnor U35489 (N_35489,N_33966,N_34377);
or U35490 (N_35490,N_32717,N_33351);
nor U35491 (N_35491,N_34100,N_34758);
and U35492 (N_35492,N_34437,N_33627);
nor U35493 (N_35493,N_33791,N_33452);
xor U35494 (N_35494,N_32628,N_34854);
and U35495 (N_35495,N_34167,N_32872);
or U35496 (N_35496,N_32940,N_34723);
or U35497 (N_35497,N_34659,N_33408);
nand U35498 (N_35498,N_34135,N_34824);
xnor U35499 (N_35499,N_34820,N_33006);
xnor U35500 (N_35500,N_33339,N_33392);
or U35501 (N_35501,N_33421,N_32738);
nor U35502 (N_35502,N_32787,N_34455);
and U35503 (N_35503,N_34272,N_34947);
or U35504 (N_35504,N_32608,N_33346);
nand U35505 (N_35505,N_32539,N_32607);
nor U35506 (N_35506,N_33768,N_34423);
and U35507 (N_35507,N_34457,N_33955);
or U35508 (N_35508,N_33697,N_34488);
and U35509 (N_35509,N_33196,N_34796);
and U35510 (N_35510,N_33059,N_32900);
or U35511 (N_35511,N_34688,N_33946);
nor U35512 (N_35512,N_32811,N_34001);
nor U35513 (N_35513,N_34419,N_33078);
and U35514 (N_35514,N_33447,N_32817);
xnor U35515 (N_35515,N_33224,N_34741);
and U35516 (N_35516,N_34654,N_32929);
or U35517 (N_35517,N_32678,N_33467);
xor U35518 (N_35518,N_33124,N_33683);
or U35519 (N_35519,N_33988,N_34355);
and U35520 (N_35520,N_34367,N_33164);
xor U35521 (N_35521,N_32885,N_34799);
and U35522 (N_35522,N_33643,N_34672);
xor U35523 (N_35523,N_34810,N_33620);
or U35524 (N_35524,N_33150,N_32875);
xnor U35525 (N_35525,N_32819,N_34262);
nand U35526 (N_35526,N_34089,N_33259);
nand U35527 (N_35527,N_32565,N_32583);
nor U35528 (N_35528,N_33841,N_33812);
or U35529 (N_35529,N_34624,N_33509);
nand U35530 (N_35530,N_33062,N_33218);
or U35531 (N_35531,N_33846,N_33238);
and U35532 (N_35532,N_33310,N_33757);
xor U35533 (N_35533,N_33386,N_32935);
or U35534 (N_35534,N_34848,N_34934);
xnor U35535 (N_35535,N_32721,N_32842);
and U35536 (N_35536,N_34873,N_33792);
nand U35537 (N_35537,N_32692,N_33865);
nor U35538 (N_35538,N_32783,N_32688);
xor U35539 (N_35539,N_34290,N_34266);
xnor U35540 (N_35540,N_33398,N_33120);
or U35541 (N_35541,N_32718,N_33797);
nor U35542 (N_35542,N_33323,N_34264);
nand U35543 (N_35543,N_32925,N_33285);
nor U35544 (N_35544,N_34521,N_34611);
xnor U35545 (N_35545,N_33032,N_33380);
nor U35546 (N_35546,N_33246,N_34305);
or U35547 (N_35547,N_33268,N_32943);
xor U35548 (N_35548,N_33611,N_34649);
nor U35549 (N_35549,N_32704,N_33228);
or U35550 (N_35550,N_34618,N_33303);
nand U35551 (N_35551,N_32775,N_34406);
and U35552 (N_35552,N_33655,N_33063);
nor U35553 (N_35553,N_34534,N_34413);
or U35554 (N_35554,N_33283,N_34712);
and U35555 (N_35555,N_34887,N_33197);
or U35556 (N_35556,N_34733,N_33694);
and U35557 (N_35557,N_32518,N_33609);
nor U35558 (N_35558,N_33630,N_34059);
nand U35559 (N_35559,N_34573,N_34531);
nor U35560 (N_35560,N_33888,N_32815);
or U35561 (N_35561,N_34752,N_33569);
nor U35562 (N_35562,N_34938,N_33626);
or U35563 (N_35563,N_33691,N_34877);
or U35564 (N_35564,N_32746,N_33999);
or U35565 (N_35565,N_33637,N_34671);
xor U35566 (N_35566,N_34031,N_34274);
or U35567 (N_35567,N_32606,N_34030);
and U35568 (N_35568,N_33608,N_34512);
nand U35569 (N_35569,N_34268,N_32731);
xnor U35570 (N_35570,N_34077,N_33962);
or U35571 (N_35571,N_34409,N_32776);
xnor U35572 (N_35572,N_34526,N_34621);
and U35573 (N_35573,N_33836,N_34035);
and U35574 (N_35574,N_33023,N_33347);
xnor U35575 (N_35575,N_33143,N_32544);
nor U35576 (N_35576,N_32764,N_33068);
or U35577 (N_35577,N_33103,N_33060);
xor U35578 (N_35578,N_33114,N_34156);
nor U35579 (N_35579,N_34015,N_34464);
xnor U35580 (N_35580,N_34978,N_32926);
xnor U35581 (N_35581,N_33327,N_34246);
or U35582 (N_35582,N_33903,N_33502);
nand U35583 (N_35583,N_33858,N_33277);
and U35584 (N_35584,N_33284,N_32627);
or U35585 (N_35585,N_34136,N_34239);
and U35586 (N_35586,N_33041,N_33985);
or U35587 (N_35587,N_32902,N_33959);
or U35588 (N_35588,N_34626,N_32671);
or U35589 (N_35589,N_33253,N_33825);
nand U35590 (N_35590,N_33899,N_33251);
nand U35591 (N_35591,N_32941,N_34651);
or U35592 (N_35592,N_34118,N_34567);
nand U35593 (N_35593,N_33361,N_34279);
nand U35594 (N_35594,N_34370,N_33521);
xnor U35595 (N_35595,N_33473,N_34425);
and U35596 (N_35596,N_33852,N_32904);
nand U35597 (N_35597,N_32733,N_33997);
nor U35598 (N_35598,N_33119,N_34900);
xnor U35599 (N_35599,N_33666,N_34915);
and U35600 (N_35600,N_34052,N_33589);
xnor U35601 (N_35601,N_34960,N_33563);
and U35602 (N_35602,N_34715,N_33716);
or U35603 (N_35603,N_33681,N_33372);
and U35604 (N_35604,N_33583,N_33656);
xnor U35605 (N_35605,N_34811,N_34803);
or U35606 (N_35606,N_33053,N_33202);
xnor U35607 (N_35607,N_34301,N_33079);
xnor U35608 (N_35608,N_32876,N_32980);
nor U35609 (N_35609,N_32970,N_32932);
and U35610 (N_35610,N_32646,N_34117);
and U35611 (N_35611,N_33871,N_33588);
xnor U35612 (N_35612,N_34726,N_33181);
nor U35613 (N_35613,N_34163,N_34316);
xnor U35614 (N_35614,N_34554,N_34140);
and U35615 (N_35615,N_34176,N_32590);
nand U35616 (N_35616,N_33133,N_34325);
and U35617 (N_35617,N_33105,N_32537);
and U35618 (N_35618,N_34816,N_32546);
nor U35619 (N_35619,N_33823,N_34046);
xor U35620 (N_35620,N_34885,N_34711);
xor U35621 (N_35621,N_34913,N_32663);
xnor U35622 (N_35622,N_34509,N_32672);
or U35623 (N_35623,N_34505,N_32623);
nand U35624 (N_35624,N_32591,N_33880);
nor U35625 (N_35625,N_33018,N_34188);
nand U35626 (N_35626,N_34013,N_34359);
xnor U35627 (N_35627,N_34477,N_33973);
nor U35628 (N_35628,N_34812,N_34332);
or U35629 (N_35629,N_33557,N_34284);
nand U35630 (N_35630,N_33117,N_34747);
xnor U35631 (N_35631,N_33156,N_32848);
nand U35632 (N_35632,N_34650,N_32529);
and U35633 (N_35633,N_34703,N_33189);
xnor U35634 (N_35634,N_33818,N_34632);
nand U35635 (N_35635,N_33311,N_32696);
nand U35636 (N_35636,N_33489,N_33849);
nor U35637 (N_35637,N_33515,N_33861);
nand U35638 (N_35638,N_34911,N_32686);
and U35639 (N_35639,N_34705,N_34606);
and U35640 (N_35640,N_33153,N_34292);
or U35641 (N_35641,N_34055,N_33638);
nand U35642 (N_35642,N_34400,N_33312);
or U35643 (N_35643,N_34227,N_33788);
nand U35644 (N_35644,N_34120,N_34021);
or U35645 (N_35645,N_32620,N_32825);
and U35646 (N_35646,N_33902,N_34003);
and U35647 (N_35647,N_32988,N_34972);
and U35648 (N_35648,N_32936,N_33025);
or U35649 (N_35649,N_34946,N_34990);
xnor U35650 (N_35650,N_32877,N_32702);
and U35651 (N_35651,N_33304,N_34588);
nor U35652 (N_35652,N_32744,N_34254);
nand U35653 (N_35653,N_33622,N_33592);
or U35654 (N_35654,N_32798,N_33761);
nand U35655 (N_35655,N_34098,N_32553);
xor U35656 (N_35656,N_34189,N_34148);
nor U35657 (N_35657,N_33607,N_33183);
or U35658 (N_35658,N_34939,N_33116);
nor U35659 (N_35659,N_32657,N_33889);
nand U35660 (N_35660,N_34207,N_34998);
xor U35661 (N_35661,N_33020,N_32836);
xor U35662 (N_35662,N_32828,N_33095);
nor U35663 (N_35663,N_33600,N_34994);
and U35664 (N_35664,N_33331,N_33371);
xor U35665 (N_35665,N_34800,N_32782);
or U35666 (N_35666,N_32563,N_33240);
and U35667 (N_35667,N_33362,N_33987);
and U35668 (N_35668,N_34038,N_33152);
nand U35669 (N_35669,N_34841,N_34242);
and U35670 (N_35670,N_34312,N_33137);
nand U35671 (N_35671,N_33979,N_34194);
nor U35672 (N_35672,N_34463,N_33700);
or U35673 (N_35673,N_33330,N_32771);
xnor U35674 (N_35674,N_34126,N_32595);
xor U35675 (N_35675,N_33510,N_32954);
nand U35676 (N_35676,N_33545,N_34589);
and U35677 (N_35677,N_32573,N_32728);
nand U35678 (N_35678,N_32808,N_33154);
nand U35679 (N_35679,N_33783,N_33021);
xor U35680 (N_35680,N_32585,N_34199);
or U35681 (N_35681,N_34937,N_33857);
and U35682 (N_35682,N_33974,N_33326);
or U35683 (N_35683,N_34983,N_33264);
and U35684 (N_35684,N_33896,N_33354);
and U35685 (N_35685,N_32740,N_34815);
and U35686 (N_35686,N_34108,N_34302);
and U35687 (N_35687,N_33052,N_33931);
xnor U35688 (N_35688,N_33322,N_33329);
and U35689 (N_35689,N_33090,N_33491);
or U35690 (N_35690,N_33878,N_32769);
nand U35691 (N_35691,N_33044,N_34074);
xor U35692 (N_35692,N_32880,N_34575);
xnor U35693 (N_35693,N_32854,N_33516);
nor U35694 (N_35694,N_33953,N_34975);
nor U35695 (N_35695,N_33837,N_34342);
xnor U35696 (N_35696,N_34584,N_34260);
and U35697 (N_35697,N_33911,N_34830);
nor U35698 (N_35698,N_34209,N_33579);
xnor U35699 (N_35699,N_34230,N_34669);
and U35700 (N_35700,N_34604,N_34779);
and U35701 (N_35701,N_33061,N_32965);
nor U35702 (N_35702,N_33399,N_32987);
and U35703 (N_35703,N_32778,N_32682);
nor U35704 (N_35704,N_32753,N_34271);
nand U35705 (N_35705,N_32640,N_33411);
nor U35706 (N_35706,N_32715,N_34344);
nor U35707 (N_35707,N_34663,N_34394);
nand U35708 (N_35708,N_33426,N_34555);
or U35709 (N_35709,N_32622,N_33685);
xnor U35710 (N_35710,N_34220,N_33677);
nand U35711 (N_35711,N_32570,N_34065);
or U35712 (N_35712,N_34480,N_33274);
or U35713 (N_35713,N_33036,N_32773);
nor U35714 (N_35714,N_32559,N_33410);
and U35715 (N_35715,N_33900,N_34879);
and U35716 (N_35716,N_33016,N_33616);
xnor U35717 (N_35717,N_33261,N_33267);
nor U35718 (N_35718,N_34353,N_33571);
xnor U35719 (N_35719,N_34202,N_33618);
or U35720 (N_35720,N_33146,N_34754);
nor U35721 (N_35721,N_34719,N_33364);
nand U35722 (N_35722,N_33076,N_33419);
and U35723 (N_35723,N_32779,N_33674);
nor U35724 (N_35724,N_33537,N_34296);
and U35725 (N_35725,N_32660,N_33169);
xnor U35726 (N_35726,N_34000,N_33420);
xor U35727 (N_35727,N_33474,N_33390);
xnor U35728 (N_35728,N_33729,N_34451);
nand U35729 (N_35729,N_34852,N_33654);
xor U35730 (N_35730,N_34952,N_33649);
and U35731 (N_35731,N_33288,N_34868);
nand U35732 (N_35732,N_34641,N_33071);
and U35733 (N_35733,N_34245,N_33241);
nor U35734 (N_35734,N_33572,N_33042);
nor U35735 (N_35735,N_33747,N_34694);
xnor U35736 (N_35736,N_33597,N_33750);
nand U35737 (N_35737,N_32513,N_34565);
nor U35738 (N_35738,N_32818,N_33203);
xnor U35739 (N_35739,N_33517,N_34710);
xor U35740 (N_35740,N_34084,N_32683);
or U35741 (N_35741,N_33257,N_32669);
nor U35742 (N_35742,N_32886,N_33756);
xnor U35743 (N_35743,N_34619,N_34134);
xor U35744 (N_35744,N_33669,N_34476);
nand U35745 (N_35745,N_32528,N_34443);
nand U35746 (N_35746,N_34295,N_33748);
nand U35747 (N_35747,N_32510,N_33653);
and U35748 (N_35748,N_32770,N_33972);
nor U35749 (N_35749,N_33182,N_34731);
nand U35750 (N_35750,N_32785,N_33805);
xor U35751 (N_35751,N_34515,N_32959);
nor U35752 (N_35752,N_33048,N_34265);
nand U35753 (N_35753,N_33115,N_32684);
nand U35754 (N_35754,N_34745,N_34132);
nand U35755 (N_35755,N_33404,N_34896);
nor U35756 (N_35756,N_33201,N_34992);
nand U35757 (N_35757,N_33567,N_34017);
nor U35758 (N_35758,N_34595,N_32536);
or U35759 (N_35759,N_34119,N_32571);
nand U35760 (N_35760,N_33367,N_33211);
nand U35761 (N_35761,N_32991,N_34682);
and U35762 (N_35762,N_34337,N_33844);
xnor U35763 (N_35763,N_33641,N_33299);
and U35764 (N_35764,N_34919,N_34289);
or U35765 (N_35765,N_34213,N_33565);
nand U35766 (N_35766,N_33586,N_34397);
nand U35767 (N_35767,N_33262,N_34846);
nand U35768 (N_35768,N_34612,N_34323);
and U35769 (N_35769,N_34782,N_32703);
and U35770 (N_35770,N_34961,N_33185);
nor U35771 (N_35771,N_32679,N_33796);
nor U35772 (N_35772,N_32645,N_33216);
nor U35773 (N_35773,N_33086,N_33742);
nand U35774 (N_35774,N_34362,N_34340);
xor U35775 (N_35775,N_34771,N_33388);
and U35776 (N_35776,N_34674,N_34277);
and U35777 (N_35777,N_34212,N_34085);
or U35778 (N_35778,N_32633,N_33845);
and U35779 (N_35779,N_34250,N_34751);
and U35780 (N_35780,N_34630,N_33229);
xnor U35781 (N_35781,N_33356,N_33556);
xnor U35782 (N_35782,N_33977,N_34317);
nand U35783 (N_35783,N_33297,N_33782);
nand U35784 (N_35784,N_33134,N_34926);
or U35785 (N_35785,N_33300,N_33506);
nor U35786 (N_35786,N_34226,N_32747);
or U35787 (N_35787,N_33591,N_34966);
xor U35788 (N_35788,N_32711,N_34675);
nor U35789 (N_35789,N_33192,N_33416);
xor U35790 (N_35790,N_33266,N_33015);
and U35791 (N_35791,N_34838,N_34204);
nand U35792 (N_35792,N_32978,N_34971);
xnor U35793 (N_35793,N_33705,N_33073);
nand U35794 (N_35794,N_32863,N_34487);
and U35795 (N_35795,N_32974,N_33209);
nor U35796 (N_35796,N_34069,N_34373);
or U35797 (N_35797,N_33740,N_32950);
and U35798 (N_35798,N_34551,N_34927);
nor U35799 (N_35799,N_34255,N_34398);
nand U35800 (N_35800,N_34019,N_34414);
nand U35801 (N_35801,N_33239,N_32698);
xnor U35802 (N_35802,N_34249,N_34018);
or U35803 (N_35803,N_33642,N_34909);
xor U35804 (N_35804,N_32884,N_32732);
nor U35805 (N_35805,N_34587,N_33336);
nand U35806 (N_35806,N_34590,N_32730);
nor U35807 (N_35807,N_33212,N_34508);
nand U35808 (N_35808,N_32690,N_32838);
or U35809 (N_35809,N_34907,N_34666);
or U35810 (N_35810,N_33352,N_34228);
and U35811 (N_35811,N_34372,N_34985);
nor U35812 (N_35812,N_33869,N_34314);
or U35813 (N_35813,N_34047,N_32942);
nand U35814 (N_35814,N_33148,N_34656);
nor U35815 (N_35815,N_32774,N_34532);
nand U35816 (N_35816,N_33760,N_33077);
nand U35817 (N_35817,N_32763,N_33811);
and U35818 (N_35818,N_34063,N_32552);
or U35819 (N_35819,N_34062,N_33263);
nand U35820 (N_35820,N_34483,N_34640);
nor U35821 (N_35821,N_34581,N_34760);
or U35822 (N_35822,N_32567,N_33986);
or U35823 (N_35823,N_33003,N_33950);
nand U35824 (N_35824,N_33345,N_33780);
xnor U35825 (N_35825,N_32820,N_34133);
or U35826 (N_35826,N_33094,N_34687);
nand U35827 (N_35827,N_32636,N_33821);
and U35828 (N_35828,N_33220,N_33423);
and U35829 (N_35829,N_34386,N_33010);
and U35830 (N_35830,N_34256,N_34128);
xor U35831 (N_35831,N_34058,N_34388);
and U35832 (N_35832,N_33279,N_33762);
and U35833 (N_35833,N_33100,N_34730);
nor U35834 (N_35834,N_33057,N_33928);
and U35835 (N_35835,N_32624,N_33976);
nand U35836 (N_35836,N_32930,N_34977);
or U35837 (N_35837,N_34042,N_34757);
xor U35838 (N_35838,N_32833,N_34602);
and U35839 (N_35839,N_32990,N_33342);
or U35840 (N_35840,N_32576,N_33166);
nor U35841 (N_35841,N_34328,N_34169);
nor U35842 (N_35842,N_34633,N_32517);
and U35843 (N_35843,N_34324,N_33458);
and U35844 (N_35844,N_32903,N_32505);
nand U35845 (N_35845,N_32883,N_34492);
or U35846 (N_35846,N_33544,N_34076);
nand U35847 (N_35847,N_33652,N_33546);
xnor U35848 (N_35848,N_34144,N_33191);
xnor U35849 (N_35849,N_34881,N_34468);
nand U35850 (N_35850,N_34901,N_32993);
or U35851 (N_35851,N_33098,N_33413);
xor U35852 (N_35852,N_33443,N_34402);
nand U35853 (N_35853,N_34664,N_33296);
xor U35854 (N_35854,N_34653,N_33741);
nor U35855 (N_35855,N_33475,N_34127);
nor U35856 (N_35856,N_33387,N_34734);
and U35857 (N_35857,N_32956,N_34369);
xnor U35858 (N_35858,N_33550,N_34341);
and U35859 (N_35859,N_32578,N_34416);
nor U35860 (N_35860,N_34449,N_34738);
nand U35861 (N_35861,N_33316,N_34280);
nor U35862 (N_35862,N_33195,N_33235);
nor U35863 (N_35863,N_34453,N_32895);
nor U35864 (N_35864,N_34616,N_33910);
or U35865 (N_35865,N_34198,N_34548);
nand U35866 (N_35866,N_34967,N_33198);
nor U35867 (N_35867,N_32963,N_34870);
or U35868 (N_35868,N_32708,N_33820);
nor U35869 (N_35869,N_33672,N_34306);
nor U35870 (N_35870,N_34037,N_33664);
nand U35871 (N_35871,N_34917,N_34321);
nor U35872 (N_35872,N_32714,N_34281);
and U35873 (N_35873,N_33370,N_33337);
nor U35874 (N_35874,N_34435,N_32502);
nor U35875 (N_35875,N_33494,N_34049);
nor U35876 (N_35876,N_33759,N_33614);
xor U35877 (N_35877,N_34025,N_34643);
or U35878 (N_35878,N_34106,N_33624);
and U35879 (N_35879,N_34546,N_32921);
xor U35880 (N_35880,N_34608,N_34953);
nor U35881 (N_35881,N_34798,N_34203);
xnor U35882 (N_35882,N_33982,N_32918);
and U35883 (N_35883,N_34875,N_34043);
nand U35884 (N_35884,N_33952,N_33814);
nand U35885 (N_35885,N_33033,N_32916);
xor U35886 (N_35886,N_33043,N_33381);
xor U35887 (N_35887,N_32939,N_34518);
xor U35888 (N_35888,N_34549,N_33989);
or U35889 (N_35889,N_34379,N_34294);
nor U35890 (N_35890,N_32522,N_33722);
xnor U35891 (N_35891,N_33940,N_33993);
or U35892 (N_35892,N_32722,N_34269);
and U35893 (N_35893,N_34578,N_32681);
xnor U35894 (N_35894,N_32910,N_33503);
nor U35895 (N_35895,N_33919,N_33318);
or U35896 (N_35896,N_33991,N_34553);
or U35897 (N_35897,N_34774,N_34795);
and U35898 (N_35898,N_33679,N_32768);
xor U35899 (N_35899,N_33476,N_34393);
nand U35900 (N_35900,N_33621,N_32835);
and U35901 (N_35901,N_34064,N_33072);
xor U35902 (N_35902,N_33518,N_33553);
and U35903 (N_35903,N_33471,N_34580);
and U35904 (N_35904,N_34874,N_34625);
nor U35905 (N_35905,N_33859,N_33012);
nor U35906 (N_35906,N_34116,N_34174);
and U35907 (N_35907,N_33047,N_32864);
nor U35908 (N_35908,N_32924,N_34912);
and U35909 (N_35909,N_32545,N_33162);
or U35910 (N_35910,N_34769,N_32524);
xnor U35911 (N_35911,N_33929,N_33570);
xnor U35912 (N_35912,N_34023,N_33097);
xnor U35913 (N_35913,N_34842,N_33161);
or U35914 (N_35914,N_32523,N_34949);
and U35915 (N_35915,N_34944,N_32972);
xor U35916 (N_35916,N_32736,N_33680);
nand U35917 (N_35917,N_34257,N_33893);
xor U35918 (N_35918,N_34343,N_34434);
xor U35919 (N_35919,N_33551,N_34513);
nand U35920 (N_35920,N_33459,N_34045);
and U35921 (N_35921,N_32541,N_32729);
and U35922 (N_35922,N_33936,N_32927);
xnor U35923 (N_35923,N_33350,N_34441);
and U35924 (N_35924,N_33099,N_34661);
or U35925 (N_35925,N_33382,N_34087);
or U35926 (N_35926,N_33963,N_34105);
or U35927 (N_35927,N_34793,N_32966);
and U35928 (N_35928,N_34500,N_34234);
and U35929 (N_35929,N_33786,N_32515);
and U35930 (N_35930,N_34327,N_32547);
nor U35931 (N_35931,N_34159,N_32758);
nor U35932 (N_35932,N_33867,N_34190);
or U35933 (N_35933,N_33549,N_32676);
nand U35934 (N_35934,N_34570,N_34445);
xnor U35935 (N_35935,N_33412,N_33917);
or U35936 (N_35936,N_33320,N_32689);
nor U35937 (N_35937,N_34450,N_32651);
xnor U35938 (N_35938,N_33635,N_34863);
or U35939 (N_35939,N_34700,N_34522);
nand U35940 (N_35940,N_33695,N_32507);
and U35941 (N_35941,N_34354,N_34684);
nor U35942 (N_35942,N_34695,N_33717);
and U35943 (N_35943,N_32992,N_34655);
nand U35944 (N_35944,N_33763,N_33454);
or U35945 (N_35945,N_33298,N_33265);
or U35946 (N_35946,N_34210,N_34154);
and U35947 (N_35947,N_34485,N_32533);
nand U35948 (N_35948,N_32525,N_33863);
nor U35949 (N_35949,N_33301,N_33486);
nand U35950 (N_35950,N_33225,N_33754);
nand U35951 (N_35951,N_34596,N_34263);
xnor U35952 (N_35952,N_34044,N_33448);
and U35953 (N_35953,N_34347,N_33089);
or U35954 (N_35954,N_34571,N_33886);
xor U35955 (N_35955,N_33582,N_33960);
and U35956 (N_35956,N_33688,N_34054);
nand U35957 (N_35957,N_33250,N_33037);
nor U35958 (N_35958,N_32821,N_33832);
nand U35959 (N_35959,N_33445,N_34560);
nor U35960 (N_35960,N_34568,N_33733);
nand U35961 (N_35961,N_34836,N_34579);
nand U35962 (N_35962,N_34172,N_32946);
and U35963 (N_35963,N_34668,N_32984);
or U35964 (N_35964,N_32760,N_33647);
nor U35965 (N_35965,N_32795,N_32668);
nand U35966 (N_35966,N_33779,N_34753);
and U35967 (N_35967,N_34430,N_34247);
nand U35968 (N_35968,N_32945,N_34725);
and U35969 (N_35969,N_34200,N_32962);
or U35970 (N_35970,N_34742,N_34923);
xor U35971 (N_35971,N_33587,N_33714);
nor U35972 (N_35972,N_32905,N_34910);
and U35973 (N_35973,N_34857,N_34755);
and U35974 (N_35974,N_33470,N_33547);
nor U35975 (N_35975,N_34781,N_34448);
and U35976 (N_35976,N_33441,N_32958);
or U35977 (N_35977,N_34472,N_33127);
xnor U35978 (N_35978,N_33934,N_34905);
or U35979 (N_35979,N_33444,N_34080);
xor U35980 (N_35980,N_34078,N_33922);
nand U35981 (N_35981,N_34497,N_33276);
or U35982 (N_35982,N_34538,N_34662);
or U35983 (N_35983,N_33325,N_33085);
xor U35984 (N_35984,N_34559,N_34762);
nor U35985 (N_35985,N_34832,N_34205);
nor U35986 (N_35986,N_34160,N_32652);
and U35987 (N_35987,N_34436,N_33139);
or U35988 (N_35988,N_34016,N_33829);
or U35989 (N_35989,N_33713,N_32584);
nand U35990 (N_35990,N_34014,N_33478);
nor U35991 (N_35991,N_32791,N_32979);
and U35992 (N_35992,N_34410,N_33777);
nor U35993 (N_35993,N_33376,N_32759);
nand U35994 (N_35994,N_34527,N_33951);
nor U35995 (N_35995,N_32680,N_32859);
xnor U35996 (N_35996,N_33803,N_33699);
nand U35997 (N_35997,N_33483,N_34807);
and U35998 (N_35998,N_33433,N_34605);
xor U35999 (N_35999,N_33539,N_34698);
nand U36000 (N_36000,N_34139,N_34467);
xnor U36001 (N_36001,N_33633,N_34006);
nand U36002 (N_36002,N_32862,N_33145);
or U36003 (N_36003,N_32527,N_34333);
xnor U36004 (N_36004,N_32562,N_33855);
or U36005 (N_36005,N_34822,N_34475);
xnor U36006 (N_36006,N_34358,N_32788);
xnor U36007 (N_36007,N_33451,N_34235);
and U36008 (N_36008,N_34520,N_33208);
or U36009 (N_36009,N_33612,N_33944);
and U36010 (N_36010,N_34053,N_33906);
and U36011 (N_36011,N_32948,N_33034);
or U36012 (N_36012,N_33013,N_33595);
nor U36013 (N_36013,N_33573,N_32743);
nand U36014 (N_36014,N_33373,N_33843);
or U36015 (N_36015,N_32928,N_33424);
nor U36016 (N_36016,N_34371,N_33083);
nor U36017 (N_36017,N_34057,N_34620);
or U36018 (N_36018,N_34275,N_34929);
xnor U36019 (N_36019,N_34524,N_34652);
and U36020 (N_36020,N_33604,N_32829);
nand U36021 (N_36021,N_34677,N_33087);
nor U36022 (N_36022,N_34533,N_34840);
or U36023 (N_36023,N_34539,N_33130);
xnor U36024 (N_36024,N_32531,N_33415);
nor U36025 (N_36025,N_34482,N_34644);
nand U36026 (N_36026,N_33562,N_33696);
nor U36027 (N_36027,N_33531,N_32855);
or U36028 (N_36028,N_33528,N_33407);
nor U36029 (N_36029,N_34638,N_33668);
nand U36030 (N_36030,N_33469,N_33702);
or U36031 (N_36031,N_34179,N_32804);
nand U36032 (N_36032,N_32700,N_34767);
nor U36033 (N_36033,N_33378,N_34614);
xor U36034 (N_36034,N_34201,N_34598);
xnor U36035 (N_36035,N_32857,N_34601);
xor U36036 (N_36036,N_32823,N_34229);
nand U36037 (N_36037,N_33359,N_33194);
or U36038 (N_36038,N_34446,N_33002);
xor U36039 (N_36039,N_33066,N_33275);
or U36040 (N_36040,N_32564,N_33954);
or U36041 (N_36041,N_33767,N_34886);
nor U36042 (N_36042,N_33084,N_34883);
nand U36043 (N_36043,N_34253,N_32654);
nand U36044 (N_36044,N_34686,N_34785);
or U36045 (N_36045,N_33876,N_33149);
or U36046 (N_36046,N_33938,N_32887);
nor U36047 (N_36047,N_34904,N_32617);
nor U36048 (N_36048,N_34300,N_33937);
and U36049 (N_36049,N_32751,N_33088);
nor U36050 (N_36050,N_34908,N_34930);
or U36051 (N_36051,N_34940,N_34958);
nor U36052 (N_36052,N_34496,N_33281);
nand U36053 (N_36053,N_33650,N_32803);
or U36054 (N_36054,N_33639,N_33816);
xnor U36055 (N_36055,N_34060,N_33916);
nor U36056 (N_36056,N_33513,N_33223);
nand U36057 (N_36057,N_33813,N_33050);
or U36058 (N_36058,N_33490,N_33725);
and U36059 (N_36059,N_34516,N_34243);
nand U36060 (N_36060,N_34720,N_33719);
or U36061 (N_36061,N_34924,N_32693);
or U36062 (N_36062,N_32894,N_33885);
and U36063 (N_36063,N_34585,N_32976);
and U36064 (N_36064,N_32709,N_32920);
xnor U36065 (N_36065,N_33482,N_34962);
nor U36066 (N_36066,N_34871,N_33723);
nor U36067 (N_36067,N_32923,N_34701);
or U36068 (N_36068,N_33967,N_32757);
nor U36069 (N_36069,N_32694,N_34384);
or U36070 (N_36070,N_34599,N_34987);
nand U36071 (N_36071,N_34196,N_34828);
and U36072 (N_36072,N_34469,N_33248);
xnor U36073 (N_36073,N_33534,N_32618);
nor U36074 (N_36074,N_34164,N_33333);
xnor U36075 (N_36075,N_34647,N_33507);
nand U36076 (N_36076,N_33391,N_32641);
nand U36077 (N_36077,N_33975,N_33141);
nand U36078 (N_36078,N_32726,N_33163);
or U36079 (N_36079,N_34976,N_32865);
and U36080 (N_36080,N_34876,N_32638);
nor U36081 (N_36081,N_32765,N_33355);
nand U36082 (N_36082,N_34180,N_34244);
nand U36083 (N_36083,N_32727,N_34813);
xor U36084 (N_36084,N_33520,N_32511);
and U36085 (N_36085,N_33174,N_32766);
or U36086 (N_36086,N_34645,N_33864);
or U36087 (N_36087,N_34326,N_34104);
nand U36088 (N_36088,N_33512,N_32906);
or U36089 (N_36089,N_33913,N_33848);
and U36090 (N_36090,N_34995,N_34029);
nor U36091 (N_36091,N_32801,N_32508);
xor U36092 (N_36092,N_34454,N_33151);
nand U36093 (N_36093,N_33887,N_34011);
or U36094 (N_36094,N_33529,N_34166);
xnor U36095 (N_36095,N_34821,N_32741);
xnor U36096 (N_36096,N_33838,N_33605);
xor U36097 (N_36097,N_34784,N_34165);
xor U36098 (N_36098,N_34514,N_33898);
nor U36099 (N_36099,N_33594,N_34517);
or U36100 (N_36100,N_33965,N_32922);
and U36101 (N_36101,N_34320,N_33167);
xnor U36102 (N_36102,N_34797,N_32873);
nand U36103 (N_36103,N_33159,N_33110);
or U36104 (N_36104,N_33108,N_34361);
nor U36105 (N_36105,N_32975,N_33128);
xor U36106 (N_36106,N_33255,N_34153);
or U36107 (N_36107,N_33675,N_32597);
xnor U36108 (N_36108,N_34564,N_33121);
nand U36109 (N_36109,N_33045,N_33998);
xnor U36110 (N_36110,N_33406,N_34635);
and U36111 (N_36111,N_34152,N_32837);
nand U36112 (N_36112,N_33485,N_33819);
and U36113 (N_36113,N_34498,N_32635);
nor U36114 (N_36114,N_33530,N_34421);
and U36115 (N_36115,N_34866,N_34678);
nor U36116 (N_36116,N_34740,N_33244);
xnor U36117 (N_36117,N_32893,N_34387);
and U36118 (N_36118,N_34844,N_33941);
nor U36119 (N_36119,N_34859,N_32852);
or U36120 (N_36120,N_32556,N_34504);
nor U36121 (N_36121,N_33405,N_34195);
nor U36122 (N_36122,N_34808,N_33870);
or U36123 (N_36123,N_34708,N_34286);
nor U36124 (N_36124,N_32996,N_34470);
nand U36125 (N_36125,N_33628,N_32603);
and U36126 (N_36126,N_33560,N_32843);
or U36127 (N_36127,N_33418,N_34481);
xor U36128 (N_36128,N_34892,N_32814);
and U36129 (N_36129,N_34206,N_34897);
nor U36130 (N_36130,N_33873,N_32810);
or U36131 (N_36131,N_34884,N_33815);
nor U36132 (N_36132,N_33075,N_33282);
nand U36133 (N_36133,N_33924,N_34594);
nor U36134 (N_36134,N_34178,N_32762);
nand U36135 (N_36135,N_33511,N_32665);
xor U36136 (N_36136,N_33335,N_34986);
or U36137 (N_36137,N_33921,N_33170);
nand U36138 (N_36138,N_32856,N_34143);
xnor U36139 (N_36139,N_32944,N_33389);
or U36140 (N_36140,N_34685,N_33101);
or U36141 (N_36141,N_34920,N_32982);
nor U36142 (N_36142,N_33176,N_34349);
nand U36143 (N_36143,N_32748,N_33860);
and U36144 (N_36144,N_34893,N_34545);
xnor U36145 (N_36145,N_34092,N_33215);
nor U36146 (N_36146,N_33290,N_33566);
and U36147 (N_36147,N_34931,N_32648);
xnor U36148 (N_36148,N_33737,N_34658);
nor U36149 (N_36149,N_33992,N_32512);
xnor U36150 (N_36150,N_34313,N_33712);
xnor U36151 (N_36151,N_33769,N_34494);
nor U36152 (N_36152,N_33726,N_32626);
and U36153 (N_36153,N_33527,N_33498);
or U36154 (N_36154,N_34704,N_34336);
nor U36155 (N_36155,N_33368,N_33082);
nor U36156 (N_36156,N_34221,N_34683);
nand U36157 (N_36157,N_34248,N_32845);
and U36158 (N_36158,N_34600,N_33833);
xor U36159 (N_36159,N_34577,N_33555);
nor U36160 (N_36160,N_34933,N_33338);
xnor U36161 (N_36161,N_33160,N_33793);
nand U36162 (N_36162,N_32969,N_33306);
or U36163 (N_36163,N_32569,N_34827);
nor U36164 (N_36164,N_34208,N_33206);
and U36165 (N_36165,N_33615,N_33204);
nor U36166 (N_36166,N_32901,N_34145);
and U36167 (N_36167,N_34380,N_33440);
nand U36168 (N_36168,N_34158,N_34217);
and U36169 (N_36169,N_33939,N_32520);
nor U36170 (N_36170,N_33574,N_33781);
and U36171 (N_36171,N_33764,N_34819);
or U36172 (N_36172,N_34113,N_34707);
nor U36173 (N_36173,N_32521,N_34543);
and U36174 (N_36174,N_34823,N_32701);
nor U36175 (N_36175,N_32599,N_32847);
xor U36176 (N_36176,N_32866,N_32639);
xor U36177 (N_36177,N_34657,N_33138);
or U36178 (N_36178,N_33548,N_34665);
nand U36179 (N_36179,N_34378,N_33096);
and U36180 (N_36180,N_32919,N_33558);
xnor U36181 (N_36181,N_32589,N_34177);
or U36182 (N_36182,N_33165,N_32667);
nor U36183 (N_36183,N_34817,N_34473);
nand U36184 (N_36184,N_33484,N_33409);
nand U36185 (N_36185,N_32998,N_33004);
nand U36186 (N_36186,N_34181,N_34465);
or U36187 (N_36187,N_32634,N_33488);
xor U36188 (N_36188,N_34878,N_34951);
nor U36189 (N_36189,N_32951,N_34773);
and U36190 (N_36190,N_34474,N_32849);
xor U36191 (N_36191,N_33958,N_34959);
and U36192 (N_36192,N_34039,N_34329);
nor U36193 (N_36193,N_34770,N_33142);
and U36194 (N_36194,N_33882,N_33542);
xor U36195 (N_36195,N_32745,N_33175);
xnor U36196 (N_36196,N_34090,N_33125);
or U36197 (N_36197,N_34034,N_33957);
nor U36198 (N_36198,N_33453,N_34942);
or U36199 (N_36199,N_33802,N_33678);
nand U36200 (N_36200,N_34583,N_32938);
and U36201 (N_36201,N_32780,N_33049);
xnor U36202 (N_36202,N_34736,N_34982);
nor U36203 (N_36203,N_32687,N_32612);
nor U36204 (N_36204,N_32914,N_33219);
nor U36205 (N_36205,N_34185,N_33810);
nand U36206 (N_36206,N_34764,N_33602);
nand U36207 (N_36207,N_34026,N_33613);
xor U36208 (N_36208,N_32955,N_34216);
nand U36209 (N_36209,N_33051,N_33293);
xnor U36210 (N_36210,N_33945,N_34727);
nor U36211 (N_36211,N_33535,N_33258);
nand U36212 (N_36212,N_32973,N_34814);
xor U36213 (N_36213,N_32850,N_34415);
and U36214 (N_36214,N_34903,N_34331);
nand U36215 (N_36215,N_32999,N_34792);
nand U36216 (N_36216,N_33230,N_34721);
and U36217 (N_36217,N_33804,N_33109);
and U36218 (N_36218,N_34804,N_33665);
or U36219 (N_36219,N_34789,N_32949);
and U36220 (N_36220,N_33610,N_34670);
nand U36221 (N_36221,N_34537,N_32650);
or U36222 (N_36222,N_32677,N_34756);
xnor U36223 (N_36223,N_34495,N_33207);
nor U36224 (N_36224,N_34607,N_34102);
and U36225 (N_36225,N_33830,N_34562);
nor U36226 (N_36226,N_32917,N_34921);
or U36227 (N_36227,N_34330,N_33171);
and U36228 (N_36228,N_34928,N_32826);
xnor U36229 (N_36229,N_33112,N_33314);
or U36230 (N_36230,N_34005,N_34825);
nand U36231 (N_36231,N_34835,N_32934);
xor U36232 (N_36232,N_33775,N_34950);
xnor U36233 (N_36233,N_32705,N_33402);
and U36234 (N_36234,N_34311,N_33994);
and U36235 (N_36235,N_33932,N_32908);
or U36236 (N_36236,N_34697,N_33568);
nor U36237 (N_36237,N_32960,N_34932);
xor U36238 (N_36238,N_33883,N_34110);
nor U36239 (N_36239,N_34511,N_33334);
or U36240 (N_36240,N_32947,N_32551);
and U36241 (N_36241,N_33842,N_34689);
nor U36242 (N_36242,N_34963,N_33817);
nand U36243 (N_36243,N_32878,N_33738);
xor U36244 (N_36244,N_33834,N_33554);
or U36245 (N_36245,N_33926,N_34010);
xor U36246 (N_36246,N_34334,N_34186);
xor U36247 (N_36247,N_34557,N_32805);
xnor U36248 (N_36248,N_33131,N_34251);
nor U36249 (N_36249,N_34258,N_34346);
nor U36250 (N_36250,N_33294,N_33571);
and U36251 (N_36251,N_33172,N_34433);
xor U36252 (N_36252,N_33685,N_32608);
or U36253 (N_36253,N_33478,N_32948);
and U36254 (N_36254,N_34267,N_32831);
xor U36255 (N_36255,N_33370,N_34241);
nor U36256 (N_36256,N_32666,N_33016);
or U36257 (N_36257,N_34298,N_33851);
nor U36258 (N_36258,N_32847,N_33573);
or U36259 (N_36259,N_34704,N_34416);
nor U36260 (N_36260,N_34221,N_33846);
or U36261 (N_36261,N_33450,N_34510);
and U36262 (N_36262,N_34598,N_32833);
xnor U36263 (N_36263,N_33057,N_34373);
or U36264 (N_36264,N_34200,N_33078);
or U36265 (N_36265,N_32704,N_34557);
or U36266 (N_36266,N_32877,N_33241);
and U36267 (N_36267,N_33586,N_34766);
nor U36268 (N_36268,N_33924,N_33351);
nand U36269 (N_36269,N_34497,N_32917);
nor U36270 (N_36270,N_32702,N_34239);
or U36271 (N_36271,N_34818,N_33445);
and U36272 (N_36272,N_34451,N_34763);
nand U36273 (N_36273,N_34102,N_32884);
xnor U36274 (N_36274,N_34553,N_34481);
nand U36275 (N_36275,N_32639,N_33244);
nor U36276 (N_36276,N_33217,N_34162);
nand U36277 (N_36277,N_32846,N_33893);
nand U36278 (N_36278,N_32861,N_33909);
and U36279 (N_36279,N_32858,N_33951);
nand U36280 (N_36280,N_32503,N_32667);
nand U36281 (N_36281,N_33703,N_34819);
nor U36282 (N_36282,N_33801,N_32726);
xnor U36283 (N_36283,N_34043,N_33752);
and U36284 (N_36284,N_34259,N_34319);
xnor U36285 (N_36285,N_32619,N_34057);
xor U36286 (N_36286,N_32909,N_34155);
nand U36287 (N_36287,N_34310,N_34002);
nor U36288 (N_36288,N_33792,N_33257);
xnor U36289 (N_36289,N_33681,N_34113);
or U36290 (N_36290,N_32728,N_32667);
or U36291 (N_36291,N_32831,N_32658);
and U36292 (N_36292,N_33248,N_33261);
xnor U36293 (N_36293,N_33849,N_33942);
or U36294 (N_36294,N_34927,N_34958);
nand U36295 (N_36295,N_32902,N_33600);
nor U36296 (N_36296,N_34579,N_33965);
nor U36297 (N_36297,N_32717,N_34917);
nand U36298 (N_36298,N_33903,N_34376);
xnor U36299 (N_36299,N_33752,N_34072);
nor U36300 (N_36300,N_32616,N_33238);
and U36301 (N_36301,N_34189,N_33770);
or U36302 (N_36302,N_32929,N_34036);
and U36303 (N_36303,N_34359,N_34144);
or U36304 (N_36304,N_32618,N_34927);
nand U36305 (N_36305,N_32699,N_33111);
xnor U36306 (N_36306,N_34669,N_32797);
nand U36307 (N_36307,N_34373,N_34280);
or U36308 (N_36308,N_33801,N_32968);
and U36309 (N_36309,N_34931,N_33921);
nand U36310 (N_36310,N_32868,N_32984);
and U36311 (N_36311,N_33655,N_33700);
and U36312 (N_36312,N_33479,N_34653);
nand U36313 (N_36313,N_34685,N_33056);
xor U36314 (N_36314,N_34108,N_34708);
nand U36315 (N_36315,N_32937,N_33700);
and U36316 (N_36316,N_32947,N_33129);
or U36317 (N_36317,N_34663,N_33420);
or U36318 (N_36318,N_33273,N_33007);
nor U36319 (N_36319,N_34595,N_34007);
nand U36320 (N_36320,N_34420,N_32690);
xor U36321 (N_36321,N_32962,N_34384);
or U36322 (N_36322,N_34757,N_34507);
nor U36323 (N_36323,N_32978,N_34849);
nand U36324 (N_36324,N_34678,N_34816);
nand U36325 (N_36325,N_34758,N_34183);
and U36326 (N_36326,N_33847,N_33623);
and U36327 (N_36327,N_34227,N_34932);
xor U36328 (N_36328,N_34745,N_34205);
or U36329 (N_36329,N_32609,N_34974);
and U36330 (N_36330,N_33444,N_32991);
or U36331 (N_36331,N_34537,N_32873);
xor U36332 (N_36332,N_34287,N_33740);
and U36333 (N_36333,N_34212,N_32811);
nand U36334 (N_36334,N_33822,N_32834);
or U36335 (N_36335,N_32815,N_33081);
nand U36336 (N_36336,N_34518,N_32687);
nand U36337 (N_36337,N_32874,N_32611);
or U36338 (N_36338,N_34271,N_34619);
xor U36339 (N_36339,N_32554,N_34071);
and U36340 (N_36340,N_33596,N_34984);
xnor U36341 (N_36341,N_34483,N_34611);
nand U36342 (N_36342,N_34905,N_34390);
xor U36343 (N_36343,N_34541,N_34507);
xor U36344 (N_36344,N_34477,N_34751);
or U36345 (N_36345,N_32807,N_33952);
xnor U36346 (N_36346,N_33974,N_34482);
and U36347 (N_36347,N_32847,N_33328);
nand U36348 (N_36348,N_32626,N_33989);
nand U36349 (N_36349,N_32716,N_33138);
or U36350 (N_36350,N_33652,N_33136);
and U36351 (N_36351,N_33196,N_34762);
nand U36352 (N_36352,N_33688,N_32540);
nand U36353 (N_36353,N_34533,N_34087);
nor U36354 (N_36354,N_32840,N_34406);
xor U36355 (N_36355,N_34407,N_33524);
nor U36356 (N_36356,N_33367,N_33601);
nor U36357 (N_36357,N_33462,N_32654);
or U36358 (N_36358,N_33928,N_33886);
or U36359 (N_36359,N_34792,N_33022);
xnor U36360 (N_36360,N_34478,N_33848);
and U36361 (N_36361,N_32797,N_34002);
or U36362 (N_36362,N_33324,N_33467);
or U36363 (N_36363,N_34440,N_34179);
nand U36364 (N_36364,N_34906,N_33021);
and U36365 (N_36365,N_32580,N_33017);
nand U36366 (N_36366,N_34617,N_33944);
or U36367 (N_36367,N_32500,N_34519);
or U36368 (N_36368,N_32917,N_34990);
or U36369 (N_36369,N_34433,N_33728);
or U36370 (N_36370,N_32504,N_33789);
nor U36371 (N_36371,N_33070,N_33740);
and U36372 (N_36372,N_32945,N_34506);
and U36373 (N_36373,N_34147,N_33787);
nor U36374 (N_36374,N_32813,N_34502);
and U36375 (N_36375,N_32981,N_33780);
and U36376 (N_36376,N_34212,N_33679);
or U36377 (N_36377,N_33469,N_34518);
xor U36378 (N_36378,N_34660,N_34161);
nor U36379 (N_36379,N_34130,N_32861);
nor U36380 (N_36380,N_33349,N_33558);
and U36381 (N_36381,N_33882,N_33597);
nor U36382 (N_36382,N_34694,N_32987);
and U36383 (N_36383,N_33157,N_34585);
and U36384 (N_36384,N_34836,N_33622);
xnor U36385 (N_36385,N_32923,N_34562);
nand U36386 (N_36386,N_33824,N_34602);
or U36387 (N_36387,N_32697,N_34357);
nor U36388 (N_36388,N_34142,N_34838);
xnor U36389 (N_36389,N_34368,N_32955);
and U36390 (N_36390,N_34121,N_33314);
xnor U36391 (N_36391,N_33891,N_34550);
nor U36392 (N_36392,N_33473,N_33166);
xnor U36393 (N_36393,N_33667,N_34996);
or U36394 (N_36394,N_33940,N_33138);
or U36395 (N_36395,N_32888,N_34844);
or U36396 (N_36396,N_34219,N_32852);
or U36397 (N_36397,N_33786,N_33806);
xnor U36398 (N_36398,N_32775,N_34460);
or U36399 (N_36399,N_34113,N_33464);
and U36400 (N_36400,N_34185,N_34114);
xnor U36401 (N_36401,N_33588,N_34649);
nand U36402 (N_36402,N_33491,N_33144);
or U36403 (N_36403,N_33839,N_34723);
and U36404 (N_36404,N_34993,N_34968);
and U36405 (N_36405,N_32972,N_34734);
or U36406 (N_36406,N_34634,N_32924);
nor U36407 (N_36407,N_32994,N_32847);
nand U36408 (N_36408,N_34234,N_34900);
nand U36409 (N_36409,N_33667,N_32523);
and U36410 (N_36410,N_33884,N_32950);
nor U36411 (N_36411,N_33001,N_33245);
xor U36412 (N_36412,N_34879,N_33493);
or U36413 (N_36413,N_34817,N_34930);
xor U36414 (N_36414,N_33227,N_33542);
or U36415 (N_36415,N_33732,N_32946);
nor U36416 (N_36416,N_33128,N_34643);
nor U36417 (N_36417,N_33774,N_34741);
and U36418 (N_36418,N_34619,N_33061);
nor U36419 (N_36419,N_34138,N_34345);
and U36420 (N_36420,N_34734,N_32934);
xnor U36421 (N_36421,N_33811,N_34910);
and U36422 (N_36422,N_33242,N_33454);
nand U36423 (N_36423,N_32909,N_34061);
nand U36424 (N_36424,N_32623,N_32536);
or U36425 (N_36425,N_33155,N_34206);
nor U36426 (N_36426,N_33924,N_34203);
and U36427 (N_36427,N_33324,N_33214);
or U36428 (N_36428,N_33282,N_34062);
and U36429 (N_36429,N_33653,N_34282);
nand U36430 (N_36430,N_32513,N_33826);
and U36431 (N_36431,N_34357,N_33192);
nand U36432 (N_36432,N_33978,N_34470);
nand U36433 (N_36433,N_32795,N_33432);
and U36434 (N_36434,N_33541,N_34657);
xor U36435 (N_36435,N_34971,N_33016);
or U36436 (N_36436,N_34029,N_34211);
nor U36437 (N_36437,N_32735,N_34876);
nor U36438 (N_36438,N_34579,N_33097);
or U36439 (N_36439,N_33403,N_32510);
or U36440 (N_36440,N_34866,N_33908);
and U36441 (N_36441,N_32537,N_33572);
nand U36442 (N_36442,N_33579,N_34685);
nand U36443 (N_36443,N_33552,N_33973);
or U36444 (N_36444,N_33588,N_34090);
and U36445 (N_36445,N_33312,N_34904);
nand U36446 (N_36446,N_34444,N_34343);
and U36447 (N_36447,N_32650,N_32846);
or U36448 (N_36448,N_34101,N_33489);
and U36449 (N_36449,N_33394,N_33016);
or U36450 (N_36450,N_34352,N_33729);
xnor U36451 (N_36451,N_34491,N_34897);
nor U36452 (N_36452,N_34320,N_33240);
nand U36453 (N_36453,N_34364,N_34960);
nand U36454 (N_36454,N_34036,N_33857);
and U36455 (N_36455,N_34718,N_33706);
and U36456 (N_36456,N_34255,N_33511);
nor U36457 (N_36457,N_34073,N_34027);
or U36458 (N_36458,N_33814,N_33108);
and U36459 (N_36459,N_32760,N_33134);
and U36460 (N_36460,N_34968,N_34130);
nand U36461 (N_36461,N_34090,N_32581);
and U36462 (N_36462,N_33474,N_33691);
nand U36463 (N_36463,N_34967,N_33987);
nor U36464 (N_36464,N_34894,N_33896);
and U36465 (N_36465,N_33114,N_34118);
nor U36466 (N_36466,N_33670,N_33700);
and U36467 (N_36467,N_34224,N_32891);
and U36468 (N_36468,N_33204,N_34382);
or U36469 (N_36469,N_32913,N_34112);
and U36470 (N_36470,N_33088,N_34753);
nor U36471 (N_36471,N_32921,N_33421);
and U36472 (N_36472,N_33605,N_33765);
nand U36473 (N_36473,N_34725,N_33622);
and U36474 (N_36474,N_33072,N_34088);
nand U36475 (N_36475,N_34956,N_33558);
and U36476 (N_36476,N_32586,N_32791);
xnor U36477 (N_36477,N_33599,N_32504);
and U36478 (N_36478,N_33375,N_33250);
nand U36479 (N_36479,N_33619,N_32704);
and U36480 (N_36480,N_32988,N_34760);
xor U36481 (N_36481,N_33380,N_33106);
or U36482 (N_36482,N_34958,N_33060);
xnor U36483 (N_36483,N_33142,N_34673);
nand U36484 (N_36484,N_33401,N_34815);
and U36485 (N_36485,N_33138,N_32955);
nand U36486 (N_36486,N_33469,N_33503);
nand U36487 (N_36487,N_34386,N_34379);
nand U36488 (N_36488,N_33346,N_33413);
nor U36489 (N_36489,N_32985,N_34973);
and U36490 (N_36490,N_34881,N_32538);
or U36491 (N_36491,N_33028,N_34023);
or U36492 (N_36492,N_34177,N_34594);
and U36493 (N_36493,N_33656,N_34772);
and U36494 (N_36494,N_33870,N_32519);
and U36495 (N_36495,N_32862,N_34645);
nor U36496 (N_36496,N_33421,N_33598);
or U36497 (N_36497,N_33596,N_32980);
nor U36498 (N_36498,N_34289,N_33982);
nand U36499 (N_36499,N_32920,N_34868);
or U36500 (N_36500,N_33604,N_34483);
or U36501 (N_36501,N_34694,N_33405);
and U36502 (N_36502,N_33763,N_32545);
xor U36503 (N_36503,N_33163,N_34838);
xnor U36504 (N_36504,N_32960,N_33546);
nand U36505 (N_36505,N_34994,N_34029);
nand U36506 (N_36506,N_32852,N_34598);
or U36507 (N_36507,N_32639,N_33973);
or U36508 (N_36508,N_33703,N_34246);
and U36509 (N_36509,N_33110,N_33436);
nand U36510 (N_36510,N_34779,N_34783);
nand U36511 (N_36511,N_34931,N_34754);
nand U36512 (N_36512,N_34182,N_34712);
and U36513 (N_36513,N_34913,N_33770);
nor U36514 (N_36514,N_33924,N_32585);
and U36515 (N_36515,N_33475,N_33693);
nand U36516 (N_36516,N_33769,N_34808);
and U36517 (N_36517,N_34428,N_32540);
or U36518 (N_36518,N_34009,N_32610);
or U36519 (N_36519,N_34353,N_32714);
nand U36520 (N_36520,N_33169,N_34078);
and U36521 (N_36521,N_34788,N_33630);
and U36522 (N_36522,N_32738,N_33334);
xor U36523 (N_36523,N_33791,N_33946);
or U36524 (N_36524,N_33164,N_33966);
nand U36525 (N_36525,N_33244,N_33007);
nor U36526 (N_36526,N_34595,N_34332);
and U36527 (N_36527,N_33771,N_33233);
nor U36528 (N_36528,N_34624,N_34472);
nor U36529 (N_36529,N_33981,N_33568);
or U36530 (N_36530,N_34616,N_33534);
and U36531 (N_36531,N_32747,N_32567);
and U36532 (N_36532,N_34232,N_33220);
nor U36533 (N_36533,N_33476,N_32854);
nand U36534 (N_36534,N_34110,N_34619);
or U36535 (N_36535,N_34740,N_33230);
or U36536 (N_36536,N_34650,N_33629);
xor U36537 (N_36537,N_33158,N_34144);
or U36538 (N_36538,N_32880,N_34914);
and U36539 (N_36539,N_34420,N_33523);
or U36540 (N_36540,N_34866,N_33590);
and U36541 (N_36541,N_33491,N_32969);
nand U36542 (N_36542,N_34286,N_33144);
nor U36543 (N_36543,N_33808,N_33290);
nor U36544 (N_36544,N_32992,N_34066);
and U36545 (N_36545,N_32896,N_34537);
nand U36546 (N_36546,N_34688,N_33276);
and U36547 (N_36547,N_33341,N_34955);
nor U36548 (N_36548,N_34242,N_34587);
nand U36549 (N_36549,N_33949,N_33494);
nand U36550 (N_36550,N_33513,N_33969);
nand U36551 (N_36551,N_33452,N_34124);
or U36552 (N_36552,N_34925,N_33711);
xor U36553 (N_36553,N_34903,N_34593);
and U36554 (N_36554,N_34903,N_32937);
and U36555 (N_36555,N_33762,N_34256);
xnor U36556 (N_36556,N_33113,N_34493);
nand U36557 (N_36557,N_33148,N_33815);
nand U36558 (N_36558,N_34914,N_34056);
and U36559 (N_36559,N_34700,N_32910);
or U36560 (N_36560,N_34807,N_34005);
nor U36561 (N_36561,N_33124,N_34281);
nand U36562 (N_36562,N_33543,N_33932);
nand U36563 (N_36563,N_34763,N_33947);
or U36564 (N_36564,N_33556,N_34015);
or U36565 (N_36565,N_34186,N_33855);
and U36566 (N_36566,N_33109,N_32628);
or U36567 (N_36567,N_34795,N_34369);
nor U36568 (N_36568,N_33127,N_33357);
or U36569 (N_36569,N_34473,N_34448);
nor U36570 (N_36570,N_34199,N_32746);
xor U36571 (N_36571,N_33139,N_33774);
xor U36572 (N_36572,N_34047,N_34728);
nor U36573 (N_36573,N_32540,N_33967);
nor U36574 (N_36574,N_34758,N_34419);
or U36575 (N_36575,N_33669,N_34034);
nand U36576 (N_36576,N_33600,N_34132);
and U36577 (N_36577,N_34602,N_33519);
xnor U36578 (N_36578,N_32501,N_33118);
nor U36579 (N_36579,N_33144,N_34873);
xor U36580 (N_36580,N_34869,N_32879);
xnor U36581 (N_36581,N_33644,N_34807);
nor U36582 (N_36582,N_33717,N_34721);
nor U36583 (N_36583,N_34807,N_33719);
nand U36584 (N_36584,N_34441,N_33091);
xor U36585 (N_36585,N_34802,N_33794);
nand U36586 (N_36586,N_33693,N_32597);
and U36587 (N_36587,N_34754,N_33508);
and U36588 (N_36588,N_33309,N_33901);
and U36589 (N_36589,N_33665,N_34748);
nor U36590 (N_36590,N_33071,N_34508);
xor U36591 (N_36591,N_34880,N_34045);
nor U36592 (N_36592,N_34453,N_32805);
nand U36593 (N_36593,N_33636,N_33052);
and U36594 (N_36594,N_32730,N_34291);
or U36595 (N_36595,N_34641,N_34247);
or U36596 (N_36596,N_34526,N_32677);
and U36597 (N_36597,N_34613,N_34523);
or U36598 (N_36598,N_34104,N_32879);
nand U36599 (N_36599,N_34508,N_34363);
nor U36600 (N_36600,N_34910,N_34272);
and U36601 (N_36601,N_33846,N_32622);
or U36602 (N_36602,N_33265,N_33224);
or U36603 (N_36603,N_34406,N_33100);
xnor U36604 (N_36604,N_33917,N_34275);
xor U36605 (N_36605,N_34611,N_33157);
xnor U36606 (N_36606,N_32668,N_33863);
nor U36607 (N_36607,N_34823,N_33067);
nand U36608 (N_36608,N_33780,N_33155);
and U36609 (N_36609,N_33931,N_33780);
nand U36610 (N_36610,N_34683,N_33928);
nor U36611 (N_36611,N_34372,N_34893);
nor U36612 (N_36612,N_33395,N_33414);
xor U36613 (N_36613,N_33579,N_34245);
and U36614 (N_36614,N_33315,N_34720);
xnor U36615 (N_36615,N_34727,N_33339);
and U36616 (N_36616,N_32697,N_33134);
nor U36617 (N_36617,N_33055,N_33277);
and U36618 (N_36618,N_32719,N_32816);
or U36619 (N_36619,N_34980,N_34260);
nand U36620 (N_36620,N_34455,N_34298);
and U36621 (N_36621,N_33193,N_33049);
or U36622 (N_36622,N_32979,N_33849);
and U36623 (N_36623,N_33586,N_33115);
and U36624 (N_36624,N_34572,N_33251);
nor U36625 (N_36625,N_32573,N_34837);
nor U36626 (N_36626,N_32527,N_33419);
xor U36627 (N_36627,N_33186,N_34081);
and U36628 (N_36628,N_32849,N_33839);
xnor U36629 (N_36629,N_34010,N_32597);
and U36630 (N_36630,N_34016,N_33823);
nor U36631 (N_36631,N_33512,N_33582);
and U36632 (N_36632,N_34373,N_34177);
or U36633 (N_36633,N_34555,N_34363);
or U36634 (N_36634,N_32995,N_32719);
xor U36635 (N_36635,N_34696,N_34211);
and U36636 (N_36636,N_33157,N_32866);
nor U36637 (N_36637,N_34796,N_34919);
nor U36638 (N_36638,N_34405,N_33002);
or U36639 (N_36639,N_33704,N_32802);
nor U36640 (N_36640,N_34587,N_33510);
nand U36641 (N_36641,N_33292,N_33661);
or U36642 (N_36642,N_34023,N_33351);
nor U36643 (N_36643,N_34382,N_34541);
nor U36644 (N_36644,N_34573,N_34672);
and U36645 (N_36645,N_34295,N_34428);
or U36646 (N_36646,N_33441,N_34394);
nor U36647 (N_36647,N_34288,N_33962);
nor U36648 (N_36648,N_33392,N_34410);
or U36649 (N_36649,N_32991,N_33590);
or U36650 (N_36650,N_32833,N_33774);
xnor U36651 (N_36651,N_34703,N_34154);
nand U36652 (N_36652,N_32585,N_33099);
nor U36653 (N_36653,N_34441,N_33288);
xor U36654 (N_36654,N_34678,N_34561);
and U36655 (N_36655,N_34787,N_34169);
nand U36656 (N_36656,N_34387,N_34646);
nor U36657 (N_36657,N_34787,N_34299);
nand U36658 (N_36658,N_32702,N_33840);
nor U36659 (N_36659,N_33906,N_34243);
and U36660 (N_36660,N_33112,N_32862);
and U36661 (N_36661,N_34967,N_33308);
xnor U36662 (N_36662,N_34904,N_32893);
xor U36663 (N_36663,N_34280,N_34627);
nor U36664 (N_36664,N_33755,N_33779);
nor U36665 (N_36665,N_34342,N_33576);
nor U36666 (N_36666,N_34539,N_34574);
nor U36667 (N_36667,N_34258,N_33573);
xnor U36668 (N_36668,N_32718,N_33395);
nor U36669 (N_36669,N_32735,N_33693);
xnor U36670 (N_36670,N_33705,N_34365);
nor U36671 (N_36671,N_32726,N_32613);
nand U36672 (N_36672,N_33708,N_32831);
or U36673 (N_36673,N_33969,N_33787);
or U36674 (N_36674,N_34025,N_32907);
or U36675 (N_36675,N_33279,N_34168);
and U36676 (N_36676,N_34343,N_33971);
and U36677 (N_36677,N_32777,N_34065);
and U36678 (N_36678,N_33418,N_33556);
xnor U36679 (N_36679,N_32970,N_33725);
and U36680 (N_36680,N_33923,N_32986);
xor U36681 (N_36681,N_34915,N_34393);
xnor U36682 (N_36682,N_33435,N_32729);
xor U36683 (N_36683,N_34407,N_33354);
nor U36684 (N_36684,N_33360,N_32834);
or U36685 (N_36685,N_33553,N_33471);
or U36686 (N_36686,N_33109,N_32778);
nor U36687 (N_36687,N_33047,N_33065);
and U36688 (N_36688,N_32531,N_32752);
nor U36689 (N_36689,N_32709,N_34577);
nor U36690 (N_36690,N_32579,N_33730);
nor U36691 (N_36691,N_33601,N_33278);
xnor U36692 (N_36692,N_34334,N_34572);
or U36693 (N_36693,N_32722,N_32911);
nand U36694 (N_36694,N_33659,N_33056);
and U36695 (N_36695,N_33569,N_34340);
nor U36696 (N_36696,N_34909,N_33391);
xnor U36697 (N_36697,N_34838,N_33279);
and U36698 (N_36698,N_33756,N_34269);
nor U36699 (N_36699,N_33070,N_33114);
nor U36700 (N_36700,N_33732,N_33517);
or U36701 (N_36701,N_34861,N_34138);
nor U36702 (N_36702,N_33023,N_34242);
nor U36703 (N_36703,N_34006,N_33454);
nor U36704 (N_36704,N_34040,N_34998);
xnor U36705 (N_36705,N_33680,N_32537);
or U36706 (N_36706,N_33443,N_33707);
xor U36707 (N_36707,N_34923,N_32749);
or U36708 (N_36708,N_33624,N_34987);
nand U36709 (N_36709,N_33901,N_33630);
xor U36710 (N_36710,N_33172,N_33283);
nand U36711 (N_36711,N_34458,N_32627);
nand U36712 (N_36712,N_33603,N_33520);
or U36713 (N_36713,N_34151,N_34908);
and U36714 (N_36714,N_33249,N_34677);
xnor U36715 (N_36715,N_32566,N_34301);
nor U36716 (N_36716,N_33497,N_32848);
nor U36717 (N_36717,N_33234,N_34084);
nor U36718 (N_36718,N_33059,N_33076);
and U36719 (N_36719,N_34060,N_34953);
and U36720 (N_36720,N_34933,N_34239);
or U36721 (N_36721,N_34578,N_33336);
or U36722 (N_36722,N_34786,N_33832);
nor U36723 (N_36723,N_33785,N_33249);
nand U36724 (N_36724,N_33049,N_34877);
or U36725 (N_36725,N_34339,N_34741);
or U36726 (N_36726,N_34523,N_33216);
xnor U36727 (N_36727,N_34751,N_33291);
or U36728 (N_36728,N_34055,N_33860);
xnor U36729 (N_36729,N_33971,N_34345);
nor U36730 (N_36730,N_34802,N_33002);
and U36731 (N_36731,N_33973,N_34565);
nor U36732 (N_36732,N_33707,N_34949);
nor U36733 (N_36733,N_33806,N_32688);
or U36734 (N_36734,N_33774,N_34064);
and U36735 (N_36735,N_34771,N_34749);
nor U36736 (N_36736,N_32706,N_34434);
and U36737 (N_36737,N_33290,N_34152);
nand U36738 (N_36738,N_34442,N_34137);
nand U36739 (N_36739,N_33259,N_33650);
nor U36740 (N_36740,N_34287,N_34364);
xor U36741 (N_36741,N_34503,N_34097);
xor U36742 (N_36742,N_34907,N_33250);
nand U36743 (N_36743,N_33430,N_34975);
xnor U36744 (N_36744,N_33940,N_34209);
nand U36745 (N_36745,N_33547,N_33618);
and U36746 (N_36746,N_33976,N_32963);
xnor U36747 (N_36747,N_33076,N_32535);
nor U36748 (N_36748,N_34754,N_33606);
and U36749 (N_36749,N_34725,N_34113);
and U36750 (N_36750,N_34944,N_34850);
nand U36751 (N_36751,N_34027,N_34771);
xnor U36752 (N_36752,N_34215,N_32615);
or U36753 (N_36753,N_33644,N_34057);
nand U36754 (N_36754,N_33755,N_34883);
nor U36755 (N_36755,N_33958,N_33479);
xnor U36756 (N_36756,N_33457,N_34727);
nor U36757 (N_36757,N_34618,N_34964);
and U36758 (N_36758,N_34009,N_33525);
nand U36759 (N_36759,N_34650,N_32621);
xor U36760 (N_36760,N_32519,N_34378);
or U36761 (N_36761,N_32718,N_33283);
nor U36762 (N_36762,N_32768,N_34883);
nor U36763 (N_36763,N_34610,N_32629);
or U36764 (N_36764,N_34775,N_34169);
nor U36765 (N_36765,N_33805,N_32780);
xor U36766 (N_36766,N_33108,N_34026);
nand U36767 (N_36767,N_33929,N_33133);
and U36768 (N_36768,N_34813,N_34425);
nor U36769 (N_36769,N_34166,N_32985);
nor U36770 (N_36770,N_34884,N_33675);
nor U36771 (N_36771,N_32741,N_32539);
and U36772 (N_36772,N_34246,N_32963);
nand U36773 (N_36773,N_32695,N_33040);
nand U36774 (N_36774,N_32774,N_33813);
nand U36775 (N_36775,N_33271,N_34217);
or U36776 (N_36776,N_33712,N_33907);
and U36777 (N_36777,N_32792,N_34307);
or U36778 (N_36778,N_33789,N_33576);
or U36779 (N_36779,N_34534,N_34590);
nand U36780 (N_36780,N_34085,N_34106);
xnor U36781 (N_36781,N_33629,N_33509);
or U36782 (N_36782,N_33524,N_34308);
and U36783 (N_36783,N_33362,N_32756);
and U36784 (N_36784,N_33582,N_34199);
and U36785 (N_36785,N_34257,N_34527);
nor U36786 (N_36786,N_34179,N_34793);
or U36787 (N_36787,N_34053,N_33069);
and U36788 (N_36788,N_33585,N_32810);
nand U36789 (N_36789,N_34874,N_33859);
nand U36790 (N_36790,N_33957,N_34889);
nand U36791 (N_36791,N_33304,N_34383);
and U36792 (N_36792,N_33922,N_34034);
or U36793 (N_36793,N_32886,N_33392);
or U36794 (N_36794,N_32868,N_33231);
and U36795 (N_36795,N_32794,N_32935);
and U36796 (N_36796,N_34693,N_34249);
or U36797 (N_36797,N_34462,N_33916);
nor U36798 (N_36798,N_34347,N_33459);
nor U36799 (N_36799,N_34791,N_33438);
nand U36800 (N_36800,N_32558,N_32726);
xnor U36801 (N_36801,N_34101,N_33875);
nor U36802 (N_36802,N_32725,N_34902);
or U36803 (N_36803,N_33294,N_33916);
and U36804 (N_36804,N_34575,N_34679);
nand U36805 (N_36805,N_32772,N_32917);
xnor U36806 (N_36806,N_33041,N_33543);
and U36807 (N_36807,N_33458,N_33010);
nand U36808 (N_36808,N_33873,N_34624);
nand U36809 (N_36809,N_34880,N_34793);
and U36810 (N_36810,N_34108,N_34965);
nor U36811 (N_36811,N_32626,N_33752);
and U36812 (N_36812,N_33414,N_33158);
or U36813 (N_36813,N_33225,N_33668);
nand U36814 (N_36814,N_33812,N_34918);
nor U36815 (N_36815,N_32996,N_33435);
xor U36816 (N_36816,N_33072,N_34949);
xor U36817 (N_36817,N_33772,N_33727);
and U36818 (N_36818,N_34498,N_32659);
xnor U36819 (N_36819,N_33099,N_33330);
xnor U36820 (N_36820,N_34187,N_34148);
xnor U36821 (N_36821,N_33441,N_33106);
xor U36822 (N_36822,N_33273,N_33973);
and U36823 (N_36823,N_33158,N_33633);
nand U36824 (N_36824,N_34156,N_34937);
and U36825 (N_36825,N_32523,N_34290);
and U36826 (N_36826,N_32577,N_34873);
xor U36827 (N_36827,N_34829,N_33506);
and U36828 (N_36828,N_33975,N_34403);
nor U36829 (N_36829,N_34794,N_33737);
nor U36830 (N_36830,N_34501,N_33069);
nor U36831 (N_36831,N_34715,N_33627);
nor U36832 (N_36832,N_34957,N_33992);
nand U36833 (N_36833,N_34283,N_33391);
and U36834 (N_36834,N_34823,N_32514);
nor U36835 (N_36835,N_34797,N_34003);
xnor U36836 (N_36836,N_34752,N_34893);
nor U36837 (N_36837,N_32988,N_34299);
nand U36838 (N_36838,N_34869,N_34300);
nand U36839 (N_36839,N_33225,N_32723);
and U36840 (N_36840,N_33637,N_34960);
or U36841 (N_36841,N_33761,N_33956);
nor U36842 (N_36842,N_33164,N_32905);
nand U36843 (N_36843,N_33232,N_33526);
and U36844 (N_36844,N_34447,N_34415);
and U36845 (N_36845,N_33410,N_32872);
or U36846 (N_36846,N_32666,N_34037);
nand U36847 (N_36847,N_33901,N_32590);
nand U36848 (N_36848,N_32653,N_33641);
or U36849 (N_36849,N_34454,N_32586);
nand U36850 (N_36850,N_33768,N_33694);
nor U36851 (N_36851,N_33507,N_34067);
nand U36852 (N_36852,N_32955,N_33481);
nand U36853 (N_36853,N_34311,N_32751);
or U36854 (N_36854,N_33100,N_34324);
nor U36855 (N_36855,N_34448,N_33472);
nand U36856 (N_36856,N_33240,N_34310);
and U36857 (N_36857,N_34656,N_33308);
nor U36858 (N_36858,N_32851,N_33271);
xor U36859 (N_36859,N_32985,N_34922);
and U36860 (N_36860,N_33092,N_32880);
nand U36861 (N_36861,N_33233,N_34625);
nor U36862 (N_36862,N_34222,N_33055);
nand U36863 (N_36863,N_33266,N_34209);
or U36864 (N_36864,N_34097,N_34732);
nand U36865 (N_36865,N_33045,N_34795);
nor U36866 (N_36866,N_33386,N_34178);
nor U36867 (N_36867,N_32583,N_33657);
nand U36868 (N_36868,N_33966,N_33616);
xor U36869 (N_36869,N_34966,N_33170);
or U36870 (N_36870,N_34279,N_34373);
and U36871 (N_36871,N_34083,N_34948);
and U36872 (N_36872,N_34407,N_33281);
nor U36873 (N_36873,N_33900,N_32611);
and U36874 (N_36874,N_32895,N_33709);
nor U36875 (N_36875,N_34235,N_34489);
nor U36876 (N_36876,N_33255,N_34197);
or U36877 (N_36877,N_33223,N_33854);
and U36878 (N_36878,N_33915,N_32747);
and U36879 (N_36879,N_33970,N_33529);
nand U36880 (N_36880,N_33241,N_32745);
nor U36881 (N_36881,N_33656,N_33299);
xor U36882 (N_36882,N_32825,N_32947);
or U36883 (N_36883,N_34200,N_34318);
nor U36884 (N_36884,N_34797,N_34977);
or U36885 (N_36885,N_32715,N_33776);
xor U36886 (N_36886,N_33436,N_34739);
nor U36887 (N_36887,N_32655,N_32968);
and U36888 (N_36888,N_32925,N_34317);
nand U36889 (N_36889,N_34813,N_32972);
and U36890 (N_36890,N_34652,N_33345);
nand U36891 (N_36891,N_34802,N_34386);
xnor U36892 (N_36892,N_33619,N_33088);
nand U36893 (N_36893,N_34641,N_32718);
or U36894 (N_36894,N_34989,N_34619);
nand U36895 (N_36895,N_33110,N_32801);
or U36896 (N_36896,N_34130,N_33247);
nor U36897 (N_36897,N_32533,N_34156);
nor U36898 (N_36898,N_34337,N_33962);
and U36899 (N_36899,N_34137,N_34315);
nor U36900 (N_36900,N_34164,N_33878);
xnor U36901 (N_36901,N_32997,N_33174);
xnor U36902 (N_36902,N_32654,N_32535);
nor U36903 (N_36903,N_32917,N_33707);
nand U36904 (N_36904,N_33748,N_32925);
xnor U36905 (N_36905,N_33457,N_33805);
xor U36906 (N_36906,N_32667,N_34461);
nand U36907 (N_36907,N_34712,N_34320);
nor U36908 (N_36908,N_33896,N_33719);
nand U36909 (N_36909,N_33404,N_33053);
nor U36910 (N_36910,N_33149,N_33466);
xor U36911 (N_36911,N_32527,N_34532);
nand U36912 (N_36912,N_33531,N_34537);
and U36913 (N_36913,N_34797,N_33040);
xnor U36914 (N_36914,N_33096,N_34249);
xor U36915 (N_36915,N_32777,N_33859);
nand U36916 (N_36916,N_34631,N_33746);
nor U36917 (N_36917,N_34398,N_34897);
nor U36918 (N_36918,N_34271,N_33039);
and U36919 (N_36919,N_34798,N_33312);
nor U36920 (N_36920,N_34817,N_33483);
xnor U36921 (N_36921,N_32619,N_34462);
or U36922 (N_36922,N_34594,N_34353);
nand U36923 (N_36923,N_33492,N_34953);
nor U36924 (N_36924,N_34961,N_34578);
nand U36925 (N_36925,N_34485,N_33075);
nor U36926 (N_36926,N_34548,N_34105);
nor U36927 (N_36927,N_32504,N_32767);
nor U36928 (N_36928,N_32691,N_33426);
or U36929 (N_36929,N_34189,N_32785);
nand U36930 (N_36930,N_33385,N_34327);
nor U36931 (N_36931,N_34252,N_34913);
or U36932 (N_36932,N_34872,N_33514);
nand U36933 (N_36933,N_32883,N_33939);
or U36934 (N_36934,N_33669,N_33852);
nor U36935 (N_36935,N_32763,N_32843);
nor U36936 (N_36936,N_32944,N_33883);
nand U36937 (N_36937,N_33785,N_33076);
and U36938 (N_36938,N_34025,N_34999);
and U36939 (N_36939,N_34094,N_32805);
or U36940 (N_36940,N_33290,N_33887);
xnor U36941 (N_36941,N_34403,N_34304);
nor U36942 (N_36942,N_33197,N_33255);
and U36943 (N_36943,N_34891,N_34355);
and U36944 (N_36944,N_32740,N_34833);
nand U36945 (N_36945,N_32911,N_34606);
and U36946 (N_36946,N_33372,N_33985);
nor U36947 (N_36947,N_33142,N_34176);
xor U36948 (N_36948,N_33728,N_33354);
nand U36949 (N_36949,N_34481,N_34649);
nor U36950 (N_36950,N_34624,N_34367);
or U36951 (N_36951,N_32676,N_33447);
xnor U36952 (N_36952,N_33793,N_34249);
nor U36953 (N_36953,N_34653,N_34788);
nor U36954 (N_36954,N_33612,N_34354);
or U36955 (N_36955,N_34151,N_32647);
and U36956 (N_36956,N_34011,N_34753);
or U36957 (N_36957,N_34901,N_34973);
nor U36958 (N_36958,N_33427,N_34609);
or U36959 (N_36959,N_33465,N_34550);
and U36960 (N_36960,N_32623,N_33753);
xor U36961 (N_36961,N_33256,N_34102);
nor U36962 (N_36962,N_32532,N_32608);
xnor U36963 (N_36963,N_33450,N_33911);
nor U36964 (N_36964,N_34133,N_34573);
or U36965 (N_36965,N_34657,N_33012);
and U36966 (N_36966,N_33883,N_33277);
and U36967 (N_36967,N_34272,N_32715);
or U36968 (N_36968,N_33699,N_34481);
nor U36969 (N_36969,N_32888,N_33154);
and U36970 (N_36970,N_33521,N_34778);
or U36971 (N_36971,N_33424,N_34807);
nand U36972 (N_36972,N_34051,N_32836);
nor U36973 (N_36973,N_34693,N_34958);
nor U36974 (N_36974,N_32965,N_33260);
or U36975 (N_36975,N_33621,N_34561);
nor U36976 (N_36976,N_34208,N_33683);
nor U36977 (N_36977,N_34373,N_32682);
or U36978 (N_36978,N_34385,N_34151);
xnor U36979 (N_36979,N_34424,N_34185);
or U36980 (N_36980,N_33167,N_34733);
or U36981 (N_36981,N_34974,N_33283);
nor U36982 (N_36982,N_33600,N_33146);
nor U36983 (N_36983,N_32787,N_34236);
or U36984 (N_36984,N_33590,N_33665);
xor U36985 (N_36985,N_34004,N_33119);
nand U36986 (N_36986,N_33786,N_34924);
xnor U36987 (N_36987,N_34034,N_34423);
xnor U36988 (N_36988,N_34712,N_32549);
and U36989 (N_36989,N_32533,N_33325);
and U36990 (N_36990,N_33865,N_33851);
nor U36991 (N_36991,N_34446,N_33478);
and U36992 (N_36992,N_32611,N_34208);
nor U36993 (N_36993,N_34873,N_32935);
or U36994 (N_36994,N_33246,N_34447);
and U36995 (N_36995,N_34120,N_33600);
and U36996 (N_36996,N_33448,N_32563);
nand U36997 (N_36997,N_34761,N_32591);
nor U36998 (N_36998,N_32822,N_33187);
xor U36999 (N_36999,N_32904,N_34551);
nor U37000 (N_37000,N_34063,N_32879);
nand U37001 (N_37001,N_34457,N_33438);
nand U37002 (N_37002,N_34372,N_32830);
nand U37003 (N_37003,N_33299,N_32660);
xnor U37004 (N_37004,N_34820,N_33336);
and U37005 (N_37005,N_33038,N_34601);
and U37006 (N_37006,N_33048,N_34860);
xor U37007 (N_37007,N_32556,N_32712);
nor U37008 (N_37008,N_34687,N_34664);
or U37009 (N_37009,N_34086,N_32578);
nand U37010 (N_37010,N_33510,N_33556);
or U37011 (N_37011,N_33437,N_34901);
xnor U37012 (N_37012,N_33172,N_32797);
and U37013 (N_37013,N_33120,N_34700);
or U37014 (N_37014,N_33126,N_33544);
xnor U37015 (N_37015,N_34540,N_33690);
xnor U37016 (N_37016,N_33595,N_34072);
xor U37017 (N_37017,N_32690,N_34980);
and U37018 (N_37018,N_34422,N_32732);
and U37019 (N_37019,N_34888,N_33886);
nand U37020 (N_37020,N_33697,N_33149);
nand U37021 (N_37021,N_32821,N_33800);
and U37022 (N_37022,N_32879,N_33209);
and U37023 (N_37023,N_32511,N_33075);
or U37024 (N_37024,N_33395,N_33704);
or U37025 (N_37025,N_33434,N_33626);
xor U37026 (N_37026,N_32656,N_34890);
or U37027 (N_37027,N_33710,N_32887);
xnor U37028 (N_37028,N_32685,N_32871);
xnor U37029 (N_37029,N_34238,N_34294);
nor U37030 (N_37030,N_34992,N_33490);
and U37031 (N_37031,N_33068,N_34810);
and U37032 (N_37032,N_33513,N_33027);
nand U37033 (N_37033,N_33181,N_33892);
nand U37034 (N_37034,N_34945,N_33520);
nand U37035 (N_37035,N_33604,N_33815);
nand U37036 (N_37036,N_34812,N_33333);
nand U37037 (N_37037,N_33527,N_33429);
xnor U37038 (N_37038,N_33198,N_34933);
nand U37039 (N_37039,N_33634,N_33548);
nand U37040 (N_37040,N_34278,N_34579);
or U37041 (N_37041,N_34479,N_32789);
nand U37042 (N_37042,N_32767,N_34769);
nand U37043 (N_37043,N_33861,N_34692);
and U37044 (N_37044,N_34942,N_34964);
nor U37045 (N_37045,N_33555,N_33213);
and U37046 (N_37046,N_33494,N_32878);
and U37047 (N_37047,N_33481,N_33811);
or U37048 (N_37048,N_34836,N_34058);
or U37049 (N_37049,N_33368,N_34252);
nor U37050 (N_37050,N_33695,N_33748);
nor U37051 (N_37051,N_32961,N_34564);
xnor U37052 (N_37052,N_32997,N_33872);
or U37053 (N_37053,N_34975,N_32564);
and U37054 (N_37054,N_34151,N_32854);
nand U37055 (N_37055,N_32965,N_34897);
or U37056 (N_37056,N_34024,N_33996);
nand U37057 (N_37057,N_34854,N_34051);
or U37058 (N_37058,N_34988,N_34658);
nand U37059 (N_37059,N_34364,N_34503);
and U37060 (N_37060,N_34470,N_34840);
or U37061 (N_37061,N_34722,N_33055);
or U37062 (N_37062,N_32678,N_34307);
nor U37063 (N_37063,N_33657,N_34145);
and U37064 (N_37064,N_34581,N_33131);
xor U37065 (N_37065,N_33195,N_34260);
nor U37066 (N_37066,N_34851,N_34398);
nor U37067 (N_37067,N_34611,N_34676);
and U37068 (N_37068,N_33066,N_32972);
xor U37069 (N_37069,N_34073,N_34942);
and U37070 (N_37070,N_34702,N_34826);
xor U37071 (N_37071,N_34120,N_33959);
xnor U37072 (N_37072,N_32863,N_33720);
or U37073 (N_37073,N_32737,N_34267);
and U37074 (N_37074,N_34226,N_32627);
xor U37075 (N_37075,N_34805,N_33597);
nor U37076 (N_37076,N_34363,N_34476);
nor U37077 (N_37077,N_34653,N_32957);
or U37078 (N_37078,N_34607,N_34260);
and U37079 (N_37079,N_33559,N_33764);
and U37080 (N_37080,N_32790,N_32884);
nor U37081 (N_37081,N_33416,N_34215);
and U37082 (N_37082,N_34012,N_32954);
or U37083 (N_37083,N_33975,N_33460);
and U37084 (N_37084,N_33479,N_33444);
nand U37085 (N_37085,N_34568,N_34452);
nor U37086 (N_37086,N_33315,N_33346);
xnor U37087 (N_37087,N_32666,N_33011);
and U37088 (N_37088,N_32902,N_33753);
nor U37089 (N_37089,N_33360,N_34249);
xor U37090 (N_37090,N_33586,N_33227);
nand U37091 (N_37091,N_33304,N_32562);
xor U37092 (N_37092,N_33141,N_34542);
and U37093 (N_37093,N_33291,N_33264);
xnor U37094 (N_37094,N_33509,N_33638);
xor U37095 (N_37095,N_33678,N_34521);
nor U37096 (N_37096,N_34338,N_34270);
xor U37097 (N_37097,N_33206,N_32692);
nand U37098 (N_37098,N_34116,N_33298);
nand U37099 (N_37099,N_34637,N_33741);
xnor U37100 (N_37100,N_33603,N_34452);
nand U37101 (N_37101,N_32644,N_33016);
nor U37102 (N_37102,N_34944,N_34080);
nand U37103 (N_37103,N_32555,N_34626);
xnor U37104 (N_37104,N_34906,N_34846);
and U37105 (N_37105,N_32714,N_34935);
or U37106 (N_37106,N_34926,N_34983);
nand U37107 (N_37107,N_34050,N_34082);
or U37108 (N_37108,N_34721,N_33109);
and U37109 (N_37109,N_34422,N_32742);
xnor U37110 (N_37110,N_34738,N_34657);
nor U37111 (N_37111,N_34831,N_33008);
nor U37112 (N_37112,N_32918,N_33796);
nand U37113 (N_37113,N_34228,N_33574);
xnor U37114 (N_37114,N_32968,N_34857);
and U37115 (N_37115,N_34798,N_34473);
and U37116 (N_37116,N_33703,N_33178);
xor U37117 (N_37117,N_34177,N_34737);
nand U37118 (N_37118,N_33939,N_34820);
or U37119 (N_37119,N_33157,N_33083);
nand U37120 (N_37120,N_33022,N_33774);
or U37121 (N_37121,N_33068,N_34774);
nand U37122 (N_37122,N_34443,N_34641);
and U37123 (N_37123,N_33948,N_34799);
and U37124 (N_37124,N_33679,N_33049);
and U37125 (N_37125,N_34291,N_33555);
nand U37126 (N_37126,N_33662,N_33382);
xor U37127 (N_37127,N_32655,N_34740);
or U37128 (N_37128,N_34630,N_32976);
or U37129 (N_37129,N_34236,N_33355);
or U37130 (N_37130,N_34101,N_33100);
xnor U37131 (N_37131,N_34546,N_32928);
and U37132 (N_37132,N_33517,N_32744);
or U37133 (N_37133,N_33875,N_33964);
nand U37134 (N_37134,N_32576,N_32514);
xnor U37135 (N_37135,N_33898,N_33720);
nor U37136 (N_37136,N_33781,N_33569);
and U37137 (N_37137,N_33038,N_33295);
xnor U37138 (N_37138,N_33589,N_34241);
nand U37139 (N_37139,N_32534,N_33560);
nor U37140 (N_37140,N_33921,N_33494);
and U37141 (N_37141,N_33359,N_34865);
and U37142 (N_37142,N_34982,N_32701);
and U37143 (N_37143,N_33702,N_33068);
nor U37144 (N_37144,N_34121,N_33574);
xor U37145 (N_37145,N_32576,N_33089);
nor U37146 (N_37146,N_33812,N_33695);
nand U37147 (N_37147,N_34135,N_32507);
nand U37148 (N_37148,N_34074,N_34294);
and U37149 (N_37149,N_32576,N_34467);
xnor U37150 (N_37150,N_34891,N_32875);
and U37151 (N_37151,N_34027,N_32901);
nand U37152 (N_37152,N_33029,N_33085);
nor U37153 (N_37153,N_33366,N_33869);
nand U37154 (N_37154,N_33135,N_34348);
nand U37155 (N_37155,N_33065,N_33834);
nand U37156 (N_37156,N_33434,N_32642);
xnor U37157 (N_37157,N_34953,N_34979);
nand U37158 (N_37158,N_32978,N_34409);
and U37159 (N_37159,N_33873,N_33960);
nor U37160 (N_37160,N_33667,N_33468);
or U37161 (N_37161,N_32614,N_33229);
and U37162 (N_37162,N_34792,N_33915);
or U37163 (N_37163,N_33078,N_33358);
and U37164 (N_37164,N_33661,N_33227);
nor U37165 (N_37165,N_34017,N_32783);
and U37166 (N_37166,N_32889,N_34181);
or U37167 (N_37167,N_33751,N_34776);
xor U37168 (N_37168,N_33010,N_33198);
or U37169 (N_37169,N_34744,N_33555);
and U37170 (N_37170,N_34842,N_33964);
xnor U37171 (N_37171,N_33247,N_34721);
and U37172 (N_37172,N_34490,N_33082);
and U37173 (N_37173,N_33496,N_33383);
nor U37174 (N_37174,N_32906,N_34788);
nand U37175 (N_37175,N_34495,N_34157);
or U37176 (N_37176,N_34047,N_34441);
or U37177 (N_37177,N_33297,N_32559);
nor U37178 (N_37178,N_33449,N_32617);
and U37179 (N_37179,N_34365,N_32590);
nand U37180 (N_37180,N_33162,N_34572);
or U37181 (N_37181,N_32975,N_34272);
nand U37182 (N_37182,N_33194,N_32844);
and U37183 (N_37183,N_32937,N_34160);
or U37184 (N_37184,N_33683,N_33735);
xor U37185 (N_37185,N_34597,N_34055);
and U37186 (N_37186,N_33868,N_33421);
and U37187 (N_37187,N_33551,N_33117);
nor U37188 (N_37188,N_34950,N_34057);
xor U37189 (N_37189,N_33107,N_33658);
or U37190 (N_37190,N_33664,N_34103);
xnor U37191 (N_37191,N_34956,N_32615);
nand U37192 (N_37192,N_32731,N_34572);
xor U37193 (N_37193,N_33523,N_33751);
nand U37194 (N_37194,N_33424,N_34077);
or U37195 (N_37195,N_32599,N_34283);
and U37196 (N_37196,N_34618,N_34006);
and U37197 (N_37197,N_33059,N_33830);
nor U37198 (N_37198,N_32977,N_33067);
and U37199 (N_37199,N_33816,N_33487);
and U37200 (N_37200,N_34162,N_33992);
nor U37201 (N_37201,N_34091,N_32774);
xnor U37202 (N_37202,N_33774,N_33305);
and U37203 (N_37203,N_33200,N_32625);
nor U37204 (N_37204,N_32726,N_33279);
or U37205 (N_37205,N_34364,N_32820);
and U37206 (N_37206,N_33086,N_34170);
and U37207 (N_37207,N_34820,N_32623);
or U37208 (N_37208,N_34798,N_34437);
and U37209 (N_37209,N_34395,N_33877);
nor U37210 (N_37210,N_32524,N_32835);
nor U37211 (N_37211,N_34796,N_33415);
nor U37212 (N_37212,N_34727,N_34994);
or U37213 (N_37213,N_33875,N_34678);
xnor U37214 (N_37214,N_33512,N_33387);
or U37215 (N_37215,N_33126,N_34170);
and U37216 (N_37216,N_34553,N_32622);
and U37217 (N_37217,N_33264,N_33891);
and U37218 (N_37218,N_33536,N_34749);
and U37219 (N_37219,N_33526,N_34451);
xor U37220 (N_37220,N_33025,N_32736);
or U37221 (N_37221,N_34744,N_33600);
nand U37222 (N_37222,N_33735,N_32901);
xnor U37223 (N_37223,N_34152,N_32535);
nand U37224 (N_37224,N_33541,N_33222);
or U37225 (N_37225,N_32669,N_33682);
and U37226 (N_37226,N_34524,N_33229);
or U37227 (N_37227,N_32828,N_34750);
and U37228 (N_37228,N_34200,N_34084);
nand U37229 (N_37229,N_34542,N_33541);
nand U37230 (N_37230,N_33548,N_34185);
and U37231 (N_37231,N_34786,N_34667);
nand U37232 (N_37232,N_34453,N_34900);
and U37233 (N_37233,N_34726,N_34768);
or U37234 (N_37234,N_33033,N_33209);
nand U37235 (N_37235,N_34101,N_33907);
nor U37236 (N_37236,N_33421,N_34366);
nand U37237 (N_37237,N_33096,N_33961);
or U37238 (N_37238,N_34021,N_34123);
nand U37239 (N_37239,N_33171,N_33579);
and U37240 (N_37240,N_34450,N_32901);
nand U37241 (N_37241,N_32605,N_34347);
nor U37242 (N_37242,N_34504,N_33534);
or U37243 (N_37243,N_33813,N_34819);
nor U37244 (N_37244,N_34678,N_34340);
nand U37245 (N_37245,N_34981,N_34451);
nor U37246 (N_37246,N_33954,N_34503);
or U37247 (N_37247,N_33376,N_34528);
xor U37248 (N_37248,N_32811,N_34278);
nor U37249 (N_37249,N_34531,N_34677);
nand U37250 (N_37250,N_34473,N_33198);
and U37251 (N_37251,N_32510,N_34370);
nor U37252 (N_37252,N_32852,N_34220);
xor U37253 (N_37253,N_34093,N_34071);
and U37254 (N_37254,N_34225,N_33747);
xor U37255 (N_37255,N_33183,N_33085);
nand U37256 (N_37256,N_34196,N_32808);
nand U37257 (N_37257,N_33221,N_32850);
or U37258 (N_37258,N_33573,N_34986);
nand U37259 (N_37259,N_34279,N_34242);
xor U37260 (N_37260,N_34503,N_32808);
nand U37261 (N_37261,N_34639,N_34186);
or U37262 (N_37262,N_33682,N_34317);
nand U37263 (N_37263,N_34815,N_34169);
xnor U37264 (N_37264,N_34479,N_33424);
nor U37265 (N_37265,N_33329,N_33052);
or U37266 (N_37266,N_32521,N_32648);
xor U37267 (N_37267,N_34415,N_34265);
nand U37268 (N_37268,N_33272,N_34967);
nor U37269 (N_37269,N_34603,N_33468);
nor U37270 (N_37270,N_32588,N_34813);
and U37271 (N_37271,N_32635,N_34220);
or U37272 (N_37272,N_33061,N_34086);
nand U37273 (N_37273,N_34383,N_33609);
or U37274 (N_37274,N_33239,N_32890);
xor U37275 (N_37275,N_33323,N_34709);
nor U37276 (N_37276,N_34213,N_32675);
xor U37277 (N_37277,N_34339,N_33262);
xnor U37278 (N_37278,N_34679,N_34721);
xnor U37279 (N_37279,N_33894,N_34523);
nand U37280 (N_37280,N_33582,N_33409);
xnor U37281 (N_37281,N_33135,N_33824);
or U37282 (N_37282,N_33767,N_32860);
or U37283 (N_37283,N_33114,N_33244);
and U37284 (N_37284,N_33452,N_32783);
or U37285 (N_37285,N_34092,N_34296);
or U37286 (N_37286,N_34258,N_33483);
or U37287 (N_37287,N_32849,N_33238);
xor U37288 (N_37288,N_32894,N_33032);
or U37289 (N_37289,N_33842,N_33243);
nand U37290 (N_37290,N_34481,N_34081);
xnor U37291 (N_37291,N_34507,N_34902);
and U37292 (N_37292,N_32903,N_33712);
xor U37293 (N_37293,N_34524,N_34297);
nand U37294 (N_37294,N_34722,N_34984);
and U37295 (N_37295,N_34102,N_32581);
or U37296 (N_37296,N_34108,N_34657);
and U37297 (N_37297,N_34906,N_33918);
and U37298 (N_37298,N_34251,N_33925);
xnor U37299 (N_37299,N_32951,N_34870);
xnor U37300 (N_37300,N_32694,N_34529);
and U37301 (N_37301,N_32883,N_33365);
nand U37302 (N_37302,N_33930,N_32932);
and U37303 (N_37303,N_34773,N_32746);
and U37304 (N_37304,N_33563,N_33003);
nor U37305 (N_37305,N_34200,N_32759);
and U37306 (N_37306,N_32754,N_33932);
nor U37307 (N_37307,N_33301,N_34851);
nand U37308 (N_37308,N_34440,N_34259);
or U37309 (N_37309,N_33123,N_33769);
and U37310 (N_37310,N_34588,N_34341);
nor U37311 (N_37311,N_32850,N_34909);
nor U37312 (N_37312,N_32571,N_32609);
nor U37313 (N_37313,N_34785,N_34655);
or U37314 (N_37314,N_33630,N_34008);
and U37315 (N_37315,N_34594,N_34250);
nand U37316 (N_37316,N_33151,N_34139);
and U37317 (N_37317,N_33273,N_33965);
xnor U37318 (N_37318,N_32551,N_34055);
nand U37319 (N_37319,N_33825,N_33345);
nand U37320 (N_37320,N_34804,N_34159);
nand U37321 (N_37321,N_34823,N_32654);
or U37322 (N_37322,N_33264,N_33491);
nor U37323 (N_37323,N_33241,N_34583);
and U37324 (N_37324,N_34489,N_32856);
nand U37325 (N_37325,N_33847,N_33921);
or U37326 (N_37326,N_33602,N_32666);
and U37327 (N_37327,N_34457,N_32586);
nand U37328 (N_37328,N_33322,N_33407);
or U37329 (N_37329,N_32572,N_33430);
nand U37330 (N_37330,N_34238,N_34489);
or U37331 (N_37331,N_33099,N_34001);
nand U37332 (N_37332,N_32688,N_34311);
nor U37333 (N_37333,N_32520,N_32906);
nor U37334 (N_37334,N_32621,N_33168);
nor U37335 (N_37335,N_34368,N_33711);
xor U37336 (N_37336,N_34414,N_32851);
or U37337 (N_37337,N_33310,N_33438);
and U37338 (N_37338,N_33600,N_33114);
xnor U37339 (N_37339,N_33957,N_33928);
and U37340 (N_37340,N_33326,N_34002);
nand U37341 (N_37341,N_34140,N_34193);
nand U37342 (N_37342,N_33330,N_33298);
and U37343 (N_37343,N_33615,N_34159);
nand U37344 (N_37344,N_32794,N_34698);
nor U37345 (N_37345,N_34839,N_34637);
xnor U37346 (N_37346,N_34709,N_32736);
nand U37347 (N_37347,N_33266,N_34418);
nor U37348 (N_37348,N_34061,N_33147);
and U37349 (N_37349,N_33206,N_34486);
nand U37350 (N_37350,N_33479,N_33880);
and U37351 (N_37351,N_34450,N_32929);
and U37352 (N_37352,N_32759,N_32956);
nor U37353 (N_37353,N_33026,N_33905);
xnor U37354 (N_37354,N_34159,N_32585);
xnor U37355 (N_37355,N_33750,N_34577);
nor U37356 (N_37356,N_32659,N_34400);
xor U37357 (N_37357,N_34601,N_34235);
and U37358 (N_37358,N_34635,N_32576);
and U37359 (N_37359,N_34760,N_32930);
xnor U37360 (N_37360,N_34766,N_32642);
nand U37361 (N_37361,N_32561,N_33205);
or U37362 (N_37362,N_33514,N_33954);
nor U37363 (N_37363,N_34448,N_33773);
or U37364 (N_37364,N_33557,N_33968);
nor U37365 (N_37365,N_33165,N_33897);
or U37366 (N_37366,N_34412,N_33636);
nor U37367 (N_37367,N_33898,N_32837);
nor U37368 (N_37368,N_33462,N_33554);
nand U37369 (N_37369,N_34373,N_33399);
or U37370 (N_37370,N_34395,N_33811);
nor U37371 (N_37371,N_33352,N_32922);
nand U37372 (N_37372,N_33370,N_34297);
xnor U37373 (N_37373,N_33110,N_33849);
or U37374 (N_37374,N_33825,N_34292);
xnor U37375 (N_37375,N_33302,N_34856);
and U37376 (N_37376,N_33699,N_33032);
nand U37377 (N_37377,N_33364,N_34684);
or U37378 (N_37378,N_33754,N_33035);
nand U37379 (N_37379,N_33693,N_33565);
and U37380 (N_37380,N_33307,N_34474);
and U37381 (N_37381,N_33205,N_33436);
xor U37382 (N_37382,N_34117,N_34923);
and U37383 (N_37383,N_33756,N_32927);
and U37384 (N_37384,N_34313,N_32793);
nand U37385 (N_37385,N_34333,N_33683);
nor U37386 (N_37386,N_33665,N_34164);
or U37387 (N_37387,N_32834,N_34259);
xor U37388 (N_37388,N_34274,N_32745);
or U37389 (N_37389,N_32691,N_34805);
nor U37390 (N_37390,N_33337,N_33518);
nor U37391 (N_37391,N_32721,N_34930);
nor U37392 (N_37392,N_33109,N_32726);
or U37393 (N_37393,N_34109,N_33286);
xnor U37394 (N_37394,N_34430,N_33789);
nand U37395 (N_37395,N_34228,N_34218);
nand U37396 (N_37396,N_32781,N_32787);
nand U37397 (N_37397,N_34248,N_34701);
and U37398 (N_37398,N_34852,N_33909);
nand U37399 (N_37399,N_33824,N_34479);
nor U37400 (N_37400,N_34907,N_33051);
nand U37401 (N_37401,N_32676,N_33237);
or U37402 (N_37402,N_33750,N_33524);
and U37403 (N_37403,N_34442,N_34517);
or U37404 (N_37404,N_34128,N_34126);
or U37405 (N_37405,N_32768,N_32644);
and U37406 (N_37406,N_33476,N_32676);
xor U37407 (N_37407,N_33852,N_34562);
nor U37408 (N_37408,N_32586,N_34990);
nor U37409 (N_37409,N_34800,N_33575);
nand U37410 (N_37410,N_34353,N_33786);
and U37411 (N_37411,N_32638,N_32795);
or U37412 (N_37412,N_34555,N_33558);
nand U37413 (N_37413,N_34887,N_33411);
and U37414 (N_37414,N_33624,N_34361);
xnor U37415 (N_37415,N_34829,N_33790);
and U37416 (N_37416,N_33563,N_33737);
or U37417 (N_37417,N_33163,N_33682);
or U37418 (N_37418,N_34436,N_33267);
nand U37419 (N_37419,N_33201,N_34983);
nand U37420 (N_37420,N_33548,N_34414);
and U37421 (N_37421,N_34947,N_32998);
nand U37422 (N_37422,N_33526,N_34650);
xnor U37423 (N_37423,N_34735,N_32582);
nor U37424 (N_37424,N_34842,N_33756);
nor U37425 (N_37425,N_34671,N_33201);
nand U37426 (N_37426,N_32763,N_32991);
or U37427 (N_37427,N_33765,N_33992);
nand U37428 (N_37428,N_34883,N_34413);
nand U37429 (N_37429,N_33090,N_33519);
xor U37430 (N_37430,N_33097,N_34559);
xnor U37431 (N_37431,N_33182,N_34324);
or U37432 (N_37432,N_34041,N_34030);
nor U37433 (N_37433,N_32763,N_34584);
and U37434 (N_37434,N_34956,N_34415);
nor U37435 (N_37435,N_34584,N_34266);
nor U37436 (N_37436,N_32571,N_33175);
or U37437 (N_37437,N_34143,N_34345);
xnor U37438 (N_37438,N_33566,N_34054);
and U37439 (N_37439,N_34849,N_32612);
nand U37440 (N_37440,N_33870,N_32500);
xnor U37441 (N_37441,N_34811,N_33243);
nor U37442 (N_37442,N_33284,N_34916);
and U37443 (N_37443,N_32679,N_34391);
xnor U37444 (N_37444,N_34967,N_34682);
nand U37445 (N_37445,N_34384,N_33023);
or U37446 (N_37446,N_32516,N_32911);
xnor U37447 (N_37447,N_32853,N_33986);
or U37448 (N_37448,N_33837,N_32881);
xor U37449 (N_37449,N_34739,N_33121);
nor U37450 (N_37450,N_32999,N_34613);
xor U37451 (N_37451,N_33463,N_33220);
nor U37452 (N_37452,N_32809,N_32893);
nand U37453 (N_37453,N_34835,N_34129);
and U37454 (N_37454,N_33599,N_32610);
or U37455 (N_37455,N_34268,N_32567);
nand U37456 (N_37456,N_33108,N_33527);
and U37457 (N_37457,N_33308,N_33151);
and U37458 (N_37458,N_34326,N_34966);
nand U37459 (N_37459,N_34849,N_33112);
nor U37460 (N_37460,N_33687,N_34826);
and U37461 (N_37461,N_33582,N_33361);
nor U37462 (N_37462,N_34771,N_33435);
or U37463 (N_37463,N_34224,N_33215);
and U37464 (N_37464,N_32895,N_33303);
nand U37465 (N_37465,N_34538,N_34369);
xor U37466 (N_37466,N_33561,N_33216);
or U37467 (N_37467,N_34160,N_32671);
and U37468 (N_37468,N_32655,N_34027);
nor U37469 (N_37469,N_33775,N_34479);
or U37470 (N_37470,N_34994,N_33063);
or U37471 (N_37471,N_34189,N_34489);
or U37472 (N_37472,N_33348,N_33963);
or U37473 (N_37473,N_33463,N_32816);
nor U37474 (N_37474,N_33743,N_32684);
and U37475 (N_37475,N_33123,N_34523);
nand U37476 (N_37476,N_32938,N_32790);
nand U37477 (N_37477,N_32978,N_32523);
and U37478 (N_37478,N_34879,N_32695);
nor U37479 (N_37479,N_32510,N_34348);
or U37480 (N_37480,N_32781,N_32960);
or U37481 (N_37481,N_34922,N_33467);
nand U37482 (N_37482,N_33863,N_34269);
and U37483 (N_37483,N_33526,N_34129);
or U37484 (N_37484,N_33726,N_33238);
and U37485 (N_37485,N_33578,N_33525);
nor U37486 (N_37486,N_33916,N_34516);
xor U37487 (N_37487,N_34917,N_33292);
or U37488 (N_37488,N_32927,N_33577);
nor U37489 (N_37489,N_34679,N_34077);
and U37490 (N_37490,N_33655,N_34972);
nand U37491 (N_37491,N_33638,N_34465);
nor U37492 (N_37492,N_33219,N_33857);
nor U37493 (N_37493,N_34323,N_34025);
nor U37494 (N_37494,N_33265,N_32602);
and U37495 (N_37495,N_32769,N_34447);
xor U37496 (N_37496,N_33475,N_34754);
nand U37497 (N_37497,N_34886,N_33582);
or U37498 (N_37498,N_34705,N_33575);
nor U37499 (N_37499,N_33060,N_33687);
and U37500 (N_37500,N_35534,N_35416);
nor U37501 (N_37501,N_35602,N_35289);
and U37502 (N_37502,N_35294,N_36549);
xor U37503 (N_37503,N_36631,N_35048);
nand U37504 (N_37504,N_35234,N_35514);
or U37505 (N_37505,N_36965,N_36306);
nand U37506 (N_37506,N_36402,N_35722);
or U37507 (N_37507,N_35035,N_37092);
nand U37508 (N_37508,N_37183,N_36228);
xor U37509 (N_37509,N_35355,N_35475);
xnor U37510 (N_37510,N_37000,N_37303);
nand U37511 (N_37511,N_35821,N_36997);
and U37512 (N_37512,N_37395,N_37279);
and U37513 (N_37513,N_37456,N_37075);
or U37514 (N_37514,N_36481,N_36167);
and U37515 (N_37515,N_35948,N_36084);
nor U37516 (N_37516,N_35756,N_35606);
and U37517 (N_37517,N_37149,N_35467);
or U37518 (N_37518,N_37043,N_35211);
nand U37519 (N_37519,N_35703,N_36671);
nand U37520 (N_37520,N_35445,N_36243);
nor U37521 (N_37521,N_36685,N_37473);
nand U37522 (N_37522,N_36390,N_36598);
and U37523 (N_37523,N_35666,N_36363);
or U37524 (N_37524,N_37041,N_35548);
nand U37525 (N_37525,N_36908,N_37181);
nor U37526 (N_37526,N_37009,N_37046);
xor U37527 (N_37527,N_37492,N_36160);
xor U37528 (N_37528,N_35000,N_35997);
nand U37529 (N_37529,N_36054,N_35581);
nor U37530 (N_37530,N_36576,N_36017);
and U37531 (N_37531,N_36772,N_37047);
nand U37532 (N_37532,N_36894,N_36127);
nand U37533 (N_37533,N_36784,N_36162);
and U37534 (N_37534,N_35743,N_35681);
or U37535 (N_37535,N_35377,N_36432);
and U37536 (N_37536,N_37246,N_35600);
or U37537 (N_37537,N_37158,N_36220);
xnor U37538 (N_37538,N_35442,N_36603);
xor U37539 (N_37539,N_35668,N_36821);
xnor U37540 (N_37540,N_36526,N_36666);
xnor U37541 (N_37541,N_37272,N_35674);
xnor U37542 (N_37542,N_37162,N_35178);
nor U37543 (N_37543,N_37485,N_36977);
nand U37544 (N_37544,N_36878,N_36869);
xor U37545 (N_37545,N_35777,N_35111);
nand U37546 (N_37546,N_35582,N_36022);
and U37547 (N_37547,N_35784,N_35345);
and U37548 (N_37548,N_36128,N_36214);
nand U37549 (N_37549,N_36699,N_35274);
xnor U37550 (N_37550,N_35932,N_36504);
and U37551 (N_37551,N_35151,N_35812);
and U37552 (N_37552,N_35335,N_36523);
xor U37553 (N_37553,N_36799,N_37171);
or U37554 (N_37554,N_36832,N_37103);
and U37555 (N_37555,N_35008,N_35736);
and U37556 (N_37556,N_37267,N_35109);
nand U37557 (N_37557,N_36328,N_37418);
or U37558 (N_37558,N_36650,N_36672);
xor U37559 (N_37559,N_36495,N_36572);
nor U37560 (N_37560,N_35305,N_36736);
nor U37561 (N_37561,N_35291,N_36122);
nand U37562 (N_37562,N_35626,N_36461);
nand U37563 (N_37563,N_36825,N_35086);
or U37564 (N_37564,N_36662,N_35707);
or U37565 (N_37565,N_35299,N_36260);
nand U37566 (N_37566,N_36134,N_35292);
nor U37567 (N_37567,N_36048,N_35911);
or U37568 (N_37568,N_36651,N_35120);
nor U37569 (N_37569,N_35861,N_35860);
nor U37570 (N_37570,N_35824,N_36993);
nand U37571 (N_37571,N_37381,N_37433);
xor U37572 (N_37572,N_36853,N_36342);
nor U37573 (N_37573,N_36268,N_36452);
nor U37574 (N_37574,N_36326,N_36300);
xor U37575 (N_37575,N_37141,N_36680);
nand U37576 (N_37576,N_36779,N_35916);
nor U37577 (N_37577,N_37196,N_35568);
and U37578 (N_37578,N_36880,N_36205);
and U37579 (N_37579,N_35934,N_35701);
and U37580 (N_37580,N_37403,N_36034);
or U37581 (N_37581,N_35883,N_35608);
and U37582 (N_37582,N_35100,N_36348);
and U37583 (N_37583,N_36884,N_37203);
or U37584 (N_37584,N_36798,N_37010);
and U37585 (N_37585,N_35767,N_36212);
xnor U37586 (N_37586,N_35036,N_35301);
and U37587 (N_37587,N_35659,N_37087);
or U37588 (N_37588,N_35448,N_35819);
and U37589 (N_37589,N_37057,N_36778);
xnor U37590 (N_37590,N_37461,N_36294);
or U37591 (N_37591,N_35715,N_35252);
nand U37592 (N_37592,N_37095,N_35167);
nand U37593 (N_37593,N_37253,N_35363);
and U37594 (N_37594,N_35544,N_36286);
nand U37595 (N_37595,N_37412,N_36618);
nor U37596 (N_37596,N_35906,N_35254);
nand U37597 (N_37597,N_36824,N_37054);
or U37598 (N_37598,N_36649,N_37232);
nor U37599 (N_37599,N_37289,N_36972);
and U37600 (N_37600,N_35327,N_37310);
nor U37601 (N_37601,N_36942,N_36040);
and U37602 (N_37602,N_35638,N_35936);
nor U37603 (N_37603,N_37135,N_36979);
and U37604 (N_37604,N_36907,N_35221);
and U37605 (N_37605,N_36404,N_35399);
or U37606 (N_37606,N_36709,N_37308);
nor U37607 (N_37607,N_36705,N_37191);
nand U37608 (N_37608,N_35712,N_35170);
nand U37609 (N_37609,N_35610,N_36609);
nor U37610 (N_37610,N_35910,N_37265);
nor U37611 (N_37611,N_37346,N_36640);
xor U37612 (N_37612,N_36104,N_36539);
xor U37613 (N_37613,N_36937,N_36746);
nor U37614 (N_37614,N_36371,N_36531);
and U37615 (N_37615,N_35218,N_35622);
or U37616 (N_37616,N_35951,N_35116);
xnor U37617 (N_37617,N_37388,N_35280);
or U37618 (N_37618,N_35466,N_35907);
and U37619 (N_37619,N_35527,N_36773);
xnor U37620 (N_37620,N_36453,N_35990);
nor U37621 (N_37621,N_36958,N_36612);
nor U37622 (N_37622,N_35310,N_36164);
xor U37623 (N_37623,N_36838,N_35238);
nand U37624 (N_37624,N_36020,N_36053);
xor U37625 (N_37625,N_35770,N_37404);
or U37626 (N_37626,N_36497,N_35323);
or U37627 (N_37627,N_36849,N_35727);
nor U37628 (N_37628,N_36403,N_37490);
xor U37629 (N_37629,N_36026,N_36817);
nor U37630 (N_37630,N_37173,N_37193);
nand U37631 (N_37631,N_36322,N_36590);
and U37632 (N_37632,N_36716,N_36614);
and U37633 (N_37633,N_35437,N_37122);
or U37634 (N_37634,N_37013,N_36629);
xnor U37635 (N_37635,N_35615,N_36941);
or U37636 (N_37636,N_35944,N_35156);
nand U37637 (N_37637,N_36419,N_36482);
and U37638 (N_37638,N_37157,N_37164);
and U37639 (N_37639,N_36242,N_36414);
nand U37640 (N_37640,N_37263,N_35556);
xor U37641 (N_37641,N_36006,N_36186);
nand U37642 (N_37642,N_37194,N_36987);
nand U37643 (N_37643,N_35746,N_36063);
and U37644 (N_37644,N_35801,N_35235);
nor U37645 (N_37645,N_36559,N_35020);
and U37646 (N_37646,N_36510,N_37179);
nand U37647 (N_37647,N_35478,N_36912);
nand U37648 (N_37648,N_35764,N_35364);
or U37649 (N_37649,N_36265,N_35950);
nand U37650 (N_37650,N_35422,N_37148);
nand U37651 (N_37651,N_36333,N_37423);
or U37652 (N_37652,N_37118,N_36693);
nand U37653 (N_37653,N_36873,N_35137);
xor U37654 (N_37654,N_35952,N_35820);
and U37655 (N_37655,N_36995,N_35441);
or U37656 (N_37656,N_37133,N_35477);
nor U37657 (N_37657,N_35044,N_36928);
nor U37658 (N_37658,N_35631,N_35888);
or U37659 (N_37659,N_35644,N_35553);
nor U37660 (N_37660,N_35033,N_35434);
and U37661 (N_37661,N_36168,N_37331);
and U37662 (N_37662,N_35172,N_35693);
and U37663 (N_37663,N_36715,N_35967);
and U37664 (N_37664,N_37190,N_37094);
nor U37665 (N_37665,N_36280,N_36145);
nand U37666 (N_37666,N_35256,N_37254);
and U37667 (N_37667,N_35584,N_35190);
xnor U37668 (N_37668,N_35068,N_36089);
nor U37669 (N_37669,N_35460,N_35830);
nor U37670 (N_37670,N_35285,N_35601);
xnor U37671 (N_37671,N_36289,N_37019);
nand U37672 (N_37672,N_36253,N_35128);
or U37673 (N_37673,N_35419,N_36565);
nor U37674 (N_37674,N_35253,N_36855);
nand U37675 (N_37675,N_35745,N_36094);
xor U37676 (N_37676,N_36115,N_36172);
nand U37677 (N_37677,N_35829,N_35516);
xor U37678 (N_37678,N_36037,N_36811);
or U37679 (N_37679,N_36386,N_36501);
nor U37680 (N_37680,N_35426,N_37322);
or U37681 (N_37681,N_36223,N_37342);
and U37682 (N_37682,N_35920,N_35270);
nor U37683 (N_37683,N_36263,N_37305);
xor U37684 (N_37684,N_37031,N_35108);
xnor U37685 (N_37685,N_35430,N_36763);
and U37686 (N_37686,N_36702,N_37393);
nand U37687 (N_37687,N_36126,N_35667);
and U37688 (N_37688,N_36573,N_36370);
xor U37689 (N_37689,N_37207,N_37335);
or U37690 (N_37690,N_35134,N_36428);
or U37691 (N_37691,N_36235,N_35841);
or U37692 (N_37692,N_37291,N_37273);
nor U37693 (N_37693,N_36888,N_35457);
xor U37694 (N_37694,N_36233,N_37338);
nand U37695 (N_37695,N_35979,N_36443);
and U37696 (N_37696,N_37449,N_35902);
nor U37697 (N_37697,N_35655,N_36456);
nand U37698 (N_37698,N_36589,N_36733);
xnor U37699 (N_37699,N_35236,N_35896);
and U37700 (N_37700,N_37442,N_35941);
and U37701 (N_37701,N_36157,N_36473);
xnor U37702 (N_37702,N_35069,N_36871);
nor U37703 (N_37703,N_35873,N_35415);
nor U37704 (N_37704,N_36757,N_36295);
and U37705 (N_37705,N_35969,N_35213);
and U37706 (N_37706,N_35724,N_37287);
nor U37707 (N_37707,N_36303,N_36571);
or U37708 (N_37708,N_35398,N_35023);
nor U37709 (N_37709,N_36031,N_35507);
nand U37710 (N_37710,N_35558,N_36653);
nor U37711 (N_37711,N_36926,N_35961);
or U37712 (N_37712,N_36885,N_36130);
xor U37713 (N_37713,N_35792,N_36864);
xnor U37714 (N_37714,N_36913,N_36318);
xor U37715 (N_37715,N_35031,N_36727);
or U37716 (N_37716,N_36467,N_35302);
and U37717 (N_37717,N_37216,N_35796);
and U37718 (N_37718,N_36809,N_36070);
nand U37719 (N_37719,N_37339,N_36310);
and U37720 (N_37720,N_35105,N_36132);
or U37721 (N_37721,N_35037,N_35877);
and U37722 (N_37722,N_36215,N_36551);
nand U37723 (N_37723,N_37428,N_35790);
or U37724 (N_37724,N_35275,N_36780);
nor U37725 (N_37725,N_37078,N_35114);
xor U37726 (N_37726,N_36000,N_37119);
and U37727 (N_37727,N_37438,N_36049);
or U37728 (N_37728,N_36741,N_35789);
xnor U37729 (N_37729,N_35530,N_37161);
nor U37730 (N_37730,N_36059,N_35084);
nand U37731 (N_37731,N_36848,N_37211);
nor U37732 (N_37732,N_36222,N_35443);
or U37733 (N_37733,N_35181,N_36652);
nor U37734 (N_37734,N_36607,N_36960);
and U37735 (N_37735,N_35832,N_37048);
or U37736 (N_37736,N_35099,N_35287);
nor U37737 (N_37737,N_36221,N_37470);
nand U37738 (N_37738,N_35636,N_37217);
nand U37739 (N_37739,N_36686,N_35209);
nand U37740 (N_37740,N_36337,N_37396);
xor U37741 (N_37741,N_35174,N_36892);
or U37742 (N_37742,N_35429,N_35136);
or U37743 (N_37743,N_37484,N_37415);
and U37744 (N_37744,N_36731,N_36057);
xor U37745 (N_37745,N_35480,N_35273);
nor U37746 (N_37746,N_36090,N_36250);
xnor U37747 (N_37747,N_35664,N_35407);
or U37748 (N_37748,N_35670,N_36978);
and U37749 (N_37749,N_36783,N_35642);
or U37750 (N_37750,N_36257,N_35102);
or U37751 (N_37751,N_37055,N_35577);
xnor U37752 (N_37752,N_36439,N_36350);
or U37753 (N_37753,N_35246,N_35838);
nand U37754 (N_37754,N_36216,N_36694);
or U37755 (N_37755,N_37460,N_37225);
xnor U37756 (N_37756,N_36266,N_37429);
xor U37757 (N_37757,N_35552,N_35308);
nand U37758 (N_37758,N_37283,N_36412);
nor U37759 (N_37759,N_35184,N_36341);
nand U37760 (N_37760,N_36444,N_36634);
and U37761 (N_37761,N_37070,N_36940);
nor U37762 (N_37762,N_35315,N_35669);
nand U37763 (N_37763,N_35251,N_35500);
xnor U37764 (N_37764,N_36543,N_36516);
and U37765 (N_37765,N_36635,N_35247);
xor U37766 (N_37766,N_35061,N_36546);
and U37767 (N_37767,N_35219,N_35751);
and U37768 (N_37768,N_35348,N_35683);
nor U37769 (N_37769,N_36079,N_36392);
or U37770 (N_37770,N_36959,N_35504);
and U37771 (N_37771,N_36561,N_35780);
or U37772 (N_37772,N_35818,N_36277);
nand U37773 (N_37773,N_36207,N_36088);
xor U37774 (N_37774,N_36608,N_36270);
nand U37775 (N_37775,N_35512,N_36169);
or U37776 (N_37776,N_35985,N_36105);
nand U37777 (N_37777,N_35321,N_36769);
nor U37778 (N_37778,N_36120,N_35283);
nor U37779 (N_37779,N_37378,N_35781);
or U37780 (N_37780,N_37457,N_36585);
or U37781 (N_37781,N_35090,N_36284);
nand U37782 (N_37782,N_36505,N_36045);
nor U37783 (N_37783,N_36524,N_36336);
xnor U37784 (N_37784,N_37117,N_35096);
nand U37785 (N_37785,N_35365,N_35942);
xor U37786 (N_37786,N_37407,N_35816);
and U37787 (N_37787,N_37411,N_35261);
xor U37788 (N_37788,N_35187,N_36241);
or U37789 (N_37789,N_36770,N_36624);
nor U37790 (N_37790,N_35623,N_36547);
nor U37791 (N_37791,N_36512,N_36299);
or U37792 (N_37792,N_37237,N_36592);
nor U37793 (N_37793,N_37493,N_36499);
xnor U37794 (N_37794,N_35319,N_35956);
or U37795 (N_37795,N_36999,N_36200);
or U37796 (N_37796,N_36393,N_36620);
and U37797 (N_37797,N_36171,N_36776);
nor U37798 (N_37798,N_35593,N_36570);
xor U37799 (N_37799,N_36983,N_36420);
or U37800 (N_37800,N_36834,N_36311);
nand U37801 (N_37801,N_36519,N_37402);
nor U37802 (N_37802,N_36349,N_35645);
and U37803 (N_37803,N_37389,N_36232);
and U37804 (N_37804,N_35451,N_37215);
xnor U37805 (N_37805,N_36365,N_37185);
nand U37806 (N_37806,N_35284,N_35288);
nand U37807 (N_37807,N_37027,N_35083);
or U37808 (N_37808,N_36562,N_35240);
and U37809 (N_37809,N_35266,N_37175);
or U37810 (N_37810,N_37093,N_36986);
nand U37811 (N_37811,N_35700,N_36845);
nand U37812 (N_37812,N_37421,N_36465);
nor U37813 (N_37813,N_36583,N_35171);
and U37814 (N_37814,N_35124,N_36091);
or U37815 (N_37815,N_35012,N_36545);
nand U37816 (N_37816,N_37199,N_36775);
xnor U37817 (N_37817,N_36929,N_35690);
or U37818 (N_37818,N_37123,N_35449);
nand U37819 (N_37819,N_37454,N_36179);
and U37820 (N_37820,N_36854,N_35229);
xor U37821 (N_37821,N_36496,N_37288);
nor U37822 (N_37822,N_36843,N_36271);
xnor U37823 (N_37823,N_37035,N_35324);
xor U37824 (N_37824,N_36123,N_35650);
xnor U37825 (N_37825,N_35198,N_36136);
or U37826 (N_37826,N_37317,N_37005);
and U37827 (N_37827,N_37037,N_36719);
nor U37828 (N_37828,N_37372,N_35839);
or U37829 (N_37829,N_35915,N_37437);
and U37830 (N_37830,N_35982,N_36099);
xor U37831 (N_37831,N_35971,N_35470);
or U37832 (N_37832,N_35909,N_35765);
or U37833 (N_37833,N_35567,N_36463);
or U37834 (N_37834,N_35583,N_37202);
and U37835 (N_37835,N_35616,N_36288);
xor U37836 (N_37836,N_35329,N_35991);
xor U37837 (N_37837,N_35193,N_35723);
xnor U37838 (N_37838,N_35026,N_36961);
and U37839 (N_37839,N_36982,N_35456);
nand U37840 (N_37840,N_35070,N_35905);
xor U37841 (N_37841,N_35064,N_36797);
and U37842 (N_37842,N_36755,N_35783);
and U37843 (N_37843,N_37069,N_37463);
and U37844 (N_37844,N_36760,N_36357);
nor U37845 (N_37845,N_35737,N_36395);
nand U37846 (N_37846,N_36259,N_36703);
xnor U37847 (N_37847,N_35030,N_36489);
and U37848 (N_37848,N_36938,N_35939);
nor U37849 (N_37849,N_35570,N_35479);
or U37850 (N_37850,N_37383,N_35293);
and U37851 (N_37851,N_36399,N_35395);
and U37852 (N_37852,N_35937,N_36721);
xor U37853 (N_37853,N_35244,N_35505);
nor U37854 (N_37854,N_37371,N_36007);
nor U37855 (N_37855,N_36224,N_36124);
or U37856 (N_37856,N_35047,N_36865);
nor U37857 (N_37857,N_36613,N_35027);
xor U37858 (N_37858,N_36831,N_36144);
nand U37859 (N_37859,N_35630,N_36316);
and U37860 (N_37860,N_37480,N_37462);
nor U37861 (N_37861,N_35620,N_36909);
nor U37862 (N_37862,N_36738,N_36782);
nand U37863 (N_37863,N_35633,N_35182);
xor U37864 (N_37864,N_37138,N_37356);
nand U37865 (N_37865,N_36955,N_35117);
nor U37866 (N_37866,N_37250,N_36602);
nand U37867 (N_37867,N_35898,N_37375);
nor U37868 (N_37868,N_37129,N_36035);
nand U37869 (N_37869,N_36899,N_37032);
xnor U37870 (N_37870,N_35076,N_35605);
xnor U37871 (N_37871,N_36378,N_36540);
or U37872 (N_37872,N_35032,N_36248);
nor U37873 (N_37873,N_37475,N_35005);
or U37874 (N_37874,N_36344,N_37373);
nand U37875 (N_37875,N_35797,N_37364);
or U37876 (N_37876,N_36829,N_37218);
nor U37877 (N_37877,N_37063,N_37489);
nand U37878 (N_37878,N_35579,N_36690);
and U37879 (N_37879,N_36599,N_36508);
nand U37880 (N_37880,N_36438,N_36657);
xnor U37881 (N_37881,N_35004,N_35358);
nor U37882 (N_37882,N_35122,N_35465);
or U37883 (N_37883,N_36364,N_37255);
nor U37884 (N_37884,N_36472,N_35374);
or U37885 (N_37885,N_36704,N_35250);
nor U37886 (N_37886,N_35370,N_35748);
xor U37887 (N_37887,N_37380,N_35773);
nor U37888 (N_37888,N_35540,N_37350);
xor U37889 (N_37889,N_36107,N_36138);
and U37890 (N_37890,N_36158,N_35499);
nor U37891 (N_37891,N_36033,N_35802);
nor U37892 (N_37892,N_35930,N_36837);
and U37893 (N_37893,N_36071,N_37425);
xor U37894 (N_37894,N_35594,N_37114);
nor U37895 (N_37895,N_36844,N_37086);
and U37896 (N_37896,N_35168,N_35152);
or U37897 (N_37897,N_35088,N_35191);
and U37898 (N_37898,N_36203,N_36457);
xnor U37899 (N_37899,N_36577,N_37209);
nor U37900 (N_37900,N_37174,N_36073);
or U37901 (N_37901,N_35921,N_37491);
or U37902 (N_37902,N_36711,N_35011);
or U37903 (N_37903,N_36354,N_35446);
nand U37904 (N_37904,N_37235,N_36324);
nand U37905 (N_37905,N_36581,N_35019);
nor U37906 (N_37906,N_36249,N_37286);
nor U37907 (N_37907,N_36408,N_35671);
nand U37908 (N_37908,N_35042,N_37333);
xnor U37909 (N_37909,N_35842,N_36166);
xor U37910 (N_37910,N_37224,N_35800);
and U37911 (N_37911,N_36480,N_35025);
or U37912 (N_37912,N_35320,N_35933);
nor U37913 (N_37913,N_35458,N_35613);
nor U37914 (N_37914,N_37451,N_35220);
xnor U37915 (N_37915,N_36135,N_35183);
xor U37916 (N_37916,N_35599,N_36098);
and U37917 (N_37917,N_36722,N_35834);
nand U37918 (N_37918,N_36347,N_36793);
nor U37919 (N_37919,N_35859,N_36676);
nand U37920 (N_37920,N_35337,N_35836);
and U37921 (N_37921,N_35676,N_36900);
xnor U37922 (N_37922,N_36133,N_36458);
nand U37923 (N_37923,N_36100,N_36112);
or U37924 (N_37924,N_36093,N_35227);
nor U37925 (N_37925,N_35953,N_36970);
xor U37926 (N_37926,N_37169,N_35711);
and U37927 (N_37927,N_36669,N_37068);
nor U37928 (N_37928,N_37304,N_36919);
and U37929 (N_37929,N_36725,N_35303);
nand U37930 (N_37930,N_36114,N_35014);
or U37931 (N_37931,N_35634,N_35006);
or U37932 (N_37932,N_36193,N_35994);
xor U37933 (N_37933,N_37431,N_36696);
and U37934 (N_37934,N_36184,N_35085);
nor U37935 (N_37935,N_36312,N_36963);
nand U37936 (N_37936,N_35245,N_35492);
xor U37937 (N_37937,N_35785,N_35844);
nand U37938 (N_37938,N_36542,N_36717);
and U37939 (N_37939,N_36297,N_35554);
or U37940 (N_37940,N_37444,N_35141);
nor U37941 (N_37941,N_35769,N_35641);
nand U37942 (N_37942,N_37142,N_37326);
nand U37943 (N_37943,N_37003,N_35699);
xor U37944 (N_37944,N_37296,N_35474);
nand U37945 (N_37945,N_36016,N_36827);
nor U37946 (N_37946,N_36858,N_35696);
nand U37947 (N_37947,N_36897,N_37499);
nand U37948 (N_37948,N_36234,N_37097);
nor U37949 (N_37949,N_36951,N_35388);
xnor U37950 (N_37950,N_36307,N_35535);
nand U37951 (N_37951,N_36296,N_37247);
nand U37952 (N_37952,N_37239,N_37053);
nor U37953 (N_37953,N_36957,N_35074);
xnor U37954 (N_37954,N_37021,N_35768);
xor U37955 (N_37955,N_35411,N_36125);
nor U37956 (N_37956,N_35922,N_35536);
or U37957 (N_37957,N_35139,N_37434);
xor U37958 (N_37958,N_36466,N_35351);
and U37959 (N_37959,N_35565,N_35656);
xnor U37960 (N_37960,N_35925,N_37292);
or U37961 (N_37961,N_35561,N_36424);
xnor U37962 (N_37962,N_35353,N_37422);
and U37963 (N_37963,N_36202,N_37343);
and U37964 (N_37964,N_36747,N_35945);
xnor U37965 (N_37965,N_36836,N_35709);
or U37966 (N_37966,N_36530,N_35648);
nand U37967 (N_37967,N_36014,N_36106);
nand U37968 (N_37968,N_36718,N_35519);
and U37969 (N_37969,N_35525,N_36411);
nand U37970 (N_37970,N_36385,N_35845);
or U37971 (N_37971,N_36695,N_36633);
nor U37972 (N_37972,N_36688,N_37297);
xor U37973 (N_37973,N_37345,N_36327);
nand U37974 (N_37974,N_35402,N_36058);
nand U37975 (N_37975,N_35852,N_37040);
xnor U37976 (N_37976,N_35580,N_36989);
nor U37977 (N_37977,N_36687,N_35147);
xor U37978 (N_37978,N_36377,N_35401);
or U37979 (N_37979,N_36060,N_35471);
nand U37980 (N_37980,N_36862,N_36080);
nand U37981 (N_37981,N_36161,N_35013);
nand U37982 (N_37982,N_35502,N_36692);
and U37983 (N_37983,N_36194,N_36418);
and U37984 (N_37984,N_35095,N_36677);
nand U37985 (N_37985,N_36766,N_35914);
nand U37986 (N_37986,N_37360,N_37398);
or U37987 (N_37987,N_35189,N_36964);
nand U37988 (N_37988,N_36278,N_36952);
or U37989 (N_37989,N_37245,N_36426);
nor U37990 (N_37990,N_35529,N_36500);
and U37991 (N_37991,N_36352,N_37039);
xnor U37992 (N_37992,N_37153,N_36839);
or U37993 (N_37993,N_35887,N_36367);
nor U37994 (N_37994,N_35899,N_36628);
xnor U37995 (N_37995,N_35063,N_35089);
xor U37996 (N_37996,N_37464,N_36305);
or U37997 (N_37997,N_36208,N_36729);
xnor U37998 (N_37998,N_36409,N_35977);
and U37999 (N_37999,N_35589,N_37353);
and U38000 (N_38000,N_35267,N_36018);
nor U38001 (N_38001,N_36491,N_37030);
and U38002 (N_38002,N_35998,N_35840);
or U38003 (N_38003,N_35258,N_36462);
xor U38004 (N_38004,N_35705,N_36174);
or U38005 (N_38005,N_36103,N_35002);
or U38006 (N_38006,N_36621,N_36498);
nor U38007 (N_38007,N_37015,N_37369);
nand U38008 (N_38008,N_35908,N_37394);
nand U38009 (N_38009,N_36924,N_35947);
xnor U38010 (N_38010,N_35771,N_36469);
xnor U38011 (N_38011,N_37124,N_36137);
nand U38012 (N_38012,N_37406,N_35523);
nand U38013 (N_38013,N_37004,N_35144);
nor U38014 (N_38014,N_35482,N_36786);
nand U38015 (N_38015,N_37439,N_36714);
nand U38016 (N_38016,N_35384,N_36274);
xor U38017 (N_38017,N_36896,N_35336);
xnor U38018 (N_38018,N_36507,N_37074);
xnor U38019 (N_38019,N_37089,N_35242);
nor U38020 (N_38020,N_35175,N_36047);
xor U38021 (N_38021,N_36209,N_35680);
nor U38022 (N_38022,N_37266,N_36889);
and U38023 (N_38023,N_37344,N_36802);
and U38024 (N_38024,N_35188,N_35417);
nor U38025 (N_38025,N_36373,N_37414);
and U38026 (N_38026,N_36474,N_35886);
nor U38027 (N_38027,N_36484,N_36949);
or U38028 (N_38028,N_35051,N_37012);
and U38029 (N_38029,N_36656,N_35204);
xnor U38030 (N_38030,N_37386,N_36981);
nor U38031 (N_38031,N_35381,N_35882);
nand U38032 (N_38032,N_35444,N_37337);
nand U38033 (N_38033,N_35462,N_37293);
or U38034 (N_38034,N_36191,N_35058);
and U38035 (N_38035,N_36064,N_35959);
xnor U38036 (N_38036,N_35710,N_35112);
and U38037 (N_38037,N_36732,N_36082);
nor U38038 (N_38038,N_37212,N_37387);
nand U38039 (N_38039,N_36332,N_35919);
or U38040 (N_38040,N_35776,N_35753);
nand U38041 (N_38041,N_36383,N_35538);
nand U38042 (N_38042,N_37195,N_36558);
nand U38043 (N_38043,N_35215,N_37450);
xor U38044 (N_38044,N_37182,N_35317);
or U38045 (N_38045,N_35081,N_36754);
nand U38046 (N_38046,N_35895,N_36010);
xnor U38047 (N_38047,N_37391,N_35651);
or U38048 (N_38048,N_35062,N_35103);
nor U38049 (N_38049,N_37382,N_35878);
xor U38050 (N_38050,N_36555,N_36430);
nand U38051 (N_38051,N_35604,N_37270);
nor U38052 (N_38052,N_35406,N_37099);
nand U38053 (N_38053,N_36771,N_35679);
and U38054 (N_38054,N_37177,N_36131);
and U38055 (N_38055,N_35367,N_37248);
nand U38056 (N_38056,N_36943,N_36789);
and U38057 (N_38057,N_35752,N_36143);
xnor U38058 (N_38058,N_37347,N_37260);
xnor U38059 (N_38059,N_37154,N_37051);
xor U38060 (N_38060,N_35975,N_35371);
or U38061 (N_38061,N_36116,N_36325);
nand U38062 (N_38062,N_36744,N_36441);
and U38063 (N_38063,N_36417,N_36206);
or U38064 (N_38064,N_35260,N_35420);
nor U38065 (N_38065,N_37165,N_37424);
or U38066 (N_38066,N_36340,N_36842);
nand U38067 (N_38067,N_35186,N_36991);
and U38068 (N_38068,N_35356,N_35390);
or U38069 (N_38069,N_37385,N_35207);
nor U38070 (N_38070,N_37107,N_37223);
or U38071 (N_38071,N_35409,N_36730);
nor U38072 (N_38072,N_37271,N_35903);
nor U38073 (N_38073,N_35995,N_37302);
or U38074 (N_38074,N_36734,N_36847);
nor U38075 (N_38075,N_35957,N_37363);
xnor U38076 (N_38076,N_37116,N_35657);
or U38077 (N_38077,N_36749,N_37062);
and U38078 (N_38078,N_35232,N_37445);
nand U38079 (N_38079,N_36493,N_35698);
or U38080 (N_38080,N_36345,N_35255);
xor U38081 (N_38081,N_37495,N_36196);
and U38082 (N_38082,N_37052,N_36044);
xnor U38083 (N_38083,N_37112,N_35311);
nor U38084 (N_38084,N_36487,N_35376);
nand U38085 (N_38085,N_35758,N_35243);
and U38086 (N_38086,N_36947,N_36956);
nor U38087 (N_38087,N_35009,N_35224);
nor U38088 (N_38088,N_36173,N_36587);
nand U38089 (N_38089,N_35233,N_35161);
nand U38090 (N_38090,N_35573,N_35929);
nand U38091 (N_38091,N_36360,N_37214);
and U38092 (N_38092,N_37320,N_37115);
nor U38093 (N_38093,N_36920,N_36141);
and U38094 (N_38094,N_36918,N_35986);
or U38095 (N_38095,N_35459,N_35938);
or U38096 (N_38096,N_35559,N_35996);
nor U38097 (N_38097,N_36492,N_35637);
nand U38098 (N_38098,N_35383,N_35454);
nand U38099 (N_38099,N_37334,N_36870);
xor U38100 (N_38100,N_36353,N_36910);
xor U38101 (N_38101,N_37014,N_36097);
or U38102 (N_38102,N_35725,N_35412);
and U38103 (N_38103,N_37307,N_35917);
or U38104 (N_38104,N_35891,N_35719);
nor U38105 (N_38105,N_36261,N_35546);
nand U38106 (N_38106,N_36654,N_35927);
xnor U38107 (N_38107,N_37152,N_35872);
nor U38108 (N_38108,N_36362,N_35431);
nand U38109 (N_38109,N_36976,N_36898);
nor U38110 (N_38110,N_36154,N_35588);
and U38111 (N_38111,N_36156,N_35704);
nand U38112 (N_38112,N_35726,N_35392);
nor U38113 (N_38113,N_35216,N_36813);
nand U38114 (N_38114,N_36743,N_36939);
and U38115 (N_38115,N_36753,N_37028);
nand U38116 (N_38116,N_35866,N_35098);
or U38117 (N_38117,N_36488,N_36197);
nand U38118 (N_38118,N_35993,N_35562);
nand U38119 (N_38119,N_36256,N_36092);
xor U38120 (N_38120,N_36052,N_36713);
or U38121 (N_38121,N_37130,N_37284);
xnor U38122 (N_38122,N_37413,N_36391);
and U38123 (N_38123,N_36569,N_36269);
or U38124 (N_38124,N_36019,N_37264);
or U38125 (N_38125,N_35195,N_35071);
or U38126 (N_38126,N_37453,N_35307);
and U38127 (N_38127,N_36181,N_35980);
nand U38128 (N_38128,N_36996,N_35865);
nor U38129 (N_38129,N_37064,N_37100);
xor U38130 (N_38130,N_37184,N_35279);
or U38131 (N_38131,N_35506,N_36078);
xor U38132 (N_38132,N_35387,N_35165);
or U38133 (N_38133,N_36830,N_36151);
or U38134 (N_38134,N_35574,N_37262);
and U38135 (N_38135,N_37170,N_37018);
nand U38136 (N_38136,N_35598,N_36534);
xor U38137 (N_38137,N_36851,N_35885);
nor U38138 (N_38138,N_35143,N_37351);
xnor U38139 (N_38139,N_35177,N_37497);
or U38140 (N_38140,N_37017,N_36129);
or U38141 (N_38141,N_36013,N_37455);
and U38142 (N_38142,N_35739,N_37049);
xor U38143 (N_38143,N_35849,N_37252);
nor U38144 (N_38144,N_37420,N_35349);
xnor U38145 (N_38145,N_37256,N_35359);
nor U38146 (N_38146,N_35231,N_36882);
and U38147 (N_38147,N_35791,N_36658);
nand U38148 (N_38148,N_35173,N_35596);
or U38149 (N_38149,N_37275,N_36319);
and U38150 (N_38150,N_37409,N_36623);
xnor U38151 (N_38151,N_35113,N_36720);
nor U38152 (N_38152,N_36240,N_36405);
nand U38153 (N_38153,N_37399,N_36029);
nand U38154 (N_38154,N_36283,N_35675);
or U38155 (N_38155,N_36176,N_35786);
or U38156 (N_38156,N_36074,N_36142);
nor U38157 (N_38157,N_36069,N_36264);
nand U38158 (N_38158,N_36723,N_35867);
nor U38159 (N_38159,N_35992,N_35890);
nor U38160 (N_38160,N_36591,N_37222);
and U38161 (N_38161,N_35823,N_36372);
nand U38162 (N_38162,N_35817,N_36066);
nor U38163 (N_38163,N_35230,N_36165);
nand U38164 (N_38164,N_35547,N_35793);
or U38165 (N_38165,N_36291,N_37427);
and U38166 (N_38166,N_35974,N_35847);
or U38167 (N_38167,N_35894,N_35875);
nand U38168 (N_38168,N_36262,N_36901);
nor U38169 (N_38169,N_35208,N_36678);
and U38170 (N_38170,N_36659,N_36932);
nor U38171 (N_38171,N_36933,N_35884);
or U38172 (N_38172,N_37294,N_37045);
nor U38173 (N_38173,N_35488,N_37323);
and U38174 (N_38174,N_35126,N_35837);
nor U38175 (N_38175,N_36707,N_36712);
and U38176 (N_38176,N_36663,N_37022);
nor U38177 (N_38177,N_35352,N_36803);
and U38178 (N_38178,N_35052,N_36575);
nand U38179 (N_38179,N_35397,N_36231);
nand U38180 (N_38180,N_35795,N_35868);
and U38181 (N_38181,N_37366,N_35833);
xor U38182 (N_38182,N_37023,N_35464);
nor U38183 (N_38183,N_36388,N_36544);
xor U38184 (N_38184,N_36536,N_37071);
nor U38185 (N_38185,N_36517,N_35988);
and U38186 (N_38186,N_35772,N_35121);
and U38187 (N_38187,N_35249,N_37091);
or U38188 (N_38188,N_37066,N_35379);
and U38189 (N_38189,N_37487,N_36201);
xor U38190 (N_38190,N_35271,N_35624);
or U38191 (N_38191,N_36759,N_35225);
or U38192 (N_38192,N_36389,N_35130);
and U38193 (N_38193,N_35340,N_36852);
xnor U38194 (N_38194,N_35557,N_36315);
xnor U38195 (N_38195,N_36244,N_36008);
nand U38196 (N_38196,N_35325,N_35862);
xor U38197 (N_38197,N_36293,N_36323);
nor U38198 (N_38198,N_37405,N_35652);
xnor U38199 (N_38199,N_36442,N_36229);
and U38200 (N_38200,N_37101,N_36384);
and U38201 (N_38201,N_36661,N_35427);
nand U38202 (N_38202,N_36994,N_36246);
nand U38203 (N_38203,N_36627,N_35414);
or U38204 (N_38204,N_36427,N_37230);
and U38205 (N_38205,N_37166,N_35960);
nand U38206 (N_38206,N_36974,N_36302);
nor U38207 (N_38207,N_36056,N_36227);
or U38208 (N_38208,N_35731,N_35022);
nand U38209 (N_38209,N_35732,N_35119);
nand U38210 (N_38210,N_35759,N_36067);
nor U38211 (N_38211,N_36529,N_36170);
nand U38212 (N_38212,N_36806,N_35578);
and U38213 (N_38213,N_35774,N_37113);
or U38214 (N_38214,N_36706,N_37298);
or U38215 (N_38215,N_36102,N_36610);
nand U38216 (N_38216,N_36556,N_36643);
nand U38217 (N_38217,N_35093,N_37426);
and U38218 (N_38218,N_36828,N_36485);
or U38219 (N_38219,N_36616,N_35203);
xnor U38220 (N_38220,N_36021,N_36027);
or U38221 (N_38221,N_36394,N_35591);
and U38222 (N_38222,N_35060,N_36189);
nand U38223 (N_38223,N_37436,N_35438);
nor U38224 (N_38224,N_35439,N_37083);
or U38225 (N_38225,N_35469,N_37204);
nor U38226 (N_38226,N_36579,N_37370);
or U38227 (N_38227,N_36113,N_35870);
nand U38228 (N_38228,N_36800,N_35714);
nor U38229 (N_38229,N_35024,N_36460);
xor U38230 (N_38230,N_36642,N_35799);
or U38231 (N_38231,N_35077,N_35685);
nor U38232 (N_38232,N_35738,N_35263);
nand U38233 (N_38233,N_36401,N_36810);
nor U38234 (N_38234,N_36905,N_36238);
or U38235 (N_38235,N_36515,N_35493);
xnor U38236 (N_38236,N_35963,N_36111);
nand U38237 (N_38237,N_35468,N_37261);
and U38238 (N_38238,N_37206,N_35912);
or U38239 (N_38239,N_35007,N_35094);
or U38240 (N_38240,N_35569,N_36866);
nand U38241 (N_38241,N_36509,N_36397);
xor U38242 (N_38242,N_36644,N_36304);
nand U38243 (N_38243,N_37430,N_37471);
or U38244 (N_38244,N_36043,N_36647);
xor U38245 (N_38245,N_35347,N_35706);
nor U38246 (N_38246,N_35115,N_36564);
nor U38247 (N_38247,N_37110,N_35848);
or U38248 (N_38248,N_36083,N_35741);
and U38249 (N_38249,N_36667,N_36038);
or U38250 (N_38250,N_35560,N_35972);
or U38251 (N_38251,N_35924,N_36279);
xnor U38252 (N_38252,N_37188,N_36513);
and U38253 (N_38253,N_36055,N_35179);
nor U38254 (N_38254,N_35528,N_36317);
nand U38255 (N_38255,N_35495,N_37465);
and U38256 (N_38256,N_36346,N_37340);
and U38257 (N_38257,N_35380,N_36580);
or U38258 (N_38258,N_36446,N_35043);
and U38259 (N_38259,N_35970,N_36182);
and U38260 (N_38260,N_35518,N_37236);
and U38261 (N_38261,N_37238,N_35733);
xnor U38262 (N_38262,N_35692,N_36118);
or U38263 (N_38263,N_37384,N_36664);
and U38264 (N_38264,N_36637,N_36379);
nand U38265 (N_38265,N_36902,N_36413);
or U38266 (N_38266,N_35257,N_37024);
nor U38267 (N_38267,N_36087,N_35517);
xnor U38268 (N_38268,N_37011,N_36146);
xor U38269 (N_38269,N_36765,N_37441);
nor U38270 (N_38270,N_36255,N_35433);
and U38271 (N_38271,N_35718,N_35029);
xor U38272 (N_38272,N_35286,N_36252);
nand U38273 (N_38273,N_36272,N_36946);
nand U38274 (N_38274,N_36081,N_36518);
or U38275 (N_38275,N_36433,N_36039);
nor U38276 (N_38276,N_36110,N_36198);
nor U38277 (N_38277,N_36321,N_37061);
nand U38278 (N_38278,N_37244,N_37448);
nand U38279 (N_38279,N_36872,N_35747);
and U38280 (N_38280,N_36737,N_35697);
xor U38281 (N_38281,N_35087,N_35609);
nand U38282 (N_38282,N_36971,N_35306);
nand U38283 (N_38283,N_35343,N_35125);
nand U38284 (N_38284,N_37139,N_35339);
nand U38285 (N_38285,N_36915,N_35408);
nor U38286 (N_38286,N_35539,N_35237);
and U38287 (N_38287,N_35851,N_37459);
xor U38288 (N_38288,N_36931,N_36675);
xor U38289 (N_38289,N_35603,N_37085);
or U38290 (N_38290,N_36015,N_37033);
or U38291 (N_38291,N_36740,N_36009);
xor U38292 (N_38292,N_35153,N_37219);
nor U38293 (N_38293,N_35531,N_36923);
or U38294 (N_38294,N_35269,N_35566);
nor U38295 (N_38295,N_36767,N_35809);
and U38296 (N_38296,N_36541,N_36449);
or U38297 (N_38297,N_37362,N_36606);
or U38298 (N_38298,N_36816,N_35513);
nand U38299 (N_38299,N_35369,N_36973);
nor U38300 (N_38300,N_35923,N_35522);
xnor U38301 (N_38301,N_37026,N_35555);
nand U38302 (N_38302,N_35146,N_36857);
nand U38303 (N_38303,N_35607,N_35268);
nor U38304 (N_38304,N_36930,N_35394);
xor U38305 (N_38305,N_37102,N_37276);
or U38306 (N_38306,N_37134,N_35515);
or U38307 (N_38307,N_35050,N_36121);
or U38308 (N_38308,N_36861,N_37327);
nand U38309 (N_38309,N_36101,N_36506);
and U38310 (N_38310,N_36012,N_37349);
xnor U38311 (N_38311,N_35521,N_35041);
xnor U38312 (N_38312,N_35511,N_36177);
nor U38313 (N_38313,N_36625,N_36195);
nor U38314 (N_38314,N_36180,N_35928);
nand U38315 (N_38315,N_35463,N_35131);
nor U38316 (N_38316,N_37278,N_36239);
nand U38317 (N_38317,N_37309,N_36600);
xor U38318 (N_38318,N_36927,N_35496);
and U38319 (N_38319,N_37240,N_37316);
and U38320 (N_38320,N_35375,N_35935);
nor U38321 (N_38321,N_36375,N_37200);
and U38322 (N_38322,N_37357,N_36450);
nor U38323 (N_38323,N_37306,N_37127);
nor U38324 (N_38324,N_35148,N_37330);
or U38325 (N_38325,N_36903,N_35331);
or U38326 (N_38326,N_35045,N_35501);
xor U38327 (N_38327,N_35717,N_37143);
and U38328 (N_38328,N_37432,N_35154);
and U38329 (N_38329,N_36011,N_35097);
or U38330 (N_38330,N_35808,N_35889);
xnor U38331 (N_38331,N_35092,N_35079);
and U38332 (N_38332,N_36109,N_36619);
xnor U38333 (N_38333,N_37073,N_36728);
xor U38334 (N_38334,N_36567,N_35542);
and U38335 (N_38335,N_35354,N_35524);
xor U38336 (N_38336,N_35729,N_37197);
nor U38337 (N_38337,N_35016,N_37160);
nor U38338 (N_38338,N_37125,N_36792);
nand U38339 (N_38339,N_36668,N_36374);
xnor U38340 (N_38340,N_35964,N_35180);
nor U38341 (N_38341,N_35803,N_37401);
and U38342 (N_38342,N_35775,N_36217);
nor U38343 (N_38343,N_35640,N_35621);
and U38344 (N_38344,N_35341,N_35987);
xnor U38345 (N_38345,N_35989,N_36108);
xnor U38346 (N_38346,N_35176,N_36724);
or U38347 (N_38347,N_36841,N_35366);
and U38348 (N_38348,N_37067,N_36550);
or U38349 (N_38349,N_37038,N_36376);
or U38350 (N_38350,N_36421,N_37172);
and U38351 (N_38351,N_35597,N_36726);
nor U38352 (N_38352,N_36282,N_36904);
and U38353 (N_38353,N_36292,N_36648);
or U38354 (N_38354,N_37329,N_35858);
nand U38355 (N_38355,N_36936,N_35386);
and U38356 (N_38356,N_37315,N_37150);
or U38357 (N_38357,N_37410,N_35476);
and U38358 (N_38358,N_37417,N_36178);
and U38359 (N_38359,N_37120,N_35586);
and U38360 (N_38360,N_37328,N_35708);
or U38361 (N_38361,N_36944,N_36210);
nand U38362 (N_38362,N_36086,N_36343);
nand U38363 (N_38363,N_36632,N_35695);
and U38364 (N_38364,N_36308,N_35276);
nor U38365 (N_38365,N_36990,N_36245);
xnor U38366 (N_38366,N_37106,N_37082);
or U38367 (N_38367,N_37034,N_35344);
nor U38368 (N_38368,N_37443,N_37440);
xnor U38369 (N_38369,N_37474,N_37233);
and U38370 (N_38370,N_36911,N_35684);
xor U38371 (N_38371,N_35040,N_35981);
nand U38372 (N_38372,N_36358,N_35104);
nor U38373 (N_38373,N_35067,N_36948);
nor U38374 (N_38374,N_35065,N_36790);
or U38375 (N_38375,N_37137,N_36320);
nand U38376 (N_38376,N_36636,N_36247);
nand U38377 (N_38377,N_37060,N_36490);
xor U38378 (N_38378,N_36805,N_35826);
or U38379 (N_38379,N_37282,N_37408);
nor U38380 (N_38380,N_37281,N_35034);
nand U38381 (N_38381,N_36812,N_35762);
or U38382 (N_38382,N_35755,N_37301);
nand U38383 (N_38383,N_37352,N_36204);
and U38384 (N_38384,N_37251,N_36867);
and U38385 (N_38385,N_35804,N_35421);
or U38386 (N_38386,N_36945,N_36975);
nand U38387 (N_38387,N_36883,N_37077);
xnor U38388 (N_38388,N_36820,N_37176);
and U38389 (N_38389,N_36356,N_36850);
nand U38390 (N_38390,N_36791,N_36596);
xor U38391 (N_38391,N_35132,N_36396);
nand U38392 (N_38392,N_36804,N_37231);
or U38393 (N_38393,N_36398,N_36422);
or U38394 (N_38394,N_36423,N_35672);
xor U38395 (N_38395,N_37140,N_37131);
or U38396 (N_38396,N_35159,N_36459);
xor U38397 (N_38397,N_35678,N_36298);
and U38398 (N_38398,N_37390,N_36175);
and U38399 (N_38399,N_36745,N_36258);
nor U38400 (N_38400,N_35541,N_36521);
xnor U38401 (N_38401,N_37258,N_36895);
nor U38402 (N_38402,N_37072,N_37029);
nor U38403 (N_38403,N_35158,N_37257);
or U38404 (N_38404,N_35140,N_35900);
and U38405 (N_38405,N_36742,N_37227);
xor U38406 (N_38406,N_36748,N_35815);
and U38407 (N_38407,N_37076,N_35053);
nand U38408 (N_38408,N_36552,N_36701);
or U38409 (N_38409,N_36437,N_36287);
or U38410 (N_38410,N_35893,N_36815);
and U38411 (N_38411,N_35452,N_35694);
xnor U38412 (N_38412,N_36290,N_36425);
and U38413 (N_38413,N_35687,N_36028);
nand U38414 (N_38414,N_36548,N_35491);
or U38415 (N_38415,N_37059,N_35835);
xor U38416 (N_38416,N_36199,N_36761);
and U38417 (N_38417,N_35330,N_35297);
xor U38418 (N_38418,N_37268,N_37156);
nand U38419 (N_38419,N_37295,N_37178);
or U38420 (N_38420,N_37079,N_35854);
or U38421 (N_38421,N_37065,N_35976);
or U38422 (N_38422,N_35806,N_35015);
and U38423 (N_38423,N_36140,N_35665);
and U38424 (N_38424,N_35807,N_35958);
nand U38425 (N_38425,N_37002,N_36925);
xor U38426 (N_38426,N_36301,N_36068);
nand U38427 (N_38427,N_36369,N_35897);
or U38428 (N_38428,N_35904,N_36818);
xor U38429 (N_38429,N_37458,N_36190);
xor U38430 (N_38430,N_36611,N_37104);
nor U38431 (N_38431,N_35563,N_35787);
xor U38432 (N_38432,N_35572,N_35264);
and U38433 (N_38433,N_36962,N_36594);
nor U38434 (N_38434,N_35677,N_35999);
or U38435 (N_38435,N_36479,N_35721);
nand U38436 (N_38436,N_36464,N_37168);
or U38437 (N_38437,N_36520,N_35192);
or U38438 (N_38438,N_36777,N_35805);
nor U38439 (N_38439,N_35940,N_36684);
nand U38440 (N_38440,N_36163,N_37006);
or U38441 (N_38441,N_37081,N_35425);
nor U38442 (N_38442,N_37163,N_35296);
nand U38443 (N_38443,N_35965,N_35239);
and U38444 (N_38444,N_36314,N_36708);
nor U38445 (N_38445,N_36236,N_35278);
or U38446 (N_38446,N_35856,N_35564);
or U38447 (N_38447,N_37145,N_37435);
or U38448 (N_38448,N_37277,N_35333);
or U38449 (N_38449,N_37167,N_35846);
and U38450 (N_38450,N_36478,N_36788);
and U38451 (N_38451,N_37058,N_36380);
xnor U38452 (N_38452,N_35646,N_35689);
xnor U38453 (N_38453,N_37090,N_37036);
nand U38454 (N_38454,N_37285,N_36557);
nor U38455 (N_38455,N_35473,N_36560);
nand U38456 (N_38456,N_37180,N_36468);
and U38457 (N_38457,N_35197,N_36185);
and U38458 (N_38458,N_36814,N_35635);
or U38459 (N_38459,N_36525,N_36819);
xor U38460 (N_38460,N_36455,N_35338);
and U38461 (N_38461,N_35328,N_35617);
nor U38462 (N_38462,N_36148,N_35843);
xor U38463 (N_38463,N_36921,N_35612);
nor U38464 (N_38464,N_35199,N_36077);
and U38465 (N_38465,N_36476,N_35304);
or U38466 (N_38466,N_35155,N_35049);
and U38467 (N_38467,N_35282,N_35357);
or U38468 (N_38468,N_35810,N_35202);
nand U38469 (N_38469,N_35978,N_37319);
nand U38470 (N_38470,N_36967,N_36447);
nand U38471 (N_38471,N_35322,N_36096);
xnor U38472 (N_38472,N_37483,N_35010);
nor U38473 (N_38473,N_36574,N_35760);
nor U38474 (N_38474,N_35223,N_35472);
nand U38475 (N_38475,N_35265,N_36470);
nand U38476 (N_38476,N_36906,N_36410);
xnor U38477 (N_38477,N_36494,N_36431);
nand U38478 (N_38478,N_35549,N_35537);
nor U38479 (N_38479,N_36988,N_37280);
nand U38480 (N_38480,N_36582,N_36679);
nor U38481 (N_38481,N_37007,N_37482);
xor U38482 (N_38482,N_35018,N_37321);
and U38483 (N_38483,N_35039,N_35763);
nand U38484 (N_38484,N_37241,N_35647);
nand U38485 (N_38485,N_37478,N_36638);
nand U38486 (N_38486,N_36334,N_37042);
and U38487 (N_38487,N_35326,N_36739);
or U38488 (N_38488,N_35316,N_35811);
nor U38489 (N_38489,N_36075,N_37242);
nand U38490 (N_38490,N_36758,N_35750);
or U38491 (N_38491,N_36750,N_35955);
nor U38492 (N_38492,N_35106,N_36522);
or U38493 (N_38493,N_37472,N_35481);
nor U38494 (N_38494,N_35160,N_35107);
nor U38495 (N_38495,N_35003,N_37016);
nand U38496 (N_38496,N_35662,N_35272);
or U38497 (N_38497,N_35066,N_36840);
xor U38498 (N_38498,N_35814,N_36061);
nand U38499 (N_38499,N_35614,N_35798);
or U38500 (N_38500,N_35682,N_35382);
xor U38501 (N_38501,N_36823,N_37159);
or U38502 (N_38502,N_37146,N_35461);
nand U38503 (N_38503,N_35876,N_36626);
nor U38504 (N_38504,N_37147,N_35078);
xor U38505 (N_38505,N_35073,N_36954);
or U38506 (N_38506,N_35133,N_36511);
nor U38507 (N_38507,N_35510,N_36331);
xor U38508 (N_38508,N_35135,N_36183);
nand U38509 (N_38509,N_36768,N_36950);
and U38510 (N_38510,N_35673,N_36046);
or U38511 (N_38511,N_35592,N_36072);
and U38512 (N_38512,N_35309,N_35754);
xor U38513 (N_38513,N_35571,N_35503);
and U38514 (N_38514,N_36275,N_36159);
and U38515 (N_38515,N_36764,N_35259);
or U38516 (N_38516,N_37132,N_37008);
or U38517 (N_38517,N_36604,N_35716);
or U38518 (N_38518,N_36036,N_36188);
nor U38519 (N_38519,N_36471,N_36001);
nor U38520 (N_38520,N_35545,N_37446);
nor U38521 (N_38521,N_35129,N_36601);
nor U38522 (N_38522,N_35206,N_36211);
nand U38523 (N_38523,N_36807,N_36859);
xnor U38524 (N_38524,N_35595,N_37311);
xor U38525 (N_38525,N_35713,N_35520);
nand U38526 (N_38526,N_35968,N_35788);
nand U38527 (N_38527,N_35643,N_35436);
nand U38528 (N_38528,N_35334,N_35497);
and U38529 (N_38529,N_35300,N_37025);
nor U38530 (N_38530,N_36415,N_35871);
nand U38531 (N_38531,N_35628,N_36309);
or U38532 (N_38532,N_36980,N_36691);
nand U38533 (N_38533,N_36335,N_36065);
and U38534 (N_38534,N_36095,N_36139);
nand U38535 (N_38535,N_37259,N_37332);
xor U38536 (N_38536,N_36860,N_36762);
xnor U38537 (N_38537,N_35949,N_36985);
and U38538 (N_38538,N_35779,N_35879);
and U38539 (N_38539,N_35766,N_36226);
and U38540 (N_38540,N_36881,N_35021);
xnor U38541 (N_38541,N_35028,N_35403);
xor U38542 (N_38542,N_35391,N_36683);
or U38543 (N_38543,N_35432,N_36366);
xnor U38544 (N_38544,N_36359,N_36670);
xor U38545 (N_38545,N_36794,N_36149);
nor U38546 (N_38546,N_37494,N_36890);
nor U38547 (N_38547,N_36863,N_35164);
or U38548 (N_38548,N_36003,N_36155);
and U38549 (N_38549,N_35742,N_35318);
xnor U38550 (N_38550,N_36281,N_35926);
or U38551 (N_38551,N_37210,N_36032);
nand U38552 (N_38552,N_35400,N_36554);
xnor U38553 (N_38553,N_36984,N_35057);
xnor U38554 (N_38554,N_35487,N_36527);
nand U38555 (N_38555,N_35368,N_37226);
nor U38556 (N_38556,N_35455,N_35361);
xor U38557 (N_38557,N_36254,N_37341);
nor U38558 (N_38558,N_36935,N_36796);
nor U38559 (N_38559,N_37249,N_35123);
nand U38560 (N_38560,N_36062,N_35314);
or U38561 (N_38561,N_37488,N_35405);
nand U38562 (N_38562,N_36416,N_36886);
nor U38563 (N_38563,N_36005,N_36503);
xnor U38564 (N_38564,N_37098,N_37126);
xnor U38565 (N_38565,N_36710,N_37452);
nor U38566 (N_38566,N_35295,N_37208);
nand U38567 (N_38567,N_36329,N_36187);
or U38568 (N_38568,N_35585,N_35740);
and U38569 (N_38569,N_36756,N_36514);
nor U38570 (N_38570,N_35372,N_35984);
and U38571 (N_38571,N_35649,N_36085);
xnor U38572 (N_38572,N_35418,N_36537);
nor U38573 (N_38573,N_35127,N_35508);
nor U38574 (N_38574,N_36879,N_35702);
nor U38575 (N_38575,N_36966,N_36868);
and U38576 (N_38576,N_36435,N_35618);
xor U38577 (N_38577,N_35484,N_35210);
or U38578 (N_38578,N_35590,N_37486);
and U38579 (N_38579,N_37001,N_37365);
or U38580 (N_38580,N_36225,N_37318);
or U38581 (N_38581,N_36622,N_37096);
and U38582 (N_38582,N_35551,N_35853);
or U38583 (N_38583,N_36381,N_35200);
nand U38584 (N_38584,N_36024,N_37367);
and U38585 (N_38585,N_36665,N_35625);
or U38586 (N_38586,N_35169,N_36953);
nor U38587 (N_38587,N_37358,N_36781);
xor U38588 (N_38588,N_35831,N_37243);
and U38589 (N_38589,N_37355,N_35825);
or U38590 (N_38590,N_36700,N_37469);
or U38591 (N_38591,N_35413,N_36382);
and U38592 (N_38592,N_36030,N_36351);
and U38593 (N_38593,N_36969,N_36313);
and U38594 (N_38594,N_36448,N_36891);
or U38595 (N_38595,N_36801,N_37325);
xor U38596 (N_38596,N_35241,N_36406);
xnor U38597 (N_38597,N_36646,N_35056);
or U38598 (N_38598,N_35486,N_36835);
xnor U38599 (N_38599,N_37228,N_36639);
xor U38600 (N_38600,N_35360,N_36682);
xor U38601 (N_38601,N_35072,N_35639);
nand U38602 (N_38602,N_37324,N_35735);
and U38603 (N_38603,N_37476,N_35757);
nand U38604 (N_38604,N_35205,N_37044);
nor U38605 (N_38605,N_35162,N_36856);
xor U38606 (N_38606,N_35654,N_37151);
nand U38607 (N_38607,N_36874,N_36584);
and U38608 (N_38608,N_37392,N_37136);
and U38609 (N_38609,N_35428,N_35778);
nor U38610 (N_38610,N_36330,N_36660);
nor U38611 (N_38611,N_36076,N_35720);
xnor U38612 (N_38612,N_36645,N_35761);
xnor U38613 (N_38613,N_35813,N_35954);
nand U38614 (N_38614,N_35059,N_36339);
nor U38615 (N_38615,N_36568,N_35983);
nor U38616 (N_38616,N_36597,N_37496);
xnor U38617 (N_38617,N_37050,N_37498);
xor U38618 (N_38618,N_37376,N_35686);
or U38619 (N_38619,N_35611,N_35214);
nand U38620 (N_38620,N_36630,N_35017);
and U38621 (N_38621,N_36795,N_37192);
or U38622 (N_38622,N_35157,N_35038);
and U38623 (N_38623,N_36593,N_36787);
or U38624 (N_38624,N_36041,N_35688);
nand U38625 (N_38625,N_36150,N_37274);
xnor U38626 (N_38626,N_37348,N_35913);
nor U38627 (N_38627,N_36532,N_36434);
nor U38628 (N_38628,N_37234,N_36429);
nor U38629 (N_38629,N_35312,N_35150);
or U38630 (N_38630,N_36338,N_36502);
xnor U38631 (N_38631,N_36368,N_36213);
or U38632 (N_38632,N_36451,N_36535);
nor U38633 (N_38633,N_37354,N_35226);
nor U38634 (N_38634,N_35142,N_37447);
nor U38635 (N_38635,N_36218,N_36267);
and U38636 (N_38636,N_36119,N_35262);
nand U38637 (N_38637,N_35691,N_36826);
and U38638 (N_38638,N_36833,N_35212);
or U38639 (N_38639,N_37468,N_37128);
nand U38640 (N_38640,N_35046,N_35822);
nor U38641 (N_38641,N_35346,N_37155);
or U38642 (N_38642,N_35966,N_35629);
nor U38643 (N_38643,N_35389,N_37189);
nand U38644 (N_38644,N_35145,N_37205);
nand U38645 (N_38645,N_36475,N_35332);
nand U38646 (N_38646,N_35385,N_36641);
xnor U38647 (N_38647,N_35110,N_37336);
nand U38648 (N_38648,N_37187,N_35728);
or U38649 (N_38649,N_35196,N_36454);
nor U38650 (N_38650,N_36998,N_36538);
nand U38651 (N_38651,N_36689,N_35962);
and U38652 (N_38652,N_35901,N_36595);
xnor U38653 (N_38653,N_35447,N_35055);
nand U38654 (N_38654,N_35248,N_36152);
nor U38655 (N_38655,N_35874,N_36655);
and U38656 (N_38656,N_37314,N_36846);
nand U38657 (N_38657,N_36617,N_36681);
and U38658 (N_38658,N_37080,N_37481);
and U38659 (N_38659,N_37466,N_35526);
and U38660 (N_38660,N_35658,N_35483);
or U38661 (N_38661,N_37144,N_37108);
nor U38662 (N_38662,N_37361,N_37111);
and U38663 (N_38663,N_35627,N_36147);
nor U38664 (N_38664,N_37299,N_35550);
or U38665 (N_38665,N_37467,N_36042);
and U38666 (N_38666,N_36893,N_37419);
nand U38667 (N_38667,N_37377,N_35424);
nand U38668 (N_38668,N_35850,N_36237);
nand U38669 (N_38669,N_35660,N_36355);
nand U38670 (N_38670,N_37477,N_35533);
and U38671 (N_38671,N_36968,N_37379);
xor U38672 (N_38672,N_36023,N_35489);
or U38673 (N_38673,N_35149,N_36004);
and U38674 (N_38674,N_35001,N_35734);
or U38675 (N_38675,N_37213,N_37088);
xor U38676 (N_38676,N_36051,N_36992);
nand U38677 (N_38677,N_35404,N_36553);
and U38678 (N_38678,N_35298,N_36192);
or U38679 (N_38679,N_37201,N_37220);
xor U38680 (N_38680,N_36785,N_36917);
nor U38681 (N_38681,N_37105,N_35892);
and U38682 (N_38682,N_35101,N_36483);
nand U38683 (N_38683,N_35576,N_37479);
xnor U38684 (N_38684,N_36153,N_36533);
or U38685 (N_38685,N_35485,N_36273);
or U38686 (N_38686,N_36934,N_36615);
and U38687 (N_38687,N_36002,N_35931);
nand U38688 (N_38688,N_35423,N_37056);
nand U38689 (N_38689,N_36822,N_35863);
or U38690 (N_38690,N_36566,N_36219);
or U38691 (N_38691,N_35185,N_36697);
nor U38692 (N_38692,N_36774,N_35782);
nand U38693 (N_38693,N_36875,N_35075);
or U38694 (N_38694,N_36752,N_35943);
and U38695 (N_38695,N_37269,N_37313);
and U38696 (N_38696,N_35082,N_36674);
xnor U38697 (N_38697,N_35228,N_35864);
or U38698 (N_38698,N_35091,N_35222);
nor U38699 (N_38699,N_36230,N_35661);
nor U38700 (N_38700,N_35342,N_35313);
and U38701 (N_38701,N_37312,N_36285);
nor U38702 (N_38702,N_35277,N_36916);
xnor U38703 (N_38703,N_35869,N_35435);
nand U38704 (N_38704,N_35575,N_36486);
nor U38705 (N_38705,N_37359,N_36477);
and U38706 (N_38706,N_35918,N_36400);
xor U38707 (N_38707,N_36887,N_36588);
nor U38708 (N_38708,N_37229,N_36251);
nand U38709 (N_38709,N_35973,N_36751);
nand U38710 (N_38710,N_36387,N_35281);
and U38711 (N_38711,N_35827,N_37198);
or U38712 (N_38712,N_35410,N_35378);
and U38713 (N_38713,N_36440,N_35857);
xnor U38714 (N_38714,N_35730,N_37084);
and U38715 (N_38715,N_35362,N_35490);
xor U38716 (N_38716,N_36407,N_35880);
nand U38717 (N_38717,N_35749,N_35619);
and U38718 (N_38718,N_36563,N_35054);
nor U38719 (N_38719,N_35509,N_35543);
nand U38720 (N_38720,N_35881,N_37109);
nand U38721 (N_38721,N_35118,N_36698);
or U38722 (N_38722,N_37290,N_35532);
or U38723 (N_38723,N_35744,N_35373);
nand U38724 (N_38724,N_36586,N_35855);
nor U38725 (N_38725,N_36735,N_35453);
nor U38726 (N_38726,N_35163,N_36117);
or U38727 (N_38727,N_36808,N_37186);
and U38728 (N_38728,N_36578,N_36876);
nand U38729 (N_38729,N_35653,N_35080);
and U38730 (N_38730,N_35194,N_35217);
nand U38731 (N_38731,N_36877,N_35440);
xnor U38732 (N_38732,N_37020,N_35946);
nor U38733 (N_38733,N_37416,N_36361);
and U38734 (N_38734,N_35828,N_35498);
nand U38735 (N_38735,N_37121,N_36922);
or U38736 (N_38736,N_36673,N_37400);
nand U38737 (N_38737,N_36436,N_37300);
nor U38738 (N_38738,N_36276,N_35138);
nand U38739 (N_38739,N_36025,N_36914);
and U38740 (N_38740,N_35166,N_35290);
or U38741 (N_38741,N_36050,N_37221);
nand U38742 (N_38742,N_35587,N_35393);
nor U38743 (N_38743,N_35632,N_37397);
nor U38744 (N_38744,N_35794,N_37368);
nor U38745 (N_38745,N_36445,N_35201);
xnor U38746 (N_38746,N_35450,N_35663);
xnor U38747 (N_38747,N_36605,N_35494);
or U38748 (N_38748,N_35350,N_35396);
xnor U38749 (N_38749,N_36528,N_37374);
xor U38750 (N_38750,N_35069,N_36149);
nand U38751 (N_38751,N_35673,N_36070);
or U38752 (N_38752,N_35164,N_36251);
xnor U38753 (N_38753,N_37421,N_35435);
xnor U38754 (N_38754,N_36412,N_35660);
xnor U38755 (N_38755,N_37484,N_36326);
or U38756 (N_38756,N_36729,N_36132);
nand U38757 (N_38757,N_36031,N_35009);
or U38758 (N_38758,N_36946,N_37324);
nand U38759 (N_38759,N_36409,N_36079);
nor U38760 (N_38760,N_37415,N_37140);
nand U38761 (N_38761,N_35055,N_36230);
or U38762 (N_38762,N_36333,N_35923);
nand U38763 (N_38763,N_36972,N_37327);
nand U38764 (N_38764,N_37426,N_36695);
nand U38765 (N_38765,N_36999,N_35838);
or U38766 (N_38766,N_36652,N_35386);
and U38767 (N_38767,N_37106,N_35359);
nand U38768 (N_38768,N_37462,N_36860);
xnor U38769 (N_38769,N_37207,N_36334);
nor U38770 (N_38770,N_35485,N_37140);
nor U38771 (N_38771,N_35968,N_36752);
xor U38772 (N_38772,N_36244,N_36405);
or U38773 (N_38773,N_37256,N_36292);
nor U38774 (N_38774,N_35022,N_35348);
xor U38775 (N_38775,N_37273,N_35925);
or U38776 (N_38776,N_37319,N_35819);
nor U38777 (N_38777,N_36594,N_36676);
nor U38778 (N_38778,N_35380,N_35716);
xor U38779 (N_38779,N_36069,N_35247);
nor U38780 (N_38780,N_35809,N_36708);
or U38781 (N_38781,N_35514,N_35554);
nor U38782 (N_38782,N_37108,N_36417);
and U38783 (N_38783,N_35011,N_35713);
or U38784 (N_38784,N_37139,N_36612);
and U38785 (N_38785,N_35427,N_35400);
or U38786 (N_38786,N_35307,N_36332);
nand U38787 (N_38787,N_36969,N_37148);
nand U38788 (N_38788,N_36800,N_35484);
nand U38789 (N_38789,N_36653,N_35535);
and U38790 (N_38790,N_35274,N_35110);
nand U38791 (N_38791,N_36382,N_35442);
nor U38792 (N_38792,N_35016,N_36230);
or U38793 (N_38793,N_36019,N_35651);
nor U38794 (N_38794,N_37277,N_35937);
nand U38795 (N_38795,N_36652,N_35129);
and U38796 (N_38796,N_35696,N_35837);
xor U38797 (N_38797,N_36016,N_35682);
and U38798 (N_38798,N_35081,N_35506);
and U38799 (N_38799,N_36625,N_35813);
or U38800 (N_38800,N_37156,N_35413);
nand U38801 (N_38801,N_36248,N_35705);
nand U38802 (N_38802,N_35768,N_36461);
or U38803 (N_38803,N_35968,N_37388);
and U38804 (N_38804,N_35758,N_36493);
nor U38805 (N_38805,N_36187,N_35310);
xnor U38806 (N_38806,N_36819,N_36680);
or U38807 (N_38807,N_36874,N_37400);
xnor U38808 (N_38808,N_35868,N_36691);
xnor U38809 (N_38809,N_36930,N_35068);
and U38810 (N_38810,N_35160,N_36936);
nor U38811 (N_38811,N_35920,N_36191);
nor U38812 (N_38812,N_35235,N_36011);
xnor U38813 (N_38813,N_35600,N_36516);
nand U38814 (N_38814,N_35193,N_36556);
nand U38815 (N_38815,N_37264,N_36027);
nor U38816 (N_38816,N_35977,N_35765);
or U38817 (N_38817,N_36516,N_36592);
xor U38818 (N_38818,N_35658,N_37268);
and U38819 (N_38819,N_37153,N_37478);
or U38820 (N_38820,N_35996,N_37419);
or U38821 (N_38821,N_37117,N_35699);
or U38822 (N_38822,N_36841,N_35382);
nor U38823 (N_38823,N_36286,N_37120);
and U38824 (N_38824,N_36072,N_35248);
or U38825 (N_38825,N_35585,N_36416);
and U38826 (N_38826,N_35353,N_35441);
nor U38827 (N_38827,N_35286,N_35768);
nand U38828 (N_38828,N_35589,N_37142);
nand U38829 (N_38829,N_36086,N_36493);
and U38830 (N_38830,N_35199,N_36024);
nor U38831 (N_38831,N_37223,N_37250);
nor U38832 (N_38832,N_37208,N_36614);
or U38833 (N_38833,N_36050,N_36700);
or U38834 (N_38834,N_35207,N_35959);
and U38835 (N_38835,N_35997,N_35092);
nor U38836 (N_38836,N_36751,N_35193);
and U38837 (N_38837,N_35018,N_36969);
nand U38838 (N_38838,N_35907,N_36082);
xor U38839 (N_38839,N_35125,N_35310);
and U38840 (N_38840,N_36274,N_35400);
or U38841 (N_38841,N_35662,N_37200);
and U38842 (N_38842,N_37465,N_37229);
or U38843 (N_38843,N_36621,N_36085);
nor U38844 (N_38844,N_35863,N_36091);
xnor U38845 (N_38845,N_35879,N_35568);
or U38846 (N_38846,N_36762,N_37152);
and U38847 (N_38847,N_35218,N_37276);
nor U38848 (N_38848,N_36031,N_35011);
xnor U38849 (N_38849,N_36591,N_37249);
or U38850 (N_38850,N_35520,N_36845);
xor U38851 (N_38851,N_36165,N_35873);
nor U38852 (N_38852,N_37338,N_36440);
or U38853 (N_38853,N_35599,N_35183);
nand U38854 (N_38854,N_36598,N_36467);
nor U38855 (N_38855,N_36853,N_36251);
nand U38856 (N_38856,N_36585,N_37339);
nand U38857 (N_38857,N_36543,N_35125);
or U38858 (N_38858,N_36670,N_36386);
nor U38859 (N_38859,N_37134,N_36099);
nor U38860 (N_38860,N_35618,N_35873);
nand U38861 (N_38861,N_36550,N_36526);
and U38862 (N_38862,N_35099,N_36765);
xnor U38863 (N_38863,N_35266,N_35325);
nor U38864 (N_38864,N_35135,N_37292);
nand U38865 (N_38865,N_35911,N_36891);
nor U38866 (N_38866,N_36262,N_37112);
nand U38867 (N_38867,N_37067,N_35430);
or U38868 (N_38868,N_37229,N_35925);
and U38869 (N_38869,N_35168,N_36453);
and U38870 (N_38870,N_37190,N_35239);
and U38871 (N_38871,N_35292,N_36155);
or U38872 (N_38872,N_35287,N_37173);
xnor U38873 (N_38873,N_36714,N_35072);
xnor U38874 (N_38874,N_36921,N_36409);
or U38875 (N_38875,N_37099,N_35014);
or U38876 (N_38876,N_36384,N_37261);
nand U38877 (N_38877,N_37102,N_36632);
or U38878 (N_38878,N_37089,N_36373);
nand U38879 (N_38879,N_36091,N_37361);
nor U38880 (N_38880,N_36863,N_36826);
nand U38881 (N_38881,N_35324,N_36142);
or U38882 (N_38882,N_36019,N_35846);
and U38883 (N_38883,N_35632,N_35053);
or U38884 (N_38884,N_35546,N_36465);
or U38885 (N_38885,N_35167,N_36495);
nand U38886 (N_38886,N_36845,N_35678);
or U38887 (N_38887,N_35459,N_36260);
and U38888 (N_38888,N_36013,N_36687);
nor U38889 (N_38889,N_36008,N_37352);
nor U38890 (N_38890,N_35540,N_35395);
xnor U38891 (N_38891,N_36468,N_35993);
nor U38892 (N_38892,N_37156,N_36426);
xnor U38893 (N_38893,N_37344,N_36058);
xnor U38894 (N_38894,N_35158,N_37454);
xor U38895 (N_38895,N_36225,N_35541);
nand U38896 (N_38896,N_36631,N_37361);
and U38897 (N_38897,N_35033,N_36220);
nor U38898 (N_38898,N_36285,N_37072);
or U38899 (N_38899,N_36799,N_36441);
nor U38900 (N_38900,N_37107,N_37126);
or U38901 (N_38901,N_37468,N_37405);
nor U38902 (N_38902,N_36581,N_35118);
xnor U38903 (N_38903,N_37122,N_36981);
or U38904 (N_38904,N_35989,N_36237);
nor U38905 (N_38905,N_36938,N_35859);
xnor U38906 (N_38906,N_35473,N_37449);
or U38907 (N_38907,N_36383,N_37180);
or U38908 (N_38908,N_35279,N_36613);
or U38909 (N_38909,N_35749,N_35082);
nand U38910 (N_38910,N_35002,N_35506);
or U38911 (N_38911,N_36413,N_36051);
nand U38912 (N_38912,N_36889,N_35990);
nor U38913 (N_38913,N_35272,N_35852);
xor U38914 (N_38914,N_36975,N_35436);
and U38915 (N_38915,N_36005,N_35408);
nand U38916 (N_38916,N_36018,N_36079);
nor U38917 (N_38917,N_36461,N_36260);
xor U38918 (N_38918,N_37215,N_36538);
or U38919 (N_38919,N_35774,N_35660);
nor U38920 (N_38920,N_37159,N_37464);
nor U38921 (N_38921,N_36760,N_36482);
nor U38922 (N_38922,N_36556,N_35679);
xor U38923 (N_38923,N_36374,N_35282);
nor U38924 (N_38924,N_35878,N_35280);
nor U38925 (N_38925,N_35198,N_36579);
and U38926 (N_38926,N_35649,N_35762);
and U38927 (N_38927,N_36751,N_37254);
or U38928 (N_38928,N_36339,N_36042);
xnor U38929 (N_38929,N_35871,N_36099);
and U38930 (N_38930,N_36726,N_35823);
xnor U38931 (N_38931,N_37171,N_35985);
xnor U38932 (N_38932,N_36621,N_36505);
or U38933 (N_38933,N_36820,N_36724);
or U38934 (N_38934,N_35116,N_36960);
xnor U38935 (N_38935,N_37173,N_36172);
xnor U38936 (N_38936,N_37156,N_35697);
or U38937 (N_38937,N_35202,N_35507);
xor U38938 (N_38938,N_36784,N_35595);
nor U38939 (N_38939,N_37073,N_35493);
xor U38940 (N_38940,N_37400,N_36875);
nor U38941 (N_38941,N_36071,N_36791);
nor U38942 (N_38942,N_35704,N_37092);
or U38943 (N_38943,N_37017,N_36072);
xnor U38944 (N_38944,N_36997,N_35811);
nor U38945 (N_38945,N_36357,N_35955);
or U38946 (N_38946,N_36242,N_36860);
and U38947 (N_38947,N_36691,N_35158);
or U38948 (N_38948,N_36596,N_37202);
or U38949 (N_38949,N_35170,N_35909);
xor U38950 (N_38950,N_37394,N_35786);
xnor U38951 (N_38951,N_36497,N_36947);
or U38952 (N_38952,N_36861,N_36276);
xnor U38953 (N_38953,N_35022,N_37076);
or U38954 (N_38954,N_35371,N_37395);
xnor U38955 (N_38955,N_37288,N_35674);
nor U38956 (N_38956,N_35050,N_35844);
xor U38957 (N_38957,N_36839,N_36893);
nand U38958 (N_38958,N_35384,N_36904);
xnor U38959 (N_38959,N_36790,N_35943);
nor U38960 (N_38960,N_37239,N_35107);
nor U38961 (N_38961,N_35237,N_36611);
or U38962 (N_38962,N_35969,N_36712);
or U38963 (N_38963,N_36387,N_35710);
or U38964 (N_38964,N_35923,N_35195);
nor U38965 (N_38965,N_36465,N_36867);
xnor U38966 (N_38966,N_35680,N_36273);
xor U38967 (N_38967,N_35503,N_35311);
nor U38968 (N_38968,N_37459,N_37304);
and U38969 (N_38969,N_37052,N_36614);
nor U38970 (N_38970,N_35225,N_35550);
xor U38971 (N_38971,N_35494,N_36475);
nand U38972 (N_38972,N_35781,N_36180);
and U38973 (N_38973,N_37011,N_36116);
xor U38974 (N_38974,N_35596,N_37402);
and U38975 (N_38975,N_36263,N_36728);
or U38976 (N_38976,N_36942,N_36380);
xor U38977 (N_38977,N_35087,N_35726);
xnor U38978 (N_38978,N_37405,N_36292);
nand U38979 (N_38979,N_36029,N_35149);
xnor U38980 (N_38980,N_35599,N_37269);
and U38981 (N_38981,N_35127,N_37290);
nand U38982 (N_38982,N_37490,N_37296);
nand U38983 (N_38983,N_35570,N_37396);
or U38984 (N_38984,N_36913,N_35932);
or U38985 (N_38985,N_37149,N_35942);
nand U38986 (N_38986,N_35628,N_36465);
nor U38987 (N_38987,N_36816,N_36893);
xor U38988 (N_38988,N_36836,N_35773);
nand U38989 (N_38989,N_36033,N_36230);
nor U38990 (N_38990,N_35913,N_36297);
and U38991 (N_38991,N_36654,N_36066);
xor U38992 (N_38992,N_35874,N_36948);
or U38993 (N_38993,N_37005,N_35578);
or U38994 (N_38994,N_37126,N_35941);
or U38995 (N_38995,N_36951,N_35748);
nor U38996 (N_38996,N_36471,N_35786);
nand U38997 (N_38997,N_35244,N_35728);
and U38998 (N_38998,N_36392,N_35407);
xor U38999 (N_38999,N_36262,N_37356);
nand U39000 (N_39000,N_37405,N_37170);
and U39001 (N_39001,N_37453,N_35690);
nand U39002 (N_39002,N_35068,N_35581);
or U39003 (N_39003,N_37136,N_36223);
nand U39004 (N_39004,N_35532,N_35354);
or U39005 (N_39005,N_36945,N_35068);
nor U39006 (N_39006,N_37242,N_35379);
nand U39007 (N_39007,N_35134,N_37384);
nor U39008 (N_39008,N_36452,N_36959);
nand U39009 (N_39009,N_36751,N_35338);
nor U39010 (N_39010,N_35707,N_35485);
and U39011 (N_39011,N_35329,N_35894);
and U39012 (N_39012,N_35813,N_36758);
and U39013 (N_39013,N_36201,N_36350);
or U39014 (N_39014,N_36315,N_37308);
and U39015 (N_39015,N_35503,N_37192);
and U39016 (N_39016,N_35495,N_36788);
nand U39017 (N_39017,N_35417,N_35668);
or U39018 (N_39018,N_35760,N_36197);
or U39019 (N_39019,N_36094,N_36487);
nand U39020 (N_39020,N_35944,N_35764);
nor U39021 (N_39021,N_35575,N_36183);
and U39022 (N_39022,N_36892,N_35424);
nor U39023 (N_39023,N_35785,N_35179);
nor U39024 (N_39024,N_36462,N_37378);
nand U39025 (N_39025,N_37466,N_36512);
nor U39026 (N_39026,N_37224,N_35877);
nor U39027 (N_39027,N_36787,N_35396);
and U39028 (N_39028,N_36975,N_35017);
nand U39029 (N_39029,N_36520,N_35601);
or U39030 (N_39030,N_35089,N_35683);
and U39031 (N_39031,N_36836,N_37036);
and U39032 (N_39032,N_35451,N_35321);
nand U39033 (N_39033,N_36954,N_37286);
nor U39034 (N_39034,N_36830,N_37311);
nand U39035 (N_39035,N_35991,N_36128);
xnor U39036 (N_39036,N_36639,N_36120);
and U39037 (N_39037,N_37354,N_37380);
or U39038 (N_39038,N_35160,N_36447);
nand U39039 (N_39039,N_36970,N_36976);
nor U39040 (N_39040,N_36176,N_37341);
or U39041 (N_39041,N_37430,N_35443);
xnor U39042 (N_39042,N_35954,N_37090);
and U39043 (N_39043,N_35519,N_35042);
nor U39044 (N_39044,N_37087,N_36481);
nor U39045 (N_39045,N_36428,N_36465);
nand U39046 (N_39046,N_36554,N_37078);
xnor U39047 (N_39047,N_36979,N_37384);
and U39048 (N_39048,N_37388,N_36761);
xnor U39049 (N_39049,N_35011,N_35716);
and U39050 (N_39050,N_36898,N_36201);
and U39051 (N_39051,N_37092,N_35139);
or U39052 (N_39052,N_35114,N_35884);
nor U39053 (N_39053,N_36385,N_36614);
or U39054 (N_39054,N_35169,N_35765);
and U39055 (N_39055,N_37250,N_36267);
or U39056 (N_39056,N_36924,N_36390);
and U39057 (N_39057,N_36492,N_37081);
and U39058 (N_39058,N_36507,N_36328);
nand U39059 (N_39059,N_36276,N_37203);
xnor U39060 (N_39060,N_35735,N_35999);
nand U39061 (N_39061,N_36811,N_36248);
or U39062 (N_39062,N_35111,N_37195);
and U39063 (N_39063,N_36807,N_37165);
or U39064 (N_39064,N_36828,N_36360);
and U39065 (N_39065,N_36427,N_36407);
nand U39066 (N_39066,N_35774,N_35994);
nor U39067 (N_39067,N_36210,N_36605);
or U39068 (N_39068,N_35096,N_35090);
nand U39069 (N_39069,N_36097,N_35953);
and U39070 (N_39070,N_36986,N_37492);
xor U39071 (N_39071,N_36317,N_35667);
nor U39072 (N_39072,N_37118,N_35144);
and U39073 (N_39073,N_37466,N_36033);
nor U39074 (N_39074,N_36383,N_36596);
xor U39075 (N_39075,N_35269,N_36782);
nand U39076 (N_39076,N_35592,N_35654);
nor U39077 (N_39077,N_35319,N_36214);
nand U39078 (N_39078,N_35770,N_36618);
xor U39079 (N_39079,N_35153,N_35370);
nor U39080 (N_39080,N_35370,N_36953);
nand U39081 (N_39081,N_37241,N_35397);
and U39082 (N_39082,N_37136,N_35927);
nor U39083 (N_39083,N_37272,N_35924);
or U39084 (N_39084,N_35269,N_37335);
or U39085 (N_39085,N_36475,N_35819);
or U39086 (N_39086,N_36127,N_36240);
and U39087 (N_39087,N_35614,N_35842);
or U39088 (N_39088,N_35535,N_37413);
xnor U39089 (N_39089,N_36531,N_36133);
xor U39090 (N_39090,N_35137,N_36003);
xnor U39091 (N_39091,N_36230,N_36641);
xor U39092 (N_39092,N_37441,N_36313);
nor U39093 (N_39093,N_36365,N_36764);
xor U39094 (N_39094,N_35382,N_37275);
nor U39095 (N_39095,N_36198,N_35337);
nor U39096 (N_39096,N_35632,N_36755);
or U39097 (N_39097,N_35492,N_35646);
or U39098 (N_39098,N_36582,N_36506);
xnor U39099 (N_39099,N_35793,N_35065);
xor U39100 (N_39100,N_35012,N_36534);
or U39101 (N_39101,N_36615,N_35988);
nor U39102 (N_39102,N_35049,N_37253);
and U39103 (N_39103,N_36268,N_36332);
or U39104 (N_39104,N_36168,N_36647);
xor U39105 (N_39105,N_36249,N_36932);
or U39106 (N_39106,N_35600,N_36560);
and U39107 (N_39107,N_35304,N_37347);
nand U39108 (N_39108,N_36380,N_36955);
and U39109 (N_39109,N_36276,N_35607);
nor U39110 (N_39110,N_36652,N_35679);
xor U39111 (N_39111,N_35304,N_35171);
nand U39112 (N_39112,N_36548,N_35040);
nor U39113 (N_39113,N_35467,N_36812);
nor U39114 (N_39114,N_35701,N_36842);
xor U39115 (N_39115,N_37435,N_37124);
or U39116 (N_39116,N_35295,N_36079);
nand U39117 (N_39117,N_36335,N_35058);
xnor U39118 (N_39118,N_36766,N_36824);
nand U39119 (N_39119,N_36167,N_36596);
or U39120 (N_39120,N_35944,N_37465);
or U39121 (N_39121,N_36087,N_36072);
xor U39122 (N_39122,N_35116,N_36435);
and U39123 (N_39123,N_36499,N_35277);
nor U39124 (N_39124,N_36633,N_35233);
xor U39125 (N_39125,N_36581,N_36501);
nor U39126 (N_39126,N_36025,N_35931);
xor U39127 (N_39127,N_36686,N_35773);
and U39128 (N_39128,N_37213,N_36051);
nor U39129 (N_39129,N_36388,N_35142);
or U39130 (N_39130,N_35245,N_36363);
xor U39131 (N_39131,N_35306,N_36264);
nand U39132 (N_39132,N_37331,N_37279);
xnor U39133 (N_39133,N_36891,N_37135);
nor U39134 (N_39134,N_36040,N_36715);
and U39135 (N_39135,N_37344,N_35974);
or U39136 (N_39136,N_36452,N_37212);
or U39137 (N_39137,N_36856,N_36286);
nor U39138 (N_39138,N_36020,N_35771);
or U39139 (N_39139,N_36901,N_35602);
xor U39140 (N_39140,N_36639,N_35084);
nand U39141 (N_39141,N_35607,N_36108);
xnor U39142 (N_39142,N_35218,N_35918);
and U39143 (N_39143,N_35155,N_36293);
and U39144 (N_39144,N_37330,N_35268);
xor U39145 (N_39145,N_35589,N_35877);
xnor U39146 (N_39146,N_35085,N_37139);
xnor U39147 (N_39147,N_35648,N_35824);
or U39148 (N_39148,N_35882,N_35163);
nor U39149 (N_39149,N_35773,N_36701);
or U39150 (N_39150,N_35416,N_37009);
xnor U39151 (N_39151,N_35698,N_37415);
nand U39152 (N_39152,N_36410,N_37008);
nand U39153 (N_39153,N_37333,N_37372);
nor U39154 (N_39154,N_36525,N_35645);
and U39155 (N_39155,N_35846,N_35411);
nand U39156 (N_39156,N_36838,N_35350);
or U39157 (N_39157,N_35178,N_37008);
nor U39158 (N_39158,N_37199,N_35736);
xor U39159 (N_39159,N_35570,N_37338);
or U39160 (N_39160,N_37268,N_36126);
and U39161 (N_39161,N_37113,N_35316);
nand U39162 (N_39162,N_36010,N_36297);
nor U39163 (N_39163,N_37002,N_36438);
or U39164 (N_39164,N_36579,N_36871);
or U39165 (N_39165,N_36674,N_35192);
xor U39166 (N_39166,N_37496,N_36060);
and U39167 (N_39167,N_35885,N_35286);
nand U39168 (N_39168,N_35601,N_35467);
and U39169 (N_39169,N_37437,N_35193);
nor U39170 (N_39170,N_37440,N_36936);
xnor U39171 (N_39171,N_35923,N_36023);
nor U39172 (N_39172,N_37096,N_37177);
and U39173 (N_39173,N_37118,N_36307);
or U39174 (N_39174,N_37221,N_35478);
xnor U39175 (N_39175,N_36073,N_37126);
nor U39176 (N_39176,N_36840,N_37475);
xor U39177 (N_39177,N_36768,N_36471);
nor U39178 (N_39178,N_35733,N_35497);
or U39179 (N_39179,N_35138,N_37222);
nor U39180 (N_39180,N_36140,N_37049);
and U39181 (N_39181,N_37104,N_37495);
and U39182 (N_39182,N_35091,N_36110);
or U39183 (N_39183,N_35803,N_36149);
or U39184 (N_39184,N_36234,N_36140);
nand U39185 (N_39185,N_35126,N_35376);
or U39186 (N_39186,N_36162,N_35138);
xnor U39187 (N_39187,N_35788,N_36300);
nor U39188 (N_39188,N_36472,N_36848);
nor U39189 (N_39189,N_37054,N_36367);
nand U39190 (N_39190,N_37394,N_35730);
nand U39191 (N_39191,N_35751,N_36992);
or U39192 (N_39192,N_36636,N_35491);
or U39193 (N_39193,N_37294,N_36482);
nand U39194 (N_39194,N_36558,N_37009);
nor U39195 (N_39195,N_35719,N_35248);
xor U39196 (N_39196,N_36745,N_37275);
and U39197 (N_39197,N_35952,N_35184);
and U39198 (N_39198,N_36495,N_36531);
nand U39199 (N_39199,N_36898,N_35227);
xnor U39200 (N_39200,N_35719,N_35430);
nor U39201 (N_39201,N_37447,N_36967);
nand U39202 (N_39202,N_35229,N_35598);
xor U39203 (N_39203,N_37282,N_35428);
nor U39204 (N_39204,N_35651,N_35819);
xor U39205 (N_39205,N_35753,N_36411);
or U39206 (N_39206,N_37027,N_36574);
xor U39207 (N_39207,N_35105,N_36066);
nor U39208 (N_39208,N_36283,N_36502);
nand U39209 (N_39209,N_36704,N_35509);
and U39210 (N_39210,N_36070,N_37329);
and U39211 (N_39211,N_35604,N_35581);
and U39212 (N_39212,N_35943,N_35784);
nor U39213 (N_39213,N_35256,N_36543);
nor U39214 (N_39214,N_36696,N_36576);
nor U39215 (N_39215,N_37094,N_35535);
and U39216 (N_39216,N_36025,N_36594);
nand U39217 (N_39217,N_35989,N_36833);
nor U39218 (N_39218,N_35581,N_35141);
and U39219 (N_39219,N_35523,N_35798);
xor U39220 (N_39220,N_35044,N_35475);
nand U39221 (N_39221,N_35038,N_37220);
or U39222 (N_39222,N_35471,N_35997);
or U39223 (N_39223,N_35700,N_35934);
and U39224 (N_39224,N_37068,N_36985);
or U39225 (N_39225,N_36301,N_36302);
nor U39226 (N_39226,N_36868,N_37478);
and U39227 (N_39227,N_36633,N_37341);
and U39228 (N_39228,N_36067,N_35226);
xor U39229 (N_39229,N_37016,N_36704);
xnor U39230 (N_39230,N_36383,N_36222);
nor U39231 (N_39231,N_36379,N_36225);
nor U39232 (N_39232,N_35285,N_36983);
or U39233 (N_39233,N_37290,N_35317);
or U39234 (N_39234,N_35873,N_37219);
or U39235 (N_39235,N_35102,N_35687);
or U39236 (N_39236,N_35945,N_35335);
xnor U39237 (N_39237,N_36937,N_35637);
xnor U39238 (N_39238,N_36415,N_36688);
nand U39239 (N_39239,N_37122,N_36222);
and U39240 (N_39240,N_35132,N_36734);
nor U39241 (N_39241,N_35472,N_35996);
or U39242 (N_39242,N_35113,N_35284);
xnor U39243 (N_39243,N_37166,N_36540);
nand U39244 (N_39244,N_37437,N_36580);
and U39245 (N_39245,N_37181,N_36495);
or U39246 (N_39246,N_35985,N_36267);
and U39247 (N_39247,N_35604,N_36517);
and U39248 (N_39248,N_35120,N_36184);
nor U39249 (N_39249,N_35059,N_36786);
nor U39250 (N_39250,N_36966,N_35542);
nor U39251 (N_39251,N_35237,N_36072);
or U39252 (N_39252,N_36376,N_35387);
and U39253 (N_39253,N_35599,N_35059);
and U39254 (N_39254,N_36217,N_36724);
nor U39255 (N_39255,N_36949,N_36812);
xor U39256 (N_39256,N_35089,N_35380);
or U39257 (N_39257,N_35313,N_35287);
xor U39258 (N_39258,N_37258,N_36114);
xnor U39259 (N_39259,N_36163,N_36735);
nand U39260 (N_39260,N_35793,N_36268);
and U39261 (N_39261,N_35249,N_35298);
or U39262 (N_39262,N_36493,N_37020);
and U39263 (N_39263,N_37101,N_36116);
and U39264 (N_39264,N_36464,N_35430);
or U39265 (N_39265,N_37205,N_36467);
nand U39266 (N_39266,N_36177,N_36926);
xnor U39267 (N_39267,N_35721,N_36392);
or U39268 (N_39268,N_37264,N_36279);
or U39269 (N_39269,N_37143,N_36597);
nor U39270 (N_39270,N_35507,N_35417);
and U39271 (N_39271,N_37327,N_36302);
nand U39272 (N_39272,N_37247,N_35233);
nand U39273 (N_39273,N_36747,N_36507);
and U39274 (N_39274,N_35939,N_36263);
and U39275 (N_39275,N_36751,N_36014);
and U39276 (N_39276,N_35269,N_35599);
nand U39277 (N_39277,N_35933,N_36764);
xnor U39278 (N_39278,N_35744,N_36109);
nor U39279 (N_39279,N_35667,N_36867);
or U39280 (N_39280,N_35599,N_37272);
nor U39281 (N_39281,N_36103,N_36621);
xor U39282 (N_39282,N_36759,N_35860);
or U39283 (N_39283,N_35203,N_35760);
xor U39284 (N_39284,N_35556,N_36894);
nor U39285 (N_39285,N_36764,N_35872);
nor U39286 (N_39286,N_36159,N_35204);
or U39287 (N_39287,N_37397,N_35447);
and U39288 (N_39288,N_36546,N_36429);
and U39289 (N_39289,N_37161,N_35244);
xnor U39290 (N_39290,N_35664,N_35887);
nand U39291 (N_39291,N_36813,N_35918);
nand U39292 (N_39292,N_37053,N_35904);
nand U39293 (N_39293,N_35241,N_35649);
and U39294 (N_39294,N_35678,N_36465);
nor U39295 (N_39295,N_36394,N_36596);
xor U39296 (N_39296,N_35206,N_35555);
xor U39297 (N_39297,N_36140,N_36696);
or U39298 (N_39298,N_37340,N_35892);
nand U39299 (N_39299,N_35895,N_35180);
xnor U39300 (N_39300,N_35521,N_35995);
or U39301 (N_39301,N_35082,N_35694);
nor U39302 (N_39302,N_36812,N_35153);
nand U39303 (N_39303,N_36513,N_35785);
and U39304 (N_39304,N_36212,N_35087);
or U39305 (N_39305,N_37367,N_37460);
nor U39306 (N_39306,N_35044,N_35553);
and U39307 (N_39307,N_35320,N_35642);
and U39308 (N_39308,N_36047,N_36794);
or U39309 (N_39309,N_35390,N_37488);
and U39310 (N_39310,N_36102,N_36993);
nor U39311 (N_39311,N_35509,N_35178);
or U39312 (N_39312,N_36098,N_35033);
or U39313 (N_39313,N_36610,N_37482);
and U39314 (N_39314,N_37365,N_37072);
xor U39315 (N_39315,N_35144,N_35431);
and U39316 (N_39316,N_36736,N_36719);
nor U39317 (N_39317,N_35499,N_36374);
xnor U39318 (N_39318,N_36427,N_35132);
nand U39319 (N_39319,N_35698,N_36511);
or U39320 (N_39320,N_36639,N_36931);
or U39321 (N_39321,N_36229,N_37305);
or U39322 (N_39322,N_36733,N_36177);
or U39323 (N_39323,N_36573,N_35293);
xnor U39324 (N_39324,N_35970,N_36538);
or U39325 (N_39325,N_36551,N_35188);
and U39326 (N_39326,N_36146,N_36648);
xor U39327 (N_39327,N_36494,N_36168);
nor U39328 (N_39328,N_36131,N_35064);
and U39329 (N_39329,N_36172,N_37008);
nor U39330 (N_39330,N_35496,N_35277);
xor U39331 (N_39331,N_35841,N_36895);
nand U39332 (N_39332,N_37449,N_36954);
xnor U39333 (N_39333,N_36508,N_36670);
or U39334 (N_39334,N_36923,N_36528);
and U39335 (N_39335,N_36786,N_35285);
and U39336 (N_39336,N_36053,N_36349);
xor U39337 (N_39337,N_36153,N_35071);
xnor U39338 (N_39338,N_35491,N_35705);
nor U39339 (N_39339,N_36831,N_36384);
nand U39340 (N_39340,N_35330,N_37362);
or U39341 (N_39341,N_36838,N_35493);
xnor U39342 (N_39342,N_37033,N_37136);
xor U39343 (N_39343,N_35152,N_35765);
or U39344 (N_39344,N_35945,N_37126);
and U39345 (N_39345,N_35749,N_35253);
and U39346 (N_39346,N_36840,N_36722);
xnor U39347 (N_39347,N_36761,N_36908);
nand U39348 (N_39348,N_35696,N_35201);
or U39349 (N_39349,N_35484,N_35862);
xnor U39350 (N_39350,N_36319,N_36589);
xnor U39351 (N_39351,N_35825,N_35890);
or U39352 (N_39352,N_37215,N_37320);
or U39353 (N_39353,N_36703,N_35790);
xnor U39354 (N_39354,N_35365,N_35373);
and U39355 (N_39355,N_35458,N_35077);
xnor U39356 (N_39356,N_36585,N_35917);
and U39357 (N_39357,N_35578,N_35721);
and U39358 (N_39358,N_36416,N_35033);
nand U39359 (N_39359,N_35600,N_37173);
and U39360 (N_39360,N_37435,N_36762);
nand U39361 (N_39361,N_35717,N_35558);
nand U39362 (N_39362,N_35044,N_35275);
or U39363 (N_39363,N_37481,N_37181);
and U39364 (N_39364,N_36900,N_35716);
nand U39365 (N_39365,N_35086,N_36614);
nand U39366 (N_39366,N_36945,N_35702);
or U39367 (N_39367,N_36436,N_35534);
and U39368 (N_39368,N_36800,N_37033);
and U39369 (N_39369,N_36093,N_36425);
nor U39370 (N_39370,N_35564,N_35279);
nand U39371 (N_39371,N_36389,N_35231);
nand U39372 (N_39372,N_36785,N_36906);
xor U39373 (N_39373,N_36245,N_37403);
xnor U39374 (N_39374,N_37126,N_35145);
or U39375 (N_39375,N_36763,N_35221);
xnor U39376 (N_39376,N_35426,N_36568);
nand U39377 (N_39377,N_35598,N_36604);
nand U39378 (N_39378,N_35884,N_37324);
or U39379 (N_39379,N_36336,N_36400);
or U39380 (N_39380,N_35175,N_37240);
and U39381 (N_39381,N_37473,N_35835);
or U39382 (N_39382,N_37092,N_36826);
and U39383 (N_39383,N_36128,N_35212);
and U39384 (N_39384,N_36092,N_36218);
xor U39385 (N_39385,N_36714,N_37150);
nor U39386 (N_39386,N_35284,N_35048);
and U39387 (N_39387,N_35609,N_35204);
nand U39388 (N_39388,N_37273,N_36072);
nor U39389 (N_39389,N_35765,N_36063);
or U39390 (N_39390,N_35593,N_36242);
and U39391 (N_39391,N_36767,N_37057);
nor U39392 (N_39392,N_37401,N_36796);
nand U39393 (N_39393,N_36811,N_36637);
or U39394 (N_39394,N_36508,N_37087);
nor U39395 (N_39395,N_36838,N_36126);
or U39396 (N_39396,N_37000,N_35134);
nand U39397 (N_39397,N_36704,N_35049);
xnor U39398 (N_39398,N_36807,N_35735);
and U39399 (N_39399,N_35772,N_36270);
nor U39400 (N_39400,N_36063,N_35044);
nor U39401 (N_39401,N_35458,N_37470);
nand U39402 (N_39402,N_36479,N_37297);
xor U39403 (N_39403,N_35264,N_36799);
xnor U39404 (N_39404,N_35351,N_35651);
xor U39405 (N_39405,N_36664,N_36516);
and U39406 (N_39406,N_35001,N_35521);
xnor U39407 (N_39407,N_35913,N_35332);
or U39408 (N_39408,N_36208,N_37114);
or U39409 (N_39409,N_35575,N_36778);
xor U39410 (N_39410,N_35081,N_35730);
nor U39411 (N_39411,N_37061,N_36152);
nor U39412 (N_39412,N_36157,N_35577);
and U39413 (N_39413,N_35811,N_37487);
nand U39414 (N_39414,N_37093,N_35600);
and U39415 (N_39415,N_35397,N_35271);
nor U39416 (N_39416,N_36318,N_35038);
and U39417 (N_39417,N_35248,N_36798);
or U39418 (N_39418,N_36486,N_37203);
and U39419 (N_39419,N_36386,N_37303);
xor U39420 (N_39420,N_37226,N_37097);
and U39421 (N_39421,N_36980,N_36498);
nor U39422 (N_39422,N_36200,N_36905);
or U39423 (N_39423,N_36410,N_35581);
xor U39424 (N_39424,N_35232,N_35986);
and U39425 (N_39425,N_37170,N_35414);
nor U39426 (N_39426,N_35858,N_37366);
xnor U39427 (N_39427,N_36157,N_37119);
and U39428 (N_39428,N_36374,N_37281);
nor U39429 (N_39429,N_36220,N_35120);
and U39430 (N_39430,N_36200,N_35594);
or U39431 (N_39431,N_36060,N_37369);
xnor U39432 (N_39432,N_37497,N_36159);
xor U39433 (N_39433,N_37019,N_37283);
or U39434 (N_39434,N_35898,N_36602);
or U39435 (N_39435,N_35188,N_35596);
and U39436 (N_39436,N_36082,N_35004);
nand U39437 (N_39437,N_35879,N_37151);
nor U39438 (N_39438,N_37069,N_36757);
nand U39439 (N_39439,N_36910,N_35784);
or U39440 (N_39440,N_36174,N_35362);
and U39441 (N_39441,N_36305,N_36190);
and U39442 (N_39442,N_35660,N_37240);
nor U39443 (N_39443,N_35030,N_37279);
nand U39444 (N_39444,N_36593,N_35192);
nand U39445 (N_39445,N_37138,N_36441);
and U39446 (N_39446,N_35750,N_37403);
nor U39447 (N_39447,N_35335,N_36203);
nand U39448 (N_39448,N_36682,N_36104);
and U39449 (N_39449,N_35110,N_35560);
nor U39450 (N_39450,N_35860,N_37347);
xnor U39451 (N_39451,N_36753,N_35295);
or U39452 (N_39452,N_35779,N_36625);
xnor U39453 (N_39453,N_35257,N_35685);
nor U39454 (N_39454,N_37483,N_37377);
nand U39455 (N_39455,N_36409,N_35116);
nand U39456 (N_39456,N_36631,N_35448);
xor U39457 (N_39457,N_35230,N_37439);
nand U39458 (N_39458,N_37352,N_35449);
nor U39459 (N_39459,N_36211,N_37350);
or U39460 (N_39460,N_35949,N_36161);
nand U39461 (N_39461,N_37095,N_36172);
nor U39462 (N_39462,N_37263,N_36683);
and U39463 (N_39463,N_35475,N_36617);
nand U39464 (N_39464,N_36681,N_37333);
xor U39465 (N_39465,N_36062,N_36025);
nand U39466 (N_39466,N_36475,N_36074);
and U39467 (N_39467,N_37483,N_36019);
nand U39468 (N_39468,N_36546,N_36184);
and U39469 (N_39469,N_35894,N_36572);
or U39470 (N_39470,N_36579,N_35539);
nor U39471 (N_39471,N_35021,N_36335);
or U39472 (N_39472,N_35839,N_35683);
xor U39473 (N_39473,N_35926,N_35290);
and U39474 (N_39474,N_35553,N_35952);
and U39475 (N_39475,N_35536,N_35081);
nand U39476 (N_39476,N_36751,N_35979);
xnor U39477 (N_39477,N_35162,N_36390);
xor U39478 (N_39478,N_35185,N_36980);
and U39479 (N_39479,N_36890,N_36432);
and U39480 (N_39480,N_37101,N_35790);
nor U39481 (N_39481,N_35143,N_36026);
xor U39482 (N_39482,N_35513,N_35963);
xnor U39483 (N_39483,N_36615,N_35415);
and U39484 (N_39484,N_36322,N_35092);
and U39485 (N_39485,N_37109,N_36883);
nand U39486 (N_39486,N_36313,N_37453);
or U39487 (N_39487,N_35233,N_36390);
nor U39488 (N_39488,N_35275,N_36196);
xor U39489 (N_39489,N_35186,N_37406);
and U39490 (N_39490,N_37003,N_35150);
and U39491 (N_39491,N_37115,N_36972);
nand U39492 (N_39492,N_37298,N_35955);
nor U39493 (N_39493,N_36320,N_35767);
nand U39494 (N_39494,N_35685,N_37221);
xnor U39495 (N_39495,N_36339,N_37365);
and U39496 (N_39496,N_36768,N_37109);
xor U39497 (N_39497,N_35718,N_36824);
or U39498 (N_39498,N_35882,N_37125);
nor U39499 (N_39499,N_35967,N_36438);
nor U39500 (N_39500,N_36872,N_37291);
and U39501 (N_39501,N_37403,N_37416);
nand U39502 (N_39502,N_37281,N_35739);
xor U39503 (N_39503,N_36892,N_35627);
or U39504 (N_39504,N_35766,N_36527);
nor U39505 (N_39505,N_35623,N_35914);
and U39506 (N_39506,N_36576,N_36049);
xor U39507 (N_39507,N_35089,N_37261);
and U39508 (N_39508,N_35181,N_37472);
or U39509 (N_39509,N_36820,N_36291);
or U39510 (N_39510,N_36946,N_35195);
and U39511 (N_39511,N_35928,N_37480);
or U39512 (N_39512,N_35474,N_35446);
or U39513 (N_39513,N_35798,N_35990);
nand U39514 (N_39514,N_35598,N_35723);
nand U39515 (N_39515,N_36631,N_35528);
and U39516 (N_39516,N_35843,N_35883);
nor U39517 (N_39517,N_35932,N_37062);
or U39518 (N_39518,N_35904,N_37480);
xnor U39519 (N_39519,N_35876,N_35281);
xor U39520 (N_39520,N_35260,N_35939);
or U39521 (N_39521,N_36339,N_35430);
and U39522 (N_39522,N_35251,N_35535);
nor U39523 (N_39523,N_37252,N_36068);
and U39524 (N_39524,N_36112,N_35621);
xnor U39525 (N_39525,N_36442,N_37465);
xor U39526 (N_39526,N_36845,N_37405);
nand U39527 (N_39527,N_35682,N_36345);
nor U39528 (N_39528,N_35403,N_36199);
and U39529 (N_39529,N_36110,N_37094);
nor U39530 (N_39530,N_35665,N_36709);
or U39531 (N_39531,N_35472,N_36441);
xor U39532 (N_39532,N_35484,N_37011);
or U39533 (N_39533,N_35810,N_35644);
and U39534 (N_39534,N_37399,N_37357);
nor U39535 (N_39535,N_35162,N_37194);
xor U39536 (N_39536,N_36408,N_36658);
xor U39537 (N_39537,N_36234,N_36424);
or U39538 (N_39538,N_36177,N_35824);
or U39539 (N_39539,N_35205,N_36894);
or U39540 (N_39540,N_36536,N_37345);
and U39541 (N_39541,N_35447,N_36722);
and U39542 (N_39542,N_37002,N_37051);
nand U39543 (N_39543,N_35859,N_36829);
or U39544 (N_39544,N_35275,N_36997);
or U39545 (N_39545,N_35471,N_35425);
and U39546 (N_39546,N_35309,N_35024);
or U39547 (N_39547,N_37252,N_37457);
and U39548 (N_39548,N_35993,N_36574);
nor U39549 (N_39549,N_36664,N_35715);
or U39550 (N_39550,N_36205,N_36814);
xnor U39551 (N_39551,N_36036,N_35213);
or U39552 (N_39552,N_36396,N_37261);
or U39553 (N_39553,N_37098,N_35352);
nand U39554 (N_39554,N_36573,N_36444);
and U39555 (N_39555,N_36619,N_36222);
or U39556 (N_39556,N_36528,N_35422);
or U39557 (N_39557,N_36390,N_35681);
nor U39558 (N_39558,N_37102,N_37369);
nand U39559 (N_39559,N_35483,N_37076);
xor U39560 (N_39560,N_35904,N_36714);
or U39561 (N_39561,N_36919,N_35202);
or U39562 (N_39562,N_37094,N_37238);
xnor U39563 (N_39563,N_35338,N_35555);
nor U39564 (N_39564,N_35058,N_35857);
or U39565 (N_39565,N_35672,N_36360);
nor U39566 (N_39566,N_36763,N_35758);
nand U39567 (N_39567,N_37437,N_35916);
nand U39568 (N_39568,N_35567,N_36579);
or U39569 (N_39569,N_35298,N_36959);
and U39570 (N_39570,N_35075,N_36922);
and U39571 (N_39571,N_36243,N_36033);
nand U39572 (N_39572,N_36733,N_35297);
or U39573 (N_39573,N_36124,N_35290);
xor U39574 (N_39574,N_37054,N_35277);
nand U39575 (N_39575,N_35559,N_36554);
xor U39576 (N_39576,N_35876,N_35247);
nand U39577 (N_39577,N_36659,N_36445);
and U39578 (N_39578,N_35744,N_37107);
xor U39579 (N_39579,N_35905,N_36645);
xor U39580 (N_39580,N_35132,N_36875);
nor U39581 (N_39581,N_35927,N_37147);
nor U39582 (N_39582,N_37126,N_35708);
nand U39583 (N_39583,N_35702,N_37055);
xor U39584 (N_39584,N_35140,N_36590);
nor U39585 (N_39585,N_35951,N_35752);
nor U39586 (N_39586,N_35016,N_36783);
or U39587 (N_39587,N_35947,N_37093);
nor U39588 (N_39588,N_35049,N_37078);
xor U39589 (N_39589,N_36985,N_36011);
nor U39590 (N_39590,N_35401,N_35028);
and U39591 (N_39591,N_35341,N_36024);
nand U39592 (N_39592,N_35457,N_35299);
and U39593 (N_39593,N_35665,N_35097);
nor U39594 (N_39594,N_36707,N_37219);
nand U39595 (N_39595,N_35228,N_37368);
nor U39596 (N_39596,N_35190,N_36028);
or U39597 (N_39597,N_36690,N_35970);
or U39598 (N_39598,N_35652,N_37369);
nor U39599 (N_39599,N_35629,N_36476);
or U39600 (N_39600,N_35607,N_36890);
nor U39601 (N_39601,N_35466,N_35930);
nor U39602 (N_39602,N_35496,N_35901);
xor U39603 (N_39603,N_35683,N_35644);
or U39604 (N_39604,N_37361,N_36593);
or U39605 (N_39605,N_36485,N_36507);
xor U39606 (N_39606,N_37037,N_35426);
nor U39607 (N_39607,N_36501,N_36688);
or U39608 (N_39608,N_35397,N_37041);
nor U39609 (N_39609,N_36641,N_35499);
and U39610 (N_39610,N_35164,N_36461);
nor U39611 (N_39611,N_35914,N_37263);
and U39612 (N_39612,N_37002,N_35291);
xnor U39613 (N_39613,N_35283,N_36582);
xnor U39614 (N_39614,N_37325,N_37349);
xor U39615 (N_39615,N_36130,N_37484);
and U39616 (N_39616,N_36964,N_37187);
and U39617 (N_39617,N_36146,N_37238);
and U39618 (N_39618,N_36854,N_35070);
or U39619 (N_39619,N_35197,N_36933);
or U39620 (N_39620,N_35204,N_37142);
xor U39621 (N_39621,N_36610,N_36862);
xor U39622 (N_39622,N_35987,N_36981);
and U39623 (N_39623,N_36537,N_35609);
nor U39624 (N_39624,N_37295,N_35055);
and U39625 (N_39625,N_36688,N_35252);
nor U39626 (N_39626,N_36330,N_35742);
and U39627 (N_39627,N_35133,N_36010);
nor U39628 (N_39628,N_35139,N_36930);
xor U39629 (N_39629,N_35857,N_36554);
or U39630 (N_39630,N_35201,N_35597);
xor U39631 (N_39631,N_36921,N_37204);
nand U39632 (N_39632,N_35560,N_36553);
and U39633 (N_39633,N_36034,N_36961);
and U39634 (N_39634,N_37213,N_36845);
and U39635 (N_39635,N_36790,N_36609);
and U39636 (N_39636,N_35784,N_35162);
nor U39637 (N_39637,N_36962,N_36137);
or U39638 (N_39638,N_35133,N_35735);
and U39639 (N_39639,N_36114,N_36778);
nor U39640 (N_39640,N_36422,N_36460);
nand U39641 (N_39641,N_37357,N_35910);
nand U39642 (N_39642,N_35931,N_35425);
nor U39643 (N_39643,N_37076,N_36085);
nor U39644 (N_39644,N_37231,N_36450);
nand U39645 (N_39645,N_35743,N_36317);
or U39646 (N_39646,N_35294,N_35113);
nor U39647 (N_39647,N_37430,N_35528);
xnor U39648 (N_39648,N_36512,N_35172);
and U39649 (N_39649,N_36593,N_37343);
nor U39650 (N_39650,N_35104,N_35935);
nor U39651 (N_39651,N_36070,N_36996);
xor U39652 (N_39652,N_36230,N_37017);
or U39653 (N_39653,N_35233,N_35311);
nand U39654 (N_39654,N_36526,N_36578);
or U39655 (N_39655,N_37027,N_36273);
and U39656 (N_39656,N_36298,N_35824);
nor U39657 (N_39657,N_36117,N_36719);
or U39658 (N_39658,N_35682,N_35951);
nand U39659 (N_39659,N_35947,N_37000);
xnor U39660 (N_39660,N_35082,N_36559);
nor U39661 (N_39661,N_35916,N_36107);
xnor U39662 (N_39662,N_37448,N_35747);
or U39663 (N_39663,N_36723,N_37490);
or U39664 (N_39664,N_35574,N_35272);
or U39665 (N_39665,N_35315,N_36762);
nand U39666 (N_39666,N_36383,N_36669);
and U39667 (N_39667,N_35441,N_37356);
and U39668 (N_39668,N_35535,N_35240);
xnor U39669 (N_39669,N_35336,N_37228);
or U39670 (N_39670,N_35368,N_36626);
nand U39671 (N_39671,N_36761,N_35712);
nor U39672 (N_39672,N_35373,N_35891);
nand U39673 (N_39673,N_37284,N_37148);
xor U39674 (N_39674,N_35020,N_35047);
xnor U39675 (N_39675,N_35406,N_35554);
nand U39676 (N_39676,N_35607,N_35104);
xor U39677 (N_39677,N_36937,N_35120);
xor U39678 (N_39678,N_37258,N_36858);
xnor U39679 (N_39679,N_35640,N_35681);
or U39680 (N_39680,N_35476,N_36109);
nand U39681 (N_39681,N_35390,N_35949);
or U39682 (N_39682,N_36495,N_37016);
or U39683 (N_39683,N_35982,N_36130);
xnor U39684 (N_39684,N_36763,N_35918);
nand U39685 (N_39685,N_35096,N_35673);
nor U39686 (N_39686,N_35524,N_36946);
or U39687 (N_39687,N_37025,N_36709);
nand U39688 (N_39688,N_37157,N_35897);
or U39689 (N_39689,N_35388,N_37198);
and U39690 (N_39690,N_35173,N_36178);
or U39691 (N_39691,N_35502,N_35942);
xnor U39692 (N_39692,N_36719,N_35510);
nor U39693 (N_39693,N_36870,N_36177);
nor U39694 (N_39694,N_35396,N_35040);
nor U39695 (N_39695,N_35819,N_35846);
nor U39696 (N_39696,N_36825,N_36706);
xor U39697 (N_39697,N_37214,N_35929);
or U39698 (N_39698,N_36305,N_35310);
and U39699 (N_39699,N_36618,N_35722);
nand U39700 (N_39700,N_36597,N_35046);
xnor U39701 (N_39701,N_36625,N_37158);
or U39702 (N_39702,N_36404,N_36810);
or U39703 (N_39703,N_36708,N_35687);
or U39704 (N_39704,N_36961,N_36968);
nand U39705 (N_39705,N_35373,N_36899);
xnor U39706 (N_39706,N_35292,N_35756);
or U39707 (N_39707,N_35562,N_36539);
nand U39708 (N_39708,N_35002,N_35494);
xnor U39709 (N_39709,N_35514,N_37115);
nand U39710 (N_39710,N_36709,N_35305);
nand U39711 (N_39711,N_35134,N_36773);
xnor U39712 (N_39712,N_35371,N_35198);
or U39713 (N_39713,N_37041,N_36214);
nand U39714 (N_39714,N_36044,N_35276);
nor U39715 (N_39715,N_37093,N_35551);
xnor U39716 (N_39716,N_36665,N_36351);
nor U39717 (N_39717,N_36007,N_35608);
and U39718 (N_39718,N_35277,N_35834);
and U39719 (N_39719,N_36803,N_36762);
xor U39720 (N_39720,N_37005,N_35079);
or U39721 (N_39721,N_36500,N_37173);
or U39722 (N_39722,N_36230,N_35092);
xnor U39723 (N_39723,N_35226,N_36818);
or U39724 (N_39724,N_35002,N_35273);
or U39725 (N_39725,N_36926,N_36799);
and U39726 (N_39726,N_36248,N_37452);
and U39727 (N_39727,N_36907,N_35940);
nor U39728 (N_39728,N_37058,N_35559);
nand U39729 (N_39729,N_35864,N_37184);
xnor U39730 (N_39730,N_36656,N_37201);
nor U39731 (N_39731,N_35026,N_37314);
nor U39732 (N_39732,N_36100,N_35443);
nand U39733 (N_39733,N_36385,N_36076);
nor U39734 (N_39734,N_36209,N_37495);
xnor U39735 (N_39735,N_36039,N_36006);
xor U39736 (N_39736,N_35692,N_36033);
nand U39737 (N_39737,N_35850,N_37224);
nand U39738 (N_39738,N_35679,N_37336);
nor U39739 (N_39739,N_35314,N_37204);
nor U39740 (N_39740,N_36576,N_36973);
xnor U39741 (N_39741,N_37238,N_35762);
nor U39742 (N_39742,N_36870,N_35674);
xnor U39743 (N_39743,N_36514,N_35881);
nor U39744 (N_39744,N_35456,N_35689);
nand U39745 (N_39745,N_35775,N_37363);
xnor U39746 (N_39746,N_36296,N_36735);
or U39747 (N_39747,N_36464,N_35024);
nand U39748 (N_39748,N_36584,N_36666);
and U39749 (N_39749,N_36207,N_36317);
and U39750 (N_39750,N_36490,N_36635);
nand U39751 (N_39751,N_35871,N_35119);
or U39752 (N_39752,N_37474,N_36644);
or U39753 (N_39753,N_35466,N_35980);
xor U39754 (N_39754,N_35165,N_36004);
nor U39755 (N_39755,N_36795,N_35910);
xor U39756 (N_39756,N_37281,N_36605);
nand U39757 (N_39757,N_36141,N_36906);
or U39758 (N_39758,N_36676,N_37459);
xor U39759 (N_39759,N_36365,N_35651);
or U39760 (N_39760,N_35907,N_36783);
and U39761 (N_39761,N_35134,N_36692);
and U39762 (N_39762,N_37319,N_35839);
and U39763 (N_39763,N_37495,N_37059);
or U39764 (N_39764,N_37147,N_36763);
or U39765 (N_39765,N_35311,N_37423);
or U39766 (N_39766,N_35900,N_36200);
and U39767 (N_39767,N_37170,N_36652);
and U39768 (N_39768,N_36120,N_35931);
xnor U39769 (N_39769,N_36085,N_37258);
and U39770 (N_39770,N_37286,N_36056);
xor U39771 (N_39771,N_36008,N_37394);
and U39772 (N_39772,N_36429,N_36212);
nand U39773 (N_39773,N_36286,N_36157);
nand U39774 (N_39774,N_37162,N_36080);
or U39775 (N_39775,N_36793,N_35286);
nand U39776 (N_39776,N_35199,N_35791);
and U39777 (N_39777,N_36043,N_36319);
and U39778 (N_39778,N_36900,N_35958);
and U39779 (N_39779,N_35143,N_36732);
or U39780 (N_39780,N_35480,N_37064);
and U39781 (N_39781,N_35937,N_36878);
nand U39782 (N_39782,N_36539,N_36179);
nor U39783 (N_39783,N_36247,N_36902);
nor U39784 (N_39784,N_35856,N_37114);
nand U39785 (N_39785,N_36707,N_37191);
nand U39786 (N_39786,N_36964,N_36124);
or U39787 (N_39787,N_36317,N_35886);
nand U39788 (N_39788,N_36417,N_37314);
xnor U39789 (N_39789,N_35638,N_36690);
nor U39790 (N_39790,N_37167,N_37037);
nor U39791 (N_39791,N_36895,N_35505);
and U39792 (N_39792,N_35421,N_37181);
nor U39793 (N_39793,N_36072,N_35181);
and U39794 (N_39794,N_37386,N_36512);
nand U39795 (N_39795,N_36695,N_35955);
nor U39796 (N_39796,N_35974,N_35878);
nor U39797 (N_39797,N_36480,N_36251);
xnor U39798 (N_39798,N_36767,N_35025);
nor U39799 (N_39799,N_37314,N_37191);
nand U39800 (N_39800,N_36955,N_36113);
nor U39801 (N_39801,N_36231,N_37259);
nand U39802 (N_39802,N_37217,N_36710);
or U39803 (N_39803,N_35130,N_36493);
xnor U39804 (N_39804,N_35470,N_35525);
nor U39805 (N_39805,N_36205,N_37024);
and U39806 (N_39806,N_36463,N_35929);
or U39807 (N_39807,N_36047,N_37076);
or U39808 (N_39808,N_37209,N_36515);
or U39809 (N_39809,N_36011,N_35229);
and U39810 (N_39810,N_35413,N_37332);
nor U39811 (N_39811,N_35763,N_36659);
and U39812 (N_39812,N_35249,N_37415);
and U39813 (N_39813,N_35595,N_36720);
or U39814 (N_39814,N_35633,N_37225);
xor U39815 (N_39815,N_35902,N_35623);
xnor U39816 (N_39816,N_36043,N_35766);
or U39817 (N_39817,N_37472,N_35133);
xnor U39818 (N_39818,N_36211,N_37332);
or U39819 (N_39819,N_35681,N_35987);
nand U39820 (N_39820,N_36875,N_36870);
xor U39821 (N_39821,N_36734,N_35831);
and U39822 (N_39822,N_35497,N_35095);
or U39823 (N_39823,N_36331,N_37224);
or U39824 (N_39824,N_36205,N_35320);
and U39825 (N_39825,N_36202,N_35305);
or U39826 (N_39826,N_35685,N_36432);
or U39827 (N_39827,N_37148,N_36239);
nand U39828 (N_39828,N_36629,N_35446);
and U39829 (N_39829,N_36467,N_35447);
or U39830 (N_39830,N_36855,N_37138);
nor U39831 (N_39831,N_35962,N_37318);
nor U39832 (N_39832,N_36934,N_35213);
xnor U39833 (N_39833,N_35177,N_36435);
nor U39834 (N_39834,N_36305,N_36551);
or U39835 (N_39835,N_35609,N_36124);
nand U39836 (N_39836,N_36839,N_37485);
xor U39837 (N_39837,N_36208,N_35493);
and U39838 (N_39838,N_36429,N_37108);
nand U39839 (N_39839,N_35634,N_35162);
and U39840 (N_39840,N_37232,N_35664);
or U39841 (N_39841,N_37100,N_36995);
and U39842 (N_39842,N_36698,N_35011);
nand U39843 (N_39843,N_35474,N_35914);
and U39844 (N_39844,N_36369,N_35775);
nor U39845 (N_39845,N_36340,N_35270);
and U39846 (N_39846,N_36676,N_37489);
and U39847 (N_39847,N_36137,N_35992);
nand U39848 (N_39848,N_35117,N_36473);
nand U39849 (N_39849,N_37069,N_35523);
nand U39850 (N_39850,N_35298,N_37163);
xnor U39851 (N_39851,N_35893,N_37003);
xnor U39852 (N_39852,N_36123,N_36051);
nor U39853 (N_39853,N_35590,N_35019);
and U39854 (N_39854,N_36496,N_37081);
or U39855 (N_39855,N_36646,N_37137);
nand U39856 (N_39856,N_36643,N_37256);
and U39857 (N_39857,N_37490,N_37493);
nand U39858 (N_39858,N_35592,N_37490);
xnor U39859 (N_39859,N_36767,N_36343);
or U39860 (N_39860,N_36753,N_35482);
nand U39861 (N_39861,N_35329,N_36123);
xnor U39862 (N_39862,N_36342,N_35709);
xor U39863 (N_39863,N_35098,N_35235);
xor U39864 (N_39864,N_35985,N_36654);
and U39865 (N_39865,N_36299,N_35208);
xor U39866 (N_39866,N_35394,N_36975);
and U39867 (N_39867,N_35830,N_36692);
xnor U39868 (N_39868,N_35321,N_35569);
and U39869 (N_39869,N_35313,N_37006);
or U39870 (N_39870,N_36681,N_37421);
nand U39871 (N_39871,N_36582,N_35747);
or U39872 (N_39872,N_35052,N_36839);
xor U39873 (N_39873,N_37022,N_37283);
nand U39874 (N_39874,N_36008,N_36473);
or U39875 (N_39875,N_35186,N_36898);
nand U39876 (N_39876,N_37337,N_36360);
and U39877 (N_39877,N_36639,N_35868);
nor U39878 (N_39878,N_35593,N_36172);
or U39879 (N_39879,N_37105,N_35800);
and U39880 (N_39880,N_37489,N_36356);
and U39881 (N_39881,N_37056,N_36922);
nand U39882 (N_39882,N_35483,N_35413);
and U39883 (N_39883,N_35411,N_36775);
xor U39884 (N_39884,N_36150,N_36831);
or U39885 (N_39885,N_37466,N_36459);
nand U39886 (N_39886,N_37481,N_35828);
nor U39887 (N_39887,N_35386,N_35937);
or U39888 (N_39888,N_37284,N_35437);
and U39889 (N_39889,N_36629,N_36272);
nor U39890 (N_39890,N_35967,N_37272);
nor U39891 (N_39891,N_35765,N_36548);
or U39892 (N_39892,N_36877,N_35228);
or U39893 (N_39893,N_37420,N_35197);
xor U39894 (N_39894,N_35933,N_35699);
xor U39895 (N_39895,N_35995,N_37284);
nor U39896 (N_39896,N_37309,N_37265);
or U39897 (N_39897,N_36457,N_36667);
or U39898 (N_39898,N_37143,N_35353);
and U39899 (N_39899,N_35382,N_35725);
and U39900 (N_39900,N_35241,N_37345);
xnor U39901 (N_39901,N_36740,N_35352);
or U39902 (N_39902,N_36569,N_35605);
or U39903 (N_39903,N_36004,N_35734);
or U39904 (N_39904,N_35133,N_37363);
or U39905 (N_39905,N_35096,N_36810);
nor U39906 (N_39906,N_35557,N_35007);
and U39907 (N_39907,N_35286,N_36609);
and U39908 (N_39908,N_36377,N_35894);
or U39909 (N_39909,N_37055,N_36566);
nor U39910 (N_39910,N_35234,N_36913);
nor U39911 (N_39911,N_36274,N_37346);
nand U39912 (N_39912,N_36801,N_35093);
nor U39913 (N_39913,N_35879,N_35851);
nand U39914 (N_39914,N_35066,N_35850);
nand U39915 (N_39915,N_36048,N_36901);
xor U39916 (N_39916,N_36258,N_37172);
xor U39917 (N_39917,N_36938,N_36961);
or U39918 (N_39918,N_36192,N_36024);
and U39919 (N_39919,N_36761,N_35879);
or U39920 (N_39920,N_36036,N_36904);
or U39921 (N_39921,N_35873,N_35899);
or U39922 (N_39922,N_36454,N_37359);
or U39923 (N_39923,N_37031,N_36608);
nor U39924 (N_39924,N_37491,N_37086);
and U39925 (N_39925,N_35563,N_37049);
nand U39926 (N_39926,N_36789,N_35707);
and U39927 (N_39927,N_35107,N_35900);
and U39928 (N_39928,N_35049,N_36488);
or U39929 (N_39929,N_35577,N_37257);
nor U39930 (N_39930,N_36567,N_37352);
nand U39931 (N_39931,N_36661,N_37053);
nor U39932 (N_39932,N_35180,N_35109);
or U39933 (N_39933,N_37221,N_35377);
and U39934 (N_39934,N_36269,N_36165);
xnor U39935 (N_39935,N_36793,N_36512);
nand U39936 (N_39936,N_36788,N_36297);
nand U39937 (N_39937,N_36286,N_35833);
or U39938 (N_39938,N_36135,N_37046);
nand U39939 (N_39939,N_37231,N_36453);
nor U39940 (N_39940,N_36327,N_35794);
xnor U39941 (N_39941,N_35604,N_36010);
nor U39942 (N_39942,N_35830,N_35581);
nor U39943 (N_39943,N_35704,N_37307);
nand U39944 (N_39944,N_36976,N_37032);
and U39945 (N_39945,N_36052,N_37358);
nand U39946 (N_39946,N_35303,N_35378);
and U39947 (N_39947,N_37000,N_35624);
and U39948 (N_39948,N_35539,N_36644);
or U39949 (N_39949,N_36889,N_37090);
nor U39950 (N_39950,N_35842,N_35039);
or U39951 (N_39951,N_36737,N_37061);
or U39952 (N_39952,N_36891,N_35893);
nor U39953 (N_39953,N_35944,N_36794);
nor U39954 (N_39954,N_35251,N_35741);
xor U39955 (N_39955,N_37076,N_35838);
nor U39956 (N_39956,N_35184,N_36394);
xnor U39957 (N_39957,N_35276,N_37233);
and U39958 (N_39958,N_36274,N_36157);
and U39959 (N_39959,N_36442,N_35183);
nor U39960 (N_39960,N_35171,N_37433);
nand U39961 (N_39961,N_35437,N_35098);
nor U39962 (N_39962,N_36217,N_36092);
and U39963 (N_39963,N_35561,N_35222);
nor U39964 (N_39964,N_37311,N_35922);
xnor U39965 (N_39965,N_36871,N_35652);
and U39966 (N_39966,N_36203,N_35428);
or U39967 (N_39967,N_36041,N_36652);
or U39968 (N_39968,N_36176,N_36605);
nand U39969 (N_39969,N_35445,N_36791);
and U39970 (N_39970,N_35994,N_35725);
and U39971 (N_39971,N_35644,N_37252);
or U39972 (N_39972,N_35813,N_36045);
xnor U39973 (N_39973,N_37228,N_36586);
xor U39974 (N_39974,N_36248,N_36975);
xor U39975 (N_39975,N_35106,N_36922);
or U39976 (N_39976,N_35272,N_37453);
nand U39977 (N_39977,N_35853,N_37013);
or U39978 (N_39978,N_35601,N_36759);
nor U39979 (N_39979,N_35191,N_37298);
xnor U39980 (N_39980,N_36128,N_35268);
nand U39981 (N_39981,N_35371,N_36420);
xnor U39982 (N_39982,N_35084,N_36024);
and U39983 (N_39983,N_36723,N_36872);
and U39984 (N_39984,N_35410,N_36407);
nand U39985 (N_39985,N_35621,N_35596);
and U39986 (N_39986,N_35589,N_35005);
and U39987 (N_39987,N_37059,N_35402);
or U39988 (N_39988,N_36641,N_37208);
nor U39989 (N_39989,N_37075,N_37378);
or U39990 (N_39990,N_36419,N_37105);
or U39991 (N_39991,N_36137,N_36187);
or U39992 (N_39992,N_35733,N_35271);
xor U39993 (N_39993,N_36885,N_36643);
or U39994 (N_39994,N_35123,N_35474);
and U39995 (N_39995,N_36745,N_36769);
or U39996 (N_39996,N_36197,N_37438);
and U39997 (N_39997,N_36623,N_35132);
or U39998 (N_39998,N_37197,N_36821);
xnor U39999 (N_39999,N_36867,N_36151);
or U40000 (N_40000,N_39658,N_39492);
nor U40001 (N_40001,N_38392,N_38545);
xnor U40002 (N_40002,N_38628,N_38222);
xor U40003 (N_40003,N_37720,N_38174);
nand U40004 (N_40004,N_37710,N_38340);
xnor U40005 (N_40005,N_37579,N_38923);
xnor U40006 (N_40006,N_37566,N_39606);
nor U40007 (N_40007,N_39478,N_39795);
nor U40008 (N_40008,N_39910,N_38091);
xor U40009 (N_40009,N_39394,N_38033);
nor U40010 (N_40010,N_38067,N_39716);
and U40011 (N_40011,N_38488,N_39757);
and U40012 (N_40012,N_37687,N_38990);
nor U40013 (N_40013,N_38900,N_38560);
nand U40014 (N_40014,N_38283,N_39898);
nand U40015 (N_40015,N_39413,N_39599);
nor U40016 (N_40016,N_38087,N_37778);
or U40017 (N_40017,N_39450,N_39653);
and U40018 (N_40018,N_38913,N_39887);
nor U40019 (N_40019,N_37931,N_38757);
or U40020 (N_40020,N_37986,N_38133);
or U40021 (N_40021,N_38548,N_39356);
or U40022 (N_40022,N_38458,N_39252);
or U40023 (N_40023,N_39392,N_38664);
nand U40024 (N_40024,N_38636,N_39342);
or U40025 (N_40025,N_39626,N_37998);
nor U40026 (N_40026,N_38866,N_37633);
and U40027 (N_40027,N_38165,N_39050);
nand U40028 (N_40028,N_37671,N_39748);
and U40029 (N_40029,N_38865,N_38371);
or U40030 (N_40030,N_39837,N_39359);
nand U40031 (N_40031,N_38857,N_39473);
xor U40032 (N_40032,N_39860,N_39945);
or U40033 (N_40033,N_39045,N_38201);
nand U40034 (N_40034,N_38104,N_39520);
and U40035 (N_40035,N_38424,N_37829);
or U40036 (N_40036,N_38350,N_37532);
or U40037 (N_40037,N_39237,N_37718);
or U40038 (N_40038,N_38893,N_38423);
xor U40039 (N_40039,N_37902,N_39499);
nand U40040 (N_40040,N_39210,N_39244);
xnor U40041 (N_40041,N_37760,N_38403);
nand U40042 (N_40042,N_38836,N_37933);
or U40043 (N_40043,N_38247,N_38177);
or U40044 (N_40044,N_39659,N_38998);
nand U40045 (N_40045,N_39463,N_39996);
or U40046 (N_40046,N_39515,N_39440);
nor U40047 (N_40047,N_39650,N_38784);
xnor U40048 (N_40048,N_39209,N_39435);
and U40049 (N_40049,N_39211,N_39309);
and U40050 (N_40050,N_39215,N_39028);
and U40051 (N_40051,N_37582,N_39416);
xor U40052 (N_40052,N_38872,N_38566);
or U40053 (N_40053,N_39551,N_38541);
nor U40054 (N_40054,N_39691,N_38270);
nand U40055 (N_40055,N_38769,N_37969);
nand U40056 (N_40056,N_38236,N_39897);
or U40057 (N_40057,N_39605,N_38150);
or U40058 (N_40058,N_39567,N_38980);
xnor U40059 (N_40059,N_38941,N_38504);
or U40060 (N_40060,N_38610,N_39547);
or U40061 (N_40061,N_39445,N_38513);
nor U40062 (N_40062,N_39343,N_39673);
nor U40063 (N_40063,N_37715,N_39365);
xnor U40064 (N_40064,N_37682,N_38927);
or U40065 (N_40065,N_39302,N_39339);
and U40066 (N_40066,N_38699,N_37606);
and U40067 (N_40067,N_38019,N_39188);
xor U40068 (N_40068,N_39806,N_38224);
nand U40069 (N_40069,N_39946,N_39881);
and U40070 (N_40070,N_38249,N_38752);
or U40071 (N_40071,N_37843,N_38554);
nand U40072 (N_40072,N_38729,N_39808);
xnor U40073 (N_40073,N_38844,N_39006);
nand U40074 (N_40074,N_38799,N_39337);
and U40075 (N_40075,N_39190,N_37514);
or U40076 (N_40076,N_39151,N_37925);
and U40077 (N_40077,N_37573,N_39651);
nand U40078 (N_40078,N_39744,N_38715);
xor U40079 (N_40079,N_38653,N_39117);
nand U40080 (N_40080,N_38321,N_39617);
or U40081 (N_40081,N_37636,N_38598);
nor U40082 (N_40082,N_39348,N_39448);
or U40083 (N_40083,N_38074,N_38849);
or U40084 (N_40084,N_37714,N_38027);
or U40085 (N_40085,N_39715,N_38617);
nor U40086 (N_40086,N_38240,N_38968);
nand U40087 (N_40087,N_39130,N_38470);
nor U40088 (N_40088,N_38669,N_38670);
xnor U40089 (N_40089,N_38852,N_39310);
and U40090 (N_40090,N_38901,N_38446);
xnor U40091 (N_40091,N_39055,N_38188);
nand U40092 (N_40092,N_38271,N_39402);
nor U40093 (N_40093,N_37534,N_38035);
nor U40094 (N_40094,N_39294,N_38805);
nor U40095 (N_40095,N_37736,N_37592);
xor U40096 (N_40096,N_39568,N_38313);
nand U40097 (N_40097,N_37975,N_38395);
xor U40098 (N_40098,N_37645,N_39457);
nor U40099 (N_40099,N_38544,N_38838);
or U40100 (N_40100,N_37765,N_37782);
and U40101 (N_40101,N_39851,N_37820);
nand U40102 (N_40102,N_37813,N_39307);
or U40103 (N_40103,N_37670,N_39723);
or U40104 (N_40104,N_39792,N_39060);
nand U40105 (N_40105,N_39886,N_38832);
and U40106 (N_40106,N_38023,N_38348);
nor U40107 (N_40107,N_37917,N_39855);
xor U40108 (N_40108,N_39951,N_39289);
or U40109 (N_40109,N_39238,N_37656);
nor U40110 (N_40110,N_37919,N_38984);
xor U40111 (N_40111,N_37945,N_39364);
xor U40112 (N_40112,N_39104,N_37865);
nand U40113 (N_40113,N_37642,N_38791);
and U40114 (N_40114,N_38562,N_39236);
xor U40115 (N_40115,N_38237,N_39012);
nand U40116 (N_40116,N_37801,N_37836);
and U40117 (N_40117,N_38793,N_37673);
nor U40118 (N_40118,N_38971,N_39122);
xor U40119 (N_40119,N_39720,N_39818);
nand U40120 (N_40120,N_39826,N_39193);
xnor U40121 (N_40121,N_39304,N_39553);
and U40122 (N_40122,N_39760,N_37587);
xnor U40123 (N_40123,N_37841,N_38555);
nor U40124 (N_40124,N_37542,N_39220);
and U40125 (N_40125,N_39379,N_38435);
xor U40126 (N_40126,N_38894,N_38184);
nand U40127 (N_40127,N_38020,N_39021);
nor U40128 (N_40128,N_39517,N_38116);
nor U40129 (N_40129,N_39767,N_39506);
nor U40130 (N_40130,N_38462,N_38021);
xor U40131 (N_40131,N_38648,N_39692);
nor U40132 (N_40132,N_39374,N_39809);
or U40133 (N_40133,N_38641,N_39229);
and U40134 (N_40134,N_39195,N_38082);
or U40135 (N_40135,N_39769,N_39982);
or U40136 (N_40136,N_39277,N_38552);
nor U40137 (N_40137,N_38943,N_39109);
nand U40138 (N_40138,N_39166,N_39689);
nand U40139 (N_40139,N_38070,N_38029);
and U40140 (N_40140,N_39700,N_38268);
or U40141 (N_40141,N_39829,N_37802);
xor U40142 (N_40142,N_37515,N_39439);
or U40143 (N_40143,N_38471,N_38320);
xor U40144 (N_40144,N_39059,N_39418);
nand U40145 (N_40145,N_38198,N_39447);
or U40146 (N_40146,N_39846,N_39864);
or U40147 (N_40147,N_39636,N_37740);
nand U40148 (N_40148,N_39925,N_38703);
or U40149 (N_40149,N_38260,N_38101);
xor U40150 (N_40150,N_39172,N_38454);
xor U40151 (N_40151,N_38301,N_39027);
or U40152 (N_40152,N_38154,N_38486);
nor U40153 (N_40153,N_39766,N_38468);
nor U40154 (N_40154,N_38336,N_38556);
and U40155 (N_40155,N_39398,N_39273);
and U40156 (N_40156,N_39619,N_39528);
or U40157 (N_40157,N_39383,N_38863);
and U40158 (N_40158,N_39221,N_39679);
nor U40159 (N_40159,N_37701,N_39848);
xor U40160 (N_40160,N_38211,N_39604);
xnor U40161 (N_40161,N_38727,N_38064);
xnor U40162 (N_40162,N_39154,N_38692);
and U40163 (N_40163,N_38453,N_39591);
xnor U40164 (N_40164,N_38889,N_38508);
xnor U40165 (N_40165,N_38319,N_37822);
or U40166 (N_40166,N_37855,N_39942);
and U40167 (N_40167,N_39813,N_39751);
nand U40168 (N_40168,N_38032,N_39349);
xnor U40169 (N_40169,N_38449,N_39913);
nor U40170 (N_40170,N_39624,N_38627);
nor U40171 (N_40171,N_37767,N_39698);
or U40172 (N_40172,N_38906,N_39995);
xor U40173 (N_40173,N_37950,N_38952);
xor U40174 (N_40174,N_38025,N_38584);
xnor U40175 (N_40175,N_37674,N_39859);
and U40176 (N_40176,N_37614,N_37504);
xor U40177 (N_40177,N_38714,N_39836);
nor U40178 (N_40178,N_37814,N_38347);
xnor U40179 (N_40179,N_38948,N_39754);
nand U40180 (N_40180,N_39564,N_37992);
nor U40181 (N_40181,N_39361,N_37810);
or U40182 (N_40182,N_37681,N_39589);
xor U40183 (N_40183,N_37744,N_39977);
xor U40184 (N_40184,N_39889,N_38896);
xnor U40185 (N_40185,N_39969,N_38914);
or U40186 (N_40186,N_37797,N_39404);
nand U40187 (N_40187,N_38073,N_37733);
or U40188 (N_40188,N_39911,N_37994);
nor U40189 (N_40189,N_37659,N_39683);
xnor U40190 (N_40190,N_38719,N_38051);
nand U40191 (N_40191,N_38197,N_39733);
or U40192 (N_40192,N_38975,N_38772);
xnor U40193 (N_40193,N_39346,N_39372);
xnor U40194 (N_40194,N_37741,N_39271);
nor U40195 (N_40195,N_39150,N_38839);
and U40196 (N_40196,N_38926,N_38679);
and U40197 (N_40197,N_39742,N_38089);
and U40198 (N_40198,N_38044,N_38388);
xor U40199 (N_40199,N_39077,N_38352);
and U40200 (N_40200,N_38898,N_39476);
xor U40201 (N_40201,N_37529,N_38248);
or U40202 (N_40202,N_39783,N_38345);
xnor U40203 (N_40203,N_38833,N_39876);
nand U40204 (N_40204,N_39620,N_39126);
or U40205 (N_40205,N_37964,N_38050);
xor U40206 (N_40206,N_39230,N_39407);
nand U40207 (N_40207,N_38476,N_37583);
and U40208 (N_40208,N_39994,N_39867);
nand U40209 (N_40209,N_39102,N_37804);
nor U40210 (N_40210,N_38870,N_37731);
nand U40211 (N_40211,N_38701,N_39386);
nor U40212 (N_40212,N_39196,N_39602);
and U40213 (N_40213,N_38206,N_39179);
nand U40214 (N_40214,N_38671,N_38105);
and U40215 (N_40215,N_39214,N_38531);
or U40216 (N_40216,N_38734,N_38098);
or U40217 (N_40217,N_38156,N_39991);
and U40218 (N_40218,N_37698,N_39648);
or U40219 (N_40219,N_39111,N_38092);
nor U40220 (N_40220,N_37780,N_38286);
nor U40221 (N_40221,N_39485,N_38276);
nand U40222 (N_40222,N_38176,N_38904);
nand U40223 (N_40223,N_38553,N_39707);
nor U40224 (N_40224,N_38585,N_38759);
nor U40225 (N_40225,N_39719,N_39832);
or U40226 (N_40226,N_38187,N_37869);
xnor U40227 (N_40227,N_38311,N_38589);
or U40228 (N_40228,N_39844,N_39663);
or U40229 (N_40229,N_39885,N_39108);
nor U40230 (N_40230,N_38279,N_39182);
and U40231 (N_40231,N_38643,N_39741);
xnor U40232 (N_40232,N_38414,N_38537);
xnor U40233 (N_40233,N_38473,N_39727);
and U40234 (N_40234,N_37878,N_39623);
xnor U40235 (N_40235,N_39389,N_38096);
nand U40236 (N_40236,N_38935,N_37667);
nand U40237 (N_40237,N_39764,N_38043);
nor U40238 (N_40238,N_37939,N_38078);
nand U40239 (N_40239,N_39270,N_38861);
nand U40240 (N_40240,N_39863,N_39776);
and U40241 (N_40241,N_38660,N_38517);
or U40242 (N_40242,N_37776,N_39849);
or U40243 (N_40243,N_38128,N_37511);
and U40244 (N_40244,N_38013,N_38955);
nor U40245 (N_40245,N_37952,N_39070);
or U40246 (N_40246,N_37662,N_39592);
nand U40247 (N_40247,N_39668,N_37586);
and U40248 (N_40248,N_38238,N_38951);
and U40249 (N_40249,N_38915,N_39312);
and U40250 (N_40250,N_39933,N_38293);
xnor U40251 (N_40251,N_37663,N_37892);
nand U40252 (N_40252,N_38200,N_38233);
and U40253 (N_40253,N_38743,N_37658);
nand U40254 (N_40254,N_39558,N_39814);
or U40255 (N_40255,N_38758,N_37911);
nand U40256 (N_40256,N_38110,N_37675);
nand U40257 (N_40257,N_37753,N_38017);
and U40258 (N_40258,N_39952,N_39282);
xor U40259 (N_40259,N_38426,N_38781);
nor U40260 (N_40260,N_39496,N_39538);
nor U40261 (N_40261,N_38245,N_39427);
xor U40262 (N_40262,N_37818,N_38132);
nand U40263 (N_40263,N_39118,N_37500);
nor U40264 (N_40264,N_37512,N_39762);
or U40265 (N_40265,N_37708,N_39956);
nand U40266 (N_40266,N_37697,N_39871);
xnor U40267 (N_40267,N_38377,N_38384);
and U40268 (N_40268,N_39858,N_38111);
nand U40269 (N_40269,N_39552,N_38683);
nand U40270 (N_40270,N_38645,N_39774);
nor U40271 (N_40271,N_39382,N_39548);
xnor U40272 (N_40272,N_39923,N_39239);
and U40273 (N_40273,N_38259,N_39684);
nand U40274 (N_40274,N_39395,N_39815);
and U40275 (N_40275,N_38603,N_37870);
and U40276 (N_40276,N_38393,N_38045);
xnor U40277 (N_40277,N_37948,N_37584);
nand U40278 (N_40278,N_39096,N_38356);
nor U40279 (N_40279,N_39856,N_39784);
nor U40280 (N_40280,N_38803,N_39978);
or U40281 (N_40281,N_38561,N_38478);
nor U40282 (N_40282,N_37646,N_38130);
nor U40283 (N_40283,N_38515,N_39495);
or U40284 (N_40284,N_37971,N_37580);
and U40285 (N_40285,N_37569,N_39647);
or U40286 (N_40286,N_38109,N_38001);
and U40287 (N_40287,N_39971,N_39869);
nand U40288 (N_40288,N_38563,N_37837);
xnor U40289 (N_40289,N_39474,N_39011);
or U40290 (N_40290,N_38099,N_38764);
nand U40291 (N_40291,N_37608,N_39156);
nand U40292 (N_40292,N_39823,N_38810);
and U40293 (N_40293,N_39127,N_38359);
nand U40294 (N_40294,N_38090,N_38985);
xnor U40295 (N_40295,N_37655,N_38402);
nand U40296 (N_40296,N_38809,N_38753);
nor U40297 (N_40297,N_37756,N_37862);
and U40298 (N_40298,N_37953,N_39272);
xor U40299 (N_40299,N_39283,N_38146);
xor U40300 (N_40300,N_37897,N_38256);
nor U40301 (N_40301,N_37880,N_37526);
and U40302 (N_40302,N_37947,N_38009);
xnor U40303 (N_40303,N_38298,N_39804);
nor U40304 (N_40304,N_38060,N_38246);
nor U40305 (N_40305,N_37609,N_38661);
xor U40306 (N_40306,N_39437,N_37803);
or U40307 (N_40307,N_38868,N_39828);
nand U40308 (N_40308,N_38179,N_39542);
nand U40309 (N_40309,N_38063,N_37918);
nor U40310 (N_40310,N_39953,N_39367);
or U40311 (N_40311,N_39950,N_38501);
nor U40312 (N_40312,N_37882,N_37806);
or U40313 (N_40313,N_39562,N_38333);
and U40314 (N_40314,N_39738,N_37596);
or U40315 (N_40315,N_39269,N_38351);
nand U40316 (N_40316,N_39761,N_39431);
nand U40317 (N_40317,N_39170,N_37555);
or U40318 (N_40318,N_39642,N_38071);
xnor U40319 (N_40319,N_39477,N_37591);
xor U40320 (N_40320,N_37560,N_39020);
or U40321 (N_40321,N_39390,N_37700);
nand U40322 (N_40322,N_39820,N_39879);
nand U40323 (N_40323,N_39313,N_39092);
or U40324 (N_40324,N_38826,N_39157);
xnor U40325 (N_40325,N_39696,N_38455);
nor U40326 (N_40326,N_39775,N_39622);
xnor U40327 (N_40327,N_39247,N_37699);
and U40328 (N_40328,N_38565,N_37996);
or U40329 (N_40329,N_39633,N_39600);
and U40330 (N_40330,N_37634,N_39649);
nand U40331 (N_40331,N_38235,N_39186);
or U40332 (N_40332,N_39443,N_39503);
nand U40333 (N_40333,N_38946,N_38767);
xnor U40334 (N_40334,N_39128,N_37548);
nor U40335 (N_40335,N_37775,N_39075);
or U40336 (N_40336,N_39791,N_38220);
or U40337 (N_40337,N_39922,N_37866);
nand U40338 (N_40338,N_38514,N_37688);
nand U40339 (N_40339,N_39148,N_38178);
nand U40340 (N_40340,N_39843,N_39593);
or U40341 (N_40341,N_39031,N_39992);
xor U40342 (N_40342,N_38482,N_38771);
xnor U40343 (N_40343,N_37805,N_38309);
nor U40344 (N_40344,N_38385,N_38961);
xor U40345 (N_40345,N_39613,N_38824);
or U40346 (N_40346,N_38229,N_38979);
nand U40347 (N_40347,N_38970,N_38288);
nor U40348 (N_40348,N_38251,N_37851);
and U40349 (N_40349,N_37706,N_39409);
nor U40350 (N_40350,N_38785,N_37943);
and U40351 (N_40351,N_39038,N_37976);
nand U40352 (N_40352,N_38219,N_38557);
or U40353 (N_40353,N_38570,N_39638);
or U40354 (N_40354,N_39184,N_38494);
xor U40355 (N_40355,N_39291,N_39607);
and U40356 (N_40356,N_37727,N_38795);
nor U40357 (N_40357,N_37722,N_39693);
and U40358 (N_40358,N_38192,N_38143);
nor U40359 (N_40359,N_38047,N_37728);
and U40360 (N_40360,N_38472,N_39569);
nand U40361 (N_40361,N_37867,N_38843);
nand U40362 (N_40362,N_39827,N_38149);
and U40363 (N_40363,N_39449,N_38140);
xor U40364 (N_40364,N_39773,N_38606);
and U40365 (N_40365,N_38048,N_39072);
or U40366 (N_40366,N_38993,N_39275);
and U40367 (N_40367,N_38243,N_39415);
xor U40368 (N_40368,N_38665,N_37816);
or U40369 (N_40369,N_38736,N_39159);
xor U40370 (N_40370,N_38593,N_38142);
and U40371 (N_40371,N_38499,N_37724);
nand U40372 (N_40372,N_37611,N_38439);
xnor U40373 (N_40373,N_38878,N_37677);
nor U40374 (N_40374,N_39546,N_38370);
or U40375 (N_40375,N_38728,N_38163);
and U40376 (N_40376,N_38635,N_38058);
xnor U40377 (N_40377,N_39657,N_38422);
and U40378 (N_40378,N_38848,N_39778);
or U40379 (N_40379,N_38475,N_38911);
nand U40380 (N_40380,N_38940,N_37640);
nor U40381 (N_40381,N_39177,N_38835);
nor U40382 (N_40382,N_38117,N_38888);
xor U40383 (N_40383,N_39805,N_38107);
nor U40384 (N_40384,N_39475,N_39870);
xor U40385 (N_40385,N_39281,N_39811);
nand U40386 (N_40386,N_38084,N_38062);
nor U40387 (N_40387,N_39240,N_38564);
nand U40388 (N_40388,N_38582,N_38905);
and U40389 (N_40389,N_37597,N_39680);
nor U40390 (N_40390,N_38231,N_38825);
xnor U40391 (N_40391,N_37545,N_39133);
or U40392 (N_40392,N_38658,N_39375);
and U40393 (N_40393,N_37792,N_38274);
nor U40394 (N_40394,N_38427,N_38958);
and U40395 (N_40395,N_38614,N_39037);
nand U40396 (N_40396,N_39074,N_39686);
nor U40397 (N_40397,N_39217,N_39721);
xnor U40398 (N_40398,N_39771,N_38622);
and U40399 (N_40399,N_38464,N_37556);
nand U40400 (N_40400,N_38433,N_38108);
and U40401 (N_40401,N_37785,N_39153);
nand U40402 (N_40402,N_38398,N_39107);
and U40403 (N_40403,N_39681,N_39980);
xnor U40404 (N_40404,N_38005,N_39631);
nor U40405 (N_40405,N_38459,N_39779);
and U40406 (N_40406,N_39939,N_39362);
xnor U40407 (N_40407,N_37521,N_37979);
and U40408 (N_40408,N_39878,N_39183);
xor U40409 (N_40409,N_38232,N_38208);
and U40410 (N_40410,N_39530,N_39019);
nand U40411 (N_40411,N_39326,N_39484);
nand U40412 (N_40412,N_37995,N_38652);
and U40413 (N_40413,N_38014,N_38329);
or U40414 (N_40414,N_38992,N_38944);
nand U40415 (N_40415,N_39461,N_39615);
nand U40416 (N_40416,N_39087,N_39162);
or U40417 (N_40417,N_38730,N_39938);
and U40418 (N_40418,N_37509,N_38559);
nor U40419 (N_40419,N_37729,N_37773);
nor U40420 (N_40420,N_39131,N_37513);
nand U40421 (N_40421,N_38543,N_39524);
nor U40422 (N_40422,N_38039,N_39412);
nor U40423 (N_40423,N_37752,N_39290);
or U40424 (N_40424,N_39206,N_37749);
or U40425 (N_40425,N_38738,N_38722);
xor U40426 (N_40426,N_37973,N_39486);
nor U40427 (N_40427,N_37554,N_39756);
nand U40428 (N_40428,N_38886,N_37935);
or U40429 (N_40429,N_39429,N_37871);
or U40430 (N_40430,N_39116,N_38924);
or U40431 (N_40431,N_38204,N_37980);
xnor U40432 (N_40432,N_37668,N_38252);
nand U40433 (N_40433,N_39381,N_39208);
xnor U40434 (N_40434,N_38737,N_37991);
and U40435 (N_40435,N_39202,N_38907);
nand U40436 (N_40436,N_39260,N_37557);
nor U40437 (N_40437,N_37635,N_38400);
xor U40438 (N_40438,N_39222,N_39321);
nand U40439 (N_40439,N_38195,N_38594);
nand U40440 (N_40440,N_38502,N_39594);
and U40441 (N_40441,N_38925,N_38394);
or U40442 (N_40442,N_38929,N_38429);
or U40443 (N_40443,N_39608,N_37519);
xor U40444 (N_40444,N_38157,N_38676);
and U40445 (N_40445,N_38420,N_39903);
xnor U40446 (N_40446,N_37906,N_38746);
xnor U40447 (N_40447,N_38708,N_38885);
or U40448 (N_40448,N_37666,N_39284);
or U40449 (N_40449,N_38391,N_38386);
nor U40450 (N_40450,N_37789,N_37546);
xnor U40451 (N_40451,N_39563,N_39165);
xor U40452 (N_40452,N_39100,N_38700);
and U40453 (N_40453,N_38842,N_39556);
nand U40454 (N_40454,N_38479,N_39966);
or U40455 (N_40455,N_39785,N_39598);
or U40456 (N_40456,N_37531,N_37643);
and U40457 (N_40457,N_39830,N_39161);
and U40458 (N_40458,N_37576,N_39798);
nor U40459 (N_40459,N_39353,N_38503);
nand U40460 (N_40460,N_37732,N_39295);
and U40461 (N_40461,N_38381,N_38327);
or U40462 (N_40462,N_39340,N_39009);
xnor U40463 (N_40463,N_38840,N_39574);
nor U40464 (N_40464,N_38366,N_38093);
nand U40465 (N_40465,N_37779,N_38438);
nand U40466 (N_40466,N_38171,N_38272);
and U40467 (N_40467,N_38533,N_39905);
or U40468 (N_40468,N_39501,N_39001);
xor U40469 (N_40469,N_37684,N_39333);
and U40470 (N_40470,N_38726,N_37807);
or U40471 (N_40471,N_38547,N_38638);
and U40472 (N_40472,N_37567,N_39866);
and U40473 (N_40473,N_39176,N_37510);
and U40474 (N_40474,N_38278,N_39453);
or U40475 (N_40475,N_39249,N_38762);
nor U40476 (N_40476,N_38523,N_38451);
nand U40477 (N_40477,N_37903,N_39320);
xor U40478 (N_40478,N_39373,N_38265);
xnor U40479 (N_40479,N_39618,N_38281);
nor U40480 (N_40480,N_39931,N_39169);
or U40481 (N_40481,N_38480,N_38851);
and U40482 (N_40482,N_38409,N_39914);
nand U40483 (N_40483,N_39578,N_38421);
nor U40484 (N_40484,N_39628,N_39893);
nand U40485 (N_40485,N_38602,N_37965);
xor U40486 (N_40486,N_38936,N_38713);
xor U40487 (N_40487,N_38316,N_37915);
nand U40488 (N_40488,N_39305,N_39493);
nand U40489 (N_40489,N_39197,N_37725);
nor U40490 (N_40490,N_37620,N_39264);
or U40491 (N_40491,N_38672,N_38263);
or U40492 (N_40492,N_38147,N_37578);
or U40493 (N_40493,N_39998,N_39144);
and U40494 (N_40494,N_38632,N_38330);
and U40495 (N_40495,N_38677,N_37879);
xor U40496 (N_40496,N_39311,N_38573);
xor U40497 (N_40497,N_39644,N_39895);
nor U40498 (N_40498,N_37639,N_38657);
xnor U40499 (N_40499,N_38850,N_38069);
nor U40500 (N_40500,N_38228,N_38680);
or U40501 (N_40501,N_39226,N_39511);
nor U40502 (N_40502,N_38871,N_38579);
nand U40503 (N_40503,N_37957,N_38578);
or U40504 (N_40504,N_39257,N_39227);
nor U40505 (N_40505,N_38497,N_39268);
or U40506 (N_40506,N_38396,N_38218);
and U40507 (N_40507,N_38106,N_39845);
nand U40508 (N_40508,N_39755,N_37506);
and U40509 (N_40509,N_39724,N_38798);
and U40510 (N_40510,N_39745,N_37857);
nand U40511 (N_40511,N_38322,N_39276);
nand U40512 (N_40512,N_37632,N_38416);
and U40513 (N_40513,N_37650,N_38933);
xnor U40514 (N_40514,N_38640,N_38779);
nand U40515 (N_40515,N_37913,N_39654);
nor U40516 (N_40516,N_38122,N_39335);
xor U40517 (N_40517,N_37874,N_39007);
nor U40518 (N_40518,N_39471,N_38339);
nor U40519 (N_40519,N_39094,N_39327);
and U40520 (N_40520,N_38368,N_37648);
and U40521 (N_40521,N_39747,N_37654);
and U40522 (N_40522,N_38269,N_38682);
nand U40523 (N_40523,N_38725,N_38304);
and U40524 (N_40524,N_39763,N_38306);
xnor U40525 (N_40525,N_38823,N_39173);
nand U40526 (N_40526,N_39962,N_39140);
and U40527 (N_40527,N_39076,N_39894);
or U40528 (N_40528,N_38608,N_38996);
or U40529 (N_40529,N_38406,N_37746);
and U40530 (N_40530,N_39454,N_39666);
or U40531 (N_40531,N_38469,N_38748);
xnor U40532 (N_40532,N_37678,N_39656);
and U40533 (N_40533,N_39251,N_37625);
xnor U40534 (N_40534,N_38755,N_39446);
nand U40535 (N_40535,N_38967,N_39949);
nand U40536 (N_40536,N_39699,N_37622);
and U40537 (N_40537,N_37615,N_37593);
nor U40538 (N_40538,N_39073,N_39920);
nand U40539 (N_40539,N_38877,N_39687);
nor U40540 (N_40540,N_37589,N_39396);
or U40541 (N_40541,N_38332,N_39411);
xnor U40542 (N_40542,N_38485,N_38172);
nor U40543 (N_40543,N_37936,N_39015);
nor U40544 (N_40544,N_38695,N_39155);
nor U40545 (N_40545,N_39672,N_38018);
nand U40546 (N_40546,N_38978,N_38751);
nor U40547 (N_40547,N_38942,N_38847);
xnor U40548 (N_40548,N_37844,N_39854);
nand U40549 (N_40549,N_38816,N_38509);
or U40550 (N_40550,N_38261,N_37623);
or U40551 (N_40551,N_38075,N_38328);
and U40552 (N_40552,N_38223,N_38410);
xnor U40553 (N_40553,N_39308,N_37812);
and U40554 (N_40554,N_39941,N_39125);
or U40555 (N_40555,N_37676,N_38452);
nand U40556 (N_40556,N_39089,N_37754);
xnor U40557 (N_40557,N_38634,N_39749);
nand U40558 (N_40558,N_39789,N_38745);
or U40559 (N_40559,N_38169,N_39355);
and U40560 (N_40560,N_38668,N_38954);
nand U40561 (N_40561,N_39442,N_38367);
xnor U40562 (N_40562,N_38551,N_38361);
nor U40563 (N_40563,N_38095,N_38957);
xor U40564 (N_40564,N_39233,N_38181);
xnor U40565 (N_40565,N_38766,N_39555);
nor U40566 (N_40566,N_37905,N_38953);
and U40567 (N_40567,N_38308,N_39635);
or U40568 (N_40568,N_38937,N_39835);
or U40569 (N_40569,N_38808,N_38760);
or U40570 (N_40570,N_38390,N_37949);
and U40571 (N_40571,N_38828,N_39332);
and U40572 (N_40572,N_39120,N_38477);
xor U40573 (N_40573,N_38296,N_38917);
or U40574 (N_40574,N_37924,N_38138);
nand U40575 (N_40575,N_37956,N_38819);
xor U40576 (N_40576,N_38127,N_37709);
xnor U40577 (N_40577,N_39138,N_38262);
or U40578 (N_40578,N_38897,N_39918);
or U40579 (N_40579,N_38528,N_38526);
or U40580 (N_40580,N_38160,N_39579);
and U40581 (N_40581,N_39883,N_37978);
and U40582 (N_40582,N_38633,N_38932);
nor U40583 (N_40583,N_39466,N_39572);
nand U40584 (N_40584,N_39972,N_38267);
and U40585 (N_40585,N_38405,N_37734);
nor U40586 (N_40586,N_38310,N_38052);
or U40587 (N_40587,N_39862,N_37966);
nand U40588 (N_40588,N_39421,N_39204);
nor U40589 (N_40589,N_38401,N_38704);
nand U40590 (N_40590,N_39575,N_38428);
or U40591 (N_40591,N_37577,N_39838);
nand U40592 (N_40592,N_39737,N_37751);
and U40593 (N_40593,N_39033,N_38986);
or U40594 (N_40594,N_38891,N_39507);
xor U40595 (N_40595,N_38770,N_39322);
and U40596 (N_40596,N_39388,N_38520);
or U40597 (N_40597,N_39316,N_39730);
xnor U40598 (N_40598,N_37604,N_38280);
xor U40599 (N_40599,N_38037,N_38318);
nor U40600 (N_40600,N_39796,N_39262);
nor U40601 (N_40601,N_37989,N_38830);
nand U40602 (N_40602,N_38209,N_38723);
nand U40603 (N_40603,N_38651,N_38323);
or U40604 (N_40604,N_39800,N_39831);
nand U40605 (N_40605,N_39426,N_38292);
or U40606 (N_40606,N_38436,N_39709);
and U40607 (N_40607,N_39132,N_39231);
xor U40608 (N_40608,N_38969,N_37590);
xor U40609 (N_40609,N_39225,N_38776);
or U40610 (N_40610,N_37561,N_39639);
nand U40611 (N_40611,N_39872,N_39497);
and U40612 (N_40612,N_38590,N_38711);
or U40613 (N_40613,N_39143,N_38631);
nor U40614 (N_40614,N_38010,N_37967);
nor U40615 (N_40615,N_38890,N_39018);
nor U40616 (N_40616,N_38158,N_37739);
xor U40617 (N_40617,N_39728,N_38534);
or U40618 (N_40618,N_39944,N_37755);
and U40619 (N_40619,N_37926,N_39850);
nor U40620 (N_40620,N_38615,N_38909);
and U40621 (N_40621,N_38930,N_38820);
nor U40622 (N_40622,N_37916,N_39363);
nor U40623 (N_40623,N_39039,N_39576);
xor U40624 (N_40624,N_38595,N_39430);
nand U40625 (N_40625,N_39625,N_39135);
or U40626 (N_40626,N_38445,N_39079);
and U40627 (N_40627,N_39513,N_38965);
xnor U40628 (N_40628,N_38413,N_38159);
or U40629 (N_40629,N_38383,N_38862);
nand U40630 (N_40630,N_38976,N_37602);
and U40631 (N_40631,N_39840,N_39960);
or U40632 (N_40632,N_38411,N_39637);
xor U40633 (N_40633,N_38874,N_39525);
xnor U40634 (N_40634,N_38474,N_38991);
nand U40635 (N_40635,N_38696,N_38535);
xor U40636 (N_40636,N_38380,N_39053);
and U40637 (N_40637,N_38750,N_39480);
nand U40638 (N_40638,N_38837,N_37631);
nor U40639 (N_40639,N_39250,N_39044);
and U40640 (N_40640,N_38546,N_39665);
xor U40641 (N_40641,N_37603,N_38382);
and U40642 (N_40642,N_37507,N_39403);
xor U40643 (N_40643,N_37877,N_38183);
and U40644 (N_40644,N_37988,N_38705);
nand U40645 (N_40645,N_39121,N_39677);
nand U40646 (N_40646,N_38112,N_38814);
xnor U40647 (N_40647,N_37657,N_39351);
nor U40648 (N_40648,N_39753,N_38642);
nand U40649 (N_40649,N_39301,N_38408);
or U40650 (N_40650,N_38289,N_38363);
nor U40651 (N_40651,N_37637,N_38100);
or U40652 (N_40652,N_39566,N_38539);
xor U40653 (N_40653,N_37523,N_39330);
xor U40654 (N_40654,N_39585,N_39627);
nand U40655 (N_40655,N_39425,N_37535);
xnor U40656 (N_40656,N_37768,N_38613);
nor U40657 (N_40657,N_38041,N_37941);
xor U40658 (N_40658,N_39234,N_38807);
nor U40659 (N_40659,N_39505,N_38015);
and U40660 (N_40660,N_37652,N_39702);
xnor U40661 (N_40661,N_37863,N_39216);
nand U40662 (N_40662,N_39376,N_37798);
xnor U40663 (N_40663,N_39926,N_39924);
or U40664 (N_40664,N_38550,N_39185);
nor U40665 (N_40665,N_37854,N_37600);
nor U40666 (N_40666,N_38126,N_37846);
xor U40667 (N_40667,N_38425,N_37750);
nand U40668 (N_40668,N_37575,N_38441);
xor U40669 (N_40669,N_39661,N_37845);
xnor U40670 (N_40670,N_38845,N_39772);
and U40671 (N_40671,N_39168,N_39695);
xnor U40672 (N_40672,N_37685,N_39690);
nand U40673 (N_40673,N_38285,N_38831);
nor U40674 (N_40674,N_37553,N_38055);
or U40675 (N_40675,N_39160,N_37840);
nand U40676 (N_40676,N_37672,N_37743);
or U40677 (N_40677,N_39588,N_39067);
and U40678 (N_40678,N_39857,N_39491);
nand U40679 (N_40679,N_38212,N_39023);
nand U40680 (N_40680,N_39909,N_38202);
nand U40681 (N_40681,N_38344,N_39646);
nor U40682 (N_40682,N_39224,N_37723);
or U40683 (N_40683,N_39137,N_37962);
xor U40684 (N_40684,N_38136,N_38945);
or U40685 (N_40685,N_39099,N_38568);
and U40686 (N_40686,N_38687,N_39366);
and U40687 (N_40687,N_37858,N_37895);
and U40688 (N_40688,N_38068,N_38576);
nand U40689 (N_40689,N_37679,N_38599);
and U40690 (N_40690,N_38938,N_38572);
and U40691 (N_40691,N_39360,N_38801);
nor U40692 (N_40692,N_39106,N_37737);
and U40693 (N_40693,N_38995,N_38415);
or U40694 (N_40694,N_38956,N_37644);
and U40695 (N_40695,N_38800,N_38974);
or U40696 (N_40696,N_39046,N_39119);
nor U40697 (N_40697,N_39582,N_39002);
and U40698 (N_40698,N_38299,N_39200);
and U40699 (N_40699,N_39948,N_39078);
and U40700 (N_40700,N_37501,N_39921);
nand U40701 (N_40701,N_38921,N_38153);
nand U40702 (N_40702,N_39090,N_37680);
and U40703 (N_40703,N_39865,N_38114);
or U40704 (N_40704,N_37910,N_38102);
and U40705 (N_40705,N_38806,N_38574);
nor U40706 (N_40706,N_37689,N_38855);
nand U40707 (N_40707,N_39146,N_38538);
nor U40708 (N_40708,N_39630,N_38215);
nand U40709 (N_40709,N_39152,N_37850);
xnor U40710 (N_40710,N_39817,N_38707);
or U40711 (N_40711,N_39940,N_37551);
nand U40712 (N_40712,N_37987,N_37790);
xnor U40713 (N_40713,N_37772,N_38536);
xor U40714 (N_40714,N_37503,N_38355);
xor U40715 (N_40715,N_39085,N_38518);
and U40716 (N_40716,N_37848,N_37547);
xor U40717 (N_40717,N_37664,N_38397);
nand U40718 (N_40718,N_39232,N_37524);
and U40719 (N_40719,N_37549,N_38918);
nor U40720 (N_40720,N_37891,N_38994);
and U40721 (N_40721,N_38919,N_37520);
or U40722 (N_40722,N_38307,N_38987);
or U40723 (N_40723,N_39713,N_38525);
xor U40724 (N_40724,N_37771,N_37808);
xnor U40725 (N_40725,N_39968,N_38254);
or U40726 (N_40726,N_39781,N_38569);
xnor U40727 (N_40727,N_39539,N_38241);
xor U40728 (N_40728,N_39786,N_38495);
nand U40729 (N_40729,N_39508,N_38273);
xnor U40730 (N_40730,N_39988,N_39358);
or U40731 (N_40731,N_39052,N_39334);
xor U40732 (N_40732,N_38818,N_39219);
nand U40733 (N_40733,N_38962,N_38605);
nand U40734 (N_40734,N_37968,N_37794);
or U40735 (N_40735,N_37864,N_39989);
nand U40736 (N_40736,N_38461,N_37598);
nand U40737 (N_40737,N_38655,N_38747);
nor U40738 (N_40738,N_37908,N_38369);
or U40739 (N_40739,N_39253,N_37999);
xnor U40740 (N_40740,N_39540,N_39029);
and U40741 (N_40741,N_38072,N_37970);
and U40742 (N_40742,N_39371,N_37893);
and U40743 (N_40743,N_37830,N_38490);
or U40744 (N_40744,N_39722,N_38094);
or U40745 (N_40745,N_37540,N_38856);
xnor U40746 (N_40746,N_39084,N_38681);
nand U40747 (N_40747,N_38902,N_39058);
nor U40748 (N_40748,N_39810,N_38812);
nor U40749 (N_40749,N_37559,N_37791);
and U40750 (N_40750,N_38335,N_39590);
nor U40751 (N_40751,N_39004,N_37641);
nor U40752 (N_40752,N_37638,N_38190);
nor U40753 (N_40753,N_39675,N_38662);
and U40754 (N_40754,N_39095,N_39187);
nand U40755 (N_40755,N_39103,N_37612);
and U40756 (N_40756,N_39286,N_38407);
nand U40757 (N_40757,N_37660,N_39519);
nand U40758 (N_40758,N_39054,N_38511);
and U40759 (N_40759,N_38577,N_38207);
or U40760 (N_40760,N_38131,N_39861);
nand U40761 (N_40761,N_39812,N_38596);
and U40762 (N_40762,N_37585,N_39907);
xnor U40763 (N_40763,N_39259,N_37726);
nor U40764 (N_40764,N_37624,N_39896);
nor U40765 (N_40765,N_39035,N_37885);
and U40766 (N_40766,N_39387,N_39267);
xor U40767 (N_40767,N_39498,N_39016);
nor U40768 (N_40768,N_39545,N_39017);
or U40769 (N_40769,N_39643,N_39793);
and U40770 (N_40770,N_39328,N_38880);
nor U40771 (N_40771,N_39634,N_39703);
nor U40772 (N_40772,N_38947,N_39378);
nor U40773 (N_40773,N_39990,N_37787);
nand U40774 (N_40774,N_38973,N_39408);
xnor U40775 (N_40775,N_39970,N_38028);
nor U40776 (N_40776,N_37594,N_37695);
and U40777 (N_40777,N_38685,N_39541);
nor U40778 (N_40778,N_37861,N_38777);
xnor U40779 (N_40779,N_38783,N_39422);
nand U40780 (N_40780,N_39459,N_38966);
or U40781 (N_40781,N_38981,N_39008);
or U40782 (N_40782,N_39640,N_39752);
nor U40783 (N_40783,N_39587,N_39662);
nand U40784 (N_40784,N_39465,N_38717);
xnor U40785 (N_40785,N_38081,N_39401);
nand U40786 (N_40786,N_39746,N_38226);
xor U40787 (N_40787,N_39981,N_39958);
and U40788 (N_40788,N_37839,N_38689);
and U40789 (N_40789,N_39516,N_37595);
nor U40790 (N_40790,N_39086,N_38189);
nand U40791 (N_40791,N_38586,N_37522);
or U40792 (N_40792,N_39706,N_39794);
xnor U40793 (N_40793,N_39205,N_38129);
and U40794 (N_40794,N_38694,N_37617);
nand U40795 (N_40795,N_38882,N_38697);
nor U40796 (N_40796,N_37745,N_39782);
nand U40797 (N_40797,N_39780,N_39645);
xor U40798 (N_40798,N_37946,N_38284);
and U40799 (N_40799,N_38148,N_38698);
and U40800 (N_40800,N_37537,N_39163);
nor U40801 (N_40801,N_39167,N_38379);
nand U40802 (N_40802,N_37505,N_38389);
and U40803 (N_40803,N_37610,N_39908);
xor U40804 (N_40804,N_39274,N_38827);
or U40805 (N_40805,N_39350,N_38342);
and U40806 (N_40806,N_39083,N_38086);
nor U40807 (N_40807,N_38858,N_39293);
and U40808 (N_40808,N_39428,N_38731);
nand U40809 (N_40809,N_39549,N_39354);
nand U40810 (N_40810,N_37985,N_37528);
and U40811 (N_40811,N_37572,N_38225);
or U40812 (N_40812,N_39115,N_37766);
nor U40813 (N_40813,N_38740,N_38404);
nand U40814 (N_40814,N_37920,N_39544);
xnor U40815 (N_40815,N_39609,N_38213);
nand U40816 (N_40816,N_39010,N_39192);
nand U40817 (N_40817,N_37859,N_37825);
or U40818 (N_40818,N_37856,N_37824);
and U40819 (N_40819,N_38649,N_37853);
nor U40820 (N_40820,N_37516,N_38372);
xor U40821 (N_40821,N_39705,N_38196);
nor U40822 (N_40822,N_38326,N_37811);
xnor U40823 (N_40823,N_38530,N_38647);
and U40824 (N_40824,N_38644,N_39248);
xnor U40825 (N_40825,N_38253,N_38161);
nor U40826 (N_40826,N_37651,N_39451);
and U40827 (N_40827,N_39955,N_38587);
nor U40828 (N_40828,N_39134,N_38675);
xnor U40829 (N_40829,N_37629,N_38674);
and U40830 (N_40830,N_38175,N_38629);
nand U40831 (N_40831,N_38216,N_37552);
nand U40832 (N_40832,N_37686,N_39235);
and U40833 (N_40833,N_39175,N_39488);
or U40834 (N_40834,N_39410,N_38365);
and U40835 (N_40835,N_37876,N_39957);
and U40836 (N_40836,N_38360,N_37977);
nand U40837 (N_40837,N_37799,N_39082);
xor U40838 (N_40838,N_37538,N_39688);
nand U40839 (N_40839,N_37774,N_38255);
nor U40840 (N_40840,N_39049,N_37954);
and U40841 (N_40841,N_38011,N_38173);
and U40842 (N_40842,N_37993,N_39345);
nor U40843 (N_40843,N_39258,N_39975);
or U40844 (N_40844,N_38155,N_38964);
nor U40845 (N_40845,N_37717,N_37696);
and U40846 (N_40846,N_38690,N_39877);
or U40847 (N_40847,N_39660,N_38860);
xnor U40848 (N_40848,N_38492,N_37982);
and U40849 (N_40849,N_39034,N_38763);
xor U40850 (N_40850,N_37541,N_39419);
xnor U40851 (N_40851,N_38338,N_39385);
xor U40852 (N_40852,N_38103,N_39400);
nand U40853 (N_40853,N_39030,N_39947);
and U40854 (N_40854,N_39710,N_39976);
or U40855 (N_40855,N_37544,N_38193);
or U40856 (N_40856,N_37619,N_38712);
and U40857 (N_40857,N_37661,N_37826);
and U40858 (N_40858,N_38972,N_37884);
nor U40859 (N_40859,N_38718,N_37565);
and U40860 (N_40860,N_39112,N_39565);
nand U40861 (N_40861,N_39610,N_37621);
xor U40862 (N_40862,N_39213,N_38959);
xnor U40863 (N_40863,N_37809,N_39701);
or U40864 (N_40864,N_37536,N_37889);
and U40865 (N_40865,N_39616,N_37562);
nand U40866 (N_40866,N_39056,N_39207);
xnor U40867 (N_40867,N_38295,N_39434);
nand U40868 (N_40868,N_39750,N_39819);
nor U40869 (N_40869,N_37800,N_38141);
nand U40870 (N_40870,N_38085,N_38419);
and U40871 (N_40871,N_38742,N_39993);
xor U40872 (N_40872,N_38054,N_39455);
nor U40873 (N_40873,N_37795,N_39736);
or U40874 (N_40874,N_38881,N_38950);
or U40875 (N_40875,N_38040,N_38899);
or U40876 (N_40876,N_39522,N_39839);
and U40877 (N_40877,N_37886,N_39529);
xor U40878 (N_40878,N_39297,N_38337);
xor U40879 (N_40879,N_39139,N_39347);
nor U40880 (N_40880,N_38625,N_37543);
xor U40881 (N_40881,N_38754,N_38505);
nand U40882 (N_40882,N_38512,N_38616);
and U40883 (N_40883,N_38151,N_38031);
or U40884 (N_40884,N_39014,N_39468);
or U40885 (N_40885,N_39928,N_37613);
nor U40886 (N_40886,N_39930,N_38317);
nor U40887 (N_40887,N_38305,N_39243);
and U40888 (N_40888,N_39999,N_39406);
or U40889 (N_40889,N_39263,N_39765);
or U40890 (N_40890,N_39685,N_37627);
nor U40891 (N_40891,N_39768,N_39101);
nor U40892 (N_40892,N_38873,N_37669);
or U40893 (N_40893,N_39915,N_37860);
nand U40894 (N_40894,N_39601,N_39280);
xor U40895 (N_40895,N_38797,N_39632);
nor U40896 (N_40896,N_39490,N_38691);
and U40897 (N_40897,N_39024,N_38282);
xnor U40898 (N_40898,N_38903,N_37694);
nand U40899 (N_40899,N_38732,N_37601);
xnor U40900 (N_40900,N_39129,N_39042);
nand U40901 (N_40901,N_38059,N_37934);
nand U40902 (N_40902,N_37923,N_39974);
and U40903 (N_40903,N_37571,N_37937);
and U40904 (N_40904,N_39287,N_38258);
nand U40905 (N_40905,N_38214,N_37960);
or U40906 (N_40906,N_39319,N_39833);
and U40907 (N_40907,N_39093,N_39088);
and U40908 (N_40908,N_38529,N_39417);
xor U40909 (N_40909,N_39323,N_37748);
or U40910 (N_40910,N_38867,N_37702);
nand U40911 (N_40911,N_39739,N_39081);
xnor U40912 (N_40912,N_39532,N_39325);
xnor U40913 (N_40913,N_38290,N_39664);
nand U40914 (N_40914,N_38817,N_37581);
xnor U40915 (N_40915,N_38053,N_39199);
or U40916 (N_40916,N_39369,N_39000);
xnor U40917 (N_40917,N_38314,N_38580);
nor U40918 (N_40918,N_39790,N_37683);
nand U40919 (N_40919,N_38778,N_38510);
nand U40920 (N_40920,N_38724,N_37665);
xor U40921 (N_40921,N_39420,N_39380);
nor U40922 (N_40922,N_39458,N_38834);
nor U40923 (N_40923,N_39314,N_37730);
nor U40924 (N_40924,N_38257,N_37940);
nor U40925 (N_40925,N_38354,N_38437);
nand U40926 (N_40926,N_38006,N_37705);
or U40927 (N_40927,N_39384,N_38026);
and U40928 (N_40928,N_37653,N_39441);
xor U40929 (N_40929,N_39147,N_39571);
nor U40930 (N_40930,N_39344,N_38522);
xnor U40931 (N_40931,N_39603,N_38065);
nand U40932 (N_40932,N_39489,N_38788);
or U40933 (N_40933,N_39198,N_39483);
xnor U40934 (N_40934,N_37921,N_39621);
and U40935 (N_40935,N_39278,N_39467);
nor U40936 (N_40936,N_39296,N_37539);
xnor U40937 (N_40937,N_39822,N_38939);
nor U40938 (N_40938,N_39580,N_38624);
xnor U40939 (N_40939,N_39482,N_39352);
and U40940 (N_40940,N_39080,N_39674);
nor U40941 (N_40941,N_39065,N_37757);
or U40942 (N_40942,N_38287,N_39246);
or U40943 (N_40943,N_37942,N_39570);
xnor U40944 (N_40944,N_37990,N_39494);
and U40945 (N_40945,N_39596,N_39057);
or U40946 (N_40946,N_39581,N_39370);
nor U40947 (N_40947,N_39265,N_38387);
nand U40948 (N_40948,N_39726,N_39338);
nor U40949 (N_40949,N_38056,N_37781);
and U40950 (N_40950,N_39171,N_39676);
nand U40951 (N_40951,N_39036,N_38600);
xnor U40952 (N_40952,N_38012,N_37550);
or U40953 (N_40953,N_39114,N_38234);
nand U40954 (N_40954,N_38920,N_38080);
xor U40955 (N_40955,N_39985,N_39022);
nand U40956 (N_40956,N_37983,N_37944);
nand U40957 (N_40957,N_37958,N_39005);
or U40958 (N_40958,N_38275,N_37875);
nor U40959 (N_40959,N_39189,N_37763);
xnor U40960 (N_40960,N_38620,N_39329);
and U40961 (N_40961,N_39669,N_37894);
and U40962 (N_40962,N_39967,N_37784);
and U40963 (N_40963,N_38205,N_39255);
xor U40964 (N_40964,N_37793,N_38484);
nor U40965 (N_40965,N_39456,N_37690);
nor U40966 (N_40966,N_39729,N_38024);
xnor U40967 (N_40967,N_38786,N_37525);
and U40968 (N_40968,N_39821,N_39405);
and U40969 (N_40969,N_38066,N_39853);
nor U40970 (N_40970,N_39758,N_39423);
nor U40971 (N_40971,N_38558,N_37963);
xor U40972 (N_40972,N_37761,N_38498);
nor U40973 (N_40973,N_39731,N_38217);
nand U40974 (N_40974,N_39357,N_38357);
or U40975 (N_40975,N_39097,N_37981);
nand U40976 (N_40976,N_38120,N_38650);
or U40977 (N_40977,N_38000,N_38491);
nor U40978 (N_40978,N_39912,N_39777);
and U40979 (N_40979,N_39504,N_38118);
xnor U40980 (N_40980,N_39937,N_39534);
or U40981 (N_40981,N_38022,N_39502);
nor U40982 (N_40982,N_37574,N_37712);
or U40983 (N_40983,N_38607,N_38829);
xor U40984 (N_40984,N_38678,N_38782);
and U40985 (N_40985,N_39984,N_37842);
nor U40986 (N_40986,N_39936,N_37558);
or U40987 (N_40987,N_39266,N_38506);
xor U40988 (N_40988,N_38853,N_37530);
and U40989 (N_40989,N_37721,N_39444);
xor U40990 (N_40990,N_39934,N_39397);
nand U40991 (N_40991,N_38450,N_38960);
nand U40992 (N_40992,N_38883,N_38581);
xor U40993 (N_40993,N_38716,N_39241);
nor U40994 (N_40994,N_38489,N_38399);
nand U40995 (N_40995,N_39462,N_39026);
or U40996 (N_40996,N_38802,N_38846);
nand U40997 (N_40997,N_38637,N_39929);
nand U40998 (N_40998,N_39788,N_39533);
xor U40999 (N_40999,N_39834,N_39003);
nand U41000 (N_41000,N_39048,N_38869);
and U41001 (N_41001,N_39959,N_38588);
nand U41002 (N_41002,N_37928,N_37747);
and U41003 (N_41003,N_39432,N_39717);
and U41004 (N_41004,N_38079,N_38621);
nor U41005 (N_41005,N_37896,N_38639);
nor U41006 (N_41006,N_38300,N_37616);
and U41007 (N_41007,N_39142,N_38448);
nand U41008 (N_41008,N_39174,N_38004);
and U41009 (N_41009,N_38417,N_37764);
nor U41010 (N_41010,N_39900,N_38686);
nor U41011 (N_41011,N_37887,N_39279);
xor U41012 (N_41012,N_38804,N_38418);
xor U41013 (N_41013,N_39678,N_39306);
and U41014 (N_41014,N_39510,N_37959);
or U41015 (N_41015,N_38659,N_38194);
xor U41016 (N_41016,N_38266,N_39218);
and U41017 (N_41017,N_38145,N_37888);
and U41018 (N_41018,N_38467,N_38375);
and U41019 (N_41019,N_38447,N_39943);
xnor U41020 (N_41020,N_39961,N_38430);
or U41021 (N_41021,N_38186,N_38999);
nor U41022 (N_41022,N_39557,N_38180);
nor U41023 (N_41023,N_38884,N_39368);
xor U41024 (N_41024,N_37873,N_38487);
nor U41025 (N_41025,N_38928,N_39331);
or U41026 (N_41026,N_39825,N_39318);
nand U41027 (N_41027,N_39063,N_39787);
xnor U41028 (N_41028,N_38264,N_38733);
xor U41029 (N_41029,N_39487,N_38496);
or U41030 (N_41030,N_39299,N_37831);
xor U41031 (N_41031,N_38164,N_38500);
xnor U41032 (N_41032,N_38912,N_39300);
and U41033 (N_41033,N_38739,N_39559);
nand U41034 (N_41034,N_38811,N_37849);
nand U41035 (N_41035,N_39341,N_37770);
nand U41036 (N_41036,N_38892,N_38879);
nor U41037 (N_41037,N_37817,N_39718);
and U41038 (N_41038,N_37909,N_39584);
nand U41039 (N_41039,N_39527,N_39194);
xor U41040 (N_41040,N_38007,N_39523);
or U41041 (N_41041,N_38227,N_39141);
nand U41042 (N_41042,N_37930,N_37890);
xor U41043 (N_41043,N_38916,N_39842);
or U41044 (N_41044,N_39611,N_39124);
nand U41045 (N_41045,N_38135,N_38203);
or U41046 (N_41046,N_38527,N_38376);
nor U41047 (N_41047,N_39051,N_39436);
nand U41048 (N_41048,N_37819,N_37692);
xor U41049 (N_41049,N_37703,N_39181);
nor U41050 (N_41050,N_39583,N_37881);
nor U41051 (N_41051,N_39641,N_38549);
nand U41052 (N_41052,N_37783,N_39201);
nor U41053 (N_41053,N_37533,N_38859);
nor U41054 (N_41054,N_38444,N_37738);
or U41055 (N_41055,N_38623,N_39612);
or U41056 (N_41056,N_39543,N_37626);
nor U41057 (N_41057,N_39041,N_37827);
and U41058 (N_41058,N_39759,N_39973);
or U41059 (N_41059,N_39671,N_38277);
nand U41060 (N_41060,N_38949,N_39136);
xnor U41061 (N_41061,N_37898,N_38003);
nor U41062 (N_41062,N_38654,N_39399);
or U41063 (N_41063,N_37929,N_37502);
nand U41064 (N_41064,N_38046,N_39554);
or U41065 (N_41065,N_38575,N_38325);
nand U41066 (N_41066,N_37984,N_37823);
xnor U41067 (N_41067,N_37796,N_39068);
nand U41068 (N_41068,N_37835,N_38646);
nand U41069 (N_41069,N_39514,N_39667);
and U41070 (N_41070,N_37938,N_39472);
and U41071 (N_41071,N_38790,N_38875);
xnor U41072 (N_41072,N_38210,N_38604);
or U41073 (N_41073,N_38706,N_38242);
xnor U41074 (N_41074,N_37647,N_38663);
xnor U41075 (N_41075,N_39105,N_39964);
nor U41076 (N_41076,N_39965,N_39560);
xnor U41077 (N_41077,N_39670,N_39098);
or U41078 (N_41078,N_38749,N_37517);
nor U41079 (N_41079,N_39704,N_39807);
xnor U41080 (N_41080,N_39997,N_38182);
xor U41081 (N_41081,N_37570,N_39288);
nand U41082 (N_41082,N_38813,N_39904);
or U41083 (N_41083,N_39145,N_39464);
and U41084 (N_41084,N_37707,N_39714);
xor U41085 (N_41085,N_38008,N_37716);
nor U41086 (N_41086,N_38341,N_38567);
nand U41087 (N_41087,N_38346,N_38088);
xnor U41088 (N_41088,N_38612,N_37588);
nor U41089 (N_41089,N_39597,N_38166);
nor U41090 (N_41090,N_39178,N_38144);
xor U41091 (N_41091,N_38982,N_39500);
and U41092 (N_41092,N_37951,N_39317);
xor U41093 (N_41093,N_39110,N_38864);
or U41094 (N_41094,N_39983,N_37568);
nor U41095 (N_41095,N_39526,N_37618);
nor U41096 (N_41096,N_39536,N_38294);
nand U41097 (N_41097,N_38775,N_38721);
nor U41098 (N_41098,N_39824,N_38592);
and U41099 (N_41099,N_38922,N_39452);
nand U41100 (N_41100,N_39734,N_37847);
xor U41101 (N_41101,N_39694,N_38667);
xor U41102 (N_41102,N_38331,N_39531);
nand U41103 (N_41103,N_39315,N_38373);
nand U41104 (N_41104,N_39803,N_39891);
nor U41105 (N_41105,N_37972,N_38895);
nand U41106 (N_41106,N_37758,N_38854);
or U41107 (N_41107,N_39868,N_37564);
or U41108 (N_41108,N_37912,N_38591);
nor U41109 (N_41109,N_38934,N_38097);
or U41110 (N_41110,N_38466,N_39261);
or U41111 (N_41111,N_39460,N_39916);
or U41112 (N_41112,N_38185,N_37832);
xnor U41113 (N_41113,N_38787,N_38618);
nor U41114 (N_41114,N_38125,N_37769);
and U41115 (N_41115,N_37628,N_39708);
xor U41116 (N_41116,N_37711,N_39228);
nand U41117 (N_41117,N_39062,N_39550);
nand U41118 (N_41118,N_39954,N_37833);
nor U41119 (N_41119,N_39256,N_39711);
xor U41120 (N_41120,N_37788,N_39682);
nor U41121 (N_41121,N_37872,N_38702);
xnor U41122 (N_41122,N_39424,N_38221);
xnor U41123 (N_41123,N_38684,N_39518);
nand U41124 (N_41124,N_38456,N_38822);
and U41125 (N_41125,N_39884,N_38876);
or U41126 (N_41126,N_38465,N_38666);
xnor U41127 (N_41127,N_37901,N_38815);
or U41128 (N_41128,N_39927,N_38303);
and U41129 (N_41129,N_39932,N_39573);
or U41130 (N_41130,N_39013,N_37852);
nand U41131 (N_41131,N_37834,N_38076);
nor U41132 (N_41132,N_39069,N_37883);
or U41133 (N_41133,N_39799,N_39614);
nand U41134 (N_41134,N_39245,N_38988);
and U41135 (N_41135,N_37599,N_39066);
and U41136 (N_41136,N_38619,N_38364);
or U41137 (N_41137,N_39535,N_39902);
nand U41138 (N_41138,N_38780,N_39852);
xor U41139 (N_41139,N_38735,N_37693);
and U41140 (N_41140,N_38378,N_38334);
or U41141 (N_41141,N_37907,N_38519);
nor U41142 (N_41142,N_38507,N_39586);
and U41143 (N_41143,N_38199,N_37974);
nand U41144 (N_41144,N_39223,N_38524);
xor U41145 (N_41145,N_39770,N_37914);
xor U41146 (N_41146,N_39040,N_39149);
nand U41147 (N_41147,N_38191,N_39888);
xnor U41148 (N_41148,N_38483,N_38030);
and U41149 (N_41149,N_38688,N_39655);
or U41150 (N_41150,N_37932,N_38083);
nand U41151 (N_41151,N_39847,N_37900);
or U41152 (N_41152,N_39874,N_37762);
and U41153 (N_41153,N_39841,N_38442);
nand U41154 (N_41154,N_38123,N_39433);
xnor U41155 (N_41155,N_39393,N_38963);
xnor U41156 (N_41156,N_38042,N_37838);
nand U41157 (N_41157,N_39479,N_39509);
and U41158 (N_41158,N_39732,N_39892);
nor U41159 (N_41159,N_38583,N_38358);
nor U41160 (N_41160,N_38761,N_38481);
xnor U41161 (N_41161,N_38989,N_37821);
xnor U41162 (N_41162,N_39901,N_38720);
nor U41163 (N_41163,N_38571,N_39935);
and U41164 (N_41164,N_39875,N_39123);
or U41165 (N_41165,N_39801,N_39880);
and U41166 (N_41166,N_38542,N_39324);
xnor U41167 (N_41167,N_38693,N_38841);
or U41168 (N_41168,N_39882,N_39292);
xor U41169 (N_41169,N_38134,N_38710);
nand U41170 (N_41170,N_39180,N_38521);
nor U41171 (N_41171,N_38324,N_38343);
and U41172 (N_41172,N_39629,N_39725);
nor U41173 (N_41173,N_39740,N_38789);
and U41174 (N_41174,N_38115,N_39797);
nand U41175 (N_41175,N_39043,N_38630);
nor U41176 (N_41176,N_39735,N_38119);
or U41177 (N_41177,N_38002,N_39212);
and U41178 (N_41178,N_39743,N_38460);
or U41179 (N_41179,N_38774,N_38077);
nor U41180 (N_41180,N_38463,N_39512);
and U41181 (N_41181,N_37563,N_38152);
xnor U41182 (N_41182,N_38250,N_39890);
or U41183 (N_41183,N_38887,N_38709);
or U41184 (N_41184,N_39285,N_38796);
nor U41185 (N_41185,N_37955,N_39242);
and U41186 (N_41186,N_38139,N_38061);
nor U41187 (N_41187,N_39987,N_37605);
and U41188 (N_41188,N_37719,N_37691);
or U41189 (N_41189,N_38230,N_39025);
or U41190 (N_41190,N_37742,N_38034);
and U41191 (N_41191,N_39377,N_38239);
nand U41192 (N_41192,N_38741,N_37922);
nand U41193 (N_41193,N_39071,N_37828);
nand U41194 (N_41194,N_38412,N_39899);
or U41195 (N_41195,N_38931,N_37713);
and U41196 (N_41196,N_39481,N_39303);
nand U41197 (N_41197,N_37777,N_39873);
xnor U41198 (N_41198,N_38744,N_39521);
nand U41199 (N_41199,N_37527,N_39816);
nand U41200 (N_41200,N_39917,N_38432);
and U41201 (N_41201,N_39158,N_38113);
xnor U41202 (N_41202,N_39254,N_39203);
or U41203 (N_41203,N_37630,N_39414);
nand U41204 (N_41204,N_38057,N_38673);
nand U41205 (N_41205,N_39091,N_37868);
nand U41206 (N_41206,N_39391,N_38493);
xnor U41207 (N_41207,N_38167,N_38137);
nand U41208 (N_41208,N_38315,N_38297);
nor U41209 (N_41209,N_39906,N_39595);
xnor U41210 (N_41210,N_38910,N_38302);
xor U41211 (N_41211,N_39652,N_38312);
or U41212 (N_41212,N_39032,N_39061);
and U41213 (N_41213,N_37704,N_37904);
nand U41214 (N_41214,N_39298,N_38794);
and U41215 (N_41215,N_39164,N_38765);
and U41216 (N_41216,N_37899,N_38124);
nor U41217 (N_41217,N_38440,N_38997);
or U41218 (N_41218,N_37518,N_38626);
nand U41219 (N_41219,N_38821,N_39963);
or U41220 (N_41220,N_39537,N_39047);
nand U41221 (N_41221,N_38983,N_37997);
or U41222 (N_41222,N_38362,N_38792);
xor U41223 (N_41223,N_38170,N_38756);
or U41224 (N_41224,N_38609,N_39712);
or U41225 (N_41225,N_39064,N_38291);
nor U41226 (N_41226,N_37961,N_39113);
and U41227 (N_41227,N_38374,N_39438);
nor U41228 (N_41228,N_39577,N_38168);
xor U41229 (N_41229,N_38597,N_37607);
xor U41230 (N_41230,N_38431,N_38540);
or U41231 (N_41231,N_38038,N_38121);
and U41232 (N_41232,N_38036,N_39336);
nor U41233 (N_41233,N_39697,N_37815);
xnor U41234 (N_41234,N_37508,N_38532);
xor U41235 (N_41235,N_38977,N_37786);
xor U41236 (N_41236,N_38611,N_38773);
xor U41237 (N_41237,N_38908,N_38656);
nor U41238 (N_41238,N_37649,N_39986);
or U41239 (N_41239,N_38353,N_38457);
xnor U41240 (N_41240,N_37735,N_38434);
nand U41241 (N_41241,N_39802,N_38349);
and U41242 (N_41242,N_38049,N_37927);
and U41243 (N_41243,N_39469,N_38016);
nor U41244 (N_41244,N_39979,N_37759);
nand U41245 (N_41245,N_39919,N_39561);
and U41246 (N_41246,N_39191,N_38516);
xor U41247 (N_41247,N_38244,N_38162);
nor U41248 (N_41248,N_38443,N_39470);
xnor U41249 (N_41249,N_38768,N_38601);
nand U41250 (N_41250,N_37937,N_39944);
and U41251 (N_41251,N_39502,N_38212);
nor U41252 (N_41252,N_39389,N_39503);
or U41253 (N_41253,N_39250,N_38834);
or U41254 (N_41254,N_39598,N_39130);
and U41255 (N_41255,N_39773,N_37886);
nand U41256 (N_41256,N_38839,N_38405);
and U41257 (N_41257,N_39538,N_37797);
xnor U41258 (N_41258,N_37655,N_38704);
nor U41259 (N_41259,N_37844,N_39100);
xnor U41260 (N_41260,N_37706,N_37556);
or U41261 (N_41261,N_38573,N_39826);
and U41262 (N_41262,N_39536,N_38889);
xor U41263 (N_41263,N_39645,N_39223);
xnor U41264 (N_41264,N_38322,N_39669);
xnor U41265 (N_41265,N_39474,N_38164);
nor U41266 (N_41266,N_39356,N_39741);
or U41267 (N_41267,N_39708,N_38786);
nand U41268 (N_41268,N_39280,N_39810);
or U41269 (N_41269,N_39556,N_38748);
or U41270 (N_41270,N_37839,N_39983);
xor U41271 (N_41271,N_38202,N_37646);
xor U41272 (N_41272,N_38602,N_37813);
nor U41273 (N_41273,N_38015,N_38334);
or U41274 (N_41274,N_37511,N_39203);
or U41275 (N_41275,N_39536,N_37788);
and U41276 (N_41276,N_39454,N_39549);
nor U41277 (N_41277,N_39115,N_37788);
nor U41278 (N_41278,N_38355,N_37662);
and U41279 (N_41279,N_38870,N_39085);
and U41280 (N_41280,N_38364,N_38737);
and U41281 (N_41281,N_39429,N_39780);
and U41282 (N_41282,N_39903,N_38586);
nand U41283 (N_41283,N_39983,N_39966);
nand U41284 (N_41284,N_39836,N_39353);
nor U41285 (N_41285,N_39382,N_37873);
nand U41286 (N_41286,N_38420,N_37894);
nor U41287 (N_41287,N_39131,N_38565);
nand U41288 (N_41288,N_38174,N_39155);
nand U41289 (N_41289,N_38324,N_37548);
and U41290 (N_41290,N_37840,N_39931);
and U41291 (N_41291,N_39272,N_38473);
nand U41292 (N_41292,N_39637,N_39265);
nor U41293 (N_41293,N_38303,N_39758);
and U41294 (N_41294,N_39636,N_38889);
and U41295 (N_41295,N_39396,N_37615);
nand U41296 (N_41296,N_38351,N_39020);
and U41297 (N_41297,N_37843,N_39778);
or U41298 (N_41298,N_37505,N_38678);
xor U41299 (N_41299,N_39183,N_38614);
nor U41300 (N_41300,N_39696,N_37985);
xnor U41301 (N_41301,N_37813,N_38761);
nand U41302 (N_41302,N_38072,N_38768);
or U41303 (N_41303,N_39969,N_39909);
nand U41304 (N_41304,N_38937,N_38510);
nor U41305 (N_41305,N_38036,N_39433);
nand U41306 (N_41306,N_38509,N_39920);
or U41307 (N_41307,N_38920,N_38841);
nand U41308 (N_41308,N_37620,N_38565);
and U41309 (N_41309,N_38167,N_39744);
nor U41310 (N_41310,N_38053,N_38511);
or U41311 (N_41311,N_37921,N_38717);
xnor U41312 (N_41312,N_39185,N_37754);
or U41313 (N_41313,N_39100,N_38130);
xor U41314 (N_41314,N_39850,N_38992);
xnor U41315 (N_41315,N_39132,N_38699);
xnor U41316 (N_41316,N_39490,N_37562);
xnor U41317 (N_41317,N_38261,N_39799);
and U41318 (N_41318,N_39705,N_39596);
nand U41319 (N_41319,N_38081,N_38867);
nand U41320 (N_41320,N_39986,N_38852);
xnor U41321 (N_41321,N_37791,N_39578);
or U41322 (N_41322,N_37820,N_39219);
and U41323 (N_41323,N_38977,N_39456);
xnor U41324 (N_41324,N_39527,N_38889);
xnor U41325 (N_41325,N_39806,N_38056);
nand U41326 (N_41326,N_38825,N_38028);
and U41327 (N_41327,N_38009,N_37869);
nand U41328 (N_41328,N_39212,N_39925);
nand U41329 (N_41329,N_37612,N_38417);
nor U41330 (N_41330,N_38408,N_37903);
xnor U41331 (N_41331,N_38157,N_38432);
xor U41332 (N_41332,N_37642,N_37552);
and U41333 (N_41333,N_39591,N_38474);
nand U41334 (N_41334,N_39987,N_38727);
or U41335 (N_41335,N_39385,N_38078);
nand U41336 (N_41336,N_39647,N_38828);
or U41337 (N_41337,N_38739,N_37962);
nand U41338 (N_41338,N_38971,N_39335);
or U41339 (N_41339,N_38252,N_39479);
and U41340 (N_41340,N_39031,N_39947);
nor U41341 (N_41341,N_37833,N_38101);
and U41342 (N_41342,N_39842,N_37678);
and U41343 (N_41343,N_37722,N_38409);
nand U41344 (N_41344,N_37921,N_38567);
or U41345 (N_41345,N_38126,N_38051);
xnor U41346 (N_41346,N_39221,N_37630);
xor U41347 (N_41347,N_38377,N_38280);
or U41348 (N_41348,N_38065,N_39641);
nor U41349 (N_41349,N_39013,N_38191);
and U41350 (N_41350,N_39401,N_37502);
nor U41351 (N_41351,N_39728,N_39717);
or U41352 (N_41352,N_37638,N_37633);
nand U41353 (N_41353,N_39920,N_39149);
xor U41354 (N_41354,N_37806,N_39560);
nand U41355 (N_41355,N_39819,N_39919);
nor U41356 (N_41356,N_39960,N_39598);
xnor U41357 (N_41357,N_38350,N_38398);
and U41358 (N_41358,N_39145,N_39688);
nand U41359 (N_41359,N_39482,N_39059);
nand U41360 (N_41360,N_38421,N_38518);
nand U41361 (N_41361,N_38048,N_38291);
nand U41362 (N_41362,N_37568,N_39968);
and U41363 (N_41363,N_38033,N_39880);
or U41364 (N_41364,N_38691,N_38729);
or U41365 (N_41365,N_39032,N_39122);
and U41366 (N_41366,N_39207,N_37784);
nor U41367 (N_41367,N_37648,N_38014);
nor U41368 (N_41368,N_38021,N_39116);
or U41369 (N_41369,N_38841,N_38110);
and U41370 (N_41370,N_37982,N_38239);
or U41371 (N_41371,N_38762,N_39223);
nand U41372 (N_41372,N_37998,N_39366);
and U41373 (N_41373,N_39847,N_38390);
and U41374 (N_41374,N_37713,N_38128);
xor U41375 (N_41375,N_38556,N_38725);
or U41376 (N_41376,N_39651,N_39720);
xor U41377 (N_41377,N_39655,N_37609);
and U41378 (N_41378,N_38953,N_39137);
nor U41379 (N_41379,N_37665,N_37946);
nand U41380 (N_41380,N_39779,N_39069);
or U41381 (N_41381,N_37666,N_38189);
or U41382 (N_41382,N_39282,N_39003);
xor U41383 (N_41383,N_39388,N_37954);
or U41384 (N_41384,N_37909,N_39771);
and U41385 (N_41385,N_38741,N_38250);
nand U41386 (N_41386,N_39710,N_38730);
nor U41387 (N_41387,N_39964,N_39786);
or U41388 (N_41388,N_39407,N_39182);
or U41389 (N_41389,N_39427,N_39513);
nor U41390 (N_41390,N_39219,N_39945);
and U41391 (N_41391,N_38813,N_37683);
and U41392 (N_41392,N_38873,N_38861);
xor U41393 (N_41393,N_38929,N_37503);
xnor U41394 (N_41394,N_38389,N_39060);
and U41395 (N_41395,N_39550,N_39277);
nand U41396 (N_41396,N_39702,N_38205);
nand U41397 (N_41397,N_38992,N_39223);
or U41398 (N_41398,N_39611,N_38469);
nor U41399 (N_41399,N_39708,N_39909);
and U41400 (N_41400,N_37907,N_38835);
and U41401 (N_41401,N_37612,N_38646);
nor U41402 (N_41402,N_38615,N_38295);
and U41403 (N_41403,N_39374,N_39276);
nor U41404 (N_41404,N_39097,N_39002);
and U41405 (N_41405,N_39057,N_37592);
nor U41406 (N_41406,N_37948,N_38058);
xor U41407 (N_41407,N_37570,N_37596);
nand U41408 (N_41408,N_38256,N_39292);
xor U41409 (N_41409,N_38829,N_38527);
nand U41410 (N_41410,N_39110,N_38954);
nand U41411 (N_41411,N_37795,N_39472);
xnor U41412 (N_41412,N_39537,N_38858);
or U41413 (N_41413,N_37590,N_37672);
or U41414 (N_41414,N_38174,N_37572);
nand U41415 (N_41415,N_37686,N_39061);
nand U41416 (N_41416,N_38537,N_39168);
and U41417 (N_41417,N_37945,N_38793);
or U41418 (N_41418,N_39584,N_39744);
xnor U41419 (N_41419,N_38932,N_39373);
or U41420 (N_41420,N_37761,N_38411);
xnor U41421 (N_41421,N_39565,N_38532);
xor U41422 (N_41422,N_39251,N_38461);
nor U41423 (N_41423,N_38549,N_39632);
xor U41424 (N_41424,N_38084,N_37652);
nand U41425 (N_41425,N_39612,N_39631);
xor U41426 (N_41426,N_38801,N_38665);
nor U41427 (N_41427,N_38731,N_39853);
and U41428 (N_41428,N_38409,N_39640);
nand U41429 (N_41429,N_39361,N_38295);
and U41430 (N_41430,N_37779,N_39037);
nor U41431 (N_41431,N_39402,N_37993);
or U41432 (N_41432,N_38271,N_39890);
and U41433 (N_41433,N_38333,N_38722);
nand U41434 (N_41434,N_39652,N_37814);
xor U41435 (N_41435,N_38428,N_38044);
xor U41436 (N_41436,N_37614,N_37797);
nand U41437 (N_41437,N_37828,N_38808);
or U41438 (N_41438,N_37696,N_38481);
or U41439 (N_41439,N_38894,N_38779);
and U41440 (N_41440,N_38931,N_38951);
nand U41441 (N_41441,N_38311,N_38937);
or U41442 (N_41442,N_38694,N_37767);
xor U41443 (N_41443,N_39919,N_37521);
xor U41444 (N_41444,N_39531,N_38335);
or U41445 (N_41445,N_38467,N_38294);
and U41446 (N_41446,N_38821,N_37507);
nand U41447 (N_41447,N_38891,N_38492);
and U41448 (N_41448,N_38170,N_39858);
or U41449 (N_41449,N_37642,N_38627);
xnor U41450 (N_41450,N_37719,N_38906);
or U41451 (N_41451,N_39318,N_39183);
nor U41452 (N_41452,N_38542,N_38632);
nand U41453 (N_41453,N_39758,N_39279);
and U41454 (N_41454,N_39851,N_39644);
and U41455 (N_41455,N_38731,N_37795);
nand U41456 (N_41456,N_37722,N_37976);
nand U41457 (N_41457,N_39580,N_39028);
xnor U41458 (N_41458,N_37763,N_39888);
or U41459 (N_41459,N_39848,N_38593);
nor U41460 (N_41460,N_39375,N_39427);
or U41461 (N_41461,N_39664,N_37886);
and U41462 (N_41462,N_38602,N_38795);
or U41463 (N_41463,N_39599,N_38673);
and U41464 (N_41464,N_37726,N_39463);
nand U41465 (N_41465,N_38360,N_39973);
and U41466 (N_41466,N_38395,N_39539);
nand U41467 (N_41467,N_39952,N_38680);
or U41468 (N_41468,N_37823,N_39705);
and U41469 (N_41469,N_38204,N_39029);
or U41470 (N_41470,N_38816,N_38386);
or U41471 (N_41471,N_39262,N_39517);
nand U41472 (N_41472,N_38862,N_38813);
xor U41473 (N_41473,N_37712,N_37690);
nor U41474 (N_41474,N_38770,N_39689);
and U41475 (N_41475,N_38972,N_39164);
nand U41476 (N_41476,N_39013,N_38256);
nand U41477 (N_41477,N_37531,N_38925);
nand U41478 (N_41478,N_37626,N_38160);
or U41479 (N_41479,N_38144,N_38836);
nor U41480 (N_41480,N_39290,N_39242);
nor U41481 (N_41481,N_39725,N_37979);
nor U41482 (N_41482,N_39301,N_38547);
nand U41483 (N_41483,N_38104,N_39592);
nor U41484 (N_41484,N_39344,N_39166);
and U41485 (N_41485,N_39146,N_37679);
or U41486 (N_41486,N_39477,N_39303);
nand U41487 (N_41487,N_39404,N_38868);
and U41488 (N_41488,N_38639,N_39304);
nor U41489 (N_41489,N_37792,N_39824);
or U41490 (N_41490,N_37698,N_37949);
and U41491 (N_41491,N_39268,N_37540);
nor U41492 (N_41492,N_37780,N_39728);
nor U41493 (N_41493,N_38207,N_38730);
and U41494 (N_41494,N_39027,N_38533);
and U41495 (N_41495,N_38377,N_39339);
nand U41496 (N_41496,N_38754,N_39258);
xor U41497 (N_41497,N_39961,N_38499);
or U41498 (N_41498,N_39053,N_39698);
or U41499 (N_41499,N_39881,N_38882);
xnor U41500 (N_41500,N_38832,N_37924);
nor U41501 (N_41501,N_38714,N_38848);
xor U41502 (N_41502,N_39059,N_39612);
nor U41503 (N_41503,N_39320,N_38522);
and U41504 (N_41504,N_38749,N_39167);
xor U41505 (N_41505,N_39735,N_37708);
and U41506 (N_41506,N_38992,N_39922);
xor U41507 (N_41507,N_39275,N_38838);
xnor U41508 (N_41508,N_38545,N_39616);
xnor U41509 (N_41509,N_39932,N_38206);
nor U41510 (N_41510,N_38037,N_38148);
xnor U41511 (N_41511,N_37906,N_39119);
nor U41512 (N_41512,N_37946,N_38545);
xnor U41513 (N_41513,N_38267,N_39566);
nand U41514 (N_41514,N_39095,N_38165);
nand U41515 (N_41515,N_37935,N_37999);
and U41516 (N_41516,N_39737,N_37778);
or U41517 (N_41517,N_39367,N_38938);
nand U41518 (N_41518,N_39480,N_39592);
nor U41519 (N_41519,N_39165,N_39398);
or U41520 (N_41520,N_37691,N_38879);
nand U41521 (N_41521,N_38553,N_39303);
xor U41522 (N_41522,N_38355,N_39334);
and U41523 (N_41523,N_38844,N_38625);
nor U41524 (N_41524,N_39008,N_38797);
and U41525 (N_41525,N_38515,N_38217);
nor U41526 (N_41526,N_39048,N_37950);
nand U41527 (N_41527,N_38642,N_38433);
and U41528 (N_41528,N_39076,N_37725);
nor U41529 (N_41529,N_37988,N_38436);
nand U41530 (N_41530,N_39228,N_37585);
or U41531 (N_41531,N_38591,N_38926);
xor U41532 (N_41532,N_37661,N_37533);
and U41533 (N_41533,N_38190,N_37959);
and U41534 (N_41534,N_38389,N_39620);
xnor U41535 (N_41535,N_38977,N_37556);
or U41536 (N_41536,N_38176,N_37913);
nand U41537 (N_41537,N_37521,N_37608);
or U41538 (N_41538,N_39059,N_39101);
or U41539 (N_41539,N_39776,N_39902);
or U41540 (N_41540,N_38236,N_39505);
xnor U41541 (N_41541,N_37778,N_38575);
nand U41542 (N_41542,N_39549,N_38670);
nand U41543 (N_41543,N_39842,N_39621);
xor U41544 (N_41544,N_38063,N_38052);
nor U41545 (N_41545,N_38853,N_37902);
xnor U41546 (N_41546,N_38189,N_39817);
and U41547 (N_41547,N_38448,N_37983);
xnor U41548 (N_41548,N_38610,N_38001);
xor U41549 (N_41549,N_38698,N_39948);
and U41550 (N_41550,N_39087,N_38497);
or U41551 (N_41551,N_38609,N_38111);
and U41552 (N_41552,N_38766,N_38859);
nand U41553 (N_41553,N_39374,N_38716);
nand U41554 (N_41554,N_38022,N_38073);
nand U41555 (N_41555,N_37963,N_39135);
and U41556 (N_41556,N_38988,N_39635);
or U41557 (N_41557,N_38377,N_38772);
nor U41558 (N_41558,N_38551,N_39182);
xnor U41559 (N_41559,N_39844,N_39516);
or U41560 (N_41560,N_39108,N_37642);
or U41561 (N_41561,N_39668,N_39714);
xor U41562 (N_41562,N_39597,N_37850);
and U41563 (N_41563,N_38107,N_39836);
nor U41564 (N_41564,N_37587,N_39928);
nor U41565 (N_41565,N_38521,N_38921);
nand U41566 (N_41566,N_37691,N_37828);
or U41567 (N_41567,N_39289,N_39574);
and U41568 (N_41568,N_37717,N_39469);
or U41569 (N_41569,N_37507,N_39092);
nand U41570 (N_41570,N_39471,N_37865);
or U41571 (N_41571,N_37860,N_38033);
and U41572 (N_41572,N_38562,N_37641);
or U41573 (N_41573,N_38181,N_37542);
nand U41574 (N_41574,N_39637,N_39896);
and U41575 (N_41575,N_39417,N_38660);
nor U41576 (N_41576,N_39660,N_37940);
or U41577 (N_41577,N_39027,N_38762);
and U41578 (N_41578,N_39829,N_38062);
or U41579 (N_41579,N_39386,N_37615);
xor U41580 (N_41580,N_38816,N_38339);
xor U41581 (N_41581,N_39399,N_38331);
xnor U41582 (N_41582,N_39409,N_37685);
or U41583 (N_41583,N_38432,N_39754);
and U41584 (N_41584,N_38085,N_37621);
or U41585 (N_41585,N_38759,N_39909);
and U41586 (N_41586,N_39247,N_39320);
or U41587 (N_41587,N_37884,N_38434);
xor U41588 (N_41588,N_39649,N_39962);
nor U41589 (N_41589,N_39700,N_38391);
and U41590 (N_41590,N_39068,N_38264);
nor U41591 (N_41591,N_39462,N_37745);
nor U41592 (N_41592,N_39149,N_39421);
nand U41593 (N_41593,N_38762,N_38447);
xor U41594 (N_41594,N_39359,N_37863);
and U41595 (N_41595,N_38405,N_39842);
nor U41596 (N_41596,N_38692,N_39039);
nand U41597 (N_41597,N_38420,N_37619);
or U41598 (N_41598,N_39109,N_39349);
or U41599 (N_41599,N_37553,N_37664);
nand U41600 (N_41600,N_39577,N_39648);
and U41601 (N_41601,N_37918,N_38108);
nand U41602 (N_41602,N_38416,N_39411);
nor U41603 (N_41603,N_39633,N_39458);
xnor U41604 (N_41604,N_38159,N_39915);
nor U41605 (N_41605,N_38930,N_38045);
xor U41606 (N_41606,N_38131,N_39069);
or U41607 (N_41607,N_39527,N_37872);
nand U41608 (N_41608,N_38354,N_37683);
and U41609 (N_41609,N_39829,N_39360);
nor U41610 (N_41610,N_37613,N_38802);
or U41611 (N_41611,N_39317,N_37714);
or U41612 (N_41612,N_38772,N_38839);
or U41613 (N_41613,N_38322,N_39599);
or U41614 (N_41614,N_38370,N_39469);
or U41615 (N_41615,N_37558,N_38163);
nand U41616 (N_41616,N_38854,N_38185);
nand U41617 (N_41617,N_37751,N_39728);
and U41618 (N_41618,N_39039,N_38881);
or U41619 (N_41619,N_38135,N_38241);
and U41620 (N_41620,N_39808,N_38585);
nor U41621 (N_41621,N_39305,N_39637);
xor U41622 (N_41622,N_38214,N_37595);
and U41623 (N_41623,N_38799,N_37672);
nor U41624 (N_41624,N_37795,N_39812);
nor U41625 (N_41625,N_37957,N_39926);
nand U41626 (N_41626,N_38021,N_37824);
xor U41627 (N_41627,N_37832,N_37916);
nand U41628 (N_41628,N_39229,N_39301);
xor U41629 (N_41629,N_38139,N_38396);
nand U41630 (N_41630,N_38894,N_37961);
nand U41631 (N_41631,N_39915,N_38763);
and U41632 (N_41632,N_37735,N_37521);
nand U41633 (N_41633,N_39162,N_38589);
xor U41634 (N_41634,N_39519,N_37973);
nand U41635 (N_41635,N_39678,N_39242);
nor U41636 (N_41636,N_38100,N_37550);
nand U41637 (N_41637,N_38236,N_39334);
or U41638 (N_41638,N_38137,N_37672);
or U41639 (N_41639,N_39423,N_39035);
xor U41640 (N_41640,N_38845,N_38808);
nand U41641 (N_41641,N_39584,N_38051);
nand U41642 (N_41642,N_37613,N_37695);
xor U41643 (N_41643,N_39509,N_39712);
or U41644 (N_41644,N_39556,N_39922);
nor U41645 (N_41645,N_38363,N_37798);
nand U41646 (N_41646,N_39130,N_37877);
or U41647 (N_41647,N_37698,N_38067);
and U41648 (N_41648,N_37638,N_38141);
and U41649 (N_41649,N_39004,N_37923);
or U41650 (N_41650,N_38036,N_39965);
xnor U41651 (N_41651,N_39705,N_38824);
and U41652 (N_41652,N_39054,N_39739);
or U41653 (N_41653,N_39014,N_39674);
nand U41654 (N_41654,N_38326,N_39004);
nor U41655 (N_41655,N_37799,N_39579);
or U41656 (N_41656,N_39804,N_38472);
and U41657 (N_41657,N_38159,N_39330);
nand U41658 (N_41658,N_38562,N_38704);
nor U41659 (N_41659,N_38579,N_37873);
xnor U41660 (N_41660,N_37779,N_39012);
nor U41661 (N_41661,N_37879,N_37678);
nor U41662 (N_41662,N_38265,N_38038);
and U41663 (N_41663,N_39973,N_39596);
and U41664 (N_41664,N_37763,N_39566);
and U41665 (N_41665,N_38732,N_38744);
nand U41666 (N_41666,N_38433,N_37970);
nor U41667 (N_41667,N_38170,N_39983);
nand U41668 (N_41668,N_38444,N_38733);
xor U41669 (N_41669,N_39376,N_38593);
xnor U41670 (N_41670,N_38574,N_37947);
xor U41671 (N_41671,N_39886,N_39387);
nand U41672 (N_41672,N_39610,N_38711);
nand U41673 (N_41673,N_37780,N_39420);
or U41674 (N_41674,N_38317,N_39852);
or U41675 (N_41675,N_39448,N_37907);
or U41676 (N_41676,N_38804,N_39165);
or U41677 (N_41677,N_39042,N_38949);
nand U41678 (N_41678,N_38488,N_39275);
nand U41679 (N_41679,N_39390,N_39074);
nor U41680 (N_41680,N_39023,N_39063);
or U41681 (N_41681,N_38725,N_39878);
or U41682 (N_41682,N_39042,N_39774);
or U41683 (N_41683,N_39574,N_39942);
and U41684 (N_41684,N_39868,N_39697);
nor U41685 (N_41685,N_39895,N_38280);
or U41686 (N_41686,N_39420,N_38649);
or U41687 (N_41687,N_39994,N_38659);
or U41688 (N_41688,N_39043,N_39060);
or U41689 (N_41689,N_39171,N_38042);
nor U41690 (N_41690,N_39737,N_38443);
nand U41691 (N_41691,N_37710,N_39713);
nor U41692 (N_41692,N_37578,N_39086);
nand U41693 (N_41693,N_39002,N_39015);
nor U41694 (N_41694,N_39056,N_39882);
nand U41695 (N_41695,N_38415,N_39388);
nor U41696 (N_41696,N_37755,N_37933);
nor U41697 (N_41697,N_38691,N_38766);
or U41698 (N_41698,N_37766,N_37518);
xor U41699 (N_41699,N_37623,N_37778);
nand U41700 (N_41700,N_38734,N_37927);
nand U41701 (N_41701,N_39350,N_38297);
and U41702 (N_41702,N_38563,N_39718);
nand U41703 (N_41703,N_37532,N_38494);
and U41704 (N_41704,N_38660,N_39541);
nand U41705 (N_41705,N_38595,N_38023);
or U41706 (N_41706,N_39679,N_39691);
nor U41707 (N_41707,N_38402,N_37786);
nor U41708 (N_41708,N_38633,N_37651);
nor U41709 (N_41709,N_38461,N_37947);
xnor U41710 (N_41710,N_38913,N_39171);
nand U41711 (N_41711,N_39663,N_38384);
nand U41712 (N_41712,N_37642,N_39798);
nand U41713 (N_41713,N_39910,N_37709);
nand U41714 (N_41714,N_39625,N_39740);
nor U41715 (N_41715,N_38801,N_38399);
and U41716 (N_41716,N_39042,N_38169);
nor U41717 (N_41717,N_38830,N_37821);
xnor U41718 (N_41718,N_39075,N_38209);
xor U41719 (N_41719,N_39772,N_38025);
and U41720 (N_41720,N_37978,N_37757);
nor U41721 (N_41721,N_39430,N_39996);
nand U41722 (N_41722,N_38914,N_38550);
and U41723 (N_41723,N_38100,N_38490);
or U41724 (N_41724,N_38389,N_38845);
xor U41725 (N_41725,N_38591,N_38030);
and U41726 (N_41726,N_38751,N_38425);
nand U41727 (N_41727,N_39704,N_39122);
and U41728 (N_41728,N_39985,N_38832);
xnor U41729 (N_41729,N_38733,N_38743);
nor U41730 (N_41730,N_39563,N_38940);
or U41731 (N_41731,N_38162,N_38128);
nor U41732 (N_41732,N_38462,N_38397);
nand U41733 (N_41733,N_39271,N_39313);
and U41734 (N_41734,N_38571,N_39571);
nor U41735 (N_41735,N_39917,N_38733);
xnor U41736 (N_41736,N_38488,N_38496);
nor U41737 (N_41737,N_37812,N_38075);
and U41738 (N_41738,N_37965,N_39420);
or U41739 (N_41739,N_39575,N_39063);
nor U41740 (N_41740,N_38735,N_38262);
xor U41741 (N_41741,N_39391,N_38008);
nand U41742 (N_41742,N_37689,N_39776);
xor U41743 (N_41743,N_39684,N_39913);
nand U41744 (N_41744,N_38100,N_38921);
or U41745 (N_41745,N_38956,N_39752);
nor U41746 (N_41746,N_37854,N_37880);
or U41747 (N_41747,N_38119,N_37878);
nor U41748 (N_41748,N_38425,N_38456);
xnor U41749 (N_41749,N_38428,N_38736);
nand U41750 (N_41750,N_37931,N_38233);
and U41751 (N_41751,N_38717,N_39361);
or U41752 (N_41752,N_38606,N_38303);
xor U41753 (N_41753,N_38010,N_39018);
nor U41754 (N_41754,N_37675,N_38173);
or U41755 (N_41755,N_37717,N_39484);
xor U41756 (N_41756,N_39773,N_39077);
nand U41757 (N_41757,N_39056,N_38385);
nor U41758 (N_41758,N_39260,N_38770);
or U41759 (N_41759,N_39411,N_39126);
xnor U41760 (N_41760,N_38864,N_39174);
nand U41761 (N_41761,N_37909,N_38699);
nor U41762 (N_41762,N_38708,N_39595);
and U41763 (N_41763,N_39113,N_39630);
nand U41764 (N_41764,N_38644,N_39622);
nand U41765 (N_41765,N_39921,N_37913);
nor U41766 (N_41766,N_38886,N_38127);
nor U41767 (N_41767,N_38653,N_38632);
nand U41768 (N_41768,N_37991,N_38346);
nor U41769 (N_41769,N_37747,N_39845);
or U41770 (N_41770,N_38640,N_39868);
or U41771 (N_41771,N_39148,N_39448);
nor U41772 (N_41772,N_39613,N_38255);
xnor U41773 (N_41773,N_39193,N_39210);
nand U41774 (N_41774,N_37617,N_39267);
or U41775 (N_41775,N_38218,N_38850);
nand U41776 (N_41776,N_37559,N_38646);
nand U41777 (N_41777,N_38441,N_38930);
or U41778 (N_41778,N_38256,N_38488);
or U41779 (N_41779,N_38621,N_38453);
nor U41780 (N_41780,N_37689,N_37535);
nor U41781 (N_41781,N_38401,N_37538);
nor U41782 (N_41782,N_39399,N_39580);
and U41783 (N_41783,N_39368,N_39225);
nand U41784 (N_41784,N_38402,N_38392);
nor U41785 (N_41785,N_39745,N_39506);
xor U41786 (N_41786,N_38796,N_39578);
nand U41787 (N_41787,N_39355,N_38545);
nand U41788 (N_41788,N_39948,N_38747);
xor U41789 (N_41789,N_38825,N_39102);
xnor U41790 (N_41790,N_38734,N_39422);
nand U41791 (N_41791,N_37595,N_39925);
or U41792 (N_41792,N_38210,N_38965);
xor U41793 (N_41793,N_39472,N_38006);
xor U41794 (N_41794,N_38489,N_38459);
nor U41795 (N_41795,N_38681,N_38953);
and U41796 (N_41796,N_39510,N_39444);
nor U41797 (N_41797,N_38905,N_38410);
xnor U41798 (N_41798,N_37967,N_39328);
nor U41799 (N_41799,N_37816,N_39321);
xor U41800 (N_41800,N_39213,N_39124);
nand U41801 (N_41801,N_39579,N_37960);
xnor U41802 (N_41802,N_37898,N_39279);
or U41803 (N_41803,N_38001,N_38187);
and U41804 (N_41804,N_38078,N_39754);
or U41805 (N_41805,N_39370,N_39455);
nor U41806 (N_41806,N_38714,N_38135);
and U41807 (N_41807,N_39793,N_38139);
xor U41808 (N_41808,N_37761,N_38546);
nand U41809 (N_41809,N_37533,N_38657);
or U41810 (N_41810,N_38012,N_38353);
and U41811 (N_41811,N_38835,N_38733);
xnor U41812 (N_41812,N_38755,N_39270);
and U41813 (N_41813,N_39214,N_38882);
and U41814 (N_41814,N_38689,N_39599);
nor U41815 (N_41815,N_39278,N_37524);
or U41816 (N_41816,N_38181,N_38942);
xnor U41817 (N_41817,N_37673,N_39884);
xor U41818 (N_41818,N_37902,N_37602);
xnor U41819 (N_41819,N_39263,N_39691);
xor U41820 (N_41820,N_38444,N_38698);
nor U41821 (N_41821,N_37927,N_38742);
and U41822 (N_41822,N_39703,N_38860);
nor U41823 (N_41823,N_37535,N_38855);
nand U41824 (N_41824,N_37573,N_39719);
and U41825 (N_41825,N_37557,N_39711);
nand U41826 (N_41826,N_37506,N_37848);
xnor U41827 (N_41827,N_38446,N_38090);
xor U41828 (N_41828,N_39360,N_38364);
or U41829 (N_41829,N_39226,N_39325);
nand U41830 (N_41830,N_38125,N_39502);
and U41831 (N_41831,N_39971,N_37613);
nor U41832 (N_41832,N_38269,N_38099);
and U41833 (N_41833,N_37712,N_39671);
and U41834 (N_41834,N_38863,N_38011);
nand U41835 (N_41835,N_38553,N_37604);
or U41836 (N_41836,N_38078,N_38639);
nor U41837 (N_41837,N_39292,N_38323);
xnor U41838 (N_41838,N_39435,N_37582);
or U41839 (N_41839,N_38202,N_39303);
and U41840 (N_41840,N_37666,N_39217);
xor U41841 (N_41841,N_39122,N_39246);
nor U41842 (N_41842,N_38607,N_39649);
and U41843 (N_41843,N_37533,N_39016);
or U41844 (N_41844,N_39049,N_39742);
nand U41845 (N_41845,N_39858,N_38392);
nand U41846 (N_41846,N_39609,N_39719);
nand U41847 (N_41847,N_37923,N_38313);
nor U41848 (N_41848,N_39558,N_39826);
nor U41849 (N_41849,N_39849,N_37663);
nand U41850 (N_41850,N_39084,N_38289);
or U41851 (N_41851,N_39431,N_38274);
xnor U41852 (N_41852,N_39542,N_37814);
nor U41853 (N_41853,N_38327,N_38983);
nor U41854 (N_41854,N_38137,N_39641);
nand U41855 (N_41855,N_39720,N_37764);
nand U41856 (N_41856,N_37583,N_39621);
xnor U41857 (N_41857,N_39042,N_38127);
nand U41858 (N_41858,N_38140,N_39123);
xnor U41859 (N_41859,N_38035,N_39555);
and U41860 (N_41860,N_37698,N_39528);
xor U41861 (N_41861,N_38712,N_38274);
xnor U41862 (N_41862,N_38918,N_38637);
xnor U41863 (N_41863,N_38972,N_37813);
nor U41864 (N_41864,N_39645,N_37995);
nand U41865 (N_41865,N_38143,N_39317);
and U41866 (N_41866,N_38622,N_39232);
nor U41867 (N_41867,N_38017,N_39949);
xnor U41868 (N_41868,N_37575,N_38423);
and U41869 (N_41869,N_39574,N_39889);
or U41870 (N_41870,N_38103,N_37829);
nand U41871 (N_41871,N_39099,N_37669);
nor U41872 (N_41872,N_39319,N_38768);
xor U41873 (N_41873,N_38214,N_39021);
and U41874 (N_41874,N_37823,N_38276);
xnor U41875 (N_41875,N_39709,N_39182);
nand U41876 (N_41876,N_39063,N_38981);
or U41877 (N_41877,N_37880,N_39898);
nor U41878 (N_41878,N_38530,N_37981);
nand U41879 (N_41879,N_37690,N_39999);
nor U41880 (N_41880,N_38513,N_38494);
nor U41881 (N_41881,N_38343,N_38557);
nand U41882 (N_41882,N_39926,N_37659);
and U41883 (N_41883,N_38951,N_38810);
nor U41884 (N_41884,N_38416,N_37980);
or U41885 (N_41885,N_39902,N_39886);
xor U41886 (N_41886,N_38117,N_38800);
nand U41887 (N_41887,N_39751,N_39366);
nor U41888 (N_41888,N_38176,N_39259);
xnor U41889 (N_41889,N_39196,N_38864);
and U41890 (N_41890,N_39059,N_38283);
nand U41891 (N_41891,N_38395,N_38901);
nand U41892 (N_41892,N_39238,N_39312);
and U41893 (N_41893,N_39946,N_39732);
nor U41894 (N_41894,N_39390,N_37684);
and U41895 (N_41895,N_38099,N_37731);
xor U41896 (N_41896,N_37709,N_39683);
and U41897 (N_41897,N_37829,N_39446);
xnor U41898 (N_41898,N_38323,N_39799);
and U41899 (N_41899,N_39238,N_38331);
or U41900 (N_41900,N_39824,N_38012);
and U41901 (N_41901,N_38608,N_39320);
xnor U41902 (N_41902,N_38922,N_38597);
xor U41903 (N_41903,N_39314,N_38175);
nand U41904 (N_41904,N_37792,N_39854);
or U41905 (N_41905,N_38972,N_39120);
and U41906 (N_41906,N_39066,N_37776);
nor U41907 (N_41907,N_39216,N_39680);
and U41908 (N_41908,N_39298,N_37932);
nor U41909 (N_41909,N_37736,N_37974);
nand U41910 (N_41910,N_39444,N_38254);
nor U41911 (N_41911,N_38060,N_37915);
and U41912 (N_41912,N_39141,N_38764);
xnor U41913 (N_41913,N_39488,N_38383);
xor U41914 (N_41914,N_38723,N_37900);
xor U41915 (N_41915,N_39851,N_38174);
and U41916 (N_41916,N_38868,N_39683);
nand U41917 (N_41917,N_39826,N_39971);
or U41918 (N_41918,N_38739,N_39743);
or U41919 (N_41919,N_39852,N_39164);
nand U41920 (N_41920,N_38224,N_39587);
or U41921 (N_41921,N_39622,N_38376);
nand U41922 (N_41922,N_38109,N_38415);
or U41923 (N_41923,N_38788,N_38723);
and U41924 (N_41924,N_38433,N_39129);
nand U41925 (N_41925,N_39422,N_38288);
and U41926 (N_41926,N_39144,N_39214);
nand U41927 (N_41927,N_39113,N_38984);
nand U41928 (N_41928,N_38756,N_39198);
xor U41929 (N_41929,N_38658,N_39117);
nand U41930 (N_41930,N_37633,N_38401);
nand U41931 (N_41931,N_38307,N_38821);
and U41932 (N_41932,N_37511,N_38377);
xnor U41933 (N_41933,N_39100,N_38114);
nand U41934 (N_41934,N_39724,N_39581);
or U41935 (N_41935,N_37811,N_39143);
or U41936 (N_41936,N_38200,N_37805);
nand U41937 (N_41937,N_39738,N_37680);
xnor U41938 (N_41938,N_38148,N_37551);
and U41939 (N_41939,N_39918,N_39505);
xnor U41940 (N_41940,N_38368,N_39116);
nand U41941 (N_41941,N_39304,N_39378);
xnor U41942 (N_41942,N_38746,N_38689);
and U41943 (N_41943,N_39538,N_37720);
or U41944 (N_41944,N_39800,N_39745);
or U41945 (N_41945,N_38650,N_39841);
or U41946 (N_41946,N_37563,N_39125);
and U41947 (N_41947,N_39241,N_38809);
nor U41948 (N_41948,N_39770,N_38345);
nand U41949 (N_41949,N_39835,N_39394);
nand U41950 (N_41950,N_38571,N_37932);
xnor U41951 (N_41951,N_37863,N_39850);
and U41952 (N_41952,N_39430,N_39986);
or U41953 (N_41953,N_38191,N_39603);
or U41954 (N_41954,N_37910,N_38841);
nor U41955 (N_41955,N_38175,N_39444);
xnor U41956 (N_41956,N_39657,N_37701);
nand U41957 (N_41957,N_38625,N_39497);
and U41958 (N_41958,N_38616,N_39209);
nor U41959 (N_41959,N_39779,N_39704);
and U41960 (N_41960,N_38423,N_38218);
nor U41961 (N_41961,N_38007,N_38228);
nand U41962 (N_41962,N_38992,N_39338);
and U41963 (N_41963,N_39061,N_39898);
xnor U41964 (N_41964,N_39386,N_39058);
nand U41965 (N_41965,N_38964,N_38904);
or U41966 (N_41966,N_37905,N_37839);
or U41967 (N_41967,N_39149,N_39573);
or U41968 (N_41968,N_39468,N_39826);
xor U41969 (N_41969,N_38566,N_37957);
and U41970 (N_41970,N_37766,N_39077);
xnor U41971 (N_41971,N_39116,N_38809);
nor U41972 (N_41972,N_38589,N_38956);
nor U41973 (N_41973,N_38752,N_38229);
or U41974 (N_41974,N_38585,N_39428);
xnor U41975 (N_41975,N_38571,N_37528);
and U41976 (N_41976,N_39740,N_39552);
xor U41977 (N_41977,N_38598,N_38128);
xnor U41978 (N_41978,N_38125,N_39707);
nand U41979 (N_41979,N_39330,N_37692);
and U41980 (N_41980,N_38425,N_37523);
nand U41981 (N_41981,N_39618,N_37780);
nor U41982 (N_41982,N_38293,N_39578);
nor U41983 (N_41983,N_39654,N_39703);
or U41984 (N_41984,N_39401,N_38020);
xor U41985 (N_41985,N_38318,N_38713);
or U41986 (N_41986,N_38664,N_38907);
nor U41987 (N_41987,N_39745,N_39764);
or U41988 (N_41988,N_37932,N_39855);
nand U41989 (N_41989,N_37809,N_39383);
xor U41990 (N_41990,N_38094,N_38213);
nor U41991 (N_41991,N_38033,N_37822);
or U41992 (N_41992,N_37926,N_38178);
and U41993 (N_41993,N_38187,N_37661);
nand U41994 (N_41994,N_39292,N_39841);
nand U41995 (N_41995,N_37923,N_39022);
nor U41996 (N_41996,N_39551,N_39535);
or U41997 (N_41997,N_39003,N_37832);
nand U41998 (N_41998,N_39488,N_39211);
nand U41999 (N_41999,N_39446,N_37559);
xnor U42000 (N_42000,N_39304,N_39246);
nor U42001 (N_42001,N_38041,N_38700);
or U42002 (N_42002,N_39387,N_37538);
nor U42003 (N_42003,N_38680,N_39692);
xnor U42004 (N_42004,N_39421,N_37944);
xnor U42005 (N_42005,N_39733,N_39570);
xnor U42006 (N_42006,N_39326,N_37836);
nand U42007 (N_42007,N_38765,N_38372);
nor U42008 (N_42008,N_39263,N_37942);
xnor U42009 (N_42009,N_39309,N_38254);
nand U42010 (N_42010,N_39976,N_38049);
xor U42011 (N_42011,N_38574,N_37583);
nand U42012 (N_42012,N_38737,N_39789);
and U42013 (N_42013,N_37996,N_39663);
nand U42014 (N_42014,N_39621,N_37926);
or U42015 (N_42015,N_39608,N_39147);
or U42016 (N_42016,N_38635,N_38513);
nand U42017 (N_42017,N_37974,N_39262);
nor U42018 (N_42018,N_38230,N_39757);
nor U42019 (N_42019,N_39236,N_38052);
and U42020 (N_42020,N_39789,N_38199);
or U42021 (N_42021,N_38119,N_39937);
and U42022 (N_42022,N_37893,N_39774);
or U42023 (N_42023,N_39716,N_37533);
nand U42024 (N_42024,N_38569,N_39133);
nor U42025 (N_42025,N_39754,N_38192);
or U42026 (N_42026,N_38996,N_39745);
or U42027 (N_42027,N_38380,N_38712);
xnor U42028 (N_42028,N_39006,N_39939);
or U42029 (N_42029,N_39881,N_37568);
nor U42030 (N_42030,N_39905,N_38984);
or U42031 (N_42031,N_39108,N_39794);
or U42032 (N_42032,N_39660,N_39545);
xnor U42033 (N_42033,N_38357,N_37706);
nand U42034 (N_42034,N_38780,N_38948);
or U42035 (N_42035,N_39226,N_37620);
xor U42036 (N_42036,N_38788,N_38030);
and U42037 (N_42037,N_38875,N_37797);
xnor U42038 (N_42038,N_38496,N_37685);
nand U42039 (N_42039,N_39198,N_38531);
nor U42040 (N_42040,N_39969,N_38257);
nor U42041 (N_42041,N_38697,N_38125);
or U42042 (N_42042,N_38268,N_38777);
xnor U42043 (N_42043,N_37740,N_38337);
xnor U42044 (N_42044,N_39785,N_38012);
xnor U42045 (N_42045,N_39269,N_38459);
nand U42046 (N_42046,N_37767,N_39845);
xnor U42047 (N_42047,N_38053,N_38153);
xor U42048 (N_42048,N_39366,N_39835);
nor U42049 (N_42049,N_39027,N_39565);
or U42050 (N_42050,N_38131,N_39574);
or U42051 (N_42051,N_37707,N_39666);
and U42052 (N_42052,N_38726,N_38264);
or U42053 (N_42053,N_39970,N_37868);
nand U42054 (N_42054,N_39318,N_39886);
or U42055 (N_42055,N_39785,N_37824);
or U42056 (N_42056,N_37991,N_38438);
xor U42057 (N_42057,N_38791,N_38945);
and U42058 (N_42058,N_38572,N_38722);
xnor U42059 (N_42059,N_39403,N_38052);
nand U42060 (N_42060,N_37975,N_38599);
or U42061 (N_42061,N_37515,N_38350);
or U42062 (N_42062,N_37837,N_37799);
nor U42063 (N_42063,N_39628,N_39689);
xor U42064 (N_42064,N_38962,N_38292);
or U42065 (N_42065,N_37741,N_38939);
xor U42066 (N_42066,N_38278,N_39137);
and U42067 (N_42067,N_38321,N_39784);
xor U42068 (N_42068,N_38895,N_38523);
nand U42069 (N_42069,N_37508,N_39487);
or U42070 (N_42070,N_39002,N_37515);
xor U42071 (N_42071,N_38851,N_37767);
nand U42072 (N_42072,N_39177,N_38275);
nand U42073 (N_42073,N_39453,N_38500);
nor U42074 (N_42074,N_37620,N_39243);
nor U42075 (N_42075,N_38170,N_39171);
or U42076 (N_42076,N_38567,N_39214);
and U42077 (N_42077,N_37581,N_38979);
or U42078 (N_42078,N_39984,N_39181);
xnor U42079 (N_42079,N_39565,N_37781);
or U42080 (N_42080,N_39978,N_37819);
and U42081 (N_42081,N_37599,N_39847);
or U42082 (N_42082,N_37714,N_37911);
xnor U42083 (N_42083,N_38897,N_39052);
nand U42084 (N_42084,N_37814,N_39453);
xnor U42085 (N_42085,N_37607,N_38188);
xnor U42086 (N_42086,N_39304,N_37699);
or U42087 (N_42087,N_38293,N_39708);
and U42088 (N_42088,N_39973,N_39584);
or U42089 (N_42089,N_39906,N_37510);
nor U42090 (N_42090,N_38931,N_37861);
xor U42091 (N_42091,N_37530,N_38753);
nor U42092 (N_42092,N_38792,N_39819);
nand U42093 (N_42093,N_38609,N_39335);
nand U42094 (N_42094,N_39644,N_38291);
and U42095 (N_42095,N_38150,N_38627);
nand U42096 (N_42096,N_38504,N_39573);
or U42097 (N_42097,N_38957,N_38026);
and U42098 (N_42098,N_38309,N_39235);
xnor U42099 (N_42099,N_38389,N_38554);
or U42100 (N_42100,N_37984,N_39787);
nand U42101 (N_42101,N_38911,N_37981);
nor U42102 (N_42102,N_39241,N_37611);
or U42103 (N_42103,N_38210,N_37531);
nand U42104 (N_42104,N_38736,N_39614);
or U42105 (N_42105,N_39891,N_37572);
nor U42106 (N_42106,N_38817,N_39049);
nor U42107 (N_42107,N_38518,N_39632);
or U42108 (N_42108,N_38942,N_38909);
nand U42109 (N_42109,N_38872,N_39092);
xnor U42110 (N_42110,N_38259,N_39842);
nand U42111 (N_42111,N_38288,N_39751);
nor U42112 (N_42112,N_37795,N_38414);
xnor U42113 (N_42113,N_37896,N_39610);
or U42114 (N_42114,N_38316,N_38964);
or U42115 (N_42115,N_37670,N_38704);
or U42116 (N_42116,N_39044,N_38608);
nor U42117 (N_42117,N_37542,N_38202);
or U42118 (N_42118,N_38590,N_39438);
and U42119 (N_42119,N_39312,N_37655);
and U42120 (N_42120,N_38710,N_39795);
nand U42121 (N_42121,N_38867,N_38280);
or U42122 (N_42122,N_39578,N_37755);
xor U42123 (N_42123,N_38632,N_37862);
and U42124 (N_42124,N_38785,N_39808);
nor U42125 (N_42125,N_39895,N_37840);
xnor U42126 (N_42126,N_39325,N_39668);
xor U42127 (N_42127,N_38720,N_39607);
and U42128 (N_42128,N_38170,N_39953);
nand U42129 (N_42129,N_38382,N_38392);
nor U42130 (N_42130,N_39578,N_39713);
xnor U42131 (N_42131,N_37720,N_39770);
or U42132 (N_42132,N_38929,N_38637);
nand U42133 (N_42133,N_38724,N_37562);
nor U42134 (N_42134,N_39217,N_39873);
nor U42135 (N_42135,N_39033,N_38181);
nand U42136 (N_42136,N_39858,N_38413);
nor U42137 (N_42137,N_37898,N_39706);
nor U42138 (N_42138,N_37841,N_39680);
xnor U42139 (N_42139,N_38968,N_38102);
nand U42140 (N_42140,N_39861,N_38130);
or U42141 (N_42141,N_38842,N_39334);
or U42142 (N_42142,N_38953,N_38885);
nor U42143 (N_42143,N_39397,N_39122);
nand U42144 (N_42144,N_38411,N_39285);
nor U42145 (N_42145,N_38968,N_37676);
nand U42146 (N_42146,N_37768,N_39562);
xor U42147 (N_42147,N_37853,N_37995);
nand U42148 (N_42148,N_38043,N_38601);
nand U42149 (N_42149,N_39712,N_38517);
nor U42150 (N_42150,N_39575,N_37921);
nor U42151 (N_42151,N_38638,N_38803);
nand U42152 (N_42152,N_39440,N_38504);
nand U42153 (N_42153,N_39530,N_37600);
nor U42154 (N_42154,N_38571,N_37535);
nor U42155 (N_42155,N_38291,N_39411);
nor U42156 (N_42156,N_39099,N_38824);
xor U42157 (N_42157,N_38882,N_38198);
or U42158 (N_42158,N_38276,N_37812);
and U42159 (N_42159,N_39290,N_39705);
and U42160 (N_42160,N_39253,N_39146);
xor U42161 (N_42161,N_38627,N_38426);
nor U42162 (N_42162,N_38783,N_37956);
or U42163 (N_42163,N_39219,N_38259);
or U42164 (N_42164,N_38566,N_38792);
nand U42165 (N_42165,N_38716,N_39699);
and U42166 (N_42166,N_37736,N_39572);
or U42167 (N_42167,N_39176,N_37813);
and U42168 (N_42168,N_38963,N_38414);
and U42169 (N_42169,N_39412,N_39607);
nor U42170 (N_42170,N_39558,N_38415);
and U42171 (N_42171,N_37896,N_38330);
and U42172 (N_42172,N_38132,N_38082);
nor U42173 (N_42173,N_39974,N_39057);
and U42174 (N_42174,N_39907,N_38407);
nor U42175 (N_42175,N_39167,N_39651);
nor U42176 (N_42176,N_38195,N_37677);
nand U42177 (N_42177,N_38853,N_39282);
and U42178 (N_42178,N_38780,N_39049);
nor U42179 (N_42179,N_39136,N_39959);
or U42180 (N_42180,N_37905,N_37584);
or U42181 (N_42181,N_38414,N_38757);
nor U42182 (N_42182,N_38945,N_38527);
or U42183 (N_42183,N_38546,N_39836);
nand U42184 (N_42184,N_37602,N_38389);
or U42185 (N_42185,N_39121,N_39875);
xnor U42186 (N_42186,N_39324,N_38001);
or U42187 (N_42187,N_37648,N_37581);
and U42188 (N_42188,N_37952,N_39510);
nor U42189 (N_42189,N_39305,N_39294);
xnor U42190 (N_42190,N_37666,N_39050);
or U42191 (N_42191,N_39500,N_38900);
or U42192 (N_42192,N_38028,N_38784);
or U42193 (N_42193,N_39867,N_39573);
nand U42194 (N_42194,N_39656,N_37991);
and U42195 (N_42195,N_39881,N_38487);
and U42196 (N_42196,N_37792,N_38461);
nand U42197 (N_42197,N_37556,N_37824);
xnor U42198 (N_42198,N_39706,N_37647);
or U42199 (N_42199,N_37529,N_37830);
xor U42200 (N_42200,N_38840,N_38654);
nand U42201 (N_42201,N_37637,N_38903);
nor U42202 (N_42202,N_38383,N_39175);
xor U42203 (N_42203,N_38324,N_38865);
nand U42204 (N_42204,N_38020,N_38755);
nor U42205 (N_42205,N_39453,N_38840);
or U42206 (N_42206,N_39347,N_39694);
nand U42207 (N_42207,N_38769,N_39664);
nor U42208 (N_42208,N_38226,N_38989);
or U42209 (N_42209,N_37965,N_38695);
and U42210 (N_42210,N_39781,N_39580);
or U42211 (N_42211,N_37557,N_37724);
nand U42212 (N_42212,N_38314,N_39277);
nor U42213 (N_42213,N_39800,N_39779);
or U42214 (N_42214,N_39989,N_37565);
or U42215 (N_42215,N_39597,N_37985);
or U42216 (N_42216,N_38823,N_39967);
nor U42217 (N_42217,N_37547,N_39572);
or U42218 (N_42218,N_38184,N_39114);
xnor U42219 (N_42219,N_38382,N_39599);
xor U42220 (N_42220,N_39160,N_39935);
nand U42221 (N_42221,N_39322,N_39387);
and U42222 (N_42222,N_39249,N_39059);
nor U42223 (N_42223,N_38237,N_39489);
nand U42224 (N_42224,N_37790,N_38982);
or U42225 (N_42225,N_37702,N_39731);
nor U42226 (N_42226,N_37823,N_39073);
and U42227 (N_42227,N_39020,N_38254);
xor U42228 (N_42228,N_38725,N_37770);
nor U42229 (N_42229,N_39559,N_38106);
and U42230 (N_42230,N_38125,N_37722);
nor U42231 (N_42231,N_39330,N_38480);
xnor U42232 (N_42232,N_39016,N_39202);
and U42233 (N_42233,N_37727,N_38077);
or U42234 (N_42234,N_38651,N_39061);
and U42235 (N_42235,N_38753,N_37761);
nor U42236 (N_42236,N_37703,N_38282);
nor U42237 (N_42237,N_38261,N_39256);
nand U42238 (N_42238,N_39339,N_38228);
nor U42239 (N_42239,N_38177,N_38980);
or U42240 (N_42240,N_38681,N_38831);
nor U42241 (N_42241,N_39155,N_38329);
and U42242 (N_42242,N_38706,N_39749);
nor U42243 (N_42243,N_38260,N_38805);
or U42244 (N_42244,N_38716,N_37500);
nand U42245 (N_42245,N_38917,N_38165);
nor U42246 (N_42246,N_37708,N_39428);
or U42247 (N_42247,N_37883,N_38560);
nand U42248 (N_42248,N_37935,N_39129);
or U42249 (N_42249,N_38999,N_38578);
nor U42250 (N_42250,N_38624,N_37655);
or U42251 (N_42251,N_39183,N_39994);
nor U42252 (N_42252,N_39644,N_38898);
nor U42253 (N_42253,N_39192,N_38169);
nor U42254 (N_42254,N_39488,N_38281);
xor U42255 (N_42255,N_38381,N_39797);
xnor U42256 (N_42256,N_38506,N_39915);
nand U42257 (N_42257,N_37557,N_38531);
nor U42258 (N_42258,N_37687,N_38581);
nor U42259 (N_42259,N_38362,N_38958);
nor U42260 (N_42260,N_38997,N_39211);
and U42261 (N_42261,N_38093,N_38982);
and U42262 (N_42262,N_38886,N_37980);
xor U42263 (N_42263,N_38764,N_37888);
nor U42264 (N_42264,N_37504,N_39867);
xnor U42265 (N_42265,N_39131,N_38674);
nand U42266 (N_42266,N_38806,N_39426);
and U42267 (N_42267,N_37939,N_38366);
and U42268 (N_42268,N_38293,N_38969);
nor U42269 (N_42269,N_37787,N_38460);
nor U42270 (N_42270,N_38685,N_39316);
nand U42271 (N_42271,N_38071,N_39695);
nor U42272 (N_42272,N_37687,N_38356);
xnor U42273 (N_42273,N_37842,N_38758);
or U42274 (N_42274,N_38261,N_39745);
and U42275 (N_42275,N_38221,N_37677);
or U42276 (N_42276,N_38469,N_38025);
nand U42277 (N_42277,N_39328,N_39911);
or U42278 (N_42278,N_37766,N_37752);
and U42279 (N_42279,N_39168,N_39941);
xor U42280 (N_42280,N_39651,N_38558);
or U42281 (N_42281,N_39446,N_39375);
or U42282 (N_42282,N_38888,N_38320);
nor U42283 (N_42283,N_39804,N_38448);
or U42284 (N_42284,N_39737,N_39364);
and U42285 (N_42285,N_38952,N_38164);
nand U42286 (N_42286,N_39172,N_39360);
xor U42287 (N_42287,N_38944,N_38455);
nor U42288 (N_42288,N_38140,N_37574);
nor U42289 (N_42289,N_39341,N_37690);
xor U42290 (N_42290,N_38820,N_37948);
and U42291 (N_42291,N_38660,N_38844);
xnor U42292 (N_42292,N_39255,N_39583);
or U42293 (N_42293,N_38089,N_39102);
xor U42294 (N_42294,N_37514,N_38581);
xor U42295 (N_42295,N_39771,N_37518);
or U42296 (N_42296,N_39299,N_38326);
and U42297 (N_42297,N_39938,N_37735);
nand U42298 (N_42298,N_38300,N_39229);
and U42299 (N_42299,N_37642,N_38438);
and U42300 (N_42300,N_39943,N_39739);
xor U42301 (N_42301,N_38304,N_37916);
and U42302 (N_42302,N_38632,N_38394);
nor U42303 (N_42303,N_39031,N_37597);
nand U42304 (N_42304,N_38232,N_37924);
or U42305 (N_42305,N_37791,N_39587);
and U42306 (N_42306,N_38878,N_38723);
nand U42307 (N_42307,N_37726,N_39088);
nor U42308 (N_42308,N_38415,N_38662);
nand U42309 (N_42309,N_39725,N_39438);
and U42310 (N_42310,N_37779,N_39954);
or U42311 (N_42311,N_37684,N_38079);
nand U42312 (N_42312,N_37658,N_38039);
nand U42313 (N_42313,N_39702,N_39186);
or U42314 (N_42314,N_39143,N_38429);
or U42315 (N_42315,N_38502,N_39786);
or U42316 (N_42316,N_39649,N_38088);
and U42317 (N_42317,N_37660,N_38449);
or U42318 (N_42318,N_39676,N_37990);
nand U42319 (N_42319,N_39301,N_37603);
nand U42320 (N_42320,N_37743,N_38063);
nand U42321 (N_42321,N_38131,N_38834);
xnor U42322 (N_42322,N_39474,N_38581);
nor U42323 (N_42323,N_38058,N_38961);
and U42324 (N_42324,N_38448,N_39856);
and U42325 (N_42325,N_38664,N_39458);
xnor U42326 (N_42326,N_39889,N_38210);
and U42327 (N_42327,N_37694,N_38079);
or U42328 (N_42328,N_39881,N_37770);
xor U42329 (N_42329,N_39868,N_39192);
xnor U42330 (N_42330,N_39521,N_38980);
nor U42331 (N_42331,N_37900,N_39726);
or U42332 (N_42332,N_37641,N_37691);
and U42333 (N_42333,N_39546,N_38079);
and U42334 (N_42334,N_39489,N_38640);
xor U42335 (N_42335,N_37756,N_38530);
nand U42336 (N_42336,N_39585,N_38827);
xnor U42337 (N_42337,N_37977,N_39491);
nor U42338 (N_42338,N_37951,N_38164);
or U42339 (N_42339,N_39880,N_39569);
and U42340 (N_42340,N_39786,N_37891);
xor U42341 (N_42341,N_39387,N_38233);
and U42342 (N_42342,N_38263,N_38971);
nor U42343 (N_42343,N_37898,N_37921);
nor U42344 (N_42344,N_39418,N_38638);
and U42345 (N_42345,N_39659,N_38846);
xnor U42346 (N_42346,N_38333,N_38771);
xnor U42347 (N_42347,N_39146,N_39313);
and U42348 (N_42348,N_39141,N_38364);
nor U42349 (N_42349,N_38869,N_38409);
or U42350 (N_42350,N_38660,N_37691);
nor U42351 (N_42351,N_37965,N_38963);
nor U42352 (N_42352,N_39986,N_39078);
nand U42353 (N_42353,N_39245,N_38640);
nor U42354 (N_42354,N_39050,N_38070);
nand U42355 (N_42355,N_39046,N_39973);
or U42356 (N_42356,N_37855,N_38597);
nor U42357 (N_42357,N_37857,N_38007);
and U42358 (N_42358,N_39859,N_37990);
or U42359 (N_42359,N_37778,N_37946);
nor U42360 (N_42360,N_37981,N_38865);
nor U42361 (N_42361,N_38151,N_38576);
or U42362 (N_42362,N_38135,N_39145);
nor U42363 (N_42363,N_37832,N_38443);
and U42364 (N_42364,N_38930,N_39431);
nand U42365 (N_42365,N_37945,N_39027);
or U42366 (N_42366,N_38791,N_39829);
and U42367 (N_42367,N_39866,N_39341);
xor U42368 (N_42368,N_39184,N_39661);
xnor U42369 (N_42369,N_39416,N_39910);
xor U42370 (N_42370,N_38788,N_38391);
nor U42371 (N_42371,N_37696,N_39444);
or U42372 (N_42372,N_39231,N_37517);
nand U42373 (N_42373,N_38252,N_38497);
nand U42374 (N_42374,N_37575,N_38306);
and U42375 (N_42375,N_38575,N_37919);
or U42376 (N_42376,N_38474,N_37906);
or U42377 (N_42377,N_38699,N_37783);
and U42378 (N_42378,N_38540,N_39654);
or U42379 (N_42379,N_38094,N_39483);
nand U42380 (N_42380,N_38149,N_38778);
and U42381 (N_42381,N_39556,N_37922);
nand U42382 (N_42382,N_39417,N_38749);
nor U42383 (N_42383,N_38533,N_38685);
nand U42384 (N_42384,N_37705,N_39358);
and U42385 (N_42385,N_39337,N_39886);
and U42386 (N_42386,N_38664,N_37507);
nor U42387 (N_42387,N_39056,N_38729);
xnor U42388 (N_42388,N_39885,N_37770);
and U42389 (N_42389,N_37511,N_39178);
and U42390 (N_42390,N_37782,N_38103);
nor U42391 (N_42391,N_38191,N_39886);
and U42392 (N_42392,N_39827,N_39414);
or U42393 (N_42393,N_38437,N_39544);
xnor U42394 (N_42394,N_37841,N_38791);
xnor U42395 (N_42395,N_39195,N_38639);
or U42396 (N_42396,N_37880,N_39651);
and U42397 (N_42397,N_38774,N_38595);
xnor U42398 (N_42398,N_38774,N_39081);
nand U42399 (N_42399,N_38002,N_39842);
nand U42400 (N_42400,N_39684,N_39685);
or U42401 (N_42401,N_38676,N_39925);
xor U42402 (N_42402,N_38201,N_38791);
nand U42403 (N_42403,N_38131,N_39626);
xnor U42404 (N_42404,N_37919,N_38969);
and U42405 (N_42405,N_38299,N_39254);
or U42406 (N_42406,N_38186,N_37774);
nor U42407 (N_42407,N_37719,N_38478);
xnor U42408 (N_42408,N_39200,N_37854);
xnor U42409 (N_42409,N_38496,N_37621);
nand U42410 (N_42410,N_39829,N_39925);
xor U42411 (N_42411,N_37860,N_38139);
and U42412 (N_42412,N_39877,N_39958);
nand U42413 (N_42413,N_37998,N_38226);
nor U42414 (N_42414,N_38495,N_37510);
and U42415 (N_42415,N_38569,N_39790);
nand U42416 (N_42416,N_39519,N_38468);
nor U42417 (N_42417,N_39869,N_37572);
nand U42418 (N_42418,N_39478,N_38378);
nor U42419 (N_42419,N_38164,N_38775);
nand U42420 (N_42420,N_38788,N_38222);
nor U42421 (N_42421,N_38365,N_38345);
nand U42422 (N_42422,N_38329,N_39786);
or U42423 (N_42423,N_39235,N_38206);
or U42424 (N_42424,N_39147,N_38499);
and U42425 (N_42425,N_38017,N_38212);
xnor U42426 (N_42426,N_39101,N_37942);
or U42427 (N_42427,N_38393,N_39270);
nor U42428 (N_42428,N_39244,N_39066);
xnor U42429 (N_42429,N_39810,N_37922);
and U42430 (N_42430,N_39651,N_39450);
and U42431 (N_42431,N_38843,N_39657);
or U42432 (N_42432,N_39518,N_39457);
nand U42433 (N_42433,N_38638,N_37770);
or U42434 (N_42434,N_38531,N_39518);
or U42435 (N_42435,N_38582,N_38897);
nor U42436 (N_42436,N_38955,N_39491);
and U42437 (N_42437,N_38111,N_38767);
and U42438 (N_42438,N_38952,N_38269);
xor U42439 (N_42439,N_38562,N_37609);
nor U42440 (N_42440,N_39955,N_37729);
xnor U42441 (N_42441,N_37535,N_38127);
xor U42442 (N_42442,N_39242,N_38277);
nand U42443 (N_42443,N_39350,N_37557);
or U42444 (N_42444,N_39172,N_39901);
and U42445 (N_42445,N_38078,N_39002);
or U42446 (N_42446,N_38494,N_39362);
nor U42447 (N_42447,N_38918,N_37992);
or U42448 (N_42448,N_39408,N_37806);
nand U42449 (N_42449,N_37840,N_39809);
nand U42450 (N_42450,N_39608,N_38929);
nand U42451 (N_42451,N_38293,N_39965);
xor U42452 (N_42452,N_39562,N_37891);
and U42453 (N_42453,N_38659,N_39132);
nor U42454 (N_42454,N_39168,N_38989);
and U42455 (N_42455,N_38601,N_38784);
nor U42456 (N_42456,N_38728,N_38193);
nand U42457 (N_42457,N_39012,N_38937);
or U42458 (N_42458,N_38501,N_38395);
and U42459 (N_42459,N_37792,N_38826);
nor U42460 (N_42460,N_38963,N_39324);
and U42461 (N_42461,N_39990,N_38133);
and U42462 (N_42462,N_39111,N_38301);
xor U42463 (N_42463,N_38940,N_37702);
nor U42464 (N_42464,N_39909,N_39703);
and U42465 (N_42465,N_37628,N_38521);
nor U42466 (N_42466,N_37851,N_39027);
and U42467 (N_42467,N_39496,N_39991);
nand U42468 (N_42468,N_39930,N_38096);
nand U42469 (N_42469,N_37577,N_37871);
xor U42470 (N_42470,N_37567,N_38296);
xnor U42471 (N_42471,N_38182,N_38300);
and U42472 (N_42472,N_38383,N_38517);
nor U42473 (N_42473,N_37602,N_37865);
and U42474 (N_42474,N_39873,N_39602);
xnor U42475 (N_42475,N_39053,N_39558);
and U42476 (N_42476,N_38036,N_38929);
nand U42477 (N_42477,N_38957,N_39138);
and U42478 (N_42478,N_37959,N_38634);
nor U42479 (N_42479,N_38349,N_38715);
or U42480 (N_42480,N_39691,N_39743);
and U42481 (N_42481,N_39724,N_37770);
nand U42482 (N_42482,N_37559,N_39397);
nand U42483 (N_42483,N_38382,N_39813);
nor U42484 (N_42484,N_38597,N_37562);
and U42485 (N_42485,N_39743,N_39450);
and U42486 (N_42486,N_37785,N_38240);
xnor U42487 (N_42487,N_37629,N_38907);
nor U42488 (N_42488,N_37803,N_38623);
nor U42489 (N_42489,N_39351,N_39415);
or U42490 (N_42490,N_38448,N_37668);
nand U42491 (N_42491,N_39810,N_37652);
and U42492 (N_42492,N_39868,N_37889);
xor U42493 (N_42493,N_37936,N_39316);
nor U42494 (N_42494,N_39620,N_38084);
nor U42495 (N_42495,N_38104,N_39737);
nand U42496 (N_42496,N_38639,N_38549);
xor U42497 (N_42497,N_37541,N_39303);
xor U42498 (N_42498,N_39630,N_38872);
or U42499 (N_42499,N_38745,N_38047);
nor U42500 (N_42500,N_40221,N_41293);
or U42501 (N_42501,N_40952,N_42250);
or U42502 (N_42502,N_40726,N_41365);
nor U42503 (N_42503,N_41639,N_42066);
and U42504 (N_42504,N_40733,N_41677);
or U42505 (N_42505,N_42186,N_42056);
nand U42506 (N_42506,N_40302,N_40004);
or U42507 (N_42507,N_41885,N_42285);
and U42508 (N_42508,N_42165,N_40755);
xnor U42509 (N_42509,N_41851,N_41589);
xnor U42510 (N_42510,N_40363,N_40604);
or U42511 (N_42511,N_42380,N_40329);
and U42512 (N_42512,N_42488,N_40529);
and U42513 (N_42513,N_42118,N_41600);
nor U42514 (N_42514,N_42399,N_42005);
nor U42515 (N_42515,N_41936,N_40440);
nand U42516 (N_42516,N_40069,N_40662);
nand U42517 (N_42517,N_40047,N_40818);
or U42518 (N_42518,N_41286,N_41194);
and U42519 (N_42519,N_42304,N_42158);
nor U42520 (N_42520,N_40960,N_41372);
nor U42521 (N_42521,N_42443,N_42340);
nor U42522 (N_42522,N_41797,N_40067);
and U42523 (N_42523,N_40371,N_42463);
nand U42524 (N_42524,N_42050,N_40621);
xnor U42525 (N_42525,N_40553,N_41596);
nor U42526 (N_42526,N_41711,N_40867);
nand U42527 (N_42527,N_40948,N_40296);
nand U42528 (N_42528,N_40574,N_40417);
or U42529 (N_42529,N_40066,N_40128);
and U42530 (N_42530,N_41395,N_40305);
or U42531 (N_42531,N_42052,N_41346);
nor U42532 (N_42532,N_41350,N_40289);
xor U42533 (N_42533,N_40978,N_41064);
xnor U42534 (N_42534,N_40690,N_41424);
and U42535 (N_42535,N_41602,N_41321);
and U42536 (N_42536,N_41919,N_41918);
nor U42537 (N_42537,N_42174,N_41545);
nand U42538 (N_42538,N_42494,N_42491);
nand U42539 (N_42539,N_42498,N_41567);
and U42540 (N_42540,N_42205,N_40197);
or U42541 (N_42541,N_40573,N_41893);
nand U42542 (N_42542,N_42135,N_40859);
nand U42543 (N_42543,N_42177,N_40123);
xnor U42544 (N_42544,N_42375,N_41869);
nor U42545 (N_42545,N_42295,N_42263);
nand U42546 (N_42546,N_41714,N_41543);
xor U42547 (N_42547,N_41276,N_41608);
nand U42548 (N_42548,N_41171,N_42041);
nand U42549 (N_42549,N_42253,N_40708);
or U42550 (N_42550,N_40936,N_42449);
and U42551 (N_42551,N_41322,N_42356);
and U42552 (N_42552,N_40452,N_40073);
nand U42553 (N_42553,N_41694,N_42040);
or U42554 (N_42554,N_41040,N_40202);
and U42555 (N_42555,N_40348,N_41298);
nand U42556 (N_42556,N_41411,N_40741);
and U42557 (N_42557,N_41094,N_42201);
nand U42558 (N_42558,N_42029,N_41777);
or U42559 (N_42559,N_41361,N_40837);
nor U42560 (N_42560,N_41642,N_42436);
xor U42561 (N_42561,N_40385,N_40209);
and U42562 (N_42562,N_42492,N_41228);
xor U42563 (N_42563,N_40965,N_41509);
nor U42564 (N_42564,N_41930,N_41086);
or U42565 (N_42565,N_41713,N_40118);
nand U42566 (N_42566,N_41865,N_40366);
nand U42567 (N_42567,N_41904,N_41133);
or U42568 (N_42568,N_41952,N_42230);
and U42569 (N_42569,N_42388,N_41613);
or U42570 (N_42570,N_41947,N_41754);
xor U42571 (N_42571,N_41128,N_40617);
nor U42572 (N_42572,N_40001,N_40571);
and U42573 (N_42573,N_40792,N_42339);
and U42574 (N_42574,N_40855,N_40035);
or U42575 (N_42575,N_41609,N_42358);
nand U42576 (N_42576,N_42487,N_42318);
and U42577 (N_42577,N_41465,N_40187);
and U42578 (N_42578,N_42298,N_41561);
or U42579 (N_42579,N_41867,N_40083);
nand U42580 (N_42580,N_41884,N_41192);
nor U42581 (N_42581,N_40985,N_40191);
and U42582 (N_42582,N_42261,N_41778);
xnor U42583 (N_42583,N_41481,N_41989);
nand U42584 (N_42584,N_42167,N_41646);
and U42585 (N_42585,N_42422,N_41689);
nand U42586 (N_42586,N_42014,N_42310);
nand U42587 (N_42587,N_42244,N_40237);
and U42588 (N_42588,N_40585,N_42353);
and U42589 (N_42589,N_40567,N_42107);
and U42590 (N_42590,N_41747,N_42035);
and U42591 (N_42591,N_41480,N_42227);
nand U42592 (N_42592,N_41901,N_40849);
nor U42593 (N_42593,N_40184,N_42199);
nand U42594 (N_42594,N_40010,N_40620);
nand U42595 (N_42595,N_41297,N_41837);
and U42596 (N_42596,N_42495,N_41807);
xor U42597 (N_42597,N_40103,N_42370);
nor U42598 (N_42598,N_40122,N_42018);
or U42599 (N_42599,N_40929,N_41095);
or U42600 (N_42600,N_41647,N_40771);
or U42601 (N_42601,N_41164,N_41109);
and U42602 (N_42602,N_40909,N_41058);
nand U42603 (N_42603,N_42299,N_40497);
and U42604 (N_42604,N_41287,N_41848);
and U42605 (N_42605,N_40145,N_41102);
nand U42606 (N_42606,N_40940,N_40603);
nand U42607 (N_42607,N_40976,N_41091);
xnor U42608 (N_42608,N_41431,N_40860);
and U42609 (N_42609,N_41097,N_41858);
and U42610 (N_42610,N_40381,N_40406);
and U42611 (N_42611,N_41539,N_42249);
and U42612 (N_42612,N_40404,N_40809);
nor U42613 (N_42613,N_40101,N_41055);
or U42614 (N_42614,N_40132,N_40286);
xor U42615 (N_42615,N_41850,N_40919);
nand U42616 (N_42616,N_40674,N_41116);
nand U42617 (N_42617,N_42479,N_40565);
xnor U42618 (N_42618,N_40508,N_40133);
and U42619 (N_42619,N_42334,N_41566);
and U42620 (N_42620,N_42081,N_42101);
and U42621 (N_42621,N_40550,N_40559);
nand U42622 (N_42622,N_40706,N_42307);
nor U42623 (N_42623,N_42475,N_41572);
xnor U42624 (N_42624,N_40899,N_41935);
and U42625 (N_42625,N_42465,N_41290);
nor U42626 (N_42626,N_42140,N_42028);
and U42627 (N_42627,N_41436,N_42176);
and U42628 (N_42628,N_41767,N_42218);
nor U42629 (N_42629,N_42444,N_41643);
or U42630 (N_42630,N_41597,N_40071);
nand U42631 (N_42631,N_41635,N_42226);
nor U42632 (N_42632,N_42308,N_40825);
xnor U42633 (N_42633,N_40683,N_40661);
and U42634 (N_42634,N_40396,N_42473);
nand U42635 (N_42635,N_41351,N_41854);
nand U42636 (N_42636,N_41698,N_40161);
xnor U42637 (N_42637,N_41186,N_41426);
or U42638 (N_42638,N_41299,N_42352);
nand U42639 (N_42639,N_41945,N_41666);
and U42640 (N_42640,N_41588,N_40325);
xor U42641 (N_42641,N_41779,N_41631);
or U42642 (N_42642,N_40479,N_41209);
and U42643 (N_42643,N_41576,N_41143);
and U42644 (N_42644,N_41551,N_41515);
nand U42645 (N_42645,N_42207,N_41033);
nor U42646 (N_42646,N_40776,N_41997);
or U42647 (N_42647,N_42054,N_40331);
nor U42648 (N_42648,N_41521,N_41004);
xor U42649 (N_42649,N_42431,N_40634);
nand U42650 (N_42650,N_40074,N_41870);
nand U42651 (N_42651,N_41934,N_40689);
or U42652 (N_42652,N_41111,N_40306);
and U42653 (N_42653,N_40866,N_41861);
xor U42654 (N_42654,N_42031,N_41003);
nor U42655 (N_42655,N_42115,N_40596);
nor U42656 (N_42656,N_41818,N_41451);
nand U42657 (N_42657,N_40893,N_40100);
nand U42658 (N_42658,N_40090,N_41816);
nor U42659 (N_42659,N_40416,N_40050);
nand U42660 (N_42660,N_40138,N_40005);
xor U42661 (N_42661,N_40283,N_40079);
nor U42662 (N_42662,N_40271,N_40579);
xnor U42663 (N_42663,N_41274,N_40534);
nand U42664 (N_42664,N_42113,N_41054);
xor U42665 (N_42665,N_40525,N_41916);
nand U42666 (N_42666,N_40974,N_40872);
nor U42667 (N_42667,N_40458,N_41970);
and U42668 (N_42668,N_40545,N_40943);
nand U42669 (N_42669,N_41288,N_40135);
or U42670 (N_42670,N_41814,N_41531);
or U42671 (N_42671,N_42132,N_41881);
nand U42672 (N_42672,N_41099,N_40429);
or U42673 (N_42673,N_40979,N_40334);
xor U42674 (N_42674,N_42030,N_42407);
xor U42675 (N_42675,N_40758,N_40397);
nor U42676 (N_42676,N_40147,N_42151);
and U42677 (N_42677,N_41429,N_41633);
nor U42678 (N_42678,N_40433,N_41319);
nand U42679 (N_42679,N_41315,N_41190);
nand U42680 (N_42680,N_42195,N_40402);
or U42681 (N_42681,N_41991,N_41206);
nand U42682 (N_42682,N_41441,N_40017);
xnor U42683 (N_42683,N_41360,N_42163);
or U42684 (N_42684,N_40436,N_41199);
nor U42685 (N_42685,N_42364,N_41354);
or U42686 (N_42686,N_40229,N_40712);
xnor U42687 (N_42687,N_41400,N_42266);
xnor U42688 (N_42688,N_40319,N_40554);
and U42689 (N_42689,N_42361,N_40388);
xnor U42690 (N_42690,N_42457,N_40225);
nand U42691 (N_42691,N_40057,N_41506);
nand U42692 (N_42692,N_42435,N_41502);
or U42693 (N_42693,N_41528,N_40810);
xor U42694 (N_42694,N_40645,N_41047);
and U42695 (N_42695,N_42341,N_42319);
or U42696 (N_42696,N_41002,N_41808);
and U42697 (N_42697,N_40218,N_42231);
xor U42698 (N_42698,N_40852,N_41674);
nand U42699 (N_42699,N_40387,N_40806);
xor U42700 (N_42700,N_41306,N_41087);
nand U42701 (N_42701,N_41239,N_40790);
nand U42702 (N_42702,N_40422,N_41084);
nand U42703 (N_42703,N_40921,N_42190);
or U42704 (N_42704,N_41333,N_41131);
nand U42705 (N_42705,N_41150,N_40315);
nor U42706 (N_42706,N_41847,N_40993);
nor U42707 (N_42707,N_40703,N_42099);
or U42708 (N_42708,N_40829,N_40013);
and U42709 (N_42709,N_40793,N_41686);
or U42710 (N_42710,N_40091,N_42419);
nor U42711 (N_42711,N_40130,N_42223);
nand U42712 (N_42712,N_40292,N_40544);
nand U42713 (N_42713,N_41129,N_41487);
nand U42714 (N_42714,N_41096,N_40097);
nor U42715 (N_42715,N_40176,N_40226);
and U42716 (N_42716,N_42168,N_41179);
nor U42717 (N_42717,N_42093,N_41340);
or U42718 (N_42718,N_41446,N_41103);
nand U42719 (N_42719,N_41706,N_42063);
or U42720 (N_42720,N_40380,N_40214);
and U42721 (N_42721,N_41175,N_40833);
nand U42722 (N_42722,N_40231,N_41390);
and U42723 (N_42723,N_40140,N_41853);
xnor U42724 (N_42724,N_40156,N_40175);
xor U42725 (N_42725,N_40316,N_40768);
xnor U42726 (N_42726,N_41962,N_40420);
nor U42727 (N_42727,N_41247,N_40854);
nand U42728 (N_42728,N_41599,N_41914);
xor U42729 (N_42729,N_41628,N_40558);
xnor U42730 (N_42730,N_41012,N_40610);
nand U42731 (N_42731,N_42453,N_41264);
xnor U42732 (N_42732,N_42126,N_41999);
or U42733 (N_42733,N_42330,N_41938);
and U42734 (N_42734,N_41015,N_40524);
or U42735 (N_42735,N_41011,N_41637);
xor U42736 (N_42736,N_40456,N_40644);
nor U42737 (N_42737,N_40947,N_41627);
xor U42738 (N_42738,N_40281,N_41430);
xor U42739 (N_42739,N_41972,N_40379);
xnor U42740 (N_42740,N_41392,N_41349);
and U42741 (N_42741,N_40643,N_42350);
or U42742 (N_42742,N_41219,N_40483);
and U42743 (N_42743,N_40280,N_41137);
nand U42744 (N_42744,N_41156,N_41690);
nand U42745 (N_42745,N_40834,N_40982);
or U42746 (N_42746,N_42239,N_40763);
and U42747 (N_42747,N_41335,N_42215);
nand U42748 (N_42748,N_40668,N_42152);
nor U42749 (N_42749,N_41908,N_42349);
xnor U42750 (N_42750,N_40206,N_40408);
or U42751 (N_42751,N_40638,N_40764);
nand U42752 (N_42752,N_40046,N_41035);
and U42753 (N_42753,N_42321,N_40355);
xor U42754 (N_42754,N_40200,N_42044);
or U42755 (N_42755,N_42301,N_40041);
xor U42756 (N_42756,N_41231,N_40142);
xnor U42757 (N_42757,N_42009,N_41891);
or U42758 (N_42758,N_41911,N_42104);
nor U42759 (N_42759,N_40054,N_41452);
or U42760 (N_42760,N_42120,N_41728);
nand U42761 (N_42761,N_41760,N_40060);
nor U42762 (N_42762,N_42222,N_42197);
nand U42763 (N_42763,N_40522,N_41636);
xnor U42764 (N_42764,N_41367,N_41699);
nand U42765 (N_42765,N_42480,N_40024);
xor U42766 (N_42766,N_42026,N_41553);
xor U42767 (N_42767,N_41827,N_41542);
nand U42768 (N_42768,N_40357,N_42382);
or U42769 (N_42769,N_40224,N_40770);
nand U42770 (N_42770,N_40616,N_41052);
or U42771 (N_42771,N_40779,N_41326);
xor U42772 (N_42772,N_40914,N_41163);
or U42773 (N_42773,N_42036,N_41325);
nand U42774 (N_42774,N_40595,N_42493);
or U42775 (N_42775,N_41068,N_41594);
and U42776 (N_42776,N_41022,N_42108);
nand U42777 (N_42777,N_41283,N_40879);
or U42778 (N_42778,N_41895,N_40626);
nor U42779 (N_42779,N_40392,N_42280);
and U42780 (N_42780,N_40430,N_42146);
nand U42781 (N_42781,N_41866,N_42306);
and U42782 (N_42782,N_41661,N_41927);
xnor U42783 (N_42783,N_40765,N_40031);
or U42784 (N_42784,N_40875,N_40232);
xor U42785 (N_42785,N_42440,N_42376);
xnor U42786 (N_42786,N_41267,N_40660);
nor U42787 (N_42787,N_41703,N_40169);
or U42788 (N_42788,N_40642,N_40970);
or U42789 (N_42789,N_42450,N_41341);
or U42790 (N_42790,N_40223,N_40518);
xor U42791 (N_42791,N_40020,N_40951);
and U42792 (N_42792,N_42233,N_40814);
xor U42793 (N_42793,N_40501,N_41727);
nand U42794 (N_42794,N_40888,N_41871);
or U42795 (N_42795,N_40513,N_42124);
nand U42796 (N_42796,N_42159,N_40375);
xnor U42797 (N_42797,N_40443,N_42485);
nor U42798 (N_42798,N_42008,N_41044);
and U42799 (N_42799,N_41152,N_40233);
and U42800 (N_42800,N_41393,N_41880);
and U42801 (N_42801,N_40087,N_40519);
xor U42802 (N_42802,N_41549,N_41530);
and U42803 (N_42803,N_40454,N_40516);
or U42804 (N_42804,N_41153,N_41067);
nor U42805 (N_42805,N_42225,N_40160);
nor U42806 (N_42806,N_41582,N_40431);
xor U42807 (N_42807,N_42332,N_42001);
nor U42808 (N_42808,N_40962,N_40382);
nand U42809 (N_42809,N_41332,N_41786);
and U42810 (N_42810,N_40095,N_42342);
nor U42811 (N_42811,N_42481,N_40614);
nor U42812 (N_42812,N_40533,N_40434);
nand U42813 (N_42813,N_41532,N_40900);
nor U42814 (N_42814,N_40998,N_41832);
nor U42815 (N_42815,N_41318,N_40950);
or U42816 (N_42816,N_41799,N_42068);
or U42817 (N_42817,N_40515,N_40905);
nand U42818 (N_42818,N_41277,N_41664);
xor U42819 (N_42819,N_41336,N_41774);
nor U42820 (N_42820,N_40467,N_41391);
xnor U42821 (N_42821,N_40566,N_40590);
or U42822 (N_42822,N_42128,N_40045);
or U42823 (N_42823,N_40125,N_40418);
nand U42824 (N_42824,N_40916,N_42133);
and U42825 (N_42825,N_41181,N_40575);
xor U42826 (N_42826,N_40646,N_40157);
or U42827 (N_42827,N_42461,N_40155);
or U42828 (N_42828,N_41673,N_40500);
or U42829 (N_42829,N_40742,N_42489);
or U42830 (N_42830,N_41776,N_41324);
or U42831 (N_42831,N_40170,N_40030);
nor U42832 (N_42832,N_41556,N_42393);
and U42833 (N_42833,N_42289,N_41188);
nand U42834 (N_42834,N_41671,N_40210);
and U42835 (N_42835,N_41447,N_40372);
nor U42836 (N_42836,N_42271,N_41876);
nor U42837 (N_42837,N_40048,N_42203);
and U42838 (N_42838,N_40485,N_40869);
or U42839 (N_42839,N_40400,N_40795);
and U42840 (N_42840,N_41023,N_41733);
nor U42841 (N_42841,N_41527,N_42499);
or U42842 (N_42842,N_40076,N_42095);
xnor U42843 (N_42843,N_42496,N_42402);
xor U42844 (N_42844,N_42474,N_40230);
xor U42845 (N_42845,N_41598,N_41624);
or U42846 (N_42846,N_40541,N_41289);
nor U42847 (N_42847,N_40273,N_42469);
nand U42848 (N_42848,N_42212,N_40185);
nor U42849 (N_42849,N_41043,N_41427);
nand U42850 (N_42850,N_40736,N_40267);
nor U42851 (N_42851,N_40353,N_40105);
nand U42852 (N_42852,N_40455,N_41301);
nand U42853 (N_42853,N_42413,N_41540);
nand U42854 (N_42854,N_42470,N_41712);
nor U42855 (N_42855,N_41233,N_41444);
xor U42856 (N_42856,N_41682,N_40819);
xor U42857 (N_42857,N_40877,N_41258);
nor U42858 (N_42858,N_41050,N_40242);
or U42859 (N_42859,N_42333,N_40438);
xnor U42860 (N_42860,N_42347,N_40828);
and U42861 (N_42861,N_40126,N_41960);
nor U42862 (N_42862,N_41266,N_40772);
xnor U42863 (N_42863,N_41072,N_40162);
nand U42864 (N_42864,N_41889,N_40492);
nand U42865 (N_42865,N_40012,N_41752);
xor U42866 (N_42866,N_42385,N_42114);
and U42867 (N_42867,N_40631,N_41380);
nor U42868 (N_42868,N_40411,N_41840);
or U42869 (N_42869,N_41462,N_41456);
or U42870 (N_42870,N_42170,N_41507);
nand U42871 (N_42871,N_41535,N_41735);
and U42872 (N_42872,N_40724,N_42416);
nand U42873 (N_42873,N_42377,N_40794);
and U42874 (N_42874,N_42322,N_40865);
nand U42875 (N_42875,N_41825,N_40737);
nor U42876 (N_42876,N_40168,N_41769);
or U42877 (N_42877,N_41486,N_40548);
or U42878 (N_42878,N_40040,N_41353);
xnor U42879 (N_42879,N_41739,N_41701);
and U42880 (N_42880,N_41586,N_40203);
and U42881 (N_42881,N_40992,N_40459);
nand U42882 (N_42882,N_41593,N_41753);
and U42883 (N_42883,N_41039,N_40139);
and U42884 (N_42884,N_42210,N_41987);
nand U42885 (N_42885,N_41591,N_40044);
nor U42886 (N_42886,N_41026,N_42150);
nand U42887 (N_42887,N_41676,N_40798);
or U42888 (N_42888,N_42369,N_40056);
xor U42889 (N_42889,N_41160,N_41142);
nand U42890 (N_42890,N_41278,N_40310);
and U42891 (N_42891,N_40507,N_41449);
or U42892 (N_42892,N_41510,N_42374);
nor U42893 (N_42893,N_40746,N_42346);
nand U42894 (N_42894,N_40775,N_41983);
nor U42895 (N_42895,N_42011,N_40564);
nor U42896 (N_42896,N_40208,N_41155);
nor U42897 (N_42897,N_42395,N_42111);
nor U42898 (N_42898,N_40987,N_40154);
xnor U42899 (N_42899,N_41284,N_40647);
nand U42900 (N_42900,N_41308,N_40466);
nor U42901 (N_42901,N_40425,N_42335);
xor U42902 (N_42902,N_41180,N_40527);
xor U42903 (N_42903,N_41817,N_41826);
and U42904 (N_42904,N_42315,N_40910);
and U42905 (N_42905,N_40370,N_41369);
and U42906 (N_42906,N_40212,N_42178);
xnor U42907 (N_42907,N_41083,N_41491);
nor U42908 (N_42908,N_41442,N_40999);
and U42909 (N_42909,N_40245,N_40088);
and U42910 (N_42910,N_40009,N_40247);
or U42911 (N_42911,N_42238,N_40831);
xor U42912 (N_42912,N_42235,N_41967);
nor U42913 (N_42913,N_42191,N_41580);
nand U42914 (N_42914,N_41811,N_42425);
and U42915 (N_42915,N_40704,N_40696);
and U42916 (N_42916,N_41136,N_41982);
xnor U42917 (N_42917,N_40805,N_40924);
nor U42918 (N_42918,N_41790,N_41018);
nand U42919 (N_42919,N_41587,N_40055);
or U42920 (N_42920,N_42379,N_41839);
or U42921 (N_42921,N_40469,N_40153);
nand U42922 (N_42922,N_40640,N_40716);
or U42923 (N_42923,N_42414,N_40601);
or U42924 (N_42924,N_41119,N_42468);
xnor U42925 (N_42925,N_41906,N_40748);
xnor U42926 (N_42926,N_40848,N_40781);
xor U42927 (N_42927,N_41755,N_41235);
nor U42928 (N_42928,N_40213,N_40262);
nand U42929 (N_42929,N_42070,N_40317);
nand U42930 (N_42930,N_42281,N_40065);
nor U42931 (N_42931,N_41236,N_40086);
nand U42932 (N_42932,N_41124,N_42273);
nand U42933 (N_42933,N_41526,N_41681);
nor U42934 (N_42934,N_40121,N_42433);
or U42935 (N_42935,N_41125,N_40813);
xor U42936 (N_42936,N_41743,N_41725);
nor U42937 (N_42937,N_42466,N_42452);
nand U42938 (N_42938,N_41729,N_41279);
nor U42939 (N_42939,N_41700,N_40751);
nor U42940 (N_42940,N_41595,N_40800);
or U42941 (N_42941,N_41660,N_40415);
and U42942 (N_42942,N_40925,N_41342);
or U42943 (N_42943,N_41285,N_41557);
or U42944 (N_42944,N_42338,N_41915);
nor U42945 (N_42945,N_41494,N_40782);
or U42946 (N_42946,N_40883,N_42325);
xor U42947 (N_42947,N_41806,N_41505);
nand U42948 (N_42948,N_40769,N_40394);
nand U42949 (N_42949,N_41202,N_40785);
or U42950 (N_42950,N_40144,N_40882);
or U42951 (N_42951,N_42360,N_41484);
xor U42952 (N_42952,N_41208,N_41418);
and U42953 (N_42953,N_41630,N_40907);
nor U42954 (N_42954,N_42141,N_40219);
xnor U42955 (N_42955,N_40246,N_40842);
and U42956 (N_42956,N_41872,N_42147);
nand U42957 (N_42957,N_42269,N_40365);
and U42958 (N_42958,N_40783,N_42181);
xor U42959 (N_42959,N_41757,N_41605);
and U42960 (N_42960,N_41078,N_40270);
xnor U42961 (N_42961,N_40826,N_40450);
xnor U42962 (N_42962,N_41210,N_41773);
or U42963 (N_42963,N_41090,N_40444);
and U42964 (N_42964,N_41434,N_40498);
xor U42965 (N_42965,N_42189,N_41857);
nand U42966 (N_42966,N_41417,N_41836);
nand U42967 (N_42967,N_41016,N_41165);
nor U42968 (N_42968,N_42483,N_40847);
and U42969 (N_42969,N_40441,N_41178);
and U42970 (N_42970,N_40390,N_40840);
nand U42971 (N_42971,N_40906,N_40484);
or U42972 (N_42972,N_41842,N_40568);
or U42973 (N_42973,N_41939,N_41080);
xor U42974 (N_42974,N_40652,N_41253);
xnor U42975 (N_42975,N_41122,N_41772);
xnor U42976 (N_42976,N_41174,N_40856);
nor U42977 (N_42977,N_40099,N_41946);
nand U42978 (N_42978,N_40752,N_40131);
xor U42979 (N_42979,N_41006,N_40141);
and U42980 (N_42980,N_40523,N_41924);
nor U42981 (N_42981,N_40112,N_42192);
or U42982 (N_42982,N_40791,N_40248);
nand U42983 (N_42983,N_42272,N_41098);
nor U42984 (N_42984,N_41993,N_41620);
or U42985 (N_42985,N_40377,N_42434);
nor U42986 (N_42986,N_40384,N_41578);
nor U42987 (N_42987,N_41448,N_41450);
or U42988 (N_42988,N_41237,N_42386);
xor U42989 (N_42989,N_41262,N_40181);
or U42990 (N_42990,N_41302,N_40701);
xor U42991 (N_42991,N_42198,N_42216);
and U42992 (N_42992,N_42059,N_40051);
nor U42993 (N_42993,N_41139,N_40309);
or U42994 (N_42994,N_40014,N_40935);
or U42995 (N_42995,N_41371,N_41614);
xor U42996 (N_42996,N_41762,N_41041);
and U42997 (N_42997,N_40697,N_41245);
or U42998 (N_42998,N_42464,N_40183);
nand U42999 (N_42999,N_42034,N_41525);
nor U43000 (N_43000,N_41030,N_41413);
and U43001 (N_43001,N_40427,N_42083);
nor U43002 (N_43002,N_41246,N_41603);
or U43003 (N_43003,N_41254,N_40991);
and U43004 (N_43004,N_40760,N_42148);
or U43005 (N_43005,N_40682,N_40827);
nand U43006 (N_43006,N_41805,N_41419);
nand U43007 (N_43007,N_40026,N_41014);
xnor U43008 (N_43008,N_40722,N_40468);
or U43009 (N_43009,N_40897,N_42130);
nand U43010 (N_43010,N_41538,N_40946);
and U43011 (N_43011,N_41024,N_40510);
nand U43012 (N_43012,N_40890,N_42305);
xor U43013 (N_43013,N_42024,N_42129);
or U43014 (N_43014,N_41724,N_40773);
and U43015 (N_43015,N_41615,N_42027);
or U43016 (N_43016,N_42090,N_41965);
or U43017 (N_43017,N_40260,N_41656);
and U43018 (N_43018,N_41705,N_40398);
xor U43019 (N_43019,N_41765,N_40750);
and U43020 (N_43020,N_40675,N_41432);
and U43021 (N_43021,N_40658,N_41149);
or U43022 (N_43022,N_41337,N_41912);
or U43023 (N_43023,N_40207,N_41796);
or U43024 (N_43024,N_40109,N_40303);
xnor U43025 (N_43025,N_41892,N_41564);
or U43026 (N_43026,N_41428,N_40018);
and U43027 (N_43027,N_41453,N_42232);
xor U43028 (N_43028,N_42415,N_42408);
and U43029 (N_43029,N_40624,N_40578);
and U43030 (N_43030,N_42134,N_42096);
nor U43031 (N_43031,N_41529,N_41406);
nand U43032 (N_43032,N_42019,N_42254);
or U43033 (N_43033,N_41005,N_40104);
nor U43034 (N_43034,N_41990,N_42185);
or U43035 (N_43035,N_41117,N_41307);
or U43036 (N_43036,N_40435,N_41877);
nand U43037 (N_43037,N_40134,N_40113);
nand U43038 (N_43038,N_40146,N_42270);
and U43039 (N_43039,N_41314,N_41038);
xnor U43040 (N_43040,N_40812,N_40625);
nor U43041 (N_43041,N_41061,N_40918);
nor U43042 (N_43042,N_40033,N_40460);
or U43043 (N_43043,N_40186,N_41547);
nand U43044 (N_43044,N_42331,N_42455);
or U43045 (N_43045,N_42467,N_40725);
xor U43046 (N_43046,N_40062,N_41144);
xor U43047 (N_43047,N_41534,N_41734);
nor U43048 (N_43048,N_41381,N_40374);
nand U43049 (N_43049,N_40236,N_42314);
and U43050 (N_43050,N_41883,N_41211);
xnor U43051 (N_43051,N_40275,N_41721);
nand U43052 (N_43052,N_41672,N_41461);
nand U43053 (N_43053,N_40615,N_40971);
and U43054 (N_43054,N_41028,N_40239);
or U43055 (N_43055,N_42336,N_41845);
nand U43056 (N_43056,N_40904,N_41025);
nor U43057 (N_43057,N_40453,N_40592);
and U43058 (N_43058,N_40084,N_42098);
xor U43059 (N_43059,N_40967,N_42406);
xor U43060 (N_43060,N_40039,N_40337);
nor U43061 (N_43061,N_42069,N_42412);
or U43062 (N_43062,N_40194,N_42010);
or U43063 (N_43063,N_41255,N_41394);
nor U43064 (N_43064,N_41625,N_40820);
or U43065 (N_43065,N_40324,N_41475);
and U43066 (N_43066,N_41376,N_41785);
and U43067 (N_43067,N_42160,N_40171);
nor U43068 (N_43068,N_41242,N_40619);
nor U43069 (N_43069,N_40389,N_40294);
xnor U43070 (N_43070,N_40356,N_41546);
or U43071 (N_43071,N_41933,N_41957);
nor U43072 (N_43072,N_41844,N_40240);
or U43073 (N_43073,N_42426,N_41789);
xor U43074 (N_43074,N_41843,N_41626);
nor U43075 (N_43075,N_42061,N_41296);
or U43076 (N_43076,N_42094,N_41377);
and U43077 (N_43077,N_40011,N_41942);
xnor U43078 (N_43078,N_42396,N_41227);
or U43079 (N_43079,N_41077,N_40287);
and U43080 (N_43080,N_40917,N_40739);
nand U43081 (N_43081,N_40068,N_42065);
xor U43082 (N_43082,N_40148,N_40164);
nand U43083 (N_43083,N_41407,N_40016);
or U43084 (N_43084,N_42390,N_40841);
nand U43085 (N_43085,N_41654,N_41675);
xor U43086 (N_43086,N_41268,N_41420);
nand U43087 (N_43087,N_40709,N_42051);
xnor U43088 (N_43088,N_42193,N_40984);
or U43089 (N_43089,N_41020,N_40732);
and U43090 (N_43090,N_41878,N_40903);
and U43091 (N_43091,N_41496,N_41898);
or U43092 (N_43092,N_40612,N_40323);
or U43093 (N_43093,N_41189,N_40448);
nand U43094 (N_43094,N_40963,N_40038);
nand U43095 (N_43095,N_40478,N_40333);
nor U43096 (N_43096,N_40008,N_41311);
xnor U43097 (N_43097,N_40158,N_41683);
nand U43098 (N_43098,N_40217,N_41455);
and U43099 (N_43099,N_40403,N_41996);
nor U43100 (N_43100,N_41261,N_42240);
nor U43101 (N_43101,N_40762,N_40945);
xor U43102 (N_43102,N_41601,N_42092);
nor U43103 (N_43103,N_41222,N_41959);
nand U43104 (N_43104,N_41655,N_41387);
nand U43105 (N_43105,N_42175,N_42373);
nand U43106 (N_43106,N_40605,N_40957);
nor U43107 (N_43107,N_42076,N_40560);
nand U43108 (N_43108,N_40786,N_40740);
and U43109 (N_43109,N_40582,N_41928);
and U43110 (N_43110,N_41973,N_40421);
nand U43111 (N_43111,N_42003,N_41458);
nor U43112 (N_43112,N_42058,N_41707);
and U43113 (N_43113,N_41435,N_40972);
or U43114 (N_43114,N_40968,N_41544);
xor U43115 (N_43115,N_40407,N_40093);
nor U43116 (N_43116,N_41408,N_40969);
and U43117 (N_43117,N_41563,N_42359);
nor U43118 (N_43118,N_41177,N_40446);
xnor U43119 (N_43119,N_40539,N_42454);
or U43120 (N_43120,N_41800,N_40641);
xor U43121 (N_43121,N_41937,N_41493);
xor U43122 (N_43122,N_41995,N_40120);
nand U43123 (N_43123,N_41249,N_41313);
nor U43124 (N_43124,N_41756,N_42139);
or U43125 (N_43125,N_40717,N_41584);
nand U43126 (N_43126,N_41229,N_40659);
or U43127 (N_43127,N_42400,N_41882);
or U43128 (N_43128,N_41763,N_40472);
or U43129 (N_43129,N_40990,N_40759);
or U43130 (N_43130,N_40543,N_41438);
xor U43131 (N_43131,N_42372,N_40915);
nand U43132 (N_43132,N_41929,N_40474);
xnor U43133 (N_43133,N_41688,N_40954);
xnor U43134 (N_43134,N_42268,N_40178);
or U43135 (N_43135,N_40705,N_40892);
xor U43136 (N_43136,N_40077,N_40059);
xor U43137 (N_43137,N_41835,N_40563);
xor U43138 (N_43138,N_42155,N_41684);
nand U43139 (N_43139,N_40129,N_41108);
and U43140 (N_43140,N_40293,N_41182);
nor U43141 (N_43141,N_41490,N_40196);
nand U43142 (N_43142,N_42441,N_41104);
xnor U43143 (N_43143,N_41148,N_42057);
nand U43144 (N_43144,N_42021,N_42153);
and U43145 (N_43145,N_40639,N_40891);
or U43146 (N_43146,N_41503,N_41323);
and U43147 (N_43147,N_40072,N_41473);
nor U43148 (N_43148,N_40063,N_42445);
or U43149 (N_43149,N_41537,N_41145);
xor U43150 (N_43150,N_41250,N_40594);
xnor U43151 (N_43151,N_40119,N_42169);
nand U43152 (N_43152,N_41172,N_40731);
xor U43153 (N_43153,N_41559,N_42391);
or U43154 (N_43154,N_41645,N_40743);
nor U43155 (N_43155,N_40272,N_41048);
xor U43156 (N_43156,N_40797,N_42291);
or U43157 (N_43157,N_40803,N_41066);
nor U43158 (N_43158,N_41913,N_42246);
xor U43159 (N_43159,N_41212,N_42354);
and U43160 (N_43160,N_41941,N_40256);
nand U43161 (N_43161,N_40295,N_40670);
nand U43162 (N_43162,N_42312,N_41488);
xor U43163 (N_43163,N_41749,N_40953);
xnor U43164 (N_43164,N_40350,N_42290);
and U43165 (N_43165,N_41000,N_41888);
xor U43166 (N_43166,N_41583,N_41049);
nand U43167 (N_43167,N_40032,N_41702);
nor U43168 (N_43168,N_40958,N_40636);
nand U43169 (N_43169,N_40493,N_40927);
or U43170 (N_43170,N_40137,N_41304);
nor U43171 (N_43171,N_40025,N_41259);
nor U43172 (N_43172,N_41141,N_40844);
nand U43173 (N_43173,N_41495,N_42202);
xor U43174 (N_43174,N_41106,N_41112);
or U43175 (N_43175,N_42084,N_41986);
xor U43176 (N_43176,N_40078,N_40255);
or U43177 (N_43177,N_42293,N_40878);
and U43178 (N_43178,N_41801,N_41828);
nor U43179 (N_43179,N_41469,N_41396);
or U43180 (N_43180,N_42328,N_41670);
nor U43181 (N_43181,N_42208,N_40996);
nor U43182 (N_43182,N_41240,N_41466);
nand U43183 (N_43183,N_40308,N_41107);
nand U43184 (N_43184,N_40320,N_42460);
and U43185 (N_43185,N_40244,N_41281);
nor U43186 (N_43186,N_40496,N_41903);
nand U43187 (N_43187,N_41963,N_41401);
nand U43188 (N_43188,N_42122,N_40622);
xnor U43189 (N_43189,N_42409,N_42309);
nand U43190 (N_43190,N_40720,N_40964);
nand U43191 (N_43191,N_42430,N_40282);
or U43192 (N_43192,N_41740,N_41697);
or U43193 (N_43193,N_40824,N_41948);
nor U43194 (N_43194,N_40532,N_41606);
or U43195 (N_43195,N_40536,N_42055);
xor U43196 (N_43196,N_42172,N_40586);
or U43197 (N_43197,N_41065,N_41783);
and U43198 (N_43198,N_40506,N_42082);
nand U43199 (N_43199,N_41476,N_40473);
xnor U43200 (N_43200,N_40761,N_41485);
nor U43201 (N_43201,N_42209,N_41221);
nor U43202 (N_43202,N_40253,N_41829);
nor U43203 (N_43203,N_41981,N_40648);
or U43204 (N_43204,N_42446,N_42103);
nand U43205 (N_43205,N_40728,N_41269);
and U43206 (N_43206,N_41923,N_41650);
xor U43207 (N_43207,N_40608,N_42326);
or U43208 (N_43208,N_41374,N_41949);
nor U43209 (N_43209,N_40326,N_42410);
nor U43210 (N_43210,N_40851,N_41422);
and U43211 (N_43211,N_41479,N_42303);
nor U43212 (N_43212,N_40597,N_42085);
nor U43213 (N_43213,N_40729,N_40167);
nor U43214 (N_43214,N_40702,N_40028);
nor U43215 (N_43215,N_40193,N_41720);
nor U43216 (N_43216,N_40318,N_40581);
xor U43217 (N_43217,N_41732,N_40853);
nand U43218 (N_43218,N_42161,N_41073);
nor U43219 (N_43219,N_40557,N_41921);
or U43220 (N_43220,N_42490,N_40343);
nand U43221 (N_43221,N_42047,N_42256);
nor U43222 (N_43222,N_40114,N_41926);
xor U43223 (N_43223,N_41860,N_40949);
xnor U43224 (N_43224,N_41849,N_42345);
nand U43225 (N_43225,N_40475,N_41244);
nand U43226 (N_43226,N_40589,N_40311);
and U43227 (N_43227,N_41348,N_42329);
and U43228 (N_43228,N_40766,N_40476);
nand U43229 (N_43229,N_42043,N_40098);
and U43230 (N_43230,N_40681,N_41343);
nand U43231 (N_43231,N_41838,N_41577);
and U43232 (N_43232,N_40373,N_41792);
nand U43233 (N_43233,N_40606,N_42471);
and U43234 (N_43234,N_41223,N_41520);
nor U43235 (N_43235,N_42020,N_40555);
and U43236 (N_43236,N_41969,N_40961);
xnor U43237 (N_43237,N_40321,N_40211);
nor U43238 (N_43238,N_41273,N_40577);
nor U43239 (N_43239,N_40980,N_40426);
xor U43240 (N_43240,N_42217,N_41809);
and U43241 (N_43241,N_41402,N_41890);
and U43242 (N_43242,N_41716,N_42429);
xnor U43243 (N_43243,N_40234,N_42184);
nor U43244 (N_43244,N_40749,N_41744);
nand U43245 (N_43245,N_42127,N_42381);
nor U43246 (N_43246,N_40637,N_40463);
or U43247 (N_43247,N_40526,N_41819);
and U43248 (N_43248,N_40835,N_41305);
xnor U43249 (N_43249,N_40602,N_40023);
and U43250 (N_43250,N_40361,N_41795);
and U43251 (N_43251,N_40061,N_41295);
and U43252 (N_43252,N_41120,N_41652);
and U43253 (N_43253,N_40719,N_40499);
nor U43254 (N_43254,N_41241,N_42079);
nand U43255 (N_43255,N_41327,N_40756);
xor U43256 (N_43256,N_40836,N_41513);
xnor U43257 (N_43257,N_41185,N_40351);
nor U43258 (N_43258,N_41159,N_41517);
and U43259 (N_43259,N_40494,N_41366);
xnor U43260 (N_43260,N_42279,N_40461);
nand U43261 (N_43261,N_41616,N_40881);
and U43262 (N_43262,N_41187,N_42002);
and U43263 (N_43263,N_40386,N_41320);
and U43264 (N_43264,N_41263,N_40934);
or U43265 (N_43265,N_40538,N_42075);
and U43266 (N_43266,N_40342,N_41579);
xor U43267 (N_43267,N_42013,N_42138);
xnor U43268 (N_43268,N_41214,N_40235);
nand U43269 (N_43269,N_40364,N_42366);
or U43270 (N_43270,N_40442,N_42313);
nand U43271 (N_43271,N_41113,N_41359);
xnor U43272 (N_43272,N_40884,N_41640);
xnor U43273 (N_43273,N_42398,N_42378);
or U43274 (N_43274,N_42143,N_40058);
nand U43275 (N_43275,N_40276,N_40163);
xnor U43276 (N_43276,N_41317,N_42387);
or U43277 (N_43277,N_40199,N_41964);
nand U43278 (N_43278,N_41536,N_41330);
nand U43279 (N_43279,N_42403,N_41859);
nor U43280 (N_43280,N_40189,N_40432);
or U43281 (N_43281,N_40699,N_40789);
and U43282 (N_43282,N_40043,N_40328);
nor U43283 (N_43283,N_40676,N_40583);
and U43284 (N_43284,N_42016,N_41459);
nand U43285 (N_43285,N_40000,N_41875);
nand U43286 (N_43286,N_42458,N_41841);
xnor U43287 (N_43287,N_41812,N_40973);
nand U43288 (N_43288,N_40482,N_41470);
xor U43289 (N_43289,N_40340,N_41412);
and U43290 (N_43290,N_41704,N_40607);
nor U43291 (N_43291,N_40414,N_41339);
and U43292 (N_43292,N_40977,N_42117);
nor U43293 (N_43293,N_40599,N_42137);
nor U43294 (N_43294,N_41329,N_41533);
nand U43295 (N_43295,N_42033,N_40994);
or U43296 (N_43296,N_42362,N_41985);
nand U43297 (N_43297,N_40198,N_41680);
nand U43298 (N_43298,N_40570,N_42437);
nand U43299 (N_43299,N_41433,N_40277);
nand U43300 (N_43300,N_41425,N_40115);
or U43301 (N_43301,N_40535,N_41060);
or U43302 (N_43302,N_40052,N_41151);
nand U43303 (N_43303,N_42394,N_42200);
xor U43304 (N_43304,N_40923,N_41723);
xnor U43305 (N_43305,N_40850,N_42248);
nor U43306 (N_43306,N_41658,N_40630);
nand U43307 (N_43307,N_41669,N_41292);
or U43308 (N_43308,N_40332,N_41745);
nand U43309 (N_43309,N_41379,N_42089);
nand U43310 (N_43310,N_40393,N_41370);
nor U43311 (N_43311,N_41270,N_40687);
or U43312 (N_43312,N_42062,N_42288);
xnor U43313 (N_43313,N_40177,N_41775);
or U43314 (N_43314,N_41439,N_40383);
and U43315 (N_43315,N_41874,N_40238);
or U43316 (N_43316,N_41158,N_41830);
and U43317 (N_43317,N_41975,N_41955);
and U43318 (N_43318,N_41170,N_40243);
and U43319 (N_43319,N_40774,N_42247);
and U43320 (N_43320,N_40021,N_41310);
xnor U43321 (N_43321,N_40015,N_41498);
nand U43322 (N_43322,N_41225,N_41162);
nor U43323 (N_43323,N_40470,N_42211);
and U43324 (N_43324,N_42371,N_40744);
xnor U43325 (N_43325,N_40710,N_42131);
nand U43326 (N_43326,N_40767,N_42459);
and U43327 (N_43327,N_40959,N_41668);
or U43328 (N_43328,N_41471,N_40108);
xnor U43329 (N_43329,N_40799,N_40301);
xor U43330 (N_43330,N_40341,N_41693);
nor U43331 (N_43331,N_42311,N_40511);
nand U43332 (N_43332,N_41082,N_41944);
nor U43333 (N_43333,N_40368,N_42477);
nand U43334 (N_43334,N_41585,N_41316);
nand U43335 (N_43335,N_41251,N_41492);
and U43336 (N_43336,N_40428,N_40901);
nor U43337 (N_43337,N_40735,N_40723);
nor U43338 (N_43338,N_41758,N_40956);
and U43339 (N_43339,N_40939,N_41196);
or U43340 (N_43340,N_41331,N_41592);
nand U43341 (N_43341,N_41280,N_41731);
nor U43342 (N_43342,N_41971,N_40241);
and U43343 (N_43343,N_41771,N_40745);
or U43344 (N_43344,N_41007,N_40669);
nand U43345 (N_43345,N_40804,N_41265);
nand U43346 (N_43346,N_40490,N_40424);
xnor U43347 (N_43347,N_40488,N_41218);
nor U43348 (N_43348,N_40512,N_41489);
nand U43349 (N_43349,N_41824,N_41644);
and U43350 (N_43350,N_41910,N_40989);
nor U43351 (N_43351,N_40593,N_40465);
or U43352 (N_43352,N_41121,N_42220);
and U43353 (N_43353,N_41076,N_41403);
xor U43354 (N_43354,N_40347,N_42004);
nor U43355 (N_43355,N_40227,N_41667);
nor U43356 (N_43356,N_40546,N_40349);
xor U43357 (N_43357,N_41905,N_40106);
nand U43358 (N_43358,N_41665,N_40609);
and U43359 (N_43359,N_40336,N_41092);
nand U43360 (N_43360,N_41232,N_40694);
xnor U43361 (N_43361,N_42255,N_42145);
and U43362 (N_43362,N_41657,N_42194);
nand U43363 (N_43363,N_40304,N_41782);
nor U43364 (N_43364,N_42262,N_41037);
or U43365 (N_43365,N_41821,N_40462);
nor U43366 (N_43366,N_40808,N_42049);
xnor U43367 (N_43367,N_41979,N_41414);
xnor U43368 (N_43368,N_41730,N_40376);
or U43369 (N_43369,N_41368,N_40190);
and U43370 (N_43370,N_40216,N_41443);
nand U43371 (N_43371,N_41357,N_40672);
and U43372 (N_43372,N_40412,N_41224);
and U43373 (N_43373,N_41833,N_41612);
xor U43374 (N_43374,N_40913,N_41248);
nor U43375 (N_43375,N_41815,N_41662);
nor U43376 (N_43376,N_40780,N_40307);
xnor U43377 (N_43377,N_41070,N_40552);
and U43378 (N_43378,N_40034,N_42323);
and U43379 (N_43379,N_41260,N_40423);
nand U43380 (N_43380,N_42121,N_40623);
xnor U43381 (N_43381,N_41852,N_40359);
nor U43382 (N_43382,N_41943,N_41855);
xor U43383 (N_43383,N_40727,N_40149);
and U43384 (N_43384,N_42110,N_41925);
nand U43385 (N_43385,N_41474,N_41555);
nor U43386 (N_43386,N_40920,N_40150);
and U43387 (N_43387,N_40346,N_41863);
and U43388 (N_43388,N_41802,N_40686);
and U43389 (N_43389,N_42423,N_40908);
and U43390 (N_43390,N_42156,N_42404);
and U43391 (N_43391,N_42042,N_40401);
and U43392 (N_43392,N_40312,N_42144);
and U43393 (N_43393,N_42125,N_40693);
nor U43394 (N_43394,N_40285,N_41570);
and U43395 (N_43395,N_41127,N_42337);
nor U43396 (N_43396,N_42401,N_40437);
and U43397 (N_43397,N_41900,N_42438);
nand U43398 (N_43398,N_41617,N_41303);
nand U43399 (N_43399,N_41138,N_40327);
nand U43400 (N_43400,N_41238,N_40889);
or U43401 (N_43401,N_42242,N_41738);
and U43402 (N_43402,N_41516,N_41383);
xor U43403 (N_43403,N_41574,N_42102);
and U43404 (N_43404,N_41338,N_41213);
and U43405 (N_43405,N_41610,N_41021);
nor U43406 (N_43406,N_41123,N_41389);
nor U43407 (N_43407,N_40861,N_41750);
nand U43408 (N_43408,N_40649,N_40322);
or U43409 (N_43409,N_42053,N_40540);
nor U43410 (N_43410,N_42045,N_41766);
and U43411 (N_43411,N_40514,N_40788);
nor U43412 (N_43412,N_42405,N_42237);
and U43413 (N_43413,N_40874,N_40188);
nand U43414 (N_43414,N_41282,N_42060);
and U43415 (N_43415,N_41358,N_40143);
xor U43416 (N_43416,N_40880,N_40937);
nand U43417 (N_43417,N_42432,N_41565);
xnor U43418 (N_43418,N_40409,N_41715);
nor U43419 (N_43419,N_40222,N_42447);
nand U43420 (N_43420,N_40618,N_41201);
xnor U43421 (N_43421,N_40600,N_40955);
or U43422 (N_43422,N_40369,N_40863);
or U43423 (N_43423,N_41501,N_42276);
and U43424 (N_43424,N_41257,N_42297);
or U43425 (N_43425,N_41217,N_40807);
or U43426 (N_43426,N_41932,N_40685);
and U43427 (N_43427,N_41416,N_41722);
and U43428 (N_43428,N_40182,N_40173);
xor U43429 (N_43429,N_40085,N_40345);
nand U43430 (N_43430,N_40895,N_42420);
and U43431 (N_43431,N_41344,N_40549);
or U43432 (N_43432,N_42214,N_40263);
or U43433 (N_43433,N_42166,N_40279);
xor U43434 (N_43434,N_40339,N_40505);
xnor U43435 (N_43435,N_41053,N_41345);
nor U43436 (N_43436,N_42025,N_41791);
nor U43437 (N_43437,N_41385,N_41100);
and U43438 (N_43438,N_42164,N_40445);
nor U43439 (N_43439,N_40261,N_41764);
and U43440 (N_43440,N_41562,N_42296);
and U43441 (N_43441,N_40107,N_40111);
and U43442 (N_43442,N_40886,N_41831);
or U43443 (N_43443,N_42015,N_40489);
nand U43444 (N_43444,N_40019,N_41019);
or U43445 (N_43445,N_40254,N_40491);
nor U43446 (N_43446,N_40576,N_40885);
nor U43447 (N_43447,N_40257,N_42064);
nand U43448 (N_43448,N_40667,N_40082);
nand U43449 (N_43449,N_41405,N_42448);
nor U43450 (N_43450,N_41621,N_41203);
or U43451 (N_43451,N_40204,N_41010);
nor U43452 (N_43452,N_41445,N_41523);
nor U43453 (N_43453,N_41571,N_42351);
or U43454 (N_43454,N_42187,N_41692);
xnor U43455 (N_43455,N_41197,N_41497);
or U43456 (N_43456,N_41169,N_41966);
xor U43457 (N_43457,N_41115,N_41062);
or U43458 (N_43458,N_41718,N_41404);
xor U43459 (N_43459,N_41618,N_42157);
xnor U43460 (N_43460,N_41291,N_42265);
and U43461 (N_43461,N_42007,N_42097);
nand U43462 (N_43462,N_41472,N_41467);
nand U43463 (N_43463,N_41974,N_41183);
and U43464 (N_43464,N_41388,N_41514);
xor U43465 (N_43465,N_40757,N_41029);
and U43466 (N_43466,N_40537,N_42368);
nor U43467 (N_43467,N_40692,N_40651);
xor U43468 (N_43468,N_40081,N_40832);
nand U43469 (N_43469,N_42112,N_40700);
or U43470 (N_43470,N_41378,N_41173);
xnor U43471 (N_43471,N_40995,N_40509);
nor U43472 (N_43472,N_42006,N_41552);
or U43473 (N_43473,N_40830,N_41312);
nor U43474 (N_43474,N_41057,N_41220);
and U43475 (N_43475,N_41105,N_41622);
nand U43476 (N_43476,N_42397,N_41980);
nand U43477 (N_43477,N_40839,N_40730);
nor U43478 (N_43478,N_41719,N_42071);
and U43479 (N_43479,N_42327,N_41978);
or U43480 (N_43480,N_42106,N_40632);
nor U43481 (N_43481,N_41216,N_40003);
or U43482 (N_43482,N_41823,N_41726);
nand U43483 (N_43483,N_42317,N_40580);
xnor U43484 (N_43484,N_42243,N_42427);
nand U43485 (N_43485,N_40591,N_40269);
or U43486 (N_43486,N_41998,N_40778);
and U43487 (N_43487,N_41166,N_41887);
and U43488 (N_43488,N_40653,N_42074);
xnor U43489 (N_43489,N_41071,N_40391);
nand U43490 (N_43490,N_40556,N_41161);
or U43491 (N_43491,N_42072,N_40503);
and U43492 (N_43492,N_42428,N_40367);
and U43493 (N_43493,N_41132,N_41032);
xnor U43494 (N_43494,N_41356,N_40290);
xor U43495 (N_43495,N_40713,N_42252);
nor U43496 (N_43496,N_40598,N_40714);
or U43497 (N_43497,N_42179,N_41968);
or U43498 (N_43498,N_41632,N_40486);
nor U43499 (N_43499,N_42421,N_40922);
xnor U43500 (N_43500,N_40679,N_41902);
or U43501 (N_43501,N_41522,N_41951);
nand U43502 (N_43502,N_40698,N_41568);
or U43503 (N_43503,N_41499,N_40695);
and U43504 (N_43504,N_41560,N_41508);
or U43505 (N_43505,N_40075,N_40678);
nor U43506 (N_43506,N_40677,N_40152);
nor U43507 (N_43507,N_40796,N_41256);
xnor U43508 (N_43508,N_42389,N_41917);
nor U43509 (N_43509,N_42294,N_42224);
or U43510 (N_43510,N_40502,N_41920);
nor U43511 (N_43511,N_40931,N_40330);
nand U43512 (N_43512,N_41101,N_42100);
nor U43513 (N_43513,N_42417,N_41457);
and U43514 (N_43514,N_40811,N_41803);
nor U43515 (N_43515,N_41894,N_41984);
xor U43516 (N_43516,N_42300,N_42188);
nor U43517 (N_43517,N_40300,N_42363);
and U43518 (N_43518,N_41399,N_40932);
and U43519 (N_43519,N_41130,N_41482);
xnor U43520 (N_43520,N_41275,N_40180);
nand U43521 (N_43521,N_40288,N_42154);
xor U43522 (N_43522,N_41751,N_40439);
nand U43523 (N_43523,N_40220,N_40857);
nand U43524 (N_43524,N_40487,N_40165);
or U43525 (N_43525,N_42287,N_41687);
xnor U43526 (N_43526,N_40007,N_40053);
xor U43527 (N_43527,N_40715,N_41454);
nor U43528 (N_43528,N_40201,N_40116);
nor U43529 (N_43529,N_42245,N_40252);
nor U43530 (N_43530,N_40070,N_40378);
and U43531 (N_43531,N_41195,N_42080);
and U43532 (N_43532,N_41334,N_41382);
and U43533 (N_43533,N_41524,N_41641);
and U43534 (N_43534,N_40655,N_41961);
or U43535 (N_43535,N_41085,N_41940);
and U43536 (N_43536,N_41862,N_40734);
xor U43537 (N_43537,N_40521,N_40876);
nand U43538 (N_43538,N_41134,N_41191);
xor U43539 (N_43539,N_41079,N_40352);
nand U43540 (N_43540,N_41126,N_42032);
or U43541 (N_43541,N_41873,N_42497);
and U43542 (N_43542,N_40738,N_41176);
nor U43543 (N_43543,N_41198,N_42302);
nand U43544 (N_43544,N_40335,N_41810);
nand U43545 (N_43545,N_41074,N_41548);
or U43546 (N_43546,N_41294,N_42258);
nand U43547 (N_43547,N_42282,N_40988);
or U43548 (N_43548,N_41140,N_40042);
nor U43549 (N_43549,N_41958,N_40268);
and U43550 (N_43550,N_40249,N_40006);
xnor U43551 (N_43551,N_41864,N_41157);
or U43552 (N_43552,N_41309,N_40665);
nand U43553 (N_43553,N_42411,N_41834);
nand U43554 (N_43554,N_41386,N_42017);
nor U43555 (N_43555,N_42023,N_41009);
xnor U43556 (N_43556,N_41252,N_40802);
nor U43557 (N_43557,N_41678,N_41992);
xor U43558 (N_43558,N_41931,N_40822);
and U43559 (N_43559,N_41207,N_40258);
or U43560 (N_43560,N_42022,N_40291);
or U43561 (N_43561,N_40110,N_40360);
and U43562 (N_43562,N_41204,N_41804);
xor U43563 (N_43563,N_40464,N_42367);
nor U43564 (N_43564,N_41780,N_41976);
and U43565 (N_43565,N_40419,N_40815);
nor U43566 (N_43566,N_40821,N_41001);
nand U43567 (N_43567,N_41397,N_40941);
nor U43568 (N_43568,N_41518,N_40179);
and U43569 (N_43569,N_40457,N_40358);
nand U43570 (N_43570,N_41794,N_40721);
or U43571 (N_43571,N_42119,N_40477);
and U43572 (N_43572,N_42439,N_40022);
and U43573 (N_43573,N_40707,N_42182);
nor U43574 (N_43574,N_41147,N_41045);
nand U43575 (N_43575,N_42180,N_40981);
and U43576 (N_43576,N_42234,N_41659);
and U43577 (N_43577,N_41581,N_42267);
xor U43578 (N_43578,N_41017,N_42418);
xnor U43579 (N_43579,N_40664,N_40817);
nor U43580 (N_43580,N_41500,N_41042);
xor U43581 (N_43581,N_41634,N_40528);
nor U43582 (N_43582,N_41512,N_42344);
xor U43583 (N_43583,N_42274,N_41856);
or U43584 (N_43584,N_42136,N_42109);
xor U43585 (N_43585,N_42086,N_40274);
nor U43586 (N_43586,N_40166,N_42348);
nor U43587 (N_43587,N_40542,N_42343);
or U43588 (N_43588,N_42073,N_42142);
xnor U43589 (N_43589,N_42236,N_41056);
or U43590 (N_43590,N_42229,N_42365);
nor U43591 (N_43591,N_41742,N_41013);
nor U43592 (N_43592,N_41089,N_40520);
or U43593 (N_43593,N_42478,N_41328);
xor U43594 (N_43594,N_41737,N_42275);
xor U43595 (N_43595,N_40064,N_41897);
xnor U43596 (N_43596,N_40871,N_40395);
nand U43597 (N_43597,N_42320,N_41846);
or U43598 (N_43598,N_42424,N_40671);
xnor U43599 (N_43599,N_41623,N_40089);
nand U43600 (N_43600,N_40684,N_41347);
and U43601 (N_43601,N_40654,N_41781);
and U43602 (N_43602,N_40656,N_41468);
xor U43603 (N_43603,N_40049,N_41051);
or U43604 (N_43604,N_42213,N_42476);
xnor U43605 (N_43605,N_41748,N_40635);
and U43606 (N_43606,N_42241,N_40777);
and U43607 (N_43607,N_41770,N_42219);
and U43608 (N_43608,N_41907,N_42105);
nand U43609 (N_43609,N_42292,N_41575);
xnor U43610 (N_43610,N_42482,N_41031);
or U43611 (N_43611,N_41604,N_41922);
and U43612 (N_43612,N_42260,N_40298);
nor U43613 (N_43613,N_41558,N_41034);
and U43614 (N_43614,N_40584,N_40628);
nor U43615 (N_43615,N_40657,N_41477);
nand U43616 (N_43616,N_41573,N_40136);
nand U43617 (N_43617,N_40080,N_40399);
xnor U43618 (N_43618,N_40174,N_41896);
or U43619 (N_43619,N_41899,N_41619);
nand U43620 (N_43620,N_41663,N_42277);
nand U43621 (N_43621,N_40569,N_40688);
and U43622 (N_43622,N_40471,N_40192);
or U43623 (N_43623,N_41813,N_40870);
nor U43624 (N_43624,N_40151,N_41793);
and U43625 (N_43625,N_40092,N_40894);
nor U43626 (N_43626,N_42162,N_41036);
xnor U43627 (N_43627,N_40264,N_40299);
nor U43628 (N_43628,N_40627,N_42316);
nor U43629 (N_43629,N_40547,N_41988);
and U43630 (N_43630,N_41550,N_40611);
nand U43631 (N_43631,N_40027,N_42355);
and U43632 (N_43632,N_42462,N_40215);
nand U43633 (N_43633,N_41215,N_41478);
and U43634 (N_43634,N_40997,N_42196);
nor U43635 (N_43635,N_40926,N_40858);
nand U43636 (N_43636,N_40933,N_41653);
or U43637 (N_43637,N_40747,N_42228);
nor U43638 (N_43638,N_40344,N_40504);
xor U43639 (N_43639,N_41569,N_40845);
or U43640 (N_43640,N_42278,N_40633);
and U43641 (N_43641,N_40986,N_42257);
xor U43642 (N_43642,N_40928,N_40680);
or U43643 (N_43643,N_41384,N_40864);
nor U43644 (N_43644,N_41300,N_40447);
nor U43645 (N_43645,N_41784,N_42078);
nor U43646 (N_43646,N_41093,N_42472);
nand U43647 (N_43647,N_41421,N_41787);
nand U43648 (N_43648,N_40938,N_41788);
nor U43649 (N_43649,N_40801,N_40037);
nor U43650 (N_43650,N_40562,N_41519);
or U43651 (N_43651,N_41364,N_42442);
nand U43652 (N_43652,N_42149,N_41363);
xor U43653 (N_43653,N_41950,N_41759);
nand U43654 (N_43654,N_40846,N_42486);
nand U43655 (N_43655,N_40898,N_40036);
or U43656 (N_43656,N_40787,N_40251);
and U43657 (N_43657,N_42039,N_40711);
nand U43658 (N_43658,N_41059,N_41272);
and U43659 (N_43659,N_40265,N_42123);
xor U43660 (N_43660,N_40718,N_42392);
or U43661 (N_43661,N_41168,N_40314);
nand U43662 (N_43662,N_40002,N_41375);
nor U43663 (N_43663,N_41410,N_40449);
nand U43664 (N_43664,N_41184,N_40127);
nand U43665 (N_43665,N_41954,N_41200);
or U43666 (N_43666,N_42251,N_42286);
nand U43667 (N_43667,N_40159,N_41607);
xor U43668 (N_43668,N_40862,N_41696);
or U43669 (N_43669,N_41440,N_41373);
or U43670 (N_43670,N_41820,N_42324);
nor U43671 (N_43671,N_41437,N_40613);
and U43672 (N_43672,N_41886,N_40250);
nand U43673 (N_43673,N_40531,N_40975);
or U43674 (N_43674,N_40983,N_40673);
nor U43675 (N_43675,N_40666,N_42077);
and U43676 (N_43676,N_41046,N_40480);
and U43677 (N_43677,N_41956,N_42221);
nor U43678 (N_43678,N_40195,N_41027);
nand U43679 (N_43679,N_42183,N_40838);
xnor U43680 (N_43680,N_42046,N_42484);
or U43681 (N_43681,N_40588,N_41355);
xnor U43682 (N_43682,N_41154,N_41167);
nand U43683 (N_43683,N_42048,N_41822);
or U43684 (N_43684,N_41511,N_42088);
nor U43685 (N_43685,N_41464,N_40912);
and U43686 (N_43686,N_40313,N_40823);
xnor U43687 (N_43687,N_40297,N_42264);
nor U43688 (N_43688,N_42087,N_40663);
xor U43689 (N_43689,N_40259,N_41352);
or U43690 (N_43690,N_41709,N_42116);
or U43691 (N_43691,N_40944,N_40816);
and U43692 (N_43692,N_40117,N_42284);
nor U43693 (N_43693,N_41953,N_41114);
and U43694 (N_43694,N_41541,N_42451);
nand U43695 (N_43695,N_40551,N_41234);
nor U43696 (N_43696,N_42038,N_41695);
nand U43697 (N_43697,N_42384,N_42037);
and U43698 (N_43698,N_41504,N_41679);
xnor U43699 (N_43699,N_41362,N_41710);
nor U43700 (N_43700,N_41088,N_40629);
nor U43701 (N_43701,N_41741,N_40495);
or U43702 (N_43702,N_41691,N_40911);
nand U43703 (N_43703,N_40868,N_40284);
or U43704 (N_43704,N_41271,N_41463);
and U43705 (N_43705,N_40124,N_40410);
or U43706 (N_43706,N_40887,N_41135);
or U43707 (N_43707,N_40362,N_40873);
and U43708 (N_43708,N_42357,N_42283);
and U43709 (N_43709,N_42206,N_41075);
nand U43710 (N_43710,N_41736,N_41118);
nor U43711 (N_43711,N_40405,N_41685);
and U43712 (N_43712,N_41081,N_41879);
and U43713 (N_43713,N_42012,N_40691);
or U43714 (N_43714,N_41554,N_41409);
and U43715 (N_43715,N_41648,N_41008);
or U43716 (N_43716,N_40451,N_41651);
or U43717 (N_43717,N_41226,N_40753);
xnor U43718 (N_43718,N_41460,N_42067);
and U43719 (N_43719,N_40278,N_40413);
nand U43720 (N_43720,N_41611,N_40754);
or U43721 (N_43721,N_40896,N_40354);
or U43722 (N_43722,N_40561,N_41590);
xor U43723 (N_43723,N_40096,N_42383);
xor U43724 (N_43724,N_41483,N_41994);
or U43725 (N_43725,N_41205,N_40102);
or U43726 (N_43726,N_40843,N_40094);
nor U43727 (N_43727,N_41798,N_42204);
xnor U43728 (N_43728,N_40530,N_41146);
nand U43729 (N_43729,N_42173,N_41243);
xnor U43730 (N_43730,N_42259,N_40029);
xor U43731 (N_43731,N_41629,N_40572);
and U43732 (N_43732,N_41415,N_40587);
and U43733 (N_43733,N_41768,N_41717);
nand U43734 (N_43734,N_42456,N_41649);
and U43735 (N_43735,N_40172,N_40517);
and U43736 (N_43736,N_40266,N_41423);
and U43737 (N_43737,N_41063,N_41746);
xor U43738 (N_43738,N_41638,N_41110);
nand U43739 (N_43739,N_41069,N_40784);
nor U43740 (N_43740,N_41230,N_40650);
and U43741 (N_43741,N_41193,N_42091);
nor U43742 (N_43742,N_40930,N_40338);
or U43743 (N_43743,N_40228,N_41398);
nand U43744 (N_43744,N_40966,N_41868);
nand U43745 (N_43745,N_41761,N_41909);
or U43746 (N_43746,N_40481,N_42171);
and U43747 (N_43747,N_40902,N_42000);
and U43748 (N_43748,N_41708,N_40205);
nor U43749 (N_43749,N_40942,N_41977);
nor U43750 (N_43750,N_40883,N_40296);
and U43751 (N_43751,N_42143,N_40960);
xor U43752 (N_43752,N_41763,N_41244);
xor U43753 (N_43753,N_41956,N_41556);
nand U43754 (N_43754,N_40695,N_42108);
nor U43755 (N_43755,N_42479,N_40812);
nand U43756 (N_43756,N_40519,N_42381);
and U43757 (N_43757,N_41097,N_40135);
nand U43758 (N_43758,N_41841,N_42493);
xor U43759 (N_43759,N_41864,N_41280);
nand U43760 (N_43760,N_42112,N_40059);
nor U43761 (N_43761,N_42146,N_40380);
xnor U43762 (N_43762,N_42047,N_40134);
xnor U43763 (N_43763,N_40119,N_41424);
nor U43764 (N_43764,N_42278,N_40294);
nand U43765 (N_43765,N_41254,N_41475);
xor U43766 (N_43766,N_41998,N_41794);
or U43767 (N_43767,N_40657,N_41469);
nor U43768 (N_43768,N_40446,N_41859);
nand U43769 (N_43769,N_41299,N_41416);
or U43770 (N_43770,N_42025,N_41050);
and U43771 (N_43771,N_40399,N_42108);
xor U43772 (N_43772,N_40616,N_40439);
xnor U43773 (N_43773,N_42217,N_42038);
and U43774 (N_43774,N_42403,N_41438);
nand U43775 (N_43775,N_41713,N_41088);
xor U43776 (N_43776,N_40349,N_41868);
nor U43777 (N_43777,N_41309,N_41522);
or U43778 (N_43778,N_41755,N_42272);
and U43779 (N_43779,N_41732,N_41899);
nand U43780 (N_43780,N_41542,N_42150);
nand U43781 (N_43781,N_41844,N_41910);
and U43782 (N_43782,N_40535,N_42240);
or U43783 (N_43783,N_41215,N_41604);
and U43784 (N_43784,N_41448,N_42465);
nand U43785 (N_43785,N_41458,N_41652);
xnor U43786 (N_43786,N_41230,N_40005);
nor U43787 (N_43787,N_40099,N_40772);
nand U43788 (N_43788,N_40755,N_40039);
nand U43789 (N_43789,N_40553,N_42398);
or U43790 (N_43790,N_41789,N_42241);
xnor U43791 (N_43791,N_41666,N_42263);
and U43792 (N_43792,N_40112,N_41688);
xnor U43793 (N_43793,N_40393,N_41199);
or U43794 (N_43794,N_40932,N_41462);
nand U43795 (N_43795,N_41788,N_40240);
xnor U43796 (N_43796,N_40567,N_40326);
nor U43797 (N_43797,N_41049,N_41333);
and U43798 (N_43798,N_40300,N_40726);
or U43799 (N_43799,N_40062,N_42225);
and U43800 (N_43800,N_41750,N_41790);
and U43801 (N_43801,N_41694,N_42072);
nor U43802 (N_43802,N_42155,N_41226);
and U43803 (N_43803,N_42382,N_42107);
nand U43804 (N_43804,N_41012,N_40922);
and U43805 (N_43805,N_42126,N_41534);
or U43806 (N_43806,N_41614,N_42482);
or U43807 (N_43807,N_40398,N_42270);
nor U43808 (N_43808,N_40466,N_42235);
or U43809 (N_43809,N_40742,N_42423);
nor U43810 (N_43810,N_41756,N_41289);
xor U43811 (N_43811,N_42131,N_42007);
xor U43812 (N_43812,N_42217,N_41013);
and U43813 (N_43813,N_40331,N_41037);
xor U43814 (N_43814,N_40367,N_41044);
and U43815 (N_43815,N_42432,N_41191);
nand U43816 (N_43816,N_40427,N_40889);
nor U43817 (N_43817,N_41556,N_40344);
nand U43818 (N_43818,N_41694,N_41131);
nand U43819 (N_43819,N_42198,N_40171);
xor U43820 (N_43820,N_42262,N_40450);
nand U43821 (N_43821,N_40454,N_42023);
xor U43822 (N_43822,N_42443,N_40288);
nor U43823 (N_43823,N_40352,N_41567);
and U43824 (N_43824,N_41532,N_40363);
and U43825 (N_43825,N_40458,N_42390);
or U43826 (N_43826,N_42363,N_41887);
nor U43827 (N_43827,N_40372,N_42112);
xnor U43828 (N_43828,N_42210,N_41527);
or U43829 (N_43829,N_42133,N_42437);
or U43830 (N_43830,N_42180,N_42038);
and U43831 (N_43831,N_41985,N_41814);
and U43832 (N_43832,N_41790,N_40366);
and U43833 (N_43833,N_41953,N_41802);
and U43834 (N_43834,N_40130,N_40283);
and U43835 (N_43835,N_40678,N_41090);
nor U43836 (N_43836,N_40650,N_40865);
xnor U43837 (N_43837,N_41617,N_42278);
xor U43838 (N_43838,N_40694,N_40917);
xnor U43839 (N_43839,N_41146,N_42148);
and U43840 (N_43840,N_41006,N_41484);
xor U43841 (N_43841,N_40847,N_41280);
or U43842 (N_43842,N_42033,N_41440);
or U43843 (N_43843,N_40281,N_42413);
nand U43844 (N_43844,N_40568,N_41330);
nor U43845 (N_43845,N_40840,N_41202);
and U43846 (N_43846,N_42413,N_42301);
nand U43847 (N_43847,N_40468,N_42253);
or U43848 (N_43848,N_40283,N_40934);
or U43849 (N_43849,N_40556,N_41191);
xor U43850 (N_43850,N_41121,N_40563);
nand U43851 (N_43851,N_41244,N_40262);
nor U43852 (N_43852,N_41526,N_40344);
or U43853 (N_43853,N_42004,N_41691);
nand U43854 (N_43854,N_40567,N_42024);
nor U43855 (N_43855,N_41986,N_42494);
and U43856 (N_43856,N_40307,N_41675);
or U43857 (N_43857,N_41195,N_42108);
or U43858 (N_43858,N_42495,N_42130);
or U43859 (N_43859,N_41527,N_40968);
nor U43860 (N_43860,N_41355,N_42370);
and U43861 (N_43861,N_40702,N_41721);
xnor U43862 (N_43862,N_40172,N_41111);
or U43863 (N_43863,N_40357,N_40095);
and U43864 (N_43864,N_40571,N_42050);
nor U43865 (N_43865,N_41978,N_42283);
xnor U43866 (N_43866,N_40576,N_41370);
and U43867 (N_43867,N_42409,N_41048);
nor U43868 (N_43868,N_41868,N_41744);
nor U43869 (N_43869,N_40137,N_40993);
and U43870 (N_43870,N_41357,N_41168);
nor U43871 (N_43871,N_40476,N_40184);
xor U43872 (N_43872,N_42072,N_40206);
nand U43873 (N_43873,N_41355,N_41183);
and U43874 (N_43874,N_40236,N_41722);
nor U43875 (N_43875,N_41825,N_40743);
nor U43876 (N_43876,N_41627,N_41259);
nand U43877 (N_43877,N_42237,N_40982);
and U43878 (N_43878,N_41997,N_40607);
xnor U43879 (N_43879,N_41715,N_40247);
nor U43880 (N_43880,N_40088,N_40056);
or U43881 (N_43881,N_41875,N_40225);
or U43882 (N_43882,N_42084,N_40472);
nand U43883 (N_43883,N_42481,N_40621);
nor U43884 (N_43884,N_40187,N_40429);
xor U43885 (N_43885,N_42306,N_41463);
and U43886 (N_43886,N_41548,N_40397);
and U43887 (N_43887,N_40934,N_40277);
nor U43888 (N_43888,N_41874,N_40769);
nor U43889 (N_43889,N_40562,N_41994);
or U43890 (N_43890,N_40578,N_41102);
or U43891 (N_43891,N_41587,N_41777);
or U43892 (N_43892,N_40172,N_42217);
or U43893 (N_43893,N_41330,N_41774);
nor U43894 (N_43894,N_42201,N_40162);
nand U43895 (N_43895,N_41394,N_42069);
or U43896 (N_43896,N_40902,N_40453);
nand U43897 (N_43897,N_41882,N_41158);
xnor U43898 (N_43898,N_40874,N_40563);
or U43899 (N_43899,N_41108,N_40280);
nor U43900 (N_43900,N_41593,N_41409);
nor U43901 (N_43901,N_40674,N_41353);
nand U43902 (N_43902,N_41031,N_42472);
or U43903 (N_43903,N_41929,N_41115);
xnor U43904 (N_43904,N_41125,N_41571);
nor U43905 (N_43905,N_40336,N_41980);
xnor U43906 (N_43906,N_41424,N_42145);
xor U43907 (N_43907,N_42160,N_40855);
nor U43908 (N_43908,N_41624,N_40094);
or U43909 (N_43909,N_41726,N_41715);
and U43910 (N_43910,N_40504,N_42148);
nand U43911 (N_43911,N_40529,N_42467);
nor U43912 (N_43912,N_40300,N_40747);
nor U43913 (N_43913,N_41185,N_40280);
nand U43914 (N_43914,N_41635,N_41847);
and U43915 (N_43915,N_40425,N_41289);
xor U43916 (N_43916,N_40152,N_40535);
and U43917 (N_43917,N_42194,N_42393);
nand U43918 (N_43918,N_41479,N_42211);
xnor U43919 (N_43919,N_41991,N_42419);
xnor U43920 (N_43920,N_41628,N_40635);
nand U43921 (N_43921,N_41578,N_42436);
nand U43922 (N_43922,N_41016,N_41278);
nand U43923 (N_43923,N_40897,N_40454);
and U43924 (N_43924,N_41096,N_40422);
or U43925 (N_43925,N_42132,N_40080);
xnor U43926 (N_43926,N_40238,N_40682);
nor U43927 (N_43927,N_41835,N_42028);
or U43928 (N_43928,N_42128,N_41976);
nand U43929 (N_43929,N_41164,N_41875);
nand U43930 (N_43930,N_41043,N_40300);
nand U43931 (N_43931,N_41371,N_42289);
or U43932 (N_43932,N_40861,N_41379);
xor U43933 (N_43933,N_40174,N_41708);
xor U43934 (N_43934,N_40583,N_41410);
and U43935 (N_43935,N_41723,N_40737);
xnor U43936 (N_43936,N_42215,N_41964);
nor U43937 (N_43937,N_42396,N_41552);
nor U43938 (N_43938,N_40651,N_40020);
or U43939 (N_43939,N_42273,N_41484);
xnor U43940 (N_43940,N_40380,N_40881);
nor U43941 (N_43941,N_41821,N_42144);
and U43942 (N_43942,N_40503,N_41574);
nor U43943 (N_43943,N_42163,N_42389);
and U43944 (N_43944,N_40664,N_40129);
nor U43945 (N_43945,N_41488,N_40938);
nor U43946 (N_43946,N_40990,N_42363);
nor U43947 (N_43947,N_40046,N_41931);
nand U43948 (N_43948,N_42371,N_40989);
or U43949 (N_43949,N_40727,N_40851);
and U43950 (N_43950,N_42357,N_40386);
nor U43951 (N_43951,N_40821,N_41721);
and U43952 (N_43952,N_41952,N_41524);
xor U43953 (N_43953,N_42458,N_41584);
or U43954 (N_43954,N_40865,N_41275);
xnor U43955 (N_43955,N_41574,N_41957);
nand U43956 (N_43956,N_41681,N_42030);
or U43957 (N_43957,N_41301,N_42223);
and U43958 (N_43958,N_41606,N_41557);
and U43959 (N_43959,N_42429,N_40503);
xnor U43960 (N_43960,N_40085,N_41783);
nand U43961 (N_43961,N_42383,N_41362);
nor U43962 (N_43962,N_42458,N_40965);
nor U43963 (N_43963,N_41157,N_41286);
nor U43964 (N_43964,N_41207,N_42109);
and U43965 (N_43965,N_40293,N_40973);
xnor U43966 (N_43966,N_40147,N_40257);
nor U43967 (N_43967,N_42138,N_40226);
and U43968 (N_43968,N_41011,N_41384);
nor U43969 (N_43969,N_40436,N_41477);
nand U43970 (N_43970,N_40211,N_42416);
xor U43971 (N_43971,N_42022,N_41732);
nand U43972 (N_43972,N_40490,N_42386);
nor U43973 (N_43973,N_40923,N_40516);
xnor U43974 (N_43974,N_40825,N_42249);
and U43975 (N_43975,N_40446,N_41869);
and U43976 (N_43976,N_40619,N_41130);
or U43977 (N_43977,N_40931,N_40733);
nand U43978 (N_43978,N_41565,N_41163);
nand U43979 (N_43979,N_40552,N_41812);
or U43980 (N_43980,N_42381,N_40438);
and U43981 (N_43981,N_40480,N_41208);
nor U43982 (N_43982,N_40461,N_40416);
and U43983 (N_43983,N_40115,N_40570);
and U43984 (N_43984,N_40596,N_40578);
and U43985 (N_43985,N_41582,N_42374);
nor U43986 (N_43986,N_41022,N_42097);
or U43987 (N_43987,N_40220,N_40152);
xor U43988 (N_43988,N_40233,N_40148);
nor U43989 (N_43989,N_40324,N_41418);
and U43990 (N_43990,N_40244,N_42470);
nor U43991 (N_43991,N_41772,N_41137);
nand U43992 (N_43992,N_41240,N_41718);
nand U43993 (N_43993,N_40749,N_41348);
nand U43994 (N_43994,N_40794,N_41434);
or U43995 (N_43995,N_41183,N_40948);
nand U43996 (N_43996,N_42493,N_40467);
nand U43997 (N_43997,N_42346,N_40430);
or U43998 (N_43998,N_41052,N_41731);
or U43999 (N_43999,N_40375,N_40755);
or U44000 (N_44000,N_40359,N_41273);
nand U44001 (N_44001,N_42038,N_40179);
and U44002 (N_44002,N_40866,N_41349);
or U44003 (N_44003,N_41158,N_41008);
and U44004 (N_44004,N_40327,N_40617);
and U44005 (N_44005,N_40911,N_41831);
nor U44006 (N_44006,N_41599,N_41763);
and U44007 (N_44007,N_41860,N_40578);
nor U44008 (N_44008,N_40940,N_42094);
xor U44009 (N_44009,N_42390,N_41405);
and U44010 (N_44010,N_40831,N_42387);
nor U44011 (N_44011,N_41498,N_40906);
or U44012 (N_44012,N_42295,N_40369);
or U44013 (N_44013,N_42461,N_41483);
nand U44014 (N_44014,N_42322,N_40383);
and U44015 (N_44015,N_40166,N_41083);
nand U44016 (N_44016,N_42045,N_42048);
nand U44017 (N_44017,N_40484,N_42062);
and U44018 (N_44018,N_41779,N_40173);
nand U44019 (N_44019,N_40569,N_41641);
xnor U44020 (N_44020,N_40598,N_40939);
and U44021 (N_44021,N_40008,N_40063);
nand U44022 (N_44022,N_41052,N_41793);
or U44023 (N_44023,N_41636,N_41782);
nor U44024 (N_44024,N_41282,N_40279);
nor U44025 (N_44025,N_41240,N_41129);
xor U44026 (N_44026,N_42133,N_42294);
xor U44027 (N_44027,N_41547,N_41533);
and U44028 (N_44028,N_40090,N_42408);
or U44029 (N_44029,N_41270,N_40129);
and U44030 (N_44030,N_40119,N_41485);
nor U44031 (N_44031,N_41090,N_41122);
and U44032 (N_44032,N_41908,N_41927);
and U44033 (N_44033,N_42274,N_40081);
nor U44034 (N_44034,N_42119,N_41542);
nor U44035 (N_44035,N_41313,N_41872);
and U44036 (N_44036,N_41997,N_41125);
and U44037 (N_44037,N_40725,N_40051);
nand U44038 (N_44038,N_41383,N_41248);
or U44039 (N_44039,N_42251,N_40810);
nor U44040 (N_44040,N_42126,N_42057);
and U44041 (N_44041,N_40775,N_40528);
and U44042 (N_44042,N_41460,N_42010);
and U44043 (N_44043,N_40278,N_40914);
nand U44044 (N_44044,N_40549,N_41535);
nand U44045 (N_44045,N_41664,N_42302);
and U44046 (N_44046,N_40697,N_41742);
or U44047 (N_44047,N_40462,N_41037);
xnor U44048 (N_44048,N_40986,N_42339);
and U44049 (N_44049,N_41476,N_41785);
nand U44050 (N_44050,N_41052,N_40973);
nor U44051 (N_44051,N_42068,N_40444);
xor U44052 (N_44052,N_40175,N_40041);
nor U44053 (N_44053,N_41396,N_41107);
and U44054 (N_44054,N_40102,N_42043);
nor U44055 (N_44055,N_41788,N_41917);
or U44056 (N_44056,N_41254,N_42295);
or U44057 (N_44057,N_41684,N_41501);
or U44058 (N_44058,N_42068,N_42299);
xor U44059 (N_44059,N_41279,N_40403);
and U44060 (N_44060,N_40268,N_41008);
nor U44061 (N_44061,N_41013,N_40726);
and U44062 (N_44062,N_41030,N_40996);
xor U44063 (N_44063,N_42107,N_41423);
nand U44064 (N_44064,N_40348,N_41237);
nor U44065 (N_44065,N_41754,N_42237);
and U44066 (N_44066,N_40928,N_41691);
or U44067 (N_44067,N_42316,N_41409);
or U44068 (N_44068,N_41335,N_41138);
nand U44069 (N_44069,N_40330,N_40489);
or U44070 (N_44070,N_40777,N_41177);
or U44071 (N_44071,N_40727,N_41579);
xnor U44072 (N_44072,N_41729,N_42231);
nand U44073 (N_44073,N_40580,N_42196);
and U44074 (N_44074,N_41743,N_40573);
nor U44075 (N_44075,N_41755,N_41421);
nand U44076 (N_44076,N_40438,N_42090);
nor U44077 (N_44077,N_41473,N_40830);
nand U44078 (N_44078,N_40517,N_42330);
nand U44079 (N_44079,N_41962,N_41988);
nor U44080 (N_44080,N_41112,N_40350);
nand U44081 (N_44081,N_41299,N_40772);
nand U44082 (N_44082,N_42019,N_41451);
and U44083 (N_44083,N_40254,N_42195);
nor U44084 (N_44084,N_40373,N_40512);
or U44085 (N_44085,N_40501,N_41681);
xnor U44086 (N_44086,N_40050,N_40762);
or U44087 (N_44087,N_41431,N_41518);
nand U44088 (N_44088,N_41159,N_40617);
xnor U44089 (N_44089,N_40092,N_41846);
and U44090 (N_44090,N_41166,N_40811);
and U44091 (N_44091,N_41972,N_42334);
or U44092 (N_44092,N_40965,N_40154);
xor U44093 (N_44093,N_41881,N_42305);
nor U44094 (N_44094,N_41781,N_41897);
xor U44095 (N_44095,N_40432,N_42076);
and U44096 (N_44096,N_42153,N_40498);
or U44097 (N_44097,N_42211,N_40111);
nand U44098 (N_44098,N_41563,N_40063);
xnor U44099 (N_44099,N_40039,N_40863);
nor U44100 (N_44100,N_40677,N_41249);
and U44101 (N_44101,N_42297,N_41322);
or U44102 (N_44102,N_40024,N_42128);
xnor U44103 (N_44103,N_40514,N_40004);
nor U44104 (N_44104,N_40141,N_40908);
nand U44105 (N_44105,N_40246,N_41605);
xnor U44106 (N_44106,N_40229,N_42335);
or U44107 (N_44107,N_40649,N_41326);
and U44108 (N_44108,N_41981,N_41747);
nand U44109 (N_44109,N_40595,N_40429);
or U44110 (N_44110,N_41312,N_42235);
nand U44111 (N_44111,N_40062,N_41176);
nand U44112 (N_44112,N_41233,N_40790);
and U44113 (N_44113,N_40664,N_40985);
or U44114 (N_44114,N_42185,N_40902);
nand U44115 (N_44115,N_40014,N_40753);
or U44116 (N_44116,N_40922,N_40576);
xor U44117 (N_44117,N_40248,N_41309);
and U44118 (N_44118,N_41013,N_40860);
or U44119 (N_44119,N_41495,N_41708);
nand U44120 (N_44120,N_40890,N_40856);
or U44121 (N_44121,N_40585,N_41148);
and U44122 (N_44122,N_41428,N_42223);
and U44123 (N_44123,N_42333,N_40944);
nor U44124 (N_44124,N_40495,N_41832);
xnor U44125 (N_44125,N_40444,N_41100);
nand U44126 (N_44126,N_41142,N_42099);
and U44127 (N_44127,N_41699,N_40035);
and U44128 (N_44128,N_41581,N_42152);
or U44129 (N_44129,N_41250,N_41540);
nand U44130 (N_44130,N_40673,N_40829);
or U44131 (N_44131,N_40530,N_40739);
nand U44132 (N_44132,N_41699,N_40969);
nor U44133 (N_44133,N_41441,N_42220);
and U44134 (N_44134,N_42394,N_40559);
nand U44135 (N_44135,N_40538,N_41460);
or U44136 (N_44136,N_41762,N_40280);
and U44137 (N_44137,N_40744,N_41009);
and U44138 (N_44138,N_41468,N_41246);
or U44139 (N_44139,N_40180,N_41440);
nand U44140 (N_44140,N_41115,N_42344);
nand U44141 (N_44141,N_41330,N_41862);
and U44142 (N_44142,N_40983,N_41125);
nand U44143 (N_44143,N_41530,N_41508);
nand U44144 (N_44144,N_40159,N_40441);
or U44145 (N_44145,N_41869,N_41250);
xor U44146 (N_44146,N_40415,N_41865);
nand U44147 (N_44147,N_40153,N_41135);
and U44148 (N_44148,N_42231,N_40141);
xnor U44149 (N_44149,N_40929,N_42008);
nor U44150 (N_44150,N_42307,N_41958);
nor U44151 (N_44151,N_42187,N_40606);
and U44152 (N_44152,N_42137,N_41518);
nor U44153 (N_44153,N_41986,N_40348);
xor U44154 (N_44154,N_40284,N_41049);
and U44155 (N_44155,N_40438,N_40406);
or U44156 (N_44156,N_40671,N_40386);
xnor U44157 (N_44157,N_42208,N_41827);
and U44158 (N_44158,N_40256,N_42022);
xor U44159 (N_44159,N_41507,N_41639);
xor U44160 (N_44160,N_40117,N_40965);
nor U44161 (N_44161,N_41927,N_40094);
or U44162 (N_44162,N_42153,N_42436);
nor U44163 (N_44163,N_41130,N_41000);
nor U44164 (N_44164,N_41309,N_40235);
nor U44165 (N_44165,N_41091,N_41524);
or U44166 (N_44166,N_40047,N_40844);
nor U44167 (N_44167,N_42400,N_41728);
or U44168 (N_44168,N_42112,N_41488);
nor U44169 (N_44169,N_42094,N_40062);
and U44170 (N_44170,N_40785,N_40515);
or U44171 (N_44171,N_40537,N_42119);
or U44172 (N_44172,N_40796,N_40754);
nand U44173 (N_44173,N_41827,N_41414);
or U44174 (N_44174,N_40953,N_42296);
and U44175 (N_44175,N_41947,N_41342);
nor U44176 (N_44176,N_41325,N_42215);
nor U44177 (N_44177,N_42223,N_40709);
xor U44178 (N_44178,N_41596,N_41976);
or U44179 (N_44179,N_41595,N_40358);
or U44180 (N_44180,N_40973,N_41312);
and U44181 (N_44181,N_40274,N_40115);
xnor U44182 (N_44182,N_42174,N_40647);
nor U44183 (N_44183,N_40101,N_42214);
nand U44184 (N_44184,N_42445,N_40230);
nand U44185 (N_44185,N_41428,N_41529);
nor U44186 (N_44186,N_42370,N_40269);
or U44187 (N_44187,N_40475,N_40994);
or U44188 (N_44188,N_41729,N_41765);
nor U44189 (N_44189,N_40615,N_41572);
and U44190 (N_44190,N_41761,N_41882);
nand U44191 (N_44191,N_40429,N_41548);
nor U44192 (N_44192,N_41173,N_42465);
nand U44193 (N_44193,N_41073,N_40964);
and U44194 (N_44194,N_41958,N_40198);
nand U44195 (N_44195,N_41816,N_41128);
and U44196 (N_44196,N_40625,N_41772);
nor U44197 (N_44197,N_41402,N_41849);
or U44198 (N_44198,N_40281,N_41916);
nor U44199 (N_44199,N_41298,N_42354);
xnor U44200 (N_44200,N_40414,N_41940);
nand U44201 (N_44201,N_40945,N_41846);
and U44202 (N_44202,N_40772,N_40147);
xnor U44203 (N_44203,N_41622,N_41124);
nor U44204 (N_44204,N_40388,N_40091);
or U44205 (N_44205,N_41901,N_41588);
or U44206 (N_44206,N_42173,N_40500);
nor U44207 (N_44207,N_42044,N_41040);
nor U44208 (N_44208,N_40108,N_42478);
nand U44209 (N_44209,N_42257,N_40854);
xnor U44210 (N_44210,N_41759,N_41835);
and U44211 (N_44211,N_40159,N_42452);
nor U44212 (N_44212,N_40116,N_42494);
nor U44213 (N_44213,N_41936,N_40715);
xor U44214 (N_44214,N_42451,N_41294);
nand U44215 (N_44215,N_41136,N_40333);
nor U44216 (N_44216,N_42206,N_41222);
xnor U44217 (N_44217,N_40821,N_41356);
nor U44218 (N_44218,N_42498,N_40446);
xnor U44219 (N_44219,N_41478,N_42176);
nand U44220 (N_44220,N_42250,N_40036);
and U44221 (N_44221,N_41092,N_40395);
and U44222 (N_44222,N_41507,N_41431);
and U44223 (N_44223,N_42214,N_40471);
and U44224 (N_44224,N_40502,N_41162);
nand U44225 (N_44225,N_41209,N_41261);
and U44226 (N_44226,N_40550,N_40472);
nor U44227 (N_44227,N_42001,N_41437);
and U44228 (N_44228,N_41368,N_40296);
xor U44229 (N_44229,N_40580,N_42001);
nand U44230 (N_44230,N_40515,N_40941);
and U44231 (N_44231,N_42498,N_40490);
and U44232 (N_44232,N_40554,N_40828);
xor U44233 (N_44233,N_40334,N_40193);
and U44234 (N_44234,N_40034,N_41836);
nor U44235 (N_44235,N_42029,N_41900);
or U44236 (N_44236,N_41293,N_40148);
xnor U44237 (N_44237,N_41375,N_42186);
and U44238 (N_44238,N_40967,N_40507);
nor U44239 (N_44239,N_41524,N_40138);
nor U44240 (N_44240,N_42186,N_40529);
nor U44241 (N_44241,N_41815,N_40811);
nand U44242 (N_44242,N_40709,N_42455);
nand U44243 (N_44243,N_40003,N_40212);
nor U44244 (N_44244,N_40597,N_40003);
and U44245 (N_44245,N_42480,N_42157);
xnor U44246 (N_44246,N_41899,N_40519);
and U44247 (N_44247,N_40683,N_40633);
nand U44248 (N_44248,N_40932,N_41638);
or U44249 (N_44249,N_41465,N_40995);
nand U44250 (N_44250,N_41115,N_41831);
xor U44251 (N_44251,N_40981,N_42162);
xnor U44252 (N_44252,N_40746,N_40271);
or U44253 (N_44253,N_42010,N_41159);
and U44254 (N_44254,N_40230,N_40251);
or U44255 (N_44255,N_40303,N_41093);
and U44256 (N_44256,N_41378,N_40925);
or U44257 (N_44257,N_42108,N_41263);
and U44258 (N_44258,N_40750,N_41787);
xnor U44259 (N_44259,N_41384,N_42434);
nor U44260 (N_44260,N_41901,N_41544);
nor U44261 (N_44261,N_41829,N_42297);
nand U44262 (N_44262,N_41225,N_40332);
nor U44263 (N_44263,N_41023,N_40187);
or U44264 (N_44264,N_41012,N_40913);
xor U44265 (N_44265,N_40487,N_40561);
nor U44266 (N_44266,N_41938,N_40786);
nor U44267 (N_44267,N_40770,N_40828);
or U44268 (N_44268,N_41357,N_40906);
xnor U44269 (N_44269,N_40189,N_40345);
nor U44270 (N_44270,N_41854,N_41791);
nor U44271 (N_44271,N_42412,N_40432);
or U44272 (N_44272,N_41599,N_40569);
xor U44273 (N_44273,N_41671,N_42055);
nand U44274 (N_44274,N_41380,N_40498);
and U44275 (N_44275,N_40243,N_42267);
or U44276 (N_44276,N_40563,N_40763);
nand U44277 (N_44277,N_40974,N_42142);
and U44278 (N_44278,N_40007,N_41805);
nor U44279 (N_44279,N_41669,N_42065);
or U44280 (N_44280,N_40391,N_42155);
and U44281 (N_44281,N_40921,N_42053);
xor U44282 (N_44282,N_41690,N_42398);
and U44283 (N_44283,N_40827,N_42139);
nor U44284 (N_44284,N_41749,N_40181);
and U44285 (N_44285,N_40572,N_41544);
or U44286 (N_44286,N_40129,N_41406);
nor U44287 (N_44287,N_40313,N_40211);
or U44288 (N_44288,N_41027,N_41897);
nand U44289 (N_44289,N_42345,N_40075);
and U44290 (N_44290,N_42023,N_41383);
nor U44291 (N_44291,N_41819,N_42315);
nor U44292 (N_44292,N_41649,N_41400);
or U44293 (N_44293,N_42244,N_40800);
or U44294 (N_44294,N_41577,N_42471);
nor U44295 (N_44295,N_41987,N_40485);
nand U44296 (N_44296,N_40563,N_41610);
nand U44297 (N_44297,N_41270,N_40362);
or U44298 (N_44298,N_40492,N_41227);
nand U44299 (N_44299,N_40655,N_40760);
or U44300 (N_44300,N_42301,N_40566);
or U44301 (N_44301,N_41028,N_42321);
or U44302 (N_44302,N_42242,N_40499);
or U44303 (N_44303,N_42216,N_42090);
xnor U44304 (N_44304,N_42210,N_41732);
nor U44305 (N_44305,N_40778,N_40094);
or U44306 (N_44306,N_40360,N_41465);
nor U44307 (N_44307,N_42180,N_41762);
xnor U44308 (N_44308,N_42347,N_42402);
nand U44309 (N_44309,N_41538,N_40094);
or U44310 (N_44310,N_40293,N_42402);
or U44311 (N_44311,N_41363,N_41030);
or U44312 (N_44312,N_42381,N_40174);
nor U44313 (N_44313,N_41598,N_40936);
nor U44314 (N_44314,N_40597,N_42374);
or U44315 (N_44315,N_40862,N_41465);
xor U44316 (N_44316,N_42101,N_40397);
or U44317 (N_44317,N_41058,N_41452);
nand U44318 (N_44318,N_42164,N_41411);
nor U44319 (N_44319,N_42164,N_41805);
nor U44320 (N_44320,N_40490,N_42163);
xnor U44321 (N_44321,N_41844,N_40920);
or U44322 (N_44322,N_40312,N_41177);
nor U44323 (N_44323,N_40882,N_40225);
nor U44324 (N_44324,N_40176,N_42290);
or U44325 (N_44325,N_41539,N_41609);
xnor U44326 (N_44326,N_40432,N_41412);
nor U44327 (N_44327,N_41404,N_40849);
or U44328 (N_44328,N_40602,N_41146);
nor U44329 (N_44329,N_42459,N_42022);
nor U44330 (N_44330,N_40337,N_41919);
or U44331 (N_44331,N_40575,N_40867);
xnor U44332 (N_44332,N_41557,N_41046);
xnor U44333 (N_44333,N_42392,N_40477);
or U44334 (N_44334,N_40172,N_42330);
or U44335 (N_44335,N_40775,N_41713);
and U44336 (N_44336,N_41884,N_41505);
nand U44337 (N_44337,N_41259,N_40100);
or U44338 (N_44338,N_42432,N_42246);
nor U44339 (N_44339,N_41959,N_42328);
xnor U44340 (N_44340,N_40040,N_41739);
or U44341 (N_44341,N_41821,N_41028);
xor U44342 (N_44342,N_42356,N_42104);
and U44343 (N_44343,N_41159,N_41113);
xor U44344 (N_44344,N_42175,N_41323);
and U44345 (N_44345,N_41394,N_42376);
xor U44346 (N_44346,N_40454,N_41684);
and U44347 (N_44347,N_40215,N_42382);
nor U44348 (N_44348,N_42087,N_40135);
or U44349 (N_44349,N_40089,N_42332);
nand U44350 (N_44350,N_40328,N_40061);
nand U44351 (N_44351,N_41470,N_41792);
or U44352 (N_44352,N_41965,N_41395);
or U44353 (N_44353,N_40664,N_41392);
nand U44354 (N_44354,N_42381,N_40405);
or U44355 (N_44355,N_41951,N_41646);
and U44356 (N_44356,N_42005,N_40667);
xor U44357 (N_44357,N_41081,N_41472);
nor U44358 (N_44358,N_42477,N_41496);
nand U44359 (N_44359,N_40170,N_42329);
and U44360 (N_44360,N_41790,N_42489);
or U44361 (N_44361,N_40705,N_40783);
xnor U44362 (N_44362,N_40786,N_42327);
or U44363 (N_44363,N_40966,N_42303);
xor U44364 (N_44364,N_42127,N_40785);
and U44365 (N_44365,N_42320,N_42224);
or U44366 (N_44366,N_41036,N_41338);
xor U44367 (N_44367,N_42312,N_41332);
or U44368 (N_44368,N_40859,N_41528);
nand U44369 (N_44369,N_40314,N_40154);
and U44370 (N_44370,N_40830,N_41185);
xnor U44371 (N_44371,N_40741,N_40237);
or U44372 (N_44372,N_41460,N_41040);
xnor U44373 (N_44373,N_41916,N_40988);
or U44374 (N_44374,N_42334,N_42441);
and U44375 (N_44375,N_41955,N_42373);
xor U44376 (N_44376,N_40956,N_41750);
and U44377 (N_44377,N_41410,N_42054);
and U44378 (N_44378,N_40418,N_41421);
xnor U44379 (N_44379,N_40821,N_40942);
nand U44380 (N_44380,N_40446,N_41427);
or U44381 (N_44381,N_42474,N_40518);
or U44382 (N_44382,N_41025,N_40679);
and U44383 (N_44383,N_40787,N_42246);
and U44384 (N_44384,N_41291,N_40849);
and U44385 (N_44385,N_41297,N_41631);
and U44386 (N_44386,N_40578,N_41398);
or U44387 (N_44387,N_40044,N_40280);
nor U44388 (N_44388,N_41425,N_41038);
or U44389 (N_44389,N_41844,N_40008);
and U44390 (N_44390,N_41062,N_41998);
nand U44391 (N_44391,N_42012,N_40776);
xor U44392 (N_44392,N_41633,N_40377);
and U44393 (N_44393,N_40327,N_42454);
nor U44394 (N_44394,N_41170,N_41488);
or U44395 (N_44395,N_42403,N_40105);
nand U44396 (N_44396,N_40797,N_41423);
or U44397 (N_44397,N_40406,N_40550);
nor U44398 (N_44398,N_41365,N_42006);
or U44399 (N_44399,N_42066,N_40727);
and U44400 (N_44400,N_40911,N_40490);
nand U44401 (N_44401,N_40927,N_40480);
xnor U44402 (N_44402,N_41074,N_41356);
and U44403 (N_44403,N_42004,N_40518);
and U44404 (N_44404,N_40057,N_40777);
xnor U44405 (N_44405,N_40334,N_40431);
and U44406 (N_44406,N_41543,N_40199);
nor U44407 (N_44407,N_42138,N_40297);
and U44408 (N_44408,N_41720,N_40269);
xnor U44409 (N_44409,N_41667,N_42247);
and U44410 (N_44410,N_42104,N_40207);
nor U44411 (N_44411,N_41724,N_41227);
xnor U44412 (N_44412,N_41407,N_41919);
nor U44413 (N_44413,N_40648,N_42209);
xor U44414 (N_44414,N_41709,N_40849);
nor U44415 (N_44415,N_41359,N_42286);
or U44416 (N_44416,N_40803,N_40312);
nor U44417 (N_44417,N_40138,N_41218);
or U44418 (N_44418,N_41395,N_40645);
xor U44419 (N_44419,N_42215,N_40711);
or U44420 (N_44420,N_41679,N_40782);
or U44421 (N_44421,N_42448,N_42436);
xor U44422 (N_44422,N_40382,N_42269);
xnor U44423 (N_44423,N_40682,N_42334);
nand U44424 (N_44424,N_40332,N_42213);
xor U44425 (N_44425,N_40853,N_40628);
xnor U44426 (N_44426,N_41757,N_41851);
nand U44427 (N_44427,N_42269,N_40471);
nand U44428 (N_44428,N_40371,N_41615);
nand U44429 (N_44429,N_42001,N_41997);
or U44430 (N_44430,N_41109,N_42218);
and U44431 (N_44431,N_41649,N_40695);
nor U44432 (N_44432,N_42299,N_41284);
and U44433 (N_44433,N_41108,N_42463);
nor U44434 (N_44434,N_40105,N_41601);
nand U44435 (N_44435,N_42207,N_40129);
nor U44436 (N_44436,N_41440,N_42335);
or U44437 (N_44437,N_40220,N_41393);
nand U44438 (N_44438,N_41725,N_41442);
nand U44439 (N_44439,N_42072,N_41584);
nor U44440 (N_44440,N_40201,N_41986);
and U44441 (N_44441,N_40841,N_41119);
nor U44442 (N_44442,N_41927,N_40050);
nand U44443 (N_44443,N_40266,N_41959);
and U44444 (N_44444,N_40911,N_41213);
nand U44445 (N_44445,N_41582,N_40491);
or U44446 (N_44446,N_41340,N_41066);
and U44447 (N_44447,N_41608,N_41748);
and U44448 (N_44448,N_41559,N_41507);
xor U44449 (N_44449,N_40669,N_40081);
and U44450 (N_44450,N_41043,N_41123);
nand U44451 (N_44451,N_41431,N_42430);
or U44452 (N_44452,N_42005,N_40714);
xnor U44453 (N_44453,N_41401,N_40830);
and U44454 (N_44454,N_40129,N_42270);
nand U44455 (N_44455,N_41989,N_41737);
nor U44456 (N_44456,N_40778,N_40824);
and U44457 (N_44457,N_42285,N_42008);
nor U44458 (N_44458,N_42473,N_41503);
xnor U44459 (N_44459,N_40310,N_41059);
nor U44460 (N_44460,N_41974,N_40891);
nor U44461 (N_44461,N_40255,N_42310);
nor U44462 (N_44462,N_40905,N_40323);
xnor U44463 (N_44463,N_42146,N_40779);
nor U44464 (N_44464,N_41718,N_40228);
and U44465 (N_44465,N_40366,N_41264);
and U44466 (N_44466,N_41821,N_40025);
nor U44467 (N_44467,N_42184,N_40896);
nand U44468 (N_44468,N_40762,N_41754);
xnor U44469 (N_44469,N_42008,N_41225);
nor U44470 (N_44470,N_40497,N_41826);
nand U44471 (N_44471,N_40654,N_40697);
and U44472 (N_44472,N_40040,N_41482);
nand U44473 (N_44473,N_41530,N_42370);
nand U44474 (N_44474,N_41897,N_42035);
nand U44475 (N_44475,N_42133,N_41019);
nand U44476 (N_44476,N_41274,N_40340);
nand U44477 (N_44477,N_40473,N_41763);
xnor U44478 (N_44478,N_41890,N_40947);
nand U44479 (N_44479,N_42074,N_41484);
nand U44480 (N_44480,N_40464,N_42291);
nand U44481 (N_44481,N_40977,N_40841);
xnor U44482 (N_44482,N_40332,N_42260);
or U44483 (N_44483,N_40251,N_40659);
or U44484 (N_44484,N_41930,N_41646);
nor U44485 (N_44485,N_41251,N_40137);
or U44486 (N_44486,N_41848,N_41818);
nor U44487 (N_44487,N_41379,N_42188);
nor U44488 (N_44488,N_40490,N_41091);
xor U44489 (N_44489,N_40469,N_40032);
or U44490 (N_44490,N_40266,N_40433);
and U44491 (N_44491,N_41250,N_42442);
nand U44492 (N_44492,N_41395,N_41864);
nor U44493 (N_44493,N_41312,N_42370);
xnor U44494 (N_44494,N_42064,N_41075);
nor U44495 (N_44495,N_42072,N_40791);
nor U44496 (N_44496,N_40440,N_41680);
xor U44497 (N_44497,N_41772,N_41221);
or U44498 (N_44498,N_40247,N_40972);
or U44499 (N_44499,N_42268,N_41132);
xnor U44500 (N_44500,N_41986,N_40480);
and U44501 (N_44501,N_40776,N_41293);
xnor U44502 (N_44502,N_40238,N_40859);
nor U44503 (N_44503,N_41255,N_42276);
or U44504 (N_44504,N_40688,N_41134);
or U44505 (N_44505,N_40470,N_40706);
or U44506 (N_44506,N_41951,N_40085);
nand U44507 (N_44507,N_41923,N_40187);
or U44508 (N_44508,N_42053,N_42136);
or U44509 (N_44509,N_40130,N_41105);
or U44510 (N_44510,N_40579,N_40626);
or U44511 (N_44511,N_41427,N_40815);
nand U44512 (N_44512,N_41140,N_41163);
xor U44513 (N_44513,N_40850,N_41212);
or U44514 (N_44514,N_40831,N_41516);
nor U44515 (N_44515,N_40645,N_40696);
nor U44516 (N_44516,N_40759,N_41831);
or U44517 (N_44517,N_42383,N_40805);
or U44518 (N_44518,N_40457,N_40050);
xor U44519 (N_44519,N_40614,N_40429);
or U44520 (N_44520,N_41191,N_40340);
or U44521 (N_44521,N_41031,N_40344);
or U44522 (N_44522,N_42384,N_40615);
or U44523 (N_44523,N_41780,N_41371);
or U44524 (N_44524,N_40705,N_40370);
xnor U44525 (N_44525,N_41043,N_40942);
nand U44526 (N_44526,N_42274,N_42031);
nor U44527 (N_44527,N_42147,N_41570);
or U44528 (N_44528,N_41479,N_40600);
xnor U44529 (N_44529,N_40885,N_41556);
or U44530 (N_44530,N_41514,N_40550);
nor U44531 (N_44531,N_41983,N_42104);
xnor U44532 (N_44532,N_40871,N_41953);
and U44533 (N_44533,N_40764,N_41850);
nand U44534 (N_44534,N_40225,N_41941);
nand U44535 (N_44535,N_41436,N_41546);
and U44536 (N_44536,N_41834,N_42336);
nor U44537 (N_44537,N_42120,N_41900);
nor U44538 (N_44538,N_41636,N_40804);
and U44539 (N_44539,N_41976,N_42403);
and U44540 (N_44540,N_40339,N_40695);
or U44541 (N_44541,N_41248,N_41520);
xor U44542 (N_44542,N_40117,N_42009);
or U44543 (N_44543,N_41901,N_41509);
and U44544 (N_44544,N_40474,N_40618);
or U44545 (N_44545,N_42450,N_42050);
nand U44546 (N_44546,N_41536,N_40604);
nand U44547 (N_44547,N_42164,N_40756);
and U44548 (N_44548,N_40423,N_40762);
nor U44549 (N_44549,N_41762,N_40190);
and U44550 (N_44550,N_42118,N_41958);
and U44551 (N_44551,N_40013,N_42054);
nor U44552 (N_44552,N_40566,N_40751);
nand U44553 (N_44553,N_41474,N_41304);
and U44554 (N_44554,N_41207,N_41742);
xnor U44555 (N_44555,N_40263,N_40101);
nand U44556 (N_44556,N_42096,N_41708);
nand U44557 (N_44557,N_40824,N_41839);
nand U44558 (N_44558,N_41028,N_41266);
xor U44559 (N_44559,N_42117,N_41884);
xnor U44560 (N_44560,N_42170,N_40124);
xor U44561 (N_44561,N_41291,N_42233);
nand U44562 (N_44562,N_41552,N_40370);
or U44563 (N_44563,N_41756,N_40355);
or U44564 (N_44564,N_41059,N_41772);
nand U44565 (N_44565,N_41821,N_41311);
xor U44566 (N_44566,N_41152,N_41524);
nand U44567 (N_44567,N_40018,N_40613);
and U44568 (N_44568,N_42107,N_41919);
xnor U44569 (N_44569,N_41753,N_42371);
xor U44570 (N_44570,N_41853,N_41650);
and U44571 (N_44571,N_41237,N_42098);
xnor U44572 (N_44572,N_40489,N_41014);
or U44573 (N_44573,N_40197,N_40788);
and U44574 (N_44574,N_40189,N_41576);
xor U44575 (N_44575,N_42031,N_41713);
nand U44576 (N_44576,N_40740,N_42468);
nor U44577 (N_44577,N_42389,N_40627);
xor U44578 (N_44578,N_40674,N_41021);
nor U44579 (N_44579,N_41886,N_41502);
nor U44580 (N_44580,N_41382,N_42070);
or U44581 (N_44581,N_40260,N_40198);
nand U44582 (N_44582,N_41038,N_42305);
or U44583 (N_44583,N_40792,N_40598);
nand U44584 (N_44584,N_40230,N_40255);
and U44585 (N_44585,N_40727,N_40785);
nand U44586 (N_44586,N_40476,N_41296);
nor U44587 (N_44587,N_40959,N_40495);
and U44588 (N_44588,N_41379,N_41646);
xor U44589 (N_44589,N_41552,N_41380);
nand U44590 (N_44590,N_42369,N_41608);
and U44591 (N_44591,N_41708,N_40791);
nand U44592 (N_44592,N_42297,N_40575);
or U44593 (N_44593,N_42414,N_42114);
nand U44594 (N_44594,N_41901,N_42346);
and U44595 (N_44595,N_41110,N_41952);
or U44596 (N_44596,N_41191,N_42417);
nand U44597 (N_44597,N_40265,N_40322);
nor U44598 (N_44598,N_41815,N_40166);
nand U44599 (N_44599,N_40508,N_40797);
nor U44600 (N_44600,N_42453,N_41567);
xor U44601 (N_44601,N_41334,N_41145);
nor U44602 (N_44602,N_40674,N_40029);
nor U44603 (N_44603,N_41444,N_41156);
xor U44604 (N_44604,N_40944,N_40768);
and U44605 (N_44605,N_42397,N_41144);
and U44606 (N_44606,N_41657,N_42431);
nor U44607 (N_44607,N_40628,N_41573);
xor U44608 (N_44608,N_40564,N_41314);
xor U44609 (N_44609,N_41344,N_40800);
and U44610 (N_44610,N_41030,N_41664);
nand U44611 (N_44611,N_41275,N_41763);
nor U44612 (N_44612,N_42236,N_42006);
or U44613 (N_44613,N_41006,N_40577);
and U44614 (N_44614,N_41190,N_41484);
nand U44615 (N_44615,N_41814,N_40140);
nand U44616 (N_44616,N_42450,N_42223);
or U44617 (N_44617,N_41837,N_42267);
nand U44618 (N_44618,N_41150,N_41220);
nand U44619 (N_44619,N_40899,N_42378);
nand U44620 (N_44620,N_41394,N_41420);
or U44621 (N_44621,N_40307,N_41995);
nand U44622 (N_44622,N_40764,N_40258);
xor U44623 (N_44623,N_40008,N_41149);
and U44624 (N_44624,N_42174,N_41094);
nor U44625 (N_44625,N_41420,N_40135);
nand U44626 (N_44626,N_41318,N_40005);
or U44627 (N_44627,N_41762,N_41256);
nand U44628 (N_44628,N_42020,N_42424);
and U44629 (N_44629,N_41377,N_40215);
nand U44630 (N_44630,N_41165,N_42417);
or U44631 (N_44631,N_42000,N_41424);
nor U44632 (N_44632,N_41569,N_41722);
or U44633 (N_44633,N_41741,N_42006);
or U44634 (N_44634,N_42296,N_40195);
nand U44635 (N_44635,N_40045,N_40451);
or U44636 (N_44636,N_40191,N_41213);
nor U44637 (N_44637,N_42199,N_40583);
xnor U44638 (N_44638,N_41118,N_42498);
nand U44639 (N_44639,N_41300,N_41331);
nor U44640 (N_44640,N_41982,N_40217);
xor U44641 (N_44641,N_40160,N_40787);
xnor U44642 (N_44642,N_40593,N_41053);
and U44643 (N_44643,N_41221,N_41807);
or U44644 (N_44644,N_41857,N_40131);
nor U44645 (N_44645,N_40949,N_40669);
nor U44646 (N_44646,N_40248,N_42355);
or U44647 (N_44647,N_42405,N_41930);
xor U44648 (N_44648,N_41782,N_42189);
xor U44649 (N_44649,N_41773,N_40932);
nor U44650 (N_44650,N_42343,N_40373);
or U44651 (N_44651,N_42355,N_41312);
nand U44652 (N_44652,N_41676,N_40050);
or U44653 (N_44653,N_40661,N_40225);
and U44654 (N_44654,N_41630,N_41151);
or U44655 (N_44655,N_41246,N_41395);
xor U44656 (N_44656,N_40021,N_41351);
nand U44657 (N_44657,N_42119,N_41594);
or U44658 (N_44658,N_41549,N_40934);
and U44659 (N_44659,N_42225,N_41250);
nor U44660 (N_44660,N_41935,N_40328);
nand U44661 (N_44661,N_42257,N_41631);
nand U44662 (N_44662,N_42172,N_41263);
nand U44663 (N_44663,N_42093,N_40952);
nand U44664 (N_44664,N_40583,N_40144);
or U44665 (N_44665,N_41420,N_41397);
xor U44666 (N_44666,N_40843,N_41079);
or U44667 (N_44667,N_41977,N_40477);
nor U44668 (N_44668,N_41767,N_40196);
and U44669 (N_44669,N_41232,N_40712);
nand U44670 (N_44670,N_40088,N_41291);
or U44671 (N_44671,N_42305,N_41817);
nor U44672 (N_44672,N_40740,N_41280);
nand U44673 (N_44673,N_42375,N_42457);
nand U44674 (N_44674,N_42361,N_41083);
nor U44675 (N_44675,N_40030,N_40116);
nand U44676 (N_44676,N_40905,N_40631);
or U44677 (N_44677,N_40946,N_41901);
nor U44678 (N_44678,N_40092,N_42046);
and U44679 (N_44679,N_40956,N_41026);
nand U44680 (N_44680,N_42180,N_42362);
or U44681 (N_44681,N_40541,N_41312);
nor U44682 (N_44682,N_40802,N_41959);
nand U44683 (N_44683,N_41655,N_40586);
or U44684 (N_44684,N_41644,N_41050);
xor U44685 (N_44685,N_41903,N_41856);
nor U44686 (N_44686,N_41749,N_40737);
and U44687 (N_44687,N_42116,N_42455);
xnor U44688 (N_44688,N_41800,N_42255);
nor U44689 (N_44689,N_40594,N_41174);
nand U44690 (N_44690,N_41635,N_42187);
nor U44691 (N_44691,N_42284,N_42424);
nor U44692 (N_44692,N_42416,N_41402);
and U44693 (N_44693,N_41428,N_41963);
xnor U44694 (N_44694,N_41086,N_40742);
nor U44695 (N_44695,N_40789,N_40091);
or U44696 (N_44696,N_41608,N_41968);
nand U44697 (N_44697,N_40557,N_41345);
nand U44698 (N_44698,N_42198,N_40114);
nor U44699 (N_44699,N_42069,N_41643);
and U44700 (N_44700,N_41160,N_41449);
nor U44701 (N_44701,N_40633,N_40143);
nand U44702 (N_44702,N_40673,N_41612);
or U44703 (N_44703,N_41748,N_42378);
nand U44704 (N_44704,N_40927,N_40102);
nand U44705 (N_44705,N_40797,N_42221);
or U44706 (N_44706,N_42275,N_42124);
nand U44707 (N_44707,N_42044,N_41754);
nor U44708 (N_44708,N_42245,N_40582);
and U44709 (N_44709,N_40942,N_40020);
xnor U44710 (N_44710,N_40360,N_41137);
or U44711 (N_44711,N_40975,N_40308);
and U44712 (N_44712,N_41990,N_40702);
and U44713 (N_44713,N_42123,N_41468);
and U44714 (N_44714,N_41880,N_42035);
xor U44715 (N_44715,N_40721,N_41845);
nor U44716 (N_44716,N_41694,N_41239);
and U44717 (N_44717,N_42471,N_41272);
nand U44718 (N_44718,N_40828,N_41047);
nand U44719 (N_44719,N_42364,N_41717);
xor U44720 (N_44720,N_40845,N_41891);
xor U44721 (N_44721,N_41387,N_42066);
and U44722 (N_44722,N_41438,N_41932);
xnor U44723 (N_44723,N_40948,N_40255);
or U44724 (N_44724,N_41934,N_41984);
nor U44725 (N_44725,N_40208,N_41593);
nand U44726 (N_44726,N_41297,N_41505);
nand U44727 (N_44727,N_40028,N_40142);
nand U44728 (N_44728,N_40993,N_40504);
and U44729 (N_44729,N_41170,N_40141);
xnor U44730 (N_44730,N_40669,N_41831);
nor U44731 (N_44731,N_41298,N_41068);
or U44732 (N_44732,N_41258,N_41868);
and U44733 (N_44733,N_40129,N_40838);
nand U44734 (N_44734,N_40392,N_42348);
nor U44735 (N_44735,N_42481,N_41835);
or U44736 (N_44736,N_40877,N_40886);
xnor U44737 (N_44737,N_41803,N_41175);
nand U44738 (N_44738,N_41078,N_41416);
or U44739 (N_44739,N_42017,N_40865);
and U44740 (N_44740,N_41708,N_40461);
nor U44741 (N_44741,N_42326,N_42292);
xor U44742 (N_44742,N_41620,N_41825);
nor U44743 (N_44743,N_40609,N_40118);
or U44744 (N_44744,N_41480,N_41340);
nor U44745 (N_44745,N_40017,N_40445);
and U44746 (N_44746,N_41678,N_40505);
xor U44747 (N_44747,N_41106,N_40945);
nand U44748 (N_44748,N_41942,N_40933);
nand U44749 (N_44749,N_40822,N_40841);
xnor U44750 (N_44750,N_41225,N_42254);
nor U44751 (N_44751,N_40590,N_40975);
nor U44752 (N_44752,N_40968,N_41774);
and U44753 (N_44753,N_40021,N_40955);
nand U44754 (N_44754,N_41171,N_40334);
nor U44755 (N_44755,N_41407,N_40882);
nand U44756 (N_44756,N_40984,N_40455);
nor U44757 (N_44757,N_41712,N_41421);
and U44758 (N_44758,N_41051,N_41249);
xor U44759 (N_44759,N_40311,N_42283);
nand U44760 (N_44760,N_40377,N_41258);
nand U44761 (N_44761,N_42243,N_42469);
xor U44762 (N_44762,N_40547,N_41510);
and U44763 (N_44763,N_41577,N_42381);
or U44764 (N_44764,N_41710,N_40686);
nand U44765 (N_44765,N_40764,N_41893);
nand U44766 (N_44766,N_41414,N_41549);
and U44767 (N_44767,N_40105,N_41650);
nand U44768 (N_44768,N_41128,N_41895);
nor U44769 (N_44769,N_41985,N_42319);
nor U44770 (N_44770,N_42064,N_40884);
and U44771 (N_44771,N_42149,N_41823);
or U44772 (N_44772,N_40472,N_42464);
xor U44773 (N_44773,N_40379,N_40725);
nor U44774 (N_44774,N_42304,N_42393);
nor U44775 (N_44775,N_42083,N_41716);
or U44776 (N_44776,N_41657,N_40811);
xor U44777 (N_44777,N_41783,N_40454);
nor U44778 (N_44778,N_42491,N_41029);
nor U44779 (N_44779,N_40463,N_40162);
xnor U44780 (N_44780,N_41904,N_41921);
xor U44781 (N_44781,N_42475,N_40278);
nand U44782 (N_44782,N_40279,N_40801);
or U44783 (N_44783,N_40711,N_40786);
and U44784 (N_44784,N_42126,N_40975);
nor U44785 (N_44785,N_42265,N_40734);
or U44786 (N_44786,N_41298,N_41810);
or U44787 (N_44787,N_40659,N_40140);
or U44788 (N_44788,N_40077,N_41136);
nor U44789 (N_44789,N_41990,N_41933);
and U44790 (N_44790,N_40731,N_40613);
nor U44791 (N_44791,N_41925,N_41543);
nand U44792 (N_44792,N_40460,N_42121);
or U44793 (N_44793,N_41484,N_41157);
nor U44794 (N_44794,N_40312,N_40935);
nand U44795 (N_44795,N_40958,N_41428);
nand U44796 (N_44796,N_41557,N_42487);
or U44797 (N_44797,N_40574,N_40387);
and U44798 (N_44798,N_40193,N_41109);
and U44799 (N_44799,N_41235,N_41444);
nand U44800 (N_44800,N_40524,N_41496);
or U44801 (N_44801,N_42462,N_42100);
nand U44802 (N_44802,N_40927,N_40208);
and U44803 (N_44803,N_40036,N_40224);
and U44804 (N_44804,N_41345,N_40880);
xnor U44805 (N_44805,N_40653,N_42224);
or U44806 (N_44806,N_41272,N_41782);
or U44807 (N_44807,N_40002,N_40227);
nor U44808 (N_44808,N_41593,N_40418);
and U44809 (N_44809,N_40435,N_42430);
nand U44810 (N_44810,N_41244,N_41609);
xor U44811 (N_44811,N_42055,N_41759);
nand U44812 (N_44812,N_41605,N_40986);
nand U44813 (N_44813,N_41172,N_42107);
xnor U44814 (N_44814,N_40169,N_41641);
xnor U44815 (N_44815,N_41679,N_40492);
nor U44816 (N_44816,N_42358,N_42089);
nand U44817 (N_44817,N_40982,N_40379);
and U44818 (N_44818,N_40959,N_40383);
nor U44819 (N_44819,N_41900,N_40930);
nor U44820 (N_44820,N_41113,N_41334);
and U44821 (N_44821,N_40961,N_41488);
nor U44822 (N_44822,N_40311,N_40224);
xnor U44823 (N_44823,N_41511,N_40328);
nand U44824 (N_44824,N_42370,N_41944);
xor U44825 (N_44825,N_42384,N_41125);
xnor U44826 (N_44826,N_42099,N_40500);
or U44827 (N_44827,N_41757,N_41955);
nor U44828 (N_44828,N_41295,N_41944);
xor U44829 (N_44829,N_40299,N_41836);
and U44830 (N_44830,N_40262,N_40249);
or U44831 (N_44831,N_42407,N_42011);
xor U44832 (N_44832,N_42020,N_41273);
nand U44833 (N_44833,N_40299,N_41629);
and U44834 (N_44834,N_42294,N_41675);
and U44835 (N_44835,N_42180,N_41279);
or U44836 (N_44836,N_40889,N_41695);
nor U44837 (N_44837,N_41128,N_40257);
xor U44838 (N_44838,N_40349,N_40938);
and U44839 (N_44839,N_41266,N_41416);
xor U44840 (N_44840,N_41484,N_41375);
nand U44841 (N_44841,N_41857,N_40477);
nand U44842 (N_44842,N_41674,N_41052);
xnor U44843 (N_44843,N_40682,N_40084);
nor U44844 (N_44844,N_42035,N_40940);
nand U44845 (N_44845,N_40266,N_42168);
nand U44846 (N_44846,N_42147,N_42322);
nor U44847 (N_44847,N_40836,N_42499);
nor U44848 (N_44848,N_40360,N_41495);
or U44849 (N_44849,N_40982,N_41744);
nor U44850 (N_44850,N_41505,N_41440);
and U44851 (N_44851,N_40142,N_41321);
nor U44852 (N_44852,N_40091,N_42436);
xor U44853 (N_44853,N_42053,N_41107);
or U44854 (N_44854,N_40220,N_41255);
or U44855 (N_44855,N_40486,N_42407);
nand U44856 (N_44856,N_40686,N_42430);
xor U44857 (N_44857,N_40119,N_42238);
nor U44858 (N_44858,N_41644,N_40155);
nor U44859 (N_44859,N_40938,N_42450);
xor U44860 (N_44860,N_41920,N_40286);
or U44861 (N_44861,N_40466,N_40940);
xor U44862 (N_44862,N_41706,N_42484);
xor U44863 (N_44863,N_41520,N_41067);
or U44864 (N_44864,N_40853,N_42376);
nor U44865 (N_44865,N_40830,N_42267);
nand U44866 (N_44866,N_40552,N_41055);
xor U44867 (N_44867,N_40647,N_41729);
nor U44868 (N_44868,N_40476,N_40641);
and U44869 (N_44869,N_40186,N_42354);
or U44870 (N_44870,N_41549,N_41426);
and U44871 (N_44871,N_42077,N_42372);
and U44872 (N_44872,N_40722,N_41570);
xor U44873 (N_44873,N_40139,N_40175);
and U44874 (N_44874,N_41935,N_41357);
nor U44875 (N_44875,N_42140,N_40248);
nand U44876 (N_44876,N_41731,N_40693);
and U44877 (N_44877,N_40074,N_40225);
or U44878 (N_44878,N_42050,N_42031);
or U44879 (N_44879,N_41143,N_41436);
nand U44880 (N_44880,N_40650,N_41845);
or U44881 (N_44881,N_41986,N_40039);
nand U44882 (N_44882,N_40961,N_40914);
nor U44883 (N_44883,N_40437,N_40375);
and U44884 (N_44884,N_42205,N_41167);
nor U44885 (N_44885,N_41346,N_42482);
xnor U44886 (N_44886,N_41730,N_41098);
nand U44887 (N_44887,N_40585,N_41653);
nor U44888 (N_44888,N_42359,N_40773);
or U44889 (N_44889,N_40231,N_40143);
and U44890 (N_44890,N_41007,N_40321);
nor U44891 (N_44891,N_42066,N_42351);
and U44892 (N_44892,N_41885,N_41611);
and U44893 (N_44893,N_41627,N_41375);
nand U44894 (N_44894,N_41450,N_40110);
and U44895 (N_44895,N_40436,N_41335);
nor U44896 (N_44896,N_41935,N_40888);
and U44897 (N_44897,N_41310,N_41938);
or U44898 (N_44898,N_41299,N_40164);
xnor U44899 (N_44899,N_41971,N_41884);
and U44900 (N_44900,N_42153,N_41879);
xnor U44901 (N_44901,N_41509,N_41828);
xor U44902 (N_44902,N_40748,N_42001);
or U44903 (N_44903,N_42105,N_40022);
nor U44904 (N_44904,N_42057,N_41946);
and U44905 (N_44905,N_42011,N_41493);
or U44906 (N_44906,N_40666,N_41638);
or U44907 (N_44907,N_40424,N_41022);
nand U44908 (N_44908,N_40715,N_42469);
nor U44909 (N_44909,N_40234,N_42095);
xor U44910 (N_44910,N_40141,N_40901);
or U44911 (N_44911,N_40201,N_40233);
nor U44912 (N_44912,N_41193,N_42406);
and U44913 (N_44913,N_40033,N_41078);
and U44914 (N_44914,N_40598,N_40427);
and U44915 (N_44915,N_41048,N_41486);
and U44916 (N_44916,N_41157,N_41021);
nand U44917 (N_44917,N_42423,N_41805);
or U44918 (N_44918,N_41392,N_41835);
and U44919 (N_44919,N_41291,N_41134);
nor U44920 (N_44920,N_42233,N_41690);
nand U44921 (N_44921,N_42266,N_41686);
or U44922 (N_44922,N_41044,N_40517);
xor U44923 (N_44923,N_42349,N_40113);
or U44924 (N_44924,N_40341,N_42169);
and U44925 (N_44925,N_42465,N_40726);
or U44926 (N_44926,N_42418,N_40664);
or U44927 (N_44927,N_40578,N_41663);
nor U44928 (N_44928,N_41386,N_40630);
nand U44929 (N_44929,N_42457,N_41954);
nand U44930 (N_44930,N_40534,N_41053);
and U44931 (N_44931,N_40796,N_40769);
nor U44932 (N_44932,N_42401,N_42021);
or U44933 (N_44933,N_40061,N_41462);
nor U44934 (N_44934,N_41634,N_40367);
nand U44935 (N_44935,N_40764,N_41013);
nand U44936 (N_44936,N_41457,N_40885);
or U44937 (N_44937,N_41314,N_42384);
nand U44938 (N_44938,N_40603,N_41329);
nor U44939 (N_44939,N_40484,N_40895);
xor U44940 (N_44940,N_40289,N_41424);
nand U44941 (N_44941,N_40839,N_40401);
xnor U44942 (N_44942,N_40205,N_42067);
and U44943 (N_44943,N_41947,N_42450);
and U44944 (N_44944,N_41422,N_40104);
and U44945 (N_44945,N_40222,N_41468);
nor U44946 (N_44946,N_40851,N_40070);
nor U44947 (N_44947,N_40753,N_41301);
nand U44948 (N_44948,N_40292,N_42197);
nor U44949 (N_44949,N_40535,N_40778);
nor U44950 (N_44950,N_42438,N_40105);
and U44951 (N_44951,N_41815,N_42122);
xnor U44952 (N_44952,N_41709,N_40242);
nor U44953 (N_44953,N_41314,N_41174);
and U44954 (N_44954,N_42393,N_42219);
and U44955 (N_44955,N_40611,N_40699);
or U44956 (N_44956,N_41297,N_41381);
and U44957 (N_44957,N_40135,N_41141);
nand U44958 (N_44958,N_41040,N_40992);
or U44959 (N_44959,N_41411,N_40373);
nand U44960 (N_44960,N_41686,N_40638);
nor U44961 (N_44961,N_41896,N_42160);
or U44962 (N_44962,N_40789,N_42173);
xor U44963 (N_44963,N_42241,N_41381);
xnor U44964 (N_44964,N_41537,N_41706);
nor U44965 (N_44965,N_41820,N_40844);
and U44966 (N_44966,N_41114,N_41394);
nand U44967 (N_44967,N_40512,N_41093);
or U44968 (N_44968,N_40109,N_42146);
or U44969 (N_44969,N_40535,N_41957);
xor U44970 (N_44970,N_41511,N_40746);
nor U44971 (N_44971,N_42009,N_42368);
and U44972 (N_44972,N_41212,N_40612);
nand U44973 (N_44973,N_42076,N_40237);
xor U44974 (N_44974,N_41307,N_41238);
nand U44975 (N_44975,N_40857,N_42332);
nand U44976 (N_44976,N_41962,N_40313);
nand U44977 (N_44977,N_41898,N_40249);
nor U44978 (N_44978,N_41546,N_40112);
nor U44979 (N_44979,N_40905,N_40410);
and U44980 (N_44980,N_40729,N_41054);
nor U44981 (N_44981,N_41822,N_40722);
and U44982 (N_44982,N_41761,N_40630);
nand U44983 (N_44983,N_40931,N_40603);
and U44984 (N_44984,N_41819,N_40856);
or U44985 (N_44985,N_41316,N_41978);
and U44986 (N_44986,N_42352,N_41108);
nor U44987 (N_44987,N_40664,N_42009);
or U44988 (N_44988,N_41018,N_40207);
nor U44989 (N_44989,N_41691,N_41079);
or U44990 (N_44990,N_41873,N_41071);
and U44991 (N_44991,N_42047,N_40780);
and U44992 (N_44992,N_40486,N_41263);
nand U44993 (N_44993,N_42183,N_42137);
nand U44994 (N_44994,N_42108,N_41048);
nor U44995 (N_44995,N_41251,N_41505);
nand U44996 (N_44996,N_40324,N_40971);
nand U44997 (N_44997,N_40623,N_40610);
nor U44998 (N_44998,N_40671,N_41131);
xnor U44999 (N_44999,N_41654,N_41470);
nor U45000 (N_45000,N_43858,N_43615);
or U45001 (N_45001,N_44237,N_44012);
xor U45002 (N_45002,N_44146,N_43096);
and U45003 (N_45003,N_42655,N_44252);
nand U45004 (N_45004,N_42522,N_43048);
or U45005 (N_45005,N_43838,N_44007);
xnor U45006 (N_45006,N_43047,N_43575);
nor U45007 (N_45007,N_42727,N_44937);
or U45008 (N_45008,N_44988,N_43794);
nand U45009 (N_45009,N_44393,N_43177);
nor U45010 (N_45010,N_42913,N_44998);
and U45011 (N_45011,N_43184,N_42753);
nand U45012 (N_45012,N_43148,N_44339);
and U45013 (N_45013,N_43694,N_42578);
xnor U45014 (N_45014,N_44745,N_44197);
nor U45015 (N_45015,N_43283,N_44000);
or U45016 (N_45016,N_44497,N_43539);
xor U45017 (N_45017,N_42669,N_43917);
nand U45018 (N_45018,N_44606,N_44679);
or U45019 (N_45019,N_44288,N_44825);
nand U45020 (N_45020,N_44722,N_44730);
and U45021 (N_45021,N_42979,N_44807);
or U45022 (N_45022,N_44354,N_42666);
nor U45023 (N_45023,N_42795,N_43482);
and U45024 (N_45024,N_43278,N_42665);
xnor U45025 (N_45025,N_44250,N_44112);
or U45026 (N_45026,N_44641,N_44590);
nor U45027 (N_45027,N_43513,N_44527);
xnor U45028 (N_45028,N_43018,N_43469);
xnor U45029 (N_45029,N_44915,N_43141);
nand U45030 (N_45030,N_43679,N_43366);
xor U45031 (N_45031,N_42521,N_44892);
xor U45032 (N_45032,N_43876,N_44551);
xnor U45033 (N_45033,N_44109,N_43788);
nand U45034 (N_45034,N_44772,N_43693);
or U45035 (N_45035,N_43673,N_44259);
nand U45036 (N_45036,N_42944,N_43302);
nor U45037 (N_45037,N_43761,N_43831);
xor U45038 (N_45038,N_44689,N_44559);
nand U45039 (N_45039,N_44879,N_44852);
nand U45040 (N_45040,N_43394,N_43660);
xnor U45041 (N_45041,N_42853,N_43641);
nor U45042 (N_45042,N_44349,N_44838);
nor U45043 (N_45043,N_43455,N_44913);
nor U45044 (N_45044,N_43985,N_43465);
and U45045 (N_45045,N_44344,N_44886);
nor U45046 (N_45046,N_42626,N_43384);
and U45047 (N_45047,N_44663,N_43074);
xnor U45048 (N_45048,N_44002,N_43004);
and U45049 (N_45049,N_44413,N_44990);
or U45050 (N_45050,N_43826,N_43578);
nand U45051 (N_45051,N_43653,N_43087);
xnor U45052 (N_45052,N_43506,N_43458);
nor U45053 (N_45053,N_43981,N_43994);
xnor U45054 (N_45054,N_43582,N_42965);
and U45055 (N_45055,N_43542,N_44704);
xor U45056 (N_45056,N_44383,N_43597);
or U45057 (N_45057,N_44909,N_43421);
nor U45058 (N_45058,N_42553,N_43704);
xnor U45059 (N_45059,N_42502,N_44940);
and U45060 (N_45060,N_44900,N_42635);
or U45061 (N_45061,N_43785,N_44968);
xor U45062 (N_45062,N_44020,N_44938);
xnor U45063 (N_45063,N_43197,N_43564);
nand U45064 (N_45064,N_42875,N_43198);
nand U45065 (N_45065,N_43752,N_43897);
and U45066 (N_45066,N_43367,N_44747);
and U45067 (N_45067,N_42963,N_43452);
xnor U45068 (N_45068,N_43487,N_44669);
or U45069 (N_45069,N_42791,N_44549);
or U45070 (N_45070,N_43762,N_44717);
nor U45071 (N_45071,N_43988,N_43094);
or U45072 (N_45072,N_42611,N_44723);
nand U45073 (N_45073,N_43472,N_43676);
nand U45074 (N_45074,N_44902,N_42551);
xnor U45075 (N_45075,N_43900,N_44672);
nand U45076 (N_45076,N_43436,N_43872);
nand U45077 (N_45077,N_44552,N_43159);
or U45078 (N_45078,N_44342,N_43435);
nor U45079 (N_45079,N_43158,N_44166);
nor U45080 (N_45080,N_44743,N_44885);
xor U45081 (N_45081,N_43750,N_42878);
or U45082 (N_45082,N_44801,N_44207);
and U45083 (N_45083,N_44853,N_43282);
nor U45084 (N_45084,N_43376,N_44217);
xor U45085 (N_45085,N_44280,N_44253);
xor U45086 (N_45086,N_43360,N_43783);
or U45087 (N_45087,N_44691,N_42811);
xor U45088 (N_45088,N_43233,N_43416);
or U45089 (N_45089,N_43108,N_42579);
nor U45090 (N_45090,N_43522,N_42829);
nor U45091 (N_45091,N_44188,N_42743);
nor U45092 (N_45092,N_43816,N_42572);
and U45093 (N_45093,N_42988,N_44578);
and U45094 (N_45094,N_43150,N_44563);
and U45095 (N_45095,N_43099,N_42886);
and U45096 (N_45096,N_43927,N_43330);
nor U45097 (N_45097,N_42971,N_43844);
xor U45098 (N_45098,N_43590,N_43885);
and U45099 (N_45099,N_42636,N_44177);
nor U45100 (N_45100,N_44665,N_43447);
xor U45101 (N_45101,N_44428,N_43336);
nand U45102 (N_45102,N_44303,N_44041);
xnor U45103 (N_45103,N_42687,N_42792);
or U45104 (N_45104,N_42747,N_43772);
nor U45105 (N_45105,N_44827,N_43942);
nand U45106 (N_45106,N_44509,N_42726);
nor U45107 (N_45107,N_42667,N_42569);
or U45108 (N_45108,N_42891,N_43133);
nand U45109 (N_45109,N_44486,N_44300);
or U45110 (N_45110,N_44321,N_43378);
nand U45111 (N_45111,N_44681,N_44524);
xnor U45112 (N_45112,N_43869,N_42542);
or U45113 (N_45113,N_44986,N_44397);
nor U45114 (N_45114,N_44107,N_42748);
xor U45115 (N_45115,N_44334,N_44792);
and U45116 (N_45116,N_44036,N_43646);
xor U45117 (N_45117,N_44292,N_43424);
and U45118 (N_45118,N_43552,N_42735);
xor U45119 (N_45119,N_43996,N_43304);
and U45120 (N_45120,N_43138,N_42555);
or U45121 (N_45121,N_43587,N_43026);
or U45122 (N_45122,N_42613,N_42739);
and U45123 (N_45123,N_42856,N_42862);
nor U45124 (N_45124,N_44193,N_43683);
nand U45125 (N_45125,N_44351,N_44750);
and U45126 (N_45126,N_44184,N_43797);
nand U45127 (N_45127,N_44971,N_43556);
nor U45128 (N_45128,N_44330,N_43796);
nand U45129 (N_45129,N_44026,N_43120);
or U45130 (N_45130,N_44991,N_42616);
nand U45131 (N_45131,N_44298,N_44888);
and U45132 (N_45132,N_43489,N_44198);
nor U45133 (N_45133,N_43861,N_43616);
xor U45134 (N_45134,N_44978,N_42884);
nand U45135 (N_45135,N_43437,N_43520);
or U45136 (N_45136,N_43187,N_43977);
nor U45137 (N_45137,N_44183,N_44864);
nand U45138 (N_45138,N_43650,N_43205);
and U45139 (N_45139,N_42529,N_43260);
nor U45140 (N_45140,N_43031,N_43253);
nor U45141 (N_45141,N_44618,N_44287);
nor U45142 (N_45142,N_43540,N_43490);
nand U45143 (N_45143,N_44795,N_43083);
nand U45144 (N_45144,N_42992,N_44271);
xor U45145 (N_45145,N_42844,N_43978);
xnor U45146 (N_45146,N_43865,N_43448);
nand U45147 (N_45147,N_44963,N_44893);
nor U45148 (N_45148,N_44543,N_42648);
or U45149 (N_45149,N_44810,N_44235);
and U45150 (N_45150,N_43194,N_44710);
or U45151 (N_45151,N_44441,N_44331);
nor U45152 (N_45152,N_43393,N_42607);
nand U45153 (N_45153,N_42882,N_44013);
nand U45154 (N_45154,N_44142,N_44561);
xnor U45155 (N_45155,N_44070,N_43964);
xnor U45156 (N_45156,N_44683,N_44410);
and U45157 (N_45157,N_43944,N_43151);
xor U45158 (N_45158,N_44680,N_43212);
xnor U45159 (N_45159,N_44398,N_44180);
xnor U45160 (N_45160,N_43229,N_42679);
and U45161 (N_45161,N_42625,N_44797);
or U45162 (N_45162,N_44817,N_44975);
and U45163 (N_45163,N_44028,N_44239);
and U45164 (N_45164,N_44290,N_44139);
xnor U45165 (N_45165,N_43270,N_43288);
or U45166 (N_45166,N_44949,N_43941);
and U45167 (N_45167,N_42517,N_43668);
and U45168 (N_45168,N_44195,N_44976);
and U45169 (N_45169,N_44511,N_42817);
nor U45170 (N_45170,N_44104,N_43803);
or U45171 (N_45171,N_43059,N_42774);
nor U45172 (N_45172,N_44905,N_44100);
and U45173 (N_45173,N_42640,N_44875);
nor U45174 (N_45174,N_43396,N_43883);
nand U45175 (N_45175,N_44493,N_42771);
and U45176 (N_45176,N_44003,N_43565);
or U45177 (N_45177,N_44279,N_44094);
nand U45178 (N_45178,N_44282,N_44061);
nand U45179 (N_45179,N_43711,N_43898);
nand U45180 (N_45180,N_42563,N_44095);
nand U45181 (N_45181,N_42949,N_43459);
nand U45182 (N_45182,N_44401,N_44662);
nor U45183 (N_45183,N_43388,N_44451);
or U45184 (N_45184,N_44993,N_44008);
nand U45185 (N_45185,N_44951,N_42621);
and U45186 (N_45186,N_43736,N_43422);
nand U45187 (N_45187,N_44078,N_44794);
xnor U45188 (N_45188,N_43037,N_43918);
or U45189 (N_45189,N_42513,N_43237);
and U45190 (N_45190,N_42741,N_42860);
xnor U45191 (N_45191,N_43554,N_44631);
xnor U45192 (N_45192,N_42620,N_44501);
xnor U45193 (N_45193,N_43132,N_43182);
nand U45194 (N_45194,N_44395,N_42695);
or U45195 (N_45195,N_44160,N_42820);
nor U45196 (N_45196,N_42880,N_43579);
nor U45197 (N_45197,N_43432,N_42677);
or U45198 (N_45198,N_44033,N_43553);
xor U45199 (N_45199,N_44169,N_44345);
nor U45200 (N_45200,N_44011,N_42777);
or U45201 (N_45201,N_42518,N_43595);
or U45202 (N_45202,N_44133,N_43491);
and U45203 (N_45203,N_43107,N_42605);
xnor U45204 (N_45204,N_44128,N_44707);
or U45205 (N_45205,N_43773,N_43022);
nor U45206 (N_45206,N_42783,N_43390);
nand U45207 (N_45207,N_42705,N_44804);
nand U45208 (N_45208,N_44754,N_43933);
nand U45209 (N_45209,N_43906,N_44243);
nand U45210 (N_45210,N_43777,N_43454);
xnor U45211 (N_45211,N_42903,N_44121);
xnor U45212 (N_45212,N_44487,N_44537);
xnor U45213 (N_45213,N_42547,N_43904);
nand U45214 (N_45214,N_43881,N_44521);
or U45215 (N_45215,N_43814,N_43992);
nor U45216 (N_45216,N_43258,N_44961);
or U45217 (N_45217,N_42708,N_44332);
and U45218 (N_45218,N_42938,N_43843);
xor U45219 (N_45219,N_42769,N_43702);
nor U45220 (N_45220,N_43669,N_43257);
nor U45221 (N_45221,N_44369,N_42641);
nand U45222 (N_45222,N_42937,N_42678);
or U45223 (N_45223,N_42651,N_43852);
or U45224 (N_45224,N_43884,N_44148);
or U45225 (N_45225,N_44765,N_44067);
nor U45226 (N_45226,N_43122,N_44343);
and U45227 (N_45227,N_42656,N_44602);
nor U45228 (N_45228,N_44069,N_43223);
xnor U45229 (N_45229,N_43729,N_42653);
and U45230 (N_45230,N_44803,N_44528);
nor U45231 (N_45231,N_44314,N_44519);
nand U45232 (N_45232,N_44416,N_44620);
nor U45233 (N_45233,N_44355,N_42838);
or U45234 (N_45234,N_44582,N_42514);
xor U45235 (N_45235,N_43546,N_43382);
nand U45236 (N_45236,N_44920,N_43079);
nand U45237 (N_45237,N_43682,N_44604);
nor U45238 (N_45238,N_44305,N_42520);
xor U45239 (N_45239,N_42675,N_43611);
or U45240 (N_45240,N_44157,N_43937);
or U45241 (N_45241,N_42858,N_43834);
xnor U45242 (N_45242,N_44168,N_43536);
nor U45243 (N_45243,N_43739,N_42580);
nand U45244 (N_45244,N_43518,N_43612);
or U45245 (N_45245,N_43139,N_42558);
xnor U45246 (N_45246,N_44285,N_43244);
xnor U45247 (N_45247,N_43191,N_44945);
or U45248 (N_45248,N_44845,N_43202);
xnor U45249 (N_45249,N_43146,N_44868);
or U45250 (N_45250,N_43586,N_43281);
or U45251 (N_45251,N_42715,N_42642);
nand U45252 (N_45252,N_42849,N_43339);
xnor U45253 (N_45253,N_44498,N_43126);
nor U45254 (N_45254,N_43757,N_44014);
nand U45255 (N_45255,N_44346,N_44468);
nor U45256 (N_45256,N_44642,N_44651);
nor U45257 (N_45257,N_43189,N_44820);
and U45258 (N_45258,N_42968,N_44872);
nor U45259 (N_45259,N_43813,N_44058);
and U45260 (N_45260,N_42790,N_43080);
nand U45261 (N_45261,N_42590,N_44015);
xor U45262 (N_45262,N_44943,N_44788);
nor U45263 (N_45263,N_44350,N_44172);
nor U45264 (N_45264,N_44218,N_44671);
and U45265 (N_45265,N_43063,N_42659);
or U45266 (N_45266,N_43179,N_44075);
nand U45267 (N_45267,N_43372,N_44135);
or U45268 (N_45268,N_44956,N_43562);
xnor U45269 (N_45269,N_44673,N_43001);
nand U45270 (N_45270,N_42980,N_42505);
and U45271 (N_45271,N_42924,N_44841);
nor U45272 (N_45272,N_44771,N_44917);
and U45273 (N_45273,N_44586,N_43507);
xor U45274 (N_45274,N_44276,N_44391);
nor U45275 (N_45275,N_42951,N_43042);
or U45276 (N_45276,N_43822,N_43156);
nand U45277 (N_45277,N_43936,N_43705);
xnor U45278 (N_45278,N_44277,N_42784);
and U45279 (N_45279,N_42919,N_42909);
xor U45280 (N_45280,N_43477,N_44205);
nand U45281 (N_45281,N_42527,N_44258);
and U45282 (N_45282,N_43945,N_44857);
or U45283 (N_45283,N_42538,N_43890);
or U45284 (N_45284,N_43209,N_43916);
xnor U45285 (N_45285,N_44645,N_43867);
xor U45286 (N_45286,N_44293,N_44776);
nor U45287 (N_45287,N_43053,N_42841);
and U45288 (N_45288,N_43561,N_44221);
nor U45289 (N_45289,N_44546,N_42728);
and U45290 (N_45290,N_44781,N_43529);
xnor U45291 (N_45291,N_44783,N_43889);
nand U45292 (N_45292,N_43527,N_44286);
and U45293 (N_45293,N_44392,N_44220);
or U45294 (N_45294,N_44456,N_43555);
nand U45295 (N_45295,N_42837,N_44608);
or U45296 (N_45296,N_43038,N_44213);
nor U45297 (N_45297,N_44162,N_44127);
xor U45298 (N_45298,N_42516,N_43505);
xor U45299 (N_45299,N_42624,N_43046);
or U45300 (N_45300,N_42528,N_42916);
xnor U45301 (N_45301,N_43789,N_43450);
or U45302 (N_45302,N_44533,N_44752);
xnor U45303 (N_45303,N_43954,N_43248);
nand U45304 (N_45304,N_43817,N_44869);
nor U45305 (N_45305,N_44633,N_44903);
and U45306 (N_45306,N_43537,N_42818);
nor U45307 (N_45307,N_42706,N_44494);
nor U45308 (N_45308,N_44508,N_42638);
nand U45309 (N_45309,N_43263,N_43551);
nor U45310 (N_45310,N_42645,N_42848);
nand U45311 (N_45311,N_44840,N_43175);
nand U45312 (N_45312,N_44571,N_44137);
and U45313 (N_45313,N_43780,N_42554);
and U45314 (N_45314,N_43220,N_44698);
or U45315 (N_45315,N_42985,N_44774);
nor U45316 (N_45316,N_44726,N_43262);
nand U45317 (N_45317,N_43580,N_44315);
and U45318 (N_45318,N_44677,N_43280);
or U45319 (N_45319,N_43605,N_44040);
nand U45320 (N_45320,N_44834,N_43602);
xor U45321 (N_45321,N_44916,N_42933);
xnor U45322 (N_45322,N_42816,N_44912);
or U45323 (N_45323,N_42825,N_42894);
nor U45324 (N_45324,N_44767,N_44304);
nor U45325 (N_45325,N_44706,N_42649);
xnor U45326 (N_45326,N_43246,N_44248);
and U45327 (N_45327,N_44170,N_42597);
nor U45328 (N_45328,N_42874,N_42776);
nand U45329 (N_45329,N_43842,N_42719);
nor U45330 (N_45330,N_44402,N_44686);
nand U45331 (N_45331,N_43243,N_43925);
and U45332 (N_45332,N_42574,N_43261);
nor U45333 (N_45333,N_43828,N_44529);
nor U45334 (N_45334,N_43608,N_42914);
or U45335 (N_45335,N_44227,N_43749);
or U45336 (N_45336,N_44244,N_44340);
xor U45337 (N_45337,N_42976,N_43118);
and U45338 (N_45338,N_43603,N_43667);
nand U45339 (N_45339,N_44027,N_43017);
and U45340 (N_45340,N_42519,N_42503);
nor U45341 (N_45341,N_44714,N_44045);
nand U45342 (N_45342,N_42945,N_44042);
nand U45343 (N_45343,N_44228,N_42930);
and U45344 (N_45344,N_42699,N_43235);
nand U45345 (N_45345,N_44793,N_43703);
nor U45346 (N_45346,N_43236,N_44309);
nor U45347 (N_45347,N_42573,N_43347);
nor U45348 (N_45348,N_43741,N_42911);
xor U45349 (N_45349,N_43888,N_44576);
xor U45350 (N_45350,N_43403,N_44923);
nand U45351 (N_45351,N_43428,N_44382);
and U45352 (N_45352,N_44132,N_42960);
xnor U45353 (N_45353,N_43939,N_44769);
and U45354 (N_45354,N_42724,N_43753);
nor U45355 (N_45355,N_43170,N_43201);
nand U45356 (N_45356,N_43695,N_44921);
xor U45357 (N_45357,N_43102,N_43145);
or U45358 (N_45358,N_43592,N_43307);
xnor U45359 (N_45359,N_43274,N_43147);
xnor U45360 (N_45360,N_44557,N_44470);
nand U45361 (N_45361,N_43055,N_42509);
nor U45362 (N_45362,N_43952,N_42987);
xnor U45363 (N_45363,N_43013,N_43934);
xor U45364 (N_45364,N_44946,N_44570);
xnor U45365 (N_45365,N_43815,N_44445);
or U45366 (N_45366,N_44442,N_42530);
and U45367 (N_45367,N_44530,N_42617);
xor U45368 (N_45368,N_44152,N_43011);
or U45369 (N_45369,N_43335,N_44424);
nand U45370 (N_45370,N_44245,N_44694);
and U45371 (N_45371,N_44165,N_44405);
and U45372 (N_45372,N_43019,N_42670);
nand U45373 (N_45373,N_42959,N_43474);
nor U45374 (N_45374,N_44800,N_42566);
and U45375 (N_45375,N_42515,N_44328);
xnor U45376 (N_45376,N_44230,N_43041);
or U45377 (N_45377,N_43804,N_43610);
or U45378 (N_45378,N_44477,N_42879);
xnor U45379 (N_45379,N_43027,N_43991);
or U45380 (N_45380,N_44775,N_44046);
and U45381 (N_45381,N_44705,N_42834);
and U45382 (N_45382,N_43530,N_44667);
or U45383 (N_45383,N_42756,N_42685);
nand U45384 (N_45384,N_44194,N_44373);
nor U45385 (N_45385,N_43091,N_44174);
xnor U45386 (N_45386,N_42668,N_43143);
or U45387 (N_45387,N_44614,N_43097);
and U45388 (N_45388,N_42901,N_43446);
xnor U45389 (N_45389,N_43137,N_44777);
or U45390 (N_45390,N_42793,N_43835);
or U45391 (N_45391,N_42644,N_44336);
nor U45392 (N_45392,N_42990,N_44634);
xnor U45393 (N_45393,N_43453,N_43574);
nand U45394 (N_45394,N_43955,N_43868);
nor U45395 (N_45395,N_44550,N_42895);
or U45396 (N_45396,N_44461,N_44032);
or U45397 (N_45397,N_44755,N_44187);
nand U45398 (N_45398,N_43387,N_44272);
and U45399 (N_45399,N_43242,N_44377);
nand U45400 (N_45400,N_44080,N_42947);
and U45401 (N_45401,N_44291,N_42866);
nor U45402 (N_45402,N_43348,N_43654);
nor U45403 (N_45403,N_43217,N_42955);
xnor U45404 (N_45404,N_43128,N_43167);
xnor U45405 (N_45405,N_43320,N_43962);
xnor U45406 (N_45406,N_44646,N_42940);
nand U45407 (N_45407,N_44181,N_44721);
nand U45408 (N_45408,N_43926,N_44471);
xor U45409 (N_45409,N_44520,N_44815);
and U45410 (N_45410,N_43104,N_42592);
and U45411 (N_45411,N_43833,N_44575);
nand U45412 (N_45412,N_44644,N_44001);
or U45413 (N_45413,N_42855,N_43839);
xnor U45414 (N_45414,N_43696,N_43370);
or U45415 (N_45415,N_44363,N_42815);
xnor U45416 (N_45416,N_43853,N_44757);
nand U45417 (N_45417,N_43411,N_43986);
or U45418 (N_45418,N_44122,N_43742);
xnor U45419 (N_45419,N_44255,N_43628);
nand U45420 (N_45420,N_42754,N_44526);
nor U45421 (N_45421,N_44407,N_43043);
and U45422 (N_45422,N_42843,N_44558);
nand U45423 (N_45423,N_43328,N_42525);
and U45424 (N_45424,N_42956,N_44097);
nor U45425 (N_45425,N_44068,N_44855);
nand U45426 (N_45426,N_43358,N_44966);
xnor U45427 (N_45427,N_44199,N_44611);
or U45428 (N_45428,N_43052,N_44223);
and U45429 (N_45429,N_43599,N_43114);
or U45430 (N_45430,N_44450,N_44136);
nor U45431 (N_45431,N_42714,N_43629);
xnor U45432 (N_45432,N_42686,N_42546);
nor U45433 (N_45433,N_42552,N_42821);
or U45434 (N_45434,N_44171,N_43829);
xnor U45435 (N_45435,N_42740,N_44310);
nor U45436 (N_45436,N_44692,N_43726);
nor U45437 (N_45437,N_43002,N_44761);
xor U45438 (N_45438,N_43718,N_43830);
and U45439 (N_45439,N_43624,N_43412);
nor U45440 (N_45440,N_44832,N_44762);
nor U45441 (N_45441,N_42702,N_43334);
or U45442 (N_45442,N_44647,N_44338);
nand U45443 (N_45443,N_43979,N_43299);
or U45444 (N_45444,N_43066,N_44531);
nand U45445 (N_45445,N_42587,N_43982);
or U45446 (N_45446,N_44837,N_43313);
and U45447 (N_45447,N_43528,N_43073);
xnor U45448 (N_45448,N_44906,N_44863);
and U45449 (N_45449,N_43784,N_42845);
nor U45450 (N_45450,N_42755,N_43030);
xor U45451 (N_45451,N_43287,N_44703);
or U45452 (N_45452,N_43976,N_43371);
nor U45453 (N_45453,N_43871,N_43015);
nor U45454 (N_45454,N_44635,N_42787);
nor U45455 (N_45455,N_44584,N_43385);
or U45456 (N_45456,N_43756,N_43375);
nor U45457 (N_45457,N_44431,N_42602);
and U45458 (N_45458,N_43207,N_44742);
nand U45459 (N_45459,N_43481,N_44610);
xnor U45460 (N_45460,N_43910,N_44348);
and U45461 (N_45461,N_44770,N_42671);
or U45462 (N_45462,N_43509,N_43514);
nor U45463 (N_45463,N_43214,N_43275);
nor U45464 (N_45464,N_43819,N_44658);
or U45465 (N_45465,N_43870,N_42803);
nor U45466 (N_45466,N_42562,N_43425);
xor U45467 (N_45467,N_44836,N_43402);
or U45468 (N_45468,N_44785,N_44831);
nand U45469 (N_45469,N_44274,N_43269);
nor U45470 (N_45470,N_44403,N_43078);
nand U45471 (N_45471,N_44016,N_43631);
and U45472 (N_45472,N_42775,N_43956);
and U45473 (N_45473,N_44928,N_44466);
xnor U45474 (N_45474,N_42857,N_42900);
xor U45475 (N_45475,N_43095,N_43751);
and U45476 (N_45476,N_44118,N_44544);
and U45477 (N_45477,N_42905,N_42710);
and U45478 (N_45478,N_42681,N_44932);
nor U45479 (N_45479,N_44615,N_43659);
nand U45480 (N_45480,N_42610,N_42704);
and U45481 (N_45481,N_43319,N_42500);
nand U45482 (N_45482,N_44129,N_44994);
nand U45483 (N_45483,N_44161,N_44732);
xor U45484 (N_45484,N_44661,N_43204);
nand U45485 (N_45485,N_43406,N_44098);
or U45486 (N_45486,N_44263,N_42700);
nor U45487 (N_45487,N_43101,N_44556);
and U45488 (N_45488,N_42604,N_43632);
or U45489 (N_45489,N_43072,N_44439);
nor U45490 (N_45490,N_44091,N_43501);
nand U45491 (N_45491,N_43301,N_43305);
nand U45492 (N_45492,N_43919,N_42762);
and U45493 (N_45493,N_44084,N_42585);
nor U45494 (N_45494,N_43915,N_43677);
and U45495 (N_45495,N_43524,N_43254);
nand U45496 (N_45496,N_42745,N_44989);
nor U45497 (N_45497,N_44394,N_44265);
nor U45498 (N_45498,N_43932,N_42779);
xor U45499 (N_45499,N_43811,N_44819);
and U45500 (N_45500,N_43451,N_43764);
nand U45501 (N_45501,N_44693,N_43533);
and U45502 (N_45502,N_42615,N_43965);
and U45503 (N_45503,N_44603,N_44105);
xnor U45504 (N_45504,N_44539,N_42512);
nor U45505 (N_45505,N_42564,N_43180);
or U45506 (N_45506,N_44830,N_44948);
xnor U45507 (N_45507,N_43134,N_43731);
xnor U45508 (N_45508,N_44965,N_42723);
xnor U45509 (N_45509,N_43449,N_44835);
xnor U45510 (N_45510,N_44376,N_44596);
xor U45511 (N_45511,N_43727,N_42993);
nor U45512 (N_45512,N_42898,N_43460);
xnor U45513 (N_45513,N_43846,N_44882);
xor U45514 (N_45514,N_43178,N_44739);
xnor U45515 (N_45515,N_44478,N_44950);
and U45516 (N_45516,N_43700,N_44753);
xnor U45517 (N_45517,N_43210,N_42764);
xnor U45518 (N_45518,N_44452,N_42526);
xor U45519 (N_45519,N_44256,N_43989);
nor U45520 (N_45520,N_44799,N_43231);
nor U45521 (N_45521,N_44904,N_43276);
and U45522 (N_45522,N_44208,N_43570);
nand U45523 (N_45523,N_43559,N_43855);
nor U45524 (N_45524,N_42545,N_43443);
and U45525 (N_45525,N_43153,N_42923);
nor U45526 (N_45526,N_42922,N_44959);
xnor U45527 (N_45527,N_43050,N_42694);
xnor U45528 (N_45528,N_44476,N_44113);
and U45529 (N_45529,N_44178,N_43476);
xnor U45530 (N_45530,N_42984,N_44495);
nor U45531 (N_45531,N_43340,N_43300);
and U45532 (N_45532,N_44063,N_43531);
or U45533 (N_45533,N_43238,N_43085);
and U45534 (N_45534,N_42798,N_43787);
and U45535 (N_45535,N_44209,N_43892);
nand U45536 (N_45536,N_44126,N_43192);
or U45537 (N_45537,N_44010,N_44702);
and U45538 (N_45538,N_44572,N_43931);
xor U45539 (N_45539,N_42565,N_44787);
xor U45540 (N_45540,N_43818,N_44850);
xnor U45541 (N_45541,N_42983,N_43457);
xor U45542 (N_45542,N_44648,N_43508);
nand U45543 (N_45543,N_43566,N_44992);
nor U45544 (N_45544,N_43755,N_43226);
nand U45545 (N_45545,N_43322,N_43172);
nor U45546 (N_45546,N_43999,N_43557);
or U45547 (N_45547,N_44418,N_43003);
or U45548 (N_45548,N_43643,N_44469);
nand U45549 (N_45549,N_42995,N_44353);
nor U45550 (N_45550,N_42807,N_42556);
nor U45551 (N_45551,N_43051,N_42543);
and U45552 (N_45552,N_44432,N_43401);
nor U45553 (N_45553,N_43966,N_44908);
or U45554 (N_45554,N_44510,N_43032);
nor U45555 (N_45555,N_44577,N_43029);
and U45556 (N_45556,N_44592,N_43308);
xor U45557 (N_45557,N_43893,N_43935);
and U45558 (N_45558,N_44744,N_43639);
nand U45559 (N_45559,N_44627,N_42941);
nand U45560 (N_45560,N_43882,N_44086);
or U45561 (N_45561,N_43740,N_42634);
xor U45562 (N_45562,N_43851,N_44759);
nor U45563 (N_45563,N_42584,N_44918);
nand U45564 (N_45564,N_44434,N_43381);
nand U45565 (N_45565,N_43470,N_44878);
xnor U45566 (N_45566,N_44192,N_43856);
and U45567 (N_45567,N_43325,N_44050);
and U45568 (N_45568,N_42805,N_44052);
xor U45569 (N_45569,N_42981,N_43805);
or U45570 (N_45570,N_44238,N_42982);
nand U45571 (N_45571,N_43268,N_43351);
nor U45572 (N_45572,N_44047,N_43373);
xnor U45573 (N_45573,N_44987,N_43495);
xor U45574 (N_45574,N_43665,N_43823);
or U45575 (N_45575,N_44983,N_43464);
and U45576 (N_45576,N_43215,N_42859);
xnor U45577 (N_45577,N_43277,N_43312);
nor U45578 (N_45578,N_44430,N_43049);
nand U45579 (N_45579,N_44599,N_43583);
nor U45580 (N_45580,N_44138,N_43009);
and U45581 (N_45581,N_43368,N_42647);
nand U45582 (N_45582,N_44682,N_43316);
or U45583 (N_45583,N_43544,N_43136);
and U45584 (N_45584,N_43959,N_43329);
nand U45585 (N_45585,N_44283,N_43768);
and U45586 (N_45586,N_44833,N_44907);
nor U45587 (N_45587,N_43149,N_44140);
and U45588 (N_45588,N_44490,N_44231);
and U45589 (N_45589,N_43827,N_44360);
nor U45590 (N_45590,N_44609,N_43563);
nand U45591 (N_45591,N_43200,N_44257);
and U45592 (N_45592,N_43975,N_44624);
nor U45593 (N_45593,N_43970,N_44653);
nor U45594 (N_45594,N_43186,N_42603);
and U45595 (N_45595,N_44268,N_42827);
nor U45596 (N_45596,N_43604,N_43427);
and U45597 (N_45597,N_44896,N_44297);
and U45598 (N_45598,N_44625,N_43674);
and U45599 (N_45599,N_42977,N_42720);
and U45600 (N_45600,N_43649,N_42734);
and U45601 (N_45601,N_44039,N_42536);
nor U45602 (N_45602,N_44399,N_43591);
nor U45603 (N_45603,N_43832,N_43206);
xor U45604 (N_45604,N_43008,N_42633);
xnor U45605 (N_45605,N_44999,N_42885);
or U45606 (N_45606,N_43400,N_42760);
or U45607 (N_45607,N_43249,N_44666);
nand U45608 (N_45608,N_44370,N_44201);
nor U45609 (N_45609,N_44630,N_42800);
nand U45610 (N_45610,N_44766,N_42537);
xnor U45611 (N_45611,N_43737,N_44930);
nand U45612 (N_45612,N_43875,N_44491);
nand U45613 (N_45613,N_42583,N_42778);
nor U45614 (N_45614,N_44619,N_43199);
nor U45615 (N_45615,N_44967,N_44981);
and U45616 (N_45616,N_42888,N_42806);
nor U45617 (N_45617,N_43743,N_43719);
xnor U45618 (N_45618,N_43721,N_44085);
xor U45619 (N_45619,N_42680,N_42867);
nor U45620 (N_45620,N_42731,N_44186);
or U45621 (N_45621,N_44891,N_43098);
nand U45622 (N_45622,N_43241,N_43426);
nand U45623 (N_45623,N_43294,N_44179);
nand U45624 (N_45624,N_43100,N_44798);
nand U45625 (N_45625,N_43532,N_43560);
xor U45626 (N_45626,N_43369,N_44202);
nor U45627 (N_45627,N_44554,N_44232);
nand U45628 (N_45628,N_42618,N_42643);
or U45629 (N_45629,N_43651,N_42865);
nand U45630 (N_45630,N_44106,N_44347);
xnor U45631 (N_45631,N_43500,N_43625);
and U45632 (N_45632,N_44387,N_43093);
nor U45633 (N_45633,N_43809,N_44141);
and U45634 (N_45634,N_44087,N_44621);
nor U45635 (N_45635,N_44433,N_43543);
xor U45636 (N_45636,N_44362,N_42887);
nand U45637 (N_45637,N_43445,N_43957);
xor U45638 (N_45638,N_44089,N_43161);
and U45639 (N_45639,N_44643,N_44167);
nor U45640 (N_45640,N_43311,N_44422);
and U45641 (N_45641,N_44200,N_42629);
xnor U45642 (N_45642,N_44024,N_43894);
xor U45643 (N_45643,N_44375,N_44482);
nor U45644 (N_45644,N_43473,N_44119);
or U45645 (N_45645,N_44874,N_43801);
nor U45646 (N_45646,N_42501,N_44182);
or U45647 (N_45647,N_44261,N_44190);
xor U45648 (N_45648,N_43928,N_43293);
xnor U45649 (N_45649,N_43825,N_44583);
nand U45650 (N_45650,N_42689,N_43572);
nor U45651 (N_45651,N_43005,N_44125);
nand U45652 (N_45652,N_42835,N_44019);
or U45653 (N_45653,N_44859,N_43399);
nand U45654 (N_45654,N_43264,N_43636);
and U45655 (N_45655,N_44251,N_43671);
xnor U45656 (N_45656,N_43462,N_42920);
and U45657 (N_45657,N_44492,N_42964);
nor U45658 (N_45658,N_44613,N_43359);
and U45659 (N_45659,N_43247,N_44545);
xor U45660 (N_45660,N_43020,N_42511);
xnor U45661 (N_45661,N_43271,N_43745);
xor U45662 (N_45662,N_42535,N_44158);
and U45663 (N_45663,N_44517,N_43549);
and U45664 (N_45664,N_43732,N_42846);
nand U45665 (N_45665,N_44688,N_44307);
or U45666 (N_45666,N_42541,N_43361);
xor U45667 (N_45667,N_44738,N_43950);
nor U45668 (N_45668,N_43584,N_44485);
nand U45669 (N_45669,N_43398,N_42549);
nand U45670 (N_45670,N_43034,N_43203);
nand U45671 (N_45671,N_43848,N_43849);
or U45672 (N_45672,N_43407,N_43708);
or U45673 (N_45673,N_43039,N_44018);
nor U45674 (N_45674,N_44017,N_44598);
or U45675 (N_45675,N_43921,N_44843);
xor U45676 (N_45676,N_44404,N_43346);
xnor U45677 (N_45677,N_44972,N_42504);
xor U45678 (N_45678,N_43297,N_43324);
or U45679 (N_45679,N_43309,N_44060);
xor U45680 (N_45680,N_43769,N_42736);
xnor U45681 (N_45681,N_44318,N_44124);
nand U45682 (N_45682,N_44108,N_43800);
nand U45683 (N_45683,N_43060,N_44145);
nand U45684 (N_45684,N_44327,N_42890);
or U45685 (N_45685,N_44851,N_44448);
nor U45686 (N_45686,N_42540,N_44388);
xor U45687 (N_45687,N_43973,N_44746);
or U45688 (N_45688,N_44701,N_44789);
xnor U45689 (N_45689,N_43125,N_43902);
or U45690 (N_45690,N_44720,N_43655);
and U45691 (N_45691,N_43023,N_42507);
nor U45692 (N_45692,N_44587,N_44654);
nand U45693 (N_45693,N_43863,N_43995);
nor U45694 (N_45694,N_43227,N_43338);
and U45695 (N_45695,N_42998,N_42593);
and U45696 (N_45696,N_44581,N_44926);
and U45697 (N_45697,N_43000,N_43071);
nor U45698 (N_45698,N_44735,N_42661);
nand U45699 (N_45699,N_43901,N_44749);
xor U45700 (N_45700,N_43573,N_43692);
nand U45701 (N_45701,N_43517,N_44616);
nand U45702 (N_45702,N_43113,N_43230);
nor U45703 (N_45703,N_44737,N_42948);
nand U45704 (N_45704,N_44734,N_43345);
xor U45705 (N_45705,N_44656,N_44728);
or U45706 (N_45706,N_42524,N_44839);
or U45707 (N_45707,N_44083,N_42703);
or U45708 (N_45708,N_43240,N_44449);
xnor U45709 (N_45709,N_44374,N_44718);
or U45710 (N_45710,N_43420,N_44724);
nor U45711 (N_45711,N_44234,N_43971);
or U45712 (N_45712,N_44185,N_42799);
nor U45713 (N_45713,N_43810,N_44861);
or U45714 (N_45714,N_44871,N_42646);
xnor U45715 (N_45715,N_44573,N_44727);
nand U45716 (N_45716,N_43593,N_43010);
or U45717 (N_45717,N_44457,N_42852);
or U45718 (N_45718,N_43292,N_44591);
nand U45719 (N_45719,N_44629,N_43131);
and U45720 (N_45720,N_42658,N_42662);
nor U45721 (N_45721,N_43845,N_43774);
nor U45722 (N_45722,N_44823,N_43163);
or U45723 (N_45723,N_42966,N_44267);
or U45724 (N_45724,N_43903,N_44206);
nor U45725 (N_45725,N_42749,N_44484);
nand U45726 (N_45726,N_43609,N_43314);
nor U45727 (N_45727,N_43502,N_43333);
or U45728 (N_45728,N_43791,N_44415);
xor U45729 (N_45729,N_42869,N_44973);
and U45730 (N_45730,N_44249,N_43526);
nand U45731 (N_45731,N_44219,N_44203);
and U45732 (N_45732,N_43511,N_43211);
nor U45733 (N_45733,N_44116,N_43064);
and U45734 (N_45734,N_44709,N_43746);
nand U45735 (N_45735,N_42893,N_44323);
xnor U45736 (N_45736,N_42994,N_44412);
or U45737 (N_45737,N_43456,N_43874);
nand U45738 (N_45738,N_44472,N_44365);
or U45739 (N_45739,N_44246,N_43614);
and U45740 (N_45740,N_43441,N_43758);
nor U45741 (N_45741,N_42780,N_42839);
nand U45742 (N_45742,N_44072,N_43488);
nand U45743 (N_45743,N_43065,N_44386);
or U45744 (N_45744,N_43352,N_43601);
nor U45745 (N_45745,N_42954,N_42650);
nor U45746 (N_45746,N_44156,N_43479);
nand U45747 (N_45747,N_44821,N_43681);
nor U45748 (N_45748,N_42690,N_43648);
nand U45749 (N_45749,N_42850,N_43968);
nor U45750 (N_45750,N_43837,N_44499);
nor U45751 (N_45751,N_43613,N_43618);
nand U45752 (N_45752,N_44034,N_43983);
nor U45753 (N_45753,N_42730,N_43033);
or U45754 (N_45754,N_44154,N_43045);
nor U45755 (N_45755,N_42763,N_44480);
and U45756 (N_45756,N_43776,N_43343);
or U45757 (N_45757,N_44417,N_44927);
and U45758 (N_45758,N_43525,N_44953);
and U45759 (N_45759,N_44899,N_42896);
nor U45760 (N_45760,N_42692,N_44814);
xnor U45761 (N_45761,N_44111,N_42718);
nand U45762 (N_45762,N_44566,N_43306);
or U45763 (N_45763,N_42596,N_43878);
nor U45764 (N_45764,N_44312,N_43656);
xor U45765 (N_45765,N_43196,N_44163);
nor U45766 (N_45766,N_44296,N_43154);
xnor U45767 (N_45767,N_44044,N_43571);
and U45768 (N_45768,N_44516,N_43492);
xor U45769 (N_45769,N_44313,N_44311);
nand U45770 (N_45770,N_43841,N_43321);
or U45771 (N_45771,N_44065,N_43940);
and U45772 (N_45772,N_42926,N_43850);
or U45773 (N_45773,N_43585,N_42688);
or U45774 (N_45774,N_44035,N_44514);
nor U45775 (N_45775,N_43626,N_42707);
nor U45776 (N_45776,N_44877,N_42770);
or U45777 (N_45777,N_43647,N_43225);
or U45778 (N_45778,N_42819,N_44969);
xor U45779 (N_45779,N_42600,N_43640);
or U45780 (N_45780,N_43658,N_43596);
and U45781 (N_45781,N_44540,N_44004);
xnor U45782 (N_45782,N_44699,N_44684);
or U45783 (N_45783,N_43213,N_42716);
or U45784 (N_45784,N_44847,N_44802);
and U45785 (N_45785,N_43088,N_42586);
and U45786 (N_45786,N_44023,N_42908);
and U45787 (N_45787,N_44260,N_44411);
and U45788 (N_45788,N_43697,N_44458);
or U45789 (N_45789,N_44942,N_44278);
nand U45790 (N_45790,N_42601,N_44210);
or U45791 (N_45791,N_44224,N_43461);
nor U45792 (N_45792,N_44381,N_44030);
or U45793 (N_45793,N_44173,N_43442);
or U45794 (N_45794,N_44664,N_43541);
and U45795 (N_45795,N_42917,N_42808);
xnor U45796 (N_45796,N_43440,N_44284);
xnor U45797 (N_45797,N_42973,N_44130);
nand U45798 (N_45798,N_43598,N_43535);
or U45799 (N_45799,N_43298,N_42752);
nor U45800 (N_45800,N_44455,N_43188);
or U45801 (N_45801,N_43478,N_43483);
nor U45802 (N_45802,N_43123,N_42608);
nor U45803 (N_45803,N_43356,N_44475);
xor U45804 (N_45804,N_43405,N_43155);
nor U45805 (N_45805,N_44560,N_44057);
nor U45806 (N_45806,N_44866,N_43550);
and U45807 (N_45807,N_44924,N_44211);
xor U45808 (N_45808,N_43963,N_42544);
xor U45809 (N_45809,N_44773,N_43067);
and U45810 (N_45810,N_43891,N_43389);
or U45811 (N_45811,N_42637,N_43723);
xor U45812 (N_45812,N_43545,N_44419);
nand U45813 (N_45813,N_43621,N_42567);
or U45814 (N_45814,N_44884,N_44266);
nor U45815 (N_45815,N_43802,N_44406);
nor U45816 (N_45816,N_44955,N_44049);
or U45817 (N_45817,N_43089,N_43397);
and U45818 (N_45818,N_44222,N_42814);
and U45819 (N_45819,N_42877,N_43234);
nand U45820 (N_45820,N_43523,N_43510);
nand U45821 (N_45821,N_43896,N_44901);
or U45822 (N_45822,N_43062,N_44867);
and U45823 (N_45823,N_43516,N_44748);
or U45824 (N_45824,N_42575,N_42974);
nor U45825 (N_45825,N_43710,N_44713);
xor U45826 (N_45826,N_44786,N_43272);
nor U45827 (N_45827,N_44504,N_43357);
or U45828 (N_45828,N_44096,N_42871);
nor U45829 (N_45829,N_44565,N_43998);
nor U45830 (N_45830,N_43635,N_43859);
nor U45831 (N_45831,N_44479,N_44897);
and U45832 (N_45832,N_42691,N_43392);
and U45833 (N_45833,N_44881,N_43606);
nor U45834 (N_45834,N_44676,N_42928);
xor U45835 (N_45835,N_43862,N_43286);
or U45836 (N_45836,N_42627,N_43866);
or U45837 (N_45837,N_44502,N_44062);
and U45838 (N_45838,N_42768,N_43251);
and U45839 (N_45839,N_43577,N_44214);
or U45840 (N_45840,N_44697,N_42663);
xnor U45841 (N_45841,N_44562,N_42673);
nor U45842 (N_45842,N_44600,N_43960);
xnor U45843 (N_45843,N_44048,N_43061);
xor U45844 (N_45844,N_43337,N_42892);
nor U45845 (N_45845,N_42664,N_43716);
nor U45846 (N_45846,N_43408,N_43438);
xor U45847 (N_45847,N_44535,N_44240);
nand U45848 (N_45848,N_43657,N_43984);
nand U45849 (N_45849,N_42582,N_44957);
xor U45850 (N_45850,N_44894,N_43987);
or U45851 (N_45851,N_44880,N_44150);
or U45852 (N_45852,N_44597,N_44623);
or U45853 (N_45853,N_43162,N_44326);
or U45854 (N_45854,N_42813,N_44844);
and U45855 (N_45855,N_42872,N_43109);
and U45856 (N_45856,N_43860,N_44435);
and U45857 (N_45857,N_44637,N_44719);
and U45858 (N_45858,N_42801,N_42672);
or U45859 (N_45859,N_44532,N_44425);
nand U45860 (N_45860,N_44826,N_43734);
nand U45861 (N_45861,N_43786,N_44371);
xnor U45862 (N_45862,N_44460,N_42788);
and U45863 (N_45863,N_44674,N_43429);
nand U45864 (N_45864,N_44229,N_43070);
or U45865 (N_45865,N_43687,N_44302);
and U45866 (N_45866,N_42910,N_42684);
xnor U45867 (N_45867,N_42595,N_44408);
and U45868 (N_45868,N_44295,N_44974);
nand U45869 (N_45869,N_44446,N_44862);
xnor U45870 (N_45870,N_43793,N_44421);
and U45871 (N_45871,N_44379,N_42721);
or U45872 (N_45872,N_43116,N_43619);
or U45873 (N_45873,N_43496,N_42729);
nand U45874 (N_45874,N_43930,N_44077);
xor U45875 (N_45875,N_44670,N_44751);
or U45876 (N_45876,N_44538,N_43219);
and U45877 (N_45877,N_44131,N_43224);
xor U45878 (N_45878,N_43285,N_44088);
xnor U45879 (N_45879,N_42830,N_43142);
or U45880 (N_45880,N_43497,N_42746);
and U45881 (N_45881,N_43183,N_43265);
nand U45882 (N_45882,N_44934,N_42840);
or U45883 (N_45883,N_43824,N_43840);
and U45884 (N_45884,N_44574,N_43082);
or U45885 (N_45885,N_43947,N_44822);
nand U45886 (N_45886,N_43576,N_43086);
nor U45887 (N_45887,N_42761,N_44384);
or U45888 (N_45888,N_44505,N_43377);
nand U45889 (N_45889,N_44101,N_44225);
or U45890 (N_45890,N_43907,N_43946);
nand U45891 (N_45891,N_42810,N_44980);
or U45892 (N_45892,N_43485,N_43515);
nand U45893 (N_45893,N_43688,N_43770);
xor U45894 (N_45894,N_43686,N_42682);
or U45895 (N_45895,N_44808,N_44628);
xnor U45896 (N_45896,N_44784,N_44763);
nand U45897 (N_45897,N_43630,N_42997);
nand U45898 (N_45898,N_43444,N_42942);
and U45899 (N_45899,N_44649,N_43807);
or U45900 (N_45900,N_43808,N_44935);
nand U45901 (N_45901,N_43689,N_43327);
or U45902 (N_45902,N_43341,N_42953);
or U45903 (N_45903,N_44021,N_44895);
or U45904 (N_45904,N_43678,N_44164);
xnor U45905 (N_45905,N_43332,N_42906);
and U45906 (N_45906,N_44846,N_43548);
nor U45907 (N_45907,N_43007,N_42652);
and U45908 (N_45908,N_43912,N_44842);
nand U45909 (N_45909,N_44301,N_44396);
or U45910 (N_45910,N_44626,N_43569);
nand U45911 (N_45911,N_43433,N_43924);
xnor U45912 (N_45912,N_43836,N_42773);
and U45913 (N_45913,N_44115,N_42962);
and U45914 (N_45914,N_44473,N_43418);
and U45915 (N_45915,N_44944,N_43303);
nand U45916 (N_45916,N_43363,N_43779);
and U45917 (N_45917,N_42571,N_43208);
nor U45918 (N_45918,N_44555,N_44423);
or U45919 (N_45919,N_43058,N_43854);
and U45920 (N_45920,N_42594,N_44962);
or U45921 (N_45921,N_43068,N_44038);
or U45922 (N_45922,N_42832,N_43036);
nor U45923 (N_45923,N_43806,N_43699);
and U45924 (N_45924,N_42986,N_44352);
nand U45925 (N_45925,N_42676,N_44954);
or U45926 (N_45926,N_44650,N_43990);
nor U45927 (N_45927,N_42797,N_43266);
nand U45928 (N_45928,N_44366,N_43121);
nor U45929 (N_45929,N_42598,N_43637);
and U45930 (N_45930,N_44500,N_44372);
nor U45931 (N_45931,N_43012,N_42711);
and U45932 (N_45932,N_43404,N_42899);
and U45933 (N_45933,N_44865,N_44816);
and U45934 (N_45934,N_44593,N_42738);
and U45935 (N_45935,N_44768,N_44005);
nand U45936 (N_45936,N_44443,N_44308);
xnor U45937 (N_45937,N_42713,N_43124);
and U45938 (N_45938,N_44054,N_43318);
and U45939 (N_45939,N_43627,N_44632);
nor U45940 (N_45940,N_44189,N_44103);
and U45941 (N_45941,N_43075,N_43362);
or U45942 (N_45942,N_43475,N_43821);
nor U45943 (N_45943,N_43493,N_43430);
or U45944 (N_45944,N_42576,N_43468);
and U45945 (N_45945,N_44079,N_42589);
or U45946 (N_45946,N_42523,N_43439);
and U45947 (N_45947,N_43909,N_44568);
xor U45948 (N_45948,N_42969,N_44123);
nand U45949 (N_45949,N_43724,N_43766);
nand U45950 (N_45950,N_42570,N_43181);
xnor U45951 (N_45951,N_42609,N_42581);
nand U45952 (N_45952,N_42854,N_43484);
nor U45953 (N_45953,N_44389,N_42932);
xor U45954 (N_45954,N_43953,N_43171);
and U45955 (N_45955,N_43961,N_43798);
or U45956 (N_45956,N_43391,N_43326);
and U45957 (N_45957,N_44911,N_43165);
or U45958 (N_45958,N_43355,N_42836);
nor U45959 (N_45959,N_44678,N_44117);
nor U45960 (N_45960,N_42560,N_43763);
nor U45961 (N_45961,N_44873,N_43680);
xor U45962 (N_45962,N_43701,N_44074);
and U45963 (N_45963,N_43911,N_43016);
nand U45964 (N_45964,N_43195,N_42957);
nor U45965 (N_45965,N_44612,N_43040);
or U45966 (N_45966,N_43069,N_44977);
xnor U45967 (N_45967,N_44483,N_42864);
nor U45968 (N_45968,N_43354,N_44958);
xnor U45969 (N_45969,N_44860,N_44368);
nand U45970 (N_45970,N_43117,N_44191);
nor U45971 (N_45971,N_43331,N_44542);
or U45972 (N_45972,N_44333,N_44736);
nand U45973 (N_45973,N_44212,N_44960);
nor U45974 (N_45974,N_42732,N_43790);
xor U45975 (N_45975,N_44367,N_43232);
or U45976 (N_45976,N_43949,N_42758);
nand U45977 (N_45977,N_44159,N_43707);
or U45978 (N_45978,N_44601,N_44175);
nor U45979 (N_45979,N_44329,N_44758);
nor U45980 (N_45980,N_44507,N_44110);
or U45981 (N_45981,N_42623,N_42531);
nand U45982 (N_45982,N_43157,N_44660);
xnor U45983 (N_45983,N_44890,N_44043);
xnor U45984 (N_45984,N_44870,N_44390);
xor U45985 (N_45985,N_42881,N_42631);
xnor U45986 (N_45986,N_44939,N_43638);
nand U45987 (N_45987,N_42532,N_43886);
and U45988 (N_45988,N_42978,N_42789);
or U45989 (N_45989,N_43252,N_44503);
nor U45990 (N_45990,N_43028,N_42782);
and U45991 (N_45991,N_42950,N_44675);
nand U45992 (N_45992,N_44617,N_42907);
xor U45993 (N_45993,N_42828,N_44522);
xor U45994 (N_45994,N_44324,N_42831);
nand U45995 (N_45995,N_43600,N_42510);
nor U45996 (N_45996,N_44270,N_44782);
and U45997 (N_45997,N_43103,N_43380);
nand U45998 (N_45998,N_43938,N_44467);
nor U45999 (N_45999,N_43698,N_43905);
nor U46000 (N_46000,N_44541,N_44712);
nand U46001 (N_46001,N_44638,N_43315);
xor U46002 (N_46002,N_44447,N_43166);
nand U46003 (N_46003,N_43409,N_43922);
and U46004 (N_46004,N_43534,N_44569);
nor U46005 (N_46005,N_44809,N_44464);
nor U46006 (N_46006,N_44887,N_43383);
nor U46007 (N_46007,N_44553,N_43090);
nor U46008 (N_46008,N_43245,N_43466);
nand U46009 (N_46009,N_44585,N_43284);
nor U46010 (N_46010,N_42804,N_43144);
and U46011 (N_46011,N_43895,N_44636);
xor U46012 (N_46012,N_43415,N_43706);
or U46013 (N_46013,N_42934,N_44919);
nor U46014 (N_46014,N_42696,N_44512);
nor U46015 (N_46015,N_44829,N_43504);
xnor U46016 (N_46016,N_44729,N_42861);
and U46017 (N_46017,N_42802,N_43914);
and U46018 (N_46018,N_44828,N_43767);
nand U46019 (N_46019,N_42693,N_44548);
nand U46020 (N_46020,N_42826,N_42915);
nand U46021 (N_46021,N_43106,N_44143);
xor U46022 (N_46022,N_42654,N_42709);
or U46023 (N_46023,N_44076,N_44254);
and U46024 (N_46024,N_43413,N_44151);
or U46025 (N_46025,N_42842,N_42785);
and U46026 (N_46026,N_43712,N_43350);
nand U46027 (N_46027,N_44848,N_43353);
and U46028 (N_46028,N_43349,N_44081);
and U46029 (N_46029,N_44436,N_44813);
nand U46030 (N_46030,N_42577,N_42534);
nor U46031 (N_46031,N_44790,N_43857);
nor U46032 (N_46032,N_44687,N_44925);
nand U46033 (N_46033,N_44059,N_44595);
nor U46034 (N_46034,N_44474,N_44320);
xnor U46035 (N_46035,N_42725,N_44319);
and U46036 (N_46036,N_43958,N_43617);
nor U46037 (N_46037,N_44740,N_42588);
nor U46038 (N_46038,N_44856,N_43728);
or U46039 (N_46039,N_44715,N_43386);
and U46040 (N_46040,N_44700,N_44364);
or U46041 (N_46041,N_44964,N_42975);
nand U46042 (N_46042,N_42701,N_43077);
xor U46043 (N_46043,N_44031,N_44029);
nor U46044 (N_46044,N_42822,N_42559);
nor U46045 (N_46045,N_44525,N_44594);
nor U46046 (N_46046,N_44952,N_43943);
or U46047 (N_46047,N_42506,N_43969);
nor U46048 (N_46048,N_44931,N_44589);
or U46049 (N_46049,N_44454,N_44380);
nand U46050 (N_46050,N_42809,N_42902);
nor U46051 (N_46051,N_42533,N_44289);
nor U46052 (N_46052,N_43747,N_43168);
nor U46053 (N_46053,N_43081,N_44580);
nor U46054 (N_46054,N_44779,N_42622);
xnor U46055 (N_46055,N_44262,N_42876);
and U46056 (N_46056,N_43997,N_44708);
xnor U46057 (N_46057,N_42614,N_44995);
and U46058 (N_46058,N_44996,N_44006);
or U46059 (N_46059,N_43714,N_42868);
and U46060 (N_46060,N_43634,N_42912);
nand U46061 (N_46061,N_42796,N_43519);
or U46062 (N_46062,N_42568,N_44796);
nor U46063 (N_46063,N_44236,N_42786);
and U46064 (N_46064,N_42935,N_44997);
or U46065 (N_46065,N_44811,N_44226);
nand U46066 (N_46066,N_43913,N_42683);
nor U46067 (N_46067,N_42961,N_43498);
or U46068 (N_46068,N_44655,N_42767);
nand U46069 (N_46069,N_44073,N_42508);
nand U46070 (N_46070,N_42989,N_44933);
and U46071 (N_46071,N_42952,N_44242);
and U46072 (N_46072,N_44536,N_43419);
and U46073 (N_46073,N_44898,N_44337);
nor U46074 (N_46074,N_43645,N_42639);
nand U46075 (N_46075,N_42847,N_44275);
xnor U46076 (N_46076,N_43503,N_44306);
nand U46077 (N_46077,N_43980,N_43365);
or U46078 (N_46078,N_44147,N_43342);
nand U46079 (N_46079,N_42765,N_43054);
nor U46080 (N_46080,N_43722,N_43993);
nor U46081 (N_46081,N_43317,N_42757);
xnor U46082 (N_46082,N_43666,N_44427);
and U46083 (N_46083,N_42967,N_44579);
nand U46084 (N_46084,N_43622,N_43228);
xor U46085 (N_46085,N_43176,N_44778);
xnor U46086 (N_46086,N_43169,N_44093);
and U46087 (N_46087,N_43111,N_43771);
and U46088 (N_46088,N_42619,N_43567);
and U46089 (N_46089,N_42863,N_42918);
or U46090 (N_46090,N_44144,N_43417);
and U46091 (N_46091,N_42766,N_43967);
nand U46092 (N_46092,N_44444,N_43652);
xor U46093 (N_46093,N_43494,N_44176);
and U46094 (N_46094,N_43014,N_42557);
nand U46095 (N_46095,N_43255,N_42697);
xor U46096 (N_46096,N_43173,N_44437);
nor U46097 (N_46097,N_43279,N_44149);
and U46098 (N_46098,N_43661,N_44269);
nor U46099 (N_46099,N_44216,N_43164);
and U46100 (N_46100,N_43877,N_43152);
xnor U46101 (N_46101,N_43135,N_43644);
nand U46102 (N_46102,N_42744,N_43056);
and U46103 (N_46103,N_44696,N_44910);
xnor U46104 (N_46104,N_42632,N_42812);
and U46105 (N_46105,N_44438,N_44984);
xor U46106 (N_46106,N_44979,N_44459);
and U46107 (N_46107,N_44812,N_44273);
nor U46108 (N_46108,N_42772,N_44325);
or U46109 (N_46109,N_44356,N_42925);
nand U46110 (N_46110,N_42999,N_44341);
nand U46111 (N_46111,N_44053,N_44876);
xor U46112 (N_46112,N_44716,N_44854);
nor U46113 (N_46113,N_44564,N_43759);
xor U46114 (N_46114,N_43423,N_42591);
nor U46115 (N_46115,N_43256,N_43431);
nand U46116 (N_46116,N_43006,N_44567);
xnor U46117 (N_46117,N_43709,N_44357);
nand U46118 (N_46118,N_44515,N_43289);
or U46119 (N_46119,N_43291,N_43140);
xnor U46120 (N_46120,N_44764,N_43025);
or U46121 (N_46121,N_43765,N_44756);
and U46122 (N_46122,N_42674,N_43754);
and U46123 (N_46123,N_42737,N_42712);
xor U46124 (N_46124,N_42946,N_42722);
nor U46125 (N_46125,N_44385,N_43105);
nand U46126 (N_46126,N_42823,N_42936);
and U46127 (N_46127,N_43717,N_43267);
nor U46128 (N_46128,N_43948,N_43112);
nand U46129 (N_46129,N_44639,N_43190);
nor U46130 (N_46130,N_44941,N_42958);
or U46131 (N_46131,N_44711,N_42742);
nor U46132 (N_46132,N_43021,N_43218);
or U46133 (N_46133,N_43748,N_44090);
nand U46134 (N_46134,N_42550,N_44361);
and U46135 (N_46135,N_43471,N_43129);
xor U46136 (N_46136,N_44685,N_42921);
nand U46137 (N_46137,N_43795,N_44652);
xnor U46138 (N_46138,N_43467,N_44294);
xor U46139 (N_46139,N_44120,N_44929);
nor U46140 (N_46140,N_42781,N_44322);
nand U46141 (N_46141,N_43434,N_42612);
nor U46142 (N_46142,N_44725,N_44513);
nor U46143 (N_46143,N_44426,N_44824);
or U46144 (N_46144,N_44420,N_43735);
or U46145 (N_46145,N_44009,N_44414);
and U46146 (N_46146,N_44657,N_43672);
nand U46147 (N_46147,N_44622,N_43395);
xor U46148 (N_46148,N_42873,N_43499);
and U46149 (N_46149,N_44488,N_42698);
xor U46150 (N_46150,N_43760,N_42660);
nand U46151 (N_46151,N_43110,N_42927);
xor U46152 (N_46152,N_43035,N_44534);
nand U46153 (N_46153,N_42733,N_43044);
xnor U46154 (N_46154,N_44607,N_44695);
nor U46155 (N_46155,N_44465,N_43290);
and U46156 (N_46156,N_43799,N_43568);
nand U46157 (N_46157,N_43185,N_43160);
and U46158 (N_46158,N_43864,N_43127);
xnor U46159 (N_46159,N_43899,N_44805);
xnor U46160 (N_46160,N_43130,N_43715);
and U46161 (N_46161,N_44281,N_44489);
or U46162 (N_46162,N_44440,N_43323);
nor U46163 (N_46163,N_44153,N_43581);
and U46164 (N_46164,N_44690,N_44134);
xnor U46165 (N_46165,N_43521,N_43633);
nand U46166 (N_46166,N_43720,N_44733);
nor U46167 (N_46167,N_44731,N_44022);
nand U46168 (N_46168,N_43310,N_43295);
or U46169 (N_46169,N_43923,N_43480);
or U46170 (N_46170,N_43664,N_43344);
xor U46171 (N_46171,N_44066,N_42972);
nor U46172 (N_46172,N_43812,N_44970);
and U46173 (N_46173,N_43733,N_43778);
nor U46174 (N_46174,N_44359,N_44064);
or U46175 (N_46175,N_44741,N_44760);
nor U46176 (N_46176,N_43908,N_44668);
nor U46177 (N_46177,N_44982,N_44264);
nor U46178 (N_46178,N_44056,N_44453);
and U46179 (N_46179,N_42943,N_44889);
or U46180 (N_46180,N_44233,N_43972);
and U46181 (N_46181,N_44506,N_42561);
xnor U46182 (N_46182,N_44985,N_44780);
nor U46183 (N_46183,N_42991,N_44071);
and U46184 (N_46184,N_42599,N_42539);
nand U46185 (N_46185,N_43374,N_42851);
or U46186 (N_46186,N_44588,N_44605);
nor U46187 (N_46187,N_43847,N_43084);
nand U46188 (N_46188,N_42657,N_42883);
and U46189 (N_46189,N_44025,N_42931);
nor U46190 (N_46190,N_44092,N_43675);
nand U46191 (N_46191,N_44659,N_44055);
or U46192 (N_46192,N_44247,N_43410);
nand U46193 (N_46193,N_42939,N_43792);
nor U46194 (N_46194,N_44462,N_43119);
or U46195 (N_46195,N_44317,N_43730);
xor U46196 (N_46196,N_44335,N_43663);
nand U46197 (N_46197,N_43690,N_43092);
or U46198 (N_46198,N_43623,N_44114);
and U46199 (N_46199,N_44914,N_43222);
nand U46200 (N_46200,N_43642,N_43744);
or U46201 (N_46201,N_43820,N_44215);
or U46202 (N_46202,N_44429,N_43547);
nand U46203 (N_46203,N_42717,N_42929);
or U46204 (N_46204,N_42897,N_43379);
nand U46205 (N_46205,N_44883,N_42750);
xor U46206 (N_46206,N_43920,N_42751);
and U46207 (N_46207,N_44082,N_43782);
or U46208 (N_46208,N_43296,N_42628);
nand U46209 (N_46209,N_43662,N_43076);
nand U46210 (N_46210,N_42970,N_43880);
or U46211 (N_46211,N_43685,N_43024);
or U46212 (N_46212,N_43115,N_44496);
nand U46213 (N_46213,N_42996,N_43558);
or U46214 (N_46214,N_44051,N_42794);
nand U46215 (N_46215,N_44518,N_43887);
and U46216 (N_46216,N_43951,N_43713);
xor U46217 (N_46217,N_44640,N_43873);
nand U46218 (N_46218,N_44481,N_43929);
xnor U46219 (N_46219,N_43620,N_42548);
nor U46220 (N_46220,N_43684,N_44378);
nand U46221 (N_46221,N_43725,N_43588);
nand U46222 (N_46222,N_42833,N_44099);
and U46223 (N_46223,N_43463,N_42870);
xor U46224 (N_46224,N_42889,N_44791);
or U46225 (N_46225,N_44299,N_44102);
nand U46226 (N_46226,N_43216,N_42759);
and U46227 (N_46227,N_44196,N_43691);
xnor U46228 (N_46228,N_43974,N_43174);
nor U46229 (N_46229,N_43512,N_43057);
and U46230 (N_46230,N_43364,N_43670);
nor U46231 (N_46231,N_43414,N_44523);
or U46232 (N_46232,N_43239,N_43259);
xor U46233 (N_46233,N_44858,N_43607);
nor U46234 (N_46234,N_44547,N_43193);
nor U46235 (N_46235,N_44316,N_44806);
nand U46236 (N_46236,N_44849,N_44241);
xnor U46237 (N_46237,N_43738,N_44037);
nand U46238 (N_46238,N_43538,N_44400);
nand U46239 (N_46239,N_42606,N_42824);
and U46240 (N_46240,N_44936,N_44922);
nor U46241 (N_46241,N_43250,N_44358);
and U46242 (N_46242,N_43589,N_42630);
nand U46243 (N_46243,N_43486,N_44947);
xnor U46244 (N_46244,N_44818,N_43879);
and U46245 (N_46245,N_43594,N_43775);
or U46246 (N_46246,N_44463,N_43273);
or U46247 (N_46247,N_44409,N_44155);
xnor U46248 (N_46248,N_44204,N_43781);
nor U46249 (N_46249,N_43221,N_42904);
or U46250 (N_46250,N_43445,N_43316);
xor U46251 (N_46251,N_43381,N_44045);
xor U46252 (N_46252,N_43584,N_44788);
or U46253 (N_46253,N_43485,N_43840);
or U46254 (N_46254,N_43168,N_44644);
nor U46255 (N_46255,N_42940,N_42595);
nand U46256 (N_46256,N_43484,N_44466);
and U46257 (N_46257,N_44414,N_43619);
nor U46258 (N_46258,N_44475,N_44242);
nand U46259 (N_46259,N_44747,N_43599);
nand U46260 (N_46260,N_43861,N_44715);
or U46261 (N_46261,N_42923,N_44468);
xor U46262 (N_46262,N_44148,N_43391);
and U46263 (N_46263,N_43372,N_42685);
and U46264 (N_46264,N_44224,N_43005);
nand U46265 (N_46265,N_44032,N_43443);
xnor U46266 (N_46266,N_43886,N_44230);
or U46267 (N_46267,N_44048,N_44257);
xnor U46268 (N_46268,N_42555,N_43437);
nand U46269 (N_46269,N_43542,N_44740);
nor U46270 (N_46270,N_44145,N_44889);
xnor U46271 (N_46271,N_44964,N_42531);
xor U46272 (N_46272,N_44392,N_43865);
nand U46273 (N_46273,N_42966,N_44028);
nor U46274 (N_46274,N_43610,N_44396);
xor U46275 (N_46275,N_44923,N_43853);
and U46276 (N_46276,N_42945,N_42891);
or U46277 (N_46277,N_43953,N_44403);
and U46278 (N_46278,N_43816,N_43305);
or U46279 (N_46279,N_43440,N_42899);
nor U46280 (N_46280,N_44745,N_43461);
or U46281 (N_46281,N_43195,N_42907);
nand U46282 (N_46282,N_42715,N_43520);
and U46283 (N_46283,N_44276,N_44252);
xnor U46284 (N_46284,N_42713,N_43171);
nand U46285 (N_46285,N_43625,N_44205);
nor U46286 (N_46286,N_42920,N_44467);
xor U46287 (N_46287,N_43127,N_43046);
nand U46288 (N_46288,N_42934,N_42909);
xor U46289 (N_46289,N_44905,N_43937);
xor U46290 (N_46290,N_44652,N_44859);
xnor U46291 (N_46291,N_42554,N_42689);
or U46292 (N_46292,N_43154,N_44170);
or U46293 (N_46293,N_44274,N_43029);
or U46294 (N_46294,N_43579,N_43479);
nand U46295 (N_46295,N_43911,N_43045);
xnor U46296 (N_46296,N_42845,N_44264);
or U46297 (N_46297,N_42635,N_43668);
or U46298 (N_46298,N_43809,N_44232);
and U46299 (N_46299,N_44256,N_44813);
and U46300 (N_46300,N_44488,N_43185);
nand U46301 (N_46301,N_43940,N_44246);
nor U46302 (N_46302,N_42826,N_44093);
and U46303 (N_46303,N_44731,N_43951);
nand U46304 (N_46304,N_44781,N_42846);
and U46305 (N_46305,N_42776,N_44612);
xnor U46306 (N_46306,N_42602,N_44872);
or U46307 (N_46307,N_44742,N_44046);
and U46308 (N_46308,N_43499,N_42841);
xnor U46309 (N_46309,N_43205,N_43584);
nor U46310 (N_46310,N_43103,N_42584);
and U46311 (N_46311,N_44798,N_43380);
nand U46312 (N_46312,N_44096,N_42778);
nand U46313 (N_46313,N_43461,N_43446);
nand U46314 (N_46314,N_42674,N_43284);
xnor U46315 (N_46315,N_42738,N_44500);
xnor U46316 (N_46316,N_44466,N_42544);
nand U46317 (N_46317,N_43681,N_43903);
nand U46318 (N_46318,N_44189,N_43809);
and U46319 (N_46319,N_43140,N_44544);
nor U46320 (N_46320,N_43944,N_44227);
or U46321 (N_46321,N_43307,N_44107);
nor U46322 (N_46322,N_43867,N_42802);
nand U46323 (N_46323,N_44449,N_43691);
or U46324 (N_46324,N_44954,N_43731);
nor U46325 (N_46325,N_44618,N_44980);
or U46326 (N_46326,N_44632,N_43988);
and U46327 (N_46327,N_44771,N_43252);
xor U46328 (N_46328,N_43566,N_43476);
nor U46329 (N_46329,N_42789,N_44185);
and U46330 (N_46330,N_44736,N_44360);
nand U46331 (N_46331,N_44481,N_43768);
nor U46332 (N_46332,N_44833,N_43272);
nand U46333 (N_46333,N_44959,N_42614);
or U46334 (N_46334,N_43376,N_43588);
xor U46335 (N_46335,N_44146,N_44284);
xnor U46336 (N_46336,N_44296,N_44565);
xor U46337 (N_46337,N_44735,N_44370);
xnor U46338 (N_46338,N_44962,N_44150);
xnor U46339 (N_46339,N_43939,N_43842);
nand U46340 (N_46340,N_43547,N_43601);
nand U46341 (N_46341,N_43595,N_44772);
nand U46342 (N_46342,N_44728,N_44307);
nor U46343 (N_46343,N_44620,N_44404);
xnor U46344 (N_46344,N_42577,N_42670);
or U46345 (N_46345,N_43644,N_44489);
xor U46346 (N_46346,N_43312,N_44867);
nand U46347 (N_46347,N_44126,N_44087);
nor U46348 (N_46348,N_42644,N_44199);
xnor U46349 (N_46349,N_44469,N_43371);
or U46350 (N_46350,N_44537,N_44324);
xnor U46351 (N_46351,N_43940,N_44538);
nand U46352 (N_46352,N_42909,N_44157);
and U46353 (N_46353,N_43792,N_44556);
and U46354 (N_46354,N_44029,N_43830);
nand U46355 (N_46355,N_43014,N_44396);
and U46356 (N_46356,N_44946,N_42828);
and U46357 (N_46357,N_44360,N_43546);
nand U46358 (N_46358,N_44419,N_43331);
xor U46359 (N_46359,N_42594,N_43070);
or U46360 (N_46360,N_43966,N_43633);
xnor U46361 (N_46361,N_42701,N_43666);
nor U46362 (N_46362,N_44211,N_44503);
nor U46363 (N_46363,N_42551,N_43205);
nand U46364 (N_46364,N_42766,N_43740);
and U46365 (N_46365,N_44775,N_42559);
nor U46366 (N_46366,N_42756,N_42513);
nor U46367 (N_46367,N_44039,N_44563);
and U46368 (N_46368,N_43257,N_43239);
nand U46369 (N_46369,N_44988,N_43444);
and U46370 (N_46370,N_44155,N_44494);
nor U46371 (N_46371,N_43197,N_44938);
nand U46372 (N_46372,N_43614,N_44709);
or U46373 (N_46373,N_43425,N_43075);
xor U46374 (N_46374,N_43400,N_44711);
or U46375 (N_46375,N_44877,N_44117);
and U46376 (N_46376,N_44399,N_43037);
nor U46377 (N_46377,N_43608,N_43253);
xor U46378 (N_46378,N_44805,N_43482);
nand U46379 (N_46379,N_44163,N_44818);
or U46380 (N_46380,N_44925,N_43612);
or U46381 (N_46381,N_42960,N_43403);
nor U46382 (N_46382,N_43560,N_43710);
or U46383 (N_46383,N_44722,N_44212);
nand U46384 (N_46384,N_43319,N_44030);
and U46385 (N_46385,N_44873,N_44741);
and U46386 (N_46386,N_44893,N_43181);
xor U46387 (N_46387,N_44614,N_43328);
or U46388 (N_46388,N_44902,N_43392);
nor U46389 (N_46389,N_43781,N_44811);
or U46390 (N_46390,N_43330,N_44409);
xor U46391 (N_46391,N_42778,N_43645);
nand U46392 (N_46392,N_43636,N_43285);
and U46393 (N_46393,N_42562,N_43569);
or U46394 (N_46394,N_43678,N_43550);
xor U46395 (N_46395,N_44404,N_43295);
nand U46396 (N_46396,N_44137,N_44288);
or U46397 (N_46397,N_43173,N_43089);
xor U46398 (N_46398,N_42912,N_43415);
or U46399 (N_46399,N_43633,N_44038);
xor U46400 (N_46400,N_44719,N_43151);
and U46401 (N_46401,N_42633,N_43495);
and U46402 (N_46402,N_42897,N_44674);
nand U46403 (N_46403,N_42648,N_44318);
nand U46404 (N_46404,N_44655,N_44904);
nand U46405 (N_46405,N_44946,N_44262);
xnor U46406 (N_46406,N_43920,N_43432);
xor U46407 (N_46407,N_43867,N_42659);
xor U46408 (N_46408,N_43909,N_44356);
or U46409 (N_46409,N_43886,N_42658);
xnor U46410 (N_46410,N_42975,N_44865);
nor U46411 (N_46411,N_42650,N_44708);
nand U46412 (N_46412,N_43465,N_42894);
nor U46413 (N_46413,N_44676,N_43098);
xnor U46414 (N_46414,N_44608,N_44640);
nor U46415 (N_46415,N_43735,N_42660);
or U46416 (N_46416,N_43358,N_43010);
and U46417 (N_46417,N_44422,N_43849);
or U46418 (N_46418,N_43270,N_44830);
xor U46419 (N_46419,N_44780,N_43517);
or U46420 (N_46420,N_42562,N_44383);
nor U46421 (N_46421,N_43041,N_43365);
or U46422 (N_46422,N_43240,N_42783);
xnor U46423 (N_46423,N_42784,N_44786);
or U46424 (N_46424,N_44312,N_44170);
nor U46425 (N_46425,N_43772,N_43396);
and U46426 (N_46426,N_42981,N_44779);
nor U46427 (N_46427,N_44020,N_44659);
nor U46428 (N_46428,N_43340,N_44055);
xor U46429 (N_46429,N_44823,N_44560);
and U46430 (N_46430,N_42960,N_43292);
nor U46431 (N_46431,N_43641,N_44257);
nor U46432 (N_46432,N_43479,N_43539);
nand U46433 (N_46433,N_42840,N_43417);
nand U46434 (N_46434,N_43467,N_42969);
nor U46435 (N_46435,N_43837,N_43232);
nand U46436 (N_46436,N_44208,N_43743);
or U46437 (N_46437,N_42702,N_44293);
and U46438 (N_46438,N_43875,N_44987);
and U46439 (N_46439,N_43498,N_43205);
xnor U46440 (N_46440,N_44524,N_44104);
xor U46441 (N_46441,N_42938,N_43100);
nand U46442 (N_46442,N_43975,N_43885);
nand U46443 (N_46443,N_43877,N_44147);
nor U46444 (N_46444,N_44677,N_43753);
or U46445 (N_46445,N_44595,N_44642);
and U46446 (N_46446,N_44655,N_43602);
nand U46447 (N_46447,N_43988,N_42924);
xnor U46448 (N_46448,N_44141,N_44168);
nor U46449 (N_46449,N_43359,N_43130);
or U46450 (N_46450,N_42699,N_43150);
xnor U46451 (N_46451,N_44798,N_44298);
nand U46452 (N_46452,N_43452,N_43845);
xnor U46453 (N_46453,N_43451,N_42992);
or U46454 (N_46454,N_42676,N_44739);
nor U46455 (N_46455,N_43130,N_43429);
nor U46456 (N_46456,N_43493,N_44871);
nor U46457 (N_46457,N_43381,N_43890);
or U46458 (N_46458,N_44223,N_43628);
xor U46459 (N_46459,N_42714,N_42658);
nand U46460 (N_46460,N_42915,N_44863);
nor U46461 (N_46461,N_43527,N_43672);
nand U46462 (N_46462,N_44852,N_43723);
or U46463 (N_46463,N_43346,N_44748);
nand U46464 (N_46464,N_43775,N_43810);
nand U46465 (N_46465,N_44725,N_43350);
nor U46466 (N_46466,N_43446,N_44592);
nand U46467 (N_46467,N_44113,N_44234);
nor U46468 (N_46468,N_44392,N_44897);
nand U46469 (N_46469,N_42973,N_43043);
nand U46470 (N_46470,N_42778,N_44434);
or U46471 (N_46471,N_42724,N_43670);
nand U46472 (N_46472,N_43348,N_43010);
or U46473 (N_46473,N_44158,N_44750);
or U46474 (N_46474,N_44574,N_43024);
nor U46475 (N_46475,N_43991,N_43093);
and U46476 (N_46476,N_43387,N_43572);
xnor U46477 (N_46477,N_43697,N_43176);
and U46478 (N_46478,N_42825,N_42658);
xnor U46479 (N_46479,N_42825,N_42960);
nand U46480 (N_46480,N_44324,N_44242);
or U46481 (N_46481,N_44551,N_44233);
nor U46482 (N_46482,N_44317,N_43657);
xnor U46483 (N_46483,N_42679,N_44237);
nand U46484 (N_46484,N_43395,N_44347);
nor U46485 (N_46485,N_44656,N_44993);
nor U46486 (N_46486,N_42717,N_43329);
xor U46487 (N_46487,N_43685,N_42745);
xor U46488 (N_46488,N_42619,N_43476);
nand U46489 (N_46489,N_44536,N_44775);
nand U46490 (N_46490,N_43510,N_43558);
nand U46491 (N_46491,N_44689,N_44790);
nand U46492 (N_46492,N_44730,N_44807);
nand U46493 (N_46493,N_44666,N_44114);
and U46494 (N_46494,N_43016,N_42559);
xor U46495 (N_46495,N_44050,N_43792);
xnor U46496 (N_46496,N_42893,N_44881);
nor U46497 (N_46497,N_42526,N_44151);
and U46498 (N_46498,N_43306,N_44181);
nor U46499 (N_46499,N_44765,N_44292);
nand U46500 (N_46500,N_44806,N_43380);
or U46501 (N_46501,N_44428,N_43666);
nor U46502 (N_46502,N_43221,N_42924);
and U46503 (N_46503,N_43844,N_44650);
nor U46504 (N_46504,N_43592,N_43185);
nor U46505 (N_46505,N_44834,N_44431);
nand U46506 (N_46506,N_43136,N_43356);
nor U46507 (N_46507,N_44170,N_43636);
and U46508 (N_46508,N_44030,N_44867);
or U46509 (N_46509,N_42732,N_43306);
or U46510 (N_46510,N_42652,N_43388);
or U46511 (N_46511,N_44915,N_44242);
xnor U46512 (N_46512,N_44869,N_43867);
xor U46513 (N_46513,N_44656,N_43293);
xor U46514 (N_46514,N_43089,N_44266);
and U46515 (N_46515,N_44771,N_44036);
or U46516 (N_46516,N_43215,N_43056);
nand U46517 (N_46517,N_42522,N_44501);
nand U46518 (N_46518,N_43951,N_43240);
nand U46519 (N_46519,N_43128,N_43157);
or U46520 (N_46520,N_43654,N_43595);
and U46521 (N_46521,N_44033,N_44229);
xor U46522 (N_46522,N_44943,N_43699);
and U46523 (N_46523,N_44432,N_43798);
xnor U46524 (N_46524,N_42942,N_43277);
or U46525 (N_46525,N_43736,N_43731);
and U46526 (N_46526,N_43516,N_42983);
xor U46527 (N_46527,N_42521,N_44075);
nor U46528 (N_46528,N_42995,N_43715);
nor U46529 (N_46529,N_44013,N_43788);
or U46530 (N_46530,N_44708,N_44589);
nor U46531 (N_46531,N_43010,N_42790);
nor U46532 (N_46532,N_44255,N_43627);
and U46533 (N_46533,N_43118,N_43758);
and U46534 (N_46534,N_43561,N_43235);
or U46535 (N_46535,N_43036,N_44988);
or U46536 (N_46536,N_43873,N_43206);
or U46537 (N_46537,N_42877,N_43458);
or U46538 (N_46538,N_44952,N_44903);
xnor U46539 (N_46539,N_44708,N_42747);
or U46540 (N_46540,N_44718,N_43105);
and U46541 (N_46541,N_43606,N_44359);
xor U46542 (N_46542,N_44566,N_44276);
nand U46543 (N_46543,N_43853,N_43212);
xnor U46544 (N_46544,N_43516,N_44292);
nor U46545 (N_46545,N_43496,N_42998);
xor U46546 (N_46546,N_44298,N_43527);
nand U46547 (N_46547,N_43374,N_43662);
and U46548 (N_46548,N_44006,N_44018);
and U46549 (N_46549,N_44720,N_43345);
xnor U46550 (N_46550,N_43945,N_44492);
and U46551 (N_46551,N_44739,N_42749);
and U46552 (N_46552,N_42870,N_42628);
nand U46553 (N_46553,N_42845,N_44637);
and U46554 (N_46554,N_42743,N_43196);
nor U46555 (N_46555,N_42513,N_43957);
nor U46556 (N_46556,N_44166,N_44372);
or U46557 (N_46557,N_43431,N_43619);
and U46558 (N_46558,N_43010,N_43785);
or U46559 (N_46559,N_43500,N_43725);
xnor U46560 (N_46560,N_42707,N_44688);
xnor U46561 (N_46561,N_44021,N_42591);
xor U46562 (N_46562,N_44197,N_44579);
or U46563 (N_46563,N_42975,N_42822);
nand U46564 (N_46564,N_44244,N_42725);
nor U46565 (N_46565,N_44333,N_43520);
and U46566 (N_46566,N_44483,N_43713);
nor U46567 (N_46567,N_44823,N_44736);
xnor U46568 (N_46568,N_43746,N_44708);
nor U46569 (N_46569,N_42772,N_44615);
or U46570 (N_46570,N_44988,N_44991);
or U46571 (N_46571,N_44376,N_44017);
nand U46572 (N_46572,N_43744,N_44727);
xor U46573 (N_46573,N_44701,N_42865);
nor U46574 (N_46574,N_44088,N_44275);
xnor U46575 (N_46575,N_43245,N_42997);
or U46576 (N_46576,N_44364,N_43459);
nor U46577 (N_46577,N_42946,N_43585);
nor U46578 (N_46578,N_42527,N_43652);
xnor U46579 (N_46579,N_43827,N_43647);
nand U46580 (N_46580,N_44725,N_44556);
nand U46581 (N_46581,N_44894,N_42523);
nor U46582 (N_46582,N_44517,N_43150);
nor U46583 (N_46583,N_42816,N_44707);
xor U46584 (N_46584,N_42825,N_43165);
or U46585 (N_46585,N_44058,N_43897);
nand U46586 (N_46586,N_44481,N_43960);
xor U46587 (N_46587,N_43975,N_44740);
nor U46588 (N_46588,N_42660,N_42752);
or U46589 (N_46589,N_44302,N_44573);
nor U46590 (N_46590,N_44061,N_43332);
or U46591 (N_46591,N_43507,N_43761);
and U46592 (N_46592,N_44008,N_43641);
or U46593 (N_46593,N_44374,N_44861);
nor U46594 (N_46594,N_44361,N_43313);
and U46595 (N_46595,N_43395,N_43352);
or U46596 (N_46596,N_44168,N_43149);
nand U46597 (N_46597,N_44920,N_43671);
nand U46598 (N_46598,N_44580,N_44969);
and U46599 (N_46599,N_43186,N_44144);
nand U46600 (N_46600,N_43692,N_43799);
nor U46601 (N_46601,N_42863,N_44655);
and U46602 (N_46602,N_42536,N_42685);
nand U46603 (N_46603,N_44375,N_43061);
or U46604 (N_46604,N_43378,N_43613);
nor U46605 (N_46605,N_42901,N_43184);
xnor U46606 (N_46606,N_42746,N_44731);
xnor U46607 (N_46607,N_43804,N_43587);
or U46608 (N_46608,N_44082,N_43046);
and U46609 (N_46609,N_43893,N_44203);
nor U46610 (N_46610,N_43572,N_43449);
nand U46611 (N_46611,N_44734,N_43616);
or U46612 (N_46612,N_44212,N_43935);
nor U46613 (N_46613,N_44334,N_44760);
nor U46614 (N_46614,N_42522,N_44396);
xnor U46615 (N_46615,N_43862,N_44924);
xor U46616 (N_46616,N_43020,N_44847);
or U46617 (N_46617,N_42708,N_42636);
or U46618 (N_46618,N_42701,N_43453);
and U46619 (N_46619,N_44822,N_43306);
or U46620 (N_46620,N_44868,N_43504);
xnor U46621 (N_46621,N_44396,N_43325);
nand U46622 (N_46622,N_44715,N_44497);
and U46623 (N_46623,N_43386,N_43272);
nand U46624 (N_46624,N_43152,N_44004);
nor U46625 (N_46625,N_43273,N_43525);
and U46626 (N_46626,N_44677,N_42777);
xor U46627 (N_46627,N_43589,N_42526);
xor U46628 (N_46628,N_43640,N_44952);
and U46629 (N_46629,N_43126,N_44826);
and U46630 (N_46630,N_44026,N_43415);
nand U46631 (N_46631,N_43707,N_44161);
or U46632 (N_46632,N_42513,N_44497);
and U46633 (N_46633,N_42852,N_42811);
nor U46634 (N_46634,N_44248,N_44479);
nand U46635 (N_46635,N_42914,N_42994);
xor U46636 (N_46636,N_43046,N_44327);
xnor U46637 (N_46637,N_43258,N_43544);
nand U46638 (N_46638,N_43284,N_44426);
nor U46639 (N_46639,N_44530,N_44750);
nor U46640 (N_46640,N_42995,N_42716);
nor U46641 (N_46641,N_44252,N_42789);
nor U46642 (N_46642,N_44414,N_44107);
xnor U46643 (N_46643,N_44493,N_44575);
nor U46644 (N_46644,N_43967,N_44348);
or U46645 (N_46645,N_43042,N_44553);
xor U46646 (N_46646,N_43974,N_43595);
nor U46647 (N_46647,N_43023,N_44515);
and U46648 (N_46648,N_44403,N_44124);
nor U46649 (N_46649,N_43342,N_43475);
xor U46650 (N_46650,N_42528,N_43922);
nand U46651 (N_46651,N_44459,N_44801);
xor U46652 (N_46652,N_42578,N_42715);
nor U46653 (N_46653,N_43367,N_42562);
nor U46654 (N_46654,N_43565,N_43838);
and U46655 (N_46655,N_44636,N_44822);
xnor U46656 (N_46656,N_43319,N_44220);
or U46657 (N_46657,N_42687,N_42925);
nand U46658 (N_46658,N_43834,N_44681);
xnor U46659 (N_46659,N_42731,N_44853);
or U46660 (N_46660,N_44662,N_43922);
xnor U46661 (N_46661,N_43531,N_44469);
xor U46662 (N_46662,N_43580,N_43529);
nand U46663 (N_46663,N_44262,N_43569);
and U46664 (N_46664,N_43408,N_42568);
or U46665 (N_46665,N_43287,N_42528);
nor U46666 (N_46666,N_44125,N_44817);
or U46667 (N_46667,N_43778,N_42550);
and U46668 (N_46668,N_44863,N_44991);
nand U46669 (N_46669,N_43133,N_44355);
nand U46670 (N_46670,N_43117,N_44306);
and U46671 (N_46671,N_44679,N_44436);
xnor U46672 (N_46672,N_44891,N_43311);
and U46673 (N_46673,N_44717,N_44937);
and U46674 (N_46674,N_44990,N_42585);
nand U46675 (N_46675,N_43077,N_44249);
and U46676 (N_46676,N_43114,N_43908);
and U46677 (N_46677,N_43631,N_43627);
and U46678 (N_46678,N_42656,N_43275);
nor U46679 (N_46679,N_43715,N_43657);
and U46680 (N_46680,N_44144,N_44280);
and U46681 (N_46681,N_44545,N_44387);
and U46682 (N_46682,N_42758,N_43730);
nor U46683 (N_46683,N_43097,N_43337);
nand U46684 (N_46684,N_44489,N_43319);
or U46685 (N_46685,N_44575,N_43581);
xnor U46686 (N_46686,N_43222,N_42694);
or U46687 (N_46687,N_43889,N_44328);
nor U46688 (N_46688,N_43598,N_43591);
and U46689 (N_46689,N_44206,N_43161);
nor U46690 (N_46690,N_44375,N_43759);
or U46691 (N_46691,N_44759,N_44916);
nor U46692 (N_46692,N_42769,N_44611);
or U46693 (N_46693,N_43046,N_43776);
nand U46694 (N_46694,N_44255,N_44021);
and U46695 (N_46695,N_44560,N_42562);
nor U46696 (N_46696,N_43537,N_43771);
nor U46697 (N_46697,N_43027,N_44412);
or U46698 (N_46698,N_43283,N_43906);
nand U46699 (N_46699,N_44217,N_44069);
xor U46700 (N_46700,N_43271,N_43623);
nor U46701 (N_46701,N_44335,N_44029);
or U46702 (N_46702,N_42600,N_43149);
and U46703 (N_46703,N_42836,N_44025);
or U46704 (N_46704,N_43144,N_42792);
xnor U46705 (N_46705,N_43666,N_44893);
nor U46706 (N_46706,N_44251,N_43997);
or U46707 (N_46707,N_44926,N_44687);
or U46708 (N_46708,N_44716,N_43089);
xnor U46709 (N_46709,N_44881,N_44202);
nor U46710 (N_46710,N_42836,N_44679);
and U46711 (N_46711,N_43559,N_44787);
or U46712 (N_46712,N_42970,N_43573);
and U46713 (N_46713,N_44386,N_42869);
and U46714 (N_46714,N_42582,N_43456);
nor U46715 (N_46715,N_42754,N_44197);
xor U46716 (N_46716,N_44692,N_42662);
and U46717 (N_46717,N_43732,N_44671);
nor U46718 (N_46718,N_43858,N_43196);
nand U46719 (N_46719,N_44268,N_44088);
xor U46720 (N_46720,N_44115,N_43567);
nor U46721 (N_46721,N_43991,N_43501);
nand U46722 (N_46722,N_44189,N_43155);
nand U46723 (N_46723,N_43458,N_42670);
and U46724 (N_46724,N_44989,N_43131);
nand U46725 (N_46725,N_43083,N_43492);
nand U46726 (N_46726,N_43414,N_42514);
xor U46727 (N_46727,N_44571,N_44841);
or U46728 (N_46728,N_43483,N_42853);
or U46729 (N_46729,N_43665,N_43174);
and U46730 (N_46730,N_44388,N_43560);
or U46731 (N_46731,N_44006,N_43701);
and U46732 (N_46732,N_44093,N_44182);
or U46733 (N_46733,N_42644,N_43405);
or U46734 (N_46734,N_44056,N_43557);
and U46735 (N_46735,N_43399,N_44845);
xor U46736 (N_46736,N_43238,N_42583);
and U46737 (N_46737,N_42771,N_42787);
nand U46738 (N_46738,N_42745,N_43460);
nand U46739 (N_46739,N_42907,N_42889);
nor U46740 (N_46740,N_44422,N_44000);
xnor U46741 (N_46741,N_43939,N_44790);
xor U46742 (N_46742,N_43014,N_43487);
and U46743 (N_46743,N_43625,N_44818);
or U46744 (N_46744,N_42648,N_43314);
xor U46745 (N_46745,N_44766,N_44261);
nor U46746 (N_46746,N_44194,N_42907);
xor U46747 (N_46747,N_44089,N_43695);
nand U46748 (N_46748,N_43268,N_43906);
nand U46749 (N_46749,N_44121,N_42517);
nand U46750 (N_46750,N_43813,N_43717);
and U46751 (N_46751,N_43474,N_44288);
and U46752 (N_46752,N_43152,N_42836);
or U46753 (N_46753,N_44751,N_44834);
or U46754 (N_46754,N_42891,N_42879);
or U46755 (N_46755,N_44750,N_43718);
xnor U46756 (N_46756,N_43345,N_44829);
xnor U46757 (N_46757,N_43422,N_43366);
nor U46758 (N_46758,N_43198,N_44341);
or U46759 (N_46759,N_42520,N_42562);
or U46760 (N_46760,N_43519,N_42933);
nor U46761 (N_46761,N_43352,N_44940);
xnor U46762 (N_46762,N_42998,N_43083);
and U46763 (N_46763,N_42790,N_44238);
xnor U46764 (N_46764,N_44181,N_44047);
xnor U46765 (N_46765,N_43702,N_44621);
or U46766 (N_46766,N_43711,N_42837);
nor U46767 (N_46767,N_43009,N_43036);
xor U46768 (N_46768,N_44838,N_43928);
nor U46769 (N_46769,N_44559,N_42697);
nor U46770 (N_46770,N_43606,N_44910);
nand U46771 (N_46771,N_43867,N_44100);
and U46772 (N_46772,N_44861,N_42737);
nand U46773 (N_46773,N_43215,N_44101);
nor U46774 (N_46774,N_44530,N_44797);
and U46775 (N_46775,N_43941,N_43520);
and U46776 (N_46776,N_44221,N_43854);
and U46777 (N_46777,N_42858,N_44316);
nand U46778 (N_46778,N_43871,N_43079);
nor U46779 (N_46779,N_43899,N_43729);
or U46780 (N_46780,N_44971,N_44778);
nor U46781 (N_46781,N_43994,N_42865);
xor U46782 (N_46782,N_42791,N_42994);
xnor U46783 (N_46783,N_44307,N_42641);
nor U46784 (N_46784,N_43129,N_43939);
and U46785 (N_46785,N_42611,N_43009);
and U46786 (N_46786,N_42950,N_44701);
nand U46787 (N_46787,N_42702,N_44059);
and U46788 (N_46788,N_43057,N_43252);
or U46789 (N_46789,N_44860,N_43130);
nor U46790 (N_46790,N_44928,N_42754);
xor U46791 (N_46791,N_44923,N_43869);
and U46792 (N_46792,N_43074,N_44948);
nand U46793 (N_46793,N_44409,N_43436);
nand U46794 (N_46794,N_44862,N_44089);
xnor U46795 (N_46795,N_42672,N_43936);
xor U46796 (N_46796,N_44165,N_42847);
and U46797 (N_46797,N_44739,N_42976);
and U46798 (N_46798,N_42560,N_44011);
xor U46799 (N_46799,N_43150,N_44386);
nand U46800 (N_46800,N_44043,N_42543);
nor U46801 (N_46801,N_44808,N_44110);
xor U46802 (N_46802,N_44306,N_42960);
xor U46803 (N_46803,N_44098,N_43144);
nor U46804 (N_46804,N_44142,N_43485);
or U46805 (N_46805,N_43181,N_44999);
xnor U46806 (N_46806,N_43545,N_42639);
xor U46807 (N_46807,N_44620,N_43002);
xor U46808 (N_46808,N_44436,N_43940);
nor U46809 (N_46809,N_43755,N_43498);
xnor U46810 (N_46810,N_44724,N_44279);
and U46811 (N_46811,N_44183,N_43177);
nand U46812 (N_46812,N_44138,N_44140);
or U46813 (N_46813,N_43698,N_44060);
or U46814 (N_46814,N_44937,N_43307);
nor U46815 (N_46815,N_44010,N_44304);
nor U46816 (N_46816,N_44045,N_43050);
or U46817 (N_46817,N_44621,N_43246);
and U46818 (N_46818,N_44201,N_43774);
or U46819 (N_46819,N_43315,N_43999);
xor U46820 (N_46820,N_44043,N_43371);
xor U46821 (N_46821,N_43229,N_42534);
nor U46822 (N_46822,N_44048,N_44236);
nand U46823 (N_46823,N_44440,N_43309);
or U46824 (N_46824,N_44373,N_42764);
xor U46825 (N_46825,N_43994,N_42672);
nor U46826 (N_46826,N_43521,N_42784);
xor U46827 (N_46827,N_43203,N_44696);
and U46828 (N_46828,N_44675,N_44538);
xnor U46829 (N_46829,N_43666,N_44534);
xnor U46830 (N_46830,N_44912,N_42796);
and U46831 (N_46831,N_42972,N_44368);
and U46832 (N_46832,N_43602,N_44171);
or U46833 (N_46833,N_44791,N_43289);
xnor U46834 (N_46834,N_43880,N_42621);
and U46835 (N_46835,N_42889,N_43752);
xnor U46836 (N_46836,N_44620,N_44821);
nor U46837 (N_46837,N_43590,N_43698);
nor U46838 (N_46838,N_44501,N_44296);
nor U46839 (N_46839,N_44413,N_43657);
nand U46840 (N_46840,N_43188,N_43510);
nand U46841 (N_46841,N_43152,N_44789);
and U46842 (N_46842,N_43841,N_42593);
nand U46843 (N_46843,N_43978,N_44459);
or U46844 (N_46844,N_43387,N_43009);
nand U46845 (N_46845,N_44724,N_44874);
nor U46846 (N_46846,N_43797,N_42839);
and U46847 (N_46847,N_43702,N_44979);
and U46848 (N_46848,N_43389,N_43543);
nand U46849 (N_46849,N_43554,N_44773);
or U46850 (N_46850,N_44475,N_44208);
xnor U46851 (N_46851,N_44109,N_42696);
xor U46852 (N_46852,N_44148,N_42784);
or U46853 (N_46853,N_42583,N_44946);
nand U46854 (N_46854,N_42742,N_42933);
nor U46855 (N_46855,N_43739,N_43661);
nor U46856 (N_46856,N_43304,N_43189);
or U46857 (N_46857,N_44836,N_44203);
and U46858 (N_46858,N_43713,N_44476);
nand U46859 (N_46859,N_43505,N_42646);
nor U46860 (N_46860,N_43523,N_42841);
nand U46861 (N_46861,N_43623,N_44071);
nand U46862 (N_46862,N_44110,N_43137);
nor U46863 (N_46863,N_44140,N_43945);
and U46864 (N_46864,N_44122,N_43792);
nor U46865 (N_46865,N_44007,N_42602);
and U46866 (N_46866,N_43232,N_43595);
xor U46867 (N_46867,N_44212,N_43639);
and U46868 (N_46868,N_44828,N_42709);
or U46869 (N_46869,N_43043,N_44299);
or U46870 (N_46870,N_44631,N_43290);
or U46871 (N_46871,N_44034,N_43605);
and U46872 (N_46872,N_43813,N_44941);
nand U46873 (N_46873,N_42992,N_44053);
nor U46874 (N_46874,N_43770,N_42672);
nand U46875 (N_46875,N_43845,N_44836);
nor U46876 (N_46876,N_42741,N_44256);
xnor U46877 (N_46877,N_42816,N_42919);
xor U46878 (N_46878,N_42820,N_42982);
nand U46879 (N_46879,N_42788,N_43060);
nand U46880 (N_46880,N_43605,N_42777);
nand U46881 (N_46881,N_43932,N_44298);
nor U46882 (N_46882,N_44661,N_42588);
xnor U46883 (N_46883,N_43708,N_44617);
nand U46884 (N_46884,N_43027,N_44808);
and U46885 (N_46885,N_44611,N_42808);
and U46886 (N_46886,N_42988,N_44266);
nor U46887 (N_46887,N_43271,N_42990);
nor U46888 (N_46888,N_43987,N_44999);
and U46889 (N_46889,N_43975,N_44581);
and U46890 (N_46890,N_42697,N_43476);
nand U46891 (N_46891,N_43149,N_43335);
xor U46892 (N_46892,N_43337,N_43549);
or U46893 (N_46893,N_44085,N_43218);
nand U46894 (N_46894,N_43544,N_44522);
and U46895 (N_46895,N_44784,N_42516);
and U46896 (N_46896,N_43256,N_44978);
nor U46897 (N_46897,N_43251,N_43116);
nand U46898 (N_46898,N_44937,N_43957);
xor U46899 (N_46899,N_42512,N_43849);
nor U46900 (N_46900,N_43665,N_44198);
and U46901 (N_46901,N_43322,N_42774);
nor U46902 (N_46902,N_44984,N_44087);
and U46903 (N_46903,N_43032,N_44670);
nor U46904 (N_46904,N_44227,N_44302);
or U46905 (N_46905,N_44787,N_44611);
xnor U46906 (N_46906,N_43509,N_43329);
nor U46907 (N_46907,N_44972,N_44835);
nor U46908 (N_46908,N_42996,N_43814);
xnor U46909 (N_46909,N_42875,N_44563);
or U46910 (N_46910,N_44538,N_44705);
xor U46911 (N_46911,N_44474,N_42599);
and U46912 (N_46912,N_43460,N_44813);
and U46913 (N_46913,N_44255,N_43822);
xnor U46914 (N_46914,N_43022,N_43867);
xor U46915 (N_46915,N_43633,N_44479);
nor U46916 (N_46916,N_44698,N_43833);
xnor U46917 (N_46917,N_44606,N_43336);
and U46918 (N_46918,N_44005,N_44858);
or U46919 (N_46919,N_43998,N_44227);
xnor U46920 (N_46920,N_44378,N_42670);
or U46921 (N_46921,N_43645,N_43469);
nand U46922 (N_46922,N_43453,N_42888);
nand U46923 (N_46923,N_42633,N_42928);
nand U46924 (N_46924,N_44901,N_42524);
xor U46925 (N_46925,N_44867,N_43383);
nor U46926 (N_46926,N_43810,N_43426);
xor U46927 (N_46927,N_43839,N_42756);
xor U46928 (N_46928,N_43797,N_44606);
xor U46929 (N_46929,N_44348,N_44244);
nor U46930 (N_46930,N_43997,N_42588);
xnor U46931 (N_46931,N_43904,N_44525);
or U46932 (N_46932,N_44933,N_44331);
xor U46933 (N_46933,N_44323,N_42836);
nor U46934 (N_46934,N_42664,N_43550);
or U46935 (N_46935,N_43882,N_43344);
or U46936 (N_46936,N_44168,N_43045);
xor U46937 (N_46937,N_44067,N_43891);
nand U46938 (N_46938,N_43428,N_43423);
nand U46939 (N_46939,N_42732,N_43495);
xor U46940 (N_46940,N_43407,N_44188);
xnor U46941 (N_46941,N_43524,N_42537);
nand U46942 (N_46942,N_44368,N_42846);
or U46943 (N_46943,N_42512,N_43366);
nor U46944 (N_46944,N_44336,N_43722);
xnor U46945 (N_46945,N_44276,N_42648);
nor U46946 (N_46946,N_44380,N_43052);
xor U46947 (N_46947,N_43792,N_42876);
xor U46948 (N_46948,N_43045,N_42705);
and U46949 (N_46949,N_44834,N_44463);
nor U46950 (N_46950,N_43283,N_44290);
nor U46951 (N_46951,N_43667,N_43487);
xor U46952 (N_46952,N_44872,N_42666);
nand U46953 (N_46953,N_43459,N_43670);
xnor U46954 (N_46954,N_44787,N_43322);
and U46955 (N_46955,N_42511,N_44880);
or U46956 (N_46956,N_43088,N_44260);
or U46957 (N_46957,N_43816,N_44914);
or U46958 (N_46958,N_42868,N_44035);
or U46959 (N_46959,N_42539,N_44151);
nand U46960 (N_46960,N_43499,N_43189);
or U46961 (N_46961,N_43682,N_44298);
or U46962 (N_46962,N_44523,N_44336);
or U46963 (N_46963,N_42961,N_43323);
nor U46964 (N_46964,N_44931,N_42926);
and U46965 (N_46965,N_42932,N_42787);
and U46966 (N_46966,N_43282,N_44745);
xor U46967 (N_46967,N_44251,N_44487);
nand U46968 (N_46968,N_44572,N_44982);
or U46969 (N_46969,N_43976,N_43595);
nor U46970 (N_46970,N_43717,N_43018);
or U46971 (N_46971,N_43644,N_44491);
nand U46972 (N_46972,N_43100,N_43053);
or U46973 (N_46973,N_43643,N_44310);
nor U46974 (N_46974,N_43018,N_42551);
xor U46975 (N_46975,N_44722,N_44437);
nor U46976 (N_46976,N_43004,N_43836);
xor U46977 (N_46977,N_44605,N_44186);
and U46978 (N_46978,N_42647,N_42751);
or U46979 (N_46979,N_44179,N_44518);
xnor U46980 (N_46980,N_43353,N_44553);
and U46981 (N_46981,N_43578,N_44689);
nor U46982 (N_46982,N_44728,N_44735);
and U46983 (N_46983,N_43621,N_44980);
and U46984 (N_46984,N_44736,N_44563);
or U46985 (N_46985,N_42826,N_42545);
nor U46986 (N_46986,N_44267,N_42839);
nand U46987 (N_46987,N_43948,N_44379);
and U46988 (N_46988,N_44194,N_44511);
or U46989 (N_46989,N_43525,N_42871);
nand U46990 (N_46990,N_42514,N_44282);
nand U46991 (N_46991,N_43120,N_44383);
or U46992 (N_46992,N_42758,N_44867);
xor U46993 (N_46993,N_44197,N_44753);
xnor U46994 (N_46994,N_44425,N_44090);
xor U46995 (N_46995,N_42559,N_43195);
nor U46996 (N_46996,N_44007,N_44405);
or U46997 (N_46997,N_44038,N_42654);
and U46998 (N_46998,N_43980,N_42941);
and U46999 (N_46999,N_44013,N_44211);
nand U47000 (N_47000,N_44927,N_43565);
and U47001 (N_47001,N_43284,N_44030);
nor U47002 (N_47002,N_43704,N_42998);
or U47003 (N_47003,N_43728,N_43791);
nor U47004 (N_47004,N_43844,N_44735);
or U47005 (N_47005,N_42658,N_42889);
nand U47006 (N_47006,N_44704,N_43776);
xnor U47007 (N_47007,N_43443,N_43776);
xnor U47008 (N_47008,N_43465,N_43020);
or U47009 (N_47009,N_42724,N_43493);
nor U47010 (N_47010,N_44646,N_43137);
nand U47011 (N_47011,N_42827,N_42790);
or U47012 (N_47012,N_42780,N_43564);
and U47013 (N_47013,N_42598,N_43393);
or U47014 (N_47014,N_42651,N_44337);
or U47015 (N_47015,N_43171,N_44596);
xnor U47016 (N_47016,N_44932,N_43964);
nor U47017 (N_47017,N_44281,N_42740);
nor U47018 (N_47018,N_44023,N_44551);
and U47019 (N_47019,N_44898,N_44534);
nor U47020 (N_47020,N_42922,N_43190);
xnor U47021 (N_47021,N_43396,N_44408);
nand U47022 (N_47022,N_44682,N_43142);
xor U47023 (N_47023,N_42895,N_44454);
xor U47024 (N_47024,N_42718,N_44582);
xnor U47025 (N_47025,N_43105,N_43491);
xnor U47026 (N_47026,N_44433,N_43660);
or U47027 (N_47027,N_44901,N_44001);
or U47028 (N_47028,N_44867,N_43622);
and U47029 (N_47029,N_43906,N_43752);
and U47030 (N_47030,N_43839,N_43925);
xor U47031 (N_47031,N_43415,N_42824);
or U47032 (N_47032,N_43842,N_42534);
or U47033 (N_47033,N_42802,N_44616);
or U47034 (N_47034,N_42718,N_42867);
or U47035 (N_47035,N_44794,N_44814);
or U47036 (N_47036,N_42677,N_43807);
and U47037 (N_47037,N_44850,N_43749);
or U47038 (N_47038,N_43330,N_43251);
nor U47039 (N_47039,N_43529,N_44442);
nor U47040 (N_47040,N_44941,N_43409);
and U47041 (N_47041,N_43010,N_42546);
nor U47042 (N_47042,N_43210,N_44986);
nand U47043 (N_47043,N_44876,N_42663);
nor U47044 (N_47044,N_42811,N_42606);
xnor U47045 (N_47045,N_43401,N_42598);
xnor U47046 (N_47046,N_44215,N_43111);
nand U47047 (N_47047,N_42886,N_43011);
nand U47048 (N_47048,N_44965,N_44957);
or U47049 (N_47049,N_43511,N_43309);
xnor U47050 (N_47050,N_43355,N_43934);
xnor U47051 (N_47051,N_43953,N_42722);
or U47052 (N_47052,N_44637,N_44399);
nor U47053 (N_47053,N_43058,N_44399);
nand U47054 (N_47054,N_43607,N_44415);
nor U47055 (N_47055,N_44023,N_43735);
or U47056 (N_47056,N_44162,N_43872);
nand U47057 (N_47057,N_43347,N_44284);
xnor U47058 (N_47058,N_44730,N_44024);
xor U47059 (N_47059,N_44005,N_43011);
nor U47060 (N_47060,N_42833,N_44318);
nand U47061 (N_47061,N_42748,N_42774);
and U47062 (N_47062,N_44793,N_43251);
xnor U47063 (N_47063,N_43077,N_43811);
or U47064 (N_47064,N_44234,N_43964);
and U47065 (N_47065,N_43909,N_43356);
and U47066 (N_47066,N_43974,N_44114);
and U47067 (N_47067,N_42792,N_42794);
nand U47068 (N_47068,N_43027,N_42719);
or U47069 (N_47069,N_42545,N_43743);
xnor U47070 (N_47070,N_44514,N_44971);
nor U47071 (N_47071,N_43099,N_42840);
xnor U47072 (N_47072,N_43401,N_44959);
or U47073 (N_47073,N_43392,N_44795);
nand U47074 (N_47074,N_42842,N_43283);
nand U47075 (N_47075,N_42537,N_44995);
nor U47076 (N_47076,N_43477,N_43784);
nor U47077 (N_47077,N_42896,N_44378);
and U47078 (N_47078,N_44309,N_42613);
nand U47079 (N_47079,N_42560,N_43945);
nor U47080 (N_47080,N_43185,N_44002);
and U47081 (N_47081,N_43905,N_42760);
nor U47082 (N_47082,N_43858,N_42773);
or U47083 (N_47083,N_42914,N_44881);
nand U47084 (N_47084,N_44152,N_43352);
nand U47085 (N_47085,N_43782,N_44335);
xor U47086 (N_47086,N_43997,N_43302);
xor U47087 (N_47087,N_44778,N_44726);
or U47088 (N_47088,N_44713,N_42672);
and U47089 (N_47089,N_43666,N_42877);
or U47090 (N_47090,N_44128,N_43214);
nand U47091 (N_47091,N_43527,N_44343);
xor U47092 (N_47092,N_42541,N_44607);
nor U47093 (N_47093,N_43957,N_42986);
nand U47094 (N_47094,N_43484,N_44067);
xor U47095 (N_47095,N_44379,N_44439);
xnor U47096 (N_47096,N_44958,N_43770);
nor U47097 (N_47097,N_42886,N_42688);
nor U47098 (N_47098,N_42638,N_43671);
nor U47099 (N_47099,N_42960,N_42859);
or U47100 (N_47100,N_44662,N_44011);
or U47101 (N_47101,N_44522,N_43336);
nor U47102 (N_47102,N_43020,N_44562);
nor U47103 (N_47103,N_44183,N_44482);
xnor U47104 (N_47104,N_43805,N_42919);
xor U47105 (N_47105,N_44077,N_42695);
nand U47106 (N_47106,N_44082,N_44688);
and U47107 (N_47107,N_43761,N_43103);
and U47108 (N_47108,N_42729,N_43483);
nand U47109 (N_47109,N_44505,N_43631);
or U47110 (N_47110,N_42819,N_44330);
xor U47111 (N_47111,N_43398,N_43871);
and U47112 (N_47112,N_44219,N_44759);
xnor U47113 (N_47113,N_44640,N_42545);
nand U47114 (N_47114,N_44111,N_43895);
nand U47115 (N_47115,N_43042,N_44748);
or U47116 (N_47116,N_42817,N_43570);
nand U47117 (N_47117,N_42605,N_44732);
or U47118 (N_47118,N_44582,N_43975);
and U47119 (N_47119,N_43175,N_43469);
or U47120 (N_47120,N_44210,N_43172);
and U47121 (N_47121,N_44363,N_44395);
or U47122 (N_47122,N_43828,N_43479);
or U47123 (N_47123,N_44139,N_43774);
nor U47124 (N_47124,N_43329,N_43485);
or U47125 (N_47125,N_42517,N_42649);
or U47126 (N_47126,N_44791,N_43250);
nand U47127 (N_47127,N_42951,N_44475);
nand U47128 (N_47128,N_44349,N_42674);
nand U47129 (N_47129,N_42509,N_42751);
or U47130 (N_47130,N_44068,N_44392);
xor U47131 (N_47131,N_44319,N_43615);
nand U47132 (N_47132,N_44788,N_44030);
nor U47133 (N_47133,N_43213,N_44392);
nor U47134 (N_47134,N_43018,N_44187);
nand U47135 (N_47135,N_44344,N_43298);
xnor U47136 (N_47136,N_44835,N_42662);
or U47137 (N_47137,N_43204,N_43096);
xnor U47138 (N_47138,N_43133,N_44766);
or U47139 (N_47139,N_43608,N_43651);
nand U47140 (N_47140,N_44934,N_42924);
nor U47141 (N_47141,N_44608,N_44759);
nand U47142 (N_47142,N_43661,N_43684);
nand U47143 (N_47143,N_44307,N_44987);
xor U47144 (N_47144,N_44960,N_43573);
nand U47145 (N_47145,N_43830,N_43753);
xor U47146 (N_47146,N_44305,N_44222);
nor U47147 (N_47147,N_43204,N_44953);
xor U47148 (N_47148,N_44805,N_44881);
and U47149 (N_47149,N_43802,N_44689);
and U47150 (N_47150,N_42911,N_43937);
nor U47151 (N_47151,N_43401,N_44964);
nand U47152 (N_47152,N_43749,N_44243);
nand U47153 (N_47153,N_43152,N_44424);
or U47154 (N_47154,N_43318,N_44091);
xnor U47155 (N_47155,N_43715,N_44261);
and U47156 (N_47156,N_43020,N_42981);
or U47157 (N_47157,N_42862,N_43131);
xor U47158 (N_47158,N_43240,N_43102);
nor U47159 (N_47159,N_42791,N_43391);
nand U47160 (N_47160,N_43972,N_44673);
nand U47161 (N_47161,N_43999,N_42595);
and U47162 (N_47162,N_44708,N_43197);
nor U47163 (N_47163,N_44583,N_44002);
nand U47164 (N_47164,N_43499,N_43536);
or U47165 (N_47165,N_43129,N_44220);
or U47166 (N_47166,N_44934,N_44600);
and U47167 (N_47167,N_43785,N_42899);
or U47168 (N_47168,N_44846,N_44473);
nor U47169 (N_47169,N_43203,N_43429);
and U47170 (N_47170,N_43267,N_43610);
nor U47171 (N_47171,N_44268,N_42565);
and U47172 (N_47172,N_44354,N_43819);
or U47173 (N_47173,N_43163,N_44269);
nand U47174 (N_47174,N_44913,N_43676);
xnor U47175 (N_47175,N_44274,N_44099);
nand U47176 (N_47176,N_42519,N_43493);
xor U47177 (N_47177,N_43357,N_44194);
nand U47178 (N_47178,N_43206,N_42598);
nor U47179 (N_47179,N_43804,N_44581);
or U47180 (N_47180,N_42864,N_43679);
or U47181 (N_47181,N_42548,N_43850);
nor U47182 (N_47182,N_44456,N_42726);
nor U47183 (N_47183,N_44825,N_43565);
nand U47184 (N_47184,N_44826,N_42806);
or U47185 (N_47185,N_44745,N_44626);
xor U47186 (N_47186,N_44217,N_43494);
xnor U47187 (N_47187,N_43122,N_43751);
or U47188 (N_47188,N_44294,N_43440);
xor U47189 (N_47189,N_42862,N_44082);
or U47190 (N_47190,N_43344,N_43829);
or U47191 (N_47191,N_42687,N_43643);
and U47192 (N_47192,N_44443,N_44890);
xnor U47193 (N_47193,N_43302,N_42598);
nand U47194 (N_47194,N_43244,N_43965);
nand U47195 (N_47195,N_44137,N_43843);
xor U47196 (N_47196,N_43186,N_44125);
nor U47197 (N_47197,N_43542,N_43416);
nand U47198 (N_47198,N_44238,N_43242);
nor U47199 (N_47199,N_43081,N_42810);
xnor U47200 (N_47200,N_44779,N_43607);
xor U47201 (N_47201,N_44903,N_43072);
or U47202 (N_47202,N_44974,N_43258);
and U47203 (N_47203,N_43236,N_43811);
and U47204 (N_47204,N_42933,N_44902);
nor U47205 (N_47205,N_43828,N_43190);
or U47206 (N_47206,N_44468,N_44074);
nor U47207 (N_47207,N_43786,N_44490);
or U47208 (N_47208,N_43721,N_42524);
or U47209 (N_47209,N_43984,N_44709);
xnor U47210 (N_47210,N_43986,N_43769);
nand U47211 (N_47211,N_43026,N_42752);
and U47212 (N_47212,N_44079,N_42920);
nor U47213 (N_47213,N_43414,N_44729);
nand U47214 (N_47214,N_44977,N_44803);
nand U47215 (N_47215,N_42716,N_44496);
xor U47216 (N_47216,N_43698,N_42818);
xor U47217 (N_47217,N_43599,N_44190);
nand U47218 (N_47218,N_43176,N_43189);
and U47219 (N_47219,N_44270,N_43200);
nand U47220 (N_47220,N_43465,N_42621);
and U47221 (N_47221,N_43483,N_44617);
nand U47222 (N_47222,N_44040,N_43544);
xor U47223 (N_47223,N_43135,N_44811);
xor U47224 (N_47224,N_44529,N_43010);
or U47225 (N_47225,N_44135,N_44356);
xnor U47226 (N_47226,N_42579,N_43652);
or U47227 (N_47227,N_43344,N_44270);
or U47228 (N_47228,N_42999,N_43878);
xor U47229 (N_47229,N_43477,N_43907);
and U47230 (N_47230,N_43087,N_44178);
nor U47231 (N_47231,N_42511,N_42934);
and U47232 (N_47232,N_42768,N_44574);
nor U47233 (N_47233,N_42760,N_42684);
or U47234 (N_47234,N_44600,N_43739);
and U47235 (N_47235,N_44236,N_44347);
nor U47236 (N_47236,N_44991,N_43139);
nor U47237 (N_47237,N_43865,N_44215);
xor U47238 (N_47238,N_42603,N_42988);
nand U47239 (N_47239,N_42726,N_44976);
nor U47240 (N_47240,N_43992,N_42521);
and U47241 (N_47241,N_43962,N_43639);
and U47242 (N_47242,N_42703,N_43690);
and U47243 (N_47243,N_43550,N_44418);
and U47244 (N_47244,N_42666,N_43479);
or U47245 (N_47245,N_43294,N_43610);
xnor U47246 (N_47246,N_44821,N_43366);
nand U47247 (N_47247,N_43916,N_44034);
xnor U47248 (N_47248,N_44427,N_42828);
nor U47249 (N_47249,N_43998,N_42989);
xor U47250 (N_47250,N_44689,N_44331);
and U47251 (N_47251,N_44646,N_42918);
xnor U47252 (N_47252,N_44336,N_44460);
or U47253 (N_47253,N_43069,N_43187);
nor U47254 (N_47254,N_43943,N_42687);
and U47255 (N_47255,N_43715,N_44842);
xor U47256 (N_47256,N_44719,N_44525);
nor U47257 (N_47257,N_44857,N_42729);
and U47258 (N_47258,N_42592,N_43831);
and U47259 (N_47259,N_44747,N_44957);
xnor U47260 (N_47260,N_42617,N_42608);
or U47261 (N_47261,N_43681,N_43977);
and U47262 (N_47262,N_43005,N_44027);
and U47263 (N_47263,N_44977,N_44548);
or U47264 (N_47264,N_43927,N_44921);
nand U47265 (N_47265,N_43663,N_44787);
or U47266 (N_47266,N_44681,N_43372);
nand U47267 (N_47267,N_43539,N_42502);
xnor U47268 (N_47268,N_43729,N_43505);
and U47269 (N_47269,N_42770,N_43142);
or U47270 (N_47270,N_44277,N_43301);
nand U47271 (N_47271,N_43467,N_43107);
and U47272 (N_47272,N_44311,N_43547);
nor U47273 (N_47273,N_44895,N_42946);
nor U47274 (N_47274,N_44268,N_44084);
or U47275 (N_47275,N_42962,N_43643);
or U47276 (N_47276,N_44870,N_44251);
nand U47277 (N_47277,N_43563,N_44541);
nand U47278 (N_47278,N_44427,N_43522);
xnor U47279 (N_47279,N_43003,N_43364);
xnor U47280 (N_47280,N_44456,N_43206);
xor U47281 (N_47281,N_44435,N_43591);
or U47282 (N_47282,N_43432,N_43690);
nor U47283 (N_47283,N_44460,N_44986);
xor U47284 (N_47284,N_44095,N_44196);
xor U47285 (N_47285,N_43530,N_44324);
or U47286 (N_47286,N_44087,N_42603);
and U47287 (N_47287,N_44292,N_43047);
nand U47288 (N_47288,N_44118,N_43950);
xnor U47289 (N_47289,N_43204,N_44732);
xnor U47290 (N_47290,N_44419,N_44969);
nand U47291 (N_47291,N_44008,N_43327);
or U47292 (N_47292,N_43048,N_44062);
and U47293 (N_47293,N_42719,N_44659);
or U47294 (N_47294,N_43037,N_42548);
xor U47295 (N_47295,N_43683,N_44262);
xnor U47296 (N_47296,N_42999,N_44842);
nand U47297 (N_47297,N_44681,N_44694);
xor U47298 (N_47298,N_44982,N_44527);
nand U47299 (N_47299,N_44503,N_43271);
or U47300 (N_47300,N_44165,N_43138);
or U47301 (N_47301,N_42577,N_42875);
or U47302 (N_47302,N_44119,N_43142);
or U47303 (N_47303,N_44109,N_42955);
nand U47304 (N_47304,N_42909,N_44664);
nor U47305 (N_47305,N_44485,N_43283);
nand U47306 (N_47306,N_43463,N_44714);
or U47307 (N_47307,N_43057,N_44434);
or U47308 (N_47308,N_44234,N_44713);
xor U47309 (N_47309,N_44022,N_43750);
xor U47310 (N_47310,N_44791,N_44019);
or U47311 (N_47311,N_43317,N_43478);
or U47312 (N_47312,N_43576,N_43255);
nand U47313 (N_47313,N_43248,N_42833);
xor U47314 (N_47314,N_44342,N_42753);
and U47315 (N_47315,N_44754,N_44067);
xor U47316 (N_47316,N_44447,N_42940);
nor U47317 (N_47317,N_42824,N_44594);
nor U47318 (N_47318,N_44629,N_43124);
xnor U47319 (N_47319,N_43958,N_42980);
and U47320 (N_47320,N_43011,N_43320);
nor U47321 (N_47321,N_44511,N_42944);
nor U47322 (N_47322,N_43035,N_43480);
nand U47323 (N_47323,N_43332,N_42912);
or U47324 (N_47324,N_44013,N_44681);
nor U47325 (N_47325,N_42882,N_44181);
or U47326 (N_47326,N_43717,N_43756);
nand U47327 (N_47327,N_43323,N_42667);
nor U47328 (N_47328,N_44235,N_43553);
or U47329 (N_47329,N_44627,N_43540);
nand U47330 (N_47330,N_43289,N_43141);
nand U47331 (N_47331,N_44501,N_43661);
or U47332 (N_47332,N_43722,N_42664);
nand U47333 (N_47333,N_44672,N_44679);
or U47334 (N_47334,N_43162,N_44859);
and U47335 (N_47335,N_44147,N_43523);
nand U47336 (N_47336,N_44527,N_44041);
nand U47337 (N_47337,N_44626,N_44074);
or U47338 (N_47338,N_42538,N_42887);
nor U47339 (N_47339,N_44153,N_43153);
nand U47340 (N_47340,N_42772,N_42884);
nand U47341 (N_47341,N_44191,N_42602);
or U47342 (N_47342,N_44159,N_42760);
xnor U47343 (N_47343,N_44773,N_42658);
and U47344 (N_47344,N_43801,N_44077);
nand U47345 (N_47345,N_43256,N_43965);
or U47346 (N_47346,N_44699,N_44959);
or U47347 (N_47347,N_42987,N_44605);
and U47348 (N_47348,N_43972,N_43696);
or U47349 (N_47349,N_43971,N_42607);
nand U47350 (N_47350,N_42710,N_43349);
nand U47351 (N_47351,N_44052,N_43496);
or U47352 (N_47352,N_44804,N_44841);
nand U47353 (N_47353,N_44127,N_44403);
nor U47354 (N_47354,N_43036,N_42924);
and U47355 (N_47355,N_44221,N_42761);
and U47356 (N_47356,N_44845,N_42789);
nor U47357 (N_47357,N_44148,N_44564);
or U47358 (N_47358,N_44488,N_44582);
or U47359 (N_47359,N_43005,N_44484);
or U47360 (N_47360,N_44999,N_43359);
nand U47361 (N_47361,N_43792,N_44916);
nor U47362 (N_47362,N_42869,N_43139);
or U47363 (N_47363,N_44088,N_43021);
nor U47364 (N_47364,N_43887,N_44624);
and U47365 (N_47365,N_42952,N_44568);
xnor U47366 (N_47366,N_44014,N_44774);
nor U47367 (N_47367,N_43061,N_42555);
nand U47368 (N_47368,N_44680,N_44117);
and U47369 (N_47369,N_42619,N_44315);
nand U47370 (N_47370,N_44836,N_43439);
or U47371 (N_47371,N_42561,N_44513);
or U47372 (N_47372,N_44289,N_42708);
nor U47373 (N_47373,N_44236,N_43800);
and U47374 (N_47374,N_42749,N_44102);
xor U47375 (N_47375,N_43979,N_42954);
xor U47376 (N_47376,N_44911,N_43986);
nand U47377 (N_47377,N_44203,N_43015);
and U47378 (N_47378,N_43641,N_44695);
and U47379 (N_47379,N_43831,N_44120);
or U47380 (N_47380,N_44287,N_42952);
or U47381 (N_47381,N_43708,N_44724);
nor U47382 (N_47382,N_42929,N_43070);
nand U47383 (N_47383,N_43262,N_43948);
or U47384 (N_47384,N_44646,N_44359);
and U47385 (N_47385,N_43787,N_42719);
or U47386 (N_47386,N_44448,N_43595);
or U47387 (N_47387,N_43724,N_44379);
xor U47388 (N_47388,N_42925,N_44152);
xor U47389 (N_47389,N_44088,N_42628);
or U47390 (N_47390,N_44710,N_42604);
nand U47391 (N_47391,N_44233,N_44650);
xor U47392 (N_47392,N_44526,N_42573);
nor U47393 (N_47393,N_44478,N_44399);
nand U47394 (N_47394,N_44898,N_43851);
nand U47395 (N_47395,N_42993,N_43310);
xnor U47396 (N_47396,N_44713,N_44490);
nor U47397 (N_47397,N_44904,N_43469);
xnor U47398 (N_47398,N_43036,N_44808);
nor U47399 (N_47399,N_43438,N_42636);
nand U47400 (N_47400,N_42986,N_44436);
and U47401 (N_47401,N_42691,N_43243);
xnor U47402 (N_47402,N_44299,N_43769);
nand U47403 (N_47403,N_42907,N_43397);
xor U47404 (N_47404,N_44928,N_42544);
or U47405 (N_47405,N_44878,N_42592);
nor U47406 (N_47406,N_44150,N_44602);
or U47407 (N_47407,N_43378,N_44948);
and U47408 (N_47408,N_44233,N_44664);
nor U47409 (N_47409,N_43142,N_44440);
or U47410 (N_47410,N_44735,N_44298);
and U47411 (N_47411,N_43953,N_42702);
nand U47412 (N_47412,N_43552,N_44595);
xnor U47413 (N_47413,N_44870,N_44262);
and U47414 (N_47414,N_43962,N_43635);
nand U47415 (N_47415,N_44644,N_42719);
and U47416 (N_47416,N_44561,N_43885);
or U47417 (N_47417,N_43415,N_44702);
and U47418 (N_47418,N_43873,N_43843);
or U47419 (N_47419,N_43572,N_44867);
and U47420 (N_47420,N_42652,N_42645);
xnor U47421 (N_47421,N_43366,N_44186);
or U47422 (N_47422,N_44812,N_43205);
xor U47423 (N_47423,N_43887,N_43235);
nand U47424 (N_47424,N_44287,N_42842);
and U47425 (N_47425,N_44080,N_44928);
xnor U47426 (N_47426,N_43360,N_44795);
xor U47427 (N_47427,N_44294,N_43275);
xor U47428 (N_47428,N_44196,N_43739);
nor U47429 (N_47429,N_43697,N_44627);
or U47430 (N_47430,N_43161,N_43203);
or U47431 (N_47431,N_44510,N_42958);
or U47432 (N_47432,N_44568,N_43425);
nor U47433 (N_47433,N_44778,N_44861);
nor U47434 (N_47434,N_43027,N_44020);
nor U47435 (N_47435,N_44288,N_42672);
nand U47436 (N_47436,N_43292,N_44336);
nor U47437 (N_47437,N_43793,N_43064);
nor U47438 (N_47438,N_42521,N_43299);
xor U47439 (N_47439,N_44312,N_44203);
and U47440 (N_47440,N_42732,N_44526);
xnor U47441 (N_47441,N_43029,N_44774);
nand U47442 (N_47442,N_43082,N_44902);
nor U47443 (N_47443,N_43315,N_43222);
or U47444 (N_47444,N_44405,N_42894);
and U47445 (N_47445,N_43311,N_43539);
or U47446 (N_47446,N_44171,N_44729);
or U47447 (N_47447,N_44508,N_44213);
nand U47448 (N_47448,N_44548,N_44078);
or U47449 (N_47449,N_43680,N_44335);
nand U47450 (N_47450,N_43871,N_44596);
xnor U47451 (N_47451,N_44959,N_42559);
nand U47452 (N_47452,N_44623,N_43848);
and U47453 (N_47453,N_44103,N_44654);
xor U47454 (N_47454,N_44168,N_44761);
xor U47455 (N_47455,N_43706,N_43030);
or U47456 (N_47456,N_44196,N_44049);
and U47457 (N_47457,N_44214,N_44012);
nor U47458 (N_47458,N_44662,N_43309);
nand U47459 (N_47459,N_43592,N_43653);
xnor U47460 (N_47460,N_43102,N_42995);
xnor U47461 (N_47461,N_44746,N_42974);
nor U47462 (N_47462,N_42618,N_42919);
xor U47463 (N_47463,N_44112,N_44596);
nand U47464 (N_47464,N_44205,N_44547);
or U47465 (N_47465,N_44409,N_42989);
or U47466 (N_47466,N_43275,N_43369);
or U47467 (N_47467,N_43849,N_43371);
nor U47468 (N_47468,N_43061,N_43223);
nand U47469 (N_47469,N_42937,N_42771);
and U47470 (N_47470,N_43429,N_44016);
xnor U47471 (N_47471,N_44069,N_42942);
nor U47472 (N_47472,N_44519,N_43949);
xor U47473 (N_47473,N_42973,N_44435);
nand U47474 (N_47474,N_43304,N_43362);
nand U47475 (N_47475,N_43845,N_43953);
or U47476 (N_47476,N_43157,N_42501);
and U47477 (N_47477,N_42618,N_44549);
nand U47478 (N_47478,N_43263,N_42569);
nand U47479 (N_47479,N_42552,N_43871);
nand U47480 (N_47480,N_44610,N_44702);
xnor U47481 (N_47481,N_44430,N_44416);
and U47482 (N_47482,N_43443,N_43529);
xnor U47483 (N_47483,N_44776,N_44940);
xor U47484 (N_47484,N_44967,N_42538);
nand U47485 (N_47485,N_43821,N_43933);
and U47486 (N_47486,N_44012,N_43482);
or U47487 (N_47487,N_42585,N_42964);
xor U47488 (N_47488,N_43441,N_42513);
xor U47489 (N_47489,N_43916,N_42813);
nand U47490 (N_47490,N_44370,N_43549);
and U47491 (N_47491,N_44865,N_44871);
nor U47492 (N_47492,N_43103,N_43998);
nor U47493 (N_47493,N_44830,N_42677);
xor U47494 (N_47494,N_44783,N_42756);
xnor U47495 (N_47495,N_43787,N_42810);
and U47496 (N_47496,N_43702,N_42638);
nor U47497 (N_47497,N_44315,N_42592);
or U47498 (N_47498,N_44984,N_42872);
or U47499 (N_47499,N_42557,N_44788);
or U47500 (N_47500,N_45559,N_46302);
nor U47501 (N_47501,N_46583,N_47379);
or U47502 (N_47502,N_46428,N_46089);
and U47503 (N_47503,N_47304,N_45157);
nand U47504 (N_47504,N_47404,N_45216);
nor U47505 (N_47505,N_46957,N_45369);
nand U47506 (N_47506,N_46550,N_46275);
nor U47507 (N_47507,N_47235,N_46714);
xor U47508 (N_47508,N_46959,N_47424);
and U47509 (N_47509,N_47148,N_47043);
nand U47510 (N_47510,N_45373,N_46344);
or U47511 (N_47511,N_45043,N_46857);
nand U47512 (N_47512,N_45167,N_46338);
xnor U47513 (N_47513,N_46417,N_46877);
nor U47514 (N_47514,N_45553,N_45292);
or U47515 (N_47515,N_46538,N_45358);
and U47516 (N_47516,N_47498,N_46005);
nor U47517 (N_47517,N_47056,N_46009);
xor U47518 (N_47518,N_46331,N_45789);
and U47519 (N_47519,N_47029,N_47422);
or U47520 (N_47520,N_45323,N_45385);
or U47521 (N_47521,N_46415,N_45391);
nor U47522 (N_47522,N_45648,N_46590);
xor U47523 (N_47523,N_45131,N_46732);
nand U47524 (N_47524,N_45837,N_45341);
and U47525 (N_47525,N_47191,N_47154);
and U47526 (N_47526,N_45832,N_46214);
xor U47527 (N_47527,N_45602,N_46175);
xor U47528 (N_47528,N_46266,N_45153);
xor U47529 (N_47529,N_46473,N_47131);
and U47530 (N_47530,N_46893,N_45546);
nor U47531 (N_47531,N_45860,N_46207);
and U47532 (N_47532,N_45498,N_47409);
xor U47533 (N_47533,N_46662,N_45245);
nand U47534 (N_47534,N_47085,N_47139);
nand U47535 (N_47535,N_46357,N_46804);
nor U47536 (N_47536,N_47201,N_45692);
or U47537 (N_47537,N_45410,N_45721);
or U47538 (N_47538,N_46462,N_46416);
nor U47539 (N_47539,N_46004,N_46599);
or U47540 (N_47540,N_45405,N_45886);
nor U47541 (N_47541,N_45751,N_45384);
xor U47542 (N_47542,N_45725,N_45739);
nand U47543 (N_47543,N_45618,N_47326);
nor U47544 (N_47544,N_45701,N_46573);
and U47545 (N_47545,N_46063,N_47062);
and U47546 (N_47546,N_46655,N_46674);
or U47547 (N_47547,N_47357,N_45394);
nor U47548 (N_47548,N_45379,N_46492);
nand U47549 (N_47549,N_46845,N_45044);
xnor U47550 (N_47550,N_46101,N_46306);
and U47551 (N_47551,N_45937,N_46847);
nand U47552 (N_47552,N_46489,N_45911);
or U47553 (N_47553,N_45927,N_45423);
and U47554 (N_47554,N_47183,N_46509);
and U47555 (N_47555,N_45647,N_45241);
nand U47556 (N_47556,N_45991,N_45398);
nor U47557 (N_47557,N_45197,N_46470);
and U47558 (N_47558,N_46634,N_47297);
and U47559 (N_47559,N_46665,N_47138);
or U47560 (N_47560,N_45168,N_45668);
and U47561 (N_47561,N_46361,N_46341);
nand U47562 (N_47562,N_46374,N_45412);
or U47563 (N_47563,N_45479,N_45383);
nor U47564 (N_47564,N_45427,N_47113);
or U47565 (N_47565,N_45687,N_46825);
and U47566 (N_47566,N_47008,N_45064);
and U47567 (N_47567,N_46245,N_45998);
or U47568 (N_47568,N_46312,N_46024);
nor U47569 (N_47569,N_45762,N_47316);
and U47570 (N_47570,N_45260,N_45110);
xor U47571 (N_47571,N_47038,N_46012);
and U47572 (N_47572,N_46441,N_45255);
xnor U47573 (N_47573,N_45368,N_46111);
and U47574 (N_47574,N_46649,N_46965);
xnor U47575 (N_47575,N_46181,N_45004);
nor U47576 (N_47576,N_45801,N_46973);
or U47577 (N_47577,N_45355,N_45339);
and U47578 (N_47578,N_46713,N_46057);
nor U47579 (N_47579,N_46272,N_45092);
and U47580 (N_47580,N_46777,N_45724);
and U47581 (N_47581,N_46353,N_47408);
nor U47582 (N_47582,N_46709,N_45758);
nand U47583 (N_47583,N_47109,N_47251);
and U47584 (N_47584,N_45613,N_46586);
xor U47585 (N_47585,N_46900,N_46928);
or U47586 (N_47586,N_45024,N_46767);
xor U47587 (N_47587,N_45716,N_46797);
and U47588 (N_47588,N_46578,N_46398);
nand U47589 (N_47589,N_46535,N_46083);
nand U47590 (N_47590,N_45612,N_45809);
xor U47591 (N_47591,N_46269,N_46966);
or U47592 (N_47592,N_45015,N_46947);
or U47593 (N_47593,N_46380,N_46017);
nand U47594 (N_47594,N_46739,N_45715);
and U47595 (N_47595,N_46407,N_47112);
xor U47596 (N_47596,N_47473,N_45430);
xnor U47597 (N_47597,N_45617,N_47333);
and U47598 (N_47598,N_47100,N_47446);
xor U47599 (N_47599,N_46846,N_47023);
or U47600 (N_47600,N_46090,N_45165);
and U47601 (N_47601,N_46678,N_46533);
or U47602 (N_47602,N_46025,N_47274);
and U47603 (N_47603,N_47472,N_47164);
or U47604 (N_47604,N_46629,N_46880);
and U47605 (N_47605,N_46442,N_47240);
nand U47606 (N_47606,N_47325,N_46799);
and U47607 (N_47607,N_46860,N_46367);
and U47608 (N_47608,N_45690,N_47035);
or U47609 (N_47609,N_47250,N_46593);
or U47610 (N_47610,N_45753,N_46477);
nor U47611 (N_47611,N_47057,N_45637);
and U47612 (N_47612,N_45859,N_45088);
nand U47613 (N_47613,N_45215,N_46179);
nand U47614 (N_47614,N_46562,N_45510);
xnor U47615 (N_47615,N_46680,N_45584);
xor U47616 (N_47616,N_46018,N_45773);
nand U47617 (N_47617,N_47241,N_46482);
or U47618 (N_47618,N_46373,N_46666);
or U47619 (N_47619,N_45528,N_46029);
xnor U47620 (N_47620,N_45626,N_46079);
and U47621 (N_47621,N_47026,N_47484);
nor U47622 (N_47622,N_47301,N_45611);
nor U47623 (N_47623,N_45306,N_47342);
xnor U47624 (N_47624,N_46359,N_47175);
or U47625 (N_47625,N_45743,N_45673);
and U47626 (N_47626,N_45416,N_46886);
or U47627 (N_47627,N_45776,N_47237);
xor U47628 (N_47628,N_45091,N_46393);
or U47629 (N_47629,N_47262,N_45465);
and U47630 (N_47630,N_45760,N_45041);
or U47631 (N_47631,N_46663,N_47293);
or U47632 (N_47632,N_45467,N_46040);
xor U47633 (N_47633,N_45146,N_45922);
nor U47634 (N_47634,N_46785,N_46042);
nor U47635 (N_47635,N_46980,N_45977);
and U47636 (N_47636,N_47416,N_46828);
and U47637 (N_47637,N_46355,N_47045);
nand U47638 (N_47638,N_46244,N_46466);
nand U47639 (N_47639,N_45349,N_45399);
nor U47640 (N_47640,N_47474,N_47218);
or U47641 (N_47641,N_45095,N_46127);
xor U47642 (N_47642,N_47127,N_45303);
and U47643 (N_47643,N_47445,N_46925);
nand U47644 (N_47644,N_46391,N_46765);
nand U47645 (N_47645,N_45364,N_46324);
nor U47646 (N_47646,N_47092,N_46459);
nor U47647 (N_47647,N_45328,N_47072);
or U47648 (N_47648,N_46708,N_45771);
nand U47649 (N_47649,N_45812,N_46484);
or U47650 (N_47650,N_47343,N_45950);
nor U47651 (N_47651,N_47168,N_47341);
nand U47652 (N_47652,N_45959,N_46003);
or U47653 (N_47653,N_46611,N_46604);
or U47654 (N_47654,N_46388,N_46745);
nand U47655 (N_47655,N_46279,N_46451);
xnor U47656 (N_47656,N_47011,N_46960);
or U47657 (N_47657,N_45443,N_45824);
or U47658 (N_47658,N_45065,N_45316);
nand U47659 (N_47659,N_46653,N_45769);
xor U47660 (N_47660,N_46171,N_46351);
nor U47661 (N_47661,N_45208,N_47243);
and U47662 (N_47662,N_46330,N_45718);
and U47663 (N_47663,N_47488,N_46201);
xnor U47664 (N_47664,N_45929,N_45754);
nand U47665 (N_47665,N_46711,N_46763);
or U47666 (N_47666,N_45939,N_45264);
and U47667 (N_47667,N_45363,N_47065);
xnor U47668 (N_47668,N_47377,N_46978);
nor U47669 (N_47669,N_45908,N_46199);
and U47670 (N_47670,N_45901,N_45074);
and U47671 (N_47671,N_46735,N_45943);
nor U47672 (N_47672,N_46682,N_46722);
and U47673 (N_47673,N_45890,N_46086);
xnor U47674 (N_47674,N_46782,N_46028);
nor U47675 (N_47675,N_46951,N_45190);
and U47676 (N_47676,N_45273,N_46850);
and U47677 (N_47677,N_46651,N_45548);
and U47678 (N_47678,N_46758,N_47486);
xor U47679 (N_47679,N_46231,N_45720);
and U47680 (N_47680,N_47153,N_46370);
or U47681 (N_47681,N_45630,N_47182);
nor U47682 (N_47682,N_45144,N_46157);
xnor U47683 (N_47683,N_46793,N_47346);
nor U47684 (N_47684,N_46814,N_45121);
nor U47685 (N_47685,N_45294,N_46532);
xnor U47686 (N_47686,N_46766,N_45527);
or U47687 (N_47687,N_45324,N_45037);
xnor U47688 (N_47688,N_47388,N_45605);
xor U47689 (N_47689,N_47137,N_45244);
nor U47690 (N_47690,N_46088,N_46411);
nand U47691 (N_47691,N_47354,N_46021);
and U47692 (N_47692,N_46555,N_45981);
nand U47693 (N_47693,N_45401,N_46729);
and U47694 (N_47694,N_46723,N_45547);
or U47695 (N_47695,N_46138,N_46117);
xnor U47696 (N_47696,N_45060,N_46588);
or U47697 (N_47697,N_45788,N_46750);
nor U47698 (N_47698,N_46239,N_46639);
xor U47699 (N_47699,N_45545,N_46871);
nand U47700 (N_47700,N_45409,N_45699);
xor U47701 (N_47701,N_47222,N_46483);
nor U47702 (N_47702,N_45912,N_47294);
or U47703 (N_47703,N_45456,N_45406);
xnor U47704 (N_47704,N_45470,N_46910);
xnor U47705 (N_47705,N_46360,N_47017);
and U47706 (N_47706,N_45402,N_46582);
or U47707 (N_47707,N_45787,N_45202);
nor U47708 (N_47708,N_45969,N_46443);
or U47709 (N_47709,N_47406,N_46200);
xnor U47710 (N_47710,N_45576,N_46541);
and U47711 (N_47711,N_45028,N_47344);
xnor U47712 (N_47712,N_47075,N_46703);
nor U47713 (N_47713,N_47120,N_45100);
nand U47714 (N_47714,N_45031,N_46223);
or U47715 (N_47715,N_46511,N_47454);
nor U47716 (N_47716,N_47081,N_47387);
nor U47717 (N_47717,N_46560,N_45330);
nand U47718 (N_47718,N_47279,N_45600);
or U47719 (N_47719,N_45257,N_45047);
nand U47720 (N_47720,N_46452,N_47275);
xor U47721 (N_47721,N_46383,N_45660);
or U47722 (N_47722,N_45871,N_45185);
and U47723 (N_47723,N_45694,N_46158);
and U47724 (N_47724,N_47156,N_45039);
nand U47725 (N_47725,N_45154,N_46051);
xnor U47726 (N_47726,N_45505,N_46876);
or U47727 (N_47727,N_46206,N_45813);
and U47728 (N_47728,N_45597,N_46493);
and U47729 (N_47729,N_47369,N_46320);
nor U47730 (N_47730,N_46196,N_47185);
or U47731 (N_47731,N_45652,N_45435);
xnor U47732 (N_47732,N_47285,N_46147);
and U47733 (N_47733,N_45176,N_46997);
and U47734 (N_47734,N_45863,N_47132);
or U47735 (N_47735,N_45962,N_45841);
or U47736 (N_47736,N_45371,N_46041);
and U47737 (N_47737,N_47264,N_45920);
or U47738 (N_47738,N_47124,N_45055);
or U47739 (N_47739,N_46553,N_47210);
nor U47740 (N_47740,N_46429,N_46019);
nand U47741 (N_47741,N_47329,N_45344);
nand U47742 (N_47742,N_46805,N_46636);
and U47743 (N_47743,N_46898,N_45102);
nor U47744 (N_47744,N_45661,N_46656);
or U47745 (N_47745,N_47298,N_46971);
nor U47746 (N_47746,N_45035,N_45086);
or U47747 (N_47747,N_46068,N_46508);
xnor U47748 (N_47748,N_47128,N_45595);
and U47749 (N_47749,N_46924,N_46494);
and U47750 (N_47750,N_45437,N_47234);
or U47751 (N_47751,N_46053,N_47111);
xnor U47752 (N_47752,N_46915,N_45233);
and U47753 (N_47753,N_45938,N_46323);
nand U47754 (N_47754,N_46140,N_45223);
and U47755 (N_47755,N_45537,N_46833);
nand U47756 (N_47756,N_45089,N_46851);
xnor U47757 (N_47757,N_47090,N_46290);
nor U47758 (N_47758,N_47373,N_45270);
nand U47759 (N_47759,N_46803,N_45816);
nand U47760 (N_47760,N_46187,N_46110);
or U47761 (N_47761,N_45217,N_46549);
nand U47762 (N_47762,N_46992,N_46528);
xnor U47763 (N_47763,N_45013,N_45454);
or U47764 (N_47764,N_45307,N_45194);
and U47765 (N_47765,N_46174,N_47493);
nand U47766 (N_47766,N_47031,N_46792);
or U47767 (N_47767,N_45432,N_47073);
or U47768 (N_47768,N_46237,N_46654);
and U47769 (N_47769,N_45823,N_45562);
nand U47770 (N_47770,N_47068,N_45972);
or U47771 (N_47771,N_47088,N_47082);
nor U47772 (N_47772,N_45261,N_45935);
xor U47773 (N_47773,N_46784,N_46093);
nand U47774 (N_47774,N_45071,N_45164);
nand U47775 (N_47775,N_45606,N_46534);
nand U47776 (N_47776,N_47260,N_46645);
nor U47777 (N_47777,N_46499,N_47295);
nand U47778 (N_47778,N_46826,N_45976);
xnor U47779 (N_47779,N_47159,N_46014);
and U47780 (N_47780,N_45830,N_46585);
xor U47781 (N_47781,N_46410,N_45755);
nand U47782 (N_47782,N_46524,N_45441);
and U47783 (N_47783,N_45332,N_47423);
nand U47784 (N_47784,N_46333,N_45192);
and U47785 (N_47785,N_45212,N_46354);
and U47786 (N_47786,N_46569,N_47270);
and U47787 (N_47787,N_47115,N_47007);
or U47788 (N_47788,N_46736,N_47303);
xor U47789 (N_47789,N_46630,N_45275);
or U47790 (N_47790,N_47282,N_47228);
xor U47791 (N_47791,N_46292,N_45209);
xor U47792 (N_47792,N_47126,N_47467);
nor U47793 (N_47793,N_47225,N_45892);
nor U47794 (N_47794,N_46406,N_47310);
nand U47795 (N_47795,N_45983,N_46632);
nand U47796 (N_47796,N_45101,N_46752);
and U47797 (N_47797,N_46761,N_47477);
nor U47798 (N_47798,N_45759,N_45382);
or U47799 (N_47799,N_46184,N_46764);
and U47800 (N_47800,N_47361,N_45442);
nor U47801 (N_47801,N_45234,N_45112);
nand U47802 (N_47802,N_45675,N_45504);
nor U47803 (N_47803,N_46095,N_46781);
or U47804 (N_47804,N_46375,N_45656);
xnor U47805 (N_47805,N_45726,N_45572);
nor U47806 (N_47806,N_45654,N_47058);
or U47807 (N_47807,N_45375,N_47078);
nand U47808 (N_47808,N_45968,N_46318);
nor U47809 (N_47809,N_45431,N_46186);
nor U47810 (N_47810,N_46397,N_46707);
nor U47811 (N_47811,N_46545,N_45677);
xor U47812 (N_47812,N_46035,N_46495);
xnor U47813 (N_47813,N_47267,N_45484);
or U47814 (N_47814,N_45978,N_47483);
and U47815 (N_47815,N_45887,N_45870);
nor U47816 (N_47816,N_46901,N_45624);
nor U47817 (N_47817,N_45475,N_45151);
xor U47818 (N_47818,N_45550,N_46888);
nor U47819 (N_47819,N_46685,N_46465);
nor U47820 (N_47820,N_46246,N_46334);
xor U47821 (N_47821,N_46883,N_47321);
or U47822 (N_47822,N_45644,N_45918);
or U47823 (N_47823,N_46536,N_47340);
nand U47824 (N_47824,N_47145,N_45666);
nor U47825 (N_47825,N_45714,N_45390);
xor U47826 (N_47826,N_45985,N_47427);
nand U47827 (N_47827,N_46497,N_46621);
xor U47828 (N_47828,N_45967,N_46969);
nand U47829 (N_47829,N_47380,N_45222);
xnor U47830 (N_47830,N_47269,N_46938);
and U47831 (N_47831,N_46249,N_47229);
xor U47832 (N_47832,N_46491,N_45356);
nand U47833 (N_47833,N_46011,N_47084);
and U47834 (N_47834,N_45469,N_45609);
xnor U47835 (N_47835,N_45766,N_46046);
nand U47836 (N_47836,N_45598,N_45669);
and U47837 (N_47837,N_46675,N_46133);
or U47838 (N_47838,N_47108,N_47475);
and U47839 (N_47839,N_47273,N_45036);
nor U47840 (N_47840,N_45949,N_47413);
and U47841 (N_47841,N_46658,N_46991);
and U47842 (N_47842,N_45542,N_45061);
nand U47843 (N_47843,N_45016,N_45747);
nor U47844 (N_47844,N_47162,N_45765);
or U47845 (N_47845,N_45227,N_47444);
nand U47846 (N_47846,N_46554,N_45891);
and U47847 (N_47847,N_46501,N_45796);
and U47848 (N_47848,N_45797,N_46975);
xnor U47849 (N_47849,N_45277,N_45732);
or U47850 (N_47850,N_47047,N_47314);
and U47851 (N_47851,N_45082,N_45560);
nor U47852 (N_47852,N_46219,N_45496);
nor U47853 (N_47853,N_46844,N_47188);
and U47854 (N_47854,N_47421,N_46648);
or U47855 (N_47855,N_45184,N_46882);
and U47856 (N_47856,N_46838,N_45784);
or U47857 (N_47857,N_47307,N_46574);
xor U47858 (N_47858,N_46413,N_45070);
or U47859 (N_47859,N_47348,N_47287);
xnor U47860 (N_47860,N_45018,N_45511);
xnor U47861 (N_47861,N_45899,N_45996);
and U47862 (N_47862,N_46071,N_46027);
nand U47863 (N_47863,N_47037,N_46638);
or U47864 (N_47864,N_46864,N_46669);
nand U47865 (N_47865,N_47048,N_46762);
or U47866 (N_47866,N_46660,N_45826);
nor U47867 (N_47867,N_45638,N_47214);
or U47868 (N_47868,N_46756,N_46222);
xor U47869 (N_47869,N_45093,N_46810);
xor U47870 (N_47870,N_47117,N_45632);
or U47871 (N_47871,N_47104,N_46015);
nand U47872 (N_47872,N_47125,N_45540);
nand U47873 (N_47873,N_46316,N_46748);
nor U47874 (N_47874,N_45236,N_46788);
and U47875 (N_47875,N_45116,N_45249);
nor U47876 (N_47876,N_45495,N_45351);
and U47877 (N_47877,N_46130,N_47179);
xnor U47878 (N_47878,N_46738,N_45536);
xor U47879 (N_47879,N_46007,N_46366);
nand U47880 (N_47880,N_46801,N_45099);
and U47881 (N_47881,N_46646,N_46791);
and U47882 (N_47882,N_47398,N_45200);
nor U47883 (N_47883,N_45928,N_45767);
and U47884 (N_47884,N_47381,N_46956);
or U47885 (N_47885,N_45608,N_46036);
xnor U47886 (N_47886,N_47049,N_46432);
nor U47887 (N_47887,N_45610,N_46234);
and U47888 (N_47888,N_45695,N_46218);
and U47889 (N_47889,N_46229,N_45683);
nor U47890 (N_47890,N_45161,N_46319);
nor U47891 (N_47891,N_45325,N_46044);
and U47892 (N_47892,N_45421,N_46902);
xnor U47893 (N_47893,N_46294,N_46163);
xnor U47894 (N_47894,N_46624,N_46558);
nand U47895 (N_47895,N_47118,N_47283);
and U47896 (N_47896,N_46304,N_46233);
xor U47897 (N_47897,N_45072,N_46150);
xnor U47898 (N_47898,N_46885,N_46379);
nor U47899 (N_47899,N_45247,N_47490);
xor U47900 (N_47900,N_47364,N_45338);
xor U47901 (N_47901,N_47453,N_47323);
nand U47902 (N_47902,N_46936,N_46387);
nor U47903 (N_47903,N_46148,N_46567);
and U47904 (N_47904,N_45111,N_45951);
xor U47905 (N_47905,N_46309,N_45874);
or U47906 (N_47906,N_45974,N_46125);
and U47907 (N_47907,N_46468,N_45287);
or U47908 (N_47908,N_45625,N_46724);
and U47909 (N_47909,N_45336,N_45119);
and U47910 (N_47910,N_45982,N_46235);
nand U47911 (N_47911,N_46185,N_47407);
nor U47912 (N_47912,N_45032,N_45627);
nand U47913 (N_47913,N_46409,N_45558);
nor U47914 (N_47914,N_46620,N_46070);
or U47915 (N_47915,N_47371,N_45388);
or U47916 (N_47916,N_45376,N_46808);
and U47917 (N_47917,N_46193,N_46710);
nor U47918 (N_47918,N_46463,N_45019);
nand U47919 (N_47919,N_45880,N_45569);
nand U47920 (N_47920,N_47394,N_45136);
nor U47921 (N_47921,N_47372,N_45295);
nor U47922 (N_47922,N_45076,N_45623);
xor U47923 (N_47923,N_47060,N_46225);
nand U47924 (N_47924,N_46920,N_45803);
nand U47925 (N_47925,N_46488,N_46631);
nand U47926 (N_47926,N_46109,N_46633);
xnor U47927 (N_47927,N_46287,N_47212);
xor U47928 (N_47928,N_45159,N_45895);
and U47929 (N_47929,N_45455,N_46208);
xor U47930 (N_47930,N_46480,N_45451);
nand U47931 (N_47931,N_45898,N_45709);
or U47932 (N_47932,N_46382,N_45252);
xnor U47933 (N_47933,N_45757,N_45298);
nor U47934 (N_47934,N_46099,N_46146);
or U47935 (N_47935,N_45583,N_47174);
nand U47936 (N_47936,N_46809,N_46267);
nor U47937 (N_47937,N_46092,N_47155);
nor U47938 (N_47938,N_46173,N_45053);
or U47939 (N_47939,N_46929,N_45218);
nor U47940 (N_47940,N_45027,N_46345);
xor U47941 (N_47941,N_46356,N_45414);
nand U47942 (N_47942,N_45942,N_47176);
xor U47943 (N_47943,N_46328,N_45593);
or U47944 (N_47944,N_47206,N_47116);
xor U47945 (N_47945,N_46546,N_46265);
nor U47946 (N_47946,N_45001,N_45744);
nand U47947 (N_47947,N_47390,N_45806);
or U47948 (N_47948,N_45662,N_46444);
or U47949 (N_47949,N_46065,N_45335);
and U47950 (N_47950,N_45040,N_45490);
nand U47951 (N_47951,N_45986,N_46100);
xnor U47952 (N_47952,N_47268,N_46132);
nor U47953 (N_47953,N_47418,N_46944);
nand U47954 (N_47954,N_45655,N_45940);
xor U47955 (N_47955,N_46162,N_45820);
or U47956 (N_47956,N_45411,N_45094);
or U47957 (N_47957,N_45782,N_46757);
and U47958 (N_47958,N_47479,N_46155);
and U47959 (N_47959,N_45069,N_45728);
and U47960 (N_47960,N_47160,N_45109);
nor U47961 (N_47961,N_45987,N_46667);
or U47962 (N_47962,N_45729,N_47415);
xor U47963 (N_47963,N_46816,N_45150);
xnor U47964 (N_47964,N_45163,N_46283);
or U47965 (N_47965,N_46293,N_45667);
nand U47966 (N_47966,N_47143,N_47263);
and U47967 (N_47967,N_45183,N_45259);
nor U47968 (N_47968,N_45152,N_47368);
xor U47969 (N_47969,N_45422,N_47123);
nor U47970 (N_47970,N_45311,N_45517);
nand U47971 (N_47971,N_46295,N_46950);
nand U47972 (N_47972,N_46591,N_46539);
nand U47973 (N_47973,N_46006,N_46203);
nor U47974 (N_47974,N_47147,N_46561);
nand U47975 (N_47975,N_47338,N_46149);
or U47976 (N_47976,N_45835,N_46458);
nand U47977 (N_47977,N_46420,N_45242);
and U47978 (N_47978,N_45058,N_46075);
or U47979 (N_47979,N_46628,N_45555);
or U47980 (N_47980,N_46253,N_45734);
and U47981 (N_47981,N_45106,N_46577);
and U47982 (N_47982,N_46166,N_47265);
nor U47983 (N_47983,N_45915,N_46626);
and U47984 (N_47984,N_46114,N_46967);
nor U47985 (N_47985,N_45777,N_46342);
nand U47986 (N_47986,N_47257,N_47020);
or U47987 (N_47987,N_47334,N_46300);
nor U47988 (N_47988,N_46614,N_47499);
nor U47989 (N_47989,N_45858,N_46516);
nor U47990 (N_47990,N_46439,N_45272);
nand U47991 (N_47991,N_45062,N_47209);
xnor U47992 (N_47992,N_45127,N_45114);
nor U47993 (N_47993,N_47284,N_46815);
xnor U47994 (N_47994,N_45350,N_45657);
nand U47995 (N_47995,N_46537,N_45229);
nor U47996 (N_47996,N_46610,N_46418);
and U47997 (N_47997,N_46983,N_45741);
and U47998 (N_47998,N_45865,N_45320);
or U47999 (N_47999,N_46115,N_47157);
nand U48000 (N_48000,N_45301,N_47300);
or U48001 (N_48001,N_45457,N_45567);
nor U48002 (N_48002,N_46842,N_46453);
nand U48003 (N_48003,N_46848,N_45514);
xnor U48004 (N_48004,N_47246,N_46475);
and U48005 (N_48005,N_46371,N_46909);
and U48006 (N_48006,N_46394,N_46424);
xnor U48007 (N_48007,N_45628,N_46247);
nand U48008 (N_48008,N_45964,N_45607);
nor U48009 (N_48009,N_47315,N_45995);
xnor U48010 (N_48010,N_45961,N_45448);
xor U48011 (N_48011,N_45285,N_45195);
nor U48012 (N_48012,N_47030,N_45499);
nand U48013 (N_48013,N_46780,N_45764);
and U48014 (N_48014,N_45483,N_46422);
nor U48015 (N_48015,N_46812,N_46941);
nor U48016 (N_48016,N_46121,N_47358);
nand U48017 (N_48017,N_45965,N_47039);
and U48018 (N_48018,N_47106,N_45226);
nor U48019 (N_48019,N_46988,N_46270);
nor U48020 (N_48020,N_46178,N_46897);
nand U48021 (N_48021,N_46022,N_45855);
xnor U48022 (N_48022,N_46384,N_45571);
xnor U48023 (N_48023,N_46849,N_45370);
nor U48024 (N_48024,N_46336,N_45904);
nor U48025 (N_48025,N_46414,N_47476);
or U48026 (N_48026,N_46719,N_45296);
or U48027 (N_48027,N_45428,N_45080);
or U48028 (N_48028,N_46581,N_46995);
xor U48029 (N_48029,N_45175,N_45643);
and U48030 (N_48030,N_46113,N_45772);
nor U48031 (N_48031,N_46592,N_47050);
nor U48032 (N_48032,N_47009,N_46054);
xnor U48033 (N_48033,N_45189,N_45629);
xor U48034 (N_48034,N_45693,N_46124);
nor U48035 (N_48035,N_47091,N_45580);
xor U48036 (N_48036,N_45552,N_46182);
or U48037 (N_48037,N_46048,N_46087);
nor U48038 (N_48038,N_45481,N_46625);
and U48039 (N_48039,N_47061,N_46521);
xnor U48040 (N_48040,N_45834,N_46096);
and U48041 (N_48041,N_46519,N_45746);
or U48042 (N_48042,N_45374,N_46376);
nor U48043 (N_48043,N_47226,N_46776);
xnor U48044 (N_48044,N_45444,N_46347);
xor U48045 (N_48045,N_47232,N_45828);
nor U48046 (N_48046,N_45710,N_45649);
nand U48047 (N_48047,N_46517,N_45512);
xnor U48048 (N_48048,N_46192,N_45513);
xnor U48049 (N_48049,N_46953,N_46603);
or U48050 (N_48050,N_45237,N_47173);
xnor U48051 (N_48051,N_46152,N_45557);
and U48052 (N_48052,N_45705,N_45745);
and U48053 (N_48053,N_46362,N_46221);
nand U48054 (N_48054,N_45909,N_45284);
or U48055 (N_48055,N_46570,N_45804);
nand U48056 (N_48056,N_47345,N_45780);
nand U48057 (N_48057,N_45362,N_45377);
or U48058 (N_48058,N_45220,N_46268);
or U48059 (N_48059,N_47365,N_46856);
or U48060 (N_48060,N_45519,N_45417);
nor U48061 (N_48061,N_45487,N_47375);
nor U48062 (N_48062,N_46693,N_46032);
nor U48063 (N_48063,N_46183,N_45930);
or U48064 (N_48064,N_45524,N_45232);
or U48065 (N_48065,N_45785,N_46164);
xnor U48066 (N_48066,N_45125,N_46504);
nand U48067 (N_48067,N_47305,N_46890);
and U48068 (N_48068,N_45450,N_45360);
nor U48069 (N_48069,N_47491,N_46854);
xnor U48070 (N_48070,N_45703,N_45408);
and U48071 (N_48071,N_47277,N_47142);
or U48072 (N_48072,N_45678,N_45140);
nand U48073 (N_48073,N_47402,N_45269);
or U48074 (N_48074,N_47255,N_45997);
xnor U48075 (N_48075,N_45719,N_45476);
xor U48076 (N_48076,N_46274,N_46704);
nor U48077 (N_48077,N_45166,N_45672);
nand U48078 (N_48078,N_45581,N_47184);
nor U48079 (N_48079,N_45549,N_47448);
nand U48080 (N_48080,N_46296,N_46142);
nand U48081 (N_48081,N_45526,N_46855);
nor U48082 (N_48082,N_47291,N_46455);
and U48083 (N_48083,N_45482,N_46968);
and U48084 (N_48084,N_47299,N_46224);
or U48085 (N_48085,N_46303,N_46464);
or U48086 (N_48086,N_46659,N_46830);
or U48087 (N_48087,N_45141,N_45162);
or U48088 (N_48088,N_45913,N_47399);
xnor U48089 (N_48089,N_47386,N_46220);
or U48090 (N_48090,N_45645,N_46615);
or U48091 (N_48091,N_46060,N_46718);
nor U48092 (N_48092,N_46156,N_46419);
nor U48093 (N_48093,N_47331,N_47450);
nor U48094 (N_48094,N_46884,N_45117);
and U48095 (N_48095,N_47016,N_46120);
and U48096 (N_48096,N_46010,N_47347);
or U48097 (N_48097,N_45509,N_45591);
or U48098 (N_48098,N_46364,N_46544);
xnor U48099 (N_48099,N_45205,N_45910);
nor U48100 (N_48100,N_45354,N_46506);
and U48101 (N_48101,N_45049,N_46905);
or U48102 (N_48102,N_47494,N_45878);
and U48103 (N_48103,N_45413,N_46518);
nand U48104 (N_48104,N_46188,N_46998);
nor U48105 (N_48105,N_46552,N_46285);
nor U48106 (N_48106,N_46616,N_45621);
nor U48107 (N_48107,N_45770,N_45955);
nor U48108 (N_48108,N_46180,N_46940);
and U48109 (N_48109,N_46559,N_47089);
or U48110 (N_48110,N_45663,N_47306);
or U48111 (N_48111,N_45445,N_46346);
and U48112 (N_48112,N_45148,N_45123);
nand U48113 (N_48113,N_45274,N_45698);
or U48114 (N_48114,N_46216,N_46059);
xor U48115 (N_48115,N_46402,N_46644);
xnor U48116 (N_48116,N_45472,N_45170);
xor U48117 (N_48117,N_46587,N_45850);
xnor U48118 (N_48118,N_45808,N_46942);
nor U48119 (N_48119,N_46817,N_46731);
or U48120 (N_48120,N_46211,N_45463);
or U48121 (N_48121,N_45251,N_45497);
xor U48122 (N_48122,N_45045,N_46447);
or U48123 (N_48123,N_45786,N_46823);
and U48124 (N_48124,N_45993,N_45502);
and U48125 (N_48125,N_45419,N_46329);
nor U48126 (N_48126,N_46650,N_47054);
and U48127 (N_48127,N_45893,N_46595);
and U48128 (N_48128,N_45014,N_45817);
nand U48129 (N_48129,N_46568,N_46343);
nand U48130 (N_48130,N_45577,N_45903);
nand U48131 (N_48131,N_46705,N_45480);
nand U48132 (N_48132,N_45397,N_45635);
xor U48133 (N_48133,N_46547,N_47071);
nand U48134 (N_48134,N_46990,N_47256);
or U48135 (N_48135,N_45556,N_46987);
and U48136 (N_48136,N_45489,N_45829);
and U48137 (N_48137,N_46202,N_45266);
and U48138 (N_48138,N_47460,N_46527);
or U48139 (N_48139,N_45488,N_45319);
xor U48140 (N_48140,N_46717,N_47335);
xor U48141 (N_48141,N_46169,N_46778);
or U48142 (N_48142,N_45254,N_46820);
xor U48143 (N_48143,N_46277,N_45956);
xnor U48144 (N_48144,N_46608,N_45980);
or U48145 (N_48145,N_45516,N_45133);
and U48146 (N_48146,N_47033,N_45842);
nand U48147 (N_48147,N_45302,N_45781);
or U48148 (N_48148,N_47070,N_46543);
or U48149 (N_48149,N_46769,N_46673);
nor U48150 (N_48150,N_46259,N_46576);
nor U48151 (N_48151,N_47204,N_45877);
nand U48152 (N_48152,N_45034,N_47328);
or U48153 (N_48153,N_45544,N_46238);
xnor U48154 (N_48154,N_47302,N_46242);
or U48155 (N_48155,N_45400,N_46209);
nor U48156 (N_48156,N_45090,N_45885);
nor U48157 (N_48157,N_46490,N_47245);
xnor U48158 (N_48158,N_47005,N_47223);
nand U48159 (N_48159,N_45381,N_45833);
nand U48160 (N_48160,N_47052,N_46013);
nor U48161 (N_48161,N_45686,N_46701);
or U48162 (N_48162,N_46141,N_46106);
nand U48163 (N_48163,N_46921,N_45073);
and U48164 (N_48164,N_46425,N_46874);
and U48165 (N_48165,N_45646,N_47457);
nor U48166 (N_48166,N_46104,N_45305);
nand U48167 (N_48167,N_45876,N_46427);
nand U48168 (N_48168,N_46143,N_45946);
or U48169 (N_48169,N_45530,N_46513);
or U48170 (N_48170,N_47107,N_46779);
xnor U48171 (N_48171,N_45868,N_47028);
nor U48172 (N_48172,N_46961,N_45196);
nor U48173 (N_48173,N_46715,N_47428);
nor U48174 (N_48174,N_45822,N_47231);
nand U48175 (N_48175,N_47376,N_45641);
nor U48176 (N_48176,N_46843,N_46933);
xnor U48177 (N_48177,N_45531,N_46922);
and U48178 (N_48178,N_45113,N_47438);
xor U48179 (N_48179,N_47219,N_45160);
nand U48180 (N_48180,N_46564,N_46399);
nand U48181 (N_48181,N_46436,N_47311);
xnor U48182 (N_48182,N_46172,N_45297);
or U48183 (N_48183,N_46753,N_45945);
and U48184 (N_48184,N_46575,N_45916);
xnor U48185 (N_48185,N_46080,N_46440);
or U48186 (N_48186,N_46687,N_46474);
and U48187 (N_48187,N_45688,N_45173);
xor U48188 (N_48188,N_47004,N_47455);
nand U48189 (N_48189,N_45147,N_47410);
and U48190 (N_48190,N_46741,N_47150);
xnor U48191 (N_48191,N_45814,N_45848);
nor U48192 (N_48192,N_45315,N_47458);
and U48193 (N_48193,N_47121,N_47242);
or U48194 (N_48194,N_47435,N_45334);
or U48195 (N_48195,N_45973,N_47215);
and U48196 (N_48196,N_46525,N_46510);
nand U48197 (N_48197,N_45926,N_46911);
xor U48198 (N_48198,N_45748,N_45473);
nand U48199 (N_48199,N_47046,N_47405);
xnor U48200 (N_48200,N_45464,N_46105);
nor U48201 (N_48201,N_45799,N_46317);
or U48202 (N_48202,N_46385,N_47244);
or U48203 (N_48203,N_46526,N_46252);
nor U48204 (N_48204,N_45078,N_47393);
nand U48205 (N_48205,N_45931,N_46859);
nor U48206 (N_48206,N_46720,N_47383);
xor U48207 (N_48207,N_46496,N_46985);
nor U48208 (N_48208,N_45230,N_46563);
and U48209 (N_48209,N_46363,N_45522);
xnor U48210 (N_48210,N_47385,N_45068);
and U48211 (N_48211,N_46930,N_47098);
and U48212 (N_48212,N_47200,N_46134);
xnor U48213 (N_48213,N_45839,N_47099);
xnor U48214 (N_48214,N_45844,N_45763);
and U48215 (N_48215,N_45081,N_46067);
xnor U48216 (N_48216,N_47093,N_47066);
and U48217 (N_48217,N_47464,N_45393);
nor U48218 (N_48218,N_46031,N_46026);
xor U48219 (N_48219,N_46401,N_47161);
and U48220 (N_48220,N_47459,N_45749);
or U48221 (N_48221,N_46052,N_47140);
nor U48222 (N_48222,N_45250,N_45447);
xor U48223 (N_48223,N_45142,N_47213);
nand U48224 (N_48224,N_46212,N_45932);
nand U48225 (N_48225,N_46408,N_45988);
nand U48226 (N_48226,N_46831,N_45506);
or U48227 (N_48227,N_45966,N_46217);
nor U48228 (N_48228,N_46640,N_46123);
xor U48229 (N_48229,N_46698,N_46073);
nor U48230 (N_48230,N_45827,N_46725);
nand U48231 (N_48231,N_47286,N_46694);
and U48232 (N_48232,N_46935,N_47330);
or U48233 (N_48233,N_46282,N_46807);
nand U48234 (N_48234,N_47130,N_45790);
nor U48235 (N_48235,N_46502,N_45565);
or U48236 (N_48236,N_46264,N_47163);
nor U48237 (N_48237,N_45707,N_45840);
xnor U48238 (N_48238,N_47198,N_46500);
xnor U48239 (N_48239,N_47001,N_45389);
nand U48240 (N_48240,N_46260,N_46369);
xor U48241 (N_48241,N_47495,N_45650);
nor U48242 (N_48242,N_47227,N_45415);
nand U48243 (N_48243,N_46161,N_45894);
nand U48244 (N_48244,N_45722,N_46699);
nand U48245 (N_48245,N_47276,N_46049);
or U48246 (N_48246,N_46405,N_45616);
nand U48247 (N_48247,N_46454,N_45138);
xor U48248 (N_48248,N_47281,N_45365);
and U48249 (N_48249,N_45172,N_46899);
nor U48250 (N_48250,N_47322,N_45947);
and U48251 (N_48251,N_45994,N_46170);
or U48252 (N_48252,N_46276,N_45740);
nand U48253 (N_48253,N_45852,N_46689);
xor U48254 (N_48254,N_46594,N_47487);
nor U48255 (N_48255,N_45792,N_45665);
nand U48256 (N_48256,N_46926,N_46566);
or U48257 (N_48257,N_47094,N_47492);
nor U48258 (N_48258,N_45326,N_46580);
and U48259 (N_48259,N_46618,N_45936);
and U48260 (N_48260,N_45246,N_45021);
nor U48261 (N_48261,N_45214,N_47169);
nor U48262 (N_48262,N_46964,N_45359);
xor U48263 (N_48263,N_47144,N_45206);
nand U48264 (N_48264,N_45501,N_45906);
or U48265 (N_48265,N_46861,N_46889);
nand U48266 (N_48266,N_47151,N_46612);
nor U48267 (N_48267,N_45048,N_45924);
and U48268 (N_48268,N_45849,N_46916);
and U48269 (N_48269,N_45425,N_46084);
and U48270 (N_48270,N_47417,N_45815);
nor U48271 (N_48271,N_47485,N_47086);
nor U48272 (N_48272,N_45831,N_46337);
and U48273 (N_48273,N_46103,N_46954);
or U48274 (N_48274,N_46931,N_46230);
xor U48275 (N_48275,N_45783,N_47230);
or U48276 (N_48276,N_46875,N_45426);
xnor U48277 (N_48277,N_45439,N_46700);
nor U48278 (N_48278,N_46800,N_46085);
xnor U48279 (N_48279,N_45258,N_45367);
nand U48280 (N_48280,N_46840,N_45944);
or U48281 (N_48281,N_46198,N_46668);
nor U48282 (N_48282,N_46802,N_46751);
nand U48283 (N_48283,N_46681,N_46278);
or U48284 (N_48284,N_45601,N_46327);
or U48285 (N_48285,N_47411,N_46879);
nand U48286 (N_48286,N_45291,N_47272);
nor U48287 (N_48287,N_46118,N_45742);
nand U48288 (N_48288,N_45005,N_45124);
or U48289 (N_48289,N_45057,N_45750);
nand U48290 (N_48290,N_46986,N_46395);
or U48291 (N_48291,N_45875,N_46404);
nand U48292 (N_48292,N_46597,N_46600);
nor U48293 (N_48293,N_45696,N_46908);
or U48294 (N_48294,N_46894,N_46286);
and U48295 (N_48295,N_45529,N_45353);
nor U48296 (N_48296,N_45126,N_46904);
or U48297 (N_48297,N_47318,N_45380);
or U48298 (N_48298,N_47456,N_47103);
or U48299 (N_48299,N_45403,N_46284);
nand U48300 (N_48300,N_47384,N_45023);
nor U48301 (N_48301,N_45179,N_46435);
nor U48302 (N_48302,N_47356,N_47205);
or U48303 (N_48303,N_45271,N_45539);
or U48304 (N_48304,N_46255,N_46299);
nand U48305 (N_48305,N_45902,N_45156);
nand U48306 (N_48306,N_46258,N_45054);
nand U48307 (N_48307,N_46937,N_46572);
or U48308 (N_48308,N_47324,N_45889);
nor U48309 (N_48309,N_45468,N_45115);
or U48310 (N_48310,N_47069,N_46999);
and U48311 (N_48311,N_47259,N_45570);
and U48312 (N_48312,N_45077,N_46789);
xnor U48313 (N_48313,N_46688,N_46195);
or U48314 (N_48314,N_45281,N_45193);
nand U48315 (N_48315,N_45543,N_45596);
nand U48316 (N_48316,N_47079,N_45098);
xnor U48317 (N_48317,N_46236,N_45387);
or U48318 (N_48318,N_46637,N_45685);
and U48319 (N_48319,N_45507,N_45919);
or U48320 (N_48320,N_45299,N_46927);
xnor U48321 (N_48321,N_45000,N_46529);
or U48322 (N_48322,N_46486,N_46023);
nand U48323 (N_48323,N_47249,N_45671);
and U48324 (N_48324,N_46606,N_46873);
nand U48325 (N_48325,N_45067,N_46865);
nor U48326 (N_48326,N_45238,N_46760);
xnor U48327 (N_48327,N_45866,N_46691);
or U48328 (N_48328,N_47136,N_45992);
nand U48329 (N_48329,N_46989,N_45807);
nor U48330 (N_48330,N_46512,N_45689);
nor U48331 (N_48331,N_46852,N_46321);
xor U48332 (N_48332,N_46746,N_47360);
or U48333 (N_48333,N_45392,N_46796);
and U48334 (N_48334,N_46790,N_46949);
xnor U48335 (N_48335,N_47119,N_46098);
or U48336 (N_48336,N_45300,N_46215);
nor U48337 (N_48337,N_46878,N_45805);
nand U48338 (N_48338,N_46522,N_45104);
xnor U48339 (N_48339,N_46918,N_46016);
xnor U48340 (N_48340,N_46116,N_47289);
nand U48341 (N_48341,N_45017,N_45327);
nand U48342 (N_48342,N_46806,N_45340);
and U48343 (N_48343,N_46261,N_47165);
and U48344 (N_48344,N_46887,N_45418);
nand U48345 (N_48345,N_46273,N_45221);
or U48346 (N_48346,N_45897,N_45503);
and U48347 (N_48347,N_46795,N_46794);
and U48348 (N_48348,N_46396,N_47041);
xor U48349 (N_48349,N_47167,N_47382);
or U48350 (N_48350,N_45604,N_45587);
nand U48351 (N_48351,N_46819,N_46994);
nor U48352 (N_48352,N_47425,N_45737);
or U48353 (N_48353,N_45051,N_47105);
nor U48354 (N_48354,N_46952,N_47308);
xor U48355 (N_48355,N_46652,N_46348);
and U48356 (N_48356,N_45317,N_45843);
and U48357 (N_48357,N_46696,N_46322);
nor U48358 (N_48358,N_46122,N_45042);
nand U48359 (N_48359,N_45541,N_47166);
xor U48360 (N_48360,N_47096,N_46119);
nor U48361 (N_48361,N_46310,N_45573);
nor U48362 (N_48362,N_45551,N_45174);
and U48363 (N_48363,N_45532,N_46305);
or U48364 (N_48364,N_45105,N_45681);
and U48365 (N_48365,N_45225,N_45407);
xnor U48366 (N_48366,N_45730,N_45515);
and U48367 (N_48367,N_45429,N_47170);
nor U48368 (N_48368,N_46984,N_45564);
xnor U48369 (N_48369,N_46774,N_46702);
nand U48370 (N_48370,N_46907,N_45736);
nand U48371 (N_48371,N_46050,N_46058);
nand U48372 (N_48372,N_46129,N_45267);
nand U48373 (N_48373,N_45191,N_46870);
and U48374 (N_48374,N_46832,N_47471);
or U48375 (N_48375,N_46613,N_45007);
nand U48376 (N_48376,N_45075,N_45953);
xnor U48377 (N_48377,N_46841,N_46530);
nand U48378 (N_48378,N_47199,N_45288);
and U48379 (N_48379,N_46759,N_46176);
and U48380 (N_48380,N_46478,N_45811);
or U48381 (N_48381,N_46102,N_47396);
and U48382 (N_48382,N_45674,N_45149);
nand U48383 (N_48383,N_46313,N_46108);
nor U48384 (N_48384,N_45614,N_45186);
xor U48385 (N_48385,N_46913,N_46747);
nor U48386 (N_48386,N_47177,N_45231);
xnor U48387 (N_48387,N_45357,N_45029);
and U48388 (N_48388,N_46263,N_45658);
or U48389 (N_48389,N_45599,N_46571);
xnor U48390 (N_48390,N_46377,N_46733);
xor U48391 (N_48391,N_46449,N_46866);
xnor U48392 (N_48392,N_45970,N_45460);
nor U48393 (N_48393,N_45523,N_47401);
and U48394 (N_48394,N_46097,N_47221);
or U48395 (N_48395,N_47496,N_46020);
and U48396 (N_48396,N_45533,N_47186);
xor U48397 (N_48397,N_46551,N_45268);
nand U48398 (N_48398,N_45026,N_46479);
or U48399 (N_48399,N_46635,N_45670);
xnor U48400 (N_48400,N_45933,N_46684);
nor U48401 (N_48401,N_45706,N_45182);
nand U48402 (N_48402,N_46131,N_46039);
nand U48403 (N_48403,N_47313,N_45310);
or U48404 (N_48404,N_47392,N_46822);
nor U48405 (N_48405,N_45768,N_47064);
or U48406 (N_48406,N_45378,N_45395);
or U48407 (N_48407,N_45396,N_47192);
xnor U48408 (N_48408,N_46160,N_46556);
or U48409 (N_48409,N_45466,N_46340);
and U48410 (N_48410,N_46298,N_45914);
nand U48411 (N_48411,N_47247,N_45603);
or U48412 (N_48412,N_45491,N_46786);
or U48413 (N_48413,N_45433,N_47395);
or U48414 (N_48414,N_45046,N_47497);
and U48415 (N_48415,N_46979,N_45286);
xor U48416 (N_48416,N_45854,N_47389);
xnor U48417 (N_48417,N_45331,N_47194);
or U48418 (N_48418,N_46378,N_46837);
xor U48419 (N_48419,N_45118,N_46677);
nand U48420 (N_48420,N_45954,N_45800);
and U48421 (N_48421,N_45680,N_46783);
and U48422 (N_48422,N_46094,N_45177);
nand U48423 (N_48423,N_46456,N_47482);
nor U48424 (N_48424,N_45582,N_46892);
nand U48425 (N_48425,N_45436,N_47180);
xnor U48426 (N_48426,N_46107,N_46827);
nand U48427 (N_48427,N_46112,N_47010);
or U48428 (N_48428,N_45321,N_46540);
xnor U48429 (N_48429,N_46872,N_45424);
nand U48430 (N_48430,N_46069,N_46072);
nor U48431 (N_48431,N_47254,N_46939);
xnor U48432 (N_48432,N_47465,N_47432);
xnor U48433 (N_48433,N_45934,N_46074);
xor U48434 (N_48434,N_47436,N_46829);
nand U48435 (N_48435,N_45449,N_45702);
nor U48436 (N_48436,N_46542,N_46191);
nor U48437 (N_48437,N_46469,N_47412);
nand U48438 (N_48438,N_47040,N_46030);
or U48439 (N_48439,N_45518,N_46963);
nor U48440 (N_48440,N_45733,N_45579);
nand U48441 (N_48441,N_46461,N_46548);
and U48442 (N_48442,N_45108,N_47122);
xnor U48443 (N_48443,N_45337,N_47397);
and U48444 (N_48444,N_46514,N_46250);
and U48445 (N_48445,N_46256,N_46446);
or U48446 (N_48446,N_45723,N_45948);
or U48447 (N_48447,N_47431,N_45276);
and U48448 (N_48448,N_45989,N_46695);
nor U48449 (N_48449,N_45478,N_45003);
or U48450 (N_48450,N_47480,N_45566);
and U48451 (N_48451,N_46311,N_46037);
nor U48452 (N_48452,N_46976,N_47363);
nor U48453 (N_48453,N_46423,N_47366);
or U48454 (N_48454,N_47042,N_46948);
nor U48455 (N_48455,N_45361,N_45438);
nor U48456 (N_48456,N_46728,N_47233);
or U48457 (N_48457,N_45103,N_46798);
nand U48458 (N_48458,N_45952,N_46895);
xnor U48459 (N_48459,N_46744,N_46858);
and U48460 (N_48460,N_45862,N_46128);
nor U48461 (N_48461,N_46205,N_46770);
and U48462 (N_48462,N_46448,N_45917);
nand U48463 (N_48463,N_45957,N_47452);
nand U48464 (N_48464,N_45735,N_46487);
nor U48465 (N_48465,N_47461,N_45590);
nor U48466 (N_48466,N_46154,N_45203);
or U48467 (N_48467,N_46081,N_47006);
xnor U48468 (N_48468,N_46064,N_46692);
or U48469 (N_48469,N_45308,N_46683);
nor U48470 (N_48470,N_47196,N_47044);
nor U48471 (N_48471,N_47207,N_46934);
and U48472 (N_48472,N_45888,N_45708);
nand U48473 (N_48473,N_45290,N_47261);
xnor U48474 (N_48474,N_45554,N_47146);
xor U48475 (N_48475,N_45059,N_45143);
xor U48476 (N_48476,N_46281,N_46945);
nand U48477 (N_48477,N_45493,N_46972);
nand U48478 (N_48478,N_47271,N_45520);
nor U48479 (N_48479,N_45056,N_45063);
and U48480 (N_48480,N_47278,N_47217);
and U48481 (N_48481,N_47430,N_45896);
or U48482 (N_48482,N_45761,N_46297);
xnor U48483 (N_48483,N_47187,N_45731);
xor U48484 (N_48484,N_47463,N_47195);
and U48485 (N_48485,N_47349,N_45372);
xnor U48486 (N_48486,N_46167,N_45534);
nor U48487 (N_48487,N_45979,N_46248);
nor U48488 (N_48488,N_46139,N_45756);
xor U48489 (N_48489,N_47083,N_45158);
and U48490 (N_48490,N_45471,N_47462);
or U48491 (N_48491,N_45313,N_46917);
or U48492 (N_48492,N_45181,N_47032);
nor U48493 (N_48493,N_45738,N_45038);
nand U48494 (N_48494,N_46386,N_46903);
nor U48495 (N_48495,N_45477,N_45958);
or U48496 (N_48496,N_45006,N_46690);
or U48497 (N_48497,N_45211,N_45984);
or U48498 (N_48498,N_46734,N_46623);
or U48499 (N_48499,N_46946,N_46213);
nand U48500 (N_48500,N_47439,N_45201);
nand U48501 (N_48501,N_46598,N_46159);
xor U48502 (N_48502,N_47181,N_45352);
nor U48503 (N_48503,N_46970,N_45575);
nand U48504 (N_48504,N_46043,N_46498);
nand U48505 (N_48505,N_46262,N_46914);
xnor U48506 (N_48506,N_45128,N_47359);
and U48507 (N_48507,N_45508,N_47003);
nor U48508 (N_48508,N_46314,N_45240);
nand U48509 (N_48509,N_46165,N_46721);
nor U48510 (N_48510,N_47478,N_45461);
nand U48511 (N_48511,N_46288,N_47080);
nand U48512 (N_48512,N_47197,N_45329);
or U48513 (N_48513,N_45120,N_45265);
or U48514 (N_48514,N_46869,N_47236);
xnor U48515 (N_48515,N_46381,N_47202);
nand U48516 (N_48516,N_46974,N_45907);
or U48517 (N_48517,N_47426,N_45180);
or U48518 (N_48518,N_47002,N_47442);
or U48519 (N_48519,N_47468,N_47022);
or U48520 (N_48520,N_47374,N_46061);
or U48521 (N_48521,N_45500,N_45171);
xnor U48522 (N_48522,N_45634,N_47239);
nand U48523 (N_48523,N_46055,N_45280);
and U48524 (N_48524,N_45458,N_46289);
or U48525 (N_48525,N_45592,N_46033);
or U48526 (N_48526,N_45333,N_46962);
or U48527 (N_48527,N_45578,N_46471);
or U48528 (N_48528,N_45712,N_45107);
nand U48529 (N_48529,N_45971,N_46034);
nor U48530 (N_48530,N_47102,N_46430);
or U48531 (N_48531,N_46773,N_47352);
nand U48532 (N_48532,N_45210,N_46641);
or U48533 (N_48533,N_45052,N_45525);
xor U48534 (N_48534,N_45134,N_45079);
or U48535 (N_48535,N_46339,N_45869);
nand U48536 (N_48536,N_47021,N_46389);
nor U48537 (N_48537,N_46676,N_47135);
and U48538 (N_48538,N_46726,N_47190);
nor U48539 (N_48539,N_46056,N_47036);
nand U48540 (N_48540,N_45346,N_46605);
nand U48541 (N_48541,N_47451,N_47141);
nor U48542 (N_48542,N_46392,N_45228);
or U48543 (N_48543,N_46622,N_46350);
nand U48544 (N_48544,N_46557,N_46467);
xnor U48545 (N_48545,N_47252,N_45253);
nor U48546 (N_48546,N_46326,N_45204);
and U48547 (N_48547,N_46481,N_45050);
or U48548 (N_48548,N_47414,N_47055);
nand U48549 (N_48549,N_47400,N_45145);
xnor U48550 (N_48550,N_45188,N_46749);
xnor U48551 (N_48551,N_45453,N_45682);
and U48552 (N_48552,N_46349,N_46523);
nand U48553 (N_48553,N_46868,N_45283);
or U48554 (N_48554,N_47248,N_45129);
and U48555 (N_48555,N_47051,N_46076);
nand U48556 (N_48556,N_46421,N_46617);
and U48557 (N_48557,N_46943,N_46135);
or U48558 (N_48558,N_47019,N_45347);
nand U48559 (N_48559,N_46712,N_47440);
xor U48560 (N_48560,N_46352,N_46853);
or U48561 (N_48561,N_47133,N_46189);
nor U48562 (N_48562,N_45345,N_46520);
nand U48563 (N_48563,N_45960,N_46881);
nor U48564 (N_48564,N_45535,N_45857);
or U48565 (N_48565,N_46993,N_47447);
and U48566 (N_48566,N_45620,N_45030);
and U48567 (N_48567,N_46768,N_45921);
and U48568 (N_48568,N_46457,N_47469);
or U48569 (N_48569,N_45861,N_45821);
nand U48570 (N_48570,N_46891,N_47420);
and U48571 (N_48571,N_46485,N_45864);
xor U48572 (N_48572,N_45881,N_47337);
xnor U48573 (N_48573,N_47433,N_46579);
and U48574 (N_48574,N_46227,N_45169);
or U48575 (N_48575,N_45343,N_45083);
or U48576 (N_48576,N_47024,N_45309);
nor U48577 (N_48577,N_47025,N_45568);
nor U48578 (N_48578,N_47059,N_47312);
nor U48579 (N_48579,N_45486,N_47441);
or U48580 (N_48580,N_47134,N_47253);
nor U48581 (N_48581,N_45538,N_46602);
xor U48582 (N_48582,N_45836,N_46977);
nand U48583 (N_48583,N_46896,N_46740);
nor U48584 (N_48584,N_45187,N_45279);
and U48585 (N_48585,N_46400,N_46232);
and U48586 (N_48586,N_45009,N_46472);
nand U48587 (N_48587,N_47189,N_47403);
or U48588 (N_48588,N_47466,N_46706);
xor U48589 (N_48589,N_45856,N_47077);
xor U48590 (N_48590,N_45420,N_45492);
xor U48591 (N_48591,N_45130,N_45386);
or U48592 (N_48592,N_46958,N_46507);
or U48593 (N_48593,N_46045,N_45137);
xnor U48594 (N_48594,N_47014,N_47367);
or U48595 (N_48595,N_47110,N_46686);
nor U48596 (N_48596,N_46335,N_46426);
or U48597 (N_48597,N_45462,N_45872);
or U48598 (N_48598,N_46589,N_46515);
nor U48599 (N_48599,N_45905,N_45684);
nor U48600 (N_48600,N_45452,N_46307);
and U48601 (N_48601,N_45199,N_46254);
and U48602 (N_48602,N_46754,N_45589);
and U48603 (N_48603,N_47280,N_46584);
and U48604 (N_48604,N_45235,N_45851);
nor U48605 (N_48605,N_47419,N_47101);
xnor U48606 (N_48606,N_45282,N_46996);
and U48607 (N_48607,N_47129,N_47258);
nand U48608 (N_48608,N_45798,N_45010);
nand U48609 (N_48609,N_46824,N_47193);
and U48610 (N_48610,N_46358,N_45713);
and U48611 (N_48611,N_45791,N_46821);
or U48612 (N_48612,N_46818,N_47208);
xor U48613 (N_48613,N_47290,N_45873);
and U48614 (N_48614,N_46923,N_45615);
or U48615 (N_48615,N_46365,N_45342);
or U48616 (N_48616,N_45263,N_46047);
or U48617 (N_48617,N_45846,N_46078);
and U48618 (N_48618,N_45975,N_45795);
and U48619 (N_48619,N_47203,N_47339);
xor U48620 (N_48620,N_46664,N_45248);
nand U48621 (N_48621,N_47292,N_45132);
xnor U48622 (N_48622,N_45312,N_45727);
xnor U48623 (N_48623,N_46197,N_47288);
nor U48624 (N_48624,N_46000,N_46596);
nand U48625 (N_48625,N_46727,N_45847);
nor U48626 (N_48626,N_47353,N_47336);
xnor U48627 (N_48627,N_46315,N_46912);
and U48628 (N_48628,N_45084,N_47317);
xnor U48629 (N_48629,N_46126,N_46002);
xor U48630 (N_48630,N_47309,N_46813);
or U48631 (N_48631,N_47027,N_46647);
nor U48632 (N_48632,N_46505,N_45085);
or U48633 (N_48633,N_45882,N_46730);
and U48634 (N_48634,N_47063,N_46437);
and U48635 (N_48635,N_46368,N_45025);
xor U48636 (N_48636,N_45485,N_45818);
nor U48637 (N_48637,N_46082,N_47053);
or U48638 (N_48638,N_46670,N_46434);
or U48639 (N_48639,N_46153,N_46836);
and U48640 (N_48640,N_46412,N_45867);
and U48641 (N_48641,N_47481,N_45588);
xnor U48642 (N_48642,N_45883,N_46136);
or U48643 (N_48643,N_45853,N_45778);
or U48644 (N_48644,N_46627,N_45619);
nor U48645 (N_48645,N_45213,N_47216);
and U48646 (N_48646,N_47296,N_45012);
nor U48647 (N_48647,N_46390,N_46241);
and U48648 (N_48648,N_46243,N_45440);
or U48649 (N_48649,N_45941,N_45278);
xnor U48650 (N_48650,N_47095,N_46787);
nand U48651 (N_48651,N_45793,N_47332);
nand U48652 (N_48652,N_47211,N_45474);
nor U48653 (N_48653,N_45459,N_46503);
or U48654 (N_48654,N_45594,N_46982);
xnor U48655 (N_48655,N_45642,N_45775);
nor U48656 (N_48656,N_45155,N_46190);
or U48657 (N_48657,N_47355,N_46619);
and U48658 (N_48658,N_45900,N_45289);
or U48659 (N_48659,N_47114,N_45008);
or U48660 (N_48660,N_47097,N_46372);
and U48661 (N_48661,N_46168,N_45022);
nand U48662 (N_48662,N_45066,N_47067);
nand U48663 (N_48663,N_47378,N_46008);
and U48664 (N_48664,N_45923,N_45925);
nand U48665 (N_48665,N_47470,N_46679);
nor U48666 (N_48666,N_46038,N_46301);
xnor U48667 (N_48667,N_45819,N_46863);
nand U48668 (N_48668,N_45679,N_46228);
nor U48669 (N_48669,N_45697,N_45794);
and U48670 (N_48670,N_45139,N_46565);
and U48671 (N_48671,N_47391,N_46476);
or U48672 (N_48672,N_47362,N_46251);
nand U48673 (N_48673,N_47013,N_45636);
or U48674 (N_48674,N_46460,N_45293);
xnor U48675 (N_48675,N_45631,N_45256);
nand U48676 (N_48676,N_45633,N_46981);
and U48677 (N_48677,N_46716,N_45990);
or U48678 (N_48678,N_46271,N_47018);
nand U48679 (N_48679,N_45207,N_45838);
or U48680 (N_48680,N_46657,N_46742);
or U48681 (N_48681,N_46433,N_46144);
xnor U48682 (N_48682,N_45879,N_47178);
nand U48683 (N_48683,N_45691,N_46862);
or U48684 (N_48684,N_46151,N_47152);
and U48685 (N_48685,N_46066,N_46672);
and U48686 (N_48686,N_47171,N_45563);
and U48687 (N_48687,N_46280,N_45434);
and U48688 (N_48688,N_45561,N_45752);
or U48689 (N_48689,N_45999,N_45178);
nor U48690 (N_48690,N_46737,N_47034);
or U48691 (N_48691,N_45779,N_47087);
xnor U48692 (N_48692,N_46834,N_45096);
xor U48693 (N_48693,N_47158,N_46137);
nor U48694 (N_48694,N_46772,N_46077);
nand U48695 (N_48695,N_45717,N_45198);
or U48696 (N_48696,N_47351,N_46091);
xor U48697 (N_48697,N_45884,N_46308);
nor U48698 (N_48698,N_45243,N_46906);
or U48699 (N_48699,N_45366,N_46919);
nand U48700 (N_48700,N_45135,N_45810);
or U48701 (N_48701,N_45219,N_47224);
and U48702 (N_48702,N_46145,N_46177);
xnor U48703 (N_48703,N_47449,N_45700);
nand U48704 (N_48704,N_46194,N_47437);
xnor U48705 (N_48705,N_45622,N_45404);
and U48706 (N_48706,N_45640,N_45318);
xnor U48707 (N_48707,N_45494,N_45521);
xor U48708 (N_48708,N_47320,N_45963);
nand U48709 (N_48709,N_46642,N_45825);
or U48710 (N_48710,N_46609,N_45802);
xnor U48711 (N_48711,N_46210,N_45659);
or U48712 (N_48712,N_45224,N_45774);
nor U48713 (N_48713,N_45348,N_45639);
and U48714 (N_48714,N_46839,N_47370);
nor U48715 (N_48715,N_46835,N_47172);
and U48716 (N_48716,N_47015,N_46001);
nand U48717 (N_48717,N_45704,N_45002);
xnor U48718 (N_48718,N_47266,N_47443);
and U48719 (N_48719,N_46240,N_46811);
and U48720 (N_48720,N_46531,N_47327);
xnor U48721 (N_48721,N_47076,N_46438);
nor U48722 (N_48722,N_45664,N_46697);
or U48723 (N_48723,N_45020,N_45239);
and U48724 (N_48724,N_46607,N_46332);
and U48725 (N_48725,N_45304,N_46775);
xnor U48726 (N_48726,N_46671,N_45322);
xor U48727 (N_48727,N_47319,N_46661);
nor U48728 (N_48728,N_45087,N_46257);
nor U48729 (N_48729,N_46204,N_45446);
and U48730 (N_48730,N_47220,N_46932);
nand U48731 (N_48731,N_45122,N_45574);
or U48732 (N_48732,N_46867,N_47429);
nor U48733 (N_48733,N_45033,N_45845);
nor U48734 (N_48734,N_47434,N_47000);
nand U48735 (N_48735,N_47238,N_46643);
nand U48736 (N_48736,N_46403,N_45651);
or U48737 (N_48737,N_46771,N_46450);
or U48738 (N_48738,N_46431,N_47149);
nor U48739 (N_48739,N_45653,N_47350);
xor U48740 (N_48740,N_45585,N_46291);
and U48741 (N_48741,N_45314,N_46955);
nor U48742 (N_48742,N_45097,N_47489);
xor U48743 (N_48743,N_46325,N_45586);
or U48744 (N_48744,N_46445,N_46226);
xnor U48745 (N_48745,N_47012,N_47074);
nor U48746 (N_48746,N_45262,N_46062);
nand U48747 (N_48747,N_45676,N_45011);
or U48748 (N_48748,N_46743,N_45711);
nand U48749 (N_48749,N_46755,N_46601);
or U48750 (N_48750,N_46669,N_46707);
or U48751 (N_48751,N_47207,N_45642);
or U48752 (N_48752,N_46236,N_45034);
nor U48753 (N_48753,N_46587,N_45256);
xnor U48754 (N_48754,N_45749,N_45641);
xnor U48755 (N_48755,N_47077,N_46238);
xor U48756 (N_48756,N_45165,N_45323);
xor U48757 (N_48757,N_46497,N_46320);
and U48758 (N_48758,N_46529,N_47173);
nand U48759 (N_48759,N_45195,N_46334);
xor U48760 (N_48760,N_47237,N_47399);
nand U48761 (N_48761,N_46380,N_46959);
xor U48762 (N_48762,N_46820,N_47327);
nand U48763 (N_48763,N_46551,N_45891);
or U48764 (N_48764,N_45033,N_45299);
and U48765 (N_48765,N_45037,N_47465);
or U48766 (N_48766,N_45547,N_45859);
xnor U48767 (N_48767,N_45853,N_46834);
xor U48768 (N_48768,N_45989,N_46012);
xor U48769 (N_48769,N_46191,N_45924);
and U48770 (N_48770,N_45967,N_47433);
xnor U48771 (N_48771,N_46932,N_46701);
and U48772 (N_48772,N_45497,N_45009);
xnor U48773 (N_48773,N_46181,N_45077);
nand U48774 (N_48774,N_46418,N_47296);
or U48775 (N_48775,N_45276,N_46304);
or U48776 (N_48776,N_47067,N_46480);
or U48777 (N_48777,N_46898,N_47170);
nor U48778 (N_48778,N_45925,N_46350);
xnor U48779 (N_48779,N_46590,N_45341);
nor U48780 (N_48780,N_45406,N_46387);
nor U48781 (N_48781,N_47166,N_46200);
and U48782 (N_48782,N_46144,N_45356);
xnor U48783 (N_48783,N_46449,N_45296);
nor U48784 (N_48784,N_45100,N_46183);
or U48785 (N_48785,N_45300,N_46885);
nand U48786 (N_48786,N_45201,N_47159);
xor U48787 (N_48787,N_45684,N_47147);
nand U48788 (N_48788,N_45707,N_47427);
nor U48789 (N_48789,N_45153,N_45653);
nand U48790 (N_48790,N_46525,N_46538);
or U48791 (N_48791,N_46522,N_46577);
nand U48792 (N_48792,N_45997,N_46388);
or U48793 (N_48793,N_45730,N_45202);
xnor U48794 (N_48794,N_46497,N_45747);
and U48795 (N_48795,N_47301,N_47427);
nand U48796 (N_48796,N_45668,N_47199);
or U48797 (N_48797,N_47439,N_47196);
or U48798 (N_48798,N_46870,N_46809);
xor U48799 (N_48799,N_46764,N_45008);
nand U48800 (N_48800,N_47287,N_46694);
or U48801 (N_48801,N_45171,N_45370);
nor U48802 (N_48802,N_46146,N_45549);
nor U48803 (N_48803,N_46428,N_46813);
xnor U48804 (N_48804,N_45041,N_45298);
and U48805 (N_48805,N_45393,N_45404);
and U48806 (N_48806,N_46799,N_46245);
nor U48807 (N_48807,N_45770,N_45915);
nand U48808 (N_48808,N_45833,N_45717);
xnor U48809 (N_48809,N_46918,N_45284);
and U48810 (N_48810,N_46672,N_45418);
nor U48811 (N_48811,N_47055,N_45808);
nand U48812 (N_48812,N_46630,N_47301);
or U48813 (N_48813,N_46622,N_46506);
nand U48814 (N_48814,N_45134,N_47217);
nand U48815 (N_48815,N_45328,N_45646);
xnor U48816 (N_48816,N_46799,N_46484);
nor U48817 (N_48817,N_45317,N_46610);
or U48818 (N_48818,N_46027,N_47381);
nand U48819 (N_48819,N_45777,N_45592);
and U48820 (N_48820,N_45587,N_46544);
or U48821 (N_48821,N_45225,N_46044);
nor U48822 (N_48822,N_46953,N_46156);
nor U48823 (N_48823,N_47274,N_45343);
nand U48824 (N_48824,N_46113,N_45792);
or U48825 (N_48825,N_46104,N_46520);
nor U48826 (N_48826,N_45610,N_45320);
nor U48827 (N_48827,N_46387,N_46673);
and U48828 (N_48828,N_47422,N_46168);
nand U48829 (N_48829,N_45729,N_46146);
or U48830 (N_48830,N_45115,N_47425);
nor U48831 (N_48831,N_46295,N_47460);
or U48832 (N_48832,N_47256,N_46861);
and U48833 (N_48833,N_47078,N_45765);
nand U48834 (N_48834,N_46052,N_46656);
and U48835 (N_48835,N_46465,N_45372);
or U48836 (N_48836,N_45971,N_46393);
nand U48837 (N_48837,N_45859,N_45652);
and U48838 (N_48838,N_46547,N_46745);
nor U48839 (N_48839,N_46068,N_45718);
xnor U48840 (N_48840,N_46156,N_46319);
nor U48841 (N_48841,N_46480,N_45111);
or U48842 (N_48842,N_45203,N_47265);
and U48843 (N_48843,N_45541,N_45889);
nand U48844 (N_48844,N_45978,N_45321);
nor U48845 (N_48845,N_45383,N_46942);
or U48846 (N_48846,N_46374,N_46673);
and U48847 (N_48847,N_45169,N_46457);
xnor U48848 (N_48848,N_45535,N_45931);
xnor U48849 (N_48849,N_45775,N_45207);
nand U48850 (N_48850,N_45819,N_45738);
and U48851 (N_48851,N_45237,N_45519);
xnor U48852 (N_48852,N_45197,N_46465);
nor U48853 (N_48853,N_45527,N_46553);
xor U48854 (N_48854,N_46649,N_47376);
nand U48855 (N_48855,N_45037,N_46086);
or U48856 (N_48856,N_45509,N_47480);
nor U48857 (N_48857,N_45073,N_45709);
nor U48858 (N_48858,N_46252,N_45092);
nand U48859 (N_48859,N_45876,N_45137);
nor U48860 (N_48860,N_46442,N_45625);
nor U48861 (N_48861,N_46303,N_46233);
or U48862 (N_48862,N_45933,N_47401);
or U48863 (N_48863,N_46512,N_46171);
nor U48864 (N_48864,N_46854,N_46196);
nand U48865 (N_48865,N_46694,N_46537);
xor U48866 (N_48866,N_46381,N_45973);
xnor U48867 (N_48867,N_46755,N_45550);
nand U48868 (N_48868,N_46848,N_45500);
nor U48869 (N_48869,N_46754,N_45557);
nor U48870 (N_48870,N_46765,N_46949);
xor U48871 (N_48871,N_46286,N_46608);
and U48872 (N_48872,N_46827,N_45658);
and U48873 (N_48873,N_45421,N_46023);
nand U48874 (N_48874,N_45320,N_47479);
xor U48875 (N_48875,N_47323,N_45562);
and U48876 (N_48876,N_45284,N_47431);
xnor U48877 (N_48877,N_45970,N_45477);
or U48878 (N_48878,N_46023,N_46964);
nand U48879 (N_48879,N_45122,N_46780);
xnor U48880 (N_48880,N_47031,N_45528);
xnor U48881 (N_48881,N_46003,N_45414);
nor U48882 (N_48882,N_46317,N_45950);
xnor U48883 (N_48883,N_47248,N_46058);
and U48884 (N_48884,N_47450,N_46982);
or U48885 (N_48885,N_47282,N_46169);
and U48886 (N_48886,N_46208,N_46260);
xor U48887 (N_48887,N_45579,N_46132);
nor U48888 (N_48888,N_45150,N_45540);
nor U48889 (N_48889,N_45609,N_46297);
or U48890 (N_48890,N_47321,N_46389);
xnor U48891 (N_48891,N_45744,N_46922);
nor U48892 (N_48892,N_45756,N_45344);
xor U48893 (N_48893,N_46373,N_46861);
or U48894 (N_48894,N_47337,N_47461);
and U48895 (N_48895,N_46686,N_46239);
and U48896 (N_48896,N_46949,N_46140);
nand U48897 (N_48897,N_47120,N_45240);
nand U48898 (N_48898,N_46270,N_46487);
nor U48899 (N_48899,N_46201,N_47039);
xor U48900 (N_48900,N_47004,N_46885);
and U48901 (N_48901,N_46257,N_45488);
and U48902 (N_48902,N_46818,N_45565);
and U48903 (N_48903,N_45270,N_47086);
and U48904 (N_48904,N_46475,N_46453);
and U48905 (N_48905,N_45228,N_46418);
and U48906 (N_48906,N_46158,N_46171);
or U48907 (N_48907,N_46218,N_46788);
nor U48908 (N_48908,N_47183,N_46904);
and U48909 (N_48909,N_45570,N_46673);
nor U48910 (N_48910,N_46957,N_45107);
and U48911 (N_48911,N_45250,N_46966);
xor U48912 (N_48912,N_45951,N_47349);
xnor U48913 (N_48913,N_46088,N_46488);
xnor U48914 (N_48914,N_47386,N_46477);
or U48915 (N_48915,N_47303,N_47240);
nand U48916 (N_48916,N_45620,N_47252);
nor U48917 (N_48917,N_45595,N_46266);
or U48918 (N_48918,N_46404,N_46762);
or U48919 (N_48919,N_46483,N_45088);
nor U48920 (N_48920,N_46390,N_46634);
nor U48921 (N_48921,N_45178,N_46684);
and U48922 (N_48922,N_47494,N_45879);
xnor U48923 (N_48923,N_45250,N_46206);
or U48924 (N_48924,N_45421,N_45832);
nand U48925 (N_48925,N_45020,N_45124);
or U48926 (N_48926,N_45247,N_46563);
nand U48927 (N_48927,N_46341,N_46149);
xnor U48928 (N_48928,N_47460,N_45739);
or U48929 (N_48929,N_46433,N_47016);
nand U48930 (N_48930,N_47295,N_47285);
or U48931 (N_48931,N_46195,N_45112);
nand U48932 (N_48932,N_47030,N_45347);
or U48933 (N_48933,N_46909,N_46742);
nor U48934 (N_48934,N_47044,N_45705);
nand U48935 (N_48935,N_45811,N_46028);
and U48936 (N_48936,N_45489,N_45112);
nand U48937 (N_48937,N_45675,N_46294);
nor U48938 (N_48938,N_46007,N_46812);
xnor U48939 (N_48939,N_46487,N_45364);
or U48940 (N_48940,N_46968,N_45483);
xor U48941 (N_48941,N_47234,N_46355);
nand U48942 (N_48942,N_46737,N_45026);
or U48943 (N_48943,N_46332,N_47229);
nand U48944 (N_48944,N_45780,N_45277);
and U48945 (N_48945,N_46967,N_47089);
or U48946 (N_48946,N_47030,N_45887);
nand U48947 (N_48947,N_46275,N_47251);
or U48948 (N_48948,N_47199,N_45990);
nor U48949 (N_48949,N_46322,N_45861);
nand U48950 (N_48950,N_45253,N_47235);
xnor U48951 (N_48951,N_47372,N_46511);
nand U48952 (N_48952,N_45881,N_45266);
nand U48953 (N_48953,N_46913,N_46707);
xnor U48954 (N_48954,N_47424,N_46686);
nand U48955 (N_48955,N_46903,N_46178);
nor U48956 (N_48956,N_47474,N_45641);
nor U48957 (N_48957,N_47043,N_47280);
nor U48958 (N_48958,N_46923,N_46682);
and U48959 (N_48959,N_45307,N_45275);
and U48960 (N_48960,N_45797,N_47162);
nor U48961 (N_48961,N_45253,N_46337);
xor U48962 (N_48962,N_47171,N_47227);
nor U48963 (N_48963,N_46847,N_47187);
xnor U48964 (N_48964,N_46201,N_45734);
and U48965 (N_48965,N_45328,N_47350);
xor U48966 (N_48966,N_45177,N_46349);
nor U48967 (N_48967,N_46066,N_45554);
or U48968 (N_48968,N_47377,N_46753);
xor U48969 (N_48969,N_45014,N_46446);
nor U48970 (N_48970,N_46233,N_47099);
nand U48971 (N_48971,N_45274,N_45825);
or U48972 (N_48972,N_45836,N_46687);
or U48973 (N_48973,N_47373,N_46275);
xnor U48974 (N_48974,N_45197,N_47107);
and U48975 (N_48975,N_45065,N_45335);
nor U48976 (N_48976,N_47317,N_46729);
xor U48977 (N_48977,N_46138,N_46018);
and U48978 (N_48978,N_47301,N_46994);
nor U48979 (N_48979,N_46510,N_46609);
and U48980 (N_48980,N_47032,N_46050);
or U48981 (N_48981,N_46963,N_46333);
or U48982 (N_48982,N_46634,N_45768);
nor U48983 (N_48983,N_46581,N_46026);
nand U48984 (N_48984,N_46763,N_46807);
nor U48985 (N_48985,N_46663,N_45517);
and U48986 (N_48986,N_47384,N_45035);
xnor U48987 (N_48987,N_45326,N_46014);
xor U48988 (N_48988,N_47347,N_46953);
nand U48989 (N_48989,N_47447,N_47382);
nor U48990 (N_48990,N_46285,N_46424);
xnor U48991 (N_48991,N_46331,N_46169);
nand U48992 (N_48992,N_47037,N_46564);
nor U48993 (N_48993,N_45840,N_47126);
xor U48994 (N_48994,N_46674,N_47440);
nor U48995 (N_48995,N_47142,N_45699);
nor U48996 (N_48996,N_45904,N_46836);
and U48997 (N_48997,N_45902,N_46053);
nand U48998 (N_48998,N_45732,N_46439);
and U48999 (N_48999,N_46165,N_45214);
nand U49000 (N_49000,N_45957,N_47067);
xor U49001 (N_49001,N_45801,N_47205);
or U49002 (N_49002,N_46328,N_46625);
nand U49003 (N_49003,N_47286,N_47140);
xnor U49004 (N_49004,N_46820,N_45613);
and U49005 (N_49005,N_46906,N_46037);
and U49006 (N_49006,N_46268,N_47427);
xor U49007 (N_49007,N_45121,N_46347);
and U49008 (N_49008,N_46463,N_46482);
and U49009 (N_49009,N_45057,N_45650);
nand U49010 (N_49010,N_45492,N_46585);
nor U49011 (N_49011,N_46025,N_46698);
nand U49012 (N_49012,N_47260,N_45540);
and U49013 (N_49013,N_46260,N_45866);
nand U49014 (N_49014,N_47472,N_46337);
and U49015 (N_49015,N_45056,N_45065);
or U49016 (N_49016,N_46268,N_46889);
and U49017 (N_49017,N_46154,N_45591);
or U49018 (N_49018,N_47383,N_45087);
nand U49019 (N_49019,N_45567,N_46306);
xnor U49020 (N_49020,N_45625,N_46878);
or U49021 (N_49021,N_46890,N_45165);
xnor U49022 (N_49022,N_46028,N_45708);
nor U49023 (N_49023,N_45140,N_45213);
and U49024 (N_49024,N_47145,N_46211);
and U49025 (N_49025,N_45060,N_46082);
and U49026 (N_49026,N_47020,N_45989);
or U49027 (N_49027,N_46730,N_46738);
nand U49028 (N_49028,N_46589,N_46159);
nand U49029 (N_49029,N_45489,N_46172);
nor U49030 (N_49030,N_46412,N_46168);
nand U49031 (N_49031,N_45789,N_46579);
and U49032 (N_49032,N_46231,N_45880);
and U49033 (N_49033,N_47056,N_45379);
xor U49034 (N_49034,N_47111,N_45268);
nand U49035 (N_49035,N_46490,N_47146);
and U49036 (N_49036,N_46739,N_46404);
nor U49037 (N_49037,N_46525,N_47455);
nand U49038 (N_49038,N_46985,N_45306);
and U49039 (N_49039,N_45247,N_46920);
nand U49040 (N_49040,N_46314,N_46399);
and U49041 (N_49041,N_46136,N_46905);
nand U49042 (N_49042,N_46216,N_46923);
or U49043 (N_49043,N_46588,N_46379);
xor U49044 (N_49044,N_46031,N_45957);
xor U49045 (N_49045,N_46100,N_45899);
xor U49046 (N_49046,N_47092,N_45344);
xnor U49047 (N_49047,N_46714,N_45996);
xor U49048 (N_49048,N_45330,N_46678);
or U49049 (N_49049,N_46647,N_45521);
nor U49050 (N_49050,N_46496,N_47006);
nand U49051 (N_49051,N_45018,N_45371);
nor U49052 (N_49052,N_45984,N_47280);
nand U49053 (N_49053,N_46999,N_46125);
or U49054 (N_49054,N_46962,N_45665);
and U49055 (N_49055,N_45538,N_45012);
xor U49056 (N_49056,N_45537,N_46893);
nor U49057 (N_49057,N_47061,N_45897);
xnor U49058 (N_49058,N_45058,N_45371);
nand U49059 (N_49059,N_46033,N_46515);
and U49060 (N_49060,N_46923,N_46652);
nor U49061 (N_49061,N_45751,N_45028);
nand U49062 (N_49062,N_46141,N_46647);
nor U49063 (N_49063,N_46406,N_47301);
nor U49064 (N_49064,N_46268,N_46930);
xor U49065 (N_49065,N_46404,N_45225);
or U49066 (N_49066,N_47101,N_45071);
and U49067 (N_49067,N_46829,N_46853);
xnor U49068 (N_49068,N_47337,N_45874);
nor U49069 (N_49069,N_45409,N_45376);
xnor U49070 (N_49070,N_47071,N_46744);
xnor U49071 (N_49071,N_45046,N_47395);
xnor U49072 (N_49072,N_45772,N_45671);
and U49073 (N_49073,N_45455,N_47486);
and U49074 (N_49074,N_45783,N_46651);
nand U49075 (N_49075,N_47499,N_45284);
nand U49076 (N_49076,N_46670,N_46115);
nand U49077 (N_49077,N_45018,N_46808);
nand U49078 (N_49078,N_46497,N_45021);
nand U49079 (N_49079,N_46565,N_45015);
nand U49080 (N_49080,N_46784,N_45044);
xnor U49081 (N_49081,N_45688,N_45689);
and U49082 (N_49082,N_47281,N_46569);
nor U49083 (N_49083,N_45876,N_47296);
or U49084 (N_49084,N_45240,N_46953);
or U49085 (N_49085,N_46457,N_45289);
nand U49086 (N_49086,N_46615,N_46757);
and U49087 (N_49087,N_46324,N_45496);
xnor U49088 (N_49088,N_47478,N_46709);
and U49089 (N_49089,N_47375,N_46963);
nand U49090 (N_49090,N_46537,N_46876);
xor U49091 (N_49091,N_45629,N_45045);
nand U49092 (N_49092,N_45928,N_46289);
and U49093 (N_49093,N_46999,N_45651);
nand U49094 (N_49094,N_46664,N_45806);
xnor U49095 (N_49095,N_47190,N_45694);
nor U49096 (N_49096,N_45492,N_45449);
or U49097 (N_49097,N_45068,N_46196);
xnor U49098 (N_49098,N_47038,N_45646);
nand U49099 (N_49099,N_47208,N_47068);
nor U49100 (N_49100,N_45514,N_45713);
or U49101 (N_49101,N_46618,N_45044);
or U49102 (N_49102,N_46535,N_45436);
nor U49103 (N_49103,N_45274,N_46519);
xor U49104 (N_49104,N_45673,N_46598);
or U49105 (N_49105,N_46934,N_45891);
or U49106 (N_49106,N_45496,N_47075);
nor U49107 (N_49107,N_45594,N_47208);
or U49108 (N_49108,N_45063,N_47106);
or U49109 (N_49109,N_45292,N_46051);
nor U49110 (N_49110,N_45490,N_45203);
xor U49111 (N_49111,N_47252,N_46765);
or U49112 (N_49112,N_45982,N_45493);
xnor U49113 (N_49113,N_45729,N_46560);
or U49114 (N_49114,N_45275,N_46379);
nand U49115 (N_49115,N_47092,N_45630);
and U49116 (N_49116,N_45197,N_46782);
or U49117 (N_49117,N_46615,N_46715);
xnor U49118 (N_49118,N_45564,N_46798);
nor U49119 (N_49119,N_47018,N_45765);
nor U49120 (N_49120,N_45948,N_46309);
xnor U49121 (N_49121,N_46485,N_46396);
and U49122 (N_49122,N_46328,N_46176);
or U49123 (N_49123,N_46677,N_45083);
xnor U49124 (N_49124,N_47218,N_46464);
xnor U49125 (N_49125,N_45142,N_45795);
or U49126 (N_49126,N_46690,N_45013);
xnor U49127 (N_49127,N_45096,N_46349);
xnor U49128 (N_49128,N_45811,N_46521);
or U49129 (N_49129,N_45775,N_45432);
xnor U49130 (N_49130,N_46457,N_46340);
xor U49131 (N_49131,N_47213,N_45033);
and U49132 (N_49132,N_45087,N_46834);
nand U49133 (N_49133,N_47246,N_46398);
and U49134 (N_49134,N_45832,N_45087);
nand U49135 (N_49135,N_45374,N_47395);
nor U49136 (N_49136,N_47096,N_46505);
xor U49137 (N_49137,N_45735,N_46303);
nand U49138 (N_49138,N_45295,N_45698);
xnor U49139 (N_49139,N_45684,N_46381);
nor U49140 (N_49140,N_46930,N_45935);
nor U49141 (N_49141,N_46653,N_45050);
xnor U49142 (N_49142,N_46504,N_46826);
nor U49143 (N_49143,N_46896,N_46407);
xnor U49144 (N_49144,N_46450,N_46943);
nor U49145 (N_49145,N_46183,N_47060);
nand U49146 (N_49146,N_47131,N_45920);
xor U49147 (N_49147,N_45708,N_46711);
xnor U49148 (N_49148,N_46147,N_46558);
nor U49149 (N_49149,N_45467,N_45752);
xor U49150 (N_49150,N_47052,N_46585);
and U49151 (N_49151,N_46336,N_45671);
or U49152 (N_49152,N_45202,N_47375);
xor U49153 (N_49153,N_47206,N_47094);
or U49154 (N_49154,N_46552,N_45089);
and U49155 (N_49155,N_45237,N_47150);
and U49156 (N_49156,N_45513,N_45175);
or U49157 (N_49157,N_45965,N_45787);
and U49158 (N_49158,N_46768,N_45226);
nor U49159 (N_49159,N_47358,N_46945);
nor U49160 (N_49160,N_46271,N_45301);
or U49161 (N_49161,N_46214,N_45518);
and U49162 (N_49162,N_46597,N_46764);
or U49163 (N_49163,N_46374,N_46122);
nor U49164 (N_49164,N_46627,N_46917);
or U49165 (N_49165,N_45242,N_46411);
and U49166 (N_49166,N_45865,N_45045);
and U49167 (N_49167,N_46273,N_46826);
nand U49168 (N_49168,N_46647,N_45892);
xor U49169 (N_49169,N_47194,N_45768);
nor U49170 (N_49170,N_45955,N_45356);
and U49171 (N_49171,N_47006,N_46597);
xnor U49172 (N_49172,N_45754,N_45508);
and U49173 (N_49173,N_47009,N_45592);
or U49174 (N_49174,N_45952,N_46099);
and U49175 (N_49175,N_47180,N_47451);
or U49176 (N_49176,N_45707,N_46250);
nand U49177 (N_49177,N_46552,N_45458);
or U49178 (N_49178,N_45680,N_45847);
or U49179 (N_49179,N_47231,N_45848);
nand U49180 (N_49180,N_45021,N_46082);
nand U49181 (N_49181,N_45216,N_47334);
xnor U49182 (N_49182,N_45236,N_46636);
or U49183 (N_49183,N_47391,N_47002);
or U49184 (N_49184,N_45450,N_45668);
xor U49185 (N_49185,N_45587,N_47367);
or U49186 (N_49186,N_45838,N_45487);
xor U49187 (N_49187,N_45372,N_46155);
or U49188 (N_49188,N_45412,N_45084);
or U49189 (N_49189,N_45068,N_46630);
nand U49190 (N_49190,N_47070,N_47072);
nand U49191 (N_49191,N_45185,N_47172);
xor U49192 (N_49192,N_46645,N_45466);
nor U49193 (N_49193,N_47139,N_46298);
xor U49194 (N_49194,N_47254,N_46907);
nand U49195 (N_49195,N_47167,N_46847);
nor U49196 (N_49196,N_47227,N_45901);
or U49197 (N_49197,N_45951,N_45796);
or U49198 (N_49198,N_46616,N_47367);
nand U49199 (N_49199,N_45124,N_45600);
or U49200 (N_49200,N_46123,N_45941);
nand U49201 (N_49201,N_46922,N_46115);
nor U49202 (N_49202,N_46313,N_47418);
nor U49203 (N_49203,N_45106,N_46159);
xor U49204 (N_49204,N_45326,N_46303);
or U49205 (N_49205,N_47073,N_46965);
and U49206 (N_49206,N_46488,N_45030);
nand U49207 (N_49207,N_46867,N_46361);
nor U49208 (N_49208,N_45294,N_46771);
and U49209 (N_49209,N_46260,N_47058);
xor U49210 (N_49210,N_45591,N_45900);
or U49211 (N_49211,N_47020,N_45795);
nand U49212 (N_49212,N_45964,N_46869);
and U49213 (N_49213,N_45206,N_46921);
nand U49214 (N_49214,N_45371,N_45143);
or U49215 (N_49215,N_47236,N_47153);
or U49216 (N_49216,N_47425,N_45144);
or U49217 (N_49217,N_47003,N_46674);
and U49218 (N_49218,N_45232,N_45851);
or U49219 (N_49219,N_45972,N_45340);
nor U49220 (N_49220,N_46378,N_46900);
and U49221 (N_49221,N_45822,N_46683);
and U49222 (N_49222,N_47476,N_45051);
or U49223 (N_49223,N_46287,N_46599);
or U49224 (N_49224,N_47115,N_45806);
nor U49225 (N_49225,N_45571,N_46803);
nor U49226 (N_49226,N_45615,N_45947);
or U49227 (N_49227,N_45082,N_45067);
nand U49228 (N_49228,N_45432,N_45794);
nor U49229 (N_49229,N_45242,N_46863);
and U49230 (N_49230,N_46384,N_46239);
nand U49231 (N_49231,N_45633,N_46504);
or U49232 (N_49232,N_45854,N_45266);
xnor U49233 (N_49233,N_46587,N_47461);
nand U49234 (N_49234,N_47323,N_46222);
and U49235 (N_49235,N_47144,N_45508);
xor U49236 (N_49236,N_46968,N_46626);
or U49237 (N_49237,N_45882,N_46205);
nor U49238 (N_49238,N_47414,N_46096);
nand U49239 (N_49239,N_45272,N_45707);
and U49240 (N_49240,N_46874,N_45619);
nand U49241 (N_49241,N_47465,N_45009);
nor U49242 (N_49242,N_46392,N_47173);
nand U49243 (N_49243,N_47329,N_47309);
nand U49244 (N_49244,N_45472,N_47207);
xnor U49245 (N_49245,N_45642,N_45254);
or U49246 (N_49246,N_47198,N_45313);
xnor U49247 (N_49247,N_45937,N_47356);
or U49248 (N_49248,N_45599,N_47451);
and U49249 (N_49249,N_46571,N_45001);
and U49250 (N_49250,N_46232,N_45722);
nand U49251 (N_49251,N_46695,N_45248);
nor U49252 (N_49252,N_45005,N_47224);
or U49253 (N_49253,N_46286,N_46658);
and U49254 (N_49254,N_45599,N_47286);
nor U49255 (N_49255,N_46339,N_45088);
nor U49256 (N_49256,N_45327,N_46650);
or U49257 (N_49257,N_46807,N_46552);
nor U49258 (N_49258,N_46473,N_47167);
nor U49259 (N_49259,N_46501,N_45103);
nor U49260 (N_49260,N_45053,N_45659);
nor U49261 (N_49261,N_46061,N_46390);
nand U49262 (N_49262,N_47052,N_46567);
nor U49263 (N_49263,N_46145,N_45515);
xnor U49264 (N_49264,N_46022,N_46330);
nand U49265 (N_49265,N_45492,N_47331);
nor U49266 (N_49266,N_46963,N_45954);
xnor U49267 (N_49267,N_45622,N_45556);
and U49268 (N_49268,N_46015,N_47278);
and U49269 (N_49269,N_45411,N_45892);
or U49270 (N_49270,N_46536,N_45542);
nand U49271 (N_49271,N_45855,N_46665);
or U49272 (N_49272,N_46901,N_47241);
nand U49273 (N_49273,N_47170,N_45917);
and U49274 (N_49274,N_45836,N_46303);
and U49275 (N_49275,N_46989,N_45141);
nor U49276 (N_49276,N_47451,N_45982);
nand U49277 (N_49277,N_45414,N_45545);
nand U49278 (N_49278,N_46596,N_47364);
nor U49279 (N_49279,N_46812,N_47267);
and U49280 (N_49280,N_46939,N_45234);
xor U49281 (N_49281,N_46146,N_47350);
and U49282 (N_49282,N_45267,N_45572);
xnor U49283 (N_49283,N_45209,N_46015);
and U49284 (N_49284,N_47206,N_47455);
and U49285 (N_49285,N_46454,N_46237);
nor U49286 (N_49286,N_46118,N_46745);
nand U49287 (N_49287,N_45846,N_46263);
xnor U49288 (N_49288,N_45922,N_46648);
and U49289 (N_49289,N_45752,N_46196);
xnor U49290 (N_49290,N_45459,N_47420);
nor U49291 (N_49291,N_45553,N_45247);
xor U49292 (N_49292,N_45937,N_45139);
xnor U49293 (N_49293,N_47346,N_45788);
and U49294 (N_49294,N_45331,N_46948);
xnor U49295 (N_49295,N_46532,N_46012);
nand U49296 (N_49296,N_45827,N_46926);
and U49297 (N_49297,N_47007,N_46483);
xor U49298 (N_49298,N_46214,N_46215);
and U49299 (N_49299,N_45434,N_45933);
or U49300 (N_49300,N_46254,N_46204);
xnor U49301 (N_49301,N_46970,N_47004);
nor U49302 (N_49302,N_46620,N_46478);
nor U49303 (N_49303,N_47004,N_45908);
and U49304 (N_49304,N_46274,N_45773);
or U49305 (N_49305,N_46047,N_47486);
xor U49306 (N_49306,N_46490,N_46829);
and U49307 (N_49307,N_45636,N_46123);
nand U49308 (N_49308,N_46296,N_47019);
nor U49309 (N_49309,N_47457,N_46888);
and U49310 (N_49310,N_46067,N_46692);
nor U49311 (N_49311,N_47402,N_46782);
and U49312 (N_49312,N_45786,N_47491);
and U49313 (N_49313,N_46360,N_46104);
nand U49314 (N_49314,N_45037,N_47481);
xnor U49315 (N_49315,N_46300,N_46612);
or U49316 (N_49316,N_46062,N_45744);
xor U49317 (N_49317,N_46170,N_45414);
or U49318 (N_49318,N_45603,N_45136);
xnor U49319 (N_49319,N_47252,N_46101);
nand U49320 (N_49320,N_45110,N_47100);
nor U49321 (N_49321,N_45102,N_46747);
and U49322 (N_49322,N_46989,N_47473);
or U49323 (N_49323,N_45052,N_45852);
xnor U49324 (N_49324,N_46507,N_45205);
nand U49325 (N_49325,N_47221,N_45133);
or U49326 (N_49326,N_47346,N_46250);
nor U49327 (N_49327,N_47494,N_46909);
or U49328 (N_49328,N_46609,N_46431);
nor U49329 (N_49329,N_46523,N_46034);
nor U49330 (N_49330,N_46149,N_45209);
and U49331 (N_49331,N_46257,N_45951);
or U49332 (N_49332,N_45128,N_47081);
nand U49333 (N_49333,N_47053,N_45367);
or U49334 (N_49334,N_46419,N_46361);
nand U49335 (N_49335,N_47220,N_45751);
nand U49336 (N_49336,N_45198,N_47406);
and U49337 (N_49337,N_45351,N_45416);
nor U49338 (N_49338,N_46680,N_46575);
and U49339 (N_49339,N_47013,N_47422);
nand U49340 (N_49340,N_45687,N_46676);
or U49341 (N_49341,N_45709,N_47390);
xor U49342 (N_49342,N_47029,N_45048);
xor U49343 (N_49343,N_47057,N_46029);
nor U49344 (N_49344,N_46113,N_47026);
or U49345 (N_49345,N_47343,N_45008);
xor U49346 (N_49346,N_46841,N_45380);
nand U49347 (N_49347,N_46971,N_47077);
and U49348 (N_49348,N_45564,N_45404);
nor U49349 (N_49349,N_46681,N_45159);
and U49350 (N_49350,N_46234,N_47260);
or U49351 (N_49351,N_45802,N_46843);
and U49352 (N_49352,N_45597,N_47296);
and U49353 (N_49353,N_45178,N_46364);
or U49354 (N_49354,N_45366,N_45630);
nor U49355 (N_49355,N_47101,N_47349);
xor U49356 (N_49356,N_47181,N_46774);
and U49357 (N_49357,N_45640,N_45752);
and U49358 (N_49358,N_45926,N_46269);
nor U49359 (N_49359,N_45564,N_46107);
nand U49360 (N_49360,N_45865,N_46517);
nor U49361 (N_49361,N_46291,N_46392);
and U49362 (N_49362,N_45329,N_46195);
or U49363 (N_49363,N_45159,N_47109);
or U49364 (N_49364,N_46588,N_47408);
xor U49365 (N_49365,N_46944,N_47489);
and U49366 (N_49366,N_46357,N_46521);
nand U49367 (N_49367,N_45646,N_45694);
nand U49368 (N_49368,N_46833,N_47263);
or U49369 (N_49369,N_46249,N_46753);
nor U49370 (N_49370,N_47169,N_45163);
nor U49371 (N_49371,N_45109,N_45167);
and U49372 (N_49372,N_45793,N_45277);
xor U49373 (N_49373,N_47202,N_47156);
or U49374 (N_49374,N_45134,N_45602);
or U49375 (N_49375,N_45156,N_45086);
nor U49376 (N_49376,N_45977,N_47219);
xor U49377 (N_49377,N_45382,N_46486);
or U49378 (N_49378,N_46731,N_47138);
xor U49379 (N_49379,N_45323,N_45593);
nand U49380 (N_49380,N_45106,N_45355);
nor U49381 (N_49381,N_46316,N_45549);
nand U49382 (N_49382,N_45819,N_46244);
nor U49383 (N_49383,N_45043,N_45957);
or U49384 (N_49384,N_45588,N_47177);
xor U49385 (N_49385,N_45520,N_45856);
xor U49386 (N_49386,N_46604,N_46426);
nand U49387 (N_49387,N_45334,N_45737);
nand U49388 (N_49388,N_45153,N_45280);
nor U49389 (N_49389,N_46825,N_45031);
xnor U49390 (N_49390,N_47065,N_45101);
or U49391 (N_49391,N_46031,N_46829);
and U49392 (N_49392,N_45953,N_47385);
nand U49393 (N_49393,N_47389,N_46980);
nor U49394 (N_49394,N_46857,N_46070);
and U49395 (N_49395,N_45127,N_47066);
nand U49396 (N_49396,N_47114,N_45311);
xnor U49397 (N_49397,N_46877,N_47118);
and U49398 (N_49398,N_45176,N_46011);
xnor U49399 (N_49399,N_47370,N_45152);
and U49400 (N_49400,N_47054,N_47150);
nand U49401 (N_49401,N_45963,N_46151);
and U49402 (N_49402,N_46414,N_46764);
nor U49403 (N_49403,N_45567,N_45600);
nand U49404 (N_49404,N_47009,N_46837);
nand U49405 (N_49405,N_46967,N_46910);
xor U49406 (N_49406,N_46211,N_45012);
nand U49407 (N_49407,N_46463,N_46800);
xnor U49408 (N_49408,N_45058,N_45166);
xor U49409 (N_49409,N_46577,N_46121);
and U49410 (N_49410,N_46607,N_47257);
nor U49411 (N_49411,N_45188,N_47285);
xnor U49412 (N_49412,N_45728,N_46933);
nor U49413 (N_49413,N_46272,N_46747);
nand U49414 (N_49414,N_45070,N_45247);
nor U49415 (N_49415,N_45149,N_45103);
nand U49416 (N_49416,N_45433,N_45684);
xor U49417 (N_49417,N_46870,N_45002);
nor U49418 (N_49418,N_47290,N_45091);
nor U49419 (N_49419,N_46619,N_45703);
nand U49420 (N_49420,N_47152,N_46443);
nor U49421 (N_49421,N_46330,N_45601);
xor U49422 (N_49422,N_46148,N_45810);
nor U49423 (N_49423,N_45163,N_46831);
nor U49424 (N_49424,N_45816,N_45455);
and U49425 (N_49425,N_47308,N_45632);
nand U49426 (N_49426,N_45744,N_47190);
nand U49427 (N_49427,N_47155,N_45244);
nand U49428 (N_49428,N_45133,N_45944);
or U49429 (N_49429,N_45861,N_45522);
nand U49430 (N_49430,N_46576,N_45903);
and U49431 (N_49431,N_46173,N_46095);
and U49432 (N_49432,N_47288,N_46013);
nor U49433 (N_49433,N_47429,N_47276);
xor U49434 (N_49434,N_47231,N_45198);
and U49435 (N_49435,N_47129,N_46925);
or U49436 (N_49436,N_46253,N_45116);
xor U49437 (N_49437,N_45314,N_45716);
or U49438 (N_49438,N_47487,N_46847);
or U49439 (N_49439,N_46462,N_46329);
xnor U49440 (N_49440,N_45495,N_47014);
xor U49441 (N_49441,N_45784,N_45860);
xor U49442 (N_49442,N_46687,N_45426);
nand U49443 (N_49443,N_45148,N_45421);
nand U49444 (N_49444,N_46645,N_46227);
nor U49445 (N_49445,N_45691,N_45678);
and U49446 (N_49446,N_46091,N_45291);
or U49447 (N_49447,N_45938,N_46741);
or U49448 (N_49448,N_46002,N_47449);
and U49449 (N_49449,N_45879,N_47413);
nor U49450 (N_49450,N_47090,N_45124);
nand U49451 (N_49451,N_46989,N_45901);
and U49452 (N_49452,N_46287,N_45427);
and U49453 (N_49453,N_46918,N_45669);
nor U49454 (N_49454,N_47461,N_45258);
nor U49455 (N_49455,N_45921,N_45692);
or U49456 (N_49456,N_46661,N_47277);
nor U49457 (N_49457,N_46312,N_45007);
or U49458 (N_49458,N_45967,N_46917);
and U49459 (N_49459,N_46347,N_46754);
or U49460 (N_49460,N_46731,N_46501);
or U49461 (N_49461,N_46379,N_46213);
nor U49462 (N_49462,N_45395,N_47493);
or U49463 (N_49463,N_46570,N_45861);
nor U49464 (N_49464,N_45294,N_46868);
nor U49465 (N_49465,N_47172,N_45491);
xor U49466 (N_49466,N_46755,N_46932);
or U49467 (N_49467,N_45066,N_45942);
nor U49468 (N_49468,N_45569,N_47278);
or U49469 (N_49469,N_45040,N_47200);
nor U49470 (N_49470,N_46346,N_45754);
nand U49471 (N_49471,N_47472,N_47309);
nand U49472 (N_49472,N_45610,N_47085);
or U49473 (N_49473,N_45934,N_45685);
and U49474 (N_49474,N_45516,N_47176);
nand U49475 (N_49475,N_46352,N_46861);
xor U49476 (N_49476,N_47100,N_46523);
or U49477 (N_49477,N_45503,N_45555);
nor U49478 (N_49478,N_46042,N_45934);
and U49479 (N_49479,N_45473,N_46697);
xor U49480 (N_49480,N_46601,N_46486);
nand U49481 (N_49481,N_46130,N_46163);
nand U49482 (N_49482,N_46325,N_45171);
xor U49483 (N_49483,N_46959,N_46502);
nand U49484 (N_49484,N_47465,N_45850);
xor U49485 (N_49485,N_47238,N_46815);
and U49486 (N_49486,N_46690,N_45652);
or U49487 (N_49487,N_45545,N_45547);
nor U49488 (N_49488,N_47449,N_45441);
xor U49489 (N_49489,N_46230,N_45069);
nand U49490 (N_49490,N_46587,N_46387);
or U49491 (N_49491,N_45816,N_46942);
nand U49492 (N_49492,N_45340,N_46111);
nand U49493 (N_49493,N_47183,N_47269);
xnor U49494 (N_49494,N_45369,N_47305);
and U49495 (N_49495,N_46224,N_47300);
nand U49496 (N_49496,N_47120,N_45664);
nand U49497 (N_49497,N_46387,N_46121);
nand U49498 (N_49498,N_45006,N_47288);
nor U49499 (N_49499,N_46303,N_45161);
or U49500 (N_49500,N_47282,N_45891);
or U49501 (N_49501,N_45773,N_45878);
nor U49502 (N_49502,N_46837,N_45304);
xor U49503 (N_49503,N_45749,N_46694);
nor U49504 (N_49504,N_45085,N_46480);
nand U49505 (N_49505,N_47239,N_47475);
nor U49506 (N_49506,N_46102,N_45235);
or U49507 (N_49507,N_46390,N_45525);
nand U49508 (N_49508,N_46853,N_46258);
nand U49509 (N_49509,N_47215,N_47345);
nor U49510 (N_49510,N_46774,N_46230);
or U49511 (N_49511,N_45715,N_46411);
xor U49512 (N_49512,N_47446,N_45846);
nand U49513 (N_49513,N_46645,N_46804);
xnor U49514 (N_49514,N_45611,N_46713);
and U49515 (N_49515,N_45450,N_46756);
nand U49516 (N_49516,N_45413,N_46007);
nand U49517 (N_49517,N_45175,N_46715);
xor U49518 (N_49518,N_45753,N_46364);
xor U49519 (N_49519,N_46227,N_46789);
nand U49520 (N_49520,N_45701,N_45335);
nor U49521 (N_49521,N_45660,N_46051);
xnor U49522 (N_49522,N_46346,N_46820);
and U49523 (N_49523,N_45757,N_46865);
nand U49524 (N_49524,N_45581,N_47143);
and U49525 (N_49525,N_45490,N_47161);
xor U49526 (N_49526,N_45698,N_45321);
xnor U49527 (N_49527,N_45655,N_46957);
nand U49528 (N_49528,N_46401,N_47340);
nand U49529 (N_49529,N_45990,N_45989);
and U49530 (N_49530,N_47066,N_47315);
and U49531 (N_49531,N_45270,N_45078);
nor U49532 (N_49532,N_46888,N_45151);
or U49533 (N_49533,N_46860,N_46815);
xor U49534 (N_49534,N_47068,N_45876);
or U49535 (N_49535,N_46460,N_45055);
nand U49536 (N_49536,N_45500,N_46195);
nand U49537 (N_49537,N_46777,N_46508);
and U49538 (N_49538,N_46268,N_46042);
nor U49539 (N_49539,N_45693,N_47055);
nor U49540 (N_49540,N_46758,N_46238);
and U49541 (N_49541,N_46453,N_45142);
nor U49542 (N_49542,N_45708,N_46193);
nor U49543 (N_49543,N_45389,N_45154);
nor U49544 (N_49544,N_46102,N_45170);
or U49545 (N_49545,N_45169,N_46789);
nor U49546 (N_49546,N_45649,N_45632);
nand U49547 (N_49547,N_45567,N_46134);
nor U49548 (N_49548,N_46972,N_46387);
xnor U49549 (N_49549,N_46379,N_46614);
nor U49550 (N_49550,N_45044,N_47431);
nor U49551 (N_49551,N_46339,N_45621);
nand U49552 (N_49552,N_45494,N_46882);
nand U49553 (N_49553,N_46136,N_45740);
or U49554 (N_49554,N_45275,N_45285);
and U49555 (N_49555,N_46263,N_45902);
xnor U49556 (N_49556,N_46973,N_47121);
and U49557 (N_49557,N_45045,N_47117);
or U49558 (N_49558,N_45623,N_45931);
and U49559 (N_49559,N_46562,N_46088);
nor U49560 (N_49560,N_46534,N_45815);
and U49561 (N_49561,N_45505,N_46619);
or U49562 (N_49562,N_45974,N_45592);
nand U49563 (N_49563,N_45813,N_46392);
nand U49564 (N_49564,N_46659,N_45552);
and U49565 (N_49565,N_45852,N_45681);
xnor U49566 (N_49566,N_45777,N_45617);
or U49567 (N_49567,N_47241,N_46871);
nand U49568 (N_49568,N_45421,N_46511);
or U49569 (N_49569,N_46417,N_47067);
nor U49570 (N_49570,N_47407,N_46825);
or U49571 (N_49571,N_45946,N_45820);
xor U49572 (N_49572,N_45244,N_46423);
or U49573 (N_49573,N_46381,N_45470);
nor U49574 (N_49574,N_45988,N_45982);
nor U49575 (N_49575,N_46437,N_46313);
or U49576 (N_49576,N_46403,N_45371);
nand U49577 (N_49577,N_47012,N_47297);
or U49578 (N_49578,N_46971,N_45093);
and U49579 (N_49579,N_45590,N_46320);
nor U49580 (N_49580,N_45711,N_47380);
or U49581 (N_49581,N_45662,N_46283);
nor U49582 (N_49582,N_45734,N_47208);
and U49583 (N_49583,N_47499,N_45012);
and U49584 (N_49584,N_46671,N_45091);
xnor U49585 (N_49585,N_45528,N_45883);
or U49586 (N_49586,N_46460,N_46506);
or U49587 (N_49587,N_45591,N_46195);
nor U49588 (N_49588,N_45313,N_45741);
nor U49589 (N_49589,N_45686,N_46473);
nor U49590 (N_49590,N_46728,N_46071);
nand U49591 (N_49591,N_46302,N_45849);
xor U49592 (N_49592,N_46096,N_46536);
or U49593 (N_49593,N_46832,N_47083);
or U49594 (N_49594,N_46815,N_46201);
xor U49595 (N_49595,N_45859,N_46983);
xor U49596 (N_49596,N_46874,N_45296);
or U49597 (N_49597,N_45865,N_47105);
nor U49598 (N_49598,N_47492,N_47215);
and U49599 (N_49599,N_47158,N_47185);
and U49600 (N_49600,N_46197,N_45349);
or U49601 (N_49601,N_45643,N_45388);
nand U49602 (N_49602,N_46002,N_45871);
or U49603 (N_49603,N_46315,N_45152);
xor U49604 (N_49604,N_45075,N_47041);
nor U49605 (N_49605,N_45173,N_45471);
and U49606 (N_49606,N_47340,N_46726);
xor U49607 (N_49607,N_46986,N_45375);
nand U49608 (N_49608,N_45008,N_47110);
and U49609 (N_49609,N_46314,N_45441);
nand U49610 (N_49610,N_45707,N_47235);
and U49611 (N_49611,N_45258,N_47052);
xor U49612 (N_49612,N_45464,N_46644);
or U49613 (N_49613,N_46875,N_46592);
or U49614 (N_49614,N_47024,N_46591);
nand U49615 (N_49615,N_45652,N_45426);
and U49616 (N_49616,N_47043,N_47472);
nand U49617 (N_49617,N_46192,N_46852);
or U49618 (N_49618,N_45493,N_45701);
xnor U49619 (N_49619,N_47012,N_46297);
nor U49620 (N_49620,N_45054,N_45183);
and U49621 (N_49621,N_45776,N_45988);
and U49622 (N_49622,N_45976,N_46421);
xor U49623 (N_49623,N_47023,N_45165);
nand U49624 (N_49624,N_45006,N_45351);
or U49625 (N_49625,N_46773,N_47369);
xnor U49626 (N_49626,N_46406,N_46906);
nor U49627 (N_49627,N_45751,N_46429);
nand U49628 (N_49628,N_46078,N_46975);
or U49629 (N_49629,N_45975,N_46765);
or U49630 (N_49630,N_46556,N_47188);
or U49631 (N_49631,N_45974,N_45099);
and U49632 (N_49632,N_45423,N_46815);
and U49633 (N_49633,N_46962,N_45331);
and U49634 (N_49634,N_47421,N_45991);
nand U49635 (N_49635,N_47428,N_45557);
or U49636 (N_49636,N_45252,N_46867);
or U49637 (N_49637,N_45731,N_46535);
or U49638 (N_49638,N_45357,N_46203);
and U49639 (N_49639,N_45230,N_47256);
and U49640 (N_49640,N_45594,N_45904);
nand U49641 (N_49641,N_46304,N_47122);
or U49642 (N_49642,N_45827,N_47204);
nand U49643 (N_49643,N_47252,N_46214);
nor U49644 (N_49644,N_47264,N_45011);
nand U49645 (N_49645,N_45067,N_46603);
or U49646 (N_49646,N_45615,N_45116);
xnor U49647 (N_49647,N_46039,N_47175);
nand U49648 (N_49648,N_47170,N_45703);
nand U49649 (N_49649,N_47042,N_45158);
nor U49650 (N_49650,N_46777,N_45318);
nor U49651 (N_49651,N_45748,N_45253);
xnor U49652 (N_49652,N_45474,N_45109);
xnor U49653 (N_49653,N_46347,N_45763);
nor U49654 (N_49654,N_47224,N_45624);
nor U49655 (N_49655,N_45248,N_46556);
nor U49656 (N_49656,N_45363,N_47076);
xor U49657 (N_49657,N_46153,N_45796);
nor U49658 (N_49658,N_45965,N_45507);
nand U49659 (N_49659,N_45930,N_45951);
nand U49660 (N_49660,N_45234,N_45860);
or U49661 (N_49661,N_46711,N_45026);
xnor U49662 (N_49662,N_47159,N_46005);
and U49663 (N_49663,N_45290,N_46233);
or U49664 (N_49664,N_45820,N_47156);
or U49665 (N_49665,N_46702,N_47362);
and U49666 (N_49666,N_46069,N_45255);
nor U49667 (N_49667,N_45350,N_46909);
nand U49668 (N_49668,N_46264,N_45307);
and U49669 (N_49669,N_47034,N_45305);
nand U49670 (N_49670,N_45687,N_47062);
or U49671 (N_49671,N_45226,N_47315);
nor U49672 (N_49672,N_47260,N_47368);
nand U49673 (N_49673,N_46118,N_45555);
or U49674 (N_49674,N_45946,N_47322);
or U49675 (N_49675,N_46003,N_45673);
or U49676 (N_49676,N_46378,N_47157);
nand U49677 (N_49677,N_46799,N_45590);
nor U49678 (N_49678,N_45386,N_46195);
and U49679 (N_49679,N_46444,N_46101);
nor U49680 (N_49680,N_45881,N_46001);
or U49681 (N_49681,N_46823,N_47345);
or U49682 (N_49682,N_45559,N_46755);
and U49683 (N_49683,N_46231,N_46125);
or U49684 (N_49684,N_46544,N_45139);
and U49685 (N_49685,N_46047,N_46288);
nand U49686 (N_49686,N_45581,N_47079);
xor U49687 (N_49687,N_46823,N_45142);
nand U49688 (N_49688,N_46984,N_46923);
nor U49689 (N_49689,N_45339,N_45593);
xor U49690 (N_49690,N_46602,N_46358);
xor U49691 (N_49691,N_47474,N_47188);
nor U49692 (N_49692,N_46119,N_46114);
nor U49693 (N_49693,N_45289,N_47049);
nand U49694 (N_49694,N_45638,N_46342);
xnor U49695 (N_49695,N_46582,N_46409);
and U49696 (N_49696,N_45597,N_46015);
nand U49697 (N_49697,N_46997,N_45458);
and U49698 (N_49698,N_45348,N_46175);
nand U49699 (N_49699,N_46373,N_46159);
xnor U49700 (N_49700,N_45871,N_45563);
nand U49701 (N_49701,N_45238,N_45630);
nand U49702 (N_49702,N_45083,N_46592);
or U49703 (N_49703,N_45595,N_47258);
nor U49704 (N_49704,N_46097,N_46356);
nand U49705 (N_49705,N_46630,N_46982);
or U49706 (N_49706,N_46578,N_46986);
nand U49707 (N_49707,N_45020,N_46626);
or U49708 (N_49708,N_46846,N_45984);
nor U49709 (N_49709,N_46466,N_45281);
xnor U49710 (N_49710,N_46217,N_45145);
and U49711 (N_49711,N_45286,N_46329);
xnor U49712 (N_49712,N_46035,N_46211);
nor U49713 (N_49713,N_45675,N_46412);
or U49714 (N_49714,N_46184,N_45737);
and U49715 (N_49715,N_46299,N_45735);
xnor U49716 (N_49716,N_46078,N_46914);
nor U49717 (N_49717,N_47268,N_46104);
or U49718 (N_49718,N_47474,N_45475);
nor U49719 (N_49719,N_47313,N_46005);
nand U49720 (N_49720,N_45436,N_46044);
nor U49721 (N_49721,N_45888,N_45095);
nand U49722 (N_49722,N_45280,N_46777);
xnor U49723 (N_49723,N_46013,N_46330);
nand U49724 (N_49724,N_47003,N_45523);
or U49725 (N_49725,N_47101,N_46016);
or U49726 (N_49726,N_45667,N_46870);
and U49727 (N_49727,N_45628,N_46959);
and U49728 (N_49728,N_45616,N_46601);
nand U49729 (N_49729,N_46940,N_46735);
and U49730 (N_49730,N_45240,N_46843);
or U49731 (N_49731,N_47270,N_46977);
nor U49732 (N_49732,N_46584,N_46885);
or U49733 (N_49733,N_45075,N_46377);
xnor U49734 (N_49734,N_46974,N_46713);
and U49735 (N_49735,N_47167,N_45979);
xnor U49736 (N_49736,N_46437,N_47467);
xor U49737 (N_49737,N_45776,N_46508);
and U49738 (N_49738,N_46002,N_46250);
nor U49739 (N_49739,N_46035,N_45852);
and U49740 (N_49740,N_45152,N_46584);
nand U49741 (N_49741,N_46916,N_47452);
and U49742 (N_49742,N_47107,N_46168);
and U49743 (N_49743,N_46673,N_46084);
and U49744 (N_49744,N_45573,N_47211);
nor U49745 (N_49745,N_45190,N_46919);
xnor U49746 (N_49746,N_46519,N_46566);
nor U49747 (N_49747,N_45986,N_46941);
or U49748 (N_49748,N_46832,N_45837);
xnor U49749 (N_49749,N_46179,N_45061);
nor U49750 (N_49750,N_46311,N_46263);
nand U49751 (N_49751,N_46590,N_46865);
or U49752 (N_49752,N_46252,N_46037);
nand U49753 (N_49753,N_47188,N_46688);
nand U49754 (N_49754,N_46566,N_46521);
nand U49755 (N_49755,N_45369,N_45005);
nand U49756 (N_49756,N_46031,N_45297);
nor U49757 (N_49757,N_45322,N_47360);
or U49758 (N_49758,N_47385,N_46971);
nand U49759 (N_49759,N_47461,N_46876);
xor U49760 (N_49760,N_47029,N_47007);
and U49761 (N_49761,N_47435,N_45864);
nor U49762 (N_49762,N_47407,N_46574);
nor U49763 (N_49763,N_45198,N_47053);
or U49764 (N_49764,N_45545,N_45942);
and U49765 (N_49765,N_47196,N_46679);
or U49766 (N_49766,N_46431,N_46868);
or U49767 (N_49767,N_46247,N_45609);
nand U49768 (N_49768,N_45009,N_46307);
xor U49769 (N_49769,N_45482,N_46491);
xor U49770 (N_49770,N_47397,N_47062);
and U49771 (N_49771,N_45020,N_45616);
or U49772 (N_49772,N_47128,N_47174);
xor U49773 (N_49773,N_46479,N_46858);
xor U49774 (N_49774,N_47417,N_45527);
and U49775 (N_49775,N_46480,N_46645);
and U49776 (N_49776,N_45472,N_47196);
or U49777 (N_49777,N_46577,N_45080);
nand U49778 (N_49778,N_45842,N_47101);
xnor U49779 (N_49779,N_47221,N_45500);
or U49780 (N_49780,N_45413,N_46037);
nor U49781 (N_49781,N_45526,N_47145);
and U49782 (N_49782,N_45403,N_45556);
or U49783 (N_49783,N_46060,N_45397);
nand U49784 (N_49784,N_46880,N_45331);
xnor U49785 (N_49785,N_47315,N_45718);
and U49786 (N_49786,N_46000,N_45436);
nor U49787 (N_49787,N_45182,N_46845);
or U49788 (N_49788,N_47082,N_46055);
nand U49789 (N_49789,N_47162,N_45719);
nor U49790 (N_49790,N_46759,N_45512);
nor U49791 (N_49791,N_47264,N_46289);
nand U49792 (N_49792,N_45103,N_45476);
or U49793 (N_49793,N_46791,N_46258);
and U49794 (N_49794,N_45526,N_46608);
xor U49795 (N_49795,N_45183,N_45928);
nor U49796 (N_49796,N_45372,N_45567);
xor U49797 (N_49797,N_47294,N_45976);
or U49798 (N_49798,N_45197,N_47488);
nor U49799 (N_49799,N_45225,N_46839);
or U49800 (N_49800,N_46313,N_46370);
nand U49801 (N_49801,N_45777,N_46351);
xnor U49802 (N_49802,N_46021,N_45991);
xor U49803 (N_49803,N_45311,N_47415);
and U49804 (N_49804,N_45340,N_47077);
xnor U49805 (N_49805,N_46658,N_45320);
xor U49806 (N_49806,N_46014,N_46304);
nand U49807 (N_49807,N_45120,N_46586);
xor U49808 (N_49808,N_46373,N_47240);
and U49809 (N_49809,N_46076,N_45573);
nor U49810 (N_49810,N_47210,N_45460);
and U49811 (N_49811,N_45133,N_46170);
xor U49812 (N_49812,N_45126,N_45684);
or U49813 (N_49813,N_46608,N_45291);
and U49814 (N_49814,N_47373,N_45592);
nand U49815 (N_49815,N_45620,N_47220);
nand U49816 (N_49816,N_47161,N_45706);
nand U49817 (N_49817,N_46171,N_46210);
nor U49818 (N_49818,N_46051,N_46999);
xor U49819 (N_49819,N_46918,N_46644);
nand U49820 (N_49820,N_45554,N_45473);
or U49821 (N_49821,N_45824,N_45496);
and U49822 (N_49822,N_46177,N_45430);
xnor U49823 (N_49823,N_45964,N_45793);
nand U49824 (N_49824,N_47050,N_46064);
nor U49825 (N_49825,N_45895,N_47217);
and U49826 (N_49826,N_46736,N_46648);
nor U49827 (N_49827,N_45208,N_46735);
or U49828 (N_49828,N_45046,N_45240);
nor U49829 (N_49829,N_45193,N_45413);
xnor U49830 (N_49830,N_46993,N_45630);
nor U49831 (N_49831,N_45102,N_45986);
or U49832 (N_49832,N_45171,N_45120);
xnor U49833 (N_49833,N_45401,N_45608);
nor U49834 (N_49834,N_46944,N_46163);
nor U49835 (N_49835,N_45146,N_47068);
or U49836 (N_49836,N_46302,N_46906);
or U49837 (N_49837,N_46943,N_46013);
xnor U49838 (N_49838,N_45176,N_46775);
xor U49839 (N_49839,N_45033,N_46247);
and U49840 (N_49840,N_47355,N_47132);
nand U49841 (N_49841,N_45527,N_45949);
or U49842 (N_49842,N_47080,N_45962);
or U49843 (N_49843,N_46369,N_46901);
and U49844 (N_49844,N_46405,N_47441);
and U49845 (N_49845,N_47261,N_46079);
or U49846 (N_49846,N_46186,N_45017);
nand U49847 (N_49847,N_45247,N_45048);
nand U49848 (N_49848,N_47149,N_45622);
nor U49849 (N_49849,N_45850,N_47281);
and U49850 (N_49850,N_45508,N_46029);
nor U49851 (N_49851,N_46600,N_45543);
xor U49852 (N_49852,N_45538,N_46274);
nor U49853 (N_49853,N_46242,N_47099);
xnor U49854 (N_49854,N_45725,N_46017);
nor U49855 (N_49855,N_46647,N_46698);
xor U49856 (N_49856,N_46002,N_45317);
xor U49857 (N_49857,N_47098,N_47355);
nor U49858 (N_49858,N_46011,N_46724);
nand U49859 (N_49859,N_46756,N_46100);
nand U49860 (N_49860,N_45926,N_46800);
nor U49861 (N_49861,N_46663,N_45103);
or U49862 (N_49862,N_46485,N_46130);
xor U49863 (N_49863,N_47364,N_47378);
nand U49864 (N_49864,N_47067,N_45887);
or U49865 (N_49865,N_45161,N_46475);
xor U49866 (N_49866,N_46222,N_45753);
and U49867 (N_49867,N_47302,N_46128);
or U49868 (N_49868,N_47447,N_45159);
or U49869 (N_49869,N_46302,N_45661);
nand U49870 (N_49870,N_47286,N_46652);
nor U49871 (N_49871,N_45392,N_45099);
xor U49872 (N_49872,N_47174,N_45736);
nor U49873 (N_49873,N_45007,N_45772);
or U49874 (N_49874,N_46314,N_46922);
xor U49875 (N_49875,N_46053,N_45081);
xnor U49876 (N_49876,N_45058,N_45214);
nand U49877 (N_49877,N_46698,N_45338);
and U49878 (N_49878,N_46080,N_46797);
nor U49879 (N_49879,N_45376,N_45326);
nand U49880 (N_49880,N_46399,N_47262);
nor U49881 (N_49881,N_45395,N_45051);
nor U49882 (N_49882,N_46647,N_46391);
nor U49883 (N_49883,N_45448,N_45018);
nor U49884 (N_49884,N_45782,N_46907);
nand U49885 (N_49885,N_46376,N_45661);
and U49886 (N_49886,N_47246,N_47013);
nand U49887 (N_49887,N_46193,N_45483);
or U49888 (N_49888,N_47112,N_47307);
nand U49889 (N_49889,N_45074,N_47459);
xor U49890 (N_49890,N_47334,N_45079);
or U49891 (N_49891,N_45107,N_45277);
or U49892 (N_49892,N_46482,N_46577);
and U49893 (N_49893,N_46267,N_46112);
xor U49894 (N_49894,N_45184,N_47497);
and U49895 (N_49895,N_46118,N_46451);
and U49896 (N_49896,N_45779,N_45427);
and U49897 (N_49897,N_45964,N_47492);
nand U49898 (N_49898,N_46569,N_45067);
nand U49899 (N_49899,N_46414,N_47204);
xor U49900 (N_49900,N_45617,N_45688);
nand U49901 (N_49901,N_45433,N_46318);
and U49902 (N_49902,N_45934,N_45585);
nand U49903 (N_49903,N_45482,N_45421);
nor U49904 (N_49904,N_45621,N_45106);
and U49905 (N_49905,N_45121,N_47141);
nor U49906 (N_49906,N_45705,N_46754);
and U49907 (N_49907,N_47436,N_46714);
xor U49908 (N_49908,N_47384,N_47472);
xor U49909 (N_49909,N_46688,N_47166);
nand U49910 (N_49910,N_46162,N_47406);
xnor U49911 (N_49911,N_46227,N_45520);
nor U49912 (N_49912,N_45815,N_47144);
xnor U49913 (N_49913,N_46852,N_46504);
or U49914 (N_49914,N_45989,N_46661);
nor U49915 (N_49915,N_45879,N_46157);
nand U49916 (N_49916,N_46294,N_45608);
or U49917 (N_49917,N_45998,N_46343);
xnor U49918 (N_49918,N_47198,N_45056);
and U49919 (N_49919,N_47359,N_45614);
and U49920 (N_49920,N_47223,N_45583);
and U49921 (N_49921,N_45315,N_46698);
or U49922 (N_49922,N_45279,N_45294);
nand U49923 (N_49923,N_45093,N_46263);
nand U49924 (N_49924,N_46277,N_46732);
or U49925 (N_49925,N_45695,N_46948);
and U49926 (N_49926,N_46080,N_46238);
and U49927 (N_49927,N_46348,N_46385);
and U49928 (N_49928,N_47188,N_45971);
and U49929 (N_49929,N_45884,N_46640);
nor U49930 (N_49930,N_46034,N_46136);
and U49931 (N_49931,N_46830,N_47034);
or U49932 (N_49932,N_46711,N_46255);
xnor U49933 (N_49933,N_45868,N_45091);
or U49934 (N_49934,N_45111,N_45601);
xor U49935 (N_49935,N_46235,N_46562);
or U49936 (N_49936,N_46372,N_45719);
and U49937 (N_49937,N_46915,N_45010);
nor U49938 (N_49938,N_46885,N_46120);
nand U49939 (N_49939,N_45308,N_46527);
nand U49940 (N_49940,N_47020,N_46739);
nor U49941 (N_49941,N_47012,N_45739);
or U49942 (N_49942,N_45883,N_45711);
xnor U49943 (N_49943,N_46319,N_47241);
and U49944 (N_49944,N_46600,N_46562);
xor U49945 (N_49945,N_45288,N_47454);
nand U49946 (N_49946,N_46096,N_47404);
nor U49947 (N_49947,N_47499,N_46834);
and U49948 (N_49948,N_45251,N_46394);
or U49949 (N_49949,N_46046,N_45954);
nand U49950 (N_49950,N_45521,N_46244);
nor U49951 (N_49951,N_47238,N_47115);
or U49952 (N_49952,N_45054,N_45494);
xnor U49953 (N_49953,N_45020,N_45017);
xnor U49954 (N_49954,N_45438,N_47289);
nand U49955 (N_49955,N_46847,N_46334);
or U49956 (N_49956,N_46164,N_47373);
and U49957 (N_49957,N_46356,N_46214);
and U49958 (N_49958,N_46525,N_45975);
nand U49959 (N_49959,N_45303,N_47435);
xor U49960 (N_49960,N_46426,N_45917);
or U49961 (N_49961,N_45395,N_46134);
nand U49962 (N_49962,N_45443,N_45616);
nor U49963 (N_49963,N_46715,N_46097);
nor U49964 (N_49964,N_47492,N_45789);
and U49965 (N_49965,N_45970,N_46889);
xnor U49966 (N_49966,N_45531,N_47370);
xnor U49967 (N_49967,N_45965,N_46600);
and U49968 (N_49968,N_46729,N_47201);
nand U49969 (N_49969,N_46173,N_46828);
xor U49970 (N_49970,N_47041,N_47236);
nor U49971 (N_49971,N_45529,N_46944);
and U49972 (N_49972,N_45767,N_47001);
nor U49973 (N_49973,N_46614,N_45007);
or U49974 (N_49974,N_47186,N_47037);
nand U49975 (N_49975,N_46930,N_46336);
nand U49976 (N_49976,N_45099,N_46378);
nand U49977 (N_49977,N_47178,N_45123);
xor U49978 (N_49978,N_45633,N_46789);
xnor U49979 (N_49979,N_45311,N_46017);
and U49980 (N_49980,N_45300,N_45088);
nor U49981 (N_49981,N_46772,N_45749);
xor U49982 (N_49982,N_47137,N_45831);
xor U49983 (N_49983,N_46000,N_47179);
xnor U49984 (N_49984,N_46599,N_46261);
nand U49985 (N_49985,N_46157,N_45751);
nand U49986 (N_49986,N_46516,N_46380);
nor U49987 (N_49987,N_45094,N_47301);
xnor U49988 (N_49988,N_46489,N_46605);
or U49989 (N_49989,N_46207,N_45444);
nand U49990 (N_49990,N_45788,N_46165);
xor U49991 (N_49991,N_45503,N_45387);
nand U49992 (N_49992,N_45166,N_46769);
nand U49993 (N_49993,N_47187,N_47233);
and U49994 (N_49994,N_45565,N_46705);
nor U49995 (N_49995,N_46474,N_46784);
or U49996 (N_49996,N_46203,N_45889);
xnor U49997 (N_49997,N_46293,N_47238);
and U49998 (N_49998,N_45921,N_45803);
xnor U49999 (N_49999,N_46085,N_46231);
or UO_0 (O_0,N_49984,N_49555);
and UO_1 (O_1,N_49276,N_47997);
nand UO_2 (O_2,N_48286,N_47527);
xor UO_3 (O_3,N_48779,N_49971);
nor UO_4 (O_4,N_48381,N_47649);
nor UO_5 (O_5,N_48697,N_49037);
and UO_6 (O_6,N_47838,N_47569);
and UO_7 (O_7,N_49892,N_49197);
xor UO_8 (O_8,N_48683,N_47913);
nor UO_9 (O_9,N_48056,N_48078);
or UO_10 (O_10,N_47664,N_48397);
or UO_11 (O_11,N_49383,N_48145);
nor UO_12 (O_12,N_48144,N_47658);
nand UO_13 (O_13,N_47804,N_48458);
and UO_14 (O_14,N_48642,N_47740);
or UO_15 (O_15,N_48103,N_48036);
nand UO_16 (O_16,N_48645,N_49160);
and UO_17 (O_17,N_49060,N_47937);
nor UO_18 (O_18,N_48090,N_48715);
and UO_19 (O_19,N_48535,N_48191);
or UO_20 (O_20,N_49649,N_48083);
nand UO_21 (O_21,N_49371,N_49139);
nand UO_22 (O_22,N_48364,N_48579);
xor UO_23 (O_23,N_49247,N_49263);
or UO_24 (O_24,N_49487,N_49043);
nand UO_25 (O_25,N_48825,N_48020);
nor UO_26 (O_26,N_49729,N_49851);
nor UO_27 (O_27,N_49423,N_48299);
and UO_28 (O_28,N_49047,N_47564);
or UO_29 (O_29,N_48565,N_47511);
or UO_30 (O_30,N_47853,N_49058);
and UO_31 (O_31,N_48962,N_49538);
nor UO_32 (O_32,N_48587,N_49733);
and UO_33 (O_33,N_48210,N_47858);
xor UO_34 (O_34,N_49335,N_48102);
nor UO_35 (O_35,N_49443,N_48313);
or UO_36 (O_36,N_47681,N_49355);
nand UO_37 (O_37,N_48816,N_48915);
or UO_38 (O_38,N_48624,N_47713);
or UO_39 (O_39,N_49142,N_48067);
nor UO_40 (O_40,N_49471,N_48784);
nor UO_41 (O_41,N_49833,N_49210);
or UO_42 (O_42,N_48076,N_47826);
xor UO_43 (O_43,N_49896,N_48731);
xor UO_44 (O_44,N_47991,N_49305);
nor UO_45 (O_45,N_49457,N_49241);
nor UO_46 (O_46,N_49343,N_48686);
and UO_47 (O_47,N_49393,N_48164);
and UO_48 (O_48,N_49169,N_48442);
nor UO_49 (O_49,N_48761,N_47809);
or UO_50 (O_50,N_49829,N_49111);
and UO_51 (O_51,N_48147,N_47662);
and UO_52 (O_52,N_48319,N_47956);
or UO_53 (O_53,N_49044,N_47595);
nor UO_54 (O_54,N_49859,N_47798);
nand UO_55 (O_55,N_49634,N_48220);
nor UO_56 (O_56,N_48457,N_47519);
nor UO_57 (O_57,N_48219,N_49313);
and UO_58 (O_58,N_47601,N_48189);
and UO_59 (O_59,N_49131,N_49563);
or UO_60 (O_60,N_49928,N_48358);
nand UO_61 (O_61,N_47539,N_48621);
or UO_62 (O_62,N_49166,N_48508);
or UO_63 (O_63,N_49041,N_48992);
nand UO_64 (O_64,N_49618,N_47786);
xnor UO_65 (O_65,N_49866,N_49446);
nor UO_66 (O_66,N_49352,N_47878);
nand UO_67 (O_67,N_49643,N_48729);
and UO_68 (O_68,N_48065,N_49795);
nand UO_69 (O_69,N_48157,N_49914);
and UO_70 (O_70,N_47758,N_48389);
xnor UO_71 (O_71,N_48833,N_48818);
xnor UO_72 (O_72,N_48328,N_48085);
or UO_73 (O_73,N_48096,N_49765);
and UO_74 (O_74,N_49891,N_47558);
nor UO_75 (O_75,N_48188,N_48351);
nor UO_76 (O_76,N_48541,N_48676);
or UO_77 (O_77,N_48080,N_47801);
nand UO_78 (O_78,N_48482,N_48785);
and UO_79 (O_79,N_47966,N_49644);
xor UO_80 (O_80,N_48139,N_48542);
nor UO_81 (O_81,N_48414,N_48835);
xor UO_82 (O_82,N_47950,N_48583);
or UO_83 (O_83,N_47825,N_49484);
xnor UO_84 (O_84,N_49285,N_48589);
nand UO_85 (O_85,N_47729,N_48943);
nand UO_86 (O_86,N_48710,N_49607);
xor UO_87 (O_87,N_48502,N_49089);
and UO_88 (O_88,N_49817,N_49615);
nand UO_89 (O_89,N_47744,N_49126);
xor UO_90 (O_90,N_49539,N_48557);
xnor UO_91 (O_91,N_48994,N_48465);
xor UO_92 (O_92,N_49536,N_49448);
nor UO_93 (O_93,N_49753,N_49147);
or UO_94 (O_94,N_48913,N_48936);
or UO_95 (O_95,N_47995,N_49202);
and UO_96 (O_96,N_49402,N_49939);
or UO_97 (O_97,N_48371,N_48734);
xor UO_98 (O_98,N_49229,N_48180);
or UO_99 (O_99,N_48045,N_48217);
xnor UO_100 (O_100,N_48593,N_48807);
nand UO_101 (O_101,N_48384,N_49045);
xnor UO_102 (O_102,N_49901,N_49898);
xnor UO_103 (O_103,N_48488,N_48503);
xnor UO_104 (O_104,N_49717,N_49049);
nand UO_105 (O_105,N_49001,N_49323);
and UO_106 (O_106,N_48114,N_49957);
or UO_107 (O_107,N_48478,N_48127);
or UO_108 (O_108,N_48044,N_49426);
xnor UO_109 (O_109,N_48107,N_49944);
nor UO_110 (O_110,N_48911,N_49161);
and UO_111 (O_111,N_48693,N_47520);
nor UO_112 (O_112,N_48563,N_49728);
or UO_113 (O_113,N_48453,N_48237);
or UO_114 (O_114,N_47749,N_48880);
xor UO_115 (O_115,N_49521,N_47582);
and UO_116 (O_116,N_49057,N_48499);
or UO_117 (O_117,N_48647,N_48674);
nor UO_118 (O_118,N_49766,N_48918);
and UO_119 (O_119,N_49587,N_47884);
nand UO_120 (O_120,N_49938,N_48916);
or UO_121 (O_121,N_48419,N_48576);
nor UO_122 (O_122,N_49430,N_49948);
xnor UO_123 (O_123,N_48662,N_49080);
nor UO_124 (O_124,N_48428,N_48211);
nand UO_125 (O_125,N_49260,N_47725);
nand UO_126 (O_126,N_49257,N_47665);
or UO_127 (O_127,N_48652,N_48775);
or UO_128 (O_128,N_48518,N_48166);
or UO_129 (O_129,N_48324,N_48948);
xor UO_130 (O_130,N_49746,N_48336);
xor UO_131 (O_131,N_48214,N_49351);
or UO_132 (O_132,N_49081,N_48346);
or UO_133 (O_133,N_49922,N_49992);
and UO_134 (O_134,N_49790,N_48207);
and UO_135 (O_135,N_47975,N_48505);
nand UO_136 (O_136,N_47574,N_48736);
nand UO_137 (O_137,N_48363,N_47597);
and UO_138 (O_138,N_48746,N_48345);
and UO_139 (O_139,N_48228,N_48239);
nor UO_140 (O_140,N_48374,N_49379);
nor UO_141 (O_141,N_49706,N_47863);
xnor UO_142 (O_142,N_48754,N_48288);
nor UO_143 (O_143,N_48269,N_49592);
nor UO_144 (O_144,N_49022,N_48532);
xnor UO_145 (O_145,N_48264,N_48623);
nand UO_146 (O_146,N_48848,N_49700);
and UO_147 (O_147,N_47695,N_49871);
and UO_148 (O_148,N_48495,N_49814);
xnor UO_149 (O_149,N_48860,N_49972);
and UO_150 (O_150,N_49449,N_48243);
or UO_151 (O_151,N_48974,N_48395);
nor UO_152 (O_152,N_49902,N_49658);
xor UO_153 (O_153,N_49911,N_49533);
and UO_154 (O_154,N_48278,N_48799);
and UO_155 (O_155,N_47773,N_47948);
xnor UO_156 (O_156,N_47981,N_48872);
and UO_157 (O_157,N_48119,N_47578);
nand UO_158 (O_158,N_48850,N_48163);
or UO_159 (O_159,N_49495,N_49621);
nand UO_160 (O_160,N_48942,N_47745);
or UO_161 (O_161,N_48536,N_48577);
and UO_162 (O_162,N_47557,N_48882);
nand UO_163 (O_163,N_48982,N_47766);
nor UO_164 (O_164,N_49480,N_47603);
xnor UO_165 (O_165,N_49013,N_49106);
nand UO_166 (O_166,N_48155,N_48633);
nand UO_167 (O_167,N_49603,N_49976);
nor UO_168 (O_168,N_49693,N_48957);
nand UO_169 (O_169,N_48034,N_49418);
xnor UO_170 (O_170,N_49178,N_48466);
nand UO_171 (O_171,N_49571,N_47893);
and UO_172 (O_172,N_47661,N_49110);
or UO_173 (O_173,N_49826,N_49339);
nor UO_174 (O_174,N_48028,N_49574);
nand UO_175 (O_175,N_48740,N_49815);
nor UO_176 (O_176,N_48087,N_48448);
or UO_177 (O_177,N_49230,N_48252);
xor UO_178 (O_178,N_47521,N_48332);
xor UO_179 (O_179,N_49368,N_47886);
nor UO_180 (O_180,N_49900,N_48824);
nand UO_181 (O_181,N_47528,N_49332);
or UO_182 (O_182,N_49946,N_47618);
xor UO_183 (O_183,N_49656,N_48856);
and UO_184 (O_184,N_48149,N_48826);
xor UO_185 (O_185,N_47824,N_47954);
nor UO_186 (O_186,N_49887,N_48912);
xor UO_187 (O_187,N_49774,N_49975);
nand UO_188 (O_188,N_48434,N_49283);
nor UO_189 (O_189,N_49016,N_48801);
xnor UO_190 (O_190,N_47555,N_49444);
and UO_191 (O_191,N_49879,N_49595);
nor UO_192 (O_192,N_49077,N_48010);
and UO_193 (O_193,N_48898,N_47828);
or UO_194 (O_194,N_47978,N_47812);
nand UO_195 (O_195,N_48658,N_47694);
xnor UO_196 (O_196,N_49399,N_48939);
and UO_197 (O_197,N_49440,N_49143);
xor UO_198 (O_198,N_48981,N_49736);
xnor UO_199 (O_199,N_47711,N_47994);
and UO_200 (O_200,N_48176,N_48098);
xor UO_201 (O_201,N_49954,N_48889);
nand UO_202 (O_202,N_47670,N_49251);
nand UO_203 (O_203,N_49123,N_47945);
or UO_204 (O_204,N_47959,N_48081);
nand UO_205 (O_205,N_49342,N_49793);
or UO_206 (O_206,N_48354,N_49085);
xor UO_207 (O_207,N_47748,N_48628);
and UO_208 (O_208,N_48070,N_48162);
nor UO_209 (O_209,N_49861,N_48097);
xnor UO_210 (O_210,N_47967,N_47614);
and UO_211 (O_211,N_48935,N_48021);
and UO_212 (O_212,N_48758,N_48698);
nor UO_213 (O_213,N_48320,N_49782);
nand UO_214 (O_214,N_47859,N_49541);
or UO_215 (O_215,N_47602,N_49918);
nor UO_216 (O_216,N_48330,N_49692);
xor UO_217 (O_217,N_49345,N_49747);
and UO_218 (O_218,N_48594,N_47721);
nand UO_219 (O_219,N_48701,N_49549);
nand UO_220 (O_220,N_49006,N_49750);
nand UO_221 (O_221,N_47999,N_49577);
xnor UO_222 (O_222,N_48572,N_49562);
and UO_223 (O_223,N_47874,N_47588);
or UO_224 (O_224,N_48222,N_47780);
nor UO_225 (O_225,N_47844,N_49771);
and UO_226 (O_226,N_47833,N_49791);
or UO_227 (O_227,N_48225,N_48111);
nor UO_228 (O_228,N_49101,N_49565);
or UO_229 (O_229,N_47599,N_49714);
xnor UO_230 (O_230,N_47964,N_48894);
xnor UO_231 (O_231,N_49792,N_48735);
and UO_232 (O_232,N_49364,N_49788);
or UO_233 (O_233,N_49120,N_49174);
nor UO_234 (O_234,N_48648,N_48321);
nor UO_235 (O_235,N_48513,N_48302);
nor UO_236 (O_236,N_49214,N_48161);
xor UO_237 (O_237,N_48312,N_47732);
xnor UO_238 (O_238,N_47613,N_48040);
nand UO_239 (O_239,N_48560,N_47860);
and UO_240 (O_240,N_49801,N_48684);
xor UO_241 (O_241,N_49201,N_48411);
xnor UO_242 (O_242,N_49773,N_48368);
xor UO_243 (O_243,N_49119,N_48362);
nor UO_244 (O_244,N_49828,N_49893);
nor UO_245 (O_245,N_49684,N_47915);
nand UO_246 (O_246,N_48811,N_49924);
and UO_247 (O_247,N_48712,N_49410);
xor UO_248 (O_248,N_48875,N_47516);
and UO_249 (O_249,N_49518,N_47709);
or UO_250 (O_250,N_48013,N_47728);
xor UO_251 (O_251,N_47633,N_49496);
nor UO_252 (O_252,N_47655,N_49913);
and UO_253 (O_253,N_48803,N_47517);
and UO_254 (O_254,N_48634,N_49752);
xnor UO_255 (O_255,N_48071,N_48050);
or UO_256 (O_256,N_49504,N_48605);
and UO_257 (O_257,N_47883,N_49292);
or UO_258 (O_258,N_47796,N_49104);
or UO_259 (O_259,N_49000,N_48005);
and UO_260 (O_260,N_49376,N_48906);
nor UO_261 (O_261,N_47581,N_49370);
nand UO_262 (O_262,N_49824,N_48530);
and UO_263 (O_263,N_47876,N_48063);
and UO_264 (O_264,N_47741,N_48075);
xor UO_265 (O_265,N_48062,N_48789);
nand UO_266 (O_266,N_48487,N_47522);
nor UO_267 (O_267,N_49551,N_47787);
and UO_268 (O_268,N_47503,N_49648);
or UO_269 (O_269,N_49378,N_47577);
or UO_270 (O_270,N_47546,N_49545);
nor UO_271 (O_271,N_48490,N_48893);
xor UO_272 (O_272,N_47856,N_47944);
nand UO_273 (O_273,N_49525,N_47841);
nand UO_274 (O_274,N_49149,N_49597);
xnor UO_275 (O_275,N_47534,N_49917);
nor UO_276 (O_276,N_47712,N_47628);
or UO_277 (O_277,N_47963,N_49438);
nand UO_278 (O_278,N_49391,N_48522);
nor UO_279 (O_279,N_48598,N_47862);
nand UO_280 (O_280,N_48099,N_48471);
xnor UO_281 (O_281,N_48204,N_48938);
nor UO_282 (O_282,N_47585,N_49605);
nand UO_283 (O_283,N_49989,N_47553);
or UO_284 (O_284,N_48196,N_48223);
or UO_285 (O_285,N_48273,N_48178);
nor UO_286 (O_286,N_47783,N_48823);
and UO_287 (O_287,N_48526,N_49838);
or UO_288 (O_288,N_48254,N_47829);
nand UO_289 (O_289,N_47652,N_49482);
xor UO_290 (O_290,N_48925,N_48743);
nand UO_291 (O_291,N_48260,N_49811);
nand UO_292 (O_292,N_47907,N_48118);
or UO_293 (O_293,N_49213,N_49731);
nor UO_294 (O_294,N_48291,N_48245);
xor UO_295 (O_295,N_49337,N_47523);
and UO_296 (O_296,N_49183,N_49857);
and UO_297 (O_297,N_48016,N_48705);
and UO_298 (O_298,N_49424,N_48617);
xnor UO_299 (O_299,N_48786,N_48361);
and UO_300 (O_300,N_48827,N_48854);
nand UO_301 (O_301,N_48186,N_47998);
and UO_302 (O_302,N_48048,N_49405);
nand UO_303 (O_303,N_48311,N_48283);
xnor UO_304 (O_304,N_48940,N_48622);
and UO_305 (O_305,N_49455,N_49350);
and UO_306 (O_306,N_47639,N_48285);
or UO_307 (O_307,N_47717,N_49458);
xor UO_308 (O_308,N_48060,N_49211);
nor UO_309 (O_309,N_48663,N_49320);
or UO_310 (O_310,N_47634,N_47918);
nor UO_311 (O_311,N_49606,N_49754);
and UO_312 (O_312,N_49236,N_47762);
xnor UO_313 (O_313,N_49679,N_49435);
nand UO_314 (O_314,N_49636,N_48639);
xor UO_315 (O_315,N_48665,N_48383);
and UO_316 (O_316,N_48999,N_48206);
xnor UO_317 (O_317,N_48776,N_49908);
and UO_318 (O_318,N_49818,N_47596);
nand UO_319 (O_319,N_47903,N_49493);
nand UO_320 (O_320,N_49189,N_49272);
or UO_321 (O_321,N_49459,N_48529);
nand UO_322 (O_322,N_48768,N_48976);
or UO_323 (O_323,N_47568,N_49329);
nor UO_324 (O_324,N_49987,N_47632);
and UO_325 (O_325,N_49751,N_48104);
xor UO_326 (O_326,N_48258,N_47604);
and UO_327 (O_327,N_49532,N_49406);
and UO_328 (O_328,N_49516,N_49702);
and UO_329 (O_329,N_48279,N_47822);
nor UO_330 (O_330,N_47743,N_48304);
nor UO_331 (O_331,N_49570,N_48849);
nor UO_332 (O_332,N_49115,N_48914);
or UO_333 (O_333,N_49947,N_49601);
or UO_334 (O_334,N_48426,N_49414);
xor UO_335 (O_335,N_48408,N_49377);
and UO_336 (O_336,N_47923,N_49204);
nor UO_337 (O_337,N_48969,N_48989);
or UO_338 (O_338,N_47646,N_48130);
nand UO_339 (O_339,N_48035,N_49567);
nand UO_340 (O_340,N_48027,N_48963);
nand UO_341 (O_341,N_49387,N_47714);
nor UO_342 (O_342,N_47679,N_48991);
xor UO_343 (O_343,N_47789,N_49289);
xor UO_344 (O_344,N_49328,N_48317);
xnor UO_345 (O_345,N_47751,N_49870);
and UO_346 (O_346,N_48718,N_48524);
nor UO_347 (O_347,N_48699,N_49167);
xnor UO_348 (O_348,N_48025,N_49083);
or UO_349 (O_349,N_48570,N_49672);
nor UO_350 (O_350,N_47960,N_49097);
nor UO_351 (O_351,N_49324,N_49281);
or UO_352 (O_352,N_48432,N_48853);
or UO_353 (O_353,N_47880,N_47622);
nand UO_354 (O_354,N_48390,N_48986);
xnor UO_355 (O_355,N_49358,N_49677);
or UO_356 (O_356,N_49515,N_47754);
xor UO_357 (O_357,N_49572,N_49112);
or UO_358 (O_358,N_49962,N_49347);
nand UO_359 (O_359,N_48858,N_48772);
or UO_360 (O_360,N_49187,N_49712);
or UO_361 (O_361,N_48476,N_49895);
xnor UO_362 (O_362,N_49019,N_48667);
xnor UO_363 (O_363,N_48838,N_49092);
nand UO_364 (O_364,N_49716,N_49524);
and UO_365 (O_365,N_47708,N_49267);
or UO_366 (O_366,N_48376,N_48660);
and UO_367 (O_367,N_49326,N_48216);
nand UO_368 (O_368,N_48190,N_47691);
and UO_369 (O_369,N_49107,N_48391);
or UO_370 (O_370,N_49874,N_48564);
xnor UO_371 (O_371,N_48468,N_47624);
nand UO_372 (O_372,N_48402,N_48531);
and UO_373 (O_373,N_49735,N_49794);
or UO_374 (O_374,N_49769,N_49640);
and UO_375 (O_375,N_49958,N_49067);
nor UO_376 (O_376,N_48533,N_48668);
nor UO_377 (O_377,N_47818,N_49207);
or UO_378 (O_378,N_49689,N_49033);
nand UO_379 (O_379,N_48301,N_48296);
nand UO_380 (O_380,N_49611,N_49599);
or UO_381 (O_381,N_47502,N_48356);
nand UO_382 (O_382,N_49638,N_49614);
and UO_383 (O_383,N_47974,N_49641);
nand UO_384 (O_384,N_48763,N_47638);
xor UO_385 (O_385,N_48094,N_49153);
and UO_386 (O_386,N_49840,N_48777);
or UO_387 (O_387,N_49973,N_47952);
nor UO_388 (O_388,N_48585,N_48122);
nand UO_389 (O_389,N_47570,N_49150);
and UO_390 (O_390,N_49651,N_48923);
nand UO_391 (O_391,N_49666,N_49812);
and UO_392 (O_392,N_49743,N_49450);
or UO_393 (O_393,N_48657,N_48810);
or UO_394 (O_394,N_49505,N_48770);
nor UO_395 (O_395,N_47561,N_48360);
or UO_396 (O_396,N_48884,N_47794);
xnor UO_397 (O_397,N_49528,N_47678);
xor UO_398 (O_398,N_48876,N_49098);
and UO_399 (O_399,N_48271,N_49141);
xnor UO_400 (O_400,N_48151,N_49985);
nor UO_401 (O_401,N_49763,N_49960);
nand UO_402 (O_402,N_48394,N_48904);
nor UO_403 (O_403,N_48650,N_48444);
or UO_404 (O_404,N_49367,N_49108);
xnor UO_405 (O_405,N_47811,N_49452);
nand UO_406 (O_406,N_48109,N_48504);
xnor UO_407 (O_407,N_48227,N_49382);
nand UO_408 (O_408,N_48695,N_48694);
or UO_409 (O_409,N_49779,N_48604);
nand UO_410 (O_410,N_49520,N_47535);
nand UO_411 (O_411,N_48903,N_49749);
nand UO_412 (O_412,N_49195,N_49265);
and UO_413 (O_413,N_49600,N_49270);
and UO_414 (O_414,N_48303,N_49858);
xnor UO_415 (O_415,N_47830,N_48485);
nand UO_416 (O_416,N_49102,N_49075);
xnor UO_417 (O_417,N_48003,N_48350);
nand UO_418 (O_418,N_47879,N_49021);
or UO_419 (O_419,N_49159,N_49864);
or UO_420 (O_420,N_48741,N_48492);
xor UO_421 (O_421,N_49894,N_47593);
and UO_422 (O_422,N_48512,N_49821);
or UO_423 (O_423,N_47854,N_47898);
nand UO_424 (O_424,N_49274,N_49760);
nor UO_425 (O_425,N_48287,N_48413);
or UO_426 (O_426,N_49277,N_48846);
xor UO_427 (O_427,N_48209,N_48802);
or UO_428 (O_428,N_49401,N_49783);
and UO_429 (O_429,N_49498,N_49865);
xor UO_430 (O_430,N_48061,N_49409);
nand UO_431 (O_431,N_49117,N_48716);
or UO_432 (O_432,N_47836,N_49034);
nor UO_433 (O_433,N_48797,N_49095);
xnor UO_434 (O_434,N_49062,N_47788);
nor UO_435 (O_435,N_48297,N_48486);
nand UO_436 (O_436,N_49403,N_49961);
nand UO_437 (O_437,N_47567,N_48259);
or UO_438 (O_438,N_49990,N_49099);
nand UO_439 (O_439,N_49420,N_48412);
and UO_440 (O_440,N_49154,N_48150);
xor UO_441 (O_441,N_48129,N_48813);
xnor UO_442 (O_442,N_48138,N_47888);
or UO_443 (O_443,N_49832,N_47641);
and UO_444 (O_444,N_49408,N_48165);
xnor UO_445 (O_445,N_49696,N_47625);
or UO_446 (O_446,N_48121,N_47774);
nand UO_447 (O_447,N_49912,N_48724);
xor UO_448 (O_448,N_48202,N_48433);
nor UO_449 (O_449,N_48256,N_49278);
and UO_450 (O_450,N_47935,N_49909);
nor UO_451 (O_451,N_47510,N_49015);
nor UO_452 (O_452,N_49988,N_48774);
or UO_453 (O_453,N_48367,N_47757);
and UO_454 (O_454,N_47839,N_48461);
nand UO_455 (O_455,N_49040,N_48954);
nand UO_456 (O_456,N_48197,N_49312);
nand UO_457 (O_457,N_47654,N_49008);
nor UO_458 (O_458,N_49129,N_49823);
xor UO_459 (O_459,N_48452,N_47616);
nand UO_460 (O_460,N_48753,N_48066);
or UO_461 (O_461,N_48215,N_48318);
and UO_462 (O_462,N_49705,N_48704);
xnor UO_463 (O_463,N_49314,N_47889);
and UO_464 (O_464,N_48342,N_48403);
xnor UO_465 (O_465,N_48174,N_49558);
xor UO_466 (O_466,N_47778,N_47768);
nand UO_467 (O_467,N_48136,N_49544);
or UO_468 (O_468,N_47610,N_47667);
xor UO_469 (O_469,N_48043,N_49398);
nand UO_470 (O_470,N_48095,N_49428);
or UO_471 (O_471,N_49472,N_49168);
nor UO_472 (O_472,N_47608,N_49134);
nand UO_473 (O_473,N_49179,N_47537);
nand UO_474 (O_474,N_48140,N_49223);
nand UO_475 (O_475,N_49464,N_49439);
and UO_476 (O_476,N_49124,N_48156);
and UO_477 (O_477,N_48038,N_48000);
or UO_478 (O_478,N_49585,N_48229);
or UO_479 (O_479,N_49660,N_48806);
xnor UO_480 (O_480,N_49434,N_48110);
nand UO_481 (O_481,N_49886,N_48711);
or UO_482 (O_482,N_49392,N_47814);
xor UO_483 (O_483,N_49127,N_49056);
nand UO_484 (O_484,N_49216,N_48241);
nor UO_485 (O_485,N_49968,N_47989);
xnor UO_486 (O_486,N_48883,N_48331);
nand UO_487 (O_487,N_48298,N_48322);
nor UO_488 (O_488,N_47756,N_47802);
or UO_489 (O_489,N_48475,N_47929);
and UO_490 (O_490,N_49456,N_48544);
xnor UO_491 (O_491,N_47598,N_49629);
nand UO_492 (O_492,N_49842,N_47620);
nand UO_493 (O_493,N_49431,N_49224);
and UO_494 (O_494,N_49386,N_47781);
and UO_495 (O_495,N_48771,N_47590);
nand UO_496 (O_496,N_49986,N_49237);
nand UO_497 (O_497,N_48396,N_48105);
nor UO_498 (O_498,N_47547,N_47734);
or UO_499 (O_499,N_48902,N_49275);
or UO_500 (O_500,N_48750,N_48985);
nand UO_501 (O_501,N_49557,N_47771);
or UO_502 (O_502,N_49994,N_48423);
or UO_503 (O_503,N_49310,N_47600);
and UO_504 (O_504,N_49125,N_49959);
xor UO_505 (O_505,N_48429,N_49949);
and UO_506 (O_506,N_49385,N_48032);
or UO_507 (O_507,N_48891,N_49843);
nor UO_508 (O_508,N_47843,N_48756);
nor UO_509 (O_509,N_47936,N_48401);
and UO_510 (O_510,N_48146,N_48863);
or UO_511 (O_511,N_48548,N_48757);
or UO_512 (O_512,N_48172,N_47776);
or UO_513 (O_513,N_47563,N_48713);
or UO_514 (O_514,N_48115,N_49186);
nor UO_515 (O_515,N_48696,N_49800);
or UO_516 (O_516,N_48327,N_49720);
xor UO_517 (O_517,N_48919,N_49280);
nand UO_518 (O_518,N_47850,N_49020);
xor UO_519 (O_519,N_47791,N_48934);
and UO_520 (O_520,N_49616,N_48051);
nand UO_521 (O_521,N_49718,N_47919);
or UO_522 (O_522,N_49724,N_48603);
nand UO_523 (O_523,N_48359,N_49009);
nor UO_524 (O_524,N_48673,N_48520);
nor UO_525 (O_525,N_49703,N_48759);
nand UO_526 (O_526,N_48998,N_48479);
and UO_527 (O_527,N_47770,N_48755);
and UO_528 (O_528,N_47980,N_49789);
nor UO_529 (O_529,N_49388,N_49357);
nor UO_530 (O_530,N_49834,N_48276);
and UO_531 (O_531,N_48248,N_48555);
xor UO_532 (O_532,N_48525,N_48865);
nand UO_533 (O_533,N_48068,N_49268);
xor UO_534 (O_534,N_48128,N_49316);
or UO_535 (O_535,N_48480,N_48744);
nand UO_536 (O_536,N_47934,N_48501);
or UO_537 (O_537,N_48947,N_48878);
nor UO_538 (O_538,N_48131,N_49514);
and UO_539 (O_539,N_48385,N_47914);
nor UO_540 (O_540,N_47892,N_48946);
xnor UO_541 (O_541,N_47571,N_48590);
nor UO_542 (O_542,N_47851,N_47540);
nand UO_543 (O_543,N_49770,N_48218);
xor UO_544 (O_544,N_47746,N_49797);
or UO_545 (O_545,N_49955,N_48325);
xor UO_546 (O_546,N_49850,N_49715);
xor UO_547 (O_547,N_48778,N_48404);
xor UO_548 (O_548,N_47607,N_49476);
xnor UO_549 (O_549,N_47609,N_49273);
nor UO_550 (O_550,N_49590,N_48496);
nand UO_551 (O_551,N_48928,N_49433);
and UO_552 (O_552,N_49950,N_48773);
nor UO_553 (O_553,N_48443,N_49185);
nand UO_554 (O_554,N_49205,N_48326);
and UO_555 (O_555,N_49144,N_48931);
or UO_556 (O_556,N_49148,N_48769);
or UO_557 (O_557,N_48945,N_49921);
and UO_558 (O_558,N_49934,N_49293);
nand UO_559 (O_559,N_48233,N_47782);
and UO_560 (O_560,N_49772,N_49240);
and UO_561 (O_561,N_49635,N_49485);
nand UO_562 (O_562,N_48275,N_49624);
or UO_563 (O_563,N_49050,N_48881);
and UO_564 (O_564,N_49014,N_48493);
or UO_565 (O_565,N_47763,N_47861);
or UO_566 (O_566,N_47635,N_49301);
xor UO_567 (O_567,N_48474,N_49191);
nand UO_568 (O_568,N_49980,N_48108);
nor UO_569 (O_569,N_49356,N_49182);
or UO_570 (O_570,N_47846,N_49319);
or UO_571 (O_571,N_49349,N_49506);
nor UO_572 (O_572,N_47940,N_48049);
nand UO_573 (O_573,N_48091,N_48595);
xnor UO_574 (O_574,N_49995,N_47693);
and UO_575 (O_575,N_49053,N_48093);
and UO_576 (O_576,N_47752,N_49489);
nor UO_577 (O_577,N_48896,N_48047);
or UO_578 (O_578,N_49175,N_49055);
xor UO_579 (O_579,N_47808,N_48236);
and UO_580 (O_580,N_48077,N_49023);
xnor UO_581 (O_581,N_47925,N_49740);
xor UO_582 (O_582,N_48026,N_47819);
xnor UO_583 (O_583,N_49164,N_48888);
and UO_584 (O_584,N_49334,N_48588);
and UO_585 (O_585,N_49907,N_49529);
and UO_586 (O_586,N_48017,N_48762);
nand UO_587 (O_587,N_48447,N_48057);
or UO_588 (O_588,N_49395,N_48392);
and UO_589 (O_589,N_47984,N_49613);
nor UO_590 (O_590,N_47848,N_49425);
nor UO_591 (O_591,N_49193,N_49628);
or UO_592 (O_592,N_48831,N_49777);
nand UO_593 (O_593,N_49196,N_47986);
or UO_594 (O_594,N_49136,N_49664);
or UO_595 (O_595,N_49076,N_49872);
and UO_596 (O_596,N_49114,N_47718);
or UO_597 (O_597,N_49018,N_48721);
or UO_598 (O_598,N_49087,N_47958);
or UO_599 (O_599,N_48305,N_48250);
and UO_600 (O_600,N_49121,N_47515);
nor UO_601 (O_601,N_47891,N_49404);
and UO_602 (O_602,N_49589,N_49593);
and UO_603 (O_603,N_47663,N_49776);
nand UO_604 (O_604,N_47761,N_47894);
xor UO_605 (O_605,N_49315,N_49340);
nand UO_606 (O_606,N_48380,N_48723);
nand UO_607 (O_607,N_48470,N_49344);
and UO_608 (O_608,N_48960,N_48314);
nand UO_609 (O_609,N_47920,N_49447);
xor UO_610 (O_610,N_47855,N_48601);
nand UO_611 (O_611,N_49372,N_48289);
nand UO_612 (O_612,N_48861,N_49966);
nor UO_613 (O_613,N_48725,N_48169);
or UO_614 (O_614,N_48978,N_48899);
nand UO_615 (O_615,N_49012,N_48867);
and UO_616 (O_616,N_49155,N_48293);
nand UO_617 (O_617,N_48733,N_48440);
xnor UO_618 (O_618,N_49991,N_47526);
and UO_619 (O_619,N_49234,N_48656);
nand UO_620 (O_620,N_48739,N_48160);
xnor UO_621 (O_621,N_47985,N_49209);
nand UO_622 (O_622,N_48975,N_49899);
or UO_623 (O_623,N_48708,N_49503);
and UO_624 (O_624,N_49116,N_47881);
or UO_625 (O_625,N_48814,N_48494);
or UO_626 (O_626,N_48126,N_47704);
or UO_627 (O_627,N_48793,N_49630);
xnor UO_628 (O_628,N_49437,N_47753);
nor UO_629 (O_629,N_49411,N_48545);
xor UO_630 (O_630,N_48373,N_49497);
nor UO_631 (O_631,N_47943,N_49145);
xnor UO_632 (O_632,N_47733,N_48234);
xor UO_633 (O_633,N_47672,N_48251);
nand UO_634 (O_634,N_48459,N_49584);
and UO_635 (O_635,N_48240,N_49983);
xor UO_636 (O_636,N_48840,N_49381);
or UO_637 (O_637,N_48053,N_47559);
and UO_638 (O_638,N_48445,N_47518);
nor UO_639 (O_639,N_48566,N_48199);
and UO_640 (O_640,N_49302,N_47816);
nor UO_641 (O_641,N_47852,N_49744);
and UO_642 (O_642,N_48788,N_48968);
nor UO_643 (O_643,N_48600,N_49923);
or UO_644 (O_644,N_48198,N_49527);
or UO_645 (O_645,N_49248,N_49937);
nand UO_646 (O_646,N_47764,N_49739);
xnor UO_647 (O_647,N_48158,N_48805);
or UO_648 (O_648,N_49194,N_48266);
nand UO_649 (O_649,N_48430,N_49903);
or UO_650 (O_650,N_48926,N_49830);
nand UO_651 (O_651,N_47805,N_48714);
nor UO_652 (O_652,N_48052,N_49502);
xnor UO_653 (O_653,N_49890,N_49678);
and UO_654 (O_654,N_49192,N_48438);
nand UO_655 (O_655,N_49930,N_47700);
or UO_656 (O_656,N_47742,N_49231);
and UO_657 (O_657,N_47899,N_48661);
nand UO_658 (O_658,N_47867,N_48339);
nor UO_659 (O_659,N_49336,N_48348);
and UO_660 (O_660,N_47636,N_47686);
xor UO_661 (O_661,N_48558,N_49091);
xor UO_662 (O_662,N_49981,N_48842);
or UO_663 (O_663,N_48135,N_47703);
or UO_664 (O_664,N_48582,N_49856);
xor UO_665 (O_665,N_47775,N_48004);
or UO_666 (O_666,N_49701,N_49885);
or UO_667 (O_667,N_47823,N_49697);
xor UO_668 (O_668,N_47910,N_48574);
xor UO_669 (O_669,N_47730,N_48349);
or UO_670 (O_670,N_48001,N_48124);
or UO_671 (O_671,N_48787,N_49461);
and UO_672 (O_672,N_48455,N_49441);
and UO_673 (O_673,N_48484,N_47807);
or UO_674 (O_674,N_49509,N_48751);
xor UO_675 (O_675,N_49798,N_48864);
nor UO_676 (O_676,N_48651,N_49470);
and UO_677 (O_677,N_49477,N_49925);
nand UO_678 (O_678,N_49531,N_49079);
or UO_679 (O_679,N_49876,N_48892);
and UO_680 (O_680,N_47500,N_48516);
nor UO_681 (O_681,N_49667,N_47611);
or UO_682 (O_682,N_47922,N_48602);
nand UO_683 (O_683,N_49366,N_49492);
and UO_684 (O_684,N_49413,N_49940);
nand UO_685 (O_685,N_48082,N_48990);
and UO_686 (O_686,N_48142,N_49764);
nand UO_687 (O_687,N_47750,N_48632);
nor UO_688 (O_688,N_49952,N_48571);
or UO_689 (O_689,N_47890,N_48113);
xor UO_690 (O_690,N_49035,N_48591);
or UO_691 (O_691,N_49627,N_49369);
nand UO_692 (O_692,N_48290,N_49999);
xnor UO_693 (O_693,N_49810,N_48599);
or UO_694 (O_694,N_48552,N_48927);
nor UO_695 (O_695,N_48631,N_47584);
and UO_696 (O_696,N_49296,N_49942);
nand UO_697 (O_697,N_49258,N_48979);
nand UO_698 (O_698,N_49052,N_49246);
nand UO_699 (O_699,N_47953,N_47533);
nand UO_700 (O_700,N_49284,N_47973);
or UO_701 (O_701,N_48489,N_49064);
nand UO_702 (O_702,N_47983,N_48037);
nor UO_703 (O_703,N_49362,N_49042);
nand UO_704 (O_704,N_48556,N_49548);
xor UO_705 (O_705,N_49462,N_49762);
or UO_706 (O_706,N_48961,N_49078);
xnor UO_707 (O_707,N_49140,N_47726);
and UO_708 (O_708,N_49103,N_47871);
xor UO_709 (O_709,N_48869,N_49863);
or UO_710 (O_710,N_49619,N_49474);
xor UO_711 (O_711,N_49652,N_47735);
nor UO_712 (O_712,N_48398,N_49253);
and UO_713 (O_713,N_48167,N_48280);
xnor UO_714 (O_714,N_48970,N_49844);
or UO_715 (O_715,N_49659,N_47688);
xor UO_716 (O_716,N_47560,N_49707);
nor UO_717 (O_717,N_49725,N_49761);
or UO_718 (O_718,N_48901,N_49024);
and UO_719 (O_719,N_49825,N_47949);
and UO_720 (O_720,N_48612,N_48764);
and UO_721 (O_721,N_48427,N_48597);
and UO_722 (O_722,N_48682,N_48732);
or UO_723 (O_723,N_48510,N_48688);
xnor UO_724 (O_724,N_49082,N_49560);
xnor UO_725 (O_725,N_48836,N_48425);
or UO_726 (O_726,N_49038,N_49072);
and UO_727 (O_727,N_49726,N_49010);
or UO_728 (O_728,N_49738,N_47845);
or UO_729 (O_729,N_49757,N_48717);
nor UO_730 (O_730,N_49066,N_48382);
nor UO_731 (O_731,N_49177,N_48950);
nor UO_732 (O_732,N_47840,N_49303);
or UO_733 (O_733,N_48973,N_47849);
xnor UO_734 (O_734,N_48261,N_49602);
xnor UO_735 (O_735,N_49727,N_47544);
nor UO_736 (O_736,N_48607,N_49690);
nor UO_737 (O_737,N_49011,N_48765);
xor UO_738 (O_738,N_49564,N_48584);
nand UO_739 (O_739,N_49680,N_47615);
and UO_740 (O_740,N_49512,N_49511);
nand UO_741 (O_741,N_47842,N_49685);
nor UO_742 (O_742,N_49977,N_48137);
and UO_743 (O_743,N_48670,N_48450);
or UO_744 (O_744,N_49173,N_49483);
or UO_745 (O_745,N_49100,N_49170);
nand UO_746 (O_746,N_47911,N_49878);
xor UO_747 (O_747,N_48586,N_49742);
nand UO_748 (O_748,N_47580,N_49816);
or UO_749 (O_749,N_47543,N_48378);
nand UO_750 (O_750,N_48909,N_47673);
or UO_751 (O_751,N_49665,N_48980);
xor UO_752 (O_752,N_49778,N_49090);
nand UO_753 (O_753,N_48795,N_48534);
xor UO_754 (O_754,N_48953,N_48072);
nand UO_755 (O_755,N_48011,N_48944);
nand UO_756 (O_756,N_47579,N_47857);
nand UO_757 (O_757,N_48420,N_49453);
or UO_758 (O_758,N_48707,N_47542);
and UO_759 (O_759,N_48924,N_47685);
xor UO_760 (O_760,N_49550,N_48578);
or UO_761 (O_761,N_48205,N_48074);
xnor UO_762 (O_762,N_49534,N_49610);
and UO_763 (O_763,N_49845,N_48224);
or UO_764 (O_764,N_47731,N_47817);
or UO_765 (O_765,N_48009,N_49250);
nand UO_766 (O_766,N_48609,N_49266);
xor UO_767 (O_767,N_48562,N_47621);
nor UO_768 (O_768,N_48559,N_49561);
xnor UO_769 (O_769,N_48277,N_47548);
nor UO_770 (O_770,N_47530,N_48246);
nand UO_771 (O_771,N_48821,N_48792);
or UO_772 (O_772,N_48965,N_48431);
or UO_773 (O_773,N_49298,N_49827);
and UO_774 (O_774,N_48920,N_49804);
nor UO_775 (O_775,N_49262,N_49065);
and UO_776 (O_776,N_47606,N_48200);
and UO_777 (O_777,N_47513,N_47562);
and UO_778 (O_778,N_48690,N_48839);
and UO_779 (O_779,N_47957,N_48387);
nor UO_780 (O_780,N_49540,N_48640);
or UO_781 (O_781,N_49906,N_47933);
and UO_782 (O_782,N_49122,N_48238);
and UO_783 (O_783,N_48841,N_49623);
xor UO_784 (O_784,N_48366,N_47627);
and UO_785 (O_785,N_49451,N_49171);
xor UO_786 (O_786,N_48175,N_48073);
nor UO_787 (O_787,N_49500,N_49217);
nand UO_788 (O_788,N_48046,N_49256);
nor UO_789 (O_789,N_48952,N_48467);
nand UO_790 (O_790,N_49226,N_47928);
nand UO_791 (O_791,N_48890,N_49956);
and UO_792 (O_792,N_47506,N_48084);
nor UO_793 (O_793,N_47705,N_49422);
xor UO_794 (O_794,N_47951,N_49723);
xnor UO_795 (O_795,N_48730,N_49785);
and UO_796 (O_796,N_47968,N_49176);
and UO_797 (O_797,N_48153,N_49373);
and UO_798 (O_798,N_48832,N_47572);
and UO_799 (O_799,N_48357,N_49128);
nand UO_800 (O_800,N_48249,N_48689);
nand UO_801 (O_801,N_48726,N_47926);
nor UO_802 (O_802,N_49576,N_49622);
and UO_803 (O_803,N_49499,N_49039);
nand UO_804 (O_804,N_49396,N_48747);
or UO_805 (O_805,N_49657,N_48415);
nand UO_806 (O_806,N_48316,N_48029);
or UO_807 (O_807,N_49086,N_48677);
nor UO_808 (O_808,N_49591,N_49813);
and UO_809 (O_809,N_48949,N_48177);
nand UO_810 (O_810,N_47619,N_47955);
or UO_811 (O_811,N_48995,N_47552);
xor UO_812 (O_812,N_49219,N_47996);
nand UO_813 (O_813,N_48141,N_49048);
nor UO_814 (O_814,N_49353,N_48907);
or UO_815 (O_815,N_48812,N_47972);
or UO_816 (O_816,N_49130,N_48262);
nand UO_817 (O_817,N_48506,N_47505);
nor UO_818 (O_818,N_47739,N_48388);
xnor UO_819 (O_819,N_49609,N_48064);
and UO_820 (O_820,N_49279,N_48410);
or UO_821 (O_821,N_49882,N_48393);
or UO_822 (O_822,N_48620,N_49775);
nand UO_823 (O_823,N_49113,N_49835);
nand UO_824 (O_824,N_49547,N_49645);
nor UO_825 (O_825,N_49632,N_49029);
nor UO_826 (O_826,N_48213,N_47877);
or UO_827 (O_827,N_49904,N_48255);
nand UO_828 (O_828,N_48352,N_49007);
nor UO_829 (O_829,N_49212,N_48908);
and UO_830 (O_830,N_49568,N_48951);
and UO_831 (O_831,N_47970,N_48203);
nand UO_832 (O_832,N_49979,N_48030);
xor UO_833 (O_833,N_47916,N_47524);
nand UO_834 (O_834,N_49841,N_48507);
or UO_835 (O_835,N_49233,N_48024);
nand UO_836 (O_836,N_48292,N_48790);
nor UO_837 (O_837,N_48808,N_48646);
and UO_838 (O_838,N_48300,N_49953);
nor UO_839 (O_839,N_48267,N_48752);
nor UO_840 (O_840,N_49469,N_48727);
or UO_841 (O_841,N_48659,N_48370);
nand UO_842 (O_842,N_49163,N_47514);
nand UO_843 (O_843,N_48905,N_49978);
xnor UO_844 (O_844,N_49699,N_47979);
or UO_845 (O_845,N_48672,N_47531);
or UO_846 (O_846,N_49820,N_48315);
nand UO_847 (O_847,N_48170,N_49546);
and UO_848 (O_848,N_48956,N_49295);
or UO_849 (O_849,N_48451,N_48143);
nor UO_850 (O_850,N_47669,N_49868);
and UO_851 (O_851,N_47575,N_48421);
or UO_852 (O_852,N_48463,N_49239);
xor UO_853 (O_853,N_48800,N_47644);
nor UO_854 (O_854,N_49473,N_48794);
or UO_855 (O_855,N_49348,N_48666);
and UO_856 (O_856,N_49668,N_48691);
xnor UO_857 (O_857,N_47587,N_48272);
nor UO_858 (O_858,N_47767,N_49530);
or UO_859 (O_859,N_49397,N_48809);
nor UO_860 (O_860,N_47906,N_48817);
and UO_861 (O_861,N_48798,N_47722);
or UO_862 (O_862,N_49637,N_49290);
and UO_863 (O_863,N_48781,N_49933);
nand UO_864 (O_864,N_48638,N_47594);
and UO_865 (O_865,N_48527,N_47927);
or UO_866 (O_866,N_48575,N_49460);
nor UO_867 (O_867,N_49575,N_49732);
nand UO_868 (O_868,N_49068,N_48561);
or UO_869 (O_869,N_48154,N_47847);
and UO_870 (O_870,N_48400,N_47671);
and UO_871 (O_871,N_49831,N_49331);
xnor UO_872 (O_872,N_48728,N_49687);
or UO_873 (O_873,N_49333,N_49088);
or UO_874 (O_874,N_49282,N_49880);
nor UO_875 (O_875,N_47777,N_48406);
and UO_876 (O_876,N_47875,N_47785);
nand UO_877 (O_877,N_48791,N_48834);
and UO_878 (O_878,N_49588,N_49093);
or UO_879 (O_879,N_49661,N_49671);
or UO_880 (O_880,N_48323,N_47545);
xor UO_881 (O_881,N_47715,N_49926);
xor UO_882 (O_882,N_48208,N_47987);
and UO_883 (O_883,N_48539,N_47872);
and UO_884 (O_884,N_48469,N_48937);
xnor UO_885 (O_885,N_47866,N_49245);
and UO_886 (O_886,N_49003,N_48337);
or UO_887 (O_887,N_49756,N_49181);
nor UO_888 (O_888,N_49553,N_47626);
xor UO_889 (O_889,N_48606,N_49970);
nor UO_890 (O_890,N_47834,N_48977);
nor UO_891 (O_891,N_48551,N_49255);
xor UO_892 (O_892,N_47645,N_48796);
nor UO_893 (O_893,N_48031,N_49803);
or UO_894 (O_894,N_47696,N_48641);
xnor UO_895 (O_895,N_48619,N_48473);
or UO_896 (O_896,N_48783,N_49287);
nand UO_897 (O_897,N_49162,N_49974);
or UO_898 (O_898,N_48008,N_49243);
or UO_899 (O_899,N_48922,N_49945);
and UO_900 (O_900,N_48614,N_49165);
and UO_901 (O_901,N_48573,N_47723);
xor UO_902 (O_902,N_48329,N_49232);
nand UO_903 (O_903,N_48538,N_48232);
nand UO_904 (O_904,N_47900,N_47988);
or UO_905 (O_905,N_48221,N_47605);
nand UO_906 (O_906,N_49380,N_48611);
xor UO_907 (O_907,N_48626,N_49004);
nand UO_908 (O_908,N_48521,N_49002);
or UO_909 (O_909,N_49848,N_49552);
nor UO_910 (O_910,N_48517,N_49719);
xnor UO_911 (O_911,N_48344,N_47565);
nand UO_912 (O_912,N_47653,N_48022);
xor UO_913 (O_913,N_47909,N_49873);
or UO_914 (O_914,N_49965,N_47896);
or UO_915 (O_915,N_48333,N_49427);
or UO_916 (O_916,N_49341,N_49421);
nand UO_917 (O_917,N_47724,N_47648);
nand UO_918 (O_918,N_49199,N_48829);
xnor UO_919 (O_919,N_48500,N_49400);
nor UO_920 (O_920,N_48123,N_49318);
nand UO_921 (O_921,N_48685,N_49875);
xor UO_922 (O_922,N_48231,N_48418);
xor UO_923 (O_923,N_49620,N_47720);
or UO_924 (O_924,N_48984,N_47941);
nor UO_925 (O_925,N_48855,N_49559);
and UO_926 (O_926,N_48439,N_49784);
nand UO_927 (O_927,N_48930,N_48868);
and UO_928 (O_928,N_49235,N_49673);
nand UO_929 (O_929,N_47554,N_47736);
and UO_930 (O_930,N_49361,N_48844);
nor UO_931 (O_931,N_49436,N_49261);
nor UO_932 (O_932,N_47536,N_47623);
and UO_933 (O_933,N_47508,N_48983);
or UO_934 (O_934,N_49897,N_49695);
nor UO_935 (O_935,N_48441,N_47897);
nor UO_936 (O_936,N_47651,N_48959);
or UO_937 (O_937,N_47727,N_49626);
nand UO_938 (O_938,N_48282,N_48112);
or UO_939 (O_939,N_49180,N_49847);
nand UO_940 (O_940,N_48847,N_48171);
nor UO_941 (O_941,N_48567,N_48972);
nand UO_942 (O_942,N_47683,N_47917);
or UO_943 (O_943,N_48088,N_49969);
xor UO_944 (O_944,N_48630,N_49596);
xnor UO_945 (O_945,N_47682,N_47810);
nand UO_946 (O_946,N_49951,N_48851);
nor UO_947 (O_947,N_48887,N_49132);
nor UO_948 (O_948,N_49993,N_47697);
nor UO_949 (O_949,N_48537,N_49997);
xor UO_950 (O_950,N_49860,N_48679);
and UO_951 (O_951,N_49822,N_49869);
and UO_952 (O_952,N_47629,N_48152);
or UO_953 (O_953,N_49808,N_48616);
nand UO_954 (O_954,N_47795,N_49704);
and UO_955 (O_955,N_49005,N_47969);
xor UO_956 (O_956,N_48343,N_47902);
or UO_957 (O_957,N_48089,N_47550);
nor UO_958 (O_958,N_49074,N_48086);
and UO_959 (O_959,N_48173,N_48596);
nor UO_960 (O_960,N_48007,N_49327);
and UO_961 (O_961,N_48837,N_47837);
nor UO_962 (O_962,N_48681,N_48625);
or UO_963 (O_963,N_47719,N_48615);
nor UO_964 (O_964,N_49317,N_48120);
and UO_965 (O_965,N_47701,N_49465);
xor UO_966 (O_966,N_49407,N_48742);
xor UO_967 (O_967,N_48678,N_49787);
nand UO_968 (O_968,N_49478,N_48509);
or UO_969 (O_969,N_48580,N_48263);
nand UO_970 (O_970,N_49073,N_48644);
xor UO_971 (O_971,N_49748,N_47710);
or UO_972 (O_972,N_49802,N_47755);
and UO_973 (O_973,N_49415,N_47617);
nor UO_974 (O_974,N_48830,N_49017);
and UO_975 (O_975,N_49304,N_49069);
or UO_976 (O_976,N_48815,N_49734);
nand UO_977 (O_977,N_49517,N_49156);
or UO_978 (O_978,N_47797,N_48193);
or UO_979 (O_979,N_49583,N_48148);
nand UO_980 (O_980,N_49071,N_48675);
nor UO_981 (O_981,N_49709,N_47793);
nand UO_982 (O_982,N_47835,N_49135);
and UO_983 (O_983,N_48168,N_47961);
xnor UO_984 (O_984,N_49682,N_48967);
nand UO_985 (O_985,N_49490,N_49683);
and UO_986 (O_986,N_48702,N_48405);
nand UO_987 (O_987,N_47566,N_48528);
nand UO_988 (O_988,N_47538,N_48472);
and UO_989 (O_989,N_48116,N_49063);
and UO_990 (O_990,N_49094,N_49286);
and UO_991 (O_991,N_49708,N_47576);
nor UO_992 (O_992,N_49146,N_47684);
xnor UO_993 (O_993,N_49030,N_47992);
and UO_994 (O_994,N_48627,N_49849);
xor UO_995 (O_995,N_49242,N_49694);
xor UO_996 (O_996,N_48871,N_48244);
nand UO_997 (O_997,N_49479,N_49084);
and UO_998 (O_998,N_49598,N_48335);
xor UO_999 (O_999,N_49061,N_48353);
nor UO_1000 (O_1000,N_49311,N_48608);
nor UO_1001 (O_1001,N_48819,N_47885);
nor UO_1002 (O_1002,N_49118,N_48379);
or UO_1003 (O_1003,N_47541,N_47640);
and UO_1004 (O_1004,N_47675,N_47583);
or UO_1005 (O_1005,N_49137,N_47939);
nor UO_1006 (O_1006,N_49542,N_48106);
nor UO_1007 (O_1007,N_49513,N_47689);
nand UO_1008 (O_1008,N_48117,N_47706);
nand UO_1009 (O_1009,N_49269,N_49936);
or UO_1010 (O_1010,N_49249,N_47738);
nor UO_1011 (O_1011,N_49510,N_48828);
nand UO_1012 (O_1012,N_49837,N_48722);
xor UO_1013 (O_1013,N_48719,N_47677);
or UO_1014 (O_1014,N_47591,N_49737);
and UO_1015 (O_1015,N_49741,N_48543);
nor UO_1016 (O_1016,N_48372,N_48610);
and UO_1017 (O_1017,N_48654,N_48159);
or UO_1018 (O_1018,N_47504,N_49184);
xor UO_1019 (O_1019,N_49445,N_48235);
nand UO_1020 (O_1020,N_49781,N_48182);
nor UO_1021 (O_1021,N_49463,N_48306);
xnor UO_1022 (O_1022,N_49046,N_47772);
or UO_1023 (O_1023,N_48874,N_48692);
nand UO_1024 (O_1024,N_48958,N_49688);
xnor UO_1025 (O_1025,N_49222,N_48843);
nor UO_1026 (O_1026,N_49721,N_49220);
nand UO_1027 (O_1027,N_49647,N_48454);
or UO_1028 (O_1028,N_49096,N_49054);
or UO_1029 (O_1029,N_49554,N_49730);
nand UO_1030 (O_1030,N_48417,N_47647);
nand UO_1031 (O_1031,N_47908,N_48307);
nand UO_1032 (O_1032,N_48133,N_48709);
or UO_1033 (O_1033,N_49839,N_49862);
nor UO_1034 (O_1034,N_49759,N_48737);
xor UO_1035 (O_1035,N_49686,N_47977);
or UO_1036 (O_1036,N_49208,N_49206);
nor UO_1037 (O_1037,N_48042,N_47507);
and UO_1038 (O_1038,N_47589,N_49419);
and UO_1039 (O_1039,N_47895,N_49109);
and UO_1040 (O_1040,N_49203,N_48966);
xnor UO_1041 (O_1041,N_47765,N_48183);
nor UO_1042 (O_1042,N_49768,N_49346);
and UO_1043 (O_1043,N_49910,N_49501);
or UO_1044 (O_1044,N_49852,N_49299);
nor UO_1045 (O_1045,N_49566,N_47660);
nor UO_1046 (O_1046,N_47831,N_49654);
nor UO_1047 (O_1047,N_49288,N_47821);
or UO_1048 (O_1048,N_48917,N_48655);
xnor UO_1049 (O_1049,N_49221,N_49252);
nor UO_1050 (O_1050,N_47832,N_47938);
nor UO_1051 (O_1051,N_49569,N_49522);
or UO_1052 (O_1052,N_47769,N_48669);
nand UO_1053 (O_1053,N_48738,N_48338);
nand UO_1054 (O_1054,N_49027,N_49884);
and UO_1055 (O_1055,N_49967,N_49655);
nor UO_1056 (O_1056,N_49662,N_49919);
nand UO_1057 (O_1057,N_47930,N_48921);
nor UO_1058 (O_1058,N_49653,N_47942);
xor UO_1059 (O_1059,N_47674,N_48514);
xnor UO_1060 (O_1060,N_48422,N_48195);
nor UO_1061 (O_1061,N_48862,N_49920);
nand UO_1062 (O_1062,N_49941,N_49807);
or UO_1063 (O_1063,N_48964,N_47573);
and UO_1064 (O_1064,N_49507,N_48018);
nor UO_1065 (O_1065,N_48988,N_49579);
nand UO_1066 (O_1066,N_49586,N_49639);
or UO_1067 (O_1067,N_49523,N_49819);
xnor UO_1068 (O_1068,N_47905,N_49264);
xnor UO_1069 (O_1069,N_49454,N_47668);
xnor UO_1070 (O_1070,N_47650,N_48257);
or UO_1071 (O_1071,N_48933,N_49674);
xnor UO_1072 (O_1072,N_48635,N_48547);
and UO_1073 (O_1073,N_49254,N_48436);
and UO_1074 (O_1074,N_47656,N_48041);
xor UO_1075 (O_1075,N_48059,N_48987);
nand UO_1076 (O_1076,N_47525,N_49996);
nor UO_1077 (O_1077,N_48706,N_48274);
nand UO_1078 (O_1078,N_48002,N_49669);
and UO_1079 (O_1079,N_49432,N_47962);
xor UO_1080 (O_1080,N_48671,N_48184);
nor UO_1081 (O_1081,N_49172,N_48498);
nand UO_1082 (O_1082,N_49916,N_48932);
and UO_1083 (O_1083,N_49573,N_48748);
and UO_1084 (O_1084,N_47716,N_48900);
nand UO_1085 (O_1085,N_49508,N_47692);
nand UO_1086 (O_1086,N_49491,N_49307);
nand UO_1087 (O_1087,N_48550,N_48483);
or UO_1088 (O_1088,N_49836,N_49330);
or UO_1089 (O_1089,N_48897,N_48873);
nand UO_1090 (O_1090,N_49051,N_47551);
nor UO_1091 (O_1091,N_48511,N_48895);
nor UO_1092 (O_1092,N_49070,N_49375);
xor UO_1093 (O_1093,N_49855,N_49059);
xor UO_1094 (O_1094,N_47737,N_48446);
nor UO_1095 (O_1095,N_49582,N_48006);
nor UO_1096 (O_1096,N_48295,N_47512);
xor UO_1097 (O_1097,N_49780,N_48845);
nor UO_1098 (O_1098,N_48687,N_49556);
nor UO_1099 (O_1099,N_47921,N_48270);
and UO_1100 (O_1100,N_48132,N_49306);
xor UO_1101 (O_1101,N_48870,N_49025);
or UO_1102 (O_1102,N_49417,N_48437);
nor UO_1103 (O_1103,N_48554,N_49309);
nor UO_1104 (O_1104,N_48334,N_47759);
and UO_1105 (O_1105,N_48055,N_48247);
and UO_1106 (O_1106,N_48910,N_47698);
or UO_1107 (O_1107,N_49198,N_48546);
and UO_1108 (O_1108,N_48460,N_48416);
and UO_1109 (O_1109,N_48033,N_48185);
or UO_1110 (O_1110,N_49297,N_48859);
nand UO_1111 (O_1111,N_49374,N_48268);
xor UO_1112 (O_1112,N_48703,N_49308);
or UO_1113 (O_1113,N_47870,N_47642);
or UO_1114 (O_1114,N_49158,N_47549);
nand UO_1115 (O_1115,N_49031,N_49321);
nand UO_1116 (O_1116,N_48424,N_49681);
nor UO_1117 (O_1117,N_49036,N_49325);
xnor UO_1118 (O_1118,N_48253,N_48886);
or UO_1119 (O_1119,N_47532,N_49429);
nand UO_1120 (O_1120,N_48435,N_48782);
xor UO_1121 (O_1121,N_48643,N_48996);
nor UO_1122 (O_1122,N_47800,N_49604);
and UO_1123 (O_1123,N_49931,N_49964);
nor UO_1124 (O_1124,N_48456,N_47690);
nor UO_1125 (O_1125,N_48879,N_48749);
nand UO_1126 (O_1126,N_48125,N_49486);
xnor UO_1127 (O_1127,N_49200,N_49519);
and UO_1128 (O_1128,N_48629,N_47529);
xnor UO_1129 (O_1129,N_48745,N_49535);
nor UO_1130 (O_1130,N_48058,N_48820);
and UO_1131 (O_1131,N_48309,N_48497);
xor UO_1132 (O_1132,N_49846,N_47947);
nor UO_1133 (O_1133,N_49710,N_48310);
nor UO_1134 (O_1134,N_47869,N_49151);
and UO_1135 (O_1135,N_48265,N_49300);
nand UO_1136 (O_1136,N_49468,N_47815);
xor UO_1137 (O_1137,N_49218,N_47971);
nand UO_1138 (O_1138,N_47509,N_49028);
and UO_1139 (O_1139,N_48877,N_48613);
nor UO_1140 (O_1140,N_47586,N_47760);
nor UO_1141 (O_1141,N_47699,N_49889);
and UO_1142 (O_1142,N_49905,N_48212);
and UO_1143 (O_1143,N_47799,N_49227);
and UO_1144 (O_1144,N_49360,N_49711);
or UO_1145 (O_1145,N_48515,N_47643);
xnor UO_1146 (O_1146,N_49805,N_48519);
and UO_1147 (O_1147,N_47813,N_47790);
and UO_1148 (O_1148,N_49755,N_49481);
or UO_1149 (O_1149,N_49244,N_48885);
and UO_1150 (O_1150,N_49642,N_49883);
nor UO_1151 (O_1151,N_49675,N_49442);
xor UO_1152 (O_1152,N_49365,N_48023);
nor UO_1153 (O_1153,N_49806,N_47803);
or UO_1154 (O_1154,N_48340,N_47912);
xnor UO_1155 (O_1155,N_48092,N_48201);
or UO_1156 (O_1156,N_47687,N_49322);
nand UO_1157 (O_1157,N_47946,N_48015);
xor UO_1158 (O_1158,N_49215,N_49963);
nand UO_1159 (O_1159,N_49935,N_49650);
and UO_1160 (O_1160,N_48618,N_48700);
and UO_1161 (O_1161,N_48226,N_48866);
or UO_1162 (O_1162,N_49670,N_48341);
nor UO_1163 (O_1163,N_49271,N_48477);
nor UO_1164 (O_1164,N_48014,N_49338);
xnor UO_1165 (O_1165,N_48019,N_48822);
nor UO_1166 (O_1166,N_47631,N_48636);
or UO_1167 (O_1167,N_48369,N_48720);
nand UO_1168 (O_1168,N_47965,N_47659);
nor UO_1169 (O_1169,N_48804,N_49152);
nand UO_1170 (O_1170,N_47820,N_47707);
nor UO_1171 (O_1171,N_48242,N_48079);
or UO_1172 (O_1172,N_48054,N_48407);
nor UO_1173 (O_1173,N_47904,N_47865);
and UO_1174 (O_1174,N_48284,N_47637);
nor UO_1175 (O_1175,N_48780,N_48012);
and UO_1176 (O_1176,N_48680,N_48377);
or UO_1177 (O_1177,N_48569,N_48664);
and UO_1178 (O_1178,N_49384,N_47806);
nand UO_1179 (O_1179,N_48347,N_49594);
or UO_1180 (O_1180,N_49259,N_48101);
nor UO_1181 (O_1181,N_49157,N_49537);
nor UO_1182 (O_1182,N_49412,N_48637);
or UO_1183 (O_1183,N_48767,N_47901);
and UO_1184 (O_1184,N_49713,N_48375);
nand UO_1185 (O_1185,N_49494,N_48523);
nor UO_1186 (O_1186,N_49466,N_49612);
or UO_1187 (O_1187,N_48971,N_49467);
nand UO_1188 (O_1188,N_48069,N_47630);
xnor UO_1189 (O_1189,N_49867,N_49888);
and UO_1190 (O_1190,N_47990,N_48592);
and UO_1191 (O_1191,N_47993,N_49389);
and UO_1192 (O_1192,N_48039,N_48481);
nor UO_1193 (O_1193,N_49475,N_49722);
xor UO_1194 (O_1194,N_49786,N_48857);
and UO_1195 (O_1195,N_48549,N_48955);
xnor UO_1196 (O_1196,N_49526,N_49943);
nand UO_1197 (O_1197,N_49580,N_49758);
or UO_1198 (O_1198,N_47612,N_49663);
xor UO_1199 (O_1199,N_48281,N_47882);
nor UO_1200 (O_1200,N_47676,N_49767);
xnor UO_1201 (O_1201,N_48540,N_48464);
nand UO_1202 (O_1202,N_47702,N_47931);
nand UO_1203 (O_1203,N_49691,N_47556);
nor UO_1204 (O_1204,N_48100,N_49228);
xor UO_1205 (O_1205,N_49646,N_48386);
nand UO_1206 (O_1206,N_49363,N_49488);
nor UO_1207 (O_1207,N_47666,N_49625);
nor UO_1208 (O_1208,N_48365,N_47976);
nand UO_1209 (O_1209,N_48491,N_49578);
nand UO_1210 (O_1210,N_48653,N_48192);
and UO_1211 (O_1211,N_48760,N_49105);
xnor UO_1212 (O_1212,N_47792,N_48187);
nor UO_1213 (O_1213,N_48179,N_49633);
and UO_1214 (O_1214,N_48399,N_49676);
and UO_1215 (O_1215,N_48230,N_49026);
nand UO_1216 (O_1216,N_49359,N_48993);
and UO_1217 (O_1217,N_49032,N_47680);
xor UO_1218 (O_1218,N_49416,N_49809);
or UO_1219 (O_1219,N_48581,N_49617);
xor UO_1220 (O_1220,N_49291,N_48294);
nand UO_1221 (O_1221,N_47868,N_47657);
xor UO_1222 (O_1222,N_49796,N_49581);
xnor UO_1223 (O_1223,N_47827,N_47864);
or UO_1224 (O_1224,N_49190,N_47592);
xnor UO_1225 (O_1225,N_48355,N_49698);
xnor UO_1226 (O_1226,N_48181,N_49927);
and UO_1227 (O_1227,N_49881,N_49354);
or UO_1228 (O_1228,N_49877,N_48449);
or UO_1229 (O_1229,N_47932,N_47982);
or UO_1230 (O_1230,N_49138,N_49238);
nand UO_1231 (O_1231,N_47887,N_48649);
or UO_1232 (O_1232,N_48997,N_48941);
nor UO_1233 (O_1233,N_49631,N_49854);
and UO_1234 (O_1234,N_47779,N_49608);
and UO_1235 (O_1235,N_49394,N_49543);
xor UO_1236 (O_1236,N_48134,N_48462);
nor UO_1237 (O_1237,N_49853,N_47924);
and UO_1238 (O_1238,N_47873,N_47784);
and UO_1239 (O_1239,N_49915,N_48194);
and UO_1240 (O_1240,N_49133,N_48308);
nor UO_1241 (O_1241,N_49982,N_49745);
nor UO_1242 (O_1242,N_48409,N_47747);
or UO_1243 (O_1243,N_47501,N_48766);
or UO_1244 (O_1244,N_49225,N_48929);
xnor UO_1245 (O_1245,N_49929,N_49294);
nand UO_1246 (O_1246,N_49390,N_49998);
or UO_1247 (O_1247,N_48568,N_49188);
or UO_1248 (O_1248,N_49932,N_48852);
nand UO_1249 (O_1249,N_49799,N_48553);
or UO_1250 (O_1250,N_48946,N_48631);
xnor UO_1251 (O_1251,N_48463,N_48312);
nand UO_1252 (O_1252,N_47960,N_49828);
nand UO_1253 (O_1253,N_47981,N_49308);
xor UO_1254 (O_1254,N_48826,N_47933);
xnor UO_1255 (O_1255,N_47799,N_49277);
and UO_1256 (O_1256,N_49067,N_48316);
xor UO_1257 (O_1257,N_49824,N_48183);
nand UO_1258 (O_1258,N_48821,N_49172);
xnor UO_1259 (O_1259,N_49764,N_48823);
and UO_1260 (O_1260,N_48506,N_49028);
and UO_1261 (O_1261,N_48128,N_49905);
and UO_1262 (O_1262,N_47527,N_48084);
xor UO_1263 (O_1263,N_48143,N_48386);
nor UO_1264 (O_1264,N_48260,N_49684);
or UO_1265 (O_1265,N_49628,N_48122);
and UO_1266 (O_1266,N_49112,N_47558);
nor UO_1267 (O_1267,N_47569,N_49659);
or UO_1268 (O_1268,N_48240,N_47589);
and UO_1269 (O_1269,N_48880,N_49216);
and UO_1270 (O_1270,N_47783,N_49169);
nand UO_1271 (O_1271,N_48054,N_48088);
and UO_1272 (O_1272,N_47857,N_47775);
nor UO_1273 (O_1273,N_48837,N_47990);
and UO_1274 (O_1274,N_47531,N_49166);
nand UO_1275 (O_1275,N_48582,N_48889);
and UO_1276 (O_1276,N_48963,N_48790);
and UO_1277 (O_1277,N_47611,N_49794);
xor UO_1278 (O_1278,N_48264,N_49415);
and UO_1279 (O_1279,N_49712,N_49407);
nand UO_1280 (O_1280,N_49405,N_48188);
xnor UO_1281 (O_1281,N_48949,N_48661);
and UO_1282 (O_1282,N_48796,N_49958);
xnor UO_1283 (O_1283,N_48740,N_49083);
nand UO_1284 (O_1284,N_49840,N_48763);
or UO_1285 (O_1285,N_47550,N_47816);
and UO_1286 (O_1286,N_49634,N_49865);
or UO_1287 (O_1287,N_48920,N_47701);
or UO_1288 (O_1288,N_48545,N_49159);
nor UO_1289 (O_1289,N_48896,N_47718);
or UO_1290 (O_1290,N_48872,N_47850);
nor UO_1291 (O_1291,N_47920,N_48906);
nor UO_1292 (O_1292,N_49409,N_48979);
xor UO_1293 (O_1293,N_47688,N_49867);
nor UO_1294 (O_1294,N_49443,N_49432);
nor UO_1295 (O_1295,N_49067,N_49091);
or UO_1296 (O_1296,N_49160,N_49237);
and UO_1297 (O_1297,N_47919,N_49104);
xor UO_1298 (O_1298,N_48788,N_48255);
nand UO_1299 (O_1299,N_47694,N_48612);
nand UO_1300 (O_1300,N_49800,N_48505);
and UO_1301 (O_1301,N_49311,N_48980);
and UO_1302 (O_1302,N_49517,N_47750);
xor UO_1303 (O_1303,N_49569,N_47732);
nand UO_1304 (O_1304,N_47844,N_49930);
nand UO_1305 (O_1305,N_49927,N_47502);
and UO_1306 (O_1306,N_48775,N_47642);
nor UO_1307 (O_1307,N_49320,N_48371);
and UO_1308 (O_1308,N_49449,N_49461);
or UO_1309 (O_1309,N_49618,N_49722);
and UO_1310 (O_1310,N_49521,N_48025);
or UO_1311 (O_1311,N_48511,N_48660);
nand UO_1312 (O_1312,N_49935,N_49930);
and UO_1313 (O_1313,N_47743,N_49409);
nor UO_1314 (O_1314,N_48544,N_49400);
nand UO_1315 (O_1315,N_47939,N_49732);
xor UO_1316 (O_1316,N_49803,N_49179);
xor UO_1317 (O_1317,N_49633,N_48514);
xnor UO_1318 (O_1318,N_47682,N_49438);
or UO_1319 (O_1319,N_48518,N_48123);
or UO_1320 (O_1320,N_48314,N_48764);
or UO_1321 (O_1321,N_48420,N_48847);
nor UO_1322 (O_1322,N_48932,N_49395);
xor UO_1323 (O_1323,N_48333,N_49018);
xnor UO_1324 (O_1324,N_48847,N_48441);
nor UO_1325 (O_1325,N_47560,N_47709);
xor UO_1326 (O_1326,N_47779,N_49197);
and UO_1327 (O_1327,N_48749,N_49139);
or UO_1328 (O_1328,N_47695,N_47855);
nand UO_1329 (O_1329,N_47613,N_47744);
xor UO_1330 (O_1330,N_49337,N_48282);
or UO_1331 (O_1331,N_47746,N_47715);
nand UO_1332 (O_1332,N_48160,N_48515);
and UO_1333 (O_1333,N_49850,N_49042);
or UO_1334 (O_1334,N_49785,N_48375);
or UO_1335 (O_1335,N_48854,N_48536);
nand UO_1336 (O_1336,N_48948,N_49217);
nor UO_1337 (O_1337,N_49202,N_48561);
and UO_1338 (O_1338,N_48924,N_49620);
xor UO_1339 (O_1339,N_48605,N_48808);
and UO_1340 (O_1340,N_49752,N_49348);
xor UO_1341 (O_1341,N_49570,N_47680);
nand UO_1342 (O_1342,N_49342,N_49796);
nor UO_1343 (O_1343,N_48189,N_49641);
xor UO_1344 (O_1344,N_49360,N_47759);
xor UO_1345 (O_1345,N_49700,N_49877);
nand UO_1346 (O_1346,N_47875,N_48350);
and UO_1347 (O_1347,N_49934,N_49412);
nor UO_1348 (O_1348,N_48254,N_47688);
nor UO_1349 (O_1349,N_48565,N_49056);
nor UO_1350 (O_1350,N_47851,N_48627);
nand UO_1351 (O_1351,N_47818,N_49752);
nand UO_1352 (O_1352,N_48128,N_47616);
xnor UO_1353 (O_1353,N_49836,N_48360);
nor UO_1354 (O_1354,N_47850,N_49989);
and UO_1355 (O_1355,N_48197,N_48056);
or UO_1356 (O_1356,N_47653,N_49794);
and UO_1357 (O_1357,N_49341,N_48194);
or UO_1358 (O_1358,N_47675,N_48865);
or UO_1359 (O_1359,N_48153,N_48263);
and UO_1360 (O_1360,N_47983,N_49945);
xnor UO_1361 (O_1361,N_47762,N_47502);
or UO_1362 (O_1362,N_48304,N_49018);
nand UO_1363 (O_1363,N_47635,N_49571);
or UO_1364 (O_1364,N_49740,N_48803);
xnor UO_1365 (O_1365,N_48860,N_49916);
nor UO_1366 (O_1366,N_48917,N_49295);
and UO_1367 (O_1367,N_48477,N_49236);
or UO_1368 (O_1368,N_48424,N_48895);
xor UO_1369 (O_1369,N_48162,N_47809);
or UO_1370 (O_1370,N_49560,N_49429);
nor UO_1371 (O_1371,N_47914,N_48343);
or UO_1372 (O_1372,N_47733,N_47802);
nand UO_1373 (O_1373,N_47612,N_49860);
nor UO_1374 (O_1374,N_48171,N_48166);
nand UO_1375 (O_1375,N_47980,N_47501);
nor UO_1376 (O_1376,N_47638,N_48615);
xor UO_1377 (O_1377,N_48626,N_49483);
or UO_1378 (O_1378,N_47966,N_49846);
or UO_1379 (O_1379,N_49376,N_48413);
xnor UO_1380 (O_1380,N_49462,N_49144);
and UO_1381 (O_1381,N_47893,N_49810);
xnor UO_1382 (O_1382,N_48976,N_48144);
or UO_1383 (O_1383,N_48694,N_49662);
xnor UO_1384 (O_1384,N_48496,N_47835);
or UO_1385 (O_1385,N_48944,N_48893);
nor UO_1386 (O_1386,N_47908,N_49287);
or UO_1387 (O_1387,N_49222,N_47842);
nor UO_1388 (O_1388,N_48200,N_47576);
xnor UO_1389 (O_1389,N_49395,N_49368);
or UO_1390 (O_1390,N_47754,N_47790);
xor UO_1391 (O_1391,N_48415,N_48979);
nor UO_1392 (O_1392,N_48227,N_49445);
xnor UO_1393 (O_1393,N_47731,N_49326);
or UO_1394 (O_1394,N_48610,N_49136);
xnor UO_1395 (O_1395,N_47747,N_47961);
and UO_1396 (O_1396,N_48419,N_48499);
nor UO_1397 (O_1397,N_48231,N_47501);
nor UO_1398 (O_1398,N_47969,N_48029);
nor UO_1399 (O_1399,N_49298,N_49662);
nand UO_1400 (O_1400,N_47738,N_48137);
nand UO_1401 (O_1401,N_49497,N_48293);
nand UO_1402 (O_1402,N_48087,N_47908);
and UO_1403 (O_1403,N_48493,N_49367);
nor UO_1404 (O_1404,N_47554,N_48888);
and UO_1405 (O_1405,N_48212,N_48744);
nand UO_1406 (O_1406,N_48501,N_48197);
nand UO_1407 (O_1407,N_47840,N_48866);
nand UO_1408 (O_1408,N_48242,N_48896);
nand UO_1409 (O_1409,N_49310,N_48553);
and UO_1410 (O_1410,N_49563,N_48886);
and UO_1411 (O_1411,N_48101,N_49922);
nand UO_1412 (O_1412,N_48734,N_48053);
nand UO_1413 (O_1413,N_48636,N_47959);
xor UO_1414 (O_1414,N_48632,N_47783);
and UO_1415 (O_1415,N_48945,N_48610);
nand UO_1416 (O_1416,N_47614,N_47747);
nor UO_1417 (O_1417,N_47756,N_49493);
nor UO_1418 (O_1418,N_49321,N_47703);
and UO_1419 (O_1419,N_47675,N_47796);
or UO_1420 (O_1420,N_47701,N_48549);
nand UO_1421 (O_1421,N_47584,N_48914);
xor UO_1422 (O_1422,N_48038,N_48169);
nand UO_1423 (O_1423,N_49524,N_48675);
nand UO_1424 (O_1424,N_47858,N_49963);
nor UO_1425 (O_1425,N_48453,N_47508);
and UO_1426 (O_1426,N_49707,N_48319);
xor UO_1427 (O_1427,N_49758,N_48157);
nand UO_1428 (O_1428,N_48943,N_48135);
xnor UO_1429 (O_1429,N_49954,N_48327);
nand UO_1430 (O_1430,N_49023,N_49918);
or UO_1431 (O_1431,N_47599,N_47735);
nor UO_1432 (O_1432,N_49374,N_48924);
or UO_1433 (O_1433,N_48850,N_49506);
and UO_1434 (O_1434,N_48597,N_48949);
nor UO_1435 (O_1435,N_48888,N_47518);
xor UO_1436 (O_1436,N_49036,N_49486);
or UO_1437 (O_1437,N_49177,N_47754);
and UO_1438 (O_1438,N_48538,N_48734);
nor UO_1439 (O_1439,N_48988,N_47671);
or UO_1440 (O_1440,N_49622,N_49142);
xnor UO_1441 (O_1441,N_47564,N_48359);
nor UO_1442 (O_1442,N_48378,N_48929);
xnor UO_1443 (O_1443,N_49531,N_48126);
nor UO_1444 (O_1444,N_49204,N_47799);
and UO_1445 (O_1445,N_47890,N_49225);
nand UO_1446 (O_1446,N_49449,N_49653);
or UO_1447 (O_1447,N_48641,N_49760);
nor UO_1448 (O_1448,N_49806,N_49485);
nor UO_1449 (O_1449,N_48300,N_48095);
nand UO_1450 (O_1450,N_49172,N_48318);
xnor UO_1451 (O_1451,N_49457,N_48028);
nand UO_1452 (O_1452,N_49090,N_49748);
nor UO_1453 (O_1453,N_48421,N_49782);
nand UO_1454 (O_1454,N_47517,N_48040);
nor UO_1455 (O_1455,N_48371,N_49425);
nor UO_1456 (O_1456,N_49387,N_49998);
nand UO_1457 (O_1457,N_47791,N_47638);
nor UO_1458 (O_1458,N_48116,N_49131);
and UO_1459 (O_1459,N_48231,N_47977);
nand UO_1460 (O_1460,N_47852,N_48175);
nor UO_1461 (O_1461,N_48337,N_48848);
nor UO_1462 (O_1462,N_47897,N_49736);
xnor UO_1463 (O_1463,N_48698,N_49356);
nor UO_1464 (O_1464,N_49403,N_49873);
nor UO_1465 (O_1465,N_49265,N_47512);
or UO_1466 (O_1466,N_49202,N_48937);
and UO_1467 (O_1467,N_48917,N_49740);
nand UO_1468 (O_1468,N_49959,N_47625);
or UO_1469 (O_1469,N_47877,N_48613);
xor UO_1470 (O_1470,N_49030,N_48469);
nand UO_1471 (O_1471,N_49331,N_49728);
or UO_1472 (O_1472,N_48190,N_49788);
nand UO_1473 (O_1473,N_47783,N_48730);
nand UO_1474 (O_1474,N_47931,N_48700);
or UO_1475 (O_1475,N_49301,N_48753);
nand UO_1476 (O_1476,N_48999,N_48787);
nand UO_1477 (O_1477,N_49334,N_48122);
nor UO_1478 (O_1478,N_48875,N_48697);
nand UO_1479 (O_1479,N_48781,N_48896);
xor UO_1480 (O_1480,N_47667,N_48509);
xor UO_1481 (O_1481,N_49486,N_47791);
or UO_1482 (O_1482,N_49083,N_48550);
nand UO_1483 (O_1483,N_49311,N_49540);
nor UO_1484 (O_1484,N_48377,N_48917);
nand UO_1485 (O_1485,N_49839,N_48314);
or UO_1486 (O_1486,N_49119,N_47774);
nor UO_1487 (O_1487,N_49415,N_47767);
nand UO_1488 (O_1488,N_49747,N_49974);
and UO_1489 (O_1489,N_49745,N_48633);
or UO_1490 (O_1490,N_47999,N_48077);
and UO_1491 (O_1491,N_48445,N_49831);
xor UO_1492 (O_1492,N_49378,N_49542);
nor UO_1493 (O_1493,N_48678,N_47595);
or UO_1494 (O_1494,N_49847,N_49168);
nand UO_1495 (O_1495,N_47640,N_47987);
xor UO_1496 (O_1496,N_49208,N_48957);
or UO_1497 (O_1497,N_49130,N_47501);
and UO_1498 (O_1498,N_48238,N_49918);
and UO_1499 (O_1499,N_47540,N_48586);
nand UO_1500 (O_1500,N_47809,N_49835);
nand UO_1501 (O_1501,N_48389,N_48828);
or UO_1502 (O_1502,N_49730,N_48875);
nor UO_1503 (O_1503,N_48709,N_47739);
or UO_1504 (O_1504,N_47544,N_49932);
or UO_1505 (O_1505,N_48393,N_48585);
nor UO_1506 (O_1506,N_49892,N_47630);
and UO_1507 (O_1507,N_49751,N_48119);
xnor UO_1508 (O_1508,N_48323,N_49875);
or UO_1509 (O_1509,N_48169,N_49898);
nand UO_1510 (O_1510,N_48645,N_49933);
and UO_1511 (O_1511,N_47506,N_49960);
and UO_1512 (O_1512,N_47753,N_48718);
xor UO_1513 (O_1513,N_49913,N_49999);
and UO_1514 (O_1514,N_49191,N_48298);
or UO_1515 (O_1515,N_48382,N_49885);
or UO_1516 (O_1516,N_48528,N_49860);
nand UO_1517 (O_1517,N_47946,N_49023);
or UO_1518 (O_1518,N_47552,N_47611);
or UO_1519 (O_1519,N_48640,N_48887);
or UO_1520 (O_1520,N_48867,N_48870);
and UO_1521 (O_1521,N_48026,N_48114);
xor UO_1522 (O_1522,N_49474,N_49589);
xnor UO_1523 (O_1523,N_48270,N_48405);
or UO_1524 (O_1524,N_48524,N_49143);
nor UO_1525 (O_1525,N_48545,N_48114);
or UO_1526 (O_1526,N_48603,N_48333);
or UO_1527 (O_1527,N_49548,N_49265);
nand UO_1528 (O_1528,N_49443,N_49504);
or UO_1529 (O_1529,N_48883,N_47708);
nand UO_1530 (O_1530,N_49080,N_48405);
or UO_1531 (O_1531,N_48169,N_48998);
nand UO_1532 (O_1532,N_48925,N_48139);
or UO_1533 (O_1533,N_47660,N_48709);
or UO_1534 (O_1534,N_49665,N_49892);
xnor UO_1535 (O_1535,N_49472,N_49465);
and UO_1536 (O_1536,N_48693,N_48526);
nor UO_1537 (O_1537,N_47814,N_47968);
and UO_1538 (O_1538,N_47757,N_49375);
and UO_1539 (O_1539,N_48869,N_49867);
and UO_1540 (O_1540,N_48562,N_48007);
and UO_1541 (O_1541,N_49185,N_49523);
nand UO_1542 (O_1542,N_49291,N_47570);
nor UO_1543 (O_1543,N_47800,N_47893);
or UO_1544 (O_1544,N_48539,N_49050);
xnor UO_1545 (O_1545,N_48317,N_49225);
xor UO_1546 (O_1546,N_48749,N_49482);
nor UO_1547 (O_1547,N_49899,N_49254);
nor UO_1548 (O_1548,N_48998,N_48534);
xor UO_1549 (O_1549,N_49618,N_48683);
or UO_1550 (O_1550,N_48506,N_49048);
and UO_1551 (O_1551,N_47817,N_49301);
nor UO_1552 (O_1552,N_49801,N_47550);
and UO_1553 (O_1553,N_49617,N_48057);
and UO_1554 (O_1554,N_48293,N_49321);
or UO_1555 (O_1555,N_47551,N_49044);
and UO_1556 (O_1556,N_49641,N_49975);
or UO_1557 (O_1557,N_49254,N_47855);
and UO_1558 (O_1558,N_49534,N_48430);
xor UO_1559 (O_1559,N_49396,N_49409);
or UO_1560 (O_1560,N_49216,N_48273);
xnor UO_1561 (O_1561,N_49714,N_49487);
and UO_1562 (O_1562,N_47938,N_49290);
nand UO_1563 (O_1563,N_48362,N_49785);
or UO_1564 (O_1564,N_48002,N_47666);
nor UO_1565 (O_1565,N_48712,N_49308);
and UO_1566 (O_1566,N_47591,N_48562);
and UO_1567 (O_1567,N_48971,N_49299);
xor UO_1568 (O_1568,N_47927,N_49839);
nand UO_1569 (O_1569,N_48162,N_49049);
or UO_1570 (O_1570,N_49814,N_48669);
and UO_1571 (O_1571,N_48931,N_47587);
xnor UO_1572 (O_1572,N_47573,N_49199);
and UO_1573 (O_1573,N_49636,N_48797);
xnor UO_1574 (O_1574,N_49417,N_47706);
and UO_1575 (O_1575,N_48909,N_48946);
or UO_1576 (O_1576,N_48992,N_47904);
and UO_1577 (O_1577,N_47830,N_49529);
nor UO_1578 (O_1578,N_48034,N_47524);
and UO_1579 (O_1579,N_47755,N_48266);
and UO_1580 (O_1580,N_49986,N_49448);
or UO_1581 (O_1581,N_47892,N_48696);
and UO_1582 (O_1582,N_48378,N_48989);
or UO_1583 (O_1583,N_49887,N_47970);
xnor UO_1584 (O_1584,N_48652,N_48101);
nand UO_1585 (O_1585,N_49655,N_49011);
xnor UO_1586 (O_1586,N_47820,N_48247);
and UO_1587 (O_1587,N_48415,N_48386);
nand UO_1588 (O_1588,N_49295,N_49820);
nand UO_1589 (O_1589,N_48403,N_49157);
nand UO_1590 (O_1590,N_47654,N_47777);
xor UO_1591 (O_1591,N_47995,N_48750);
nor UO_1592 (O_1592,N_47940,N_47803);
nor UO_1593 (O_1593,N_48222,N_48865);
nor UO_1594 (O_1594,N_49167,N_48217);
and UO_1595 (O_1595,N_49509,N_49808);
nor UO_1596 (O_1596,N_48083,N_48268);
nand UO_1597 (O_1597,N_48890,N_47791);
nor UO_1598 (O_1598,N_48517,N_48117);
xnor UO_1599 (O_1599,N_49455,N_48214);
or UO_1600 (O_1600,N_47633,N_48658);
nand UO_1601 (O_1601,N_48940,N_48140);
xnor UO_1602 (O_1602,N_49868,N_48714);
xor UO_1603 (O_1603,N_48445,N_49683);
nor UO_1604 (O_1604,N_47622,N_48325);
or UO_1605 (O_1605,N_49472,N_47514);
and UO_1606 (O_1606,N_48633,N_47539);
nor UO_1607 (O_1607,N_49241,N_48206);
or UO_1608 (O_1608,N_49740,N_49854);
nand UO_1609 (O_1609,N_48473,N_47836);
nor UO_1610 (O_1610,N_49941,N_48231);
and UO_1611 (O_1611,N_49980,N_48105);
nand UO_1612 (O_1612,N_49796,N_47914);
xor UO_1613 (O_1613,N_48252,N_49965);
nor UO_1614 (O_1614,N_49298,N_48031);
nand UO_1615 (O_1615,N_48862,N_48188);
nor UO_1616 (O_1616,N_49498,N_48956);
nand UO_1617 (O_1617,N_49880,N_48210);
nand UO_1618 (O_1618,N_48415,N_49636);
or UO_1619 (O_1619,N_48274,N_49726);
and UO_1620 (O_1620,N_49113,N_49029);
nand UO_1621 (O_1621,N_48077,N_48317);
nand UO_1622 (O_1622,N_49688,N_49424);
nand UO_1623 (O_1623,N_48023,N_48516);
and UO_1624 (O_1624,N_47643,N_49739);
nor UO_1625 (O_1625,N_48438,N_47854);
and UO_1626 (O_1626,N_49588,N_49075);
xor UO_1627 (O_1627,N_49147,N_49218);
or UO_1628 (O_1628,N_47548,N_48499);
or UO_1629 (O_1629,N_49912,N_49622);
xor UO_1630 (O_1630,N_48004,N_48916);
nand UO_1631 (O_1631,N_49768,N_48497);
and UO_1632 (O_1632,N_48123,N_48461);
nand UO_1633 (O_1633,N_47534,N_49206);
xor UO_1634 (O_1634,N_49211,N_48693);
xor UO_1635 (O_1635,N_48807,N_47579);
or UO_1636 (O_1636,N_49765,N_49730);
nand UO_1637 (O_1637,N_47727,N_47818);
xnor UO_1638 (O_1638,N_48511,N_48416);
nand UO_1639 (O_1639,N_48014,N_47859);
xor UO_1640 (O_1640,N_47530,N_49796);
xnor UO_1641 (O_1641,N_49613,N_47672);
and UO_1642 (O_1642,N_48723,N_48036);
and UO_1643 (O_1643,N_48954,N_47616);
nand UO_1644 (O_1644,N_49646,N_48934);
nand UO_1645 (O_1645,N_48978,N_48144);
or UO_1646 (O_1646,N_49260,N_48093);
or UO_1647 (O_1647,N_49075,N_49416);
and UO_1648 (O_1648,N_49916,N_47774);
xnor UO_1649 (O_1649,N_48710,N_47618);
and UO_1650 (O_1650,N_48097,N_49681);
and UO_1651 (O_1651,N_48253,N_49430);
nand UO_1652 (O_1652,N_49562,N_47696);
and UO_1653 (O_1653,N_48793,N_48328);
nor UO_1654 (O_1654,N_48758,N_49247);
or UO_1655 (O_1655,N_48278,N_48372);
xnor UO_1656 (O_1656,N_49806,N_48371);
nand UO_1657 (O_1657,N_47609,N_48153);
nand UO_1658 (O_1658,N_49489,N_48366);
or UO_1659 (O_1659,N_48582,N_48910);
and UO_1660 (O_1660,N_49914,N_49597);
and UO_1661 (O_1661,N_48328,N_49967);
xor UO_1662 (O_1662,N_49947,N_48002);
and UO_1663 (O_1663,N_49212,N_49381);
and UO_1664 (O_1664,N_48147,N_49863);
xnor UO_1665 (O_1665,N_49692,N_49791);
xor UO_1666 (O_1666,N_49973,N_48026);
xnor UO_1667 (O_1667,N_49667,N_48124);
and UO_1668 (O_1668,N_49899,N_49713);
and UO_1669 (O_1669,N_48476,N_48545);
xor UO_1670 (O_1670,N_48793,N_47738);
and UO_1671 (O_1671,N_48644,N_47978);
or UO_1672 (O_1672,N_47863,N_48232);
nand UO_1673 (O_1673,N_48302,N_49384);
or UO_1674 (O_1674,N_47886,N_47691);
nand UO_1675 (O_1675,N_48993,N_49630);
and UO_1676 (O_1676,N_48241,N_48017);
or UO_1677 (O_1677,N_49103,N_47825);
and UO_1678 (O_1678,N_49061,N_47932);
nand UO_1679 (O_1679,N_48407,N_48499);
nor UO_1680 (O_1680,N_48327,N_49001);
nand UO_1681 (O_1681,N_49987,N_49914);
and UO_1682 (O_1682,N_48286,N_47844);
xor UO_1683 (O_1683,N_47531,N_49425);
nor UO_1684 (O_1684,N_48411,N_48739);
nand UO_1685 (O_1685,N_48918,N_49505);
xor UO_1686 (O_1686,N_49358,N_49647);
nand UO_1687 (O_1687,N_48260,N_47507);
xor UO_1688 (O_1688,N_48121,N_49855);
xor UO_1689 (O_1689,N_48926,N_49005);
or UO_1690 (O_1690,N_47658,N_48805);
nand UO_1691 (O_1691,N_49216,N_49050);
xnor UO_1692 (O_1692,N_49629,N_47592);
nor UO_1693 (O_1693,N_49626,N_47684);
xor UO_1694 (O_1694,N_49885,N_49560);
nor UO_1695 (O_1695,N_49776,N_47780);
and UO_1696 (O_1696,N_48841,N_49818);
xor UO_1697 (O_1697,N_49324,N_49063);
and UO_1698 (O_1698,N_49654,N_49829);
xnor UO_1699 (O_1699,N_47930,N_49479);
xnor UO_1700 (O_1700,N_48966,N_48503);
nand UO_1701 (O_1701,N_49512,N_48995);
and UO_1702 (O_1702,N_49949,N_49137);
xor UO_1703 (O_1703,N_49446,N_48564);
nand UO_1704 (O_1704,N_49036,N_47683);
or UO_1705 (O_1705,N_49630,N_49632);
nor UO_1706 (O_1706,N_49637,N_48381);
xnor UO_1707 (O_1707,N_49292,N_49413);
nor UO_1708 (O_1708,N_48327,N_49249);
or UO_1709 (O_1709,N_48851,N_49150);
nor UO_1710 (O_1710,N_49642,N_47546);
and UO_1711 (O_1711,N_48171,N_49232);
xor UO_1712 (O_1712,N_48164,N_49007);
xnor UO_1713 (O_1713,N_48971,N_49874);
nand UO_1714 (O_1714,N_48124,N_48041);
nand UO_1715 (O_1715,N_49916,N_49136);
nand UO_1716 (O_1716,N_47542,N_48120);
or UO_1717 (O_1717,N_47959,N_49140);
nand UO_1718 (O_1718,N_49083,N_49251);
or UO_1719 (O_1719,N_49565,N_48442);
nand UO_1720 (O_1720,N_48805,N_48774);
or UO_1721 (O_1721,N_48966,N_48108);
and UO_1722 (O_1722,N_48164,N_49559);
and UO_1723 (O_1723,N_48556,N_49123);
nor UO_1724 (O_1724,N_47952,N_49527);
nor UO_1725 (O_1725,N_49603,N_49709);
xnor UO_1726 (O_1726,N_48027,N_48436);
nor UO_1727 (O_1727,N_48147,N_47510);
nor UO_1728 (O_1728,N_48840,N_49637);
or UO_1729 (O_1729,N_49614,N_49904);
or UO_1730 (O_1730,N_48144,N_48614);
nand UO_1731 (O_1731,N_49660,N_49162);
and UO_1732 (O_1732,N_48895,N_48273);
nor UO_1733 (O_1733,N_49092,N_49265);
or UO_1734 (O_1734,N_49312,N_47631);
or UO_1735 (O_1735,N_47729,N_49376);
xor UO_1736 (O_1736,N_49319,N_49170);
xor UO_1737 (O_1737,N_49271,N_49182);
or UO_1738 (O_1738,N_48172,N_49268);
nor UO_1739 (O_1739,N_48858,N_49789);
or UO_1740 (O_1740,N_47928,N_47851);
nand UO_1741 (O_1741,N_49179,N_49593);
nand UO_1742 (O_1742,N_49331,N_47593);
nor UO_1743 (O_1743,N_48008,N_49594);
or UO_1744 (O_1744,N_49100,N_48924);
nor UO_1745 (O_1745,N_48520,N_47815);
and UO_1746 (O_1746,N_49846,N_47559);
xor UO_1747 (O_1747,N_49429,N_47665);
and UO_1748 (O_1748,N_47635,N_49960);
nor UO_1749 (O_1749,N_48278,N_48984);
nor UO_1750 (O_1750,N_48480,N_49354);
nand UO_1751 (O_1751,N_47873,N_48351);
or UO_1752 (O_1752,N_47552,N_47705);
xnor UO_1753 (O_1753,N_48916,N_47942);
xnor UO_1754 (O_1754,N_47961,N_47620);
or UO_1755 (O_1755,N_48408,N_47791);
xnor UO_1756 (O_1756,N_48229,N_48127);
or UO_1757 (O_1757,N_47996,N_47988);
nor UO_1758 (O_1758,N_49101,N_48615);
and UO_1759 (O_1759,N_49507,N_49746);
nand UO_1760 (O_1760,N_49156,N_49534);
nor UO_1761 (O_1761,N_48750,N_49781);
nor UO_1762 (O_1762,N_49061,N_48165);
nand UO_1763 (O_1763,N_48521,N_47668);
or UO_1764 (O_1764,N_48709,N_47985);
nand UO_1765 (O_1765,N_48328,N_48752);
and UO_1766 (O_1766,N_48751,N_47890);
xor UO_1767 (O_1767,N_49471,N_49472);
nor UO_1768 (O_1768,N_49335,N_49490);
and UO_1769 (O_1769,N_47731,N_48557);
xnor UO_1770 (O_1770,N_47928,N_47879);
or UO_1771 (O_1771,N_48735,N_49836);
nor UO_1772 (O_1772,N_48843,N_48520);
and UO_1773 (O_1773,N_48297,N_49611);
nand UO_1774 (O_1774,N_49351,N_49846);
and UO_1775 (O_1775,N_49224,N_49829);
and UO_1776 (O_1776,N_48825,N_49704);
and UO_1777 (O_1777,N_49711,N_48141);
xnor UO_1778 (O_1778,N_47875,N_49746);
or UO_1779 (O_1779,N_49284,N_49979);
nand UO_1780 (O_1780,N_49848,N_48347);
or UO_1781 (O_1781,N_48453,N_49950);
and UO_1782 (O_1782,N_49130,N_47643);
nand UO_1783 (O_1783,N_49158,N_49803);
or UO_1784 (O_1784,N_47633,N_47782);
nand UO_1785 (O_1785,N_47630,N_49507);
xnor UO_1786 (O_1786,N_48204,N_49465);
nand UO_1787 (O_1787,N_49882,N_49649);
nand UO_1788 (O_1788,N_48960,N_48149);
or UO_1789 (O_1789,N_48148,N_49350);
or UO_1790 (O_1790,N_47910,N_47967);
nand UO_1791 (O_1791,N_47641,N_49387);
nand UO_1792 (O_1792,N_49474,N_48694);
nor UO_1793 (O_1793,N_48902,N_49732);
nand UO_1794 (O_1794,N_49509,N_49239);
or UO_1795 (O_1795,N_49794,N_48560);
nand UO_1796 (O_1796,N_48280,N_48023);
or UO_1797 (O_1797,N_49021,N_47885);
nand UO_1798 (O_1798,N_49471,N_48429);
and UO_1799 (O_1799,N_47939,N_48243);
xor UO_1800 (O_1800,N_48923,N_48231);
and UO_1801 (O_1801,N_49649,N_48393);
nor UO_1802 (O_1802,N_47872,N_48748);
nor UO_1803 (O_1803,N_48949,N_47795);
xnor UO_1804 (O_1804,N_49803,N_49546);
nor UO_1805 (O_1805,N_47663,N_49291);
or UO_1806 (O_1806,N_48749,N_49193);
nand UO_1807 (O_1807,N_49360,N_47677);
nor UO_1808 (O_1808,N_49638,N_48971);
nand UO_1809 (O_1809,N_48955,N_47739);
and UO_1810 (O_1810,N_47536,N_48731);
or UO_1811 (O_1811,N_47571,N_49394);
and UO_1812 (O_1812,N_49010,N_48000);
nor UO_1813 (O_1813,N_49160,N_47769);
xor UO_1814 (O_1814,N_49165,N_48713);
nand UO_1815 (O_1815,N_49080,N_48138);
or UO_1816 (O_1816,N_49773,N_48888);
and UO_1817 (O_1817,N_48683,N_48717);
nor UO_1818 (O_1818,N_49758,N_47919);
or UO_1819 (O_1819,N_48845,N_49950);
or UO_1820 (O_1820,N_48309,N_48700);
or UO_1821 (O_1821,N_48887,N_49213);
and UO_1822 (O_1822,N_47629,N_48246);
nand UO_1823 (O_1823,N_47793,N_48152);
xnor UO_1824 (O_1824,N_48701,N_48433);
nand UO_1825 (O_1825,N_47781,N_48013);
nor UO_1826 (O_1826,N_48414,N_48905);
or UO_1827 (O_1827,N_49882,N_48890);
nor UO_1828 (O_1828,N_47982,N_49319);
nor UO_1829 (O_1829,N_49336,N_48159);
nor UO_1830 (O_1830,N_49413,N_49770);
nor UO_1831 (O_1831,N_48633,N_49601);
nor UO_1832 (O_1832,N_49142,N_49146);
or UO_1833 (O_1833,N_48895,N_49556);
or UO_1834 (O_1834,N_48854,N_47991);
xnor UO_1835 (O_1835,N_48661,N_49885);
xor UO_1836 (O_1836,N_49238,N_47577);
nor UO_1837 (O_1837,N_47773,N_49056);
nand UO_1838 (O_1838,N_49891,N_48497);
and UO_1839 (O_1839,N_48794,N_49060);
nor UO_1840 (O_1840,N_49670,N_48279);
xnor UO_1841 (O_1841,N_49436,N_49111);
and UO_1842 (O_1842,N_47679,N_48057);
and UO_1843 (O_1843,N_49488,N_48334);
nor UO_1844 (O_1844,N_48891,N_49444);
or UO_1845 (O_1845,N_48857,N_49993);
and UO_1846 (O_1846,N_49216,N_49233);
or UO_1847 (O_1847,N_49623,N_49319);
xnor UO_1848 (O_1848,N_49000,N_47893);
nand UO_1849 (O_1849,N_49334,N_47785);
or UO_1850 (O_1850,N_47799,N_48669);
and UO_1851 (O_1851,N_49579,N_49928);
nand UO_1852 (O_1852,N_49113,N_49411);
xnor UO_1853 (O_1853,N_49001,N_47539);
xor UO_1854 (O_1854,N_48131,N_48229);
nand UO_1855 (O_1855,N_48752,N_47659);
or UO_1856 (O_1856,N_49345,N_48649);
xor UO_1857 (O_1857,N_49459,N_49946);
xnor UO_1858 (O_1858,N_49149,N_49561);
xnor UO_1859 (O_1859,N_47940,N_47738);
or UO_1860 (O_1860,N_49133,N_49076);
and UO_1861 (O_1861,N_48366,N_49617);
or UO_1862 (O_1862,N_48976,N_47703);
xor UO_1863 (O_1863,N_49559,N_48992);
and UO_1864 (O_1864,N_48229,N_47668);
xor UO_1865 (O_1865,N_48559,N_47833);
or UO_1866 (O_1866,N_48590,N_49834);
nand UO_1867 (O_1867,N_49487,N_49299);
xnor UO_1868 (O_1868,N_48732,N_47516);
and UO_1869 (O_1869,N_48072,N_47576);
xor UO_1870 (O_1870,N_48670,N_47521);
nor UO_1871 (O_1871,N_48618,N_48307);
xor UO_1872 (O_1872,N_49311,N_48546);
nor UO_1873 (O_1873,N_47715,N_48012);
nor UO_1874 (O_1874,N_47856,N_48376);
and UO_1875 (O_1875,N_48633,N_49238);
and UO_1876 (O_1876,N_47523,N_49004);
xor UO_1877 (O_1877,N_49865,N_47833);
nand UO_1878 (O_1878,N_48962,N_49512);
and UO_1879 (O_1879,N_49601,N_48039);
and UO_1880 (O_1880,N_48956,N_49596);
and UO_1881 (O_1881,N_48931,N_49915);
nand UO_1882 (O_1882,N_47513,N_49802);
and UO_1883 (O_1883,N_48845,N_48096);
nor UO_1884 (O_1884,N_47544,N_48144);
and UO_1885 (O_1885,N_49157,N_48735);
nor UO_1886 (O_1886,N_48042,N_47970);
nand UO_1887 (O_1887,N_47804,N_48061);
nor UO_1888 (O_1888,N_48149,N_48647);
nor UO_1889 (O_1889,N_48824,N_47648);
nor UO_1890 (O_1890,N_47554,N_49260);
xor UO_1891 (O_1891,N_48563,N_47565);
and UO_1892 (O_1892,N_48157,N_47879);
nor UO_1893 (O_1893,N_47882,N_49228);
and UO_1894 (O_1894,N_49868,N_47891);
or UO_1895 (O_1895,N_48060,N_49434);
nand UO_1896 (O_1896,N_49216,N_48458);
nor UO_1897 (O_1897,N_49314,N_49126);
or UO_1898 (O_1898,N_48721,N_47644);
xnor UO_1899 (O_1899,N_48778,N_48869);
and UO_1900 (O_1900,N_49267,N_49095);
and UO_1901 (O_1901,N_49291,N_49160);
nand UO_1902 (O_1902,N_49363,N_49964);
xor UO_1903 (O_1903,N_48799,N_49561);
or UO_1904 (O_1904,N_48633,N_49638);
nand UO_1905 (O_1905,N_49539,N_48892);
nor UO_1906 (O_1906,N_49534,N_49620);
nand UO_1907 (O_1907,N_49738,N_47823);
xor UO_1908 (O_1908,N_47548,N_47922);
or UO_1909 (O_1909,N_49744,N_48636);
xor UO_1910 (O_1910,N_49853,N_47796);
nor UO_1911 (O_1911,N_47521,N_47651);
nand UO_1912 (O_1912,N_49676,N_49542);
xnor UO_1913 (O_1913,N_48696,N_49198);
and UO_1914 (O_1914,N_48384,N_49407);
xor UO_1915 (O_1915,N_48944,N_49392);
or UO_1916 (O_1916,N_49317,N_47955);
or UO_1917 (O_1917,N_48374,N_48000);
and UO_1918 (O_1918,N_48655,N_47528);
xnor UO_1919 (O_1919,N_48446,N_49869);
xor UO_1920 (O_1920,N_49560,N_49932);
nor UO_1921 (O_1921,N_48184,N_47895);
xor UO_1922 (O_1922,N_48054,N_48601);
xnor UO_1923 (O_1923,N_47666,N_48329);
and UO_1924 (O_1924,N_48613,N_49840);
nand UO_1925 (O_1925,N_47995,N_49130);
nor UO_1926 (O_1926,N_48602,N_48863);
and UO_1927 (O_1927,N_48875,N_48390);
xnor UO_1928 (O_1928,N_48683,N_48070);
and UO_1929 (O_1929,N_48011,N_47555);
nor UO_1930 (O_1930,N_48211,N_49039);
xnor UO_1931 (O_1931,N_49586,N_47727);
xor UO_1932 (O_1932,N_48269,N_48135);
nand UO_1933 (O_1933,N_48945,N_49742);
xor UO_1934 (O_1934,N_48281,N_48392);
xnor UO_1935 (O_1935,N_49620,N_49377);
nand UO_1936 (O_1936,N_48316,N_47742);
or UO_1937 (O_1937,N_49292,N_48987);
nor UO_1938 (O_1938,N_49136,N_48056);
nor UO_1939 (O_1939,N_49531,N_48536);
and UO_1940 (O_1940,N_48318,N_48869);
nand UO_1941 (O_1941,N_49785,N_48315);
nor UO_1942 (O_1942,N_47651,N_47798);
nor UO_1943 (O_1943,N_48494,N_47775);
or UO_1944 (O_1944,N_49881,N_47990);
or UO_1945 (O_1945,N_49195,N_49095);
nor UO_1946 (O_1946,N_48085,N_48122);
and UO_1947 (O_1947,N_47957,N_49433);
or UO_1948 (O_1948,N_49865,N_47807);
and UO_1949 (O_1949,N_49996,N_49932);
nor UO_1950 (O_1950,N_47507,N_49660);
nand UO_1951 (O_1951,N_49619,N_49876);
nor UO_1952 (O_1952,N_47649,N_48361);
nor UO_1953 (O_1953,N_47668,N_49950);
nand UO_1954 (O_1954,N_47589,N_47947);
and UO_1955 (O_1955,N_49593,N_49301);
nor UO_1956 (O_1956,N_49810,N_48657);
and UO_1957 (O_1957,N_48812,N_49103);
xor UO_1958 (O_1958,N_49040,N_48978);
nand UO_1959 (O_1959,N_47873,N_49567);
nor UO_1960 (O_1960,N_49029,N_47681);
nor UO_1961 (O_1961,N_47759,N_49740);
or UO_1962 (O_1962,N_49664,N_47940);
xnor UO_1963 (O_1963,N_48012,N_49498);
nor UO_1964 (O_1964,N_48095,N_49496);
nand UO_1965 (O_1965,N_48350,N_47890);
and UO_1966 (O_1966,N_48646,N_49924);
xor UO_1967 (O_1967,N_49670,N_47757);
and UO_1968 (O_1968,N_47769,N_48632);
nor UO_1969 (O_1969,N_49947,N_49510);
or UO_1970 (O_1970,N_48709,N_48908);
and UO_1971 (O_1971,N_47720,N_48749);
or UO_1972 (O_1972,N_49247,N_49099);
xnor UO_1973 (O_1973,N_49064,N_48804);
or UO_1974 (O_1974,N_47663,N_49638);
and UO_1975 (O_1975,N_49669,N_49713);
or UO_1976 (O_1976,N_49850,N_49500);
or UO_1977 (O_1977,N_49450,N_47595);
and UO_1978 (O_1978,N_49985,N_48383);
and UO_1979 (O_1979,N_49815,N_49834);
or UO_1980 (O_1980,N_49130,N_48652);
or UO_1981 (O_1981,N_47970,N_48914);
and UO_1982 (O_1982,N_48445,N_49441);
xor UO_1983 (O_1983,N_47794,N_48621);
xor UO_1984 (O_1984,N_48624,N_49983);
and UO_1985 (O_1985,N_49925,N_49890);
nor UO_1986 (O_1986,N_49225,N_48534);
nand UO_1987 (O_1987,N_48714,N_49077);
and UO_1988 (O_1988,N_48361,N_49598);
or UO_1989 (O_1989,N_49258,N_48445);
or UO_1990 (O_1990,N_49379,N_48500);
nand UO_1991 (O_1991,N_49826,N_49707);
or UO_1992 (O_1992,N_47850,N_49544);
or UO_1993 (O_1993,N_49024,N_47964);
or UO_1994 (O_1994,N_48854,N_47903);
xor UO_1995 (O_1995,N_48197,N_48717);
xor UO_1996 (O_1996,N_47958,N_48701);
nand UO_1997 (O_1997,N_48589,N_49894);
and UO_1998 (O_1998,N_48586,N_48175);
xor UO_1999 (O_1999,N_49440,N_48583);
xnor UO_2000 (O_2000,N_48101,N_47528);
nor UO_2001 (O_2001,N_47853,N_49768);
xnor UO_2002 (O_2002,N_48414,N_47904);
xnor UO_2003 (O_2003,N_48088,N_48196);
nor UO_2004 (O_2004,N_48462,N_47556);
nand UO_2005 (O_2005,N_48035,N_47837);
nor UO_2006 (O_2006,N_49677,N_49071);
and UO_2007 (O_2007,N_48500,N_48395);
nand UO_2008 (O_2008,N_48843,N_48739);
nor UO_2009 (O_2009,N_49435,N_48826);
nor UO_2010 (O_2010,N_47705,N_49691);
xor UO_2011 (O_2011,N_48710,N_48592);
nor UO_2012 (O_2012,N_47667,N_49627);
nor UO_2013 (O_2013,N_48607,N_48542);
xor UO_2014 (O_2014,N_48569,N_49159);
nor UO_2015 (O_2015,N_48588,N_49754);
xor UO_2016 (O_2016,N_49411,N_48525);
or UO_2017 (O_2017,N_47802,N_49328);
nand UO_2018 (O_2018,N_48038,N_48223);
or UO_2019 (O_2019,N_49566,N_49347);
nor UO_2020 (O_2020,N_48457,N_49245);
or UO_2021 (O_2021,N_49385,N_49646);
or UO_2022 (O_2022,N_48814,N_49569);
or UO_2023 (O_2023,N_49206,N_48968);
or UO_2024 (O_2024,N_48711,N_47653);
xnor UO_2025 (O_2025,N_48051,N_48768);
nor UO_2026 (O_2026,N_49325,N_49024);
and UO_2027 (O_2027,N_49130,N_48217);
nand UO_2028 (O_2028,N_48952,N_48090);
or UO_2029 (O_2029,N_48211,N_48170);
nand UO_2030 (O_2030,N_48454,N_49995);
nand UO_2031 (O_2031,N_47756,N_48219);
and UO_2032 (O_2032,N_47566,N_49656);
nor UO_2033 (O_2033,N_47518,N_48271);
or UO_2034 (O_2034,N_48571,N_47809);
nand UO_2035 (O_2035,N_47655,N_48779);
nor UO_2036 (O_2036,N_49335,N_48830);
or UO_2037 (O_2037,N_48770,N_48741);
nand UO_2038 (O_2038,N_48768,N_49332);
nand UO_2039 (O_2039,N_49955,N_48197);
xor UO_2040 (O_2040,N_49523,N_49276);
xor UO_2041 (O_2041,N_48829,N_48894);
nor UO_2042 (O_2042,N_49127,N_49678);
xor UO_2043 (O_2043,N_49185,N_47550);
and UO_2044 (O_2044,N_47800,N_48598);
nand UO_2045 (O_2045,N_48207,N_47960);
xnor UO_2046 (O_2046,N_49230,N_48719);
nand UO_2047 (O_2047,N_49093,N_49129);
or UO_2048 (O_2048,N_48054,N_48069);
xor UO_2049 (O_2049,N_48391,N_49599);
xnor UO_2050 (O_2050,N_49309,N_49724);
nor UO_2051 (O_2051,N_47639,N_49667);
or UO_2052 (O_2052,N_49387,N_47842);
and UO_2053 (O_2053,N_49594,N_49891);
xnor UO_2054 (O_2054,N_48808,N_49864);
or UO_2055 (O_2055,N_49548,N_48127);
xnor UO_2056 (O_2056,N_47829,N_48595);
or UO_2057 (O_2057,N_47998,N_48782);
and UO_2058 (O_2058,N_49972,N_49363);
nand UO_2059 (O_2059,N_48632,N_47725);
xor UO_2060 (O_2060,N_48673,N_47811);
or UO_2061 (O_2061,N_48199,N_47643);
nor UO_2062 (O_2062,N_48744,N_47530);
nor UO_2063 (O_2063,N_47643,N_48678);
or UO_2064 (O_2064,N_49430,N_48087);
or UO_2065 (O_2065,N_47685,N_48266);
xnor UO_2066 (O_2066,N_47966,N_48093);
or UO_2067 (O_2067,N_47928,N_48512);
and UO_2068 (O_2068,N_47562,N_48049);
or UO_2069 (O_2069,N_49264,N_48268);
nor UO_2070 (O_2070,N_49840,N_49243);
and UO_2071 (O_2071,N_49790,N_49893);
nand UO_2072 (O_2072,N_49141,N_47629);
and UO_2073 (O_2073,N_48638,N_47950);
nor UO_2074 (O_2074,N_47880,N_47843);
and UO_2075 (O_2075,N_47643,N_49381);
nand UO_2076 (O_2076,N_48385,N_47524);
xnor UO_2077 (O_2077,N_49355,N_48090);
nand UO_2078 (O_2078,N_48166,N_49599);
or UO_2079 (O_2079,N_47673,N_47866);
xnor UO_2080 (O_2080,N_49239,N_47549);
or UO_2081 (O_2081,N_48739,N_49582);
xnor UO_2082 (O_2082,N_49643,N_48607);
xor UO_2083 (O_2083,N_48654,N_47750);
and UO_2084 (O_2084,N_49453,N_49837);
xnor UO_2085 (O_2085,N_48867,N_49479);
nor UO_2086 (O_2086,N_47762,N_48452);
and UO_2087 (O_2087,N_49692,N_48845);
nand UO_2088 (O_2088,N_48872,N_49582);
xnor UO_2089 (O_2089,N_47687,N_49216);
or UO_2090 (O_2090,N_47577,N_47902);
nor UO_2091 (O_2091,N_47839,N_48517);
xor UO_2092 (O_2092,N_49188,N_48584);
or UO_2093 (O_2093,N_48984,N_49082);
and UO_2094 (O_2094,N_47721,N_48307);
and UO_2095 (O_2095,N_48434,N_48002);
or UO_2096 (O_2096,N_48181,N_49153);
nor UO_2097 (O_2097,N_48852,N_49586);
and UO_2098 (O_2098,N_49608,N_48280);
nor UO_2099 (O_2099,N_48062,N_47926);
nand UO_2100 (O_2100,N_49831,N_47951);
nand UO_2101 (O_2101,N_47620,N_49702);
or UO_2102 (O_2102,N_49213,N_49068);
xnor UO_2103 (O_2103,N_49129,N_49873);
and UO_2104 (O_2104,N_47930,N_48681);
or UO_2105 (O_2105,N_49619,N_48464);
and UO_2106 (O_2106,N_49134,N_48097);
nor UO_2107 (O_2107,N_48053,N_48845);
xor UO_2108 (O_2108,N_47795,N_49570);
or UO_2109 (O_2109,N_49314,N_49018);
and UO_2110 (O_2110,N_49547,N_47568);
or UO_2111 (O_2111,N_49702,N_47817);
or UO_2112 (O_2112,N_47656,N_47710);
nand UO_2113 (O_2113,N_49202,N_47765);
and UO_2114 (O_2114,N_48341,N_48086);
xnor UO_2115 (O_2115,N_49980,N_47979);
xnor UO_2116 (O_2116,N_48623,N_48236);
nand UO_2117 (O_2117,N_49137,N_48538);
nand UO_2118 (O_2118,N_49909,N_48887);
or UO_2119 (O_2119,N_48686,N_48742);
or UO_2120 (O_2120,N_47850,N_48859);
nand UO_2121 (O_2121,N_48864,N_48350);
xor UO_2122 (O_2122,N_48525,N_47937);
or UO_2123 (O_2123,N_48728,N_49257);
nand UO_2124 (O_2124,N_48131,N_48607);
nor UO_2125 (O_2125,N_48099,N_48530);
nand UO_2126 (O_2126,N_49544,N_49921);
and UO_2127 (O_2127,N_47864,N_49162);
and UO_2128 (O_2128,N_47937,N_48856);
nor UO_2129 (O_2129,N_49582,N_49180);
or UO_2130 (O_2130,N_48546,N_48515);
nor UO_2131 (O_2131,N_49854,N_49426);
and UO_2132 (O_2132,N_49842,N_47929);
nor UO_2133 (O_2133,N_48973,N_48593);
and UO_2134 (O_2134,N_47689,N_49349);
and UO_2135 (O_2135,N_49918,N_49106);
xnor UO_2136 (O_2136,N_49841,N_48888);
nand UO_2137 (O_2137,N_49554,N_48309);
nor UO_2138 (O_2138,N_48906,N_48529);
and UO_2139 (O_2139,N_49497,N_48567);
and UO_2140 (O_2140,N_48947,N_48057);
nand UO_2141 (O_2141,N_49487,N_49262);
and UO_2142 (O_2142,N_49308,N_49841);
nor UO_2143 (O_2143,N_49468,N_49915);
nor UO_2144 (O_2144,N_49188,N_49014);
or UO_2145 (O_2145,N_47942,N_47550);
nand UO_2146 (O_2146,N_47676,N_48303);
nand UO_2147 (O_2147,N_49226,N_49225);
and UO_2148 (O_2148,N_48326,N_49726);
and UO_2149 (O_2149,N_48626,N_49191);
nand UO_2150 (O_2150,N_48212,N_48234);
xor UO_2151 (O_2151,N_48288,N_47775);
nand UO_2152 (O_2152,N_49160,N_49214);
or UO_2153 (O_2153,N_49324,N_49105);
xor UO_2154 (O_2154,N_48160,N_48135);
xor UO_2155 (O_2155,N_48252,N_48160);
nand UO_2156 (O_2156,N_48522,N_47620);
nor UO_2157 (O_2157,N_49786,N_49346);
nor UO_2158 (O_2158,N_48729,N_48996);
nor UO_2159 (O_2159,N_48200,N_49572);
or UO_2160 (O_2160,N_49002,N_49851);
nor UO_2161 (O_2161,N_49944,N_48977);
nand UO_2162 (O_2162,N_47748,N_48051);
xnor UO_2163 (O_2163,N_48325,N_49507);
nor UO_2164 (O_2164,N_48888,N_47742);
nor UO_2165 (O_2165,N_49866,N_49148);
nor UO_2166 (O_2166,N_47591,N_48908);
and UO_2167 (O_2167,N_47712,N_49386);
nand UO_2168 (O_2168,N_49971,N_48706);
xnor UO_2169 (O_2169,N_49803,N_49739);
xor UO_2170 (O_2170,N_47793,N_49985);
xor UO_2171 (O_2171,N_48400,N_47779);
nand UO_2172 (O_2172,N_48817,N_49355);
or UO_2173 (O_2173,N_48304,N_49112);
xor UO_2174 (O_2174,N_48395,N_47907);
nor UO_2175 (O_2175,N_48388,N_49332);
xnor UO_2176 (O_2176,N_47552,N_47567);
xnor UO_2177 (O_2177,N_49436,N_49081);
and UO_2178 (O_2178,N_48057,N_49450);
and UO_2179 (O_2179,N_47989,N_48171);
nor UO_2180 (O_2180,N_48333,N_49847);
nor UO_2181 (O_2181,N_48602,N_47703);
nand UO_2182 (O_2182,N_48509,N_48874);
or UO_2183 (O_2183,N_47900,N_48900);
or UO_2184 (O_2184,N_49777,N_48548);
or UO_2185 (O_2185,N_49195,N_49582);
nand UO_2186 (O_2186,N_49284,N_47535);
or UO_2187 (O_2187,N_49472,N_48816);
xor UO_2188 (O_2188,N_47715,N_49704);
and UO_2189 (O_2189,N_47727,N_48528);
and UO_2190 (O_2190,N_49358,N_48791);
nor UO_2191 (O_2191,N_48719,N_47986);
and UO_2192 (O_2192,N_48413,N_48292);
nor UO_2193 (O_2193,N_47812,N_47984);
and UO_2194 (O_2194,N_49022,N_49977);
or UO_2195 (O_2195,N_48710,N_49376);
and UO_2196 (O_2196,N_48466,N_47845);
nor UO_2197 (O_2197,N_49011,N_48389);
or UO_2198 (O_2198,N_49712,N_48096);
nand UO_2199 (O_2199,N_49446,N_48709);
xnor UO_2200 (O_2200,N_49637,N_47564);
nand UO_2201 (O_2201,N_48518,N_49363);
and UO_2202 (O_2202,N_47558,N_48608);
and UO_2203 (O_2203,N_48491,N_48224);
or UO_2204 (O_2204,N_48528,N_49926);
xnor UO_2205 (O_2205,N_48429,N_49798);
or UO_2206 (O_2206,N_48141,N_47839);
or UO_2207 (O_2207,N_48321,N_48455);
or UO_2208 (O_2208,N_49716,N_48916);
nand UO_2209 (O_2209,N_49204,N_49625);
nand UO_2210 (O_2210,N_49817,N_49914);
and UO_2211 (O_2211,N_49028,N_47765);
and UO_2212 (O_2212,N_49507,N_48151);
or UO_2213 (O_2213,N_47927,N_48981);
xnor UO_2214 (O_2214,N_48606,N_48710);
nand UO_2215 (O_2215,N_48641,N_49254);
nor UO_2216 (O_2216,N_47710,N_48741);
xnor UO_2217 (O_2217,N_48093,N_47630);
and UO_2218 (O_2218,N_48705,N_49787);
nor UO_2219 (O_2219,N_49948,N_49937);
or UO_2220 (O_2220,N_48352,N_47822);
nor UO_2221 (O_2221,N_47778,N_48595);
nor UO_2222 (O_2222,N_48799,N_48986);
nand UO_2223 (O_2223,N_49004,N_48696);
or UO_2224 (O_2224,N_48675,N_49148);
nand UO_2225 (O_2225,N_48880,N_47539);
nor UO_2226 (O_2226,N_48046,N_48235);
xor UO_2227 (O_2227,N_47916,N_47668);
nand UO_2228 (O_2228,N_47560,N_47655);
xor UO_2229 (O_2229,N_48417,N_48307);
nand UO_2230 (O_2230,N_47610,N_49398);
xor UO_2231 (O_2231,N_48109,N_49661);
and UO_2232 (O_2232,N_49818,N_49987);
nand UO_2233 (O_2233,N_47837,N_47528);
nand UO_2234 (O_2234,N_49499,N_48392);
and UO_2235 (O_2235,N_49718,N_49825);
or UO_2236 (O_2236,N_49108,N_49330);
nand UO_2237 (O_2237,N_49320,N_49652);
and UO_2238 (O_2238,N_49445,N_48256);
and UO_2239 (O_2239,N_49602,N_49098);
and UO_2240 (O_2240,N_49341,N_49066);
and UO_2241 (O_2241,N_49423,N_49097);
or UO_2242 (O_2242,N_47838,N_48736);
nand UO_2243 (O_2243,N_49708,N_48705);
or UO_2244 (O_2244,N_47893,N_48173);
nor UO_2245 (O_2245,N_49163,N_49090);
and UO_2246 (O_2246,N_48945,N_47506);
and UO_2247 (O_2247,N_48595,N_49180);
nor UO_2248 (O_2248,N_49367,N_49354);
nor UO_2249 (O_2249,N_48438,N_47891);
nand UO_2250 (O_2250,N_49627,N_48413);
and UO_2251 (O_2251,N_48622,N_49942);
and UO_2252 (O_2252,N_48804,N_48683);
and UO_2253 (O_2253,N_48800,N_49133);
and UO_2254 (O_2254,N_49482,N_47769);
nor UO_2255 (O_2255,N_48862,N_48543);
and UO_2256 (O_2256,N_49435,N_49114);
xnor UO_2257 (O_2257,N_48112,N_49548);
xor UO_2258 (O_2258,N_49711,N_48099);
nor UO_2259 (O_2259,N_48747,N_49997);
or UO_2260 (O_2260,N_48374,N_49377);
xor UO_2261 (O_2261,N_48775,N_49299);
nor UO_2262 (O_2262,N_48939,N_49027);
or UO_2263 (O_2263,N_48353,N_48327);
or UO_2264 (O_2264,N_48320,N_49112);
nor UO_2265 (O_2265,N_49146,N_47928);
xor UO_2266 (O_2266,N_49149,N_49086);
and UO_2267 (O_2267,N_49033,N_49003);
nand UO_2268 (O_2268,N_49640,N_48681);
nor UO_2269 (O_2269,N_48562,N_48820);
or UO_2270 (O_2270,N_47645,N_47694);
and UO_2271 (O_2271,N_48028,N_48036);
xor UO_2272 (O_2272,N_48808,N_47934);
and UO_2273 (O_2273,N_48547,N_48733);
xor UO_2274 (O_2274,N_48259,N_48134);
and UO_2275 (O_2275,N_48707,N_49913);
and UO_2276 (O_2276,N_48000,N_47796);
or UO_2277 (O_2277,N_48375,N_48307);
and UO_2278 (O_2278,N_48484,N_48500);
xnor UO_2279 (O_2279,N_49970,N_49458);
or UO_2280 (O_2280,N_48207,N_47735);
or UO_2281 (O_2281,N_49554,N_49831);
xor UO_2282 (O_2282,N_49615,N_48118);
xnor UO_2283 (O_2283,N_48819,N_48559);
or UO_2284 (O_2284,N_48675,N_49923);
nand UO_2285 (O_2285,N_48439,N_49833);
and UO_2286 (O_2286,N_48393,N_49943);
and UO_2287 (O_2287,N_48459,N_48583);
or UO_2288 (O_2288,N_47946,N_48928);
nor UO_2289 (O_2289,N_49507,N_48747);
or UO_2290 (O_2290,N_49620,N_47887);
nand UO_2291 (O_2291,N_49685,N_47947);
nand UO_2292 (O_2292,N_47760,N_48850);
xnor UO_2293 (O_2293,N_47853,N_48781);
and UO_2294 (O_2294,N_48671,N_48021);
nand UO_2295 (O_2295,N_49366,N_47673);
nor UO_2296 (O_2296,N_48448,N_49748);
or UO_2297 (O_2297,N_49851,N_49181);
nand UO_2298 (O_2298,N_48371,N_48862);
or UO_2299 (O_2299,N_48668,N_49058);
or UO_2300 (O_2300,N_48715,N_47611);
and UO_2301 (O_2301,N_48241,N_49838);
xnor UO_2302 (O_2302,N_47947,N_49089);
and UO_2303 (O_2303,N_49979,N_49124);
xnor UO_2304 (O_2304,N_47802,N_49611);
xnor UO_2305 (O_2305,N_49599,N_49204);
and UO_2306 (O_2306,N_47604,N_49509);
nand UO_2307 (O_2307,N_49445,N_48085);
or UO_2308 (O_2308,N_48562,N_49667);
or UO_2309 (O_2309,N_49204,N_47701);
or UO_2310 (O_2310,N_48863,N_47755);
nor UO_2311 (O_2311,N_49619,N_48349);
and UO_2312 (O_2312,N_47977,N_47765);
nand UO_2313 (O_2313,N_48208,N_48376);
or UO_2314 (O_2314,N_49534,N_48393);
or UO_2315 (O_2315,N_49942,N_48754);
nand UO_2316 (O_2316,N_48974,N_48615);
or UO_2317 (O_2317,N_47611,N_49638);
nor UO_2318 (O_2318,N_49884,N_49063);
nand UO_2319 (O_2319,N_48821,N_48019);
or UO_2320 (O_2320,N_48407,N_49737);
nand UO_2321 (O_2321,N_49479,N_49556);
or UO_2322 (O_2322,N_48678,N_49202);
xor UO_2323 (O_2323,N_47832,N_47510);
xnor UO_2324 (O_2324,N_49092,N_48254);
or UO_2325 (O_2325,N_48842,N_49389);
or UO_2326 (O_2326,N_48274,N_49046);
and UO_2327 (O_2327,N_49049,N_48001);
nor UO_2328 (O_2328,N_49867,N_48229);
nor UO_2329 (O_2329,N_47631,N_47581);
and UO_2330 (O_2330,N_49977,N_48024);
xnor UO_2331 (O_2331,N_48046,N_49614);
and UO_2332 (O_2332,N_48330,N_48599);
or UO_2333 (O_2333,N_48463,N_48508);
xor UO_2334 (O_2334,N_48263,N_47774);
nand UO_2335 (O_2335,N_48561,N_49212);
or UO_2336 (O_2336,N_48305,N_49398);
xnor UO_2337 (O_2337,N_48310,N_47960);
or UO_2338 (O_2338,N_47833,N_47964);
xnor UO_2339 (O_2339,N_48133,N_49596);
or UO_2340 (O_2340,N_49301,N_48388);
nand UO_2341 (O_2341,N_49627,N_49848);
xnor UO_2342 (O_2342,N_48001,N_48374);
or UO_2343 (O_2343,N_49532,N_49164);
and UO_2344 (O_2344,N_48375,N_49208);
nor UO_2345 (O_2345,N_48700,N_49384);
or UO_2346 (O_2346,N_48146,N_49095);
or UO_2347 (O_2347,N_49420,N_47735);
and UO_2348 (O_2348,N_49589,N_49612);
nand UO_2349 (O_2349,N_49056,N_48227);
xnor UO_2350 (O_2350,N_47664,N_48805);
and UO_2351 (O_2351,N_48370,N_49388);
nor UO_2352 (O_2352,N_47763,N_47657);
xor UO_2353 (O_2353,N_48329,N_48399);
xnor UO_2354 (O_2354,N_48666,N_47517);
nor UO_2355 (O_2355,N_49878,N_49277);
xor UO_2356 (O_2356,N_49996,N_48964);
xnor UO_2357 (O_2357,N_49653,N_48067);
nand UO_2358 (O_2358,N_47693,N_49933);
or UO_2359 (O_2359,N_47972,N_49598);
xor UO_2360 (O_2360,N_48478,N_48342);
and UO_2361 (O_2361,N_49636,N_48643);
nor UO_2362 (O_2362,N_47810,N_48331);
and UO_2363 (O_2363,N_49052,N_48876);
xor UO_2364 (O_2364,N_49586,N_47848);
and UO_2365 (O_2365,N_48423,N_47555);
or UO_2366 (O_2366,N_49263,N_48702);
or UO_2367 (O_2367,N_49292,N_49851);
nor UO_2368 (O_2368,N_49391,N_48405);
nand UO_2369 (O_2369,N_48636,N_49342);
xnor UO_2370 (O_2370,N_49192,N_47745);
xor UO_2371 (O_2371,N_49754,N_48989);
and UO_2372 (O_2372,N_49933,N_47587);
or UO_2373 (O_2373,N_48887,N_47992);
nor UO_2374 (O_2374,N_48779,N_48837);
nand UO_2375 (O_2375,N_48567,N_47552);
nor UO_2376 (O_2376,N_49168,N_48415);
or UO_2377 (O_2377,N_48799,N_49569);
nor UO_2378 (O_2378,N_48187,N_48665);
and UO_2379 (O_2379,N_48978,N_49612);
or UO_2380 (O_2380,N_49806,N_48220);
nor UO_2381 (O_2381,N_48105,N_47846);
and UO_2382 (O_2382,N_47764,N_48825);
nand UO_2383 (O_2383,N_47983,N_49784);
or UO_2384 (O_2384,N_49821,N_49957);
nor UO_2385 (O_2385,N_49763,N_48493);
or UO_2386 (O_2386,N_49371,N_49054);
nand UO_2387 (O_2387,N_48270,N_49778);
xor UO_2388 (O_2388,N_47991,N_48688);
xor UO_2389 (O_2389,N_49926,N_47736);
nand UO_2390 (O_2390,N_48553,N_48483);
xnor UO_2391 (O_2391,N_49504,N_48589);
or UO_2392 (O_2392,N_48381,N_49127);
or UO_2393 (O_2393,N_49392,N_49830);
and UO_2394 (O_2394,N_48176,N_49078);
and UO_2395 (O_2395,N_48150,N_49546);
and UO_2396 (O_2396,N_49911,N_48573);
nand UO_2397 (O_2397,N_49376,N_49256);
nand UO_2398 (O_2398,N_48865,N_49183);
nor UO_2399 (O_2399,N_47667,N_49155);
nor UO_2400 (O_2400,N_48817,N_47649);
nor UO_2401 (O_2401,N_49667,N_49031);
and UO_2402 (O_2402,N_49239,N_48819);
and UO_2403 (O_2403,N_49027,N_49717);
or UO_2404 (O_2404,N_49816,N_49465);
nand UO_2405 (O_2405,N_49369,N_47852);
and UO_2406 (O_2406,N_48893,N_49191);
and UO_2407 (O_2407,N_48925,N_48329);
and UO_2408 (O_2408,N_49576,N_48129);
or UO_2409 (O_2409,N_47950,N_47875);
or UO_2410 (O_2410,N_49471,N_48136);
nor UO_2411 (O_2411,N_49773,N_48856);
and UO_2412 (O_2412,N_48541,N_47969);
or UO_2413 (O_2413,N_49843,N_49549);
and UO_2414 (O_2414,N_49222,N_48465);
nor UO_2415 (O_2415,N_48216,N_49815);
nor UO_2416 (O_2416,N_48207,N_48565);
xor UO_2417 (O_2417,N_49369,N_49115);
or UO_2418 (O_2418,N_49002,N_49019);
and UO_2419 (O_2419,N_48534,N_48850);
nand UO_2420 (O_2420,N_48097,N_48078);
and UO_2421 (O_2421,N_49019,N_48065);
xor UO_2422 (O_2422,N_47832,N_47656);
nand UO_2423 (O_2423,N_49264,N_49236);
xnor UO_2424 (O_2424,N_48663,N_48259);
or UO_2425 (O_2425,N_49920,N_47955);
or UO_2426 (O_2426,N_49000,N_49110);
or UO_2427 (O_2427,N_49145,N_47660);
and UO_2428 (O_2428,N_49281,N_48674);
xnor UO_2429 (O_2429,N_48366,N_48368);
and UO_2430 (O_2430,N_48385,N_48126);
nor UO_2431 (O_2431,N_49884,N_49589);
xnor UO_2432 (O_2432,N_48715,N_49797);
nor UO_2433 (O_2433,N_47914,N_48940);
and UO_2434 (O_2434,N_47783,N_48403);
nand UO_2435 (O_2435,N_49624,N_47559);
or UO_2436 (O_2436,N_49585,N_49990);
nor UO_2437 (O_2437,N_48871,N_48088);
xor UO_2438 (O_2438,N_49038,N_48431);
xor UO_2439 (O_2439,N_48952,N_49579);
xnor UO_2440 (O_2440,N_47734,N_48572);
or UO_2441 (O_2441,N_48441,N_48318);
or UO_2442 (O_2442,N_48583,N_47739);
and UO_2443 (O_2443,N_49601,N_48210);
nor UO_2444 (O_2444,N_49355,N_47962);
nor UO_2445 (O_2445,N_48573,N_47909);
and UO_2446 (O_2446,N_47931,N_48765);
or UO_2447 (O_2447,N_48529,N_48010);
xor UO_2448 (O_2448,N_48776,N_48260);
xnor UO_2449 (O_2449,N_49767,N_49665);
nor UO_2450 (O_2450,N_48195,N_48567);
and UO_2451 (O_2451,N_47866,N_49082);
and UO_2452 (O_2452,N_47675,N_49751);
and UO_2453 (O_2453,N_49544,N_49018);
xnor UO_2454 (O_2454,N_48122,N_49959);
or UO_2455 (O_2455,N_48269,N_48713);
and UO_2456 (O_2456,N_49553,N_49577);
xor UO_2457 (O_2457,N_48969,N_49543);
nand UO_2458 (O_2458,N_47599,N_47758);
nand UO_2459 (O_2459,N_47980,N_49731);
nor UO_2460 (O_2460,N_48165,N_49437);
and UO_2461 (O_2461,N_48568,N_48725);
xor UO_2462 (O_2462,N_47973,N_49614);
nor UO_2463 (O_2463,N_47955,N_48496);
nand UO_2464 (O_2464,N_49785,N_48788);
and UO_2465 (O_2465,N_48583,N_48000);
xor UO_2466 (O_2466,N_48195,N_47694);
nor UO_2467 (O_2467,N_49345,N_47899);
or UO_2468 (O_2468,N_48736,N_48839);
nand UO_2469 (O_2469,N_48307,N_47947);
nor UO_2470 (O_2470,N_48006,N_49082);
nand UO_2471 (O_2471,N_47861,N_48275);
or UO_2472 (O_2472,N_49684,N_47830);
and UO_2473 (O_2473,N_48560,N_48514);
or UO_2474 (O_2474,N_47641,N_49769);
and UO_2475 (O_2475,N_48851,N_49493);
nand UO_2476 (O_2476,N_49299,N_48828);
xnor UO_2477 (O_2477,N_49476,N_47753);
nand UO_2478 (O_2478,N_48925,N_48090);
or UO_2479 (O_2479,N_47589,N_47571);
or UO_2480 (O_2480,N_47881,N_48189);
and UO_2481 (O_2481,N_49280,N_47943);
xor UO_2482 (O_2482,N_49315,N_48057);
or UO_2483 (O_2483,N_49248,N_48698);
xor UO_2484 (O_2484,N_48876,N_48210);
and UO_2485 (O_2485,N_49410,N_48806);
and UO_2486 (O_2486,N_47926,N_49695);
and UO_2487 (O_2487,N_49084,N_49676);
or UO_2488 (O_2488,N_49298,N_47801);
or UO_2489 (O_2489,N_47517,N_49099);
nor UO_2490 (O_2490,N_49671,N_48003);
nand UO_2491 (O_2491,N_49222,N_48408);
or UO_2492 (O_2492,N_48590,N_48848);
or UO_2493 (O_2493,N_49460,N_47590);
or UO_2494 (O_2494,N_49145,N_48388);
nor UO_2495 (O_2495,N_49009,N_47624);
nor UO_2496 (O_2496,N_48968,N_49997);
xor UO_2497 (O_2497,N_48069,N_49155);
or UO_2498 (O_2498,N_49621,N_47935);
nor UO_2499 (O_2499,N_48187,N_47617);
nand UO_2500 (O_2500,N_47995,N_49334);
xnor UO_2501 (O_2501,N_47880,N_48041);
xor UO_2502 (O_2502,N_49602,N_49542);
and UO_2503 (O_2503,N_48305,N_47925);
xor UO_2504 (O_2504,N_49473,N_48631);
xor UO_2505 (O_2505,N_48262,N_49452);
and UO_2506 (O_2506,N_49923,N_47703);
nor UO_2507 (O_2507,N_47580,N_48476);
xor UO_2508 (O_2508,N_49427,N_48205);
nor UO_2509 (O_2509,N_49134,N_48233);
nand UO_2510 (O_2510,N_47949,N_48216);
nor UO_2511 (O_2511,N_49338,N_48275);
and UO_2512 (O_2512,N_49506,N_47874);
nand UO_2513 (O_2513,N_48507,N_49322);
or UO_2514 (O_2514,N_48901,N_47795);
and UO_2515 (O_2515,N_48554,N_49467);
nor UO_2516 (O_2516,N_49860,N_48373);
nand UO_2517 (O_2517,N_49646,N_49207);
nor UO_2518 (O_2518,N_49085,N_49954);
nand UO_2519 (O_2519,N_48760,N_48255);
or UO_2520 (O_2520,N_47532,N_47990);
xnor UO_2521 (O_2521,N_49200,N_49749);
nand UO_2522 (O_2522,N_49011,N_48242);
and UO_2523 (O_2523,N_48794,N_49416);
nand UO_2524 (O_2524,N_47701,N_49373);
and UO_2525 (O_2525,N_49953,N_48226);
and UO_2526 (O_2526,N_48611,N_49336);
nand UO_2527 (O_2527,N_48976,N_48008);
or UO_2528 (O_2528,N_49720,N_48151);
or UO_2529 (O_2529,N_49303,N_49239);
or UO_2530 (O_2530,N_48483,N_49668);
nand UO_2531 (O_2531,N_49236,N_47505);
xnor UO_2532 (O_2532,N_48415,N_49184);
xnor UO_2533 (O_2533,N_49607,N_49425);
nor UO_2534 (O_2534,N_48718,N_49526);
nand UO_2535 (O_2535,N_48300,N_48312);
and UO_2536 (O_2536,N_49522,N_49090);
or UO_2537 (O_2537,N_48670,N_47927);
or UO_2538 (O_2538,N_47536,N_48457);
xor UO_2539 (O_2539,N_48847,N_49914);
nor UO_2540 (O_2540,N_49313,N_49123);
or UO_2541 (O_2541,N_48951,N_47975);
nor UO_2542 (O_2542,N_49621,N_48150);
xor UO_2543 (O_2543,N_49998,N_47783);
xor UO_2544 (O_2544,N_49664,N_49184);
nand UO_2545 (O_2545,N_47896,N_48243);
and UO_2546 (O_2546,N_48492,N_47600);
or UO_2547 (O_2547,N_48023,N_49199);
or UO_2548 (O_2548,N_49726,N_49724);
nor UO_2549 (O_2549,N_47507,N_49852);
or UO_2550 (O_2550,N_49185,N_49999);
nor UO_2551 (O_2551,N_48043,N_48507);
or UO_2552 (O_2552,N_48215,N_47848);
nor UO_2553 (O_2553,N_49595,N_48077);
nor UO_2554 (O_2554,N_49345,N_48852);
or UO_2555 (O_2555,N_49879,N_49598);
nand UO_2556 (O_2556,N_47860,N_48647);
nor UO_2557 (O_2557,N_48143,N_48033);
or UO_2558 (O_2558,N_49277,N_49513);
nor UO_2559 (O_2559,N_49350,N_49302);
xor UO_2560 (O_2560,N_47587,N_47800);
xnor UO_2561 (O_2561,N_48378,N_48117);
xor UO_2562 (O_2562,N_49009,N_47830);
and UO_2563 (O_2563,N_49527,N_48460);
or UO_2564 (O_2564,N_47863,N_49941);
xnor UO_2565 (O_2565,N_49725,N_49355);
xnor UO_2566 (O_2566,N_47728,N_48394);
xnor UO_2567 (O_2567,N_49537,N_47678);
nand UO_2568 (O_2568,N_49433,N_48649);
nand UO_2569 (O_2569,N_49100,N_48732);
or UO_2570 (O_2570,N_47656,N_48135);
and UO_2571 (O_2571,N_48966,N_49295);
nand UO_2572 (O_2572,N_48772,N_49283);
xor UO_2573 (O_2573,N_47562,N_49604);
or UO_2574 (O_2574,N_49074,N_48180);
nand UO_2575 (O_2575,N_48538,N_49122);
or UO_2576 (O_2576,N_49983,N_49273);
and UO_2577 (O_2577,N_49995,N_49859);
or UO_2578 (O_2578,N_49393,N_49216);
and UO_2579 (O_2579,N_49693,N_48979);
nor UO_2580 (O_2580,N_49740,N_48592);
or UO_2581 (O_2581,N_47920,N_48931);
nor UO_2582 (O_2582,N_47870,N_49136);
nor UO_2583 (O_2583,N_47905,N_49982);
and UO_2584 (O_2584,N_47585,N_49376);
and UO_2585 (O_2585,N_47549,N_48096);
nand UO_2586 (O_2586,N_48195,N_48060);
nand UO_2587 (O_2587,N_48261,N_47598);
nand UO_2588 (O_2588,N_47984,N_49468);
nand UO_2589 (O_2589,N_49167,N_48633);
xor UO_2590 (O_2590,N_49311,N_49475);
nand UO_2591 (O_2591,N_49515,N_48974);
xnor UO_2592 (O_2592,N_48104,N_48256);
or UO_2593 (O_2593,N_49101,N_48041);
or UO_2594 (O_2594,N_49520,N_48057);
nor UO_2595 (O_2595,N_49627,N_48532);
or UO_2596 (O_2596,N_48807,N_49175);
nand UO_2597 (O_2597,N_48012,N_49696);
nor UO_2598 (O_2598,N_47629,N_48219);
xnor UO_2599 (O_2599,N_48781,N_47640);
nor UO_2600 (O_2600,N_49560,N_48453);
nand UO_2601 (O_2601,N_48191,N_49327);
nor UO_2602 (O_2602,N_48558,N_48364);
xor UO_2603 (O_2603,N_48818,N_47713);
nand UO_2604 (O_2604,N_48694,N_49378);
nor UO_2605 (O_2605,N_47702,N_47877);
and UO_2606 (O_2606,N_48170,N_49737);
xor UO_2607 (O_2607,N_49097,N_48129);
xnor UO_2608 (O_2608,N_48186,N_49214);
nand UO_2609 (O_2609,N_49234,N_49688);
nand UO_2610 (O_2610,N_49175,N_49417);
nand UO_2611 (O_2611,N_49186,N_47621);
and UO_2612 (O_2612,N_48852,N_49564);
or UO_2613 (O_2613,N_49264,N_49306);
xor UO_2614 (O_2614,N_48998,N_49434);
xnor UO_2615 (O_2615,N_47839,N_49363);
xor UO_2616 (O_2616,N_48714,N_48441);
nor UO_2617 (O_2617,N_47718,N_47536);
nand UO_2618 (O_2618,N_47876,N_48843);
or UO_2619 (O_2619,N_48738,N_48771);
nor UO_2620 (O_2620,N_47996,N_48911);
nor UO_2621 (O_2621,N_49889,N_49466);
xnor UO_2622 (O_2622,N_48715,N_49275);
and UO_2623 (O_2623,N_48112,N_48778);
and UO_2624 (O_2624,N_49463,N_49544);
and UO_2625 (O_2625,N_49746,N_47766);
or UO_2626 (O_2626,N_48481,N_49490);
and UO_2627 (O_2627,N_48276,N_48770);
nor UO_2628 (O_2628,N_49952,N_49698);
and UO_2629 (O_2629,N_49866,N_49345);
nand UO_2630 (O_2630,N_49801,N_49543);
or UO_2631 (O_2631,N_48661,N_47503);
and UO_2632 (O_2632,N_48594,N_49872);
or UO_2633 (O_2633,N_49800,N_47561);
nor UO_2634 (O_2634,N_49749,N_48318);
xnor UO_2635 (O_2635,N_47925,N_48635);
xor UO_2636 (O_2636,N_48814,N_49615);
nand UO_2637 (O_2637,N_48305,N_48050);
and UO_2638 (O_2638,N_47648,N_47820);
nand UO_2639 (O_2639,N_48205,N_48077);
xnor UO_2640 (O_2640,N_47968,N_47690);
xnor UO_2641 (O_2641,N_47837,N_48081);
nor UO_2642 (O_2642,N_47961,N_49729);
xnor UO_2643 (O_2643,N_48263,N_47920);
xor UO_2644 (O_2644,N_49955,N_49599);
and UO_2645 (O_2645,N_47987,N_48462);
xor UO_2646 (O_2646,N_49680,N_49504);
nor UO_2647 (O_2647,N_49211,N_48672);
and UO_2648 (O_2648,N_48168,N_49505);
and UO_2649 (O_2649,N_47500,N_47538);
nand UO_2650 (O_2650,N_48087,N_49141);
nand UO_2651 (O_2651,N_48784,N_47788);
or UO_2652 (O_2652,N_47600,N_48751);
nor UO_2653 (O_2653,N_48568,N_48900);
and UO_2654 (O_2654,N_49768,N_49622);
nor UO_2655 (O_2655,N_49258,N_48388);
xnor UO_2656 (O_2656,N_48509,N_48460);
nand UO_2657 (O_2657,N_48257,N_49351);
xnor UO_2658 (O_2658,N_48420,N_48108);
and UO_2659 (O_2659,N_49523,N_47544);
nand UO_2660 (O_2660,N_47763,N_47698);
nand UO_2661 (O_2661,N_48553,N_48812);
and UO_2662 (O_2662,N_49687,N_48752);
or UO_2663 (O_2663,N_48388,N_49008);
or UO_2664 (O_2664,N_48062,N_48266);
nor UO_2665 (O_2665,N_48112,N_47620);
xnor UO_2666 (O_2666,N_49023,N_47879);
xor UO_2667 (O_2667,N_49629,N_48787);
or UO_2668 (O_2668,N_49578,N_49647);
nor UO_2669 (O_2669,N_49557,N_49494);
nand UO_2670 (O_2670,N_48907,N_49638);
or UO_2671 (O_2671,N_49015,N_49838);
and UO_2672 (O_2672,N_47837,N_47598);
and UO_2673 (O_2673,N_47631,N_48881);
xnor UO_2674 (O_2674,N_48192,N_49738);
nor UO_2675 (O_2675,N_47622,N_48348);
nor UO_2676 (O_2676,N_48806,N_49913);
nand UO_2677 (O_2677,N_49889,N_48233);
or UO_2678 (O_2678,N_48954,N_49989);
or UO_2679 (O_2679,N_49089,N_48985);
or UO_2680 (O_2680,N_47603,N_48853);
or UO_2681 (O_2681,N_48325,N_49624);
and UO_2682 (O_2682,N_49552,N_48510);
xnor UO_2683 (O_2683,N_49275,N_49083);
or UO_2684 (O_2684,N_47758,N_47869);
and UO_2685 (O_2685,N_47789,N_49140);
or UO_2686 (O_2686,N_49453,N_47904);
nand UO_2687 (O_2687,N_49072,N_49988);
nand UO_2688 (O_2688,N_48923,N_48483);
or UO_2689 (O_2689,N_48905,N_48136);
nand UO_2690 (O_2690,N_48553,N_48479);
xor UO_2691 (O_2691,N_47670,N_49784);
and UO_2692 (O_2692,N_47953,N_49426);
nor UO_2693 (O_2693,N_49110,N_49734);
or UO_2694 (O_2694,N_47854,N_49047);
or UO_2695 (O_2695,N_49702,N_49794);
and UO_2696 (O_2696,N_49973,N_47587);
nor UO_2697 (O_2697,N_47705,N_49714);
nor UO_2698 (O_2698,N_48550,N_49378);
or UO_2699 (O_2699,N_48685,N_48038);
xnor UO_2700 (O_2700,N_49519,N_49012);
xor UO_2701 (O_2701,N_48885,N_49404);
xnor UO_2702 (O_2702,N_48874,N_47893);
and UO_2703 (O_2703,N_48926,N_49900);
nand UO_2704 (O_2704,N_48751,N_49729);
nor UO_2705 (O_2705,N_47813,N_49875);
nand UO_2706 (O_2706,N_49727,N_47523);
xor UO_2707 (O_2707,N_47594,N_48237);
nand UO_2708 (O_2708,N_48878,N_49082);
or UO_2709 (O_2709,N_48605,N_48023);
nor UO_2710 (O_2710,N_48206,N_47517);
xnor UO_2711 (O_2711,N_47990,N_47880);
or UO_2712 (O_2712,N_48735,N_49853);
xnor UO_2713 (O_2713,N_49819,N_49376);
and UO_2714 (O_2714,N_47546,N_48393);
or UO_2715 (O_2715,N_47892,N_49893);
nor UO_2716 (O_2716,N_47591,N_48876);
and UO_2717 (O_2717,N_48574,N_49257);
xor UO_2718 (O_2718,N_49903,N_48399);
and UO_2719 (O_2719,N_49529,N_49838);
xnor UO_2720 (O_2720,N_49069,N_48537);
nor UO_2721 (O_2721,N_47649,N_47773);
or UO_2722 (O_2722,N_49096,N_48625);
and UO_2723 (O_2723,N_48133,N_47521);
or UO_2724 (O_2724,N_48627,N_48828);
or UO_2725 (O_2725,N_47836,N_49588);
or UO_2726 (O_2726,N_48507,N_49451);
nor UO_2727 (O_2727,N_49221,N_48288);
xor UO_2728 (O_2728,N_48687,N_47930);
and UO_2729 (O_2729,N_47505,N_49366);
or UO_2730 (O_2730,N_49922,N_48207);
nor UO_2731 (O_2731,N_47946,N_48943);
nand UO_2732 (O_2732,N_47563,N_49634);
xor UO_2733 (O_2733,N_49433,N_48641);
and UO_2734 (O_2734,N_48928,N_48763);
xnor UO_2735 (O_2735,N_48688,N_48940);
xnor UO_2736 (O_2736,N_48177,N_48064);
or UO_2737 (O_2737,N_48028,N_48152);
and UO_2738 (O_2738,N_47742,N_48707);
nor UO_2739 (O_2739,N_48459,N_47506);
xor UO_2740 (O_2740,N_49964,N_49989);
nand UO_2741 (O_2741,N_49306,N_49103);
or UO_2742 (O_2742,N_48386,N_49527);
xnor UO_2743 (O_2743,N_48754,N_48218);
xor UO_2744 (O_2744,N_49861,N_47887);
nand UO_2745 (O_2745,N_48172,N_47981);
nor UO_2746 (O_2746,N_48494,N_48719);
nand UO_2747 (O_2747,N_48818,N_47832);
nand UO_2748 (O_2748,N_48363,N_48714);
and UO_2749 (O_2749,N_49979,N_49246);
or UO_2750 (O_2750,N_49928,N_47521);
nand UO_2751 (O_2751,N_49106,N_48464);
xor UO_2752 (O_2752,N_47881,N_49758);
or UO_2753 (O_2753,N_49926,N_49061);
and UO_2754 (O_2754,N_49706,N_49544);
nand UO_2755 (O_2755,N_48714,N_48772);
or UO_2756 (O_2756,N_49859,N_47664);
or UO_2757 (O_2757,N_48953,N_49976);
xor UO_2758 (O_2758,N_49906,N_48684);
xor UO_2759 (O_2759,N_49885,N_48913);
or UO_2760 (O_2760,N_47677,N_47783);
nor UO_2761 (O_2761,N_47993,N_49216);
xor UO_2762 (O_2762,N_47982,N_48315);
and UO_2763 (O_2763,N_48345,N_49146);
or UO_2764 (O_2764,N_48403,N_48347);
xor UO_2765 (O_2765,N_49579,N_48472);
nor UO_2766 (O_2766,N_48232,N_49086);
nand UO_2767 (O_2767,N_48606,N_48061);
or UO_2768 (O_2768,N_48939,N_48199);
or UO_2769 (O_2769,N_49918,N_48457);
or UO_2770 (O_2770,N_47554,N_48708);
and UO_2771 (O_2771,N_48296,N_49083);
and UO_2772 (O_2772,N_48978,N_48429);
or UO_2773 (O_2773,N_49484,N_49614);
xor UO_2774 (O_2774,N_49698,N_48500);
nor UO_2775 (O_2775,N_49993,N_47532);
or UO_2776 (O_2776,N_48289,N_49870);
nand UO_2777 (O_2777,N_48994,N_48434);
and UO_2778 (O_2778,N_47814,N_47940);
or UO_2779 (O_2779,N_49172,N_47895);
or UO_2780 (O_2780,N_49057,N_48657);
nor UO_2781 (O_2781,N_48734,N_48105);
nand UO_2782 (O_2782,N_49320,N_49372);
nand UO_2783 (O_2783,N_47686,N_48991);
and UO_2784 (O_2784,N_48975,N_48195);
nor UO_2785 (O_2785,N_47768,N_49802);
or UO_2786 (O_2786,N_49411,N_49825);
nand UO_2787 (O_2787,N_47990,N_47558);
nor UO_2788 (O_2788,N_49037,N_47942);
and UO_2789 (O_2789,N_48373,N_48227);
xnor UO_2790 (O_2790,N_49923,N_49746);
nand UO_2791 (O_2791,N_48125,N_48138);
and UO_2792 (O_2792,N_49779,N_48890);
and UO_2793 (O_2793,N_48152,N_49061);
nand UO_2794 (O_2794,N_48222,N_49399);
nor UO_2795 (O_2795,N_49329,N_47637);
nor UO_2796 (O_2796,N_49411,N_49797);
or UO_2797 (O_2797,N_48154,N_48889);
nor UO_2798 (O_2798,N_48772,N_47802);
and UO_2799 (O_2799,N_49255,N_48865);
nand UO_2800 (O_2800,N_48660,N_48927);
nor UO_2801 (O_2801,N_49761,N_49391);
nor UO_2802 (O_2802,N_49121,N_48009);
and UO_2803 (O_2803,N_49707,N_47782);
xor UO_2804 (O_2804,N_49006,N_49792);
or UO_2805 (O_2805,N_48110,N_48093);
nor UO_2806 (O_2806,N_48913,N_48302);
nor UO_2807 (O_2807,N_49084,N_49577);
xnor UO_2808 (O_2808,N_48646,N_47794);
and UO_2809 (O_2809,N_47987,N_49054);
or UO_2810 (O_2810,N_48049,N_47528);
or UO_2811 (O_2811,N_49778,N_49394);
and UO_2812 (O_2812,N_49133,N_48620);
nand UO_2813 (O_2813,N_48794,N_48608);
or UO_2814 (O_2814,N_48380,N_48561);
nor UO_2815 (O_2815,N_47800,N_49327);
nand UO_2816 (O_2816,N_49158,N_49186);
or UO_2817 (O_2817,N_49426,N_49292);
and UO_2818 (O_2818,N_49494,N_48288);
or UO_2819 (O_2819,N_49452,N_49484);
and UO_2820 (O_2820,N_49342,N_47801);
xor UO_2821 (O_2821,N_48662,N_48267);
nand UO_2822 (O_2822,N_48280,N_47734);
nor UO_2823 (O_2823,N_48973,N_47825);
nor UO_2824 (O_2824,N_47894,N_49578);
or UO_2825 (O_2825,N_49220,N_49433);
and UO_2826 (O_2826,N_47603,N_48145);
and UO_2827 (O_2827,N_48062,N_48068);
nand UO_2828 (O_2828,N_48206,N_47781);
xnor UO_2829 (O_2829,N_49913,N_49699);
xnor UO_2830 (O_2830,N_49989,N_48849);
nor UO_2831 (O_2831,N_47769,N_48865);
nor UO_2832 (O_2832,N_47541,N_48505);
and UO_2833 (O_2833,N_49122,N_48153);
xnor UO_2834 (O_2834,N_48837,N_49281);
nand UO_2835 (O_2835,N_48058,N_48167);
nor UO_2836 (O_2836,N_49679,N_47746);
or UO_2837 (O_2837,N_47587,N_47528);
and UO_2838 (O_2838,N_49039,N_49698);
or UO_2839 (O_2839,N_48935,N_48549);
and UO_2840 (O_2840,N_48292,N_48944);
nand UO_2841 (O_2841,N_49879,N_49269);
and UO_2842 (O_2842,N_49072,N_47743);
nor UO_2843 (O_2843,N_48998,N_48613);
nor UO_2844 (O_2844,N_47571,N_49089);
nor UO_2845 (O_2845,N_48247,N_48422);
xor UO_2846 (O_2846,N_49614,N_49016);
and UO_2847 (O_2847,N_48772,N_49192);
nor UO_2848 (O_2848,N_47948,N_47637);
or UO_2849 (O_2849,N_47967,N_49477);
or UO_2850 (O_2850,N_48679,N_49885);
nand UO_2851 (O_2851,N_47826,N_49611);
and UO_2852 (O_2852,N_48284,N_48242);
nor UO_2853 (O_2853,N_48027,N_48080);
or UO_2854 (O_2854,N_48804,N_47932);
nand UO_2855 (O_2855,N_49292,N_48794);
or UO_2856 (O_2856,N_49397,N_48513);
nand UO_2857 (O_2857,N_47561,N_48044);
xor UO_2858 (O_2858,N_47653,N_48068);
or UO_2859 (O_2859,N_47870,N_48585);
nor UO_2860 (O_2860,N_48854,N_49391);
nand UO_2861 (O_2861,N_49799,N_47666);
nor UO_2862 (O_2862,N_49994,N_49493);
and UO_2863 (O_2863,N_48059,N_49263);
nor UO_2864 (O_2864,N_47971,N_49528);
nor UO_2865 (O_2865,N_49871,N_49481);
xor UO_2866 (O_2866,N_48680,N_49813);
and UO_2867 (O_2867,N_48846,N_48047);
nand UO_2868 (O_2868,N_49685,N_48762);
nor UO_2869 (O_2869,N_49554,N_47622);
nor UO_2870 (O_2870,N_49560,N_47664);
and UO_2871 (O_2871,N_49385,N_49009);
and UO_2872 (O_2872,N_49999,N_49606);
and UO_2873 (O_2873,N_47621,N_48902);
nand UO_2874 (O_2874,N_49618,N_48527);
or UO_2875 (O_2875,N_48207,N_49326);
or UO_2876 (O_2876,N_48299,N_47732);
or UO_2877 (O_2877,N_49474,N_47584);
nor UO_2878 (O_2878,N_48775,N_48564);
or UO_2879 (O_2879,N_48458,N_48831);
or UO_2880 (O_2880,N_48936,N_49922);
nand UO_2881 (O_2881,N_48061,N_49349);
and UO_2882 (O_2882,N_49338,N_49497);
xnor UO_2883 (O_2883,N_48605,N_48165);
xor UO_2884 (O_2884,N_47873,N_49082);
nor UO_2885 (O_2885,N_49565,N_48346);
nand UO_2886 (O_2886,N_49792,N_48800);
xnor UO_2887 (O_2887,N_49782,N_49696);
xnor UO_2888 (O_2888,N_48892,N_49765);
nand UO_2889 (O_2889,N_49003,N_47973);
xnor UO_2890 (O_2890,N_47617,N_48229);
nand UO_2891 (O_2891,N_49864,N_48883);
or UO_2892 (O_2892,N_48146,N_48037);
nand UO_2893 (O_2893,N_49564,N_49828);
nor UO_2894 (O_2894,N_48261,N_47552);
nor UO_2895 (O_2895,N_47566,N_49579);
nand UO_2896 (O_2896,N_48822,N_48093);
xor UO_2897 (O_2897,N_48830,N_49287);
and UO_2898 (O_2898,N_48526,N_49996);
xor UO_2899 (O_2899,N_48276,N_48352);
and UO_2900 (O_2900,N_48228,N_48303);
nand UO_2901 (O_2901,N_48451,N_48962);
nor UO_2902 (O_2902,N_49797,N_49976);
nand UO_2903 (O_2903,N_48582,N_48266);
and UO_2904 (O_2904,N_49120,N_47944);
and UO_2905 (O_2905,N_47749,N_49567);
nand UO_2906 (O_2906,N_47526,N_49633);
nor UO_2907 (O_2907,N_49588,N_49589);
xnor UO_2908 (O_2908,N_48317,N_49269);
xor UO_2909 (O_2909,N_49293,N_49268);
nor UO_2910 (O_2910,N_47518,N_47638);
and UO_2911 (O_2911,N_47873,N_49491);
and UO_2912 (O_2912,N_49134,N_49789);
and UO_2913 (O_2913,N_49336,N_47781);
and UO_2914 (O_2914,N_48367,N_48791);
and UO_2915 (O_2915,N_47579,N_48546);
and UO_2916 (O_2916,N_49015,N_49842);
and UO_2917 (O_2917,N_48793,N_47685);
and UO_2918 (O_2918,N_48509,N_47654);
nor UO_2919 (O_2919,N_48550,N_48932);
nor UO_2920 (O_2920,N_49820,N_49810);
nor UO_2921 (O_2921,N_49821,N_48927);
nor UO_2922 (O_2922,N_47894,N_47804);
nor UO_2923 (O_2923,N_47537,N_49662);
and UO_2924 (O_2924,N_49405,N_48610);
xor UO_2925 (O_2925,N_49286,N_49706);
or UO_2926 (O_2926,N_49977,N_49794);
or UO_2927 (O_2927,N_48948,N_48971);
and UO_2928 (O_2928,N_48880,N_47638);
nor UO_2929 (O_2929,N_49436,N_47549);
nand UO_2930 (O_2930,N_48162,N_48816);
and UO_2931 (O_2931,N_48586,N_48484);
and UO_2932 (O_2932,N_47603,N_49193);
nand UO_2933 (O_2933,N_47805,N_47971);
nor UO_2934 (O_2934,N_47902,N_49670);
or UO_2935 (O_2935,N_48297,N_49767);
or UO_2936 (O_2936,N_48562,N_47533);
and UO_2937 (O_2937,N_49480,N_48196);
nand UO_2938 (O_2938,N_48079,N_49543);
nor UO_2939 (O_2939,N_48039,N_48817);
and UO_2940 (O_2940,N_49822,N_49797);
nor UO_2941 (O_2941,N_47745,N_47957);
xor UO_2942 (O_2942,N_49442,N_48534);
and UO_2943 (O_2943,N_48283,N_49056);
xor UO_2944 (O_2944,N_48849,N_49875);
and UO_2945 (O_2945,N_49142,N_47686);
nand UO_2946 (O_2946,N_48095,N_48323);
nor UO_2947 (O_2947,N_49962,N_49276);
xor UO_2948 (O_2948,N_49499,N_49109);
nand UO_2949 (O_2949,N_48955,N_49194);
xnor UO_2950 (O_2950,N_48563,N_48447);
nor UO_2951 (O_2951,N_49253,N_49936);
and UO_2952 (O_2952,N_48329,N_47820);
nor UO_2953 (O_2953,N_47760,N_49130);
nand UO_2954 (O_2954,N_49124,N_48457);
nor UO_2955 (O_2955,N_48056,N_49493);
xor UO_2956 (O_2956,N_47830,N_48733);
or UO_2957 (O_2957,N_47789,N_47565);
xnor UO_2958 (O_2958,N_49551,N_48815);
or UO_2959 (O_2959,N_48647,N_49366);
and UO_2960 (O_2960,N_47708,N_49151);
or UO_2961 (O_2961,N_47914,N_47509);
nand UO_2962 (O_2962,N_47755,N_49189);
xnor UO_2963 (O_2963,N_48381,N_48027);
and UO_2964 (O_2964,N_49434,N_47835);
or UO_2965 (O_2965,N_49080,N_48210);
nor UO_2966 (O_2966,N_48976,N_48314);
or UO_2967 (O_2967,N_49752,N_48628);
and UO_2968 (O_2968,N_49165,N_49365);
and UO_2969 (O_2969,N_49289,N_47654);
xnor UO_2970 (O_2970,N_49782,N_49302);
xor UO_2971 (O_2971,N_48535,N_49228);
nand UO_2972 (O_2972,N_49399,N_48456);
nand UO_2973 (O_2973,N_49177,N_49391);
or UO_2974 (O_2974,N_49426,N_49558);
and UO_2975 (O_2975,N_48093,N_48756);
nor UO_2976 (O_2976,N_49693,N_48937);
nand UO_2977 (O_2977,N_48507,N_48032);
or UO_2978 (O_2978,N_49340,N_48667);
and UO_2979 (O_2979,N_48628,N_48558);
or UO_2980 (O_2980,N_48429,N_49366);
nand UO_2981 (O_2981,N_49999,N_48932);
and UO_2982 (O_2982,N_49647,N_47850);
xnor UO_2983 (O_2983,N_49988,N_49506);
or UO_2984 (O_2984,N_48294,N_49806);
or UO_2985 (O_2985,N_49278,N_49917);
nand UO_2986 (O_2986,N_47566,N_49551);
nor UO_2987 (O_2987,N_48116,N_49582);
xor UO_2988 (O_2988,N_49447,N_48270);
and UO_2989 (O_2989,N_49691,N_47890);
or UO_2990 (O_2990,N_49689,N_49251);
and UO_2991 (O_2991,N_48887,N_48613);
nor UO_2992 (O_2992,N_49370,N_48659);
nand UO_2993 (O_2993,N_47976,N_47814);
or UO_2994 (O_2994,N_48745,N_48119);
xnor UO_2995 (O_2995,N_48771,N_47593);
xnor UO_2996 (O_2996,N_48495,N_48982);
and UO_2997 (O_2997,N_49953,N_49976);
or UO_2998 (O_2998,N_47879,N_48095);
nand UO_2999 (O_2999,N_49975,N_49321);
xnor UO_3000 (O_3000,N_47642,N_48540);
xor UO_3001 (O_3001,N_49935,N_49122);
or UO_3002 (O_3002,N_48717,N_47957);
and UO_3003 (O_3003,N_47678,N_49812);
or UO_3004 (O_3004,N_48159,N_48163);
xor UO_3005 (O_3005,N_48351,N_49444);
nor UO_3006 (O_3006,N_49128,N_47872);
nor UO_3007 (O_3007,N_49365,N_49037);
or UO_3008 (O_3008,N_47785,N_47503);
or UO_3009 (O_3009,N_49729,N_49395);
nand UO_3010 (O_3010,N_49388,N_48783);
nor UO_3011 (O_3011,N_48933,N_49421);
or UO_3012 (O_3012,N_47854,N_49466);
nor UO_3013 (O_3013,N_49865,N_48419);
xor UO_3014 (O_3014,N_48522,N_48596);
xnor UO_3015 (O_3015,N_49731,N_47689);
or UO_3016 (O_3016,N_47562,N_48574);
nor UO_3017 (O_3017,N_49874,N_48072);
or UO_3018 (O_3018,N_49064,N_48452);
or UO_3019 (O_3019,N_49974,N_47889);
nor UO_3020 (O_3020,N_49557,N_47837);
or UO_3021 (O_3021,N_47651,N_49404);
nor UO_3022 (O_3022,N_48105,N_47500);
and UO_3023 (O_3023,N_47561,N_49358);
or UO_3024 (O_3024,N_48168,N_49239);
xor UO_3025 (O_3025,N_49820,N_48632);
nor UO_3026 (O_3026,N_49969,N_49292);
nor UO_3027 (O_3027,N_48732,N_48016);
nand UO_3028 (O_3028,N_49738,N_47938);
and UO_3029 (O_3029,N_49368,N_49437);
nor UO_3030 (O_3030,N_48523,N_48489);
nor UO_3031 (O_3031,N_49547,N_48554);
and UO_3032 (O_3032,N_47517,N_48571);
and UO_3033 (O_3033,N_48895,N_49224);
nor UO_3034 (O_3034,N_48396,N_49392);
and UO_3035 (O_3035,N_49358,N_48127);
or UO_3036 (O_3036,N_49353,N_48277);
xor UO_3037 (O_3037,N_47805,N_48308);
nand UO_3038 (O_3038,N_48446,N_48582);
or UO_3039 (O_3039,N_47911,N_49395);
and UO_3040 (O_3040,N_48357,N_47935);
nor UO_3041 (O_3041,N_48642,N_48278);
or UO_3042 (O_3042,N_48156,N_47896);
nor UO_3043 (O_3043,N_48791,N_49899);
xnor UO_3044 (O_3044,N_48985,N_49950);
nor UO_3045 (O_3045,N_49911,N_49368);
nor UO_3046 (O_3046,N_48373,N_48438);
or UO_3047 (O_3047,N_49298,N_49443);
and UO_3048 (O_3048,N_49812,N_48901);
or UO_3049 (O_3049,N_49081,N_48988);
and UO_3050 (O_3050,N_47609,N_48906);
xor UO_3051 (O_3051,N_49559,N_48571);
nand UO_3052 (O_3052,N_49914,N_49540);
nor UO_3053 (O_3053,N_49182,N_48210);
and UO_3054 (O_3054,N_49851,N_47589);
nor UO_3055 (O_3055,N_48703,N_47541);
nand UO_3056 (O_3056,N_48356,N_49092);
or UO_3057 (O_3057,N_49970,N_48571);
xor UO_3058 (O_3058,N_49411,N_49767);
or UO_3059 (O_3059,N_49857,N_49861);
nand UO_3060 (O_3060,N_49045,N_48987);
or UO_3061 (O_3061,N_48084,N_48595);
xor UO_3062 (O_3062,N_49143,N_49575);
nor UO_3063 (O_3063,N_49537,N_47681);
nand UO_3064 (O_3064,N_49399,N_47556);
nand UO_3065 (O_3065,N_47974,N_48564);
xnor UO_3066 (O_3066,N_49426,N_48097);
or UO_3067 (O_3067,N_49664,N_47581);
or UO_3068 (O_3068,N_49312,N_49397);
nand UO_3069 (O_3069,N_49267,N_49295);
or UO_3070 (O_3070,N_49235,N_49858);
and UO_3071 (O_3071,N_48186,N_47890);
nand UO_3072 (O_3072,N_49253,N_49701);
nor UO_3073 (O_3073,N_49335,N_48651);
nand UO_3074 (O_3074,N_48539,N_49095);
and UO_3075 (O_3075,N_49075,N_48197);
nor UO_3076 (O_3076,N_48049,N_48354);
or UO_3077 (O_3077,N_48285,N_49945);
or UO_3078 (O_3078,N_48367,N_49960);
or UO_3079 (O_3079,N_48711,N_49923);
nand UO_3080 (O_3080,N_48252,N_49906);
nand UO_3081 (O_3081,N_49052,N_48735);
or UO_3082 (O_3082,N_49239,N_48067);
nand UO_3083 (O_3083,N_49255,N_48094);
xnor UO_3084 (O_3084,N_49862,N_48940);
and UO_3085 (O_3085,N_49346,N_47592);
xor UO_3086 (O_3086,N_48898,N_47668);
or UO_3087 (O_3087,N_48142,N_48374);
nor UO_3088 (O_3088,N_48375,N_48519);
nand UO_3089 (O_3089,N_47924,N_47673);
or UO_3090 (O_3090,N_47732,N_49034);
nor UO_3091 (O_3091,N_48580,N_47670);
nand UO_3092 (O_3092,N_49912,N_48069);
and UO_3093 (O_3093,N_48721,N_48578);
nand UO_3094 (O_3094,N_49035,N_49001);
nand UO_3095 (O_3095,N_49350,N_47606);
nor UO_3096 (O_3096,N_48783,N_48414);
and UO_3097 (O_3097,N_49933,N_49514);
nor UO_3098 (O_3098,N_49355,N_49751);
nor UO_3099 (O_3099,N_48333,N_48051);
xnor UO_3100 (O_3100,N_49858,N_48624);
and UO_3101 (O_3101,N_47891,N_48340);
and UO_3102 (O_3102,N_48361,N_48145);
nand UO_3103 (O_3103,N_47788,N_48503);
and UO_3104 (O_3104,N_48533,N_49630);
nor UO_3105 (O_3105,N_49573,N_48642);
xor UO_3106 (O_3106,N_49636,N_49274);
nor UO_3107 (O_3107,N_47827,N_49613);
xnor UO_3108 (O_3108,N_47978,N_49362);
nand UO_3109 (O_3109,N_48934,N_49052);
or UO_3110 (O_3110,N_48391,N_49057);
nand UO_3111 (O_3111,N_49682,N_49789);
and UO_3112 (O_3112,N_48543,N_47623);
or UO_3113 (O_3113,N_49780,N_49706);
or UO_3114 (O_3114,N_48961,N_49571);
xnor UO_3115 (O_3115,N_48074,N_49384);
and UO_3116 (O_3116,N_47508,N_49635);
xor UO_3117 (O_3117,N_49807,N_48857);
and UO_3118 (O_3118,N_49606,N_49808);
nand UO_3119 (O_3119,N_48031,N_49715);
xor UO_3120 (O_3120,N_48161,N_47678);
nand UO_3121 (O_3121,N_47564,N_48140);
nand UO_3122 (O_3122,N_49877,N_47579);
nand UO_3123 (O_3123,N_48501,N_47753);
nand UO_3124 (O_3124,N_49078,N_49255);
nor UO_3125 (O_3125,N_48265,N_48066);
xor UO_3126 (O_3126,N_47569,N_48844);
nor UO_3127 (O_3127,N_48519,N_49353);
or UO_3128 (O_3128,N_48313,N_49576);
nand UO_3129 (O_3129,N_48154,N_48056);
and UO_3130 (O_3130,N_48044,N_48946);
and UO_3131 (O_3131,N_49625,N_47780);
nand UO_3132 (O_3132,N_49826,N_48323);
and UO_3133 (O_3133,N_49222,N_48222);
nand UO_3134 (O_3134,N_48611,N_47734);
xor UO_3135 (O_3135,N_49298,N_47974);
and UO_3136 (O_3136,N_47808,N_47809);
or UO_3137 (O_3137,N_49856,N_48010);
nand UO_3138 (O_3138,N_47736,N_47884);
or UO_3139 (O_3139,N_49984,N_49705);
xnor UO_3140 (O_3140,N_49064,N_47812);
xor UO_3141 (O_3141,N_49506,N_47563);
nand UO_3142 (O_3142,N_49974,N_48378);
xor UO_3143 (O_3143,N_48627,N_48044);
nand UO_3144 (O_3144,N_47838,N_48948);
nor UO_3145 (O_3145,N_48490,N_48219);
or UO_3146 (O_3146,N_48123,N_48946);
nand UO_3147 (O_3147,N_47753,N_48674);
and UO_3148 (O_3148,N_48791,N_49600);
or UO_3149 (O_3149,N_47523,N_48655);
nand UO_3150 (O_3150,N_49553,N_48743);
or UO_3151 (O_3151,N_49040,N_48660);
and UO_3152 (O_3152,N_47505,N_47896);
and UO_3153 (O_3153,N_49994,N_49977);
nor UO_3154 (O_3154,N_48635,N_47696);
or UO_3155 (O_3155,N_49386,N_49469);
nor UO_3156 (O_3156,N_48665,N_49522);
nand UO_3157 (O_3157,N_48633,N_48658);
xor UO_3158 (O_3158,N_47634,N_49666);
nor UO_3159 (O_3159,N_49717,N_49419);
nand UO_3160 (O_3160,N_49881,N_47612);
nand UO_3161 (O_3161,N_47688,N_48589);
nand UO_3162 (O_3162,N_48913,N_48945);
and UO_3163 (O_3163,N_47555,N_48063);
nor UO_3164 (O_3164,N_49457,N_48863);
nor UO_3165 (O_3165,N_48496,N_49351);
nor UO_3166 (O_3166,N_47914,N_49150);
xnor UO_3167 (O_3167,N_49583,N_49132);
and UO_3168 (O_3168,N_49542,N_47531);
or UO_3169 (O_3169,N_48708,N_49385);
and UO_3170 (O_3170,N_48149,N_49191);
nand UO_3171 (O_3171,N_48358,N_49857);
nand UO_3172 (O_3172,N_48239,N_48873);
xor UO_3173 (O_3173,N_47912,N_49421);
nor UO_3174 (O_3174,N_49257,N_47841);
and UO_3175 (O_3175,N_49355,N_48217);
and UO_3176 (O_3176,N_49444,N_48635);
xnor UO_3177 (O_3177,N_47545,N_47542);
and UO_3178 (O_3178,N_47903,N_48120);
or UO_3179 (O_3179,N_49897,N_49641);
nor UO_3180 (O_3180,N_47976,N_48969);
or UO_3181 (O_3181,N_47750,N_49266);
and UO_3182 (O_3182,N_47927,N_48828);
nand UO_3183 (O_3183,N_49157,N_47950);
or UO_3184 (O_3184,N_47690,N_49739);
or UO_3185 (O_3185,N_48339,N_47507);
nor UO_3186 (O_3186,N_49104,N_49912);
nor UO_3187 (O_3187,N_49187,N_48917);
and UO_3188 (O_3188,N_48761,N_49515);
and UO_3189 (O_3189,N_48218,N_49864);
or UO_3190 (O_3190,N_48773,N_49473);
or UO_3191 (O_3191,N_48518,N_47805);
and UO_3192 (O_3192,N_49149,N_47632);
and UO_3193 (O_3193,N_47980,N_49935);
or UO_3194 (O_3194,N_47561,N_49306);
and UO_3195 (O_3195,N_49458,N_49560);
or UO_3196 (O_3196,N_48352,N_49289);
nand UO_3197 (O_3197,N_49696,N_49353);
nor UO_3198 (O_3198,N_49648,N_48653);
nand UO_3199 (O_3199,N_49222,N_48161);
and UO_3200 (O_3200,N_49200,N_49935);
xnor UO_3201 (O_3201,N_48574,N_49526);
or UO_3202 (O_3202,N_49851,N_48576);
nor UO_3203 (O_3203,N_48714,N_49651);
and UO_3204 (O_3204,N_47623,N_47592);
xor UO_3205 (O_3205,N_49827,N_48092);
nor UO_3206 (O_3206,N_49903,N_48057);
xor UO_3207 (O_3207,N_49772,N_49316);
or UO_3208 (O_3208,N_49034,N_49468);
nand UO_3209 (O_3209,N_48091,N_49332);
or UO_3210 (O_3210,N_47510,N_48942);
nor UO_3211 (O_3211,N_48876,N_47848);
xor UO_3212 (O_3212,N_48514,N_48104);
and UO_3213 (O_3213,N_48954,N_48682);
xnor UO_3214 (O_3214,N_49157,N_48051);
and UO_3215 (O_3215,N_48028,N_47783);
nand UO_3216 (O_3216,N_49330,N_49517);
xnor UO_3217 (O_3217,N_48853,N_47806);
nor UO_3218 (O_3218,N_47782,N_47780);
nor UO_3219 (O_3219,N_47811,N_48213);
nand UO_3220 (O_3220,N_48170,N_48592);
xnor UO_3221 (O_3221,N_49024,N_48985);
nand UO_3222 (O_3222,N_47805,N_48387);
or UO_3223 (O_3223,N_48923,N_47664);
nand UO_3224 (O_3224,N_47853,N_48617);
nor UO_3225 (O_3225,N_47613,N_47797);
nand UO_3226 (O_3226,N_49690,N_49529);
nor UO_3227 (O_3227,N_47656,N_47553);
nor UO_3228 (O_3228,N_48916,N_48353);
or UO_3229 (O_3229,N_48004,N_48287);
nor UO_3230 (O_3230,N_49115,N_49616);
nor UO_3231 (O_3231,N_48803,N_49525);
or UO_3232 (O_3232,N_48301,N_48592);
or UO_3233 (O_3233,N_48273,N_48942);
or UO_3234 (O_3234,N_48144,N_48103);
nor UO_3235 (O_3235,N_48076,N_48219);
nand UO_3236 (O_3236,N_48718,N_48366);
xnor UO_3237 (O_3237,N_47856,N_49315);
nor UO_3238 (O_3238,N_47577,N_47784);
xor UO_3239 (O_3239,N_49059,N_48038);
nor UO_3240 (O_3240,N_49017,N_47557);
nand UO_3241 (O_3241,N_47597,N_49479);
or UO_3242 (O_3242,N_48407,N_48050);
or UO_3243 (O_3243,N_49626,N_48951);
xor UO_3244 (O_3244,N_48948,N_47641);
and UO_3245 (O_3245,N_49543,N_48566);
xnor UO_3246 (O_3246,N_49481,N_48954);
and UO_3247 (O_3247,N_48670,N_49244);
nand UO_3248 (O_3248,N_48982,N_49884);
nand UO_3249 (O_3249,N_48232,N_49090);
nor UO_3250 (O_3250,N_48311,N_47806);
and UO_3251 (O_3251,N_48976,N_48819);
and UO_3252 (O_3252,N_49921,N_49347);
nor UO_3253 (O_3253,N_49967,N_49729);
nand UO_3254 (O_3254,N_49347,N_47735);
xnor UO_3255 (O_3255,N_48985,N_48227);
nor UO_3256 (O_3256,N_49637,N_47788);
nand UO_3257 (O_3257,N_49760,N_47830);
xnor UO_3258 (O_3258,N_49748,N_48794);
xor UO_3259 (O_3259,N_49310,N_47529);
nand UO_3260 (O_3260,N_48801,N_48891);
nand UO_3261 (O_3261,N_48274,N_47852);
nand UO_3262 (O_3262,N_49564,N_47578);
or UO_3263 (O_3263,N_48413,N_49453);
and UO_3264 (O_3264,N_47795,N_49907);
nand UO_3265 (O_3265,N_47563,N_48855);
or UO_3266 (O_3266,N_49896,N_49445);
or UO_3267 (O_3267,N_48821,N_47831);
xor UO_3268 (O_3268,N_49124,N_47530);
or UO_3269 (O_3269,N_48355,N_49111);
xor UO_3270 (O_3270,N_49573,N_49403);
nand UO_3271 (O_3271,N_48413,N_49857);
nand UO_3272 (O_3272,N_48434,N_49477);
xor UO_3273 (O_3273,N_48997,N_49335);
or UO_3274 (O_3274,N_47534,N_49203);
nand UO_3275 (O_3275,N_47609,N_48001);
xor UO_3276 (O_3276,N_49420,N_49494);
nor UO_3277 (O_3277,N_47795,N_49275);
and UO_3278 (O_3278,N_48618,N_48627);
nor UO_3279 (O_3279,N_48745,N_48774);
nand UO_3280 (O_3280,N_47929,N_48264);
nor UO_3281 (O_3281,N_48463,N_48719);
nor UO_3282 (O_3282,N_49745,N_48193);
and UO_3283 (O_3283,N_49375,N_49100);
xnor UO_3284 (O_3284,N_48254,N_49904);
xor UO_3285 (O_3285,N_48791,N_49118);
nand UO_3286 (O_3286,N_49926,N_48564);
or UO_3287 (O_3287,N_48777,N_49303);
nor UO_3288 (O_3288,N_48114,N_49834);
nor UO_3289 (O_3289,N_49199,N_47913);
xnor UO_3290 (O_3290,N_48724,N_49993);
or UO_3291 (O_3291,N_49586,N_49145);
or UO_3292 (O_3292,N_48985,N_47815);
and UO_3293 (O_3293,N_49835,N_47711);
and UO_3294 (O_3294,N_47647,N_48760);
xnor UO_3295 (O_3295,N_48711,N_47729);
nand UO_3296 (O_3296,N_49449,N_48010);
and UO_3297 (O_3297,N_48608,N_47684);
nor UO_3298 (O_3298,N_49857,N_48692);
nor UO_3299 (O_3299,N_47531,N_49129);
xnor UO_3300 (O_3300,N_49581,N_49711);
xor UO_3301 (O_3301,N_48291,N_47551);
xor UO_3302 (O_3302,N_49204,N_48662);
nor UO_3303 (O_3303,N_49567,N_48686);
nand UO_3304 (O_3304,N_48416,N_47506);
xnor UO_3305 (O_3305,N_48435,N_49713);
nor UO_3306 (O_3306,N_49280,N_48067);
nor UO_3307 (O_3307,N_49000,N_49417);
nand UO_3308 (O_3308,N_47565,N_49345);
or UO_3309 (O_3309,N_47780,N_48797);
or UO_3310 (O_3310,N_49340,N_48624);
nand UO_3311 (O_3311,N_48180,N_49929);
xnor UO_3312 (O_3312,N_49251,N_49330);
nand UO_3313 (O_3313,N_48796,N_47617);
nand UO_3314 (O_3314,N_48897,N_49330);
or UO_3315 (O_3315,N_49112,N_49020);
nor UO_3316 (O_3316,N_47724,N_48231);
nand UO_3317 (O_3317,N_48891,N_49888);
nand UO_3318 (O_3318,N_48928,N_49575);
or UO_3319 (O_3319,N_49126,N_49142);
or UO_3320 (O_3320,N_48982,N_49424);
nand UO_3321 (O_3321,N_48808,N_47831);
xnor UO_3322 (O_3322,N_47982,N_49208);
xor UO_3323 (O_3323,N_47903,N_47697);
nand UO_3324 (O_3324,N_48984,N_49203);
and UO_3325 (O_3325,N_48450,N_48172);
nand UO_3326 (O_3326,N_49642,N_47586);
or UO_3327 (O_3327,N_47590,N_47575);
nand UO_3328 (O_3328,N_48985,N_48865);
and UO_3329 (O_3329,N_48611,N_49826);
xor UO_3330 (O_3330,N_47883,N_49547);
nand UO_3331 (O_3331,N_48399,N_49136);
nand UO_3332 (O_3332,N_49944,N_49434);
and UO_3333 (O_3333,N_49526,N_49653);
nor UO_3334 (O_3334,N_48915,N_49913);
nor UO_3335 (O_3335,N_49917,N_48540);
nand UO_3336 (O_3336,N_49668,N_47776);
and UO_3337 (O_3337,N_47534,N_49954);
or UO_3338 (O_3338,N_48206,N_48350);
nand UO_3339 (O_3339,N_49313,N_48119);
and UO_3340 (O_3340,N_49737,N_48323);
nand UO_3341 (O_3341,N_49023,N_49485);
and UO_3342 (O_3342,N_48556,N_49186);
and UO_3343 (O_3343,N_47865,N_49034);
or UO_3344 (O_3344,N_49930,N_48840);
nor UO_3345 (O_3345,N_49586,N_48542);
nand UO_3346 (O_3346,N_48758,N_48459);
nand UO_3347 (O_3347,N_49772,N_47683);
and UO_3348 (O_3348,N_48360,N_48325);
and UO_3349 (O_3349,N_48127,N_48849);
or UO_3350 (O_3350,N_49198,N_49478);
and UO_3351 (O_3351,N_48710,N_49092);
nor UO_3352 (O_3352,N_49665,N_47906);
and UO_3353 (O_3353,N_48020,N_47897);
xor UO_3354 (O_3354,N_49821,N_47625);
or UO_3355 (O_3355,N_48873,N_48088);
nor UO_3356 (O_3356,N_49918,N_49365);
nand UO_3357 (O_3357,N_48104,N_49765);
nor UO_3358 (O_3358,N_49120,N_48283);
xnor UO_3359 (O_3359,N_49835,N_47529);
and UO_3360 (O_3360,N_49800,N_47587);
nor UO_3361 (O_3361,N_49666,N_47999);
nor UO_3362 (O_3362,N_48581,N_48983);
nor UO_3363 (O_3363,N_49530,N_48072);
nor UO_3364 (O_3364,N_48975,N_48405);
or UO_3365 (O_3365,N_48450,N_48519);
nand UO_3366 (O_3366,N_49718,N_49795);
nor UO_3367 (O_3367,N_49500,N_48984);
or UO_3368 (O_3368,N_48211,N_48568);
nand UO_3369 (O_3369,N_48592,N_48337);
xnor UO_3370 (O_3370,N_48204,N_49178);
nor UO_3371 (O_3371,N_49051,N_49994);
nand UO_3372 (O_3372,N_49498,N_47558);
nand UO_3373 (O_3373,N_48857,N_47871);
xor UO_3374 (O_3374,N_49425,N_49697);
and UO_3375 (O_3375,N_48661,N_49676);
nand UO_3376 (O_3376,N_49314,N_48794);
xnor UO_3377 (O_3377,N_49878,N_48445);
nand UO_3378 (O_3378,N_47933,N_49831);
or UO_3379 (O_3379,N_49654,N_47513);
nor UO_3380 (O_3380,N_48606,N_48641);
nor UO_3381 (O_3381,N_49461,N_48886);
or UO_3382 (O_3382,N_47928,N_48227);
nor UO_3383 (O_3383,N_49804,N_48278);
and UO_3384 (O_3384,N_49490,N_48755);
or UO_3385 (O_3385,N_49838,N_47699);
nor UO_3386 (O_3386,N_47557,N_49504);
nand UO_3387 (O_3387,N_49263,N_49017);
or UO_3388 (O_3388,N_48814,N_48139);
and UO_3389 (O_3389,N_49429,N_49319);
nand UO_3390 (O_3390,N_48301,N_48495);
or UO_3391 (O_3391,N_47697,N_48281);
or UO_3392 (O_3392,N_48754,N_49832);
and UO_3393 (O_3393,N_49049,N_49564);
xnor UO_3394 (O_3394,N_49236,N_47586);
or UO_3395 (O_3395,N_48838,N_48974);
nor UO_3396 (O_3396,N_49916,N_49781);
nor UO_3397 (O_3397,N_47983,N_49465);
or UO_3398 (O_3398,N_49894,N_48917);
or UO_3399 (O_3399,N_48521,N_48215);
nor UO_3400 (O_3400,N_48387,N_48500);
xnor UO_3401 (O_3401,N_49522,N_49963);
xnor UO_3402 (O_3402,N_48498,N_48090);
nand UO_3403 (O_3403,N_48017,N_48130);
xor UO_3404 (O_3404,N_49853,N_49165);
nand UO_3405 (O_3405,N_48937,N_49924);
nor UO_3406 (O_3406,N_49909,N_49115);
nor UO_3407 (O_3407,N_47845,N_49666);
nand UO_3408 (O_3408,N_49983,N_47946);
or UO_3409 (O_3409,N_47834,N_48415);
and UO_3410 (O_3410,N_49179,N_48649);
or UO_3411 (O_3411,N_47810,N_49088);
xnor UO_3412 (O_3412,N_49910,N_47689);
nand UO_3413 (O_3413,N_48943,N_49325);
and UO_3414 (O_3414,N_49120,N_49501);
xor UO_3415 (O_3415,N_49581,N_48252);
nand UO_3416 (O_3416,N_49328,N_48611);
and UO_3417 (O_3417,N_49910,N_49446);
or UO_3418 (O_3418,N_48958,N_47703);
xor UO_3419 (O_3419,N_47537,N_49420);
nand UO_3420 (O_3420,N_49788,N_48242);
xnor UO_3421 (O_3421,N_49235,N_49559);
xnor UO_3422 (O_3422,N_47785,N_48644);
or UO_3423 (O_3423,N_49877,N_48931);
nand UO_3424 (O_3424,N_49755,N_48333);
nor UO_3425 (O_3425,N_49650,N_48752);
and UO_3426 (O_3426,N_49474,N_49267);
nor UO_3427 (O_3427,N_49500,N_49099);
xnor UO_3428 (O_3428,N_48951,N_48436);
nand UO_3429 (O_3429,N_48288,N_49145);
xor UO_3430 (O_3430,N_49419,N_49114);
nor UO_3431 (O_3431,N_47880,N_49849);
nor UO_3432 (O_3432,N_49741,N_48059);
xnor UO_3433 (O_3433,N_49700,N_47519);
xor UO_3434 (O_3434,N_48615,N_47665);
nor UO_3435 (O_3435,N_48316,N_48025);
nand UO_3436 (O_3436,N_47879,N_48577);
and UO_3437 (O_3437,N_48111,N_49966);
or UO_3438 (O_3438,N_49733,N_49213);
and UO_3439 (O_3439,N_49845,N_47938);
nand UO_3440 (O_3440,N_47651,N_48604);
nor UO_3441 (O_3441,N_48125,N_49652);
and UO_3442 (O_3442,N_47740,N_49639);
xor UO_3443 (O_3443,N_47523,N_49451);
and UO_3444 (O_3444,N_48364,N_49088);
nor UO_3445 (O_3445,N_47735,N_49743);
xnor UO_3446 (O_3446,N_49487,N_49255);
xor UO_3447 (O_3447,N_49281,N_48202);
or UO_3448 (O_3448,N_49008,N_49408);
nor UO_3449 (O_3449,N_47842,N_49328);
and UO_3450 (O_3450,N_48171,N_48493);
xor UO_3451 (O_3451,N_48130,N_48075);
xor UO_3452 (O_3452,N_48879,N_48234);
nor UO_3453 (O_3453,N_49894,N_48829);
nor UO_3454 (O_3454,N_47772,N_47983);
nor UO_3455 (O_3455,N_48729,N_47915);
nor UO_3456 (O_3456,N_49694,N_48726);
or UO_3457 (O_3457,N_47973,N_49209);
xnor UO_3458 (O_3458,N_47631,N_49822);
xnor UO_3459 (O_3459,N_48634,N_47834);
nand UO_3460 (O_3460,N_49389,N_48552);
nand UO_3461 (O_3461,N_49342,N_48028);
xor UO_3462 (O_3462,N_49910,N_48554);
or UO_3463 (O_3463,N_49927,N_48593);
or UO_3464 (O_3464,N_47541,N_47893);
or UO_3465 (O_3465,N_48251,N_48208);
nand UO_3466 (O_3466,N_49345,N_48711);
or UO_3467 (O_3467,N_48968,N_47643);
and UO_3468 (O_3468,N_49365,N_48970);
or UO_3469 (O_3469,N_48534,N_48952);
nor UO_3470 (O_3470,N_48037,N_48048);
nand UO_3471 (O_3471,N_48728,N_48789);
nor UO_3472 (O_3472,N_48696,N_47720);
nand UO_3473 (O_3473,N_49957,N_48520);
xor UO_3474 (O_3474,N_49161,N_48352);
nor UO_3475 (O_3475,N_48089,N_48410);
nor UO_3476 (O_3476,N_49617,N_49053);
nand UO_3477 (O_3477,N_47903,N_48501);
nor UO_3478 (O_3478,N_48618,N_48012);
nand UO_3479 (O_3479,N_48513,N_47884);
xor UO_3480 (O_3480,N_47796,N_48020);
and UO_3481 (O_3481,N_48746,N_48644);
nor UO_3482 (O_3482,N_49757,N_49515);
nand UO_3483 (O_3483,N_48229,N_49337);
nand UO_3484 (O_3484,N_48546,N_48269);
and UO_3485 (O_3485,N_48164,N_49650);
and UO_3486 (O_3486,N_48313,N_49908);
and UO_3487 (O_3487,N_48482,N_48664);
xnor UO_3488 (O_3488,N_49890,N_47846);
or UO_3489 (O_3489,N_48129,N_49177);
or UO_3490 (O_3490,N_48865,N_48477);
or UO_3491 (O_3491,N_49201,N_49074);
nor UO_3492 (O_3492,N_47790,N_48944);
xnor UO_3493 (O_3493,N_48166,N_49620);
nor UO_3494 (O_3494,N_49900,N_48972);
nor UO_3495 (O_3495,N_48802,N_49973);
and UO_3496 (O_3496,N_47777,N_48343);
nor UO_3497 (O_3497,N_49171,N_48459);
xor UO_3498 (O_3498,N_49761,N_47617);
nor UO_3499 (O_3499,N_48857,N_49026);
xnor UO_3500 (O_3500,N_47571,N_48967);
or UO_3501 (O_3501,N_48233,N_47932);
and UO_3502 (O_3502,N_49765,N_49514);
nand UO_3503 (O_3503,N_48448,N_48919);
or UO_3504 (O_3504,N_48729,N_49447);
nor UO_3505 (O_3505,N_48369,N_48956);
or UO_3506 (O_3506,N_47685,N_48027);
nor UO_3507 (O_3507,N_48969,N_47548);
or UO_3508 (O_3508,N_49712,N_49841);
nor UO_3509 (O_3509,N_49581,N_48959);
nor UO_3510 (O_3510,N_47792,N_47640);
nor UO_3511 (O_3511,N_49075,N_48618);
and UO_3512 (O_3512,N_49319,N_48235);
xnor UO_3513 (O_3513,N_48103,N_48222);
nor UO_3514 (O_3514,N_49598,N_47825);
and UO_3515 (O_3515,N_47858,N_48176);
nand UO_3516 (O_3516,N_48394,N_49343);
nor UO_3517 (O_3517,N_47948,N_48937);
and UO_3518 (O_3518,N_49131,N_49188);
nand UO_3519 (O_3519,N_47503,N_49615);
xor UO_3520 (O_3520,N_48157,N_49671);
and UO_3521 (O_3521,N_48548,N_47756);
and UO_3522 (O_3522,N_47787,N_48149);
or UO_3523 (O_3523,N_49351,N_49483);
nand UO_3524 (O_3524,N_48052,N_49525);
or UO_3525 (O_3525,N_49751,N_48086);
nand UO_3526 (O_3526,N_49475,N_47733);
xor UO_3527 (O_3527,N_48741,N_47623);
xor UO_3528 (O_3528,N_48276,N_48687);
nand UO_3529 (O_3529,N_47568,N_48216);
nor UO_3530 (O_3530,N_48978,N_49567);
nor UO_3531 (O_3531,N_49732,N_48361);
nor UO_3532 (O_3532,N_47508,N_47592);
nand UO_3533 (O_3533,N_48059,N_49364);
or UO_3534 (O_3534,N_48391,N_47930);
and UO_3535 (O_3535,N_49121,N_49583);
and UO_3536 (O_3536,N_47553,N_48995);
nor UO_3537 (O_3537,N_49671,N_48608);
and UO_3538 (O_3538,N_48984,N_48491);
nand UO_3539 (O_3539,N_49143,N_49191);
or UO_3540 (O_3540,N_49703,N_48351);
and UO_3541 (O_3541,N_49472,N_47540);
xor UO_3542 (O_3542,N_48518,N_49385);
and UO_3543 (O_3543,N_48721,N_48060);
nand UO_3544 (O_3544,N_49417,N_47873);
and UO_3545 (O_3545,N_49255,N_49281);
or UO_3546 (O_3546,N_48272,N_49959);
xor UO_3547 (O_3547,N_49596,N_48726);
or UO_3548 (O_3548,N_48860,N_48042);
and UO_3549 (O_3549,N_47825,N_47696);
and UO_3550 (O_3550,N_47921,N_47575);
or UO_3551 (O_3551,N_48625,N_49327);
or UO_3552 (O_3552,N_48086,N_47888);
nand UO_3553 (O_3553,N_49870,N_48026);
nor UO_3554 (O_3554,N_48480,N_48401);
and UO_3555 (O_3555,N_47925,N_49127);
xnor UO_3556 (O_3556,N_49543,N_48603);
nand UO_3557 (O_3557,N_49062,N_47871);
nand UO_3558 (O_3558,N_47587,N_48426);
or UO_3559 (O_3559,N_47999,N_48962);
and UO_3560 (O_3560,N_49596,N_47985);
and UO_3561 (O_3561,N_49131,N_48661);
nor UO_3562 (O_3562,N_48821,N_47691);
xnor UO_3563 (O_3563,N_48887,N_49433);
nand UO_3564 (O_3564,N_48428,N_48535);
xnor UO_3565 (O_3565,N_48189,N_49133);
nor UO_3566 (O_3566,N_47541,N_49306);
nand UO_3567 (O_3567,N_49947,N_49330);
and UO_3568 (O_3568,N_47547,N_47858);
or UO_3569 (O_3569,N_48410,N_48672);
nand UO_3570 (O_3570,N_48556,N_49898);
nor UO_3571 (O_3571,N_47925,N_48868);
xor UO_3572 (O_3572,N_49433,N_48985);
xnor UO_3573 (O_3573,N_48252,N_48285);
or UO_3574 (O_3574,N_49913,N_49503);
xor UO_3575 (O_3575,N_48488,N_48965);
and UO_3576 (O_3576,N_49367,N_48807);
and UO_3577 (O_3577,N_47763,N_49741);
and UO_3578 (O_3578,N_47863,N_48094);
and UO_3579 (O_3579,N_48313,N_47893);
nand UO_3580 (O_3580,N_48091,N_47968);
xor UO_3581 (O_3581,N_47844,N_48268);
xnor UO_3582 (O_3582,N_48537,N_49407);
or UO_3583 (O_3583,N_48328,N_47839);
nor UO_3584 (O_3584,N_48754,N_48918);
or UO_3585 (O_3585,N_49570,N_49235);
nand UO_3586 (O_3586,N_48770,N_49552);
nand UO_3587 (O_3587,N_48703,N_49723);
nand UO_3588 (O_3588,N_47580,N_49221);
nand UO_3589 (O_3589,N_49063,N_48311);
xnor UO_3590 (O_3590,N_49458,N_49687);
and UO_3591 (O_3591,N_49484,N_49763);
and UO_3592 (O_3592,N_48706,N_49187);
or UO_3593 (O_3593,N_48873,N_48678);
or UO_3594 (O_3594,N_49330,N_49424);
xor UO_3595 (O_3595,N_49840,N_48788);
or UO_3596 (O_3596,N_48774,N_47945);
nor UO_3597 (O_3597,N_49617,N_49151);
or UO_3598 (O_3598,N_47791,N_48034);
nand UO_3599 (O_3599,N_48248,N_48238);
nor UO_3600 (O_3600,N_48364,N_47552);
or UO_3601 (O_3601,N_48715,N_49335);
or UO_3602 (O_3602,N_48847,N_49785);
nor UO_3603 (O_3603,N_48762,N_49077);
xnor UO_3604 (O_3604,N_48321,N_48989);
xnor UO_3605 (O_3605,N_48441,N_47889);
or UO_3606 (O_3606,N_48577,N_48824);
or UO_3607 (O_3607,N_49451,N_47852);
or UO_3608 (O_3608,N_47818,N_47760);
nor UO_3609 (O_3609,N_48714,N_49187);
nor UO_3610 (O_3610,N_47970,N_49123);
or UO_3611 (O_3611,N_47937,N_47610);
and UO_3612 (O_3612,N_48196,N_48869);
nand UO_3613 (O_3613,N_49403,N_49662);
and UO_3614 (O_3614,N_48207,N_48287);
xor UO_3615 (O_3615,N_49324,N_48837);
nand UO_3616 (O_3616,N_49928,N_48148);
or UO_3617 (O_3617,N_49736,N_47693);
or UO_3618 (O_3618,N_47920,N_49480);
or UO_3619 (O_3619,N_48483,N_49589);
nor UO_3620 (O_3620,N_47897,N_48429);
xnor UO_3621 (O_3621,N_48487,N_47979);
xor UO_3622 (O_3622,N_48772,N_49528);
or UO_3623 (O_3623,N_48149,N_47981);
or UO_3624 (O_3624,N_48171,N_49615);
and UO_3625 (O_3625,N_48948,N_49021);
or UO_3626 (O_3626,N_49509,N_49789);
xor UO_3627 (O_3627,N_49045,N_48355);
or UO_3628 (O_3628,N_48472,N_49041);
xor UO_3629 (O_3629,N_48685,N_49505);
xnor UO_3630 (O_3630,N_47879,N_47745);
nor UO_3631 (O_3631,N_47542,N_49801);
xnor UO_3632 (O_3632,N_49351,N_49269);
nor UO_3633 (O_3633,N_47803,N_48343);
or UO_3634 (O_3634,N_48596,N_47671);
nor UO_3635 (O_3635,N_48253,N_48262);
nor UO_3636 (O_3636,N_47861,N_49510);
nand UO_3637 (O_3637,N_49288,N_48665);
and UO_3638 (O_3638,N_48208,N_49053);
xor UO_3639 (O_3639,N_48340,N_48576);
nor UO_3640 (O_3640,N_49016,N_48226);
and UO_3641 (O_3641,N_48966,N_49151);
and UO_3642 (O_3642,N_47588,N_49757);
and UO_3643 (O_3643,N_48785,N_48469);
nand UO_3644 (O_3644,N_48953,N_48335);
or UO_3645 (O_3645,N_49959,N_47730);
and UO_3646 (O_3646,N_48515,N_49985);
or UO_3647 (O_3647,N_49199,N_48221);
and UO_3648 (O_3648,N_49079,N_48767);
nand UO_3649 (O_3649,N_48259,N_47880);
or UO_3650 (O_3650,N_49206,N_48953);
and UO_3651 (O_3651,N_48637,N_49772);
and UO_3652 (O_3652,N_48960,N_49788);
nor UO_3653 (O_3653,N_48974,N_49856);
nand UO_3654 (O_3654,N_47934,N_49330);
nand UO_3655 (O_3655,N_49848,N_49649);
or UO_3656 (O_3656,N_49359,N_47929);
xor UO_3657 (O_3657,N_49419,N_49321);
nor UO_3658 (O_3658,N_49132,N_49248);
or UO_3659 (O_3659,N_48263,N_49434);
xnor UO_3660 (O_3660,N_48059,N_49325);
or UO_3661 (O_3661,N_48394,N_49687);
nand UO_3662 (O_3662,N_48035,N_49986);
nand UO_3663 (O_3663,N_48772,N_49904);
xnor UO_3664 (O_3664,N_47608,N_48289);
nand UO_3665 (O_3665,N_48952,N_48564);
xor UO_3666 (O_3666,N_47897,N_47503);
xnor UO_3667 (O_3667,N_47859,N_49193);
nor UO_3668 (O_3668,N_47769,N_47677);
nand UO_3669 (O_3669,N_47707,N_48964);
nand UO_3670 (O_3670,N_47706,N_49325);
and UO_3671 (O_3671,N_47592,N_49533);
or UO_3672 (O_3672,N_48765,N_48299);
nand UO_3673 (O_3673,N_48101,N_48951);
nand UO_3674 (O_3674,N_48184,N_49242);
xnor UO_3675 (O_3675,N_48703,N_47663);
or UO_3676 (O_3676,N_48546,N_49887);
nor UO_3677 (O_3677,N_49838,N_49537);
nor UO_3678 (O_3678,N_48412,N_48377);
or UO_3679 (O_3679,N_49831,N_49486);
nand UO_3680 (O_3680,N_47501,N_48122);
nor UO_3681 (O_3681,N_47671,N_48203);
nor UO_3682 (O_3682,N_49852,N_48456);
or UO_3683 (O_3683,N_48453,N_49252);
nand UO_3684 (O_3684,N_47769,N_49273);
xnor UO_3685 (O_3685,N_47803,N_47939);
nor UO_3686 (O_3686,N_49416,N_48204);
nand UO_3687 (O_3687,N_48952,N_49176);
nor UO_3688 (O_3688,N_49498,N_48889);
and UO_3689 (O_3689,N_48234,N_48486);
xnor UO_3690 (O_3690,N_48374,N_49269);
or UO_3691 (O_3691,N_48472,N_48081);
nand UO_3692 (O_3692,N_49638,N_48644);
nor UO_3693 (O_3693,N_48349,N_47623);
xnor UO_3694 (O_3694,N_47925,N_47501);
nand UO_3695 (O_3695,N_49864,N_49528);
nand UO_3696 (O_3696,N_48829,N_49543);
or UO_3697 (O_3697,N_48929,N_47842);
nor UO_3698 (O_3698,N_49657,N_49230);
nor UO_3699 (O_3699,N_49794,N_48954);
xor UO_3700 (O_3700,N_47743,N_48063);
or UO_3701 (O_3701,N_49737,N_49672);
nor UO_3702 (O_3702,N_48618,N_48378);
xor UO_3703 (O_3703,N_47842,N_48881);
nand UO_3704 (O_3704,N_49095,N_49676);
nand UO_3705 (O_3705,N_47712,N_48692);
and UO_3706 (O_3706,N_48030,N_48325);
nor UO_3707 (O_3707,N_49008,N_47880);
and UO_3708 (O_3708,N_48044,N_49598);
nand UO_3709 (O_3709,N_49351,N_48176);
nand UO_3710 (O_3710,N_48946,N_48516);
nand UO_3711 (O_3711,N_49769,N_47833);
nand UO_3712 (O_3712,N_48282,N_48148);
nand UO_3713 (O_3713,N_47622,N_48015);
nor UO_3714 (O_3714,N_48192,N_47701);
nor UO_3715 (O_3715,N_48713,N_48191);
nand UO_3716 (O_3716,N_48936,N_48324);
xnor UO_3717 (O_3717,N_49353,N_49139);
and UO_3718 (O_3718,N_48838,N_49771);
nor UO_3719 (O_3719,N_48511,N_47801);
xnor UO_3720 (O_3720,N_47978,N_49580);
nand UO_3721 (O_3721,N_47754,N_49692);
nor UO_3722 (O_3722,N_49949,N_48048);
or UO_3723 (O_3723,N_49016,N_49484);
or UO_3724 (O_3724,N_48127,N_48473);
or UO_3725 (O_3725,N_49849,N_47516);
nand UO_3726 (O_3726,N_49357,N_47916);
xnor UO_3727 (O_3727,N_48642,N_47827);
nor UO_3728 (O_3728,N_48314,N_48128);
xor UO_3729 (O_3729,N_48261,N_49408);
nand UO_3730 (O_3730,N_47864,N_49834);
and UO_3731 (O_3731,N_48600,N_47772);
and UO_3732 (O_3732,N_48282,N_48888);
nor UO_3733 (O_3733,N_49008,N_49241);
and UO_3734 (O_3734,N_49674,N_49466);
nand UO_3735 (O_3735,N_48494,N_49855);
xnor UO_3736 (O_3736,N_48654,N_47714);
xnor UO_3737 (O_3737,N_49322,N_48588);
or UO_3738 (O_3738,N_49184,N_48128);
and UO_3739 (O_3739,N_48484,N_48169);
nor UO_3740 (O_3740,N_49120,N_48478);
nand UO_3741 (O_3741,N_48547,N_48658);
xnor UO_3742 (O_3742,N_49090,N_49592);
xor UO_3743 (O_3743,N_48623,N_47693);
or UO_3744 (O_3744,N_49430,N_47822);
and UO_3745 (O_3745,N_49485,N_48565);
nand UO_3746 (O_3746,N_47782,N_48184);
nor UO_3747 (O_3747,N_47578,N_48265);
or UO_3748 (O_3748,N_49050,N_47619);
nor UO_3749 (O_3749,N_48548,N_47780);
or UO_3750 (O_3750,N_48050,N_48601);
xnor UO_3751 (O_3751,N_49189,N_49502);
nor UO_3752 (O_3752,N_47993,N_48181);
and UO_3753 (O_3753,N_49218,N_49559);
nor UO_3754 (O_3754,N_49982,N_49906);
or UO_3755 (O_3755,N_49095,N_48885);
xnor UO_3756 (O_3756,N_49988,N_49695);
and UO_3757 (O_3757,N_49031,N_49763);
or UO_3758 (O_3758,N_49830,N_48288);
or UO_3759 (O_3759,N_49345,N_49296);
nand UO_3760 (O_3760,N_49280,N_47988);
nor UO_3761 (O_3761,N_49363,N_48252);
nand UO_3762 (O_3762,N_48677,N_49295);
xor UO_3763 (O_3763,N_48215,N_47892);
nor UO_3764 (O_3764,N_49639,N_48106);
and UO_3765 (O_3765,N_48330,N_47853);
nand UO_3766 (O_3766,N_48011,N_49955);
and UO_3767 (O_3767,N_48787,N_47835);
nand UO_3768 (O_3768,N_49563,N_49140);
nand UO_3769 (O_3769,N_48103,N_49890);
or UO_3770 (O_3770,N_48444,N_47709);
nand UO_3771 (O_3771,N_48651,N_49266);
nor UO_3772 (O_3772,N_49307,N_49492);
xor UO_3773 (O_3773,N_49678,N_48106);
or UO_3774 (O_3774,N_49253,N_48345);
nor UO_3775 (O_3775,N_48071,N_48046);
or UO_3776 (O_3776,N_49645,N_49497);
nand UO_3777 (O_3777,N_49945,N_47510);
and UO_3778 (O_3778,N_47949,N_47830);
xor UO_3779 (O_3779,N_49112,N_49017);
xor UO_3780 (O_3780,N_48885,N_47827);
xnor UO_3781 (O_3781,N_49704,N_49690);
nand UO_3782 (O_3782,N_47919,N_49006);
and UO_3783 (O_3783,N_48999,N_48509);
nor UO_3784 (O_3784,N_47795,N_47517);
or UO_3785 (O_3785,N_49590,N_48242);
or UO_3786 (O_3786,N_49843,N_49751);
xor UO_3787 (O_3787,N_49995,N_48543);
nand UO_3788 (O_3788,N_48108,N_49870);
or UO_3789 (O_3789,N_49380,N_47621);
and UO_3790 (O_3790,N_48170,N_47627);
or UO_3791 (O_3791,N_48542,N_48133);
nor UO_3792 (O_3792,N_49045,N_48397);
and UO_3793 (O_3793,N_49934,N_48319);
xnor UO_3794 (O_3794,N_47768,N_48036);
nand UO_3795 (O_3795,N_49201,N_49061);
or UO_3796 (O_3796,N_48580,N_49344);
nor UO_3797 (O_3797,N_47838,N_47836);
or UO_3798 (O_3798,N_49213,N_48210);
xnor UO_3799 (O_3799,N_48508,N_49107);
or UO_3800 (O_3800,N_49147,N_48973);
nor UO_3801 (O_3801,N_47548,N_49018);
nand UO_3802 (O_3802,N_49375,N_48338);
nor UO_3803 (O_3803,N_48136,N_49582);
nand UO_3804 (O_3804,N_49643,N_49067);
and UO_3805 (O_3805,N_48368,N_48197);
and UO_3806 (O_3806,N_48223,N_48194);
xnor UO_3807 (O_3807,N_49582,N_49697);
nand UO_3808 (O_3808,N_48570,N_48026);
and UO_3809 (O_3809,N_48077,N_48527);
nor UO_3810 (O_3810,N_49721,N_49086);
and UO_3811 (O_3811,N_47954,N_47697);
and UO_3812 (O_3812,N_49968,N_47716);
and UO_3813 (O_3813,N_49617,N_48266);
nand UO_3814 (O_3814,N_48768,N_49473);
xor UO_3815 (O_3815,N_48969,N_49116);
nand UO_3816 (O_3816,N_47585,N_48988);
and UO_3817 (O_3817,N_48614,N_48265);
xnor UO_3818 (O_3818,N_48382,N_49218);
nand UO_3819 (O_3819,N_47911,N_49795);
nand UO_3820 (O_3820,N_48874,N_48057);
xnor UO_3821 (O_3821,N_48800,N_48375);
nand UO_3822 (O_3822,N_49125,N_48856);
xor UO_3823 (O_3823,N_48114,N_49519);
or UO_3824 (O_3824,N_49503,N_48435);
nor UO_3825 (O_3825,N_48052,N_48649);
xnor UO_3826 (O_3826,N_48402,N_49215);
nor UO_3827 (O_3827,N_49317,N_48442);
and UO_3828 (O_3828,N_49072,N_48729);
xnor UO_3829 (O_3829,N_49326,N_49904);
nand UO_3830 (O_3830,N_48009,N_48186);
and UO_3831 (O_3831,N_49165,N_49013);
xnor UO_3832 (O_3832,N_49228,N_49080);
or UO_3833 (O_3833,N_47909,N_48184);
xnor UO_3834 (O_3834,N_47876,N_47807);
nor UO_3835 (O_3835,N_48490,N_48495);
nand UO_3836 (O_3836,N_49391,N_48536);
or UO_3837 (O_3837,N_49566,N_48625);
or UO_3838 (O_3838,N_49903,N_49152);
nand UO_3839 (O_3839,N_48920,N_49070);
nor UO_3840 (O_3840,N_47951,N_47632);
nand UO_3841 (O_3841,N_48779,N_49112);
and UO_3842 (O_3842,N_49069,N_49921);
nand UO_3843 (O_3843,N_48757,N_49331);
or UO_3844 (O_3844,N_47777,N_48159);
nor UO_3845 (O_3845,N_48915,N_48167);
xor UO_3846 (O_3846,N_48584,N_48473);
xor UO_3847 (O_3847,N_48477,N_49795);
nand UO_3848 (O_3848,N_49681,N_48814);
and UO_3849 (O_3849,N_47710,N_47929);
nand UO_3850 (O_3850,N_47563,N_49994);
and UO_3851 (O_3851,N_48429,N_48736);
and UO_3852 (O_3852,N_48028,N_47633);
nand UO_3853 (O_3853,N_48624,N_47717);
and UO_3854 (O_3854,N_47934,N_49885);
or UO_3855 (O_3855,N_48408,N_49181);
and UO_3856 (O_3856,N_47828,N_47858);
xor UO_3857 (O_3857,N_48949,N_49837);
xor UO_3858 (O_3858,N_49205,N_49344);
or UO_3859 (O_3859,N_48488,N_48820);
or UO_3860 (O_3860,N_48640,N_47507);
xor UO_3861 (O_3861,N_49526,N_47934);
nand UO_3862 (O_3862,N_49318,N_48929);
nor UO_3863 (O_3863,N_48605,N_47640);
or UO_3864 (O_3864,N_48151,N_48779);
xnor UO_3865 (O_3865,N_48280,N_48000);
xnor UO_3866 (O_3866,N_49169,N_49601);
or UO_3867 (O_3867,N_48301,N_48236);
nand UO_3868 (O_3868,N_48134,N_49177);
and UO_3869 (O_3869,N_47568,N_48516);
and UO_3870 (O_3870,N_49807,N_48709);
and UO_3871 (O_3871,N_48117,N_48430);
xor UO_3872 (O_3872,N_49128,N_48714);
nand UO_3873 (O_3873,N_47728,N_48599);
nor UO_3874 (O_3874,N_49151,N_48322);
xnor UO_3875 (O_3875,N_49292,N_48291);
nor UO_3876 (O_3876,N_48401,N_48922);
nand UO_3877 (O_3877,N_48282,N_49323);
xor UO_3878 (O_3878,N_48996,N_49247);
or UO_3879 (O_3879,N_48930,N_49246);
and UO_3880 (O_3880,N_48149,N_48821);
and UO_3881 (O_3881,N_48247,N_49986);
nand UO_3882 (O_3882,N_49147,N_48573);
nor UO_3883 (O_3883,N_48292,N_49429);
and UO_3884 (O_3884,N_48832,N_48410);
and UO_3885 (O_3885,N_48572,N_49043);
xor UO_3886 (O_3886,N_48212,N_48793);
nor UO_3887 (O_3887,N_47535,N_48416);
xnor UO_3888 (O_3888,N_48948,N_49453);
nand UO_3889 (O_3889,N_49685,N_49834);
or UO_3890 (O_3890,N_47957,N_47697);
and UO_3891 (O_3891,N_48177,N_48420);
and UO_3892 (O_3892,N_49645,N_47573);
xnor UO_3893 (O_3893,N_49619,N_49795);
or UO_3894 (O_3894,N_47929,N_48810);
nor UO_3895 (O_3895,N_48876,N_48847);
nor UO_3896 (O_3896,N_48585,N_49393);
and UO_3897 (O_3897,N_49739,N_48838);
xnor UO_3898 (O_3898,N_49118,N_48370);
or UO_3899 (O_3899,N_48620,N_48738);
nor UO_3900 (O_3900,N_49498,N_48500);
and UO_3901 (O_3901,N_49959,N_48728);
nand UO_3902 (O_3902,N_48664,N_49492);
or UO_3903 (O_3903,N_48862,N_48273);
nand UO_3904 (O_3904,N_49736,N_49960);
nand UO_3905 (O_3905,N_49105,N_49220);
xor UO_3906 (O_3906,N_49400,N_48320);
nand UO_3907 (O_3907,N_49816,N_48762);
or UO_3908 (O_3908,N_49559,N_48474);
nor UO_3909 (O_3909,N_48709,N_48630);
nand UO_3910 (O_3910,N_49616,N_49498);
nand UO_3911 (O_3911,N_49110,N_49796);
and UO_3912 (O_3912,N_47547,N_48261);
xnor UO_3913 (O_3913,N_49386,N_47532);
and UO_3914 (O_3914,N_47778,N_47981);
or UO_3915 (O_3915,N_48430,N_49466);
or UO_3916 (O_3916,N_47771,N_48034);
and UO_3917 (O_3917,N_48774,N_49233);
and UO_3918 (O_3918,N_49797,N_47925);
or UO_3919 (O_3919,N_49343,N_49047);
nor UO_3920 (O_3920,N_47888,N_48458);
xor UO_3921 (O_3921,N_48477,N_47787);
nor UO_3922 (O_3922,N_47895,N_47525);
nor UO_3923 (O_3923,N_48706,N_48369);
nand UO_3924 (O_3924,N_49482,N_49831);
and UO_3925 (O_3925,N_48656,N_49312);
nand UO_3926 (O_3926,N_48419,N_48885);
nand UO_3927 (O_3927,N_48367,N_48238);
and UO_3928 (O_3928,N_49660,N_48494);
xor UO_3929 (O_3929,N_49924,N_47625);
or UO_3930 (O_3930,N_47904,N_48053);
xor UO_3931 (O_3931,N_49373,N_48738);
or UO_3932 (O_3932,N_49846,N_49434);
and UO_3933 (O_3933,N_48881,N_49274);
nor UO_3934 (O_3934,N_49710,N_49681);
nor UO_3935 (O_3935,N_48220,N_49915);
or UO_3936 (O_3936,N_49802,N_49275);
nor UO_3937 (O_3937,N_49071,N_49318);
and UO_3938 (O_3938,N_48506,N_49277);
or UO_3939 (O_3939,N_47557,N_48378);
and UO_3940 (O_3940,N_47937,N_48540);
nand UO_3941 (O_3941,N_47899,N_49360);
and UO_3942 (O_3942,N_47786,N_48746);
nor UO_3943 (O_3943,N_48675,N_48028);
nand UO_3944 (O_3944,N_49135,N_49761);
nor UO_3945 (O_3945,N_48282,N_48082);
nor UO_3946 (O_3946,N_48415,N_48271);
nand UO_3947 (O_3947,N_47673,N_49070);
nor UO_3948 (O_3948,N_48872,N_49052);
xnor UO_3949 (O_3949,N_48210,N_49797);
nand UO_3950 (O_3950,N_49509,N_49028);
or UO_3951 (O_3951,N_48109,N_49199);
nand UO_3952 (O_3952,N_49380,N_49484);
nand UO_3953 (O_3953,N_48415,N_49752);
xnor UO_3954 (O_3954,N_48894,N_49132);
xor UO_3955 (O_3955,N_49103,N_48884);
or UO_3956 (O_3956,N_48567,N_48850);
and UO_3957 (O_3957,N_49618,N_48422);
nand UO_3958 (O_3958,N_49421,N_47899);
nand UO_3959 (O_3959,N_48689,N_49113);
nand UO_3960 (O_3960,N_47575,N_47706);
nor UO_3961 (O_3961,N_48630,N_49379);
or UO_3962 (O_3962,N_49832,N_49587);
and UO_3963 (O_3963,N_49331,N_49114);
or UO_3964 (O_3964,N_49124,N_49000);
xnor UO_3965 (O_3965,N_49901,N_49284);
or UO_3966 (O_3966,N_48178,N_48046);
nor UO_3967 (O_3967,N_48409,N_47732);
and UO_3968 (O_3968,N_49821,N_48833);
or UO_3969 (O_3969,N_49402,N_49721);
nor UO_3970 (O_3970,N_49879,N_48421);
or UO_3971 (O_3971,N_48624,N_48412);
xor UO_3972 (O_3972,N_49699,N_48879);
xor UO_3973 (O_3973,N_49990,N_49857);
nand UO_3974 (O_3974,N_49331,N_49411);
or UO_3975 (O_3975,N_48015,N_49864);
nor UO_3976 (O_3976,N_48364,N_47907);
xnor UO_3977 (O_3977,N_49045,N_49862);
xnor UO_3978 (O_3978,N_49900,N_47661);
nand UO_3979 (O_3979,N_47940,N_48371);
nand UO_3980 (O_3980,N_49217,N_47875);
xor UO_3981 (O_3981,N_48583,N_48800);
or UO_3982 (O_3982,N_49223,N_48347);
nand UO_3983 (O_3983,N_49269,N_48275);
xnor UO_3984 (O_3984,N_48785,N_48486);
nor UO_3985 (O_3985,N_47555,N_47978);
or UO_3986 (O_3986,N_47522,N_49815);
and UO_3987 (O_3987,N_47937,N_48547);
or UO_3988 (O_3988,N_49794,N_48973);
xor UO_3989 (O_3989,N_48160,N_49171);
and UO_3990 (O_3990,N_48324,N_48332);
and UO_3991 (O_3991,N_48602,N_48105);
and UO_3992 (O_3992,N_49489,N_48137);
xor UO_3993 (O_3993,N_49685,N_48466);
nor UO_3994 (O_3994,N_47953,N_47937);
nor UO_3995 (O_3995,N_47931,N_49387);
nand UO_3996 (O_3996,N_47960,N_49037);
or UO_3997 (O_3997,N_47815,N_49856);
nor UO_3998 (O_3998,N_48109,N_47880);
and UO_3999 (O_3999,N_47568,N_49507);
nand UO_4000 (O_4000,N_48336,N_48397);
xnor UO_4001 (O_4001,N_49698,N_48654);
nor UO_4002 (O_4002,N_48593,N_48013);
and UO_4003 (O_4003,N_48383,N_48947);
and UO_4004 (O_4004,N_48582,N_48144);
or UO_4005 (O_4005,N_47802,N_48918);
nor UO_4006 (O_4006,N_47557,N_48081);
nor UO_4007 (O_4007,N_48375,N_47618);
nor UO_4008 (O_4008,N_48660,N_47971);
xor UO_4009 (O_4009,N_48422,N_48566);
or UO_4010 (O_4010,N_47510,N_48144);
xnor UO_4011 (O_4011,N_49342,N_49791);
xor UO_4012 (O_4012,N_49356,N_48026);
nor UO_4013 (O_4013,N_48286,N_47723);
nand UO_4014 (O_4014,N_48325,N_49740);
nor UO_4015 (O_4015,N_48903,N_49787);
xnor UO_4016 (O_4016,N_47830,N_49445);
and UO_4017 (O_4017,N_48315,N_48460);
and UO_4018 (O_4018,N_49171,N_48203);
nand UO_4019 (O_4019,N_49211,N_49756);
xnor UO_4020 (O_4020,N_49088,N_49073);
nor UO_4021 (O_4021,N_47855,N_48025);
nand UO_4022 (O_4022,N_48670,N_49459);
and UO_4023 (O_4023,N_48108,N_48737);
xor UO_4024 (O_4024,N_48388,N_49882);
nand UO_4025 (O_4025,N_48191,N_48013);
and UO_4026 (O_4026,N_49556,N_48785);
nand UO_4027 (O_4027,N_48501,N_49038);
or UO_4028 (O_4028,N_49070,N_49220);
nor UO_4029 (O_4029,N_49024,N_48091);
or UO_4030 (O_4030,N_49293,N_48809);
xnor UO_4031 (O_4031,N_48822,N_49700);
nand UO_4032 (O_4032,N_48972,N_49834);
nor UO_4033 (O_4033,N_49143,N_49740);
xor UO_4034 (O_4034,N_49007,N_49844);
or UO_4035 (O_4035,N_49403,N_49986);
xor UO_4036 (O_4036,N_49637,N_48141);
nor UO_4037 (O_4037,N_49297,N_48893);
nor UO_4038 (O_4038,N_48813,N_47781);
and UO_4039 (O_4039,N_49418,N_48868);
or UO_4040 (O_4040,N_47649,N_48527);
and UO_4041 (O_4041,N_47859,N_48326);
or UO_4042 (O_4042,N_48543,N_49546);
and UO_4043 (O_4043,N_49713,N_47503);
nand UO_4044 (O_4044,N_48771,N_48465);
xnor UO_4045 (O_4045,N_48638,N_48757);
xor UO_4046 (O_4046,N_49408,N_48744);
or UO_4047 (O_4047,N_48143,N_49573);
or UO_4048 (O_4048,N_48609,N_47860);
and UO_4049 (O_4049,N_49292,N_48173);
nand UO_4050 (O_4050,N_48088,N_49660);
xnor UO_4051 (O_4051,N_49821,N_49373);
xnor UO_4052 (O_4052,N_49274,N_49556);
xnor UO_4053 (O_4053,N_49370,N_49341);
nor UO_4054 (O_4054,N_47714,N_49052);
nor UO_4055 (O_4055,N_49316,N_48214);
and UO_4056 (O_4056,N_49704,N_49803);
xnor UO_4057 (O_4057,N_48148,N_48485);
xnor UO_4058 (O_4058,N_48104,N_48749);
xor UO_4059 (O_4059,N_47641,N_48397);
or UO_4060 (O_4060,N_49710,N_49177);
xor UO_4061 (O_4061,N_48518,N_49102);
or UO_4062 (O_4062,N_48166,N_48389);
xor UO_4063 (O_4063,N_47777,N_48807);
nand UO_4064 (O_4064,N_48241,N_48038);
xor UO_4065 (O_4065,N_48789,N_49719);
nor UO_4066 (O_4066,N_47856,N_49407);
nor UO_4067 (O_4067,N_49630,N_48469);
and UO_4068 (O_4068,N_49032,N_49446);
nand UO_4069 (O_4069,N_48519,N_49558);
nor UO_4070 (O_4070,N_48056,N_48997);
and UO_4071 (O_4071,N_48489,N_49564);
xor UO_4072 (O_4072,N_49184,N_47752);
and UO_4073 (O_4073,N_49130,N_47681);
and UO_4074 (O_4074,N_49577,N_48154);
nor UO_4075 (O_4075,N_48725,N_48796);
xnor UO_4076 (O_4076,N_48342,N_49033);
nor UO_4077 (O_4077,N_48028,N_48365);
xnor UO_4078 (O_4078,N_49665,N_48523);
xnor UO_4079 (O_4079,N_47823,N_48124);
nor UO_4080 (O_4080,N_48678,N_49966);
and UO_4081 (O_4081,N_48629,N_49344);
xnor UO_4082 (O_4082,N_48988,N_48319);
and UO_4083 (O_4083,N_48451,N_47998);
and UO_4084 (O_4084,N_48966,N_47637);
xnor UO_4085 (O_4085,N_48120,N_48906);
nor UO_4086 (O_4086,N_49233,N_48119);
nor UO_4087 (O_4087,N_49636,N_48541);
nand UO_4088 (O_4088,N_49609,N_47624);
xor UO_4089 (O_4089,N_49357,N_49456);
and UO_4090 (O_4090,N_48898,N_49396);
nor UO_4091 (O_4091,N_49230,N_47968);
or UO_4092 (O_4092,N_49204,N_48289);
nand UO_4093 (O_4093,N_47543,N_49605);
nor UO_4094 (O_4094,N_48558,N_48519);
or UO_4095 (O_4095,N_48578,N_48701);
nor UO_4096 (O_4096,N_47791,N_47923);
xnor UO_4097 (O_4097,N_48038,N_49899);
or UO_4098 (O_4098,N_49560,N_49129);
and UO_4099 (O_4099,N_47827,N_47624);
or UO_4100 (O_4100,N_49972,N_48357);
nor UO_4101 (O_4101,N_48682,N_47984);
nor UO_4102 (O_4102,N_47667,N_47534);
or UO_4103 (O_4103,N_49888,N_49913);
nand UO_4104 (O_4104,N_48983,N_47805);
nand UO_4105 (O_4105,N_49801,N_49649);
nand UO_4106 (O_4106,N_48001,N_48037);
and UO_4107 (O_4107,N_49401,N_48111);
nor UO_4108 (O_4108,N_47633,N_47767);
nor UO_4109 (O_4109,N_48913,N_49048);
nand UO_4110 (O_4110,N_48947,N_48626);
nor UO_4111 (O_4111,N_48157,N_48100);
nor UO_4112 (O_4112,N_48027,N_48956);
or UO_4113 (O_4113,N_49347,N_49552);
nand UO_4114 (O_4114,N_49373,N_49555);
and UO_4115 (O_4115,N_48085,N_49244);
nor UO_4116 (O_4116,N_48263,N_48994);
nor UO_4117 (O_4117,N_49948,N_49512);
nand UO_4118 (O_4118,N_49581,N_47547);
or UO_4119 (O_4119,N_49166,N_49193);
or UO_4120 (O_4120,N_48732,N_47597);
nor UO_4121 (O_4121,N_48994,N_49434);
nor UO_4122 (O_4122,N_48388,N_48526);
and UO_4123 (O_4123,N_49574,N_49078);
or UO_4124 (O_4124,N_48338,N_47537);
nor UO_4125 (O_4125,N_48618,N_49373);
xnor UO_4126 (O_4126,N_49292,N_49380);
or UO_4127 (O_4127,N_48056,N_48152);
or UO_4128 (O_4128,N_48892,N_48998);
nor UO_4129 (O_4129,N_47946,N_47643);
xor UO_4130 (O_4130,N_48164,N_48922);
nor UO_4131 (O_4131,N_49476,N_49197);
and UO_4132 (O_4132,N_47901,N_48222);
and UO_4133 (O_4133,N_48827,N_48455);
and UO_4134 (O_4134,N_49534,N_48614);
nand UO_4135 (O_4135,N_48321,N_49100);
and UO_4136 (O_4136,N_47500,N_47893);
nor UO_4137 (O_4137,N_49034,N_47936);
nand UO_4138 (O_4138,N_49567,N_48330);
and UO_4139 (O_4139,N_48777,N_48378);
xor UO_4140 (O_4140,N_47894,N_47884);
nor UO_4141 (O_4141,N_47541,N_49305);
nand UO_4142 (O_4142,N_47747,N_47657);
or UO_4143 (O_4143,N_49651,N_49012);
and UO_4144 (O_4144,N_49898,N_47889);
or UO_4145 (O_4145,N_49695,N_49564);
or UO_4146 (O_4146,N_48066,N_47600);
xnor UO_4147 (O_4147,N_48672,N_49835);
xnor UO_4148 (O_4148,N_49982,N_48307);
nand UO_4149 (O_4149,N_48823,N_49576);
xnor UO_4150 (O_4150,N_48520,N_49231);
nand UO_4151 (O_4151,N_49175,N_49410);
or UO_4152 (O_4152,N_48900,N_47985);
nor UO_4153 (O_4153,N_48864,N_48539);
and UO_4154 (O_4154,N_48676,N_49686);
nor UO_4155 (O_4155,N_47796,N_49769);
nor UO_4156 (O_4156,N_47667,N_48665);
xnor UO_4157 (O_4157,N_48148,N_48182);
and UO_4158 (O_4158,N_49907,N_48700);
nor UO_4159 (O_4159,N_48377,N_49860);
nor UO_4160 (O_4160,N_49659,N_48956);
nor UO_4161 (O_4161,N_49779,N_49492);
or UO_4162 (O_4162,N_49424,N_48926);
xnor UO_4163 (O_4163,N_48865,N_48669);
xor UO_4164 (O_4164,N_48676,N_48113);
and UO_4165 (O_4165,N_47625,N_48758);
nor UO_4166 (O_4166,N_49307,N_49529);
xnor UO_4167 (O_4167,N_49134,N_47545);
and UO_4168 (O_4168,N_48804,N_49257);
xor UO_4169 (O_4169,N_49514,N_48658);
or UO_4170 (O_4170,N_49299,N_47668);
or UO_4171 (O_4171,N_49728,N_48690);
xnor UO_4172 (O_4172,N_49405,N_48641);
xnor UO_4173 (O_4173,N_47592,N_48604);
xor UO_4174 (O_4174,N_49718,N_48605);
or UO_4175 (O_4175,N_48684,N_49027);
nor UO_4176 (O_4176,N_48285,N_48015);
and UO_4177 (O_4177,N_49470,N_49910);
nand UO_4178 (O_4178,N_47774,N_49754);
or UO_4179 (O_4179,N_49267,N_48805);
nor UO_4180 (O_4180,N_48861,N_48677);
nor UO_4181 (O_4181,N_48920,N_48280);
or UO_4182 (O_4182,N_49676,N_47572);
nor UO_4183 (O_4183,N_48030,N_48606);
nand UO_4184 (O_4184,N_47728,N_47755);
and UO_4185 (O_4185,N_47740,N_49506);
nor UO_4186 (O_4186,N_49467,N_49025);
nand UO_4187 (O_4187,N_48690,N_48501);
or UO_4188 (O_4188,N_48570,N_49157);
xor UO_4189 (O_4189,N_49126,N_48871);
xnor UO_4190 (O_4190,N_48395,N_49076);
or UO_4191 (O_4191,N_49302,N_47566);
xor UO_4192 (O_4192,N_49942,N_49706);
nor UO_4193 (O_4193,N_48801,N_49538);
xnor UO_4194 (O_4194,N_48736,N_48791);
nand UO_4195 (O_4195,N_47696,N_48936);
nand UO_4196 (O_4196,N_48977,N_48940);
nor UO_4197 (O_4197,N_48188,N_49485);
or UO_4198 (O_4198,N_49718,N_47747);
or UO_4199 (O_4199,N_49124,N_47761);
nand UO_4200 (O_4200,N_48616,N_49742);
or UO_4201 (O_4201,N_49970,N_49217);
or UO_4202 (O_4202,N_49678,N_49004);
nor UO_4203 (O_4203,N_49843,N_48800);
xnor UO_4204 (O_4204,N_47632,N_47616);
or UO_4205 (O_4205,N_48908,N_47553);
and UO_4206 (O_4206,N_49792,N_49017);
and UO_4207 (O_4207,N_49104,N_49427);
nor UO_4208 (O_4208,N_49394,N_48162);
or UO_4209 (O_4209,N_48043,N_48148);
or UO_4210 (O_4210,N_48793,N_47524);
or UO_4211 (O_4211,N_49038,N_49530);
nand UO_4212 (O_4212,N_49298,N_48803);
or UO_4213 (O_4213,N_49418,N_48798);
nand UO_4214 (O_4214,N_47501,N_48785);
xnor UO_4215 (O_4215,N_48871,N_48583);
xnor UO_4216 (O_4216,N_47852,N_49393);
nand UO_4217 (O_4217,N_48621,N_48107);
or UO_4218 (O_4218,N_49258,N_49873);
xnor UO_4219 (O_4219,N_48322,N_48621);
nand UO_4220 (O_4220,N_49230,N_48437);
nand UO_4221 (O_4221,N_49390,N_48502);
nor UO_4222 (O_4222,N_47544,N_48749);
or UO_4223 (O_4223,N_47659,N_47866);
xnor UO_4224 (O_4224,N_47985,N_49388);
nand UO_4225 (O_4225,N_49741,N_49824);
and UO_4226 (O_4226,N_49023,N_49299);
and UO_4227 (O_4227,N_48136,N_48341);
nor UO_4228 (O_4228,N_48908,N_48299);
nor UO_4229 (O_4229,N_47744,N_47909);
nand UO_4230 (O_4230,N_48202,N_47781);
nand UO_4231 (O_4231,N_48736,N_48543);
nor UO_4232 (O_4232,N_48047,N_48817);
and UO_4233 (O_4233,N_48329,N_48095);
or UO_4234 (O_4234,N_49208,N_48383);
nor UO_4235 (O_4235,N_47650,N_49096);
nor UO_4236 (O_4236,N_49704,N_48391);
nand UO_4237 (O_4237,N_48898,N_47882);
xnor UO_4238 (O_4238,N_48653,N_49826);
xnor UO_4239 (O_4239,N_49629,N_48213);
or UO_4240 (O_4240,N_49791,N_48677);
nand UO_4241 (O_4241,N_48263,N_48337);
and UO_4242 (O_4242,N_49410,N_49756);
xor UO_4243 (O_4243,N_49099,N_47641);
nand UO_4244 (O_4244,N_48942,N_49763);
nor UO_4245 (O_4245,N_49733,N_49457);
nand UO_4246 (O_4246,N_49253,N_48946);
xor UO_4247 (O_4247,N_49347,N_49582);
nand UO_4248 (O_4248,N_47633,N_48279);
nor UO_4249 (O_4249,N_48665,N_48052);
nand UO_4250 (O_4250,N_47757,N_48085);
or UO_4251 (O_4251,N_48503,N_48663);
or UO_4252 (O_4252,N_48644,N_47754);
nor UO_4253 (O_4253,N_49033,N_49591);
and UO_4254 (O_4254,N_48832,N_47897);
nor UO_4255 (O_4255,N_48633,N_47571);
xor UO_4256 (O_4256,N_47639,N_48077);
or UO_4257 (O_4257,N_48425,N_49815);
or UO_4258 (O_4258,N_48910,N_49914);
nand UO_4259 (O_4259,N_48011,N_49141);
xor UO_4260 (O_4260,N_48475,N_48483);
nand UO_4261 (O_4261,N_48694,N_47631);
nand UO_4262 (O_4262,N_49907,N_49123);
nand UO_4263 (O_4263,N_49606,N_49280);
nand UO_4264 (O_4264,N_49009,N_49038);
and UO_4265 (O_4265,N_49941,N_49891);
nand UO_4266 (O_4266,N_47783,N_47924);
and UO_4267 (O_4267,N_47801,N_49292);
nand UO_4268 (O_4268,N_48075,N_48876);
and UO_4269 (O_4269,N_49158,N_47999);
nand UO_4270 (O_4270,N_48431,N_47510);
nand UO_4271 (O_4271,N_49231,N_48703);
nand UO_4272 (O_4272,N_48650,N_49050);
nor UO_4273 (O_4273,N_49605,N_49119);
xor UO_4274 (O_4274,N_48288,N_49181);
and UO_4275 (O_4275,N_47952,N_47849);
nand UO_4276 (O_4276,N_48501,N_49528);
xnor UO_4277 (O_4277,N_49354,N_48902);
xor UO_4278 (O_4278,N_48894,N_48670);
nand UO_4279 (O_4279,N_49487,N_49547);
or UO_4280 (O_4280,N_48104,N_49800);
xor UO_4281 (O_4281,N_48196,N_48698);
xnor UO_4282 (O_4282,N_48999,N_48132);
nor UO_4283 (O_4283,N_48759,N_48766);
xor UO_4284 (O_4284,N_47736,N_49845);
xnor UO_4285 (O_4285,N_48061,N_47524);
and UO_4286 (O_4286,N_48527,N_48758);
or UO_4287 (O_4287,N_49780,N_49709);
and UO_4288 (O_4288,N_49791,N_48433);
nor UO_4289 (O_4289,N_48484,N_47787);
nand UO_4290 (O_4290,N_49547,N_48390);
nor UO_4291 (O_4291,N_49872,N_49800);
and UO_4292 (O_4292,N_48785,N_49256);
xor UO_4293 (O_4293,N_49241,N_49430);
and UO_4294 (O_4294,N_49761,N_48374);
xnor UO_4295 (O_4295,N_49179,N_49110);
nor UO_4296 (O_4296,N_47780,N_49364);
xnor UO_4297 (O_4297,N_48465,N_49756);
and UO_4298 (O_4298,N_49679,N_49540);
nor UO_4299 (O_4299,N_48625,N_49323);
nor UO_4300 (O_4300,N_47739,N_47552);
xnor UO_4301 (O_4301,N_48813,N_49374);
or UO_4302 (O_4302,N_48245,N_49903);
and UO_4303 (O_4303,N_47774,N_49250);
nand UO_4304 (O_4304,N_48167,N_47770);
xnor UO_4305 (O_4305,N_47821,N_47626);
nand UO_4306 (O_4306,N_47789,N_49729);
or UO_4307 (O_4307,N_49476,N_49586);
or UO_4308 (O_4308,N_47894,N_47859);
nand UO_4309 (O_4309,N_48083,N_47759);
nand UO_4310 (O_4310,N_47556,N_49367);
nor UO_4311 (O_4311,N_49639,N_47778);
or UO_4312 (O_4312,N_48572,N_49722);
xnor UO_4313 (O_4313,N_49282,N_47893);
nor UO_4314 (O_4314,N_47860,N_49377);
nor UO_4315 (O_4315,N_49895,N_47578);
xor UO_4316 (O_4316,N_49704,N_48426);
and UO_4317 (O_4317,N_48857,N_48912);
nand UO_4318 (O_4318,N_48742,N_48070);
xnor UO_4319 (O_4319,N_49532,N_48536);
xor UO_4320 (O_4320,N_47560,N_49435);
xor UO_4321 (O_4321,N_48966,N_48357);
or UO_4322 (O_4322,N_48848,N_48704);
nor UO_4323 (O_4323,N_48722,N_49820);
and UO_4324 (O_4324,N_47524,N_48930);
nor UO_4325 (O_4325,N_47945,N_49415);
xor UO_4326 (O_4326,N_48279,N_48885);
nand UO_4327 (O_4327,N_48650,N_49878);
and UO_4328 (O_4328,N_48172,N_47721);
nor UO_4329 (O_4329,N_48292,N_49132);
and UO_4330 (O_4330,N_49436,N_48094);
or UO_4331 (O_4331,N_49279,N_49111);
nand UO_4332 (O_4332,N_49148,N_47612);
or UO_4333 (O_4333,N_47684,N_48811);
nand UO_4334 (O_4334,N_48833,N_48383);
and UO_4335 (O_4335,N_49070,N_48851);
or UO_4336 (O_4336,N_48597,N_48923);
nand UO_4337 (O_4337,N_49480,N_49268);
or UO_4338 (O_4338,N_49476,N_49303);
and UO_4339 (O_4339,N_48220,N_48669);
xor UO_4340 (O_4340,N_48835,N_49694);
nand UO_4341 (O_4341,N_48214,N_48616);
xnor UO_4342 (O_4342,N_48942,N_49928);
nor UO_4343 (O_4343,N_48171,N_47653);
xor UO_4344 (O_4344,N_48171,N_49220);
and UO_4345 (O_4345,N_49918,N_48187);
xor UO_4346 (O_4346,N_49927,N_48025);
nand UO_4347 (O_4347,N_49949,N_49110);
or UO_4348 (O_4348,N_49528,N_48626);
xnor UO_4349 (O_4349,N_49804,N_49308);
or UO_4350 (O_4350,N_48936,N_49693);
or UO_4351 (O_4351,N_48161,N_47668);
nand UO_4352 (O_4352,N_48901,N_48559);
and UO_4353 (O_4353,N_47603,N_47566);
nand UO_4354 (O_4354,N_48213,N_49152);
nand UO_4355 (O_4355,N_48582,N_48982);
xnor UO_4356 (O_4356,N_48972,N_49781);
or UO_4357 (O_4357,N_49220,N_49141);
or UO_4358 (O_4358,N_48925,N_47791);
nor UO_4359 (O_4359,N_49110,N_48717);
nand UO_4360 (O_4360,N_48959,N_49802);
xnor UO_4361 (O_4361,N_49419,N_48784);
nor UO_4362 (O_4362,N_49351,N_48538);
xnor UO_4363 (O_4363,N_48478,N_48353);
or UO_4364 (O_4364,N_49536,N_49907);
xnor UO_4365 (O_4365,N_48943,N_47958);
xor UO_4366 (O_4366,N_49706,N_47980);
nand UO_4367 (O_4367,N_48577,N_47633);
xnor UO_4368 (O_4368,N_49802,N_48639);
nand UO_4369 (O_4369,N_49479,N_49635);
or UO_4370 (O_4370,N_49111,N_49005);
or UO_4371 (O_4371,N_48937,N_48320);
nor UO_4372 (O_4372,N_48676,N_49421);
or UO_4373 (O_4373,N_48137,N_48982);
xnor UO_4374 (O_4374,N_47998,N_48955);
nand UO_4375 (O_4375,N_48933,N_48420);
nand UO_4376 (O_4376,N_49633,N_48777);
nand UO_4377 (O_4377,N_48552,N_48858);
xor UO_4378 (O_4378,N_47981,N_48081);
nor UO_4379 (O_4379,N_48352,N_48448);
nand UO_4380 (O_4380,N_49040,N_48443);
nor UO_4381 (O_4381,N_48938,N_49295);
or UO_4382 (O_4382,N_49442,N_48119);
and UO_4383 (O_4383,N_48912,N_49881);
nand UO_4384 (O_4384,N_49002,N_49192);
nor UO_4385 (O_4385,N_49688,N_48827);
nand UO_4386 (O_4386,N_49601,N_49308);
xnor UO_4387 (O_4387,N_47913,N_47956);
nor UO_4388 (O_4388,N_49935,N_48579);
and UO_4389 (O_4389,N_49246,N_49356);
or UO_4390 (O_4390,N_49380,N_48128);
or UO_4391 (O_4391,N_49146,N_48019);
and UO_4392 (O_4392,N_49211,N_48450);
and UO_4393 (O_4393,N_49853,N_48307);
nand UO_4394 (O_4394,N_49221,N_49845);
nand UO_4395 (O_4395,N_48646,N_47604);
or UO_4396 (O_4396,N_49283,N_48128);
or UO_4397 (O_4397,N_48939,N_49863);
nor UO_4398 (O_4398,N_48046,N_49520);
xnor UO_4399 (O_4399,N_48564,N_49586);
nand UO_4400 (O_4400,N_48223,N_47796);
or UO_4401 (O_4401,N_48984,N_49872);
nand UO_4402 (O_4402,N_49944,N_48757);
xor UO_4403 (O_4403,N_48296,N_49054);
nor UO_4404 (O_4404,N_49227,N_48927);
xnor UO_4405 (O_4405,N_49661,N_48037);
nor UO_4406 (O_4406,N_48573,N_48445);
nor UO_4407 (O_4407,N_49407,N_48916);
xnor UO_4408 (O_4408,N_48966,N_49246);
nand UO_4409 (O_4409,N_49983,N_47837);
nor UO_4410 (O_4410,N_48560,N_49919);
xor UO_4411 (O_4411,N_48392,N_49666);
nor UO_4412 (O_4412,N_47986,N_49408);
and UO_4413 (O_4413,N_48790,N_48140);
and UO_4414 (O_4414,N_49748,N_49497);
nor UO_4415 (O_4415,N_47741,N_47859);
or UO_4416 (O_4416,N_48912,N_48580);
or UO_4417 (O_4417,N_47615,N_48144);
xor UO_4418 (O_4418,N_47585,N_48559);
nor UO_4419 (O_4419,N_49395,N_47513);
and UO_4420 (O_4420,N_48813,N_47658);
xnor UO_4421 (O_4421,N_48191,N_49864);
nand UO_4422 (O_4422,N_47896,N_48887);
xnor UO_4423 (O_4423,N_49478,N_48559);
xnor UO_4424 (O_4424,N_49274,N_48783);
nor UO_4425 (O_4425,N_47515,N_49409);
and UO_4426 (O_4426,N_49859,N_47639);
xnor UO_4427 (O_4427,N_49352,N_49876);
or UO_4428 (O_4428,N_48207,N_49360);
xor UO_4429 (O_4429,N_48706,N_48529);
nor UO_4430 (O_4430,N_49589,N_49243);
xor UO_4431 (O_4431,N_47936,N_49245);
nand UO_4432 (O_4432,N_48641,N_49675);
nand UO_4433 (O_4433,N_49958,N_49543);
nand UO_4434 (O_4434,N_47716,N_48915);
or UO_4435 (O_4435,N_49684,N_47977);
xor UO_4436 (O_4436,N_48141,N_48243);
and UO_4437 (O_4437,N_48969,N_48930);
or UO_4438 (O_4438,N_49576,N_49945);
xor UO_4439 (O_4439,N_49866,N_48960);
nor UO_4440 (O_4440,N_49760,N_48671);
nor UO_4441 (O_4441,N_49020,N_49265);
nand UO_4442 (O_4442,N_48153,N_48195);
or UO_4443 (O_4443,N_49338,N_48089);
nand UO_4444 (O_4444,N_48679,N_48469);
or UO_4445 (O_4445,N_47830,N_49766);
nor UO_4446 (O_4446,N_49450,N_48185);
nor UO_4447 (O_4447,N_49812,N_49198);
and UO_4448 (O_4448,N_48889,N_49566);
xnor UO_4449 (O_4449,N_49387,N_48631);
and UO_4450 (O_4450,N_47510,N_48439);
nor UO_4451 (O_4451,N_47644,N_47943);
nand UO_4452 (O_4452,N_49589,N_49925);
xor UO_4453 (O_4453,N_48289,N_48191);
nor UO_4454 (O_4454,N_49753,N_48042);
and UO_4455 (O_4455,N_48270,N_48636);
nand UO_4456 (O_4456,N_49019,N_47897);
or UO_4457 (O_4457,N_49318,N_47801);
and UO_4458 (O_4458,N_47994,N_48222);
nand UO_4459 (O_4459,N_48368,N_47879);
nand UO_4460 (O_4460,N_48421,N_48341);
and UO_4461 (O_4461,N_48817,N_48807);
and UO_4462 (O_4462,N_49432,N_47925);
nor UO_4463 (O_4463,N_49118,N_48466);
nor UO_4464 (O_4464,N_48706,N_48638);
xnor UO_4465 (O_4465,N_48278,N_48195);
nor UO_4466 (O_4466,N_49136,N_49296);
nor UO_4467 (O_4467,N_47885,N_48425);
or UO_4468 (O_4468,N_48894,N_49978);
nor UO_4469 (O_4469,N_49433,N_48905);
and UO_4470 (O_4470,N_47982,N_48778);
nand UO_4471 (O_4471,N_49736,N_49430);
nor UO_4472 (O_4472,N_49711,N_48088);
nor UO_4473 (O_4473,N_47866,N_49490);
and UO_4474 (O_4474,N_49514,N_49571);
nor UO_4475 (O_4475,N_48149,N_49931);
nor UO_4476 (O_4476,N_48486,N_47660);
nor UO_4477 (O_4477,N_48579,N_48045);
xnor UO_4478 (O_4478,N_47596,N_48918);
nand UO_4479 (O_4479,N_49250,N_47767);
or UO_4480 (O_4480,N_48369,N_48065);
and UO_4481 (O_4481,N_48495,N_48803);
and UO_4482 (O_4482,N_48764,N_48237);
nor UO_4483 (O_4483,N_49352,N_48720);
xnor UO_4484 (O_4484,N_49124,N_48728);
xnor UO_4485 (O_4485,N_48027,N_48217);
nor UO_4486 (O_4486,N_48381,N_49329);
and UO_4487 (O_4487,N_49637,N_48126);
xnor UO_4488 (O_4488,N_49550,N_48677);
nor UO_4489 (O_4489,N_49284,N_47659);
and UO_4490 (O_4490,N_49323,N_48537);
nand UO_4491 (O_4491,N_47548,N_48653);
or UO_4492 (O_4492,N_47666,N_47855);
and UO_4493 (O_4493,N_48839,N_47593);
or UO_4494 (O_4494,N_48549,N_49323);
and UO_4495 (O_4495,N_49813,N_48665);
nand UO_4496 (O_4496,N_49983,N_49228);
and UO_4497 (O_4497,N_49594,N_49339);
or UO_4498 (O_4498,N_49912,N_47543);
xnor UO_4499 (O_4499,N_48978,N_49152);
or UO_4500 (O_4500,N_48739,N_48619);
or UO_4501 (O_4501,N_47937,N_49979);
nand UO_4502 (O_4502,N_49031,N_49245);
xor UO_4503 (O_4503,N_48081,N_47554);
nand UO_4504 (O_4504,N_49639,N_49958);
xnor UO_4505 (O_4505,N_47567,N_48258);
xor UO_4506 (O_4506,N_49509,N_47999);
xnor UO_4507 (O_4507,N_47761,N_48193);
nand UO_4508 (O_4508,N_49826,N_49139);
nor UO_4509 (O_4509,N_49919,N_49416);
xnor UO_4510 (O_4510,N_48441,N_48959);
or UO_4511 (O_4511,N_47729,N_48997);
xor UO_4512 (O_4512,N_48012,N_48351);
nand UO_4513 (O_4513,N_48999,N_49505);
nor UO_4514 (O_4514,N_47727,N_49102);
nand UO_4515 (O_4515,N_49198,N_47967);
and UO_4516 (O_4516,N_48327,N_49380);
nor UO_4517 (O_4517,N_48274,N_49473);
and UO_4518 (O_4518,N_49218,N_49427);
nor UO_4519 (O_4519,N_47814,N_48277);
and UO_4520 (O_4520,N_48019,N_48152);
nor UO_4521 (O_4521,N_47983,N_49906);
and UO_4522 (O_4522,N_48723,N_47588);
or UO_4523 (O_4523,N_48015,N_48370);
nand UO_4524 (O_4524,N_48751,N_48188);
xor UO_4525 (O_4525,N_47822,N_47567);
and UO_4526 (O_4526,N_48791,N_49523);
or UO_4527 (O_4527,N_49900,N_49498);
xnor UO_4528 (O_4528,N_49445,N_48865);
nor UO_4529 (O_4529,N_47661,N_49628);
xor UO_4530 (O_4530,N_49385,N_49695);
xnor UO_4531 (O_4531,N_47626,N_49986);
nor UO_4532 (O_4532,N_48923,N_48262);
xnor UO_4533 (O_4533,N_48457,N_49111);
or UO_4534 (O_4534,N_48341,N_49235);
xor UO_4535 (O_4535,N_49251,N_47785);
xnor UO_4536 (O_4536,N_48951,N_48848);
nand UO_4537 (O_4537,N_48209,N_48281);
nor UO_4538 (O_4538,N_49668,N_49404);
or UO_4539 (O_4539,N_48691,N_49912);
nand UO_4540 (O_4540,N_48919,N_49521);
nand UO_4541 (O_4541,N_48259,N_49324);
or UO_4542 (O_4542,N_47759,N_48788);
and UO_4543 (O_4543,N_49971,N_48291);
xnor UO_4544 (O_4544,N_47609,N_48846);
nor UO_4545 (O_4545,N_49348,N_49708);
xnor UO_4546 (O_4546,N_49829,N_49611);
nor UO_4547 (O_4547,N_49828,N_48460);
nor UO_4548 (O_4548,N_49985,N_47690);
xor UO_4549 (O_4549,N_49243,N_48148);
nand UO_4550 (O_4550,N_47957,N_49714);
nor UO_4551 (O_4551,N_47694,N_48703);
or UO_4552 (O_4552,N_47968,N_47890);
nor UO_4553 (O_4553,N_47542,N_48295);
nand UO_4554 (O_4554,N_49997,N_49052);
xor UO_4555 (O_4555,N_48033,N_48686);
xnor UO_4556 (O_4556,N_49122,N_48417);
nand UO_4557 (O_4557,N_49784,N_49581);
and UO_4558 (O_4558,N_48736,N_49629);
xnor UO_4559 (O_4559,N_48908,N_49346);
nand UO_4560 (O_4560,N_47702,N_49702);
xnor UO_4561 (O_4561,N_48823,N_49096);
or UO_4562 (O_4562,N_48364,N_48347);
nor UO_4563 (O_4563,N_49063,N_48217);
and UO_4564 (O_4564,N_48173,N_49071);
and UO_4565 (O_4565,N_48052,N_47667);
and UO_4566 (O_4566,N_49204,N_47810);
nand UO_4567 (O_4567,N_48613,N_48512);
and UO_4568 (O_4568,N_49630,N_49169);
and UO_4569 (O_4569,N_48606,N_49323);
nand UO_4570 (O_4570,N_49143,N_49855);
and UO_4571 (O_4571,N_48898,N_47850);
nor UO_4572 (O_4572,N_49977,N_48639);
and UO_4573 (O_4573,N_48008,N_49657);
or UO_4574 (O_4574,N_48129,N_49039);
or UO_4575 (O_4575,N_47574,N_48913);
or UO_4576 (O_4576,N_48670,N_48527);
and UO_4577 (O_4577,N_48926,N_49413);
xnor UO_4578 (O_4578,N_48510,N_49442);
and UO_4579 (O_4579,N_49297,N_48458);
nor UO_4580 (O_4580,N_49821,N_48061);
or UO_4581 (O_4581,N_49949,N_47672);
xor UO_4582 (O_4582,N_49599,N_47622);
or UO_4583 (O_4583,N_48712,N_48131);
nand UO_4584 (O_4584,N_47551,N_48987);
and UO_4585 (O_4585,N_48718,N_48408);
xor UO_4586 (O_4586,N_47791,N_47901);
or UO_4587 (O_4587,N_48711,N_49954);
xor UO_4588 (O_4588,N_48110,N_49751);
and UO_4589 (O_4589,N_47918,N_48557);
nor UO_4590 (O_4590,N_48074,N_49946);
nor UO_4591 (O_4591,N_47610,N_48370);
or UO_4592 (O_4592,N_49619,N_48821);
nor UO_4593 (O_4593,N_47682,N_47599);
xnor UO_4594 (O_4594,N_49921,N_48966);
nand UO_4595 (O_4595,N_48311,N_48775);
nor UO_4596 (O_4596,N_47956,N_49915);
or UO_4597 (O_4597,N_49079,N_47651);
or UO_4598 (O_4598,N_47837,N_48734);
or UO_4599 (O_4599,N_49072,N_47849);
nor UO_4600 (O_4600,N_49556,N_48747);
and UO_4601 (O_4601,N_48540,N_49885);
and UO_4602 (O_4602,N_49512,N_48417);
and UO_4603 (O_4603,N_48036,N_48570);
and UO_4604 (O_4604,N_48504,N_49645);
xnor UO_4605 (O_4605,N_49545,N_49638);
or UO_4606 (O_4606,N_47876,N_49425);
xnor UO_4607 (O_4607,N_49307,N_48695);
xor UO_4608 (O_4608,N_49144,N_49635);
and UO_4609 (O_4609,N_48879,N_49425);
nor UO_4610 (O_4610,N_48275,N_48161);
and UO_4611 (O_4611,N_49724,N_49177);
and UO_4612 (O_4612,N_47872,N_47527);
xnor UO_4613 (O_4613,N_48290,N_49810);
xor UO_4614 (O_4614,N_48726,N_47959);
nand UO_4615 (O_4615,N_49869,N_48657);
nor UO_4616 (O_4616,N_48251,N_48509);
nor UO_4617 (O_4617,N_48755,N_49223);
and UO_4618 (O_4618,N_47628,N_49728);
nor UO_4619 (O_4619,N_49919,N_49807);
nand UO_4620 (O_4620,N_49469,N_47593);
xnor UO_4621 (O_4621,N_48014,N_48800);
xnor UO_4622 (O_4622,N_47562,N_48522);
or UO_4623 (O_4623,N_48257,N_49740);
and UO_4624 (O_4624,N_49798,N_49642);
nor UO_4625 (O_4625,N_49803,N_48448);
and UO_4626 (O_4626,N_48524,N_48271);
xor UO_4627 (O_4627,N_48292,N_48112);
xnor UO_4628 (O_4628,N_49288,N_48556);
nor UO_4629 (O_4629,N_47578,N_49131);
nor UO_4630 (O_4630,N_49402,N_47565);
nand UO_4631 (O_4631,N_48761,N_48280);
and UO_4632 (O_4632,N_47870,N_49857);
and UO_4633 (O_4633,N_48231,N_49226);
xor UO_4634 (O_4634,N_49615,N_49077);
xnor UO_4635 (O_4635,N_48722,N_47900);
or UO_4636 (O_4636,N_49768,N_47690);
nand UO_4637 (O_4637,N_48555,N_47595);
or UO_4638 (O_4638,N_49073,N_48732);
or UO_4639 (O_4639,N_49473,N_49735);
nor UO_4640 (O_4640,N_47765,N_47595);
or UO_4641 (O_4641,N_47658,N_49397);
nor UO_4642 (O_4642,N_47894,N_48856);
or UO_4643 (O_4643,N_49553,N_48455);
nand UO_4644 (O_4644,N_48292,N_49501);
or UO_4645 (O_4645,N_47700,N_48546);
nand UO_4646 (O_4646,N_49717,N_48100);
xor UO_4647 (O_4647,N_47692,N_47785);
nor UO_4648 (O_4648,N_47673,N_49012);
nor UO_4649 (O_4649,N_49403,N_47823);
xnor UO_4650 (O_4650,N_49885,N_48058);
nand UO_4651 (O_4651,N_48695,N_49373);
and UO_4652 (O_4652,N_48980,N_48751);
nor UO_4653 (O_4653,N_49405,N_48960);
nand UO_4654 (O_4654,N_48654,N_47743);
nor UO_4655 (O_4655,N_49162,N_48364);
nor UO_4656 (O_4656,N_48649,N_48048);
and UO_4657 (O_4657,N_47900,N_49512);
xor UO_4658 (O_4658,N_48994,N_48383);
and UO_4659 (O_4659,N_48850,N_49057);
nor UO_4660 (O_4660,N_49031,N_47819);
and UO_4661 (O_4661,N_48988,N_47853);
and UO_4662 (O_4662,N_48048,N_48862);
xnor UO_4663 (O_4663,N_49170,N_48407);
and UO_4664 (O_4664,N_49648,N_49224);
nor UO_4665 (O_4665,N_49666,N_48123);
xor UO_4666 (O_4666,N_48747,N_48419);
or UO_4667 (O_4667,N_48159,N_49742);
nor UO_4668 (O_4668,N_49580,N_49668);
or UO_4669 (O_4669,N_48138,N_49967);
xor UO_4670 (O_4670,N_49389,N_49898);
or UO_4671 (O_4671,N_48279,N_47565);
and UO_4672 (O_4672,N_48560,N_48132);
nor UO_4673 (O_4673,N_48249,N_48119);
xor UO_4674 (O_4674,N_48951,N_49175);
xor UO_4675 (O_4675,N_49426,N_48694);
or UO_4676 (O_4676,N_47720,N_49639);
nor UO_4677 (O_4677,N_48908,N_48770);
or UO_4678 (O_4678,N_49049,N_48669);
or UO_4679 (O_4679,N_49817,N_48839);
and UO_4680 (O_4680,N_48101,N_48362);
nor UO_4681 (O_4681,N_48410,N_47712);
or UO_4682 (O_4682,N_47523,N_47652);
and UO_4683 (O_4683,N_48981,N_49493);
and UO_4684 (O_4684,N_48019,N_48631);
nor UO_4685 (O_4685,N_47735,N_49790);
nand UO_4686 (O_4686,N_47506,N_47836);
nand UO_4687 (O_4687,N_47557,N_49793);
or UO_4688 (O_4688,N_47791,N_49837);
nand UO_4689 (O_4689,N_48236,N_47735);
nand UO_4690 (O_4690,N_49761,N_48217);
or UO_4691 (O_4691,N_48723,N_48854);
or UO_4692 (O_4692,N_49798,N_47801);
xor UO_4693 (O_4693,N_48626,N_48058);
and UO_4694 (O_4694,N_47595,N_47749);
nand UO_4695 (O_4695,N_48934,N_49400);
and UO_4696 (O_4696,N_47766,N_47922);
or UO_4697 (O_4697,N_47905,N_48017);
nand UO_4698 (O_4698,N_49601,N_49232);
and UO_4699 (O_4699,N_47988,N_48369);
or UO_4700 (O_4700,N_49054,N_48044);
and UO_4701 (O_4701,N_48937,N_49872);
nor UO_4702 (O_4702,N_49480,N_47747);
or UO_4703 (O_4703,N_48092,N_48273);
xnor UO_4704 (O_4704,N_49480,N_48149);
nor UO_4705 (O_4705,N_47892,N_48526);
and UO_4706 (O_4706,N_49898,N_49896);
nor UO_4707 (O_4707,N_47859,N_48753);
xor UO_4708 (O_4708,N_49131,N_47556);
nand UO_4709 (O_4709,N_49387,N_48340);
nand UO_4710 (O_4710,N_49543,N_48749);
xor UO_4711 (O_4711,N_49222,N_49933);
and UO_4712 (O_4712,N_48113,N_49360);
xnor UO_4713 (O_4713,N_48588,N_49787);
xnor UO_4714 (O_4714,N_48911,N_49785);
and UO_4715 (O_4715,N_47560,N_48731);
nor UO_4716 (O_4716,N_49737,N_48236);
xnor UO_4717 (O_4717,N_49026,N_48649);
or UO_4718 (O_4718,N_48395,N_49712);
xor UO_4719 (O_4719,N_48155,N_49186);
or UO_4720 (O_4720,N_49488,N_48035);
nand UO_4721 (O_4721,N_48052,N_49016);
and UO_4722 (O_4722,N_47794,N_49850);
nand UO_4723 (O_4723,N_48481,N_48997);
xnor UO_4724 (O_4724,N_49022,N_47540);
nand UO_4725 (O_4725,N_48623,N_48095);
xor UO_4726 (O_4726,N_49441,N_49501);
xnor UO_4727 (O_4727,N_48307,N_49270);
nor UO_4728 (O_4728,N_47601,N_48855);
and UO_4729 (O_4729,N_49965,N_48084);
xor UO_4730 (O_4730,N_49748,N_48648);
nand UO_4731 (O_4731,N_48254,N_49064);
xor UO_4732 (O_4732,N_48290,N_48182);
xnor UO_4733 (O_4733,N_47941,N_48494);
nand UO_4734 (O_4734,N_48546,N_49622);
nor UO_4735 (O_4735,N_49532,N_47747);
and UO_4736 (O_4736,N_48348,N_48127);
nor UO_4737 (O_4737,N_48012,N_48832);
nor UO_4738 (O_4738,N_49889,N_49880);
nor UO_4739 (O_4739,N_49013,N_47501);
xor UO_4740 (O_4740,N_47562,N_49788);
nand UO_4741 (O_4741,N_47805,N_49605);
nand UO_4742 (O_4742,N_48706,N_48111);
xnor UO_4743 (O_4743,N_49083,N_47648);
and UO_4744 (O_4744,N_48979,N_48912);
xnor UO_4745 (O_4745,N_48153,N_47924);
nand UO_4746 (O_4746,N_49034,N_49925);
and UO_4747 (O_4747,N_49553,N_48805);
nand UO_4748 (O_4748,N_48332,N_49040);
nor UO_4749 (O_4749,N_49116,N_49542);
xnor UO_4750 (O_4750,N_49527,N_49922);
xnor UO_4751 (O_4751,N_49962,N_47579);
nand UO_4752 (O_4752,N_48833,N_48104);
and UO_4753 (O_4753,N_48057,N_49431);
xnor UO_4754 (O_4754,N_48020,N_47712);
nand UO_4755 (O_4755,N_48654,N_49001);
or UO_4756 (O_4756,N_48089,N_49109);
or UO_4757 (O_4757,N_48171,N_48520);
xnor UO_4758 (O_4758,N_47722,N_48519);
nand UO_4759 (O_4759,N_48205,N_49791);
nand UO_4760 (O_4760,N_49768,N_49547);
or UO_4761 (O_4761,N_48884,N_48591);
nand UO_4762 (O_4762,N_48540,N_48034);
and UO_4763 (O_4763,N_48956,N_48891);
xnor UO_4764 (O_4764,N_49301,N_48574);
xor UO_4765 (O_4765,N_48229,N_48934);
nand UO_4766 (O_4766,N_49362,N_48404);
and UO_4767 (O_4767,N_48182,N_49194);
and UO_4768 (O_4768,N_48968,N_48532);
nand UO_4769 (O_4769,N_48749,N_47882);
and UO_4770 (O_4770,N_48030,N_49023);
or UO_4771 (O_4771,N_49504,N_49355);
and UO_4772 (O_4772,N_49876,N_49631);
xnor UO_4773 (O_4773,N_48142,N_47944);
or UO_4774 (O_4774,N_47803,N_48422);
xor UO_4775 (O_4775,N_48817,N_47669);
xnor UO_4776 (O_4776,N_48638,N_47707);
and UO_4777 (O_4777,N_47869,N_48811);
nand UO_4778 (O_4778,N_49309,N_49345);
or UO_4779 (O_4779,N_48877,N_49900);
nor UO_4780 (O_4780,N_49949,N_48131);
or UO_4781 (O_4781,N_48676,N_47632);
and UO_4782 (O_4782,N_47740,N_47960);
or UO_4783 (O_4783,N_48016,N_48639);
nand UO_4784 (O_4784,N_47619,N_49017);
nand UO_4785 (O_4785,N_49452,N_49722);
nand UO_4786 (O_4786,N_47846,N_49998);
nor UO_4787 (O_4787,N_48483,N_48188);
xnor UO_4788 (O_4788,N_49387,N_49869);
xnor UO_4789 (O_4789,N_48196,N_48793);
nand UO_4790 (O_4790,N_48113,N_48265);
nand UO_4791 (O_4791,N_47599,N_48665);
nand UO_4792 (O_4792,N_49614,N_49296);
nand UO_4793 (O_4793,N_47505,N_49753);
nor UO_4794 (O_4794,N_49291,N_48647);
nand UO_4795 (O_4795,N_48693,N_48599);
and UO_4796 (O_4796,N_47893,N_49012);
and UO_4797 (O_4797,N_49038,N_48057);
nand UO_4798 (O_4798,N_49009,N_48945);
nor UO_4799 (O_4799,N_49596,N_48114);
xor UO_4800 (O_4800,N_47520,N_49429);
and UO_4801 (O_4801,N_48510,N_48208);
and UO_4802 (O_4802,N_49296,N_48253);
or UO_4803 (O_4803,N_49696,N_49400);
nand UO_4804 (O_4804,N_49674,N_49685);
or UO_4805 (O_4805,N_47683,N_48877);
nor UO_4806 (O_4806,N_47874,N_48575);
xor UO_4807 (O_4807,N_48761,N_49766);
xor UO_4808 (O_4808,N_49231,N_47613);
xor UO_4809 (O_4809,N_49946,N_47616);
and UO_4810 (O_4810,N_48581,N_47673);
xor UO_4811 (O_4811,N_47576,N_47920);
nand UO_4812 (O_4812,N_49702,N_47849);
xnor UO_4813 (O_4813,N_48405,N_49300);
xnor UO_4814 (O_4814,N_47728,N_48232);
nor UO_4815 (O_4815,N_48451,N_49811);
xnor UO_4816 (O_4816,N_49678,N_48479);
nor UO_4817 (O_4817,N_48909,N_48918);
nor UO_4818 (O_4818,N_48086,N_49954);
nor UO_4819 (O_4819,N_49118,N_48721);
xnor UO_4820 (O_4820,N_49754,N_48600);
or UO_4821 (O_4821,N_48485,N_48447);
or UO_4822 (O_4822,N_47794,N_47814);
and UO_4823 (O_4823,N_47834,N_48088);
and UO_4824 (O_4824,N_49080,N_47640);
nand UO_4825 (O_4825,N_48071,N_48376);
and UO_4826 (O_4826,N_49958,N_48006);
xnor UO_4827 (O_4827,N_49763,N_48045);
xnor UO_4828 (O_4828,N_47713,N_48863);
or UO_4829 (O_4829,N_48601,N_49718);
and UO_4830 (O_4830,N_47685,N_49336);
xnor UO_4831 (O_4831,N_48887,N_48078);
or UO_4832 (O_4832,N_48097,N_49268);
nor UO_4833 (O_4833,N_48753,N_49025);
nor UO_4834 (O_4834,N_47540,N_48674);
xor UO_4835 (O_4835,N_47980,N_49064);
nand UO_4836 (O_4836,N_48915,N_47964);
or UO_4837 (O_4837,N_48238,N_48853);
nand UO_4838 (O_4838,N_48101,N_48819);
xor UO_4839 (O_4839,N_49022,N_47591);
nand UO_4840 (O_4840,N_48523,N_48580);
nor UO_4841 (O_4841,N_49315,N_48892);
or UO_4842 (O_4842,N_47913,N_48163);
nor UO_4843 (O_4843,N_48725,N_49460);
xor UO_4844 (O_4844,N_47595,N_49290);
xor UO_4845 (O_4845,N_48505,N_47699);
and UO_4846 (O_4846,N_49850,N_47556);
and UO_4847 (O_4847,N_48550,N_49913);
xor UO_4848 (O_4848,N_49823,N_49532);
and UO_4849 (O_4849,N_49473,N_47733);
nor UO_4850 (O_4850,N_47800,N_47598);
or UO_4851 (O_4851,N_49202,N_49574);
and UO_4852 (O_4852,N_47968,N_47994);
nor UO_4853 (O_4853,N_48774,N_48113);
or UO_4854 (O_4854,N_49838,N_49530);
and UO_4855 (O_4855,N_49796,N_49530);
nand UO_4856 (O_4856,N_49266,N_49250);
xnor UO_4857 (O_4857,N_49901,N_49902);
xnor UO_4858 (O_4858,N_49619,N_49720);
and UO_4859 (O_4859,N_48883,N_49063);
xnor UO_4860 (O_4860,N_48734,N_48539);
and UO_4861 (O_4861,N_49875,N_49090);
or UO_4862 (O_4862,N_47655,N_49288);
xor UO_4863 (O_4863,N_49575,N_48141);
xnor UO_4864 (O_4864,N_47782,N_47707);
xnor UO_4865 (O_4865,N_49214,N_47727);
nand UO_4866 (O_4866,N_48505,N_47555);
or UO_4867 (O_4867,N_48178,N_47828);
nand UO_4868 (O_4868,N_47717,N_48688);
nor UO_4869 (O_4869,N_49370,N_47590);
nor UO_4870 (O_4870,N_48708,N_48538);
and UO_4871 (O_4871,N_49663,N_49107);
and UO_4872 (O_4872,N_48227,N_48658);
or UO_4873 (O_4873,N_48395,N_47673);
or UO_4874 (O_4874,N_49255,N_47926);
nor UO_4875 (O_4875,N_49569,N_48603);
nand UO_4876 (O_4876,N_48508,N_47722);
or UO_4877 (O_4877,N_49370,N_47869);
nand UO_4878 (O_4878,N_49476,N_48349);
xnor UO_4879 (O_4879,N_49386,N_47586);
nand UO_4880 (O_4880,N_47589,N_47878);
or UO_4881 (O_4881,N_48179,N_47796);
and UO_4882 (O_4882,N_48384,N_49235);
or UO_4883 (O_4883,N_49163,N_49342);
nand UO_4884 (O_4884,N_49196,N_48123);
nand UO_4885 (O_4885,N_48825,N_49313);
xnor UO_4886 (O_4886,N_48414,N_49704);
xor UO_4887 (O_4887,N_48788,N_47765);
and UO_4888 (O_4888,N_48954,N_49328);
nand UO_4889 (O_4889,N_48467,N_49811);
or UO_4890 (O_4890,N_49110,N_49953);
nor UO_4891 (O_4891,N_48922,N_48422);
xnor UO_4892 (O_4892,N_48130,N_47830);
xor UO_4893 (O_4893,N_49342,N_48211);
xor UO_4894 (O_4894,N_48012,N_49950);
or UO_4895 (O_4895,N_47575,N_47596);
nand UO_4896 (O_4896,N_48318,N_48403);
nor UO_4897 (O_4897,N_48047,N_48418);
nor UO_4898 (O_4898,N_49551,N_49145);
nor UO_4899 (O_4899,N_49582,N_48633);
nand UO_4900 (O_4900,N_47941,N_47663);
nand UO_4901 (O_4901,N_47524,N_49007);
xnor UO_4902 (O_4902,N_47950,N_48209);
or UO_4903 (O_4903,N_49364,N_49991);
nand UO_4904 (O_4904,N_49349,N_49741);
and UO_4905 (O_4905,N_48920,N_49947);
and UO_4906 (O_4906,N_48653,N_47996);
nand UO_4907 (O_4907,N_48840,N_49013);
nor UO_4908 (O_4908,N_48993,N_48341);
nand UO_4909 (O_4909,N_48448,N_48601);
xor UO_4910 (O_4910,N_47670,N_48339);
or UO_4911 (O_4911,N_48714,N_47849);
and UO_4912 (O_4912,N_49739,N_49085);
nand UO_4913 (O_4913,N_49716,N_48197);
nor UO_4914 (O_4914,N_47986,N_47502);
nand UO_4915 (O_4915,N_48246,N_47919);
xnor UO_4916 (O_4916,N_48620,N_48772);
nand UO_4917 (O_4917,N_47995,N_49324);
and UO_4918 (O_4918,N_49498,N_49886);
xnor UO_4919 (O_4919,N_49186,N_47614);
nand UO_4920 (O_4920,N_48534,N_48088);
xnor UO_4921 (O_4921,N_49436,N_48577);
xnor UO_4922 (O_4922,N_48516,N_48243);
or UO_4923 (O_4923,N_48012,N_49733);
nor UO_4924 (O_4924,N_49061,N_48127);
nand UO_4925 (O_4925,N_48555,N_48549);
and UO_4926 (O_4926,N_49018,N_48720);
xnor UO_4927 (O_4927,N_49461,N_48646);
nor UO_4928 (O_4928,N_48043,N_49360);
nand UO_4929 (O_4929,N_48627,N_48000);
nand UO_4930 (O_4930,N_49739,N_48632);
xnor UO_4931 (O_4931,N_49481,N_47510);
xor UO_4932 (O_4932,N_49958,N_49345);
xnor UO_4933 (O_4933,N_47924,N_49253);
nand UO_4934 (O_4934,N_48534,N_48868);
nor UO_4935 (O_4935,N_49854,N_48639);
xnor UO_4936 (O_4936,N_47818,N_47527);
nand UO_4937 (O_4937,N_49453,N_48006);
or UO_4938 (O_4938,N_49570,N_48599);
or UO_4939 (O_4939,N_49881,N_49078);
or UO_4940 (O_4940,N_49410,N_49805);
nor UO_4941 (O_4941,N_48145,N_48515);
xnor UO_4942 (O_4942,N_49146,N_48089);
nor UO_4943 (O_4943,N_48123,N_48486);
nand UO_4944 (O_4944,N_49893,N_49125);
nor UO_4945 (O_4945,N_47693,N_47530);
and UO_4946 (O_4946,N_49073,N_48881);
and UO_4947 (O_4947,N_48745,N_49680);
xnor UO_4948 (O_4948,N_48763,N_49607);
nand UO_4949 (O_4949,N_49006,N_49809);
xor UO_4950 (O_4950,N_47559,N_48679);
xor UO_4951 (O_4951,N_48019,N_48969);
nor UO_4952 (O_4952,N_47824,N_49807);
and UO_4953 (O_4953,N_48588,N_48559);
and UO_4954 (O_4954,N_47789,N_47520);
or UO_4955 (O_4955,N_48326,N_48164);
and UO_4956 (O_4956,N_49684,N_49246);
and UO_4957 (O_4957,N_47799,N_49100);
and UO_4958 (O_4958,N_49082,N_48307);
nor UO_4959 (O_4959,N_49690,N_49443);
xor UO_4960 (O_4960,N_48902,N_48414);
nand UO_4961 (O_4961,N_49875,N_49844);
xor UO_4962 (O_4962,N_48880,N_49345);
and UO_4963 (O_4963,N_48319,N_47829);
nand UO_4964 (O_4964,N_49780,N_48098);
nor UO_4965 (O_4965,N_48430,N_49339);
nand UO_4966 (O_4966,N_48582,N_48165);
xor UO_4967 (O_4967,N_49004,N_49076);
and UO_4968 (O_4968,N_48539,N_49612);
nand UO_4969 (O_4969,N_47902,N_49490);
or UO_4970 (O_4970,N_47709,N_49924);
and UO_4971 (O_4971,N_48687,N_47903);
nand UO_4972 (O_4972,N_48303,N_47723);
nor UO_4973 (O_4973,N_48691,N_48098);
and UO_4974 (O_4974,N_49944,N_49697);
nand UO_4975 (O_4975,N_49803,N_49893);
and UO_4976 (O_4976,N_49021,N_49787);
or UO_4977 (O_4977,N_48443,N_48065);
and UO_4978 (O_4978,N_48978,N_49811);
xor UO_4979 (O_4979,N_47637,N_48494);
xnor UO_4980 (O_4980,N_49634,N_49987);
or UO_4981 (O_4981,N_48553,N_49531);
nor UO_4982 (O_4982,N_47753,N_48841);
xor UO_4983 (O_4983,N_49717,N_48190);
nor UO_4984 (O_4984,N_48521,N_48434);
or UO_4985 (O_4985,N_49030,N_49443);
or UO_4986 (O_4986,N_49144,N_49189);
nor UO_4987 (O_4987,N_48038,N_49557);
nor UO_4988 (O_4988,N_48259,N_48208);
nand UO_4989 (O_4989,N_49910,N_48719);
or UO_4990 (O_4990,N_49091,N_48468);
nor UO_4991 (O_4991,N_48108,N_47763);
and UO_4992 (O_4992,N_48227,N_49625);
and UO_4993 (O_4993,N_48538,N_49775);
nor UO_4994 (O_4994,N_49267,N_48491);
and UO_4995 (O_4995,N_49936,N_48466);
or UO_4996 (O_4996,N_49581,N_49815);
nor UO_4997 (O_4997,N_48463,N_49646);
and UO_4998 (O_4998,N_49283,N_48734);
nor UO_4999 (O_4999,N_47698,N_48058);
endmodule