module basic_3000_30000_3500_6_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1316,In_2958);
and U1 (N_1,In_323,In_207);
and U2 (N_2,In_991,In_347);
and U3 (N_3,In_1488,In_729);
and U4 (N_4,In_2237,In_1778);
nand U5 (N_5,In_1032,In_2143);
nand U6 (N_6,In_1255,In_2541);
and U7 (N_7,In_2447,In_1320);
nand U8 (N_8,In_496,In_1214);
or U9 (N_9,In_1241,In_448);
nand U10 (N_10,In_380,In_953);
nor U11 (N_11,In_523,In_2966);
nand U12 (N_12,In_2062,In_1556);
and U13 (N_13,In_1981,In_295);
nor U14 (N_14,In_583,In_2863);
nand U15 (N_15,In_2654,In_130);
or U16 (N_16,In_1597,In_1650);
or U17 (N_17,In_2262,In_132);
or U18 (N_18,In_518,In_1667);
nand U19 (N_19,In_1949,In_1194);
nand U20 (N_20,In_1141,In_279);
or U21 (N_21,In_2699,In_2683);
nor U22 (N_22,In_670,In_1232);
nor U23 (N_23,In_1852,In_71);
nor U24 (N_24,In_170,In_504);
nand U25 (N_25,In_1847,In_2770);
nand U26 (N_26,In_2599,In_2805);
and U27 (N_27,In_1441,In_1383);
nor U28 (N_28,In_1156,In_2038);
or U29 (N_29,In_482,In_1358);
or U30 (N_30,In_1076,In_2222);
nand U31 (N_31,In_2276,In_2955);
nand U32 (N_32,In_1388,In_2943);
and U33 (N_33,In_882,In_1581);
or U34 (N_34,In_928,In_686);
nor U35 (N_35,In_1716,In_1897);
nor U36 (N_36,In_8,In_2421);
nand U37 (N_37,In_1630,In_2025);
or U38 (N_38,In_1702,In_1038);
and U39 (N_39,In_2641,In_575);
nand U40 (N_40,In_2383,In_341);
nor U41 (N_41,In_2175,In_2295);
or U42 (N_42,In_2497,In_2921);
nor U43 (N_43,In_1152,In_233);
nand U44 (N_44,In_2328,In_1363);
and U45 (N_45,In_338,In_2407);
and U46 (N_46,In_1309,In_1013);
and U47 (N_47,In_423,In_663);
nand U48 (N_48,In_36,In_321);
or U49 (N_49,In_1012,In_2564);
or U50 (N_50,In_318,In_1052);
xnor U51 (N_51,In_1522,In_1535);
nor U52 (N_52,In_960,In_319);
nand U53 (N_53,In_1059,In_501);
nor U54 (N_54,In_2484,In_2493);
nand U55 (N_55,In_1960,In_846);
nor U56 (N_56,In_1478,In_2610);
or U57 (N_57,In_2259,In_1935);
or U58 (N_58,In_82,In_2186);
or U59 (N_59,In_20,In_2913);
nand U60 (N_60,In_111,In_2481);
nand U61 (N_61,In_1396,In_1503);
nor U62 (N_62,In_393,In_906);
nand U63 (N_63,In_1860,In_488);
nor U64 (N_64,In_700,In_2364);
nand U65 (N_65,In_577,In_2324);
nand U66 (N_66,In_2495,In_1527);
nand U67 (N_67,In_1861,In_241);
nor U68 (N_68,In_2064,In_2539);
nor U69 (N_69,In_181,In_2831);
and U70 (N_70,In_2692,In_2666);
nand U71 (N_71,In_838,In_1516);
nand U72 (N_72,In_356,In_376);
and U73 (N_73,In_1323,In_7);
nand U74 (N_74,In_2629,In_203);
and U75 (N_75,In_1885,In_1364);
nand U76 (N_76,In_1741,In_2631);
and U77 (N_77,In_653,In_1372);
nor U78 (N_78,In_1898,In_2698);
nand U79 (N_79,In_1709,In_1896);
and U80 (N_80,In_751,In_1017);
or U81 (N_81,In_2331,In_2658);
and U82 (N_82,In_2679,In_461);
and U83 (N_83,In_183,In_146);
nand U84 (N_84,In_238,In_1464);
and U85 (N_85,In_1746,In_320);
nor U86 (N_86,In_1791,In_1979);
and U87 (N_87,In_1412,In_1728);
nand U88 (N_88,In_1835,In_1924);
nand U89 (N_89,In_1011,In_337);
nand U90 (N_90,In_721,In_497);
or U91 (N_91,In_41,In_1116);
or U92 (N_92,In_1457,In_1439);
nor U93 (N_93,In_1287,In_2884);
and U94 (N_94,In_680,In_1449);
and U95 (N_95,In_192,In_1656);
and U96 (N_96,In_528,In_2147);
nand U97 (N_97,In_2243,In_1227);
and U98 (N_98,In_788,In_1124);
or U99 (N_99,In_1968,In_1657);
and U100 (N_100,In_1181,In_939);
and U101 (N_101,In_1917,In_2305);
and U102 (N_102,In_2487,In_2846);
nor U103 (N_103,In_1054,In_2338);
or U104 (N_104,In_120,In_901);
or U105 (N_105,In_976,In_24);
nand U106 (N_106,In_1334,In_2090);
and U107 (N_107,In_268,In_2317);
and U108 (N_108,In_2581,In_2720);
and U109 (N_109,In_1212,In_2194);
nand U110 (N_110,In_1675,In_1224);
nor U111 (N_111,In_2053,In_2323);
and U112 (N_112,In_1873,In_1617);
and U113 (N_113,In_956,In_1515);
nand U114 (N_114,In_2440,In_1958);
nand U115 (N_115,In_2207,In_1405);
or U116 (N_116,In_764,In_2393);
nor U117 (N_117,In_2466,In_437);
xor U118 (N_118,In_1109,In_2802);
or U119 (N_119,In_1566,In_1);
nor U120 (N_120,In_848,In_2696);
nor U121 (N_121,In_1520,In_1739);
and U122 (N_122,In_981,In_2069);
nor U123 (N_123,In_1421,In_2675);
and U124 (N_124,In_1609,In_1631);
nor U125 (N_125,In_163,In_1558);
nor U126 (N_126,In_2568,In_2617);
or U127 (N_127,In_2188,In_2330);
nor U128 (N_128,In_2479,In_1679);
nor U129 (N_129,In_2915,In_1344);
nor U130 (N_130,In_2063,In_2678);
xor U131 (N_131,In_656,In_463);
and U132 (N_132,In_1285,In_821);
and U133 (N_133,In_2359,In_405);
nand U134 (N_134,In_880,In_629);
and U135 (N_135,In_2174,In_313);
nor U136 (N_136,In_407,In_761);
and U137 (N_137,In_1254,In_562);
and U138 (N_138,In_718,In_2711);
or U139 (N_139,In_2755,In_2146);
and U140 (N_140,In_839,In_1889);
and U141 (N_141,In_119,In_2280);
or U142 (N_142,In_2343,In_2990);
nor U143 (N_143,In_1502,In_1524);
nand U144 (N_144,In_414,In_974);
and U145 (N_145,In_93,In_280);
and U146 (N_146,In_209,In_2847);
nor U147 (N_147,In_449,In_638);
nand U148 (N_148,In_322,In_1654);
and U149 (N_149,In_576,In_516);
nand U150 (N_150,In_1559,In_2505);
nand U151 (N_151,In_2042,In_1508);
nand U152 (N_152,In_2577,In_277);
nand U153 (N_153,In_1833,In_1962);
nand U154 (N_154,In_2432,In_1993);
nor U155 (N_155,In_1411,In_1711);
nor U156 (N_156,In_2853,In_2782);
and U157 (N_157,In_1967,In_1242);
or U158 (N_158,In_2234,In_315);
nand U159 (N_159,In_1366,In_554);
nor U160 (N_160,In_1591,In_1643);
or U161 (N_161,In_2307,In_1918);
nor U162 (N_162,In_1223,In_881);
or U163 (N_163,In_102,In_1348);
nor U164 (N_164,In_2303,In_1909);
and U165 (N_165,In_2904,In_858);
or U166 (N_166,In_2832,In_929);
nand U167 (N_167,In_2368,In_1910);
nand U168 (N_168,In_1990,In_2521);
or U169 (N_169,In_1063,In_2443);
nand U170 (N_170,In_2257,In_1921);
or U171 (N_171,In_1121,In_73);
nor U172 (N_172,In_2185,In_1066);
and U173 (N_173,In_895,In_1901);
nand U174 (N_174,In_246,In_2034);
and U175 (N_175,In_2604,In_401);
nand U176 (N_176,In_440,In_1519);
nand U177 (N_177,In_1186,In_1273);
and U178 (N_178,In_1932,In_2653);
or U179 (N_179,In_2879,In_2972);
and U180 (N_180,In_1282,In_2089);
nor U181 (N_181,In_1119,In_1030);
nor U182 (N_182,In_2296,In_1072);
nor U183 (N_183,In_77,In_2530);
or U184 (N_184,In_1367,In_1178);
or U185 (N_185,In_1151,In_2714);
and U186 (N_186,In_2367,In_2784);
and U187 (N_187,In_2967,In_525);
or U188 (N_188,In_478,In_914);
nand U189 (N_189,In_2489,In_1134);
and U190 (N_190,In_2474,In_2544);
nand U191 (N_191,In_735,In_616);
or U192 (N_192,In_1331,In_1983);
nor U193 (N_193,In_1532,In_1837);
and U194 (N_194,In_2642,In_1089);
nor U195 (N_195,In_2223,In_775);
and U196 (N_196,In_972,In_35);
or U197 (N_197,In_652,In_1740);
nand U198 (N_198,In_983,In_2420);
or U199 (N_199,In_624,In_544);
and U200 (N_200,In_1380,In_74);
nor U201 (N_201,In_1601,In_211);
or U202 (N_202,In_2938,In_2003);
nand U203 (N_203,In_526,In_2468);
nand U204 (N_204,In_2289,In_1568);
nand U205 (N_205,In_2900,In_1482);
nand U206 (N_206,In_1341,In_1187);
nor U207 (N_207,In_874,In_2817);
and U208 (N_208,In_1813,In_2217);
nor U209 (N_209,In_685,In_1957);
or U210 (N_210,In_2140,In_2159);
and U211 (N_211,In_2115,In_298);
or U212 (N_212,In_1096,In_2632);
nand U213 (N_213,In_455,In_2964);
or U214 (N_214,In_1942,In_794);
nand U215 (N_215,In_1928,In_1705);
nand U216 (N_216,In_699,In_187);
nor U217 (N_217,In_458,In_600);
or U218 (N_218,In_1540,In_2937);
and U219 (N_219,In_1080,In_987);
and U220 (N_220,In_2485,In_1298);
nand U221 (N_221,In_2464,In_2412);
nor U222 (N_222,In_493,In_2781);
xor U223 (N_223,In_2872,In_2744);
and U224 (N_224,In_2706,In_2139);
nand U225 (N_225,In_314,In_2814);
and U226 (N_226,In_456,In_509);
or U227 (N_227,In_1701,In_459);
nor U228 (N_228,In_539,In_1599);
or U229 (N_229,In_1284,In_1459);
nor U230 (N_230,In_2794,In_1004);
nand U231 (N_231,In_2138,In_1218);
nor U232 (N_232,In_495,In_2538);
nand U233 (N_233,In_2766,In_1948);
nor U234 (N_234,In_1826,In_2970);
nand U235 (N_235,In_1770,In_408);
and U236 (N_236,In_1259,In_2860);
nor U237 (N_237,In_58,In_2342);
nor U238 (N_238,In_1700,In_2601);
and U239 (N_239,In_473,In_2912);
nand U240 (N_240,In_2780,In_2561);
and U241 (N_241,In_310,In_2216);
or U242 (N_242,In_2974,In_2645);
or U243 (N_243,In_1678,In_2812);
or U244 (N_244,In_1755,In_2015);
nor U245 (N_245,In_222,In_1822);
or U246 (N_246,In_253,In_1048);
nand U247 (N_247,In_2401,In_911);
and U248 (N_248,In_2154,In_167);
and U249 (N_249,In_2997,In_1868);
and U250 (N_250,In_918,In_2946);
and U251 (N_251,In_2056,In_326);
nor U252 (N_252,In_951,In_390);
or U253 (N_253,In_2681,In_1359);
nand U254 (N_254,In_164,In_2459);
and U255 (N_255,In_113,In_1712);
and U256 (N_256,In_2861,In_4);
or U257 (N_257,In_195,In_1000);
and U258 (N_258,In_244,In_1723);
nand U259 (N_259,In_2792,In_864);
and U260 (N_260,In_845,In_2798);
or U261 (N_261,In_1317,In_2369);
xor U262 (N_262,In_1021,In_898);
and U263 (N_263,In_2523,In_1192);
nor U264 (N_264,In_522,In_768);
nor U265 (N_265,In_300,In_2700);
nand U266 (N_266,In_1451,In_840);
or U267 (N_267,In_1913,In_273);
nand U268 (N_268,In_2287,In_732);
or U269 (N_269,In_1694,In_83);
nor U270 (N_270,In_2131,In_2293);
or U271 (N_271,In_153,In_2932);
nor U272 (N_272,In_2179,In_627);
nand U273 (N_273,In_127,In_1114);
nor U274 (N_274,In_2624,In_177);
nand U275 (N_275,In_2928,In_1773);
and U276 (N_276,In_2375,In_349);
and U277 (N_277,In_2156,In_2124);
or U278 (N_278,In_235,In_6);
nor U279 (N_279,In_806,In_1277);
nand U280 (N_280,In_1229,In_1789);
and U281 (N_281,In_2376,In_2987);
nand U282 (N_282,In_1008,In_2619);
nor U283 (N_283,In_1257,In_945);
and U284 (N_284,In_173,In_2907);
or U285 (N_285,In_849,In_919);
nand U286 (N_286,In_419,In_1279);
nand U287 (N_287,In_573,In_1984);
nand U288 (N_288,In_667,In_1870);
and U289 (N_289,In_902,In_2811);
nand U290 (N_290,In_1768,In_859);
or U291 (N_291,In_1454,In_1416);
or U292 (N_292,In_0,In_2400);
xnor U293 (N_293,In_494,In_558);
nor U294 (N_294,In_382,In_2476);
and U295 (N_295,In_2540,In_2739);
nand U296 (N_296,In_400,In_2646);
and U297 (N_297,In_1668,In_65);
nor U298 (N_298,In_725,In_1304);
nor U299 (N_299,In_276,In_1293);
or U300 (N_300,In_62,In_1049);
nand U301 (N_301,In_2892,In_1531);
nand U302 (N_302,In_891,In_2531);
nor U303 (N_303,In_876,In_538);
nor U304 (N_304,In_2751,In_61);
nand U305 (N_305,In_1009,In_1560);
nor U306 (N_306,In_13,In_2233);
nand U307 (N_307,In_483,In_487);
or U308 (N_308,In_2051,In_2891);
nand U309 (N_309,In_801,In_2697);
nand U310 (N_310,In_2193,In_863);
nor U311 (N_311,In_1002,In_1828);
nor U312 (N_312,In_66,In_1533);
and U313 (N_313,In_1809,In_1043);
or U314 (N_314,In_2123,In_1238);
xnor U315 (N_315,In_1148,In_142);
nand U316 (N_316,In_17,In_2933);
nor U317 (N_317,In_787,In_1975);
and U318 (N_318,In_293,In_451);
nor U319 (N_319,In_1857,In_1829);
and U320 (N_320,In_2086,In_1300);
nand U321 (N_321,In_590,In_2041);
nor U322 (N_322,In_2591,In_500);
nor U323 (N_323,In_2837,In_1904);
and U324 (N_324,In_2727,In_1107);
xnor U325 (N_325,In_1624,In_1360);
and U326 (N_326,In_422,In_2026);
or U327 (N_327,In_1613,In_2512);
and U328 (N_328,In_2985,In_893);
or U329 (N_329,In_1602,In_827);
or U330 (N_330,In_2880,In_1862);
nand U331 (N_331,In_1506,In_2477);
nand U332 (N_332,In_740,In_1492);
or U333 (N_333,In_2644,In_604);
nand U334 (N_334,In_202,In_770);
nand U335 (N_335,In_1839,In_1351);
and U336 (N_336,In_543,In_831);
nand U337 (N_337,In_2450,In_2993);
and U338 (N_338,In_189,In_2475);
or U339 (N_339,In_2524,In_2265);
and U340 (N_340,In_2701,In_2463);
nand U341 (N_341,In_2906,In_1274);
nor U342 (N_342,In_1940,In_1501);
nand U343 (N_343,In_1154,In_224);
or U344 (N_344,In_1045,In_585);
and U345 (N_345,In_2453,In_379);
and U346 (N_346,In_2118,In_1169);
or U347 (N_347,In_677,In_1737);
and U348 (N_348,In_2559,In_598);
nor U349 (N_349,In_1426,In_2326);
nand U350 (N_350,In_560,In_2592);
nand U351 (N_351,In_535,In_2918);
and U352 (N_352,In_2862,In_1925);
nor U353 (N_353,In_671,In_1088);
nand U354 (N_354,In_1163,In_1068);
nor U355 (N_355,In_890,In_2554);
or U356 (N_356,In_2874,In_143);
nor U357 (N_357,In_1562,In_2660);
and U358 (N_358,In_1382,In_2796);
nor U359 (N_359,In_48,In_1338);
nor U360 (N_360,In_852,In_2048);
nor U361 (N_361,In_1903,In_1097);
and U362 (N_362,In_2602,In_2612);
nand U363 (N_363,In_1295,In_1754);
nand U364 (N_364,In_989,In_1392);
nor U365 (N_365,In_923,In_348);
and U366 (N_366,In_709,In_582);
nor U367 (N_367,In_2529,In_2353);
and U368 (N_368,In_2441,In_1135);
nor U369 (N_369,In_92,In_851);
or U370 (N_370,In_1687,In_373);
and U371 (N_371,In_622,In_1954);
nand U372 (N_372,In_2002,In_1168);
nor U373 (N_373,In_2079,In_1757);
nor U374 (N_374,In_2398,In_1725);
or U375 (N_375,In_2325,In_1371);
nand U376 (N_376,In_672,In_2108);
nor U377 (N_377,In_809,In_1391);
or U378 (N_378,In_578,In_2881);
and U379 (N_379,In_1406,In_332);
nand U380 (N_380,In_1931,In_80);
or U381 (N_381,In_947,In_1093);
and U382 (N_382,In_225,In_1950);
or U383 (N_383,In_269,In_1007);
and U384 (N_384,In_2870,In_2598);
and U385 (N_385,In_2828,In_530);
and U386 (N_386,In_1393,In_780);
and U387 (N_387,In_1251,In_2865);
nor U388 (N_388,In_28,In_648);
and U389 (N_389,In_2647,In_613);
and U390 (N_390,In_1646,In_2926);
nand U391 (N_391,In_2190,In_2843);
nor U392 (N_392,In_1500,In_2998);
and U393 (N_393,In_257,In_1291);
or U394 (N_394,In_1666,In_2472);
and U395 (N_395,In_820,In_1445);
nor U396 (N_396,In_2702,In_1022);
nor U397 (N_397,In_2999,In_1537);
nor U398 (N_398,In_1638,In_2099);
or U399 (N_399,In_1016,In_2348);
or U400 (N_400,In_2885,In_2894);
nor U401 (N_401,In_1422,In_1081);
or U402 (N_402,In_1235,In_1926);
nor U403 (N_403,In_602,In_210);
or U404 (N_404,In_247,In_1131);
nor U405 (N_405,In_1892,In_1819);
nor U406 (N_406,In_2284,In_108);
nor U407 (N_407,In_1489,In_229);
and U408 (N_408,In_1497,In_157);
nand U409 (N_409,In_1884,In_264);
or U410 (N_410,In_2868,In_2120);
nor U411 (N_411,In_1404,In_2600);
and U412 (N_412,In_49,In_1051);
nor U413 (N_413,In_2016,In_2403);
nor U414 (N_414,In_2628,In_129);
and U415 (N_415,In_2141,In_200);
nor U416 (N_416,In_570,In_620);
and U417 (N_417,In_1683,In_2001);
or U418 (N_418,In_1108,In_1792);
nor U419 (N_419,In_160,In_666);
xor U420 (N_420,In_1197,In_1015);
nand U421 (N_421,In_2183,In_2925);
nand U422 (N_422,In_1225,In_1234);
and U423 (N_423,In_1024,In_191);
and U424 (N_424,In_2742,In_2327);
or U425 (N_425,In_900,In_2801);
nand U426 (N_426,In_542,In_1461);
or U427 (N_427,In_2431,In_2571);
or U428 (N_428,In_2731,In_2576);
nor U429 (N_429,In_1120,In_1525);
and U430 (N_430,In_2068,In_2256);
nand U431 (N_431,In_1673,In_2589);
or U432 (N_432,In_2844,In_2128);
or U433 (N_433,In_2806,In_1982);
nand U434 (N_434,In_2236,In_1243);
or U435 (N_435,In_2671,In_1173);
and U436 (N_436,In_2335,In_541);
or U437 (N_437,In_1794,In_2077);
nor U438 (N_438,In_536,In_559);
or U439 (N_439,In_1644,In_2558);
and U440 (N_440,In_2830,In_1487);
and U441 (N_441,In_1322,In_932);
and U442 (N_442,In_2028,In_2310);
nor U443 (N_443,In_1659,In_2685);
nor U444 (N_444,In_2840,In_2643);
nor U445 (N_445,In_674,In_1872);
and U446 (N_446,In_2515,In_937);
nand U447 (N_447,In_2674,In_1155);
nand U448 (N_448,In_1713,In_2729);
and U449 (N_449,In_252,In_1945);
or U450 (N_450,In_1217,In_426);
and U451 (N_451,In_694,In_232);
or U452 (N_452,In_823,In_118);
or U453 (N_453,In_1625,In_2212);
nor U454 (N_454,In_2130,In_812);
nor U455 (N_455,In_2867,In_1340);
or U456 (N_456,In_1026,In_841);
or U457 (N_457,In_2756,In_383);
or U458 (N_458,In_29,In_2723);
or U459 (N_459,In_2341,In_1423);
nand U460 (N_460,In_1463,In_219);
or U461 (N_461,In_1018,In_297);
and U462 (N_462,In_464,In_773);
and U463 (N_463,In_2979,In_1425);
nand U464 (N_464,In_114,In_660);
or U465 (N_465,In_545,In_769);
nor U466 (N_466,In_579,In_2730);
or U467 (N_467,In_2980,In_2808);
nor U468 (N_468,In_1696,In_2842);
and U469 (N_469,In_2292,In_2081);
nor U470 (N_470,In_2164,In_634);
nor U471 (N_471,In_135,In_2785);
or U472 (N_472,In_1832,In_563);
xnor U473 (N_473,In_2267,In_978);
or U474 (N_474,In_1133,In_2890);
nor U475 (N_475,In_1965,In_2804);
and U476 (N_476,In_871,In_2772);
or U477 (N_477,In_1398,In_2752);
and U478 (N_478,In_1572,In_954);
and U479 (N_479,In_1479,In_2300);
nor U480 (N_480,In_619,In_2834);
and U481 (N_481,In_1495,In_2247);
nor U482 (N_482,In_1389,In_2114);
or U483 (N_483,In_762,In_333);
and U484 (N_484,In_1653,In_2542);
nand U485 (N_485,In_2594,In_100);
xor U486 (N_486,In_2722,In_2461);
and U487 (N_487,In_218,In_1112);
or U488 (N_488,In_979,In_1484);
nor U489 (N_489,In_1571,In_2931);
and U490 (N_490,In_359,In_2119);
and U491 (N_491,In_1838,In_1978);
nor U492 (N_492,In_1056,In_137);
nor U493 (N_493,In_2226,In_1786);
nor U494 (N_494,In_1268,In_772);
and U495 (N_495,In_2649,In_1321);
and U496 (N_496,In_457,In_2430);
nand U497 (N_497,In_1377,In_655);
and U498 (N_498,In_2774,In_2910);
nor U499 (N_499,In_1199,In_2920);
or U500 (N_500,In_766,In_1150);
or U501 (N_501,In_1036,In_1598);
nor U502 (N_502,In_1325,In_1719);
nand U503 (N_503,In_1210,In_1900);
nand U504 (N_504,In_1458,In_2651);
and U505 (N_505,In_121,In_1470);
nand U506 (N_506,In_1266,In_1205);
nor U507 (N_507,In_2178,In_39);
nand U508 (N_508,In_1628,In_870);
or U509 (N_509,In_687,In_2365);
or U510 (N_510,In_1887,In_1939);
or U511 (N_511,In_2791,In_950);
nand U512 (N_512,In_917,In_2195);
or U513 (N_513,In_2390,In_728);
nand U514 (N_514,In_308,In_973);
nor U515 (N_515,In_2127,In_964);
nor U516 (N_516,In_1866,In_1437);
or U517 (N_517,In_1697,In_328);
nand U518 (N_518,In_2315,In_2426);
or U519 (N_519,In_1991,In_564);
or U520 (N_520,In_2503,In_1677);
and U521 (N_521,In_242,In_2302);
xor U522 (N_522,In_2082,In_2737);
nand U523 (N_523,In_2715,In_606);
and U524 (N_524,In_944,In_290);
or U525 (N_525,In_2513,In_1289);
nand U526 (N_526,In_443,In_2029);
nand U527 (N_527,In_262,In_626);
nor U528 (N_528,In_2471,In_1247);
nand U529 (N_529,In_485,In_2169);
nor U530 (N_530,In_519,In_2725);
and U531 (N_531,In_2112,In_703);
nor U532 (N_532,In_599,In_669);
or U533 (N_533,In_1606,In_1082);
and U534 (N_534,In_2281,In_1246);
or U535 (N_535,In_800,In_2919);
nor U536 (N_536,In_1128,In_2627);
xnor U537 (N_537,In_2935,In_2519);
nor U538 (N_538,In_1762,In_2707);
nand U539 (N_539,In_1167,In_172);
or U540 (N_540,In_2268,In_2829);
nor U541 (N_541,In_1637,In_588);
or U542 (N_542,In_2903,In_75);
nor U543 (N_543,In_2445,In_1550);
or U544 (N_544,In_757,In_466);
nor U545 (N_545,In_2011,In_208);
nand U546 (N_546,In_1662,In_2961);
nor U547 (N_547,In_294,In_1742);
and U548 (N_548,In_1339,In_2940);
nor U549 (N_549,In_551,In_2747);
and U550 (N_550,In_1118,In_139);
and U551 (N_551,In_52,In_126);
nor U552 (N_552,In_116,In_834);
and U553 (N_553,In_650,In_2635);
nor U554 (N_554,In_2623,In_2067);
and U555 (N_555,In_1104,In_912);
nor U556 (N_556,In_970,In_631);
and U557 (N_557,In_549,In_1435);
and U558 (N_558,In_1810,In_2873);
xor U559 (N_559,In_1122,In_1191);
and U560 (N_560,In_367,In_1584);
xor U561 (N_561,In_2827,In_425);
and U562 (N_562,In_2374,In_508);
nand U563 (N_563,In_591,In_1305);
and U564 (N_564,In_915,In_1816);
nor U565 (N_565,In_2930,In_360);
nand U566 (N_566,In_186,In_2270);
and U567 (N_567,In_417,In_597);
nor U568 (N_568,In_2822,In_1596);
or U569 (N_569,In_514,In_1966);
or U570 (N_570,In_1270,In_2992);
and U571 (N_571,In_2984,In_2013);
or U572 (N_572,In_1882,In_1410);
and U573 (N_573,In_2311,In_1438);
nor U574 (N_574,In_2360,In_2444);
nand U575 (N_575,In_1185,In_611);
and U576 (N_576,In_1142,In_1297);
and U577 (N_577,In_2486,In_1061);
and U578 (N_578,In_1171,In_2469);
and U579 (N_579,In_2934,In_311);
nor U580 (N_580,In_1684,In_1450);
nor U581 (N_581,In_2963,In_30);
nor U582 (N_582,In_1621,In_339);
and U583 (N_583,In_2117,In_1718);
or U584 (N_584,In_2250,In_2269);
or U585 (N_585,In_2818,In_1342);
and U586 (N_586,In_2137,In_665);
or U587 (N_587,In_87,In_1845);
nor U588 (N_588,In_850,In_1446);
or U589 (N_589,In_995,In_2264);
nor U590 (N_590,In_1874,In_2640);
nor U591 (N_591,In_1782,In_742);
nand U592 (N_592,In_696,In_1374);
or U593 (N_593,In_467,In_134);
nor U594 (N_594,In_644,In_1370);
nand U595 (N_595,In_2550,In_2261);
nor U596 (N_596,In_2357,In_817);
or U597 (N_597,In_819,In_2951);
xnor U598 (N_598,In_291,In_771);
nor U599 (N_599,In_2319,In_505);
and U600 (N_600,In_2387,In_1823);
and U601 (N_601,In_353,In_2496);
and U602 (N_602,In_1400,In_1849);
nor U603 (N_603,In_1064,In_2528);
and U604 (N_604,In_595,In_2012);
nor U605 (N_605,In_2162,In_479);
nand U606 (N_606,In_2150,In_2165);
nand U607 (N_607,In_2522,In_1269);
or U608 (N_608,In_2975,In_2982);
or U609 (N_609,In_765,In_2911);
nor U610 (N_610,In_1985,In_2916);
and U611 (N_611,In_835,In_1264);
nor U612 (N_612,In_1206,In_1390);
or U613 (N_613,In_2093,In_690);
nor U614 (N_614,In_2449,In_1611);
and U615 (N_615,In_2621,In_125);
nor U616 (N_616,In_2351,In_1256);
nand U617 (N_617,In_1756,In_2996);
nor U618 (N_618,In_1956,In_2848);
nor U619 (N_619,In_1039,In_2201);
or U620 (N_620,In_2346,In_10);
and U621 (N_621,In_2251,In_2121);
or U622 (N_622,In_894,In_506);
or U623 (N_623,In_1751,In_1615);
nor U624 (N_624,In_2952,In_1938);
nand U625 (N_625,In_1165,In_2914);
or U626 (N_626,In_1147,In_305);
nand U627 (N_627,In_2241,In_1290);
and U628 (N_628,In_2976,In_1442);
or U629 (N_629,In_865,In_1361);
nor U630 (N_630,In_1117,In_1005);
nand U631 (N_631,In_1726,In_2525);
or U632 (N_632,In_1804,In_1475);
xor U633 (N_633,In_2995,In_2710);
nand U634 (N_634,In_2083,In_1505);
and U635 (N_635,In_2494,In_2149);
nand U636 (N_636,In_1731,In_1564);
or U637 (N_637,In_2578,In_1840);
or U638 (N_638,In_713,In_2102);
and U639 (N_639,In_1020,In_2570);
nor U640 (N_640,In_774,In_1094);
or U641 (N_641,In_1162,In_975);
nor U642 (N_642,In_1262,In_1477);
and U643 (N_643,In_708,In_1843);
and U644 (N_644,In_352,In_808);
nand U645 (N_645,In_1933,In_2759);
and U646 (N_646,In_688,In_1929);
or U647 (N_647,In_2436,In_1760);
and U648 (N_648,In_2684,In_2392);
and U649 (N_649,In_1415,In_1028);
nand U650 (N_650,In_2422,In_1436);
nor U651 (N_651,In_1201,In_57);
nand U652 (N_652,In_1448,In_1570);
or U653 (N_653,In_1612,In_197);
and U654 (N_654,In_1399,In_2010);
nor U655 (N_655,In_1720,In_2452);
or U656 (N_656,In_998,In_2562);
nor U657 (N_657,In_580,In_1552);
and U658 (N_658,In_1146,In_1357);
nor U659 (N_659,In_424,In_930);
and U660 (N_660,In_1953,In_370);
and U661 (N_661,In_1444,In_2498);
nand U662 (N_662,In_2517,In_2586);
nor U663 (N_663,In_2071,In_2689);
and U664 (N_664,In_22,In_1772);
nand U665 (N_665,In_1207,In_1513);
nand U666 (N_666,In_1378,In_1787);
nor U667 (N_667,In_1541,In_1626);
nand U668 (N_668,In_1517,In_2111);
nor U669 (N_669,In_1176,In_1785);
and U670 (N_670,In_1417,In_2414);
nand U671 (N_671,In_346,In_384);
nand U672 (N_672,In_196,In_101);
nor U673 (N_673,In_1595,In_1419);
nand U674 (N_674,In_1691,In_1174);
xor U675 (N_675,In_2661,In_147);
nand U676 (N_676,In_2682,In_784);
nor U677 (N_677,In_452,In_434);
nor U678 (N_678,In_1802,In_2616);
and U679 (N_679,In_1641,In_1911);
and U680 (N_680,In_396,In_1999);
nand U681 (N_681,In_43,In_465);
nor U682 (N_682,In_1623,In_1672);
nand U683 (N_683,In_2388,In_1443);
or U684 (N_684,In_2213,In_1906);
nor U685 (N_685,In_2386,In_1230);
or U686 (N_686,In_53,In_2394);
nand U687 (N_687,In_441,In_2446);
and U688 (N_688,In_2978,In_1029);
and U689 (N_689,In_1512,In_2786);
or U690 (N_690,In_909,In_1428);
nand U691 (N_691,In_391,In_566);
and U692 (N_692,In_1518,In_737);
nor U693 (N_693,In_96,In_2363);
nand U694 (N_694,In_1160,In_2883);
nor U695 (N_695,In_2084,In_418);
nand U696 (N_696,In_1510,In_1542);
and U697 (N_697,In_2332,In_2799);
and U698 (N_698,In_1777,In_2936);
and U699 (N_699,In_1111,In_736);
or U700 (N_700,In_968,In_682);
or U701 (N_701,In_807,In_1546);
nor U702 (N_702,In_2434,In_2429);
nand U703 (N_703,In_2245,In_1491);
and U704 (N_704,In_115,In_23);
nor U705 (N_705,In_2301,In_683);
nor U706 (N_706,In_412,In_97);
nor U707 (N_707,In_1137,In_883);
and U708 (N_708,In_2080,In_715);
or U709 (N_709,In_427,In_1708);
or U710 (N_710,In_908,In_532);
nor U711 (N_711,In_2775,In_1663);
nand U712 (N_712,In_796,In_2275);
nand U713 (N_713,In_2704,In_741);
and U714 (N_714,In_275,In_37);
and U715 (N_715,In_2969,In_2362);
and U716 (N_716,In_91,In_861);
nand U717 (N_717,In_879,In_304);
and U718 (N_718,In_2983,In_2285);
nor U719 (N_719,In_1473,In_2864);
nor U720 (N_720,In_1507,In_59);
nand U721 (N_721,In_1252,In_621);
or U722 (N_722,In_2740,In_309);
and U723 (N_723,In_1115,In_714);
or U724 (N_724,In_2070,In_2957);
and U725 (N_725,In_2196,In_1250);
and U726 (N_726,In_38,In_402);
or U727 (N_727,In_178,In_223);
nor U728 (N_728,In_1614,In_316);
and U729 (N_729,In_1164,In_357);
or U730 (N_730,In_174,In_702);
nand U731 (N_731,In_2630,In_42);
and U732 (N_732,In_892,In_1182);
nand U733 (N_733,In_1042,In_2815);
and U734 (N_734,In_397,In_1196);
and U735 (N_735,In_2052,In_517);
nand U736 (N_736,In_2516,In_1329);
nand U737 (N_737,In_695,In_986);
nand U738 (N_738,In_1577,In_1858);
nor U739 (N_739,In_2942,In_2546);
xor U740 (N_740,In_633,In_2856);
nand U741 (N_741,In_2609,In_941);
and U742 (N_742,In_220,In_1905);
and U743 (N_743,In_2361,In_299);
and U744 (N_744,In_2889,In_240);
nor U745 (N_745,In_81,In_1337);
and U746 (N_746,In_2355,In_548);
nand U747 (N_747,In_64,In_2793);
or U748 (N_748,In_1046,In_1433);
nand U749 (N_749,In_1099,In_366);
nand U750 (N_750,In_2717,In_2694);
nor U751 (N_751,In_1468,In_1352);
and U752 (N_752,In_1652,In_2344);
and U753 (N_753,In_550,In_375);
and U754 (N_754,In_490,In_603);
nor U755 (N_755,In_2572,In_2232);
and U756 (N_756,In_1343,In_2457);
nor U757 (N_757,In_842,In_1769);
or U758 (N_758,In_2354,In_574);
and U759 (N_759,In_1172,In_1616);
and U760 (N_760,In_288,In_529);
nand U761 (N_761,In_475,In_1766);
nor U762 (N_762,In_40,In_1579);
nor U763 (N_763,In_1159,In_1538);
nand U764 (N_764,In_369,In_2905);
nand U765 (N_765,In_836,In_1863);
and U766 (N_766,In_2819,In_2074);
or U767 (N_767,In_2425,In_1745);
and U768 (N_768,In_2569,In_1281);
nor U769 (N_769,In_783,In_711);
nor U770 (N_770,In_428,In_1302);
nand U771 (N_771,In_1472,In_1240);
or U772 (N_772,In_1811,In_1569);
and U773 (N_773,In_2278,In_557);
or U774 (N_774,In_569,In_2833);
or U775 (N_775,In_758,In_2769);
nor U776 (N_776,In_1453,In_2339);
or U777 (N_777,In_44,In_813);
nor U778 (N_778,In_996,In_2838);
or U779 (N_779,In_2887,In_2379);
and U780 (N_780,In_1307,In_141);
nand U781 (N_781,In_2413,In_2650);
and U782 (N_782,In_1248,In_1069);
nand U783 (N_783,In_698,In_1336);
or U784 (N_784,In_2136,In_2043);
or U785 (N_785,In_2283,In_1190);
nor U786 (N_786,In_2022,In_2585);
nor U787 (N_787,In_828,In_2072);
and U788 (N_788,In_1886,In_2058);
and U789 (N_789,In_1669,In_1824);
nand U790 (N_790,In_2500,In_2210);
nor U791 (N_791,In_1161,In_2116);
or U792 (N_792,In_2314,In_837);
nor U793 (N_793,In_925,In_1549);
or U794 (N_794,In_1044,In_188);
nand U795 (N_795,In_1970,In_2321);
or U796 (N_796,In_250,In_2032);
nand U797 (N_797,In_961,In_2007);
nand U798 (N_798,In_776,In_1314);
or U799 (N_799,In_98,In_317);
or U800 (N_800,In_2672,In_263);
or U801 (N_801,In_2396,In_1895);
and U802 (N_802,In_1130,In_767);
nor U803 (N_803,In_133,In_1554);
and U804 (N_804,In_2033,In_1655);
or U805 (N_805,In_1634,In_520);
nand U806 (N_806,In_2758,In_1031);
nand U807 (N_807,In_1447,In_888);
nor U808 (N_808,In_1743,In_2606);
nand U809 (N_809,In_2157,In_2050);
and U810 (N_810,In_2986,In_601);
nor U811 (N_811,In_511,In_1179);
and U812 (N_812,In_862,In_106);
nor U813 (N_813,In_2549,In_2555);
or U814 (N_814,In_2206,In_1375);
nand U815 (N_815,In_237,In_2773);
and U816 (N_816,In_1353,In_2688);
nor U817 (N_817,In_2734,In_857);
and U818 (N_818,In_748,In_1681);
nor U819 (N_819,In_2133,In_990);
and U820 (N_820,In_2040,In_2945);
and U821 (N_821,In_630,In_1890);
xnor U822 (N_822,In_1110,In_658);
nor U823 (N_823,In_1927,In_1587);
nand U824 (N_824,In_2556,In_9);
and U825 (N_825,In_999,In_2006);
or U826 (N_826,In_274,In_1511);
and U827 (N_827,In_1424,In_1600);
nand U828 (N_828,In_962,In_1765);
nor U829 (N_829,In_2732,In_2470);
or U830 (N_830,In_980,In_2181);
nand U831 (N_831,In_1914,In_2252);
and U832 (N_832,In_1095,In_2994);
and U833 (N_833,In_938,In_112);
nand U834 (N_834,In_2227,In_1629);
and U835 (N_835,In_701,In_1260);
nand U836 (N_836,In_720,In_1465);
nand U837 (N_837,In_1651,In_2356);
nor U838 (N_838,In_2142,In_1221);
nor U839 (N_839,In_343,In_2854);
nor U840 (N_840,In_1070,In_2208);
nor U841 (N_841,In_969,In_474);
nor U842 (N_842,In_1867,In_1692);
or U843 (N_843,In_1394,In_334);
or U844 (N_844,In_1047,In_1864);
nand U845 (N_845,In_872,In_1261);
and U846 (N_846,In_1006,In_738);
or U847 (N_847,In_1427,In_1807);
nor U848 (N_848,In_1964,In_791);
nor U849 (N_849,In_2852,In_2480);
nor U850 (N_850,In_110,In_489);
or U851 (N_851,In_2184,In_2230);
or U852 (N_852,In_2105,In_462);
and U853 (N_853,In_1812,In_676);
nor U854 (N_854,In_1721,In_659);
nor U855 (N_855,In_406,In_722);
or U856 (N_856,In_2417,In_1732);
and U857 (N_857,In_1418,In_411);
nand U858 (N_858,In_1649,In_2845);
nor U859 (N_859,In_194,In_1476);
and U860 (N_860,In_1034,In_1271);
or U861 (N_861,In_589,In_949);
and U862 (N_862,In_1553,In_1222);
nand U863 (N_863,In_33,In_2762);
nor U864 (N_864,In_734,In_802);
or U865 (N_865,In_2304,In_484);
or U866 (N_866,In_1145,In_916);
or U867 (N_867,In_1313,In_1919);
and U868 (N_868,In_2622,In_387);
and U869 (N_869,In_2927,In_377);
and U870 (N_870,In_1781,In_430);
nor U871 (N_871,In_749,In_2333);
nor U872 (N_872,In_212,In_204);
and U873 (N_873,In_581,In_2145);
nor U874 (N_874,In_1499,In_2776);
and U875 (N_875,In_786,In_1075);
and U876 (N_876,In_2663,In_267);
or U877 (N_877,In_1930,In_2000);
or U878 (N_878,In_2866,In_2132);
and U879 (N_879,In_1706,In_2826);
nand U880 (N_880,In_2438,In_2377);
nor U881 (N_881,In_2547,In_847);
and U882 (N_882,In_2030,In_2771);
or U883 (N_883,In_2152,In_2385);
nand U884 (N_884,In_816,In_2395);
nand U885 (N_885,In_977,In_635);
nand U886 (N_886,In_442,In_1125);
or U887 (N_887,In_491,In_2126);
or U888 (N_888,In_1748,In_1310);
or U889 (N_889,In_2765,In_1296);
or U890 (N_890,In_1283,In_1774);
xnor U891 (N_891,In_454,In_1783);
and U892 (N_892,In_2096,In_810);
nor U893 (N_893,In_2423,In_1879);
or U894 (N_894,In_404,In_1001);
nand U895 (N_895,In_1177,In_1263);
nor U896 (N_896,In_1202,In_2106);
nand U897 (N_897,In_661,In_2271);
or U898 (N_898,In_2560,In_94);
nor U899 (N_899,In_124,In_896);
nand U900 (N_900,In_826,In_1326);
or U901 (N_901,In_1203,In_1526);
and U902 (N_902,In_2655,In_636);
or U903 (N_903,In_2871,In_2253);
or U904 (N_904,In_1189,In_271);
nor U905 (N_905,In_935,In_1324);
xnor U906 (N_906,In_2306,In_395);
and U907 (N_907,In_2221,In_168);
or U908 (N_908,In_355,In_1775);
nand U909 (N_909,In_1355,In_1086);
nor U910 (N_910,In_2764,In_926);
nand U911 (N_911,In_351,In_2337);
or U912 (N_912,In_1971,In_855);
and U913 (N_913,In_2745,In_617);
or U914 (N_914,In_2638,In_270);
and U915 (N_915,In_1618,In_1485);
and U916 (N_916,In_1312,In_50);
and U917 (N_917,In_646,In_649);
or U918 (N_918,In_259,In_803);
nor U919 (N_919,In_152,In_2902);
and U920 (N_920,In_524,In_988);
or U921 (N_921,In_2135,In_2005);
or U922 (N_922,In_2878,In_1180);
nor U923 (N_923,In_432,In_2633);
and U924 (N_924,In_760,In_913);
or U925 (N_925,In_1545,In_151);
or U926 (N_926,In_507,In_2950);
or U927 (N_927,In_1466,In_150);
or U928 (N_928,In_1193,In_272);
or U929 (N_929,In_371,In_2266);
or U930 (N_930,In_2670,In_1943);
nand U931 (N_931,In_1561,In_1386);
and U932 (N_932,In_1140,In_1384);
nor U933 (N_933,In_873,In_824);
nor U934 (N_934,In_435,In_2708);
nand U935 (N_935,In_32,In_2166);
and U936 (N_936,In_1682,In_1620);
nand U937 (N_937,In_2509,In_1977);
and U938 (N_938,In_889,In_2255);
and U939 (N_939,In_1237,In_503);
and U940 (N_940,In_1795,In_1841);
and U941 (N_941,In_2962,In_2553);
nor U942 (N_942,In_2308,In_1846);
and U943 (N_943,In_733,In_707);
nor U944 (N_944,In_931,In_510);
nand U945 (N_945,In_70,In_2948);
or U946 (N_946,In_1267,In_2397);
nor U947 (N_947,In_957,In_2151);
and U948 (N_948,In_1092,In_1530);
or U949 (N_949,In_2218,In_2718);
or U950 (N_950,In_2204,In_1258);
nor U951 (N_951,In_2,In_284);
nor U952 (N_952,In_1856,In_415);
and U953 (N_953,In_2567,In_2242);
nand U954 (N_954,In_67,In_2092);
or U955 (N_955,In_2019,In_1753);
and U956 (N_956,In_2789,In_2366);
nand U957 (N_957,In_1853,In_2691);
nor U958 (N_958,In_2191,In_1771);
and U959 (N_959,In_95,In_2239);
or U960 (N_960,In_712,In_11);
nor U961 (N_961,In_1607,In_1200);
nand U962 (N_962,In_1633,In_25);
nor U963 (N_963,In_1994,In_2309);
or U964 (N_964,In_450,In_1308);
nor U965 (N_965,In_2597,In_1183);
and U966 (N_966,In_1209,In_1403);
and U967 (N_967,In_1632,In_618);
nand U968 (N_968,In_2192,In_2988);
or U969 (N_969,In_921,In_1215);
or U970 (N_970,In_1912,In_433);
nand U971 (N_971,In_2076,In_641);
nor U972 (N_972,In_2656,In_1585);
nand U973 (N_973,In_2371,In_421);
nor U974 (N_974,In_531,In_2219);
nand U975 (N_975,In_1636,In_292);
nand U976 (N_976,In_2380,In_2405);
nand U977 (N_977,In_2543,In_1854);
and U978 (N_978,In_790,In_1504);
and U979 (N_979,In_1588,In_1236);
or U980 (N_980,In_759,In_1455);
or U981 (N_981,In_2097,In_2465);
nand U982 (N_982,In_662,In_1231);
and U983 (N_983,In_922,In_2736);
or U984 (N_984,In_2810,In_521);
and U985 (N_985,In_78,In_266);
nand U986 (N_986,In_1995,In_1825);
nand U987 (N_987,In_2566,In_2618);
nand U988 (N_988,In_1536,In_607);
or U989 (N_989,In_1494,In_2214);
nor U990 (N_990,In_1565,In_2761);
or U991 (N_991,In_2790,In_1060);
nor U992 (N_992,In_679,In_1544);
nor U993 (N_993,In_833,In_1622);
and U994 (N_994,In_2841,In_1788);
nor U995 (N_995,In_567,In_2875);
nand U996 (N_996,In_1480,In_1126);
nor U997 (N_997,In_201,In_905);
and U998 (N_998,In_156,In_190);
or U999 (N_999,In_2263,In_1409);
nand U1000 (N_1000,In_2502,In_2336);
nor U1001 (N_1001,In_261,In_403);
nand U1002 (N_1002,In_866,In_182);
or U1003 (N_1003,In_2424,In_1714);
and U1004 (N_1004,In_1689,In_2835);
nand U1005 (N_1005,In_2020,In_1915);
nand U1006 (N_1006,In_2258,In_2291);
nor U1007 (N_1007,In_2066,In_537);
nor U1008 (N_1008,In_2411,In_1635);
xor U1009 (N_1009,In_654,In_1972);
or U1010 (N_1010,In_213,In_2896);
nor U1011 (N_1011,In_2224,In_684);
or U1012 (N_1012,In_1963,In_1376);
nand U1013 (N_1013,In_1195,In_1685);
and U1014 (N_1014,In_256,In_47);
and U1015 (N_1015,In_512,In_2809);
nor U1016 (N_1016,In_445,In_1647);
nor U1017 (N_1017,In_85,In_2608);
and U1018 (N_1018,In_2588,In_2248);
nor U1019 (N_1019,In_540,In_1065);
nor U1020 (N_1020,In_1875,In_2573);
or U1021 (N_1021,In_2659,In_239);
nand U1022 (N_1022,In_673,In_2803);
or U1023 (N_1023,In_2709,In_342);
or U1024 (N_1024,In_1851,In_1799);
and U1025 (N_1025,In_2478,In_1961);
nor U1026 (N_1026,In_2055,In_1836);
nor U1027 (N_1027,In_2381,In_940);
or U1028 (N_1028,In_2746,In_2733);
or U1029 (N_1029,In_2605,In_2548);
or U1030 (N_1030,In_27,In_2406);
nor U1031 (N_1031,In_854,In_169);
or U1032 (N_1032,In_410,In_2017);
or U1033 (N_1033,In_1878,In_34);
nand U1034 (N_1034,In_260,In_1103);
nor U1035 (N_1035,In_825,In_2850);
and U1036 (N_1036,In_1100,In_1605);
nand U1037 (N_1037,In_1085,In_289);
or U1038 (N_1038,In_1820,In_2316);
nand U1039 (N_1039,In_345,In_2593);
nand U1040 (N_1040,In_2460,In_385);
and U1041 (N_1041,In_1639,In_587);
and U1042 (N_1042,In_2482,In_1211);
and U1043 (N_1043,In_2075,In_2753);
nand U1044 (N_1044,In_327,In_55);
nand U1045 (N_1045,In_2297,In_2676);
and U1046 (N_1046,In_2582,In_1175);
nor U1047 (N_1047,In_255,In_792);
or U1048 (N_1048,In_2855,In_1402);
nor U1049 (N_1049,In_1365,In_1157);
or U1050 (N_1050,In_1969,In_2091);
nor U1051 (N_1051,In_214,In_2167);
or U1052 (N_1052,In_99,In_2049);
or U1053 (N_1053,In_1429,In_691);
and U1054 (N_1054,In_553,In_2488);
and U1055 (N_1055,In_2954,In_2209);
and U1056 (N_1056,In_2402,In_2754);
and U1057 (N_1057,In_2607,In_2536);
or U1058 (N_1058,In_1881,In_651);
nor U1059 (N_1059,In_2886,In_1947);
nand U1060 (N_1060,In_2200,In_2225);
nand U1061 (N_1061,In_1865,In_645);
nor U1062 (N_1062,In_2277,In_1132);
nor U1063 (N_1063,In_1474,In_1582);
nand U1064 (N_1064,In_1780,In_1498);
or U1065 (N_1065,In_1997,In_924);
and U1066 (N_1066,In_21,In_1430);
or U1067 (N_1067,In_1239,In_2220);
and U1068 (N_1068,In_228,In_1699);
nand U1069 (N_1069,In_1356,In_2176);
or U1070 (N_1070,In_1362,In_2504);
nor U1071 (N_1071,In_470,In_1521);
xnor U1072 (N_1072,In_234,In_1922);
or U1073 (N_1073,In_1204,In_336);
nand U1074 (N_1074,In_1091,In_2272);
and U1075 (N_1075,In_1703,In_176);
or U1076 (N_1076,In_593,In_2596);
nand U1077 (N_1077,In_920,In_2849);
and U1078 (N_1078,In_1276,In_572);
or U1079 (N_1079,In_1003,In_2189);
and U1080 (N_1080,In_1575,In_2705);
nand U1081 (N_1081,In_1330,In_1951);
and U1082 (N_1082,In_933,In_1916);
nand U1083 (N_1083,In_2626,In_1735);
and U1084 (N_1084,In_1041,In_868);
nor U1085 (N_1085,In_1084,In_389);
or U1086 (N_1086,In_447,In_1462);
nor U1087 (N_1087,In_1319,In_1288);
xor U1088 (N_1088,In_2535,In_608);
nand U1089 (N_1089,In_2249,In_2448);
and U1090 (N_1090,In_283,In_1037);
nand U1091 (N_1091,In_1888,In_236);
or U1092 (N_1092,In_307,In_1413);
or U1093 (N_1093,In_1452,In_887);
nor U1094 (N_1094,In_2839,In_249);
and U1095 (N_1095,In_469,In_692);
or U1096 (N_1096,In_1345,In_2059);
and U1097 (N_1097,In_1434,In_1481);
and U1098 (N_1098,In_1648,In_2027);
nor U1099 (N_1099,In_1349,In_2037);
nand U1100 (N_1100,In_2583,In_3);
xor U1101 (N_1101,In_1548,In_2767);
nor U1102 (N_1102,In_444,In_1019);
and U1103 (N_1103,In_1050,In_1827);
nand U1104 (N_1104,In_1055,In_664);
or U1105 (N_1105,In_867,In_1397);
and U1106 (N_1106,In_1779,In_745);
nand U1107 (N_1107,In_2078,In_843);
nand U1108 (N_1108,In_2113,In_2563);
or U1109 (N_1109,In_2254,In_2246);
and U1110 (N_1110,In_329,In_18);
or U1111 (N_1111,In_1381,In_2960);
nand U1112 (N_1112,In_2197,In_2282);
nand U1113 (N_1113,In_217,In_984);
and U1114 (N_1114,In_1859,In_1908);
and U1115 (N_1115,In_254,In_668);
nor U1116 (N_1116,In_109,In_2898);
or U1117 (N_1117,In_2795,In_1233);
nand U1118 (N_1118,In_16,In_612);
and U1119 (N_1119,In_897,In_1642);
nand U1120 (N_1120,In_2876,In_361);
or U1121 (N_1121,In_1576,In_994);
or U1122 (N_1122,In_90,In_1883);
or U1123 (N_1123,In_198,In_2575);
and U1124 (N_1124,In_2897,In_1105);
and U1125 (N_1125,In_1589,In_372);
nor U1126 (N_1126,In_2320,In_2895);
or U1127 (N_1127,In_2821,In_2743);
or U1128 (N_1128,In_331,In_2953);
and U1129 (N_1129,In_1661,In_1848);
nor U1130 (N_1130,In_1123,In_148);
nand U1131 (N_1131,In_723,In_1079);
nor U1132 (N_1132,In_2807,In_1936);
nor U1133 (N_1133,In_966,In_312);
nand U1134 (N_1134,In_584,In_2155);
or U1135 (N_1135,In_779,In_1136);
nand U1136 (N_1136,In_2345,In_68);
nand U1137 (N_1137,In_60,In_2687);
nand U1138 (N_1138,In_2490,In_468);
or U1139 (N_1139,In_184,In_165);
nand U1140 (N_1140,In_1249,In_199);
or U1141 (N_1141,In_1035,In_205);
nand U1142 (N_1142,In_446,In_640);
or U1143 (N_1143,In_2163,In_2313);
nand U1144 (N_1144,In_1674,In_2047);
nor U1145 (N_1145,In_2101,In_1808);
and U1146 (N_1146,In_811,In_1790);
or U1147 (N_1147,In_533,In_2614);
nand U1148 (N_1148,In_1941,In_2669);
nor U1149 (N_1149,In_609,In_2391);
nor U1150 (N_1150,In_2668,In_643);
nor U1151 (N_1151,In_614,In_2923);
or U1152 (N_1152,In_499,In_1057);
xnor U1153 (N_1153,In_1869,In_1850);
or U1154 (N_1154,In_1335,In_56);
or U1155 (N_1155,In_744,In_1272);
or U1156 (N_1156,In_2760,In_1660);
and U1157 (N_1157,In_2274,In_1299);
and U1158 (N_1158,In_2158,In_628);
or U1159 (N_1159,In_2888,In_2035);
nor U1160 (N_1160,In_2939,In_789);
nand U1161 (N_1161,In_2947,In_1087);
nor U1162 (N_1162,In_2153,In_1750);
nor U1163 (N_1163,In_693,In_2018);
nor U1164 (N_1164,In_1469,In_2109);
nor U1165 (N_1165,In_2172,In_2735);
and U1166 (N_1166,In_2882,In_2435);
nor U1167 (N_1167,In_747,In_103);
nand U1168 (N_1168,In_936,In_2527);
nor U1169 (N_1169,In_1759,In_1486);
nor U1170 (N_1170,In_1834,In_1734);
and U1171 (N_1171,In_1855,In_2057);
or U1172 (N_1172,In_2298,In_438);
nor U1173 (N_1173,In_778,In_1686);
nand U1174 (N_1174,In_1138,In_704);
or U1175 (N_1175,In_1385,In_2777);
and U1176 (N_1176,In_1027,In_2273);
nand U1177 (N_1177,In_2851,In_2372);
and U1178 (N_1178,In_2823,In_777);
xnor U1179 (N_1179,In_2748,In_2713);
nor U1180 (N_1180,In_1129,In_561);
or U1181 (N_1181,In_2389,In_2427);
nand U1182 (N_1182,In_869,In_1143);
or U1183 (N_1183,In_2728,In_754);
or U1184 (N_1184,In_830,In_1831);
nor U1185 (N_1185,In_1493,In_1294);
and U1186 (N_1186,In_1744,In_2378);
or U1187 (N_1187,In_1220,In_689);
nor U1188 (N_1188,In_1986,In_1722);
nand U1189 (N_1189,In_2473,In_2182);
nand U1190 (N_1190,In_2415,In_1752);
or U1191 (N_1191,In_1664,In_1670);
nand U1192 (N_1192,In_2202,In_642);
nand U1193 (N_1193,In_2750,In_340);
nand U1194 (N_1194,In_2712,In_2973);
nor U1195 (N_1195,In_2603,In_2171);
or U1196 (N_1196,In_1608,In_1555);
nand U1197 (N_1197,In_2557,In_1893);
or U1198 (N_1198,In_632,In_1275);
or U1199 (N_1199,In_1528,In_15);
and U1200 (N_1200,In_1593,In_1704);
and U1201 (N_1201,In_1603,In_623);
nor U1202 (N_1202,In_2595,In_963);
and U1203 (N_1203,In_1265,In_230);
and U1204 (N_1204,In_1534,In_927);
nor U1205 (N_1205,In_1127,In_1583);
and U1206 (N_1206,In_1369,In_104);
or U1207 (N_1207,In_2508,In_2580);
and U1208 (N_1208,In_63,In_2721);
or U1209 (N_1209,In_287,In_2763);
or U1210 (N_1210,In_409,In_1899);
nor U1211 (N_1211,In_2716,In_785);
nor U1212 (N_1212,In_1698,In_556);
nor U1213 (N_1213,In_615,In_2180);
nor U1214 (N_1214,In_2587,In_571);
and U1215 (N_1215,In_875,In_1153);
and U1216 (N_1216,In_2404,In_416);
nor U1217 (N_1217,In_1184,In_460);
nor U1218 (N_1218,In_730,In_2008);
or U1219 (N_1219,In_149,In_2329);
nor U1220 (N_1220,In_2098,In_705);
nand U1221 (N_1221,In_471,In_2511);
nand U1222 (N_1222,In_1102,In_2825);
nor U1223 (N_1223,In_486,In_1573);
or U1224 (N_1224,In_675,In_2507);
and U1225 (N_1225,In_2514,In_1989);
nand U1226 (N_1226,In_1311,In_179);
nor U1227 (N_1227,In_2499,In_472);
and U1228 (N_1228,In_381,In_136);
nor U1229 (N_1229,In_1467,In_79);
nand U1230 (N_1230,In_2959,In_637);
nor U1231 (N_1231,In_2778,In_1580);
or U1232 (N_1232,In_2877,In_625);
and U1233 (N_1233,In_350,In_2813);
nand U1234 (N_1234,In_2662,In_1871);
or U1235 (N_1235,In_2122,In_2648);
nand U1236 (N_1236,In_1101,In_131);
nor U1237 (N_1237,In_227,In_2168);
and U1238 (N_1238,In_1974,In_185);
or U1239 (N_1239,In_2103,In_818);
and U1240 (N_1240,In_2044,In_2370);
nor U1241 (N_1241,In_719,In_2611);
nor U1242 (N_1242,In_2613,In_2088);
nand U1243 (N_1243,In_2665,In_1842);
or U1244 (N_1244,In_1729,In_1219);
nand U1245 (N_1245,In_325,In_2467);
or U1246 (N_1246,In_752,In_1198);
nor U1247 (N_1247,In_2322,In_1724);
nor U1248 (N_1248,In_1149,In_1395);
or U1249 (N_1249,In_799,In_1078);
nand U1250 (N_1250,In_502,In_971);
nand U1251 (N_1251,In_324,In_750);
nor U1252 (N_1252,In_2977,In_2358);
nor U1253 (N_1253,In_1551,In_1894);
or U1254 (N_1254,In_2492,In_476);
nor U1255 (N_1255,In_2491,In_330);
and U1256 (N_1256,In_1327,In_2014);
nand U1257 (N_1257,In_731,In_1431);
or U1258 (N_1258,In_2299,In_756);
and U1259 (N_1259,In_2039,In_2636);
and U1260 (N_1260,In_2211,In_2726);
or U1261 (N_1261,In_386,In_2203);
nor U1262 (N_1262,In_1815,In_477);
and U1263 (N_1263,In_2061,In_1158);
xor U1264 (N_1264,In_1278,In_1332);
or U1265 (N_1265,In_72,In_610);
and U1266 (N_1266,In_2820,In_1880);
and U1267 (N_1267,In_122,In_1067);
nor U1268 (N_1268,In_1793,In_19);
nor U1269 (N_1269,In_1539,In_2408);
or U1270 (N_1270,In_2458,In_2352);
and U1271 (N_1271,In_155,In_534);
or U1272 (N_1272,In_565,In_586);
or U1273 (N_1273,In_251,In_955);
nand U1274 (N_1274,In_2981,In_2824);
and U1275 (N_1275,In_2104,In_2664);
and U1276 (N_1276,In_362,In_5);
and U1277 (N_1277,In_431,In_2419);
or U1278 (N_1278,In_2545,In_814);
nor U1279 (N_1279,In_2652,In_1767);
nand U1280 (N_1280,In_706,In_388);
nor U1281 (N_1281,In_763,In_453);
nor U1282 (N_1282,In_2198,In_2418);
nor U1283 (N_1283,In_1784,In_54);
nand U1284 (N_1284,In_248,In_1695);
nand U1285 (N_1285,In_161,In_1071);
and U1286 (N_1286,In_1801,In_46);
nor U1287 (N_1287,In_1213,In_2107);
nand U1288 (N_1288,In_394,In_1301);
or U1289 (N_1289,In_2565,In_1098);
nor U1290 (N_1290,In_805,In_2483);
and U1291 (N_1291,In_1944,In_2349);
nor U1292 (N_1292,In_1645,In_1693);
nor U1293 (N_1293,In_1496,In_2533);
nand U1294 (N_1294,In_1658,In_1315);
and U1295 (N_1295,In_1514,In_2526);
nor U1296 (N_1296,In_885,In_2693);
and U1297 (N_1297,In_513,In_138);
and U1298 (N_1298,In_596,In_128);
nand U1299 (N_1299,In_1578,In_1876);
and U1300 (N_1300,In_2215,In_592);
nor U1301 (N_1301,In_378,In_832);
nand U1302 (N_1302,In_2695,In_605);
and U1303 (N_1303,In_958,In_1797);
and U1304 (N_1304,In_2779,In_2110);
and U1305 (N_1305,In_2318,In_547);
or U1306 (N_1306,In_681,In_2288);
or U1307 (N_1307,In_2085,In_1988);
nand U1308 (N_1308,In_154,In_2579);
and U1309 (N_1309,In_26,In_1937);
nor U1310 (N_1310,In_2087,In_1920);
and U1311 (N_1311,In_2004,In_877);
or U1312 (N_1312,In_1354,In_1347);
nand U1313 (N_1313,In_2677,In_2031);
nor U1314 (N_1314,In_1627,In_286);
or U1315 (N_1315,In_1776,In_2073);
nand U1316 (N_1316,In_993,In_2228);
and U1317 (N_1317,In_1460,In_985);
or U1318 (N_1318,In_2667,In_1216);
nor U1319 (N_1319,In_1798,In_1073);
and U1320 (N_1320,In_258,In_1303);
xor U1321 (N_1321,In_1952,In_1077);
or U1322 (N_1322,In_2046,In_2518);
nand U1323 (N_1323,In_1318,In_739);
nor U1324 (N_1324,In_302,In_2506);
and U1325 (N_1325,In_2908,In_2205);
or U1326 (N_1326,In_2590,In_1053);
nand U1327 (N_1327,In_2836,In_1710);
xnor U1328 (N_1328,In_2433,In_1074);
nor U1329 (N_1329,In_1738,In_1800);
xnor U1330 (N_1330,In_2173,In_1590);
nand U1331 (N_1331,In_2615,In_1033);
nor U1332 (N_1332,In_2454,In_354);
nand U1333 (N_1333,In_639,In_546);
and U1334 (N_1334,In_2065,In_2334);
or U1335 (N_1335,In_2534,In_296);
nand U1336 (N_1336,In_358,In_2520);
or U1337 (N_1337,In_1490,In_1736);
nand U1338 (N_1338,In_1640,In_1747);
xor U1339 (N_1339,In_2949,In_89);
or U1340 (N_1340,In_1306,In_884);
or U1341 (N_1341,In_1228,In_144);
or U1342 (N_1342,In_2637,In_934);
nand U1343 (N_1343,In_76,In_1226);
and U1344 (N_1344,In_2024,In_724);
nand U1345 (N_1345,In_2989,In_175);
nor U1346 (N_1346,In_2857,In_910);
nand U1347 (N_1347,In_2456,In_1350);
and U1348 (N_1348,In_2170,In_1749);
and U1349 (N_1349,In_1902,In_853);
nor U1350 (N_1350,In_1976,In_2161);
nor U1351 (N_1351,In_815,In_2312);
nor U1352 (N_1352,In_2100,In_1333);
or U1353 (N_1353,In_2229,In_206);
nor U1354 (N_1354,In_2416,In_1844);
nor U1355 (N_1355,In_84,In_1715);
nand U1356 (N_1356,In_2922,In_1758);
nand U1357 (N_1357,In_344,In_123);
nor U1358 (N_1358,In_145,In_2657);
or U1359 (N_1359,In_301,In_2279);
nand U1360 (N_1360,In_2373,In_1401);
nand U1361 (N_1361,In_907,In_1923);
nand U1362 (N_1362,In_1062,In_2294);
or U1363 (N_1363,In_2455,In_1529);
nor U1364 (N_1364,In_943,In_2574);
and U1365 (N_1365,In_88,In_1420);
xor U1366 (N_1366,In_2968,In_1891);
nor U1367 (N_1367,In_2749,In_1139);
or U1368 (N_1368,In_2235,In_1610);
nand U1369 (N_1369,In_2240,In_1796);
nor U1370 (N_1370,In_829,In_959);
and U1371 (N_1371,In_2187,In_1604);
nand U1372 (N_1372,In_117,In_480);
nor U1373 (N_1373,In_657,In_1707);
nor U1374 (N_1374,In_2350,In_2634);
nor U1375 (N_1375,In_903,In_140);
nor U1376 (N_1376,In_844,In_2800);
nand U1377 (N_1377,In_2510,In_1818);
and U1378 (N_1378,In_717,In_31);
nor U1379 (N_1379,In_2290,In_413);
and U1380 (N_1380,In_2741,In_2738);
nand U1381 (N_1381,In_2023,In_1830);
and U1382 (N_1382,In_1557,In_1166);
or U1383 (N_1383,In_285,In_2462);
and U1384 (N_1384,In_399,In_2384);
nand U1385 (N_1385,In_2045,In_86);
or U1386 (N_1386,In_2286,In_2869);
or U1387 (N_1387,In_992,In_2941);
nor U1388 (N_1388,In_1727,In_105);
or U1389 (N_1389,In_2021,In_2009);
and U1390 (N_1390,In_1877,In_1025);
nand U1391 (N_1391,In_568,In_265);
nand U1392 (N_1392,In_797,In_2244);
and U1393 (N_1393,In_678,In_243);
or U1394 (N_1394,In_697,In_1292);
nand U1395 (N_1395,In_2924,In_1690);
nand U1396 (N_1396,In_281,In_727);
nand U1397 (N_1397,In_965,In_2901);
nand U1398 (N_1398,In_335,In_2768);
or U1399 (N_1399,In_1761,In_1432);
and U1400 (N_1400,In_420,In_804);
nand U1401 (N_1401,In_1763,In_1023);
and U1402 (N_1402,In_429,In_2686);
nor U1403 (N_1403,In_793,In_1764);
and U1404 (N_1404,In_2944,In_2788);
nor U1405 (N_1405,In_2036,In_1574);
and U1406 (N_1406,In_1244,In_1543);
nor U1407 (N_1407,In_2893,In_798);
or U1408 (N_1408,In_216,In_726);
nor U1409 (N_1409,In_527,In_2148);
and U1410 (N_1410,In_368,In_1680);
nand U1411 (N_1411,In_2439,In_2451);
nand U1412 (N_1412,In_1806,In_2537);
and U1413 (N_1413,In_2409,In_2552);
nand U1414 (N_1414,In_392,In_374);
or U1415 (N_1415,In_1987,In_2260);
nor U1416 (N_1416,In_946,In_2787);
nand U1417 (N_1417,In_2956,In_997);
nor U1418 (N_1418,In_1286,In_1907);
or U1419 (N_1419,In_1671,In_2160);
and U1420 (N_1420,In_2797,In_2917);
nor U1421 (N_1421,In_1328,In_180);
or U1422 (N_1422,In_860,In_1407);
and U1423 (N_1423,In_2347,In_481);
nand U1424 (N_1424,In_2399,In_1805);
or U1425 (N_1425,In_1058,In_1245);
and U1426 (N_1426,In_303,In_1821);
and U1427 (N_1427,In_2584,In_746);
nor U1428 (N_1428,In_1483,In_1509);
nand U1429 (N_1429,In_2783,In_2620);
and U1430 (N_1430,In_2909,In_193);
or U1431 (N_1431,In_2437,In_1973);
nor U1432 (N_1432,In_1188,In_1992);
nand U1433 (N_1433,In_878,In_226);
or U1434 (N_1434,In_948,In_2410);
and U1435 (N_1435,In_439,In_2719);
or U1436 (N_1436,In_1586,In_1387);
or U1437 (N_1437,In_2929,In_2340);
or U1438 (N_1438,In_1083,In_1379);
nand U1439 (N_1439,In_1523,In_158);
and U1440 (N_1440,In_492,In_1665);
nand U1441 (N_1441,In_166,In_594);
and U1442 (N_1442,In_967,In_1106);
nor U1443 (N_1443,In_1408,In_1010);
nand U1444 (N_1444,In_171,In_1090);
nor U1445 (N_1445,In_1547,In_753);
or U1446 (N_1446,In_1346,In_2965);
or U1447 (N_1447,In_2680,In_1934);
nand U1448 (N_1448,In_2428,In_107);
nand U1449 (N_1449,In_552,In_647);
and U1450 (N_1450,In_1817,In_1208);
and U1451 (N_1451,In_2238,In_2971);
nor U1452 (N_1452,In_2442,In_982);
and U1453 (N_1453,In_886,In_2095);
xor U1454 (N_1454,In_1414,In_1014);
nor U1455 (N_1455,In_69,In_1440);
and U1456 (N_1456,In_1980,In_1368);
nand U1457 (N_1457,In_1688,In_365);
nand U1458 (N_1458,In_952,In_2703);
or U1459 (N_1459,In_2673,In_1456);
nand U1460 (N_1460,In_782,In_1373);
nor U1461 (N_1461,In_2199,In_2551);
nand U1462 (N_1462,In_215,In_159);
or U1463 (N_1463,In_2144,In_716);
nor U1464 (N_1464,In_2054,In_555);
or U1465 (N_1465,In_1955,In_515);
or U1466 (N_1466,In_2858,In_278);
and U1467 (N_1467,In_498,In_1998);
nor U1468 (N_1468,In_795,In_2134);
nor U1469 (N_1469,In_306,In_2177);
nor U1470 (N_1470,In_1253,In_2382);
nand U1471 (N_1471,In_162,In_436);
nor U1472 (N_1472,In_1733,In_2231);
nand U1473 (N_1473,In_2859,In_1676);
nand U1474 (N_1474,In_1619,In_12);
and U1475 (N_1475,In_1717,In_51);
nand U1476 (N_1476,In_1592,In_1567);
or U1477 (N_1477,In_1144,In_2816);
or U1478 (N_1478,In_1594,In_2757);
and U1479 (N_1479,In_2899,In_899);
or U1480 (N_1480,In_1280,In_2639);
nor U1481 (N_1481,In_2129,In_45);
nand U1482 (N_1482,In_1959,In_1170);
nor U1483 (N_1483,In_364,In_363);
nand U1484 (N_1484,In_2724,In_2991);
nand U1485 (N_1485,In_1730,In_942);
nor U1486 (N_1486,In_398,In_231);
and U1487 (N_1487,In_2690,In_2532);
and U1488 (N_1488,In_2625,In_221);
nor U1489 (N_1489,In_2125,In_2501);
and U1490 (N_1490,In_245,In_14);
and U1491 (N_1491,In_710,In_1996);
nor U1492 (N_1492,In_1040,In_1803);
nor U1493 (N_1493,In_1814,In_282);
nand U1494 (N_1494,In_822,In_2060);
and U1495 (N_1495,In_904,In_1946);
or U1496 (N_1496,In_1563,In_856);
or U1497 (N_1497,In_755,In_781);
nor U1498 (N_1498,In_743,In_1113);
nor U1499 (N_1499,In_1471,In_2094);
nand U1500 (N_1500,In_1010,In_1830);
nor U1501 (N_1501,In_890,In_250);
nand U1502 (N_1502,In_356,In_2724);
or U1503 (N_1503,In_424,In_2475);
nand U1504 (N_1504,In_2879,In_1615);
nand U1505 (N_1505,In_2603,In_655);
nand U1506 (N_1506,In_2848,In_886);
nor U1507 (N_1507,In_428,In_960);
or U1508 (N_1508,In_1206,In_1665);
nor U1509 (N_1509,In_2063,In_2315);
or U1510 (N_1510,In_2349,In_2823);
and U1511 (N_1511,In_1200,In_2816);
or U1512 (N_1512,In_2664,In_938);
or U1513 (N_1513,In_1584,In_2646);
and U1514 (N_1514,In_1385,In_305);
nand U1515 (N_1515,In_927,In_1841);
nor U1516 (N_1516,In_559,In_2191);
or U1517 (N_1517,In_2802,In_609);
nor U1518 (N_1518,In_2910,In_701);
nand U1519 (N_1519,In_298,In_96);
or U1520 (N_1520,In_2481,In_1219);
nand U1521 (N_1521,In_1334,In_2460);
or U1522 (N_1522,In_2566,In_659);
and U1523 (N_1523,In_921,In_2339);
nand U1524 (N_1524,In_1854,In_548);
nand U1525 (N_1525,In_2418,In_998);
nand U1526 (N_1526,In_849,In_2590);
nor U1527 (N_1527,In_190,In_628);
nand U1528 (N_1528,In_2150,In_2094);
nand U1529 (N_1529,In_347,In_829);
nand U1530 (N_1530,In_909,In_1501);
or U1531 (N_1531,In_1435,In_1689);
and U1532 (N_1532,In_554,In_908);
or U1533 (N_1533,In_1318,In_2454);
or U1534 (N_1534,In_2579,In_2211);
nand U1535 (N_1535,In_1444,In_2833);
nor U1536 (N_1536,In_1080,In_2467);
xor U1537 (N_1537,In_2121,In_2635);
or U1538 (N_1538,In_2624,In_227);
and U1539 (N_1539,In_1853,In_2291);
or U1540 (N_1540,In_2228,In_1554);
and U1541 (N_1541,In_2132,In_2584);
nor U1542 (N_1542,In_1094,In_1365);
nand U1543 (N_1543,In_342,In_2199);
and U1544 (N_1544,In_748,In_2880);
nand U1545 (N_1545,In_2830,In_1789);
or U1546 (N_1546,In_2393,In_2612);
or U1547 (N_1547,In_828,In_1835);
nand U1548 (N_1548,In_582,In_411);
and U1549 (N_1549,In_2159,In_879);
nor U1550 (N_1550,In_1598,In_787);
or U1551 (N_1551,In_1414,In_173);
and U1552 (N_1552,In_1150,In_2327);
nand U1553 (N_1553,In_775,In_1087);
nor U1554 (N_1554,In_2824,In_41);
and U1555 (N_1555,In_376,In_2499);
nor U1556 (N_1556,In_494,In_1571);
and U1557 (N_1557,In_2843,In_2820);
and U1558 (N_1558,In_777,In_1517);
or U1559 (N_1559,In_949,In_257);
xnor U1560 (N_1560,In_106,In_1154);
or U1561 (N_1561,In_1227,In_2385);
nor U1562 (N_1562,In_437,In_1370);
nand U1563 (N_1563,In_2187,In_2578);
nand U1564 (N_1564,In_2018,In_381);
and U1565 (N_1565,In_633,In_1433);
xor U1566 (N_1566,In_1491,In_977);
and U1567 (N_1567,In_1544,In_1848);
and U1568 (N_1568,In_2746,In_1946);
nand U1569 (N_1569,In_2175,In_736);
nand U1570 (N_1570,In_1274,In_1883);
nor U1571 (N_1571,In_1789,In_1518);
nand U1572 (N_1572,In_1989,In_2567);
nor U1573 (N_1573,In_2294,In_1418);
nand U1574 (N_1574,In_1724,In_1768);
nor U1575 (N_1575,In_949,In_1129);
and U1576 (N_1576,In_2651,In_840);
or U1577 (N_1577,In_858,In_432);
nor U1578 (N_1578,In_2062,In_2452);
nand U1579 (N_1579,In_356,In_837);
nand U1580 (N_1580,In_1866,In_1378);
and U1581 (N_1581,In_2859,In_1675);
nor U1582 (N_1582,In_562,In_1024);
or U1583 (N_1583,In_2716,In_788);
and U1584 (N_1584,In_2917,In_1689);
nand U1585 (N_1585,In_2440,In_953);
and U1586 (N_1586,In_1906,In_2393);
nand U1587 (N_1587,In_650,In_512);
nor U1588 (N_1588,In_79,In_1893);
or U1589 (N_1589,In_1667,In_1205);
nor U1590 (N_1590,In_642,In_980);
and U1591 (N_1591,In_2610,In_2149);
and U1592 (N_1592,In_674,In_1467);
or U1593 (N_1593,In_1269,In_2654);
nor U1594 (N_1594,In_603,In_621);
and U1595 (N_1595,In_510,In_2728);
nand U1596 (N_1596,In_1483,In_1801);
or U1597 (N_1597,In_711,In_1447);
and U1598 (N_1598,In_1537,In_2965);
nand U1599 (N_1599,In_2891,In_2353);
nand U1600 (N_1600,In_2728,In_243);
nand U1601 (N_1601,In_2051,In_1268);
nor U1602 (N_1602,In_1064,In_2267);
nor U1603 (N_1603,In_1129,In_2708);
nand U1604 (N_1604,In_2513,In_2867);
and U1605 (N_1605,In_1639,In_488);
nor U1606 (N_1606,In_564,In_819);
nand U1607 (N_1607,In_2783,In_89);
nor U1608 (N_1608,In_2408,In_1262);
nor U1609 (N_1609,In_2443,In_1734);
nand U1610 (N_1610,In_1644,In_959);
and U1611 (N_1611,In_1752,In_1172);
nor U1612 (N_1612,In_1678,In_499);
nand U1613 (N_1613,In_985,In_2747);
and U1614 (N_1614,In_2816,In_798);
nor U1615 (N_1615,In_2856,In_1227);
nor U1616 (N_1616,In_398,In_1912);
and U1617 (N_1617,In_2808,In_1833);
nor U1618 (N_1618,In_1213,In_2949);
and U1619 (N_1619,In_2822,In_1850);
nand U1620 (N_1620,In_166,In_1099);
nand U1621 (N_1621,In_760,In_1288);
and U1622 (N_1622,In_1733,In_2815);
nor U1623 (N_1623,In_2246,In_2859);
nand U1624 (N_1624,In_1013,In_43);
nor U1625 (N_1625,In_1208,In_783);
nand U1626 (N_1626,In_820,In_1039);
nand U1627 (N_1627,In_751,In_807);
nor U1628 (N_1628,In_2410,In_2414);
nand U1629 (N_1629,In_145,In_1177);
and U1630 (N_1630,In_152,In_1776);
and U1631 (N_1631,In_1166,In_2087);
or U1632 (N_1632,In_1016,In_2616);
or U1633 (N_1633,In_376,In_41);
nor U1634 (N_1634,In_499,In_2620);
and U1635 (N_1635,In_500,In_2241);
and U1636 (N_1636,In_2273,In_2603);
and U1637 (N_1637,In_986,In_2285);
nor U1638 (N_1638,In_768,In_2661);
nor U1639 (N_1639,In_1224,In_1588);
and U1640 (N_1640,In_1266,In_683);
or U1641 (N_1641,In_2161,In_1043);
nand U1642 (N_1642,In_1602,In_243);
or U1643 (N_1643,In_216,In_2518);
or U1644 (N_1644,In_2404,In_820);
xnor U1645 (N_1645,In_2139,In_2198);
and U1646 (N_1646,In_1928,In_599);
nor U1647 (N_1647,In_496,In_205);
nor U1648 (N_1648,In_1674,In_517);
nand U1649 (N_1649,In_2282,In_81);
or U1650 (N_1650,In_1415,In_1614);
nor U1651 (N_1651,In_844,In_329);
and U1652 (N_1652,In_14,In_284);
nor U1653 (N_1653,In_211,In_2873);
or U1654 (N_1654,In_557,In_689);
or U1655 (N_1655,In_356,In_1724);
nor U1656 (N_1656,In_1159,In_2869);
xor U1657 (N_1657,In_2583,In_1951);
nand U1658 (N_1658,In_606,In_1738);
and U1659 (N_1659,In_10,In_1769);
and U1660 (N_1660,In_2687,In_1947);
and U1661 (N_1661,In_911,In_2973);
or U1662 (N_1662,In_1936,In_2197);
nand U1663 (N_1663,In_501,In_686);
or U1664 (N_1664,In_1260,In_780);
or U1665 (N_1665,In_2407,In_1682);
nor U1666 (N_1666,In_2619,In_1334);
nand U1667 (N_1667,In_2755,In_1514);
nand U1668 (N_1668,In_455,In_2012);
and U1669 (N_1669,In_1351,In_276);
and U1670 (N_1670,In_1147,In_1734);
nand U1671 (N_1671,In_1119,In_2104);
and U1672 (N_1672,In_1102,In_2839);
and U1673 (N_1673,In_639,In_1436);
nand U1674 (N_1674,In_2255,In_1463);
or U1675 (N_1675,In_1680,In_1070);
and U1676 (N_1676,In_2847,In_1156);
and U1677 (N_1677,In_324,In_2986);
and U1678 (N_1678,In_720,In_1595);
nand U1679 (N_1679,In_2457,In_1316);
nand U1680 (N_1680,In_1060,In_2022);
nor U1681 (N_1681,In_250,In_2280);
and U1682 (N_1682,In_2062,In_318);
nor U1683 (N_1683,In_2081,In_1928);
and U1684 (N_1684,In_1736,In_2040);
nand U1685 (N_1685,In_2976,In_1778);
and U1686 (N_1686,In_2447,In_2884);
nor U1687 (N_1687,In_2295,In_2014);
or U1688 (N_1688,In_198,In_2617);
and U1689 (N_1689,In_1127,In_1206);
and U1690 (N_1690,In_1438,In_1279);
nand U1691 (N_1691,In_2522,In_1743);
nand U1692 (N_1692,In_875,In_223);
or U1693 (N_1693,In_2526,In_1925);
nand U1694 (N_1694,In_2660,In_1822);
or U1695 (N_1695,In_2476,In_155);
nand U1696 (N_1696,In_1866,In_2456);
or U1697 (N_1697,In_1782,In_2294);
xnor U1698 (N_1698,In_7,In_2185);
nand U1699 (N_1699,In_89,In_2206);
nor U1700 (N_1700,In_118,In_475);
nand U1701 (N_1701,In_1370,In_1545);
nor U1702 (N_1702,In_24,In_2746);
nand U1703 (N_1703,In_2413,In_1310);
nor U1704 (N_1704,In_30,In_1928);
nor U1705 (N_1705,In_1551,In_960);
nor U1706 (N_1706,In_2098,In_698);
nor U1707 (N_1707,In_258,In_1655);
or U1708 (N_1708,In_2702,In_1848);
nand U1709 (N_1709,In_1362,In_2587);
nor U1710 (N_1710,In_218,In_1514);
nor U1711 (N_1711,In_384,In_2797);
nor U1712 (N_1712,In_2817,In_2233);
nand U1713 (N_1713,In_1761,In_2832);
and U1714 (N_1714,In_2951,In_1029);
nand U1715 (N_1715,In_61,In_377);
and U1716 (N_1716,In_2584,In_2761);
xnor U1717 (N_1717,In_685,In_1541);
and U1718 (N_1718,In_1864,In_435);
nand U1719 (N_1719,In_684,In_2182);
or U1720 (N_1720,In_1977,In_1620);
nand U1721 (N_1721,In_2495,In_1209);
nand U1722 (N_1722,In_2203,In_2003);
nand U1723 (N_1723,In_446,In_2208);
nand U1724 (N_1724,In_328,In_1205);
nor U1725 (N_1725,In_2274,In_312);
nor U1726 (N_1726,In_1133,In_1239);
and U1727 (N_1727,In_282,In_84);
and U1728 (N_1728,In_573,In_1949);
or U1729 (N_1729,In_1911,In_2023);
nor U1730 (N_1730,In_106,In_1342);
and U1731 (N_1731,In_28,In_2510);
nand U1732 (N_1732,In_2226,In_2219);
and U1733 (N_1733,In_2355,In_114);
or U1734 (N_1734,In_1888,In_123);
or U1735 (N_1735,In_2923,In_1299);
nor U1736 (N_1736,In_929,In_1529);
nand U1737 (N_1737,In_1222,In_708);
nor U1738 (N_1738,In_2178,In_2378);
nand U1739 (N_1739,In_446,In_2709);
nor U1740 (N_1740,In_1152,In_2926);
and U1741 (N_1741,In_1037,In_205);
or U1742 (N_1742,In_2135,In_1578);
or U1743 (N_1743,In_2417,In_58);
or U1744 (N_1744,In_2968,In_2148);
or U1745 (N_1745,In_1383,In_1148);
nand U1746 (N_1746,In_1759,In_1872);
or U1747 (N_1747,In_310,In_2792);
nor U1748 (N_1748,In_589,In_1363);
nand U1749 (N_1749,In_1456,In_1148);
nand U1750 (N_1750,In_18,In_634);
nand U1751 (N_1751,In_495,In_2070);
nand U1752 (N_1752,In_2343,In_579);
nor U1753 (N_1753,In_2229,In_1623);
or U1754 (N_1754,In_503,In_2301);
nor U1755 (N_1755,In_887,In_429);
nand U1756 (N_1756,In_1216,In_191);
and U1757 (N_1757,In_2429,In_412);
and U1758 (N_1758,In_2794,In_1800);
nand U1759 (N_1759,In_1410,In_1587);
nor U1760 (N_1760,In_1178,In_580);
and U1761 (N_1761,In_1278,In_1779);
or U1762 (N_1762,In_920,In_2038);
nand U1763 (N_1763,In_361,In_2183);
nor U1764 (N_1764,In_1480,In_933);
nand U1765 (N_1765,In_1760,In_2157);
or U1766 (N_1766,In_119,In_2016);
nor U1767 (N_1767,In_2675,In_1081);
nor U1768 (N_1768,In_929,In_969);
nand U1769 (N_1769,In_1345,In_114);
and U1770 (N_1770,In_123,In_1830);
nand U1771 (N_1771,In_1999,In_864);
nor U1772 (N_1772,In_249,In_2795);
nor U1773 (N_1773,In_882,In_2425);
nor U1774 (N_1774,In_1090,In_2887);
or U1775 (N_1775,In_213,In_1224);
or U1776 (N_1776,In_2130,In_1888);
nor U1777 (N_1777,In_1347,In_1629);
or U1778 (N_1778,In_2594,In_1735);
nor U1779 (N_1779,In_1513,In_957);
xnor U1780 (N_1780,In_1061,In_1476);
nor U1781 (N_1781,In_1867,In_191);
nor U1782 (N_1782,In_1532,In_2612);
or U1783 (N_1783,In_2424,In_787);
or U1784 (N_1784,In_1966,In_376);
or U1785 (N_1785,In_1683,In_555);
nor U1786 (N_1786,In_2781,In_2848);
or U1787 (N_1787,In_1611,In_199);
or U1788 (N_1788,In_1691,In_2769);
nand U1789 (N_1789,In_2111,In_2415);
and U1790 (N_1790,In_651,In_1879);
nor U1791 (N_1791,In_824,In_2218);
nor U1792 (N_1792,In_841,In_2261);
and U1793 (N_1793,In_1948,In_796);
or U1794 (N_1794,In_339,In_2810);
xnor U1795 (N_1795,In_2782,In_1193);
and U1796 (N_1796,In_1402,In_1425);
or U1797 (N_1797,In_152,In_2661);
and U1798 (N_1798,In_1632,In_2623);
nand U1799 (N_1799,In_1497,In_1028);
or U1800 (N_1800,In_2726,In_2435);
nand U1801 (N_1801,In_2014,In_2992);
or U1802 (N_1802,In_1083,In_1077);
or U1803 (N_1803,In_2584,In_1357);
or U1804 (N_1804,In_1176,In_2478);
or U1805 (N_1805,In_1136,In_1806);
xnor U1806 (N_1806,In_1076,In_1680);
or U1807 (N_1807,In_1828,In_2325);
and U1808 (N_1808,In_2822,In_471);
and U1809 (N_1809,In_1461,In_1227);
nand U1810 (N_1810,In_2836,In_2251);
and U1811 (N_1811,In_330,In_2810);
nand U1812 (N_1812,In_106,In_168);
nand U1813 (N_1813,In_1698,In_1012);
nand U1814 (N_1814,In_1821,In_808);
nor U1815 (N_1815,In_98,In_281);
and U1816 (N_1816,In_783,In_2648);
nor U1817 (N_1817,In_2779,In_888);
nor U1818 (N_1818,In_2459,In_2753);
nor U1819 (N_1819,In_785,In_1006);
nor U1820 (N_1820,In_859,In_1036);
or U1821 (N_1821,In_2371,In_1442);
nor U1822 (N_1822,In_1926,In_1384);
nor U1823 (N_1823,In_791,In_1769);
nor U1824 (N_1824,In_1748,In_2727);
nor U1825 (N_1825,In_867,In_1405);
and U1826 (N_1826,In_1196,In_2227);
nor U1827 (N_1827,In_862,In_833);
nor U1828 (N_1828,In_623,In_1924);
nand U1829 (N_1829,In_2424,In_2674);
nand U1830 (N_1830,In_2320,In_197);
and U1831 (N_1831,In_2846,In_1892);
and U1832 (N_1832,In_2842,In_742);
nor U1833 (N_1833,In_2338,In_347);
nor U1834 (N_1834,In_2484,In_936);
or U1835 (N_1835,In_98,In_2602);
or U1836 (N_1836,In_469,In_575);
or U1837 (N_1837,In_1801,In_1009);
and U1838 (N_1838,In_282,In_1046);
or U1839 (N_1839,In_392,In_676);
xor U1840 (N_1840,In_1729,In_199);
nor U1841 (N_1841,In_2794,In_368);
nor U1842 (N_1842,In_2172,In_372);
nor U1843 (N_1843,In_2071,In_2771);
or U1844 (N_1844,In_553,In_1898);
or U1845 (N_1845,In_2599,In_2777);
or U1846 (N_1846,In_537,In_2065);
and U1847 (N_1847,In_1157,In_32);
nand U1848 (N_1848,In_556,In_1347);
nor U1849 (N_1849,In_2407,In_309);
and U1850 (N_1850,In_2696,In_943);
and U1851 (N_1851,In_1579,In_2825);
and U1852 (N_1852,In_1335,In_2878);
or U1853 (N_1853,In_63,In_1038);
or U1854 (N_1854,In_1635,In_279);
nor U1855 (N_1855,In_2330,In_1341);
or U1856 (N_1856,In_728,In_995);
nor U1857 (N_1857,In_850,In_1851);
or U1858 (N_1858,In_2162,In_389);
nand U1859 (N_1859,In_525,In_2268);
and U1860 (N_1860,In_2668,In_2947);
nand U1861 (N_1861,In_1982,In_2156);
and U1862 (N_1862,In_2219,In_2586);
or U1863 (N_1863,In_1726,In_2823);
nor U1864 (N_1864,In_1374,In_2402);
nand U1865 (N_1865,In_838,In_1654);
and U1866 (N_1866,In_2398,In_2420);
or U1867 (N_1867,In_1667,In_2016);
and U1868 (N_1868,In_496,In_88);
and U1869 (N_1869,In_1948,In_2808);
nand U1870 (N_1870,In_835,In_1066);
nand U1871 (N_1871,In_1350,In_636);
or U1872 (N_1872,In_2023,In_700);
or U1873 (N_1873,In_332,In_1354);
nor U1874 (N_1874,In_1442,In_329);
nor U1875 (N_1875,In_80,In_510);
or U1876 (N_1876,In_613,In_2173);
or U1877 (N_1877,In_1891,In_515);
nand U1878 (N_1878,In_1972,In_210);
or U1879 (N_1879,In_1112,In_2776);
or U1880 (N_1880,In_2376,In_2178);
nor U1881 (N_1881,In_828,In_2690);
nor U1882 (N_1882,In_2946,In_1543);
nor U1883 (N_1883,In_1173,In_544);
nor U1884 (N_1884,In_758,In_1926);
or U1885 (N_1885,In_591,In_799);
or U1886 (N_1886,In_496,In_1582);
and U1887 (N_1887,In_2487,In_1184);
nor U1888 (N_1888,In_2553,In_510);
or U1889 (N_1889,In_1396,In_2199);
or U1890 (N_1890,In_592,In_2045);
or U1891 (N_1891,In_1038,In_364);
nor U1892 (N_1892,In_2645,In_2320);
and U1893 (N_1893,In_1258,In_1745);
nor U1894 (N_1894,In_2822,In_2197);
or U1895 (N_1895,In_2410,In_1097);
and U1896 (N_1896,In_718,In_1932);
nand U1897 (N_1897,In_281,In_295);
and U1898 (N_1898,In_1832,In_1434);
and U1899 (N_1899,In_2829,In_1389);
nand U1900 (N_1900,In_1809,In_492);
and U1901 (N_1901,In_509,In_2270);
or U1902 (N_1902,In_151,In_1194);
and U1903 (N_1903,In_727,In_81);
and U1904 (N_1904,In_2891,In_2662);
or U1905 (N_1905,In_2795,In_2102);
and U1906 (N_1906,In_989,In_1703);
nand U1907 (N_1907,In_1051,In_1472);
or U1908 (N_1908,In_1086,In_2610);
nor U1909 (N_1909,In_57,In_461);
nor U1910 (N_1910,In_1562,In_2101);
or U1911 (N_1911,In_2198,In_2526);
nor U1912 (N_1912,In_2771,In_2045);
or U1913 (N_1913,In_1982,In_1870);
nor U1914 (N_1914,In_2021,In_2323);
or U1915 (N_1915,In_2487,In_1346);
nor U1916 (N_1916,In_1463,In_6);
nor U1917 (N_1917,In_2307,In_1206);
and U1918 (N_1918,In_2381,In_2340);
and U1919 (N_1919,In_2840,In_2173);
nand U1920 (N_1920,In_1388,In_169);
or U1921 (N_1921,In_749,In_2366);
nand U1922 (N_1922,In_2340,In_1473);
or U1923 (N_1923,In_2231,In_9);
and U1924 (N_1924,In_84,In_2002);
nand U1925 (N_1925,In_1828,In_2581);
nor U1926 (N_1926,In_2201,In_1363);
or U1927 (N_1927,In_196,In_492);
nor U1928 (N_1928,In_98,In_1798);
nand U1929 (N_1929,In_933,In_70);
nor U1930 (N_1930,In_1782,In_149);
nand U1931 (N_1931,In_1553,In_796);
and U1932 (N_1932,In_2615,In_1485);
nand U1933 (N_1933,In_617,In_354);
and U1934 (N_1934,In_334,In_2812);
and U1935 (N_1935,In_407,In_1131);
nor U1936 (N_1936,In_137,In_2892);
or U1937 (N_1937,In_2842,In_2751);
nor U1938 (N_1938,In_2765,In_922);
or U1939 (N_1939,In_2162,In_446);
and U1940 (N_1940,In_580,In_2269);
nor U1941 (N_1941,In_343,In_2838);
nand U1942 (N_1942,In_771,In_351);
nor U1943 (N_1943,In_2745,In_2299);
nor U1944 (N_1944,In_2428,In_1162);
and U1945 (N_1945,In_743,In_1452);
nand U1946 (N_1946,In_2128,In_2662);
nand U1947 (N_1947,In_2985,In_2015);
nand U1948 (N_1948,In_1337,In_415);
or U1949 (N_1949,In_286,In_947);
nand U1950 (N_1950,In_2605,In_2452);
nor U1951 (N_1951,In_518,In_386);
and U1952 (N_1952,In_1945,In_1796);
nand U1953 (N_1953,In_1715,In_2736);
nor U1954 (N_1954,In_2722,In_1041);
or U1955 (N_1955,In_1465,In_1002);
nand U1956 (N_1956,In_162,In_1614);
nand U1957 (N_1957,In_981,In_393);
or U1958 (N_1958,In_2166,In_1734);
nand U1959 (N_1959,In_346,In_1285);
or U1960 (N_1960,In_667,In_382);
or U1961 (N_1961,In_1493,In_950);
nand U1962 (N_1962,In_2657,In_2165);
nor U1963 (N_1963,In_545,In_469);
nand U1964 (N_1964,In_1301,In_99);
and U1965 (N_1965,In_1623,In_2950);
nand U1966 (N_1966,In_2428,In_2276);
nor U1967 (N_1967,In_2196,In_2810);
nand U1968 (N_1968,In_2155,In_2508);
nor U1969 (N_1969,In_412,In_443);
and U1970 (N_1970,In_1686,In_529);
and U1971 (N_1971,In_2496,In_292);
and U1972 (N_1972,In_1558,In_409);
nor U1973 (N_1973,In_517,In_2044);
or U1974 (N_1974,In_1108,In_1470);
nor U1975 (N_1975,In_520,In_954);
nor U1976 (N_1976,In_1572,In_1101);
nand U1977 (N_1977,In_933,In_1100);
nor U1978 (N_1978,In_123,In_1678);
nor U1979 (N_1979,In_645,In_489);
nand U1980 (N_1980,In_13,In_1658);
and U1981 (N_1981,In_2003,In_486);
or U1982 (N_1982,In_530,In_1343);
nand U1983 (N_1983,In_368,In_2237);
and U1984 (N_1984,In_1985,In_2117);
nand U1985 (N_1985,In_2002,In_645);
or U1986 (N_1986,In_758,In_1428);
or U1987 (N_1987,In_1387,In_2508);
nand U1988 (N_1988,In_2320,In_943);
or U1989 (N_1989,In_618,In_120);
nand U1990 (N_1990,In_2478,In_154);
nand U1991 (N_1991,In_2465,In_660);
nor U1992 (N_1992,In_2310,In_2391);
nor U1993 (N_1993,In_2463,In_2921);
nor U1994 (N_1994,In_1874,In_8);
or U1995 (N_1995,In_46,In_2121);
nor U1996 (N_1996,In_459,In_2273);
nand U1997 (N_1997,In_70,In_732);
nor U1998 (N_1998,In_583,In_1686);
and U1999 (N_1999,In_2812,In_631);
and U2000 (N_2000,In_1012,In_1482);
and U2001 (N_2001,In_2480,In_979);
nor U2002 (N_2002,In_2688,In_2473);
nand U2003 (N_2003,In_1771,In_546);
nand U2004 (N_2004,In_304,In_1254);
nor U2005 (N_2005,In_1361,In_468);
or U2006 (N_2006,In_1711,In_1363);
nand U2007 (N_2007,In_1924,In_2593);
and U2008 (N_2008,In_2778,In_258);
nand U2009 (N_2009,In_2502,In_12);
nor U2010 (N_2010,In_1382,In_1584);
nor U2011 (N_2011,In_982,In_2728);
nor U2012 (N_2012,In_553,In_1055);
nand U2013 (N_2013,In_1678,In_1589);
nor U2014 (N_2014,In_2495,In_584);
nor U2015 (N_2015,In_1783,In_953);
nand U2016 (N_2016,In_76,In_421);
and U2017 (N_2017,In_1137,In_2261);
nand U2018 (N_2018,In_1928,In_1261);
or U2019 (N_2019,In_1360,In_2012);
nand U2020 (N_2020,In_2488,In_2815);
xnor U2021 (N_2021,In_159,In_114);
nand U2022 (N_2022,In_859,In_2633);
nor U2023 (N_2023,In_2786,In_479);
and U2024 (N_2024,In_2986,In_2135);
and U2025 (N_2025,In_64,In_1316);
or U2026 (N_2026,In_1215,In_363);
nor U2027 (N_2027,In_2347,In_1026);
or U2028 (N_2028,In_2604,In_1063);
and U2029 (N_2029,In_687,In_1300);
and U2030 (N_2030,In_994,In_557);
nor U2031 (N_2031,In_545,In_2386);
and U2032 (N_2032,In_1098,In_211);
or U2033 (N_2033,In_1472,In_66);
nor U2034 (N_2034,In_2773,In_969);
nand U2035 (N_2035,In_872,In_1987);
nor U2036 (N_2036,In_1760,In_2444);
nand U2037 (N_2037,In_2954,In_493);
nand U2038 (N_2038,In_243,In_453);
or U2039 (N_2039,In_78,In_1480);
and U2040 (N_2040,In_1874,In_2250);
nor U2041 (N_2041,In_467,In_2506);
or U2042 (N_2042,In_2958,In_455);
and U2043 (N_2043,In_2939,In_422);
nand U2044 (N_2044,In_548,In_1818);
nor U2045 (N_2045,In_2929,In_1304);
nand U2046 (N_2046,In_44,In_1516);
and U2047 (N_2047,In_965,In_2072);
nand U2048 (N_2048,In_983,In_1127);
nand U2049 (N_2049,In_2565,In_1455);
nand U2050 (N_2050,In_2730,In_2205);
and U2051 (N_2051,In_2375,In_2090);
nand U2052 (N_2052,In_343,In_745);
nand U2053 (N_2053,In_651,In_2653);
or U2054 (N_2054,In_2807,In_2309);
and U2055 (N_2055,In_1898,In_139);
nand U2056 (N_2056,In_164,In_1618);
nor U2057 (N_2057,In_1115,In_1941);
or U2058 (N_2058,In_1882,In_1436);
nor U2059 (N_2059,In_345,In_2703);
and U2060 (N_2060,In_2540,In_2883);
nor U2061 (N_2061,In_504,In_2260);
and U2062 (N_2062,In_791,In_2645);
or U2063 (N_2063,In_2134,In_1002);
or U2064 (N_2064,In_1378,In_1857);
and U2065 (N_2065,In_1311,In_1470);
nand U2066 (N_2066,In_1478,In_1329);
or U2067 (N_2067,In_1060,In_1061);
and U2068 (N_2068,In_775,In_1528);
and U2069 (N_2069,In_1001,In_1743);
nand U2070 (N_2070,In_2755,In_2474);
and U2071 (N_2071,In_356,In_2780);
and U2072 (N_2072,In_15,In_552);
and U2073 (N_2073,In_1221,In_2165);
xnor U2074 (N_2074,In_1557,In_1704);
or U2075 (N_2075,In_1157,In_2537);
nand U2076 (N_2076,In_406,In_402);
nand U2077 (N_2077,In_1215,In_2512);
nand U2078 (N_2078,In_1491,In_578);
and U2079 (N_2079,In_1014,In_345);
nor U2080 (N_2080,In_2286,In_2046);
nand U2081 (N_2081,In_496,In_76);
nand U2082 (N_2082,In_1463,In_1905);
nand U2083 (N_2083,In_208,In_1286);
and U2084 (N_2084,In_523,In_1206);
and U2085 (N_2085,In_1726,In_654);
and U2086 (N_2086,In_1209,In_2067);
nor U2087 (N_2087,In_456,In_2111);
or U2088 (N_2088,In_219,In_1585);
nand U2089 (N_2089,In_1521,In_458);
nand U2090 (N_2090,In_1418,In_2068);
nand U2091 (N_2091,In_1491,In_1673);
nor U2092 (N_2092,In_1825,In_1708);
nand U2093 (N_2093,In_1109,In_2081);
and U2094 (N_2094,In_847,In_1878);
nand U2095 (N_2095,In_851,In_2845);
and U2096 (N_2096,In_2348,In_2471);
or U2097 (N_2097,In_431,In_1254);
nor U2098 (N_2098,In_2283,In_1455);
nand U2099 (N_2099,In_2334,In_1164);
nand U2100 (N_2100,In_585,In_458);
and U2101 (N_2101,In_2729,In_1913);
and U2102 (N_2102,In_2484,In_1666);
and U2103 (N_2103,In_1400,In_2454);
or U2104 (N_2104,In_2510,In_1551);
nand U2105 (N_2105,In_2642,In_572);
and U2106 (N_2106,In_1683,In_2053);
nor U2107 (N_2107,In_1359,In_1367);
and U2108 (N_2108,In_1356,In_610);
or U2109 (N_2109,In_2898,In_1897);
nand U2110 (N_2110,In_278,In_616);
nor U2111 (N_2111,In_577,In_596);
and U2112 (N_2112,In_932,In_2549);
or U2113 (N_2113,In_1492,In_1137);
nor U2114 (N_2114,In_1300,In_1616);
nor U2115 (N_2115,In_1758,In_2082);
or U2116 (N_2116,In_2382,In_1572);
or U2117 (N_2117,In_2488,In_1663);
or U2118 (N_2118,In_1776,In_1495);
and U2119 (N_2119,In_2516,In_710);
nor U2120 (N_2120,In_881,In_2314);
nor U2121 (N_2121,In_1716,In_2267);
or U2122 (N_2122,In_1806,In_2794);
nand U2123 (N_2123,In_198,In_1400);
or U2124 (N_2124,In_2018,In_1676);
and U2125 (N_2125,In_546,In_2682);
nand U2126 (N_2126,In_2464,In_523);
or U2127 (N_2127,In_2745,In_1105);
nor U2128 (N_2128,In_2853,In_714);
nor U2129 (N_2129,In_1710,In_2838);
nor U2130 (N_2130,In_57,In_232);
and U2131 (N_2131,In_1454,In_176);
and U2132 (N_2132,In_2114,In_2212);
nor U2133 (N_2133,In_2091,In_2080);
and U2134 (N_2134,In_1259,In_2162);
nor U2135 (N_2135,In_2143,In_634);
and U2136 (N_2136,In_2344,In_2422);
nor U2137 (N_2137,In_541,In_1494);
or U2138 (N_2138,In_271,In_1933);
and U2139 (N_2139,In_498,In_1027);
or U2140 (N_2140,In_1159,In_284);
nand U2141 (N_2141,In_626,In_2156);
or U2142 (N_2142,In_1139,In_706);
nor U2143 (N_2143,In_2001,In_779);
nand U2144 (N_2144,In_335,In_1444);
nor U2145 (N_2145,In_1475,In_2291);
or U2146 (N_2146,In_850,In_1671);
nand U2147 (N_2147,In_638,In_2912);
nor U2148 (N_2148,In_176,In_1253);
or U2149 (N_2149,In_2787,In_2868);
nand U2150 (N_2150,In_2419,In_1983);
nor U2151 (N_2151,In_696,In_2662);
or U2152 (N_2152,In_1155,In_2683);
or U2153 (N_2153,In_162,In_270);
and U2154 (N_2154,In_418,In_1545);
nor U2155 (N_2155,In_459,In_1256);
nand U2156 (N_2156,In_1231,In_278);
nand U2157 (N_2157,In_2795,In_1395);
or U2158 (N_2158,In_2855,In_1816);
xor U2159 (N_2159,In_1489,In_195);
or U2160 (N_2160,In_1778,In_1384);
or U2161 (N_2161,In_437,In_1367);
or U2162 (N_2162,In_563,In_1899);
nor U2163 (N_2163,In_241,In_280);
or U2164 (N_2164,In_326,In_1868);
nor U2165 (N_2165,In_2945,In_1379);
xnor U2166 (N_2166,In_2876,In_46);
or U2167 (N_2167,In_2219,In_2718);
nor U2168 (N_2168,In_1700,In_2135);
nand U2169 (N_2169,In_2200,In_813);
or U2170 (N_2170,In_303,In_77);
xor U2171 (N_2171,In_2451,In_1999);
nand U2172 (N_2172,In_2937,In_2913);
nor U2173 (N_2173,In_320,In_1063);
or U2174 (N_2174,In_1667,In_2627);
nand U2175 (N_2175,In_1330,In_1253);
or U2176 (N_2176,In_2437,In_1810);
and U2177 (N_2177,In_2139,In_2541);
nand U2178 (N_2178,In_868,In_588);
nand U2179 (N_2179,In_1747,In_791);
and U2180 (N_2180,In_919,In_1710);
nor U2181 (N_2181,In_1465,In_2577);
nor U2182 (N_2182,In_2145,In_2273);
and U2183 (N_2183,In_2650,In_1348);
nand U2184 (N_2184,In_778,In_2646);
nand U2185 (N_2185,In_740,In_104);
nand U2186 (N_2186,In_1026,In_2382);
nand U2187 (N_2187,In_2560,In_322);
nand U2188 (N_2188,In_2027,In_2630);
and U2189 (N_2189,In_2561,In_406);
nand U2190 (N_2190,In_1738,In_1225);
xor U2191 (N_2191,In_2017,In_2213);
nand U2192 (N_2192,In_2141,In_1984);
nand U2193 (N_2193,In_160,In_365);
nand U2194 (N_2194,In_1983,In_2431);
xnor U2195 (N_2195,In_2985,In_1047);
and U2196 (N_2196,In_2827,In_2465);
or U2197 (N_2197,In_2905,In_1500);
or U2198 (N_2198,In_1741,In_2854);
and U2199 (N_2199,In_2649,In_1562);
nor U2200 (N_2200,In_816,In_457);
or U2201 (N_2201,In_2182,In_2996);
and U2202 (N_2202,In_1104,In_1868);
and U2203 (N_2203,In_344,In_1599);
nor U2204 (N_2204,In_1613,In_578);
nor U2205 (N_2205,In_2600,In_1406);
and U2206 (N_2206,In_804,In_584);
and U2207 (N_2207,In_989,In_741);
nor U2208 (N_2208,In_2674,In_1173);
nor U2209 (N_2209,In_2356,In_2702);
nand U2210 (N_2210,In_2610,In_2530);
nor U2211 (N_2211,In_895,In_1452);
or U2212 (N_2212,In_814,In_212);
nand U2213 (N_2213,In_405,In_2805);
nor U2214 (N_2214,In_2577,In_719);
or U2215 (N_2215,In_933,In_419);
and U2216 (N_2216,In_2889,In_1421);
and U2217 (N_2217,In_2597,In_2393);
nand U2218 (N_2218,In_128,In_2329);
or U2219 (N_2219,In_1523,In_888);
nor U2220 (N_2220,In_528,In_2434);
nor U2221 (N_2221,In_1437,In_2872);
nor U2222 (N_2222,In_2675,In_2810);
or U2223 (N_2223,In_1577,In_631);
or U2224 (N_2224,In_1994,In_2628);
or U2225 (N_2225,In_1423,In_2506);
nand U2226 (N_2226,In_1970,In_2936);
or U2227 (N_2227,In_989,In_340);
and U2228 (N_2228,In_2370,In_227);
nand U2229 (N_2229,In_2842,In_43);
nand U2230 (N_2230,In_699,In_2295);
nand U2231 (N_2231,In_2399,In_1015);
nand U2232 (N_2232,In_1605,In_2666);
and U2233 (N_2233,In_1745,In_228);
nand U2234 (N_2234,In_1299,In_2358);
nand U2235 (N_2235,In_2601,In_2205);
nand U2236 (N_2236,In_889,In_2119);
nor U2237 (N_2237,In_1006,In_2855);
nand U2238 (N_2238,In_236,In_2226);
nor U2239 (N_2239,In_2520,In_2106);
and U2240 (N_2240,In_645,In_1000);
or U2241 (N_2241,In_708,In_1358);
or U2242 (N_2242,In_1983,In_585);
and U2243 (N_2243,In_339,In_913);
or U2244 (N_2244,In_1829,In_2825);
and U2245 (N_2245,In_2949,In_975);
nor U2246 (N_2246,In_1464,In_976);
nand U2247 (N_2247,In_2132,In_2434);
nand U2248 (N_2248,In_1767,In_885);
nor U2249 (N_2249,In_1049,In_353);
nand U2250 (N_2250,In_591,In_1456);
nor U2251 (N_2251,In_1327,In_1366);
and U2252 (N_2252,In_2976,In_2769);
nand U2253 (N_2253,In_1353,In_1702);
or U2254 (N_2254,In_2185,In_2676);
or U2255 (N_2255,In_1979,In_110);
or U2256 (N_2256,In_2152,In_189);
nand U2257 (N_2257,In_68,In_1173);
nor U2258 (N_2258,In_2228,In_1210);
or U2259 (N_2259,In_2067,In_2488);
or U2260 (N_2260,In_1442,In_1843);
nand U2261 (N_2261,In_2061,In_173);
and U2262 (N_2262,In_2540,In_1274);
or U2263 (N_2263,In_1006,In_1766);
and U2264 (N_2264,In_1860,In_857);
nor U2265 (N_2265,In_2076,In_1312);
nor U2266 (N_2266,In_209,In_145);
or U2267 (N_2267,In_1921,In_1388);
or U2268 (N_2268,In_251,In_227);
or U2269 (N_2269,In_1218,In_832);
nor U2270 (N_2270,In_125,In_1287);
nand U2271 (N_2271,In_2046,In_2322);
nor U2272 (N_2272,In_1725,In_576);
xor U2273 (N_2273,In_1885,In_862);
and U2274 (N_2274,In_418,In_83);
or U2275 (N_2275,In_1763,In_1011);
or U2276 (N_2276,In_527,In_116);
nand U2277 (N_2277,In_177,In_623);
nand U2278 (N_2278,In_2753,In_2919);
nor U2279 (N_2279,In_624,In_2762);
and U2280 (N_2280,In_572,In_1848);
and U2281 (N_2281,In_476,In_1803);
xnor U2282 (N_2282,In_2454,In_1401);
and U2283 (N_2283,In_853,In_2013);
or U2284 (N_2284,In_2441,In_2406);
and U2285 (N_2285,In_67,In_1650);
and U2286 (N_2286,In_108,In_1679);
nand U2287 (N_2287,In_2219,In_2508);
or U2288 (N_2288,In_2827,In_1122);
or U2289 (N_2289,In_1153,In_1213);
nor U2290 (N_2290,In_1675,In_1518);
and U2291 (N_2291,In_2712,In_477);
or U2292 (N_2292,In_1049,In_2849);
or U2293 (N_2293,In_319,In_315);
xor U2294 (N_2294,In_1875,In_2303);
or U2295 (N_2295,In_273,In_933);
nand U2296 (N_2296,In_71,In_2194);
or U2297 (N_2297,In_2807,In_1850);
nor U2298 (N_2298,In_1405,In_2458);
or U2299 (N_2299,In_2351,In_1253);
and U2300 (N_2300,In_2052,In_2594);
nor U2301 (N_2301,In_81,In_398);
or U2302 (N_2302,In_2036,In_508);
nor U2303 (N_2303,In_2887,In_1634);
or U2304 (N_2304,In_2786,In_2926);
nand U2305 (N_2305,In_213,In_2030);
nor U2306 (N_2306,In_1694,In_2964);
nand U2307 (N_2307,In_1139,In_44);
and U2308 (N_2308,In_1644,In_884);
and U2309 (N_2309,In_1314,In_2644);
and U2310 (N_2310,In_1386,In_1382);
or U2311 (N_2311,In_629,In_2545);
and U2312 (N_2312,In_273,In_2620);
nand U2313 (N_2313,In_1561,In_837);
or U2314 (N_2314,In_1786,In_281);
and U2315 (N_2315,In_1135,In_2566);
nor U2316 (N_2316,In_1791,In_1700);
and U2317 (N_2317,In_1781,In_1113);
nor U2318 (N_2318,In_1045,In_2270);
and U2319 (N_2319,In_988,In_1961);
or U2320 (N_2320,In_2275,In_2249);
nand U2321 (N_2321,In_964,In_2290);
nand U2322 (N_2322,In_980,In_1936);
nand U2323 (N_2323,In_667,In_204);
or U2324 (N_2324,In_2227,In_1429);
nor U2325 (N_2325,In_587,In_2676);
nand U2326 (N_2326,In_2642,In_1002);
xor U2327 (N_2327,In_5,In_1033);
and U2328 (N_2328,In_356,In_673);
nor U2329 (N_2329,In_1291,In_2613);
or U2330 (N_2330,In_2574,In_330);
xor U2331 (N_2331,In_2179,In_2037);
nor U2332 (N_2332,In_2482,In_233);
and U2333 (N_2333,In_2773,In_260);
and U2334 (N_2334,In_207,In_1999);
and U2335 (N_2335,In_825,In_2662);
nor U2336 (N_2336,In_2659,In_1329);
or U2337 (N_2337,In_1161,In_2362);
nand U2338 (N_2338,In_1467,In_266);
or U2339 (N_2339,In_2436,In_1038);
nand U2340 (N_2340,In_310,In_984);
and U2341 (N_2341,In_70,In_41);
or U2342 (N_2342,In_2724,In_121);
nand U2343 (N_2343,In_1557,In_1326);
nand U2344 (N_2344,In_813,In_1663);
and U2345 (N_2345,In_2871,In_1144);
or U2346 (N_2346,In_1675,In_761);
nand U2347 (N_2347,In_2060,In_937);
nor U2348 (N_2348,In_1111,In_2092);
or U2349 (N_2349,In_2478,In_2390);
nand U2350 (N_2350,In_2715,In_1457);
nor U2351 (N_2351,In_1477,In_1953);
or U2352 (N_2352,In_1698,In_2837);
nor U2353 (N_2353,In_420,In_2184);
and U2354 (N_2354,In_1160,In_1841);
nand U2355 (N_2355,In_401,In_2197);
and U2356 (N_2356,In_620,In_2707);
and U2357 (N_2357,In_950,In_943);
nand U2358 (N_2358,In_2030,In_2275);
and U2359 (N_2359,In_2108,In_1942);
or U2360 (N_2360,In_1468,In_2684);
nand U2361 (N_2361,In_2565,In_2631);
and U2362 (N_2362,In_2660,In_1849);
xor U2363 (N_2363,In_994,In_2809);
nand U2364 (N_2364,In_1875,In_1865);
or U2365 (N_2365,In_482,In_1397);
or U2366 (N_2366,In_363,In_1081);
and U2367 (N_2367,In_560,In_2158);
nand U2368 (N_2368,In_361,In_885);
and U2369 (N_2369,In_1172,In_51);
nor U2370 (N_2370,In_1014,In_1310);
and U2371 (N_2371,In_2889,In_1686);
and U2372 (N_2372,In_1232,In_685);
nor U2373 (N_2373,In_2204,In_2643);
nor U2374 (N_2374,In_2952,In_2505);
nand U2375 (N_2375,In_540,In_2726);
nand U2376 (N_2376,In_99,In_1015);
nand U2377 (N_2377,In_1865,In_2752);
nand U2378 (N_2378,In_2339,In_1148);
or U2379 (N_2379,In_1680,In_989);
nor U2380 (N_2380,In_1999,In_1955);
or U2381 (N_2381,In_437,In_2061);
and U2382 (N_2382,In_2136,In_409);
and U2383 (N_2383,In_1103,In_1856);
nor U2384 (N_2384,In_2021,In_402);
nand U2385 (N_2385,In_309,In_920);
or U2386 (N_2386,In_835,In_2350);
nand U2387 (N_2387,In_2034,In_1133);
and U2388 (N_2388,In_2894,In_2608);
nand U2389 (N_2389,In_731,In_2545);
xor U2390 (N_2390,In_109,In_2788);
nor U2391 (N_2391,In_983,In_2681);
or U2392 (N_2392,In_1605,In_985);
nand U2393 (N_2393,In_59,In_2085);
nand U2394 (N_2394,In_2830,In_1354);
nand U2395 (N_2395,In_2733,In_2052);
nand U2396 (N_2396,In_1324,In_2504);
nand U2397 (N_2397,In_1428,In_856);
nand U2398 (N_2398,In_2822,In_668);
nand U2399 (N_2399,In_2406,In_2402);
or U2400 (N_2400,In_501,In_1269);
nor U2401 (N_2401,In_1476,In_2370);
and U2402 (N_2402,In_544,In_677);
and U2403 (N_2403,In_1981,In_2492);
nor U2404 (N_2404,In_2126,In_1057);
nand U2405 (N_2405,In_1514,In_2265);
and U2406 (N_2406,In_2955,In_1416);
nor U2407 (N_2407,In_2534,In_196);
or U2408 (N_2408,In_1150,In_2989);
nor U2409 (N_2409,In_1882,In_864);
or U2410 (N_2410,In_1257,In_2928);
nand U2411 (N_2411,In_2853,In_2804);
nor U2412 (N_2412,In_1793,In_2497);
and U2413 (N_2413,In_1583,In_1952);
or U2414 (N_2414,In_45,In_352);
and U2415 (N_2415,In_1591,In_1589);
or U2416 (N_2416,In_2949,In_289);
nand U2417 (N_2417,In_1581,In_1524);
nand U2418 (N_2418,In_2830,In_1991);
nand U2419 (N_2419,In_2542,In_2974);
nand U2420 (N_2420,In_49,In_181);
nor U2421 (N_2421,In_309,In_961);
or U2422 (N_2422,In_1777,In_1881);
or U2423 (N_2423,In_958,In_1668);
and U2424 (N_2424,In_360,In_1708);
nand U2425 (N_2425,In_1866,In_2173);
and U2426 (N_2426,In_784,In_690);
or U2427 (N_2427,In_2708,In_141);
and U2428 (N_2428,In_434,In_1730);
and U2429 (N_2429,In_1083,In_1151);
nand U2430 (N_2430,In_1192,In_806);
nor U2431 (N_2431,In_2818,In_2252);
or U2432 (N_2432,In_1686,In_918);
or U2433 (N_2433,In_2416,In_2745);
nor U2434 (N_2434,In_82,In_1437);
and U2435 (N_2435,In_1563,In_15);
or U2436 (N_2436,In_437,In_1705);
nand U2437 (N_2437,In_2776,In_1587);
and U2438 (N_2438,In_2616,In_2230);
nor U2439 (N_2439,In_2133,In_691);
nand U2440 (N_2440,In_1454,In_2283);
nand U2441 (N_2441,In_157,In_337);
nand U2442 (N_2442,In_1117,In_1891);
nor U2443 (N_2443,In_388,In_2178);
nor U2444 (N_2444,In_319,In_1218);
nor U2445 (N_2445,In_2528,In_1262);
or U2446 (N_2446,In_2597,In_1583);
nand U2447 (N_2447,In_902,In_1538);
or U2448 (N_2448,In_2162,In_2873);
nand U2449 (N_2449,In_2401,In_697);
or U2450 (N_2450,In_261,In_2251);
and U2451 (N_2451,In_2874,In_2319);
nand U2452 (N_2452,In_1830,In_1642);
and U2453 (N_2453,In_2642,In_1731);
nor U2454 (N_2454,In_2416,In_2614);
or U2455 (N_2455,In_1462,In_539);
nor U2456 (N_2456,In_1054,In_257);
nor U2457 (N_2457,In_1814,In_1209);
or U2458 (N_2458,In_732,In_918);
nand U2459 (N_2459,In_2526,In_2839);
or U2460 (N_2460,In_1879,In_1419);
nand U2461 (N_2461,In_1539,In_1956);
and U2462 (N_2462,In_2576,In_2428);
and U2463 (N_2463,In_707,In_1574);
nor U2464 (N_2464,In_1991,In_2082);
nand U2465 (N_2465,In_2900,In_2533);
nand U2466 (N_2466,In_2866,In_227);
or U2467 (N_2467,In_436,In_37);
or U2468 (N_2468,In_2950,In_676);
nor U2469 (N_2469,In_266,In_1265);
and U2470 (N_2470,In_2306,In_900);
nor U2471 (N_2471,In_2712,In_1617);
or U2472 (N_2472,In_1616,In_11);
nor U2473 (N_2473,In_1347,In_408);
nor U2474 (N_2474,In_1865,In_2894);
nor U2475 (N_2475,In_453,In_509);
or U2476 (N_2476,In_1945,In_582);
and U2477 (N_2477,In_2033,In_1560);
nand U2478 (N_2478,In_1215,In_1108);
nand U2479 (N_2479,In_2658,In_2909);
nand U2480 (N_2480,In_597,In_738);
xnor U2481 (N_2481,In_1000,In_710);
or U2482 (N_2482,In_178,In_2344);
and U2483 (N_2483,In_1735,In_2716);
nor U2484 (N_2484,In_2804,In_2065);
and U2485 (N_2485,In_1275,In_1788);
nor U2486 (N_2486,In_746,In_1069);
nor U2487 (N_2487,In_2556,In_1767);
nor U2488 (N_2488,In_1559,In_425);
nand U2489 (N_2489,In_1355,In_2667);
or U2490 (N_2490,In_788,In_1250);
and U2491 (N_2491,In_115,In_2271);
and U2492 (N_2492,In_1933,In_850);
or U2493 (N_2493,In_2203,In_699);
nand U2494 (N_2494,In_2630,In_1632);
nand U2495 (N_2495,In_2767,In_833);
nor U2496 (N_2496,In_709,In_309);
and U2497 (N_2497,In_975,In_674);
nand U2498 (N_2498,In_1394,In_2886);
nor U2499 (N_2499,In_1448,In_1293);
nand U2500 (N_2500,In_2090,In_1983);
nor U2501 (N_2501,In_2668,In_2885);
nand U2502 (N_2502,In_2126,In_1922);
and U2503 (N_2503,In_1531,In_2147);
nor U2504 (N_2504,In_433,In_1270);
and U2505 (N_2505,In_2151,In_156);
and U2506 (N_2506,In_1166,In_2696);
and U2507 (N_2507,In_509,In_1246);
or U2508 (N_2508,In_1102,In_1596);
and U2509 (N_2509,In_630,In_2988);
nor U2510 (N_2510,In_472,In_2563);
and U2511 (N_2511,In_1045,In_2191);
nor U2512 (N_2512,In_2699,In_2325);
and U2513 (N_2513,In_1257,In_665);
nand U2514 (N_2514,In_2006,In_717);
and U2515 (N_2515,In_1709,In_617);
nand U2516 (N_2516,In_1491,In_1012);
or U2517 (N_2517,In_681,In_1993);
nand U2518 (N_2518,In_1977,In_534);
nand U2519 (N_2519,In_871,In_877);
or U2520 (N_2520,In_2687,In_1905);
nor U2521 (N_2521,In_2951,In_2972);
nand U2522 (N_2522,In_2310,In_1951);
nand U2523 (N_2523,In_2621,In_1956);
nand U2524 (N_2524,In_2574,In_2179);
nor U2525 (N_2525,In_2281,In_366);
nor U2526 (N_2526,In_1105,In_1761);
or U2527 (N_2527,In_1271,In_1540);
and U2528 (N_2528,In_279,In_209);
nand U2529 (N_2529,In_354,In_208);
or U2530 (N_2530,In_1922,In_489);
or U2531 (N_2531,In_399,In_956);
nand U2532 (N_2532,In_1100,In_1052);
nor U2533 (N_2533,In_9,In_1437);
and U2534 (N_2534,In_1790,In_1039);
nor U2535 (N_2535,In_2798,In_1043);
and U2536 (N_2536,In_1964,In_1835);
nor U2537 (N_2537,In_2039,In_1948);
nor U2538 (N_2538,In_1503,In_2223);
nand U2539 (N_2539,In_2069,In_1698);
nand U2540 (N_2540,In_973,In_486);
nand U2541 (N_2541,In_1528,In_1218);
xnor U2542 (N_2542,In_2554,In_2142);
nand U2543 (N_2543,In_467,In_353);
and U2544 (N_2544,In_2732,In_2464);
nor U2545 (N_2545,In_1746,In_724);
xor U2546 (N_2546,In_2555,In_832);
or U2547 (N_2547,In_1754,In_1825);
and U2548 (N_2548,In_1752,In_1014);
or U2549 (N_2549,In_77,In_2110);
nor U2550 (N_2550,In_1033,In_346);
nor U2551 (N_2551,In_364,In_2030);
or U2552 (N_2552,In_2639,In_908);
or U2553 (N_2553,In_1993,In_1484);
xnor U2554 (N_2554,In_2991,In_153);
nand U2555 (N_2555,In_2545,In_1938);
nor U2556 (N_2556,In_1515,In_1254);
and U2557 (N_2557,In_454,In_438);
and U2558 (N_2558,In_2839,In_2841);
and U2559 (N_2559,In_2336,In_2061);
nand U2560 (N_2560,In_1645,In_1362);
or U2561 (N_2561,In_147,In_2253);
or U2562 (N_2562,In_2058,In_2574);
or U2563 (N_2563,In_549,In_2468);
or U2564 (N_2564,In_2103,In_2710);
or U2565 (N_2565,In_983,In_1208);
or U2566 (N_2566,In_701,In_2157);
and U2567 (N_2567,In_2983,In_2970);
nand U2568 (N_2568,In_686,In_1336);
and U2569 (N_2569,In_593,In_477);
nor U2570 (N_2570,In_2891,In_632);
nand U2571 (N_2571,In_56,In_671);
nor U2572 (N_2572,In_253,In_1762);
nand U2573 (N_2573,In_1900,In_1465);
nor U2574 (N_2574,In_527,In_230);
and U2575 (N_2575,In_118,In_2264);
or U2576 (N_2576,In_221,In_166);
nor U2577 (N_2577,In_549,In_1995);
nor U2578 (N_2578,In_2753,In_824);
or U2579 (N_2579,In_1898,In_570);
and U2580 (N_2580,In_2083,In_319);
and U2581 (N_2581,In_218,In_2112);
or U2582 (N_2582,In_1845,In_2070);
nand U2583 (N_2583,In_2337,In_1791);
nor U2584 (N_2584,In_1636,In_2044);
and U2585 (N_2585,In_1647,In_99);
nand U2586 (N_2586,In_2132,In_1970);
nand U2587 (N_2587,In_2906,In_1508);
and U2588 (N_2588,In_947,In_199);
and U2589 (N_2589,In_1171,In_2295);
nor U2590 (N_2590,In_147,In_1701);
nand U2591 (N_2591,In_2755,In_2206);
nand U2592 (N_2592,In_1357,In_406);
or U2593 (N_2593,In_1481,In_2337);
nand U2594 (N_2594,In_1649,In_1841);
or U2595 (N_2595,In_1361,In_436);
and U2596 (N_2596,In_288,In_396);
and U2597 (N_2597,In_1647,In_2999);
nor U2598 (N_2598,In_644,In_1947);
nand U2599 (N_2599,In_490,In_1430);
nand U2600 (N_2600,In_2419,In_2709);
or U2601 (N_2601,In_925,In_639);
nand U2602 (N_2602,In_1259,In_609);
nor U2603 (N_2603,In_787,In_1984);
nand U2604 (N_2604,In_2108,In_1401);
nand U2605 (N_2605,In_1581,In_959);
nand U2606 (N_2606,In_2907,In_1568);
and U2607 (N_2607,In_2550,In_2427);
or U2608 (N_2608,In_1379,In_1729);
or U2609 (N_2609,In_2069,In_2894);
nand U2610 (N_2610,In_2497,In_1299);
nor U2611 (N_2611,In_1735,In_364);
and U2612 (N_2612,In_2254,In_227);
nor U2613 (N_2613,In_5,In_44);
nor U2614 (N_2614,In_2768,In_2720);
and U2615 (N_2615,In_245,In_1183);
and U2616 (N_2616,In_2844,In_495);
nand U2617 (N_2617,In_2234,In_2073);
nand U2618 (N_2618,In_738,In_1310);
xor U2619 (N_2619,In_821,In_1602);
nand U2620 (N_2620,In_661,In_1120);
and U2621 (N_2621,In_2789,In_274);
nor U2622 (N_2622,In_1610,In_56);
nor U2623 (N_2623,In_687,In_242);
or U2624 (N_2624,In_2510,In_768);
or U2625 (N_2625,In_611,In_693);
nand U2626 (N_2626,In_1409,In_1347);
nor U2627 (N_2627,In_2343,In_1759);
nand U2628 (N_2628,In_1439,In_2447);
nor U2629 (N_2629,In_2323,In_2666);
nand U2630 (N_2630,In_1835,In_1541);
or U2631 (N_2631,In_2103,In_144);
nor U2632 (N_2632,In_2566,In_56);
nor U2633 (N_2633,In_1406,In_1820);
and U2634 (N_2634,In_992,In_1977);
or U2635 (N_2635,In_1654,In_546);
and U2636 (N_2636,In_2904,In_2775);
nor U2637 (N_2637,In_93,In_713);
or U2638 (N_2638,In_787,In_2020);
nor U2639 (N_2639,In_2014,In_1246);
or U2640 (N_2640,In_375,In_1332);
nor U2641 (N_2641,In_1928,In_1575);
and U2642 (N_2642,In_2143,In_2424);
nor U2643 (N_2643,In_1739,In_246);
nor U2644 (N_2644,In_2054,In_2308);
nand U2645 (N_2645,In_1989,In_1595);
nor U2646 (N_2646,In_1493,In_709);
nor U2647 (N_2647,In_2329,In_1782);
and U2648 (N_2648,In_1530,In_1891);
xor U2649 (N_2649,In_759,In_160);
and U2650 (N_2650,In_1571,In_2807);
nor U2651 (N_2651,In_2327,In_1306);
and U2652 (N_2652,In_2209,In_1067);
and U2653 (N_2653,In_966,In_790);
and U2654 (N_2654,In_1117,In_2435);
and U2655 (N_2655,In_173,In_2198);
and U2656 (N_2656,In_1369,In_2832);
nand U2657 (N_2657,In_2471,In_669);
nor U2658 (N_2658,In_1654,In_2640);
nand U2659 (N_2659,In_220,In_1823);
or U2660 (N_2660,In_49,In_400);
and U2661 (N_2661,In_641,In_671);
and U2662 (N_2662,In_2420,In_279);
nor U2663 (N_2663,In_1707,In_767);
nand U2664 (N_2664,In_243,In_2226);
and U2665 (N_2665,In_2729,In_478);
nand U2666 (N_2666,In_2817,In_1425);
nor U2667 (N_2667,In_2220,In_25);
and U2668 (N_2668,In_2805,In_2696);
nor U2669 (N_2669,In_684,In_1869);
nand U2670 (N_2670,In_1418,In_547);
nand U2671 (N_2671,In_629,In_2201);
and U2672 (N_2672,In_930,In_2402);
nand U2673 (N_2673,In_2085,In_692);
nor U2674 (N_2674,In_308,In_2151);
and U2675 (N_2675,In_2501,In_2662);
nand U2676 (N_2676,In_2627,In_2113);
nand U2677 (N_2677,In_1980,In_2552);
nand U2678 (N_2678,In_2270,In_2418);
nor U2679 (N_2679,In_2902,In_1814);
and U2680 (N_2680,In_2996,In_1459);
and U2681 (N_2681,In_1278,In_2643);
nor U2682 (N_2682,In_1950,In_1867);
nand U2683 (N_2683,In_451,In_2911);
or U2684 (N_2684,In_1153,In_2698);
nand U2685 (N_2685,In_2806,In_465);
nand U2686 (N_2686,In_2155,In_8);
nor U2687 (N_2687,In_1617,In_2864);
or U2688 (N_2688,In_1162,In_688);
or U2689 (N_2689,In_1164,In_2961);
nor U2690 (N_2690,In_1366,In_2531);
nand U2691 (N_2691,In_136,In_242);
and U2692 (N_2692,In_318,In_798);
nand U2693 (N_2693,In_1348,In_1660);
and U2694 (N_2694,In_2357,In_1296);
and U2695 (N_2695,In_1614,In_1900);
nand U2696 (N_2696,In_762,In_2610);
nand U2697 (N_2697,In_2125,In_943);
and U2698 (N_2698,In_2346,In_2861);
nor U2699 (N_2699,In_1711,In_2910);
nand U2700 (N_2700,In_2699,In_1990);
or U2701 (N_2701,In_576,In_2457);
or U2702 (N_2702,In_2526,In_1677);
xor U2703 (N_2703,In_1466,In_1074);
nor U2704 (N_2704,In_2651,In_512);
and U2705 (N_2705,In_823,In_598);
and U2706 (N_2706,In_2016,In_1642);
or U2707 (N_2707,In_2821,In_1415);
and U2708 (N_2708,In_2056,In_2267);
and U2709 (N_2709,In_2760,In_2623);
nor U2710 (N_2710,In_1110,In_1959);
nand U2711 (N_2711,In_421,In_1779);
nor U2712 (N_2712,In_1054,In_2546);
or U2713 (N_2713,In_1567,In_910);
or U2714 (N_2714,In_998,In_1523);
nand U2715 (N_2715,In_1719,In_1558);
or U2716 (N_2716,In_2064,In_1367);
or U2717 (N_2717,In_547,In_1758);
nand U2718 (N_2718,In_1483,In_2558);
nor U2719 (N_2719,In_1971,In_740);
or U2720 (N_2720,In_2582,In_357);
nand U2721 (N_2721,In_2607,In_1006);
nor U2722 (N_2722,In_1387,In_1710);
nor U2723 (N_2723,In_1829,In_2495);
and U2724 (N_2724,In_1062,In_549);
and U2725 (N_2725,In_1165,In_553);
and U2726 (N_2726,In_1851,In_2547);
and U2727 (N_2727,In_1972,In_389);
and U2728 (N_2728,In_2844,In_2749);
and U2729 (N_2729,In_2570,In_2347);
nand U2730 (N_2730,In_503,In_1369);
or U2731 (N_2731,In_751,In_1317);
and U2732 (N_2732,In_1269,In_1192);
and U2733 (N_2733,In_2348,In_1471);
nor U2734 (N_2734,In_2617,In_423);
nor U2735 (N_2735,In_2708,In_1135);
nor U2736 (N_2736,In_316,In_231);
or U2737 (N_2737,In_929,In_2454);
or U2738 (N_2738,In_1477,In_2366);
nor U2739 (N_2739,In_748,In_1740);
nand U2740 (N_2740,In_2341,In_200);
xor U2741 (N_2741,In_1878,In_2725);
nor U2742 (N_2742,In_786,In_284);
and U2743 (N_2743,In_2047,In_1993);
nand U2744 (N_2744,In_1191,In_195);
nor U2745 (N_2745,In_2820,In_1298);
and U2746 (N_2746,In_429,In_145);
nor U2747 (N_2747,In_1078,In_2238);
or U2748 (N_2748,In_2642,In_2117);
and U2749 (N_2749,In_2935,In_2744);
nand U2750 (N_2750,In_759,In_163);
and U2751 (N_2751,In_1557,In_151);
nor U2752 (N_2752,In_2604,In_2978);
and U2753 (N_2753,In_956,In_2677);
nor U2754 (N_2754,In_2200,In_2268);
or U2755 (N_2755,In_1124,In_60);
and U2756 (N_2756,In_2223,In_1556);
nor U2757 (N_2757,In_727,In_2676);
or U2758 (N_2758,In_155,In_2318);
and U2759 (N_2759,In_2583,In_1266);
or U2760 (N_2760,In_1014,In_1938);
nor U2761 (N_2761,In_1066,In_2665);
nand U2762 (N_2762,In_2519,In_2735);
and U2763 (N_2763,In_1283,In_2280);
nand U2764 (N_2764,In_1741,In_1665);
nand U2765 (N_2765,In_1795,In_598);
nand U2766 (N_2766,In_777,In_813);
or U2767 (N_2767,In_225,In_1227);
nor U2768 (N_2768,In_1338,In_994);
nor U2769 (N_2769,In_1298,In_1039);
or U2770 (N_2770,In_2832,In_961);
and U2771 (N_2771,In_1687,In_499);
nor U2772 (N_2772,In_2342,In_765);
or U2773 (N_2773,In_2609,In_2838);
and U2774 (N_2774,In_783,In_1148);
nor U2775 (N_2775,In_965,In_409);
or U2776 (N_2776,In_232,In_2600);
nand U2777 (N_2777,In_28,In_441);
and U2778 (N_2778,In_1069,In_2679);
xnor U2779 (N_2779,In_766,In_2605);
or U2780 (N_2780,In_685,In_1932);
nor U2781 (N_2781,In_2755,In_1653);
or U2782 (N_2782,In_2158,In_444);
nand U2783 (N_2783,In_838,In_1846);
nor U2784 (N_2784,In_1125,In_359);
nand U2785 (N_2785,In_1872,In_1399);
nor U2786 (N_2786,In_73,In_2667);
nor U2787 (N_2787,In_798,In_1073);
and U2788 (N_2788,In_2306,In_706);
and U2789 (N_2789,In_289,In_64);
nor U2790 (N_2790,In_2721,In_1867);
nand U2791 (N_2791,In_2020,In_2643);
and U2792 (N_2792,In_2031,In_2378);
and U2793 (N_2793,In_1912,In_1608);
or U2794 (N_2794,In_188,In_522);
and U2795 (N_2795,In_1056,In_534);
nor U2796 (N_2796,In_126,In_2938);
nand U2797 (N_2797,In_1135,In_1274);
or U2798 (N_2798,In_2086,In_1567);
or U2799 (N_2799,In_2516,In_308);
nand U2800 (N_2800,In_1424,In_1999);
nand U2801 (N_2801,In_2232,In_2203);
nor U2802 (N_2802,In_178,In_2380);
nand U2803 (N_2803,In_2950,In_2301);
nor U2804 (N_2804,In_2607,In_1835);
nand U2805 (N_2805,In_721,In_2383);
nor U2806 (N_2806,In_50,In_1952);
or U2807 (N_2807,In_2424,In_174);
nor U2808 (N_2808,In_1122,In_2779);
nor U2809 (N_2809,In_2536,In_2438);
and U2810 (N_2810,In_1455,In_1238);
nor U2811 (N_2811,In_2566,In_573);
or U2812 (N_2812,In_76,In_757);
nor U2813 (N_2813,In_2277,In_577);
nand U2814 (N_2814,In_1781,In_2956);
nand U2815 (N_2815,In_1944,In_867);
or U2816 (N_2816,In_2219,In_1974);
and U2817 (N_2817,In_2340,In_933);
nand U2818 (N_2818,In_1796,In_2468);
or U2819 (N_2819,In_2899,In_2890);
nand U2820 (N_2820,In_1683,In_2501);
nor U2821 (N_2821,In_556,In_461);
nand U2822 (N_2822,In_847,In_1671);
nand U2823 (N_2823,In_1756,In_2216);
and U2824 (N_2824,In_1370,In_478);
nand U2825 (N_2825,In_1066,In_876);
and U2826 (N_2826,In_1271,In_2009);
nor U2827 (N_2827,In_937,In_2531);
nor U2828 (N_2828,In_653,In_1916);
and U2829 (N_2829,In_1255,In_1706);
nor U2830 (N_2830,In_839,In_2644);
nor U2831 (N_2831,In_2118,In_1350);
and U2832 (N_2832,In_332,In_901);
and U2833 (N_2833,In_476,In_2526);
nor U2834 (N_2834,In_2750,In_2837);
and U2835 (N_2835,In_2693,In_1452);
and U2836 (N_2836,In_506,In_327);
nor U2837 (N_2837,In_731,In_2831);
and U2838 (N_2838,In_2754,In_1935);
and U2839 (N_2839,In_2249,In_750);
or U2840 (N_2840,In_1013,In_1138);
and U2841 (N_2841,In_997,In_371);
or U2842 (N_2842,In_1284,In_2993);
nor U2843 (N_2843,In_1105,In_758);
and U2844 (N_2844,In_2387,In_2515);
and U2845 (N_2845,In_2642,In_2617);
nand U2846 (N_2846,In_2315,In_1677);
nor U2847 (N_2847,In_2403,In_1720);
nor U2848 (N_2848,In_1358,In_1296);
nand U2849 (N_2849,In_55,In_891);
and U2850 (N_2850,In_1253,In_828);
or U2851 (N_2851,In_886,In_2784);
or U2852 (N_2852,In_1671,In_2800);
or U2853 (N_2853,In_2728,In_2582);
nand U2854 (N_2854,In_2960,In_109);
nand U2855 (N_2855,In_1056,In_583);
or U2856 (N_2856,In_2278,In_532);
nand U2857 (N_2857,In_515,In_1087);
or U2858 (N_2858,In_1201,In_1213);
and U2859 (N_2859,In_2523,In_2584);
or U2860 (N_2860,In_17,In_229);
nor U2861 (N_2861,In_169,In_1084);
nand U2862 (N_2862,In_592,In_271);
nor U2863 (N_2863,In_2082,In_908);
nor U2864 (N_2864,In_2592,In_1050);
or U2865 (N_2865,In_460,In_586);
nor U2866 (N_2866,In_1319,In_1555);
and U2867 (N_2867,In_2402,In_508);
nor U2868 (N_2868,In_228,In_417);
and U2869 (N_2869,In_1332,In_805);
nor U2870 (N_2870,In_2323,In_662);
and U2871 (N_2871,In_1887,In_2406);
nand U2872 (N_2872,In_1565,In_2177);
nand U2873 (N_2873,In_1623,In_2652);
nor U2874 (N_2874,In_1196,In_2596);
nor U2875 (N_2875,In_1421,In_1828);
nand U2876 (N_2876,In_1019,In_1011);
nand U2877 (N_2877,In_2775,In_1315);
xnor U2878 (N_2878,In_232,In_2798);
nor U2879 (N_2879,In_2607,In_1894);
nor U2880 (N_2880,In_332,In_2555);
and U2881 (N_2881,In_417,In_352);
and U2882 (N_2882,In_149,In_1236);
and U2883 (N_2883,In_1031,In_571);
or U2884 (N_2884,In_214,In_1275);
xor U2885 (N_2885,In_2977,In_2038);
nor U2886 (N_2886,In_1902,In_2876);
and U2887 (N_2887,In_1754,In_965);
and U2888 (N_2888,In_29,In_2560);
or U2889 (N_2889,In_1854,In_907);
or U2890 (N_2890,In_1809,In_239);
nor U2891 (N_2891,In_1970,In_2154);
nand U2892 (N_2892,In_1089,In_1942);
or U2893 (N_2893,In_1158,In_23);
nand U2894 (N_2894,In_2913,In_1533);
or U2895 (N_2895,In_1968,In_225);
xnor U2896 (N_2896,In_1062,In_1746);
or U2897 (N_2897,In_2033,In_2869);
xnor U2898 (N_2898,In_334,In_1438);
nand U2899 (N_2899,In_1869,In_1669);
nand U2900 (N_2900,In_995,In_1857);
nor U2901 (N_2901,In_1292,In_57);
nor U2902 (N_2902,In_16,In_2176);
nor U2903 (N_2903,In_372,In_1728);
and U2904 (N_2904,In_257,In_447);
and U2905 (N_2905,In_801,In_2440);
or U2906 (N_2906,In_2574,In_2951);
and U2907 (N_2907,In_1281,In_507);
nor U2908 (N_2908,In_1935,In_1389);
and U2909 (N_2909,In_2911,In_2008);
nor U2910 (N_2910,In_1133,In_916);
nand U2911 (N_2911,In_881,In_2735);
nand U2912 (N_2912,In_2641,In_161);
and U2913 (N_2913,In_1155,In_2310);
nand U2914 (N_2914,In_1799,In_2868);
or U2915 (N_2915,In_825,In_53);
and U2916 (N_2916,In_2172,In_706);
nor U2917 (N_2917,In_2922,In_2393);
or U2918 (N_2918,In_1064,In_1962);
nor U2919 (N_2919,In_2552,In_1003);
nand U2920 (N_2920,In_795,In_940);
nand U2921 (N_2921,In_638,In_2521);
and U2922 (N_2922,In_2133,In_1203);
and U2923 (N_2923,In_1940,In_1676);
and U2924 (N_2924,In_2222,In_189);
and U2925 (N_2925,In_2207,In_1413);
or U2926 (N_2926,In_265,In_1372);
nor U2927 (N_2927,In_2494,In_2599);
nor U2928 (N_2928,In_268,In_2400);
xor U2929 (N_2929,In_576,In_2742);
and U2930 (N_2930,In_2090,In_633);
or U2931 (N_2931,In_24,In_1945);
nand U2932 (N_2932,In_2874,In_1439);
nand U2933 (N_2933,In_2209,In_1987);
nand U2934 (N_2934,In_1305,In_2715);
nand U2935 (N_2935,In_398,In_2671);
nor U2936 (N_2936,In_1527,In_1432);
or U2937 (N_2937,In_2170,In_1861);
nor U2938 (N_2938,In_485,In_2781);
and U2939 (N_2939,In_1372,In_2432);
nand U2940 (N_2940,In_396,In_1309);
nand U2941 (N_2941,In_2583,In_2067);
and U2942 (N_2942,In_2695,In_2815);
or U2943 (N_2943,In_2024,In_1416);
nor U2944 (N_2944,In_788,In_342);
nor U2945 (N_2945,In_1020,In_2989);
and U2946 (N_2946,In_1503,In_2346);
and U2947 (N_2947,In_790,In_1507);
nor U2948 (N_2948,In_589,In_1212);
or U2949 (N_2949,In_1187,In_2127);
nand U2950 (N_2950,In_719,In_823);
nor U2951 (N_2951,In_1693,In_978);
nor U2952 (N_2952,In_2258,In_1040);
nor U2953 (N_2953,In_86,In_478);
nor U2954 (N_2954,In_562,In_325);
or U2955 (N_2955,In_264,In_2367);
nor U2956 (N_2956,In_1103,In_954);
nand U2957 (N_2957,In_2236,In_2048);
or U2958 (N_2958,In_1278,In_74);
nor U2959 (N_2959,In_1341,In_459);
nand U2960 (N_2960,In_1908,In_1347);
nor U2961 (N_2961,In_2741,In_2409);
nand U2962 (N_2962,In_1742,In_1330);
nand U2963 (N_2963,In_2716,In_2411);
or U2964 (N_2964,In_909,In_1482);
or U2965 (N_2965,In_2532,In_2698);
or U2966 (N_2966,In_420,In_1326);
nand U2967 (N_2967,In_638,In_373);
or U2968 (N_2968,In_2979,In_2347);
and U2969 (N_2969,In_2251,In_759);
nor U2970 (N_2970,In_2491,In_1863);
xor U2971 (N_2971,In_2367,In_2765);
nor U2972 (N_2972,In_1346,In_2686);
nor U2973 (N_2973,In_2465,In_1825);
or U2974 (N_2974,In_515,In_1111);
or U2975 (N_2975,In_2782,In_626);
or U2976 (N_2976,In_2199,In_397);
nand U2977 (N_2977,In_911,In_572);
or U2978 (N_2978,In_1566,In_2128);
or U2979 (N_2979,In_1602,In_1843);
and U2980 (N_2980,In_2912,In_878);
or U2981 (N_2981,In_2584,In_2156);
nand U2982 (N_2982,In_2310,In_25);
nor U2983 (N_2983,In_1001,In_2421);
and U2984 (N_2984,In_736,In_47);
or U2985 (N_2985,In_704,In_1928);
nor U2986 (N_2986,In_633,In_1870);
nor U2987 (N_2987,In_1279,In_847);
and U2988 (N_2988,In_2227,In_605);
and U2989 (N_2989,In_1906,In_1825);
nand U2990 (N_2990,In_693,In_538);
nor U2991 (N_2991,In_1426,In_2570);
or U2992 (N_2992,In_938,In_665);
or U2993 (N_2993,In_773,In_518);
or U2994 (N_2994,In_2227,In_955);
or U2995 (N_2995,In_2896,In_1108);
nor U2996 (N_2996,In_1933,In_1051);
nor U2997 (N_2997,In_2352,In_2421);
and U2998 (N_2998,In_2575,In_1701);
or U2999 (N_2999,In_751,In_1253);
nor U3000 (N_3000,In_807,In_2464);
or U3001 (N_3001,In_1609,In_1445);
and U3002 (N_3002,In_62,In_2076);
nor U3003 (N_3003,In_837,In_938);
or U3004 (N_3004,In_530,In_2103);
nand U3005 (N_3005,In_2875,In_679);
and U3006 (N_3006,In_1801,In_470);
and U3007 (N_3007,In_2316,In_2492);
nor U3008 (N_3008,In_2723,In_249);
or U3009 (N_3009,In_2166,In_1363);
nand U3010 (N_3010,In_147,In_1011);
or U3011 (N_3011,In_1303,In_2455);
nor U3012 (N_3012,In_2275,In_1055);
nand U3013 (N_3013,In_2299,In_1438);
nand U3014 (N_3014,In_2503,In_2705);
nand U3015 (N_3015,In_943,In_1460);
nand U3016 (N_3016,In_1828,In_1530);
nand U3017 (N_3017,In_1191,In_2480);
nand U3018 (N_3018,In_2019,In_2414);
nand U3019 (N_3019,In_78,In_738);
nor U3020 (N_3020,In_2326,In_206);
and U3021 (N_3021,In_2796,In_1894);
nand U3022 (N_3022,In_2048,In_600);
nand U3023 (N_3023,In_62,In_1576);
or U3024 (N_3024,In_612,In_2580);
and U3025 (N_3025,In_2872,In_563);
or U3026 (N_3026,In_331,In_1299);
and U3027 (N_3027,In_265,In_1730);
and U3028 (N_3028,In_2245,In_2990);
nand U3029 (N_3029,In_1,In_2332);
and U3030 (N_3030,In_2092,In_1595);
nand U3031 (N_3031,In_2838,In_2118);
or U3032 (N_3032,In_2284,In_1641);
or U3033 (N_3033,In_1824,In_296);
or U3034 (N_3034,In_1950,In_2575);
nor U3035 (N_3035,In_2062,In_2727);
or U3036 (N_3036,In_1616,In_1712);
and U3037 (N_3037,In_1485,In_540);
nor U3038 (N_3038,In_2475,In_1470);
or U3039 (N_3039,In_2255,In_1912);
and U3040 (N_3040,In_1417,In_2097);
or U3041 (N_3041,In_532,In_2752);
and U3042 (N_3042,In_2721,In_1673);
nand U3043 (N_3043,In_2373,In_640);
nand U3044 (N_3044,In_1796,In_2200);
or U3045 (N_3045,In_1548,In_1690);
and U3046 (N_3046,In_2928,In_874);
or U3047 (N_3047,In_627,In_2265);
or U3048 (N_3048,In_1023,In_2242);
nand U3049 (N_3049,In_148,In_965);
nand U3050 (N_3050,In_1290,In_2849);
and U3051 (N_3051,In_1053,In_2940);
nor U3052 (N_3052,In_138,In_528);
nand U3053 (N_3053,In_865,In_2574);
nor U3054 (N_3054,In_2860,In_833);
nor U3055 (N_3055,In_563,In_1990);
nand U3056 (N_3056,In_2466,In_2231);
nor U3057 (N_3057,In_1525,In_2051);
and U3058 (N_3058,In_2392,In_926);
nor U3059 (N_3059,In_1357,In_2511);
or U3060 (N_3060,In_275,In_1510);
nand U3061 (N_3061,In_2798,In_1635);
and U3062 (N_3062,In_1953,In_106);
nor U3063 (N_3063,In_637,In_1870);
nor U3064 (N_3064,In_2438,In_476);
nand U3065 (N_3065,In_2774,In_755);
nor U3066 (N_3066,In_592,In_2668);
nand U3067 (N_3067,In_133,In_688);
and U3068 (N_3068,In_1217,In_2457);
nor U3069 (N_3069,In_885,In_1361);
and U3070 (N_3070,In_1554,In_2301);
nand U3071 (N_3071,In_2551,In_196);
or U3072 (N_3072,In_275,In_2112);
nand U3073 (N_3073,In_1630,In_2554);
nor U3074 (N_3074,In_1474,In_144);
or U3075 (N_3075,In_667,In_43);
and U3076 (N_3076,In_2390,In_727);
or U3077 (N_3077,In_2070,In_2854);
and U3078 (N_3078,In_2435,In_2141);
nand U3079 (N_3079,In_347,In_345);
and U3080 (N_3080,In_1029,In_1854);
and U3081 (N_3081,In_2730,In_1836);
nor U3082 (N_3082,In_2275,In_2806);
nor U3083 (N_3083,In_2832,In_1273);
nor U3084 (N_3084,In_2001,In_1820);
and U3085 (N_3085,In_2480,In_2416);
nand U3086 (N_3086,In_2406,In_1625);
and U3087 (N_3087,In_937,In_2839);
or U3088 (N_3088,In_24,In_380);
nand U3089 (N_3089,In_2946,In_1725);
nand U3090 (N_3090,In_802,In_1201);
nor U3091 (N_3091,In_698,In_2310);
or U3092 (N_3092,In_230,In_848);
and U3093 (N_3093,In_2248,In_2584);
or U3094 (N_3094,In_2599,In_2395);
nand U3095 (N_3095,In_293,In_753);
nor U3096 (N_3096,In_2046,In_2202);
nor U3097 (N_3097,In_2261,In_510);
nor U3098 (N_3098,In_2989,In_438);
or U3099 (N_3099,In_1285,In_2621);
nand U3100 (N_3100,In_918,In_823);
nor U3101 (N_3101,In_2730,In_2763);
nand U3102 (N_3102,In_598,In_1588);
nor U3103 (N_3103,In_818,In_447);
nor U3104 (N_3104,In_1484,In_1232);
xnor U3105 (N_3105,In_310,In_1174);
nand U3106 (N_3106,In_485,In_1126);
and U3107 (N_3107,In_1280,In_276);
or U3108 (N_3108,In_508,In_296);
and U3109 (N_3109,In_2868,In_2176);
nor U3110 (N_3110,In_1867,In_365);
nand U3111 (N_3111,In_2888,In_2423);
nand U3112 (N_3112,In_926,In_85);
or U3113 (N_3113,In_823,In_1483);
or U3114 (N_3114,In_2844,In_1239);
nand U3115 (N_3115,In_2331,In_1081);
nor U3116 (N_3116,In_2130,In_2714);
nor U3117 (N_3117,In_1058,In_2474);
nor U3118 (N_3118,In_2047,In_1263);
and U3119 (N_3119,In_1644,In_2696);
and U3120 (N_3120,In_1914,In_1738);
nand U3121 (N_3121,In_1537,In_1399);
and U3122 (N_3122,In_2022,In_2259);
and U3123 (N_3123,In_2602,In_1766);
and U3124 (N_3124,In_666,In_1379);
or U3125 (N_3125,In_2221,In_546);
or U3126 (N_3126,In_1924,In_328);
nor U3127 (N_3127,In_2842,In_2045);
or U3128 (N_3128,In_1998,In_1276);
or U3129 (N_3129,In_2903,In_1064);
and U3130 (N_3130,In_2794,In_2206);
and U3131 (N_3131,In_606,In_2747);
or U3132 (N_3132,In_1529,In_830);
nor U3133 (N_3133,In_1472,In_1229);
or U3134 (N_3134,In_2069,In_2619);
nand U3135 (N_3135,In_2601,In_195);
and U3136 (N_3136,In_1365,In_1218);
nor U3137 (N_3137,In_421,In_1572);
nor U3138 (N_3138,In_1511,In_817);
nand U3139 (N_3139,In_498,In_855);
or U3140 (N_3140,In_1179,In_1990);
nor U3141 (N_3141,In_1561,In_125);
nor U3142 (N_3142,In_973,In_609);
or U3143 (N_3143,In_1082,In_524);
or U3144 (N_3144,In_757,In_2721);
nor U3145 (N_3145,In_651,In_2714);
nor U3146 (N_3146,In_2290,In_446);
or U3147 (N_3147,In_2682,In_1445);
or U3148 (N_3148,In_1596,In_1486);
nand U3149 (N_3149,In_1954,In_2761);
nor U3150 (N_3150,In_64,In_1273);
and U3151 (N_3151,In_78,In_1166);
or U3152 (N_3152,In_904,In_861);
and U3153 (N_3153,In_2724,In_2631);
nor U3154 (N_3154,In_324,In_2311);
and U3155 (N_3155,In_2344,In_2067);
or U3156 (N_3156,In_1782,In_1764);
and U3157 (N_3157,In_1722,In_614);
and U3158 (N_3158,In_1328,In_243);
nand U3159 (N_3159,In_552,In_2899);
nor U3160 (N_3160,In_757,In_1560);
or U3161 (N_3161,In_2391,In_1049);
nor U3162 (N_3162,In_1869,In_1971);
nor U3163 (N_3163,In_362,In_1369);
and U3164 (N_3164,In_2310,In_1807);
and U3165 (N_3165,In_2213,In_844);
nand U3166 (N_3166,In_692,In_1346);
nor U3167 (N_3167,In_1575,In_2010);
nand U3168 (N_3168,In_2984,In_2927);
and U3169 (N_3169,In_2742,In_2320);
nor U3170 (N_3170,In_1738,In_2164);
or U3171 (N_3171,In_917,In_2877);
or U3172 (N_3172,In_2860,In_2723);
nand U3173 (N_3173,In_2169,In_801);
nand U3174 (N_3174,In_2482,In_2563);
nand U3175 (N_3175,In_1246,In_451);
and U3176 (N_3176,In_463,In_7);
and U3177 (N_3177,In_1768,In_1818);
and U3178 (N_3178,In_1877,In_1711);
and U3179 (N_3179,In_1805,In_1684);
or U3180 (N_3180,In_651,In_2577);
nand U3181 (N_3181,In_1597,In_2063);
xnor U3182 (N_3182,In_2527,In_122);
and U3183 (N_3183,In_2836,In_1495);
nor U3184 (N_3184,In_847,In_2808);
and U3185 (N_3185,In_2849,In_2428);
nor U3186 (N_3186,In_2629,In_2021);
nor U3187 (N_3187,In_1458,In_906);
and U3188 (N_3188,In_738,In_430);
nor U3189 (N_3189,In_1448,In_196);
and U3190 (N_3190,In_548,In_1688);
or U3191 (N_3191,In_1897,In_1186);
and U3192 (N_3192,In_1759,In_451);
nor U3193 (N_3193,In_61,In_390);
or U3194 (N_3194,In_1738,In_2873);
or U3195 (N_3195,In_2077,In_936);
or U3196 (N_3196,In_1936,In_1606);
nand U3197 (N_3197,In_710,In_180);
nand U3198 (N_3198,In_739,In_9);
or U3199 (N_3199,In_1291,In_2239);
and U3200 (N_3200,In_447,In_1076);
or U3201 (N_3201,In_1081,In_612);
nor U3202 (N_3202,In_1164,In_2103);
or U3203 (N_3203,In_848,In_1272);
or U3204 (N_3204,In_1765,In_37);
nor U3205 (N_3205,In_2398,In_1550);
and U3206 (N_3206,In_1009,In_2703);
and U3207 (N_3207,In_1648,In_1045);
nor U3208 (N_3208,In_2157,In_1362);
or U3209 (N_3209,In_1809,In_597);
nor U3210 (N_3210,In_2737,In_2463);
or U3211 (N_3211,In_253,In_2226);
and U3212 (N_3212,In_640,In_2563);
and U3213 (N_3213,In_2395,In_2837);
or U3214 (N_3214,In_2939,In_2040);
nand U3215 (N_3215,In_1253,In_1898);
and U3216 (N_3216,In_754,In_242);
nand U3217 (N_3217,In_2701,In_2147);
and U3218 (N_3218,In_1009,In_2402);
nand U3219 (N_3219,In_2977,In_1753);
and U3220 (N_3220,In_2502,In_1735);
nor U3221 (N_3221,In_1358,In_1497);
nor U3222 (N_3222,In_240,In_1406);
nor U3223 (N_3223,In_314,In_2812);
nand U3224 (N_3224,In_2180,In_1414);
nand U3225 (N_3225,In_2200,In_1162);
nand U3226 (N_3226,In_580,In_2116);
and U3227 (N_3227,In_902,In_1493);
nor U3228 (N_3228,In_2156,In_2676);
or U3229 (N_3229,In_1784,In_857);
nand U3230 (N_3230,In_1214,In_1776);
or U3231 (N_3231,In_2601,In_2948);
nand U3232 (N_3232,In_2206,In_2025);
nor U3233 (N_3233,In_2388,In_2712);
and U3234 (N_3234,In_1532,In_2315);
or U3235 (N_3235,In_1880,In_2271);
and U3236 (N_3236,In_1432,In_46);
nor U3237 (N_3237,In_2942,In_2251);
nand U3238 (N_3238,In_1317,In_1713);
nor U3239 (N_3239,In_1972,In_1184);
and U3240 (N_3240,In_436,In_2940);
nand U3241 (N_3241,In_1360,In_2930);
or U3242 (N_3242,In_858,In_2411);
or U3243 (N_3243,In_1223,In_1290);
and U3244 (N_3244,In_2065,In_1364);
nand U3245 (N_3245,In_1081,In_450);
or U3246 (N_3246,In_448,In_2176);
or U3247 (N_3247,In_2420,In_1267);
or U3248 (N_3248,In_2832,In_1387);
nor U3249 (N_3249,In_1342,In_1023);
nor U3250 (N_3250,In_2997,In_415);
nor U3251 (N_3251,In_2083,In_1062);
and U3252 (N_3252,In_1178,In_2922);
or U3253 (N_3253,In_785,In_997);
nand U3254 (N_3254,In_1531,In_1341);
and U3255 (N_3255,In_1245,In_2799);
or U3256 (N_3256,In_406,In_771);
or U3257 (N_3257,In_1174,In_2065);
and U3258 (N_3258,In_430,In_1216);
and U3259 (N_3259,In_2902,In_851);
nand U3260 (N_3260,In_199,In_2444);
nor U3261 (N_3261,In_1664,In_335);
and U3262 (N_3262,In_139,In_662);
nor U3263 (N_3263,In_2140,In_1191);
and U3264 (N_3264,In_2730,In_1826);
nor U3265 (N_3265,In_2740,In_1521);
and U3266 (N_3266,In_619,In_490);
or U3267 (N_3267,In_2076,In_2333);
and U3268 (N_3268,In_529,In_1512);
and U3269 (N_3269,In_1372,In_2096);
or U3270 (N_3270,In_2147,In_1483);
nand U3271 (N_3271,In_1024,In_2463);
nor U3272 (N_3272,In_2611,In_1581);
nand U3273 (N_3273,In_2739,In_2192);
and U3274 (N_3274,In_2759,In_2618);
nor U3275 (N_3275,In_887,In_112);
and U3276 (N_3276,In_504,In_1156);
nor U3277 (N_3277,In_2215,In_2108);
or U3278 (N_3278,In_1086,In_761);
nand U3279 (N_3279,In_2124,In_781);
nor U3280 (N_3280,In_2232,In_1560);
and U3281 (N_3281,In_151,In_1376);
and U3282 (N_3282,In_744,In_1630);
nor U3283 (N_3283,In_2628,In_1065);
nand U3284 (N_3284,In_202,In_2470);
nor U3285 (N_3285,In_2135,In_1145);
nor U3286 (N_3286,In_2382,In_1953);
and U3287 (N_3287,In_2,In_1343);
and U3288 (N_3288,In_448,In_69);
and U3289 (N_3289,In_2410,In_1506);
nor U3290 (N_3290,In_1095,In_1091);
nand U3291 (N_3291,In_2418,In_2805);
and U3292 (N_3292,In_1995,In_1888);
nor U3293 (N_3293,In_1309,In_821);
or U3294 (N_3294,In_1639,In_2283);
nor U3295 (N_3295,In_1518,In_1679);
nor U3296 (N_3296,In_1879,In_1819);
or U3297 (N_3297,In_702,In_322);
and U3298 (N_3298,In_1800,In_2411);
or U3299 (N_3299,In_114,In_245);
and U3300 (N_3300,In_1010,In_1307);
or U3301 (N_3301,In_2580,In_241);
or U3302 (N_3302,In_2151,In_1947);
or U3303 (N_3303,In_496,In_946);
nor U3304 (N_3304,In_249,In_1016);
or U3305 (N_3305,In_1422,In_1516);
and U3306 (N_3306,In_762,In_2765);
nand U3307 (N_3307,In_1600,In_582);
and U3308 (N_3308,In_15,In_2892);
nand U3309 (N_3309,In_1689,In_2139);
nand U3310 (N_3310,In_825,In_1935);
and U3311 (N_3311,In_1182,In_538);
or U3312 (N_3312,In_1745,In_1739);
nand U3313 (N_3313,In_1131,In_1650);
or U3314 (N_3314,In_1916,In_1074);
and U3315 (N_3315,In_2098,In_1880);
nand U3316 (N_3316,In_1908,In_9);
or U3317 (N_3317,In_818,In_226);
nor U3318 (N_3318,In_2220,In_375);
nor U3319 (N_3319,In_940,In_1149);
or U3320 (N_3320,In_2434,In_2069);
and U3321 (N_3321,In_1392,In_2222);
nand U3322 (N_3322,In_50,In_731);
or U3323 (N_3323,In_2441,In_676);
xnor U3324 (N_3324,In_1693,In_1489);
xnor U3325 (N_3325,In_1006,In_2180);
nand U3326 (N_3326,In_1976,In_2833);
nor U3327 (N_3327,In_1300,In_2228);
and U3328 (N_3328,In_1064,In_432);
nor U3329 (N_3329,In_2696,In_1327);
nand U3330 (N_3330,In_869,In_92);
nor U3331 (N_3331,In_1172,In_1963);
or U3332 (N_3332,In_2200,In_675);
or U3333 (N_3333,In_2884,In_2604);
and U3334 (N_3334,In_2040,In_220);
nand U3335 (N_3335,In_1139,In_312);
or U3336 (N_3336,In_2543,In_2275);
nor U3337 (N_3337,In_322,In_1785);
and U3338 (N_3338,In_985,In_2209);
or U3339 (N_3339,In_2995,In_2459);
and U3340 (N_3340,In_469,In_124);
or U3341 (N_3341,In_2956,In_597);
nor U3342 (N_3342,In_2590,In_507);
nor U3343 (N_3343,In_2129,In_13);
and U3344 (N_3344,In_269,In_627);
or U3345 (N_3345,In_2229,In_227);
nand U3346 (N_3346,In_218,In_1902);
nor U3347 (N_3347,In_1941,In_2579);
nand U3348 (N_3348,In_905,In_2855);
nor U3349 (N_3349,In_1684,In_1037);
nor U3350 (N_3350,In_2370,In_842);
nor U3351 (N_3351,In_1147,In_778);
nor U3352 (N_3352,In_481,In_353);
nor U3353 (N_3353,In_532,In_1793);
and U3354 (N_3354,In_1363,In_1462);
nor U3355 (N_3355,In_1083,In_55);
nor U3356 (N_3356,In_130,In_2678);
nor U3357 (N_3357,In_348,In_2123);
nand U3358 (N_3358,In_38,In_634);
and U3359 (N_3359,In_2178,In_879);
nand U3360 (N_3360,In_1770,In_230);
and U3361 (N_3361,In_2848,In_1006);
nand U3362 (N_3362,In_759,In_2260);
nor U3363 (N_3363,In_2685,In_813);
xnor U3364 (N_3364,In_1486,In_684);
and U3365 (N_3365,In_2783,In_955);
and U3366 (N_3366,In_2435,In_256);
nand U3367 (N_3367,In_1813,In_252);
and U3368 (N_3368,In_2809,In_2911);
nor U3369 (N_3369,In_2029,In_1878);
nand U3370 (N_3370,In_1727,In_1251);
nand U3371 (N_3371,In_1315,In_2873);
nand U3372 (N_3372,In_217,In_1561);
nor U3373 (N_3373,In_1194,In_2615);
and U3374 (N_3374,In_941,In_2273);
nand U3375 (N_3375,In_618,In_1151);
nor U3376 (N_3376,In_980,In_95);
nand U3377 (N_3377,In_1213,In_2556);
or U3378 (N_3378,In_1233,In_1301);
nand U3379 (N_3379,In_6,In_1116);
or U3380 (N_3380,In_2111,In_1099);
nor U3381 (N_3381,In_1031,In_292);
nor U3382 (N_3382,In_896,In_2182);
xnor U3383 (N_3383,In_259,In_1486);
and U3384 (N_3384,In_403,In_2694);
nor U3385 (N_3385,In_1665,In_623);
and U3386 (N_3386,In_532,In_230);
nand U3387 (N_3387,In_308,In_1712);
nand U3388 (N_3388,In_247,In_818);
nand U3389 (N_3389,In_2498,In_2406);
or U3390 (N_3390,In_2744,In_2217);
and U3391 (N_3391,In_1956,In_2890);
nand U3392 (N_3392,In_2586,In_1658);
nor U3393 (N_3393,In_303,In_2128);
nor U3394 (N_3394,In_1483,In_1404);
nand U3395 (N_3395,In_551,In_97);
nor U3396 (N_3396,In_544,In_1947);
and U3397 (N_3397,In_1772,In_420);
nor U3398 (N_3398,In_2592,In_2381);
or U3399 (N_3399,In_1383,In_1780);
and U3400 (N_3400,In_1364,In_255);
or U3401 (N_3401,In_2825,In_2192);
nand U3402 (N_3402,In_1647,In_146);
or U3403 (N_3403,In_1189,In_2113);
nor U3404 (N_3404,In_123,In_2135);
or U3405 (N_3405,In_491,In_2574);
nor U3406 (N_3406,In_2456,In_2325);
and U3407 (N_3407,In_1682,In_467);
and U3408 (N_3408,In_1620,In_1133);
and U3409 (N_3409,In_1488,In_1760);
or U3410 (N_3410,In_798,In_514);
nor U3411 (N_3411,In_1162,In_2077);
or U3412 (N_3412,In_722,In_1566);
nor U3413 (N_3413,In_1932,In_1618);
nand U3414 (N_3414,In_1159,In_898);
and U3415 (N_3415,In_1552,In_2531);
xnor U3416 (N_3416,In_2280,In_2822);
nand U3417 (N_3417,In_597,In_2048);
or U3418 (N_3418,In_877,In_1573);
nor U3419 (N_3419,In_1530,In_2155);
nor U3420 (N_3420,In_40,In_494);
or U3421 (N_3421,In_2291,In_2654);
nor U3422 (N_3422,In_414,In_733);
nor U3423 (N_3423,In_2794,In_944);
or U3424 (N_3424,In_2651,In_91);
or U3425 (N_3425,In_390,In_83);
nor U3426 (N_3426,In_2706,In_2540);
and U3427 (N_3427,In_655,In_2767);
or U3428 (N_3428,In_14,In_326);
and U3429 (N_3429,In_221,In_2535);
nand U3430 (N_3430,In_1741,In_520);
or U3431 (N_3431,In_2404,In_568);
or U3432 (N_3432,In_539,In_1552);
or U3433 (N_3433,In_808,In_2706);
or U3434 (N_3434,In_1327,In_2656);
or U3435 (N_3435,In_1519,In_231);
nor U3436 (N_3436,In_2617,In_1625);
nor U3437 (N_3437,In_614,In_2793);
nand U3438 (N_3438,In_153,In_765);
nand U3439 (N_3439,In_2436,In_35);
nor U3440 (N_3440,In_2365,In_2217);
and U3441 (N_3441,In_380,In_591);
and U3442 (N_3442,In_2438,In_1752);
and U3443 (N_3443,In_2682,In_1412);
and U3444 (N_3444,In_145,In_1547);
nand U3445 (N_3445,In_206,In_1915);
nand U3446 (N_3446,In_2271,In_2220);
and U3447 (N_3447,In_1858,In_424);
or U3448 (N_3448,In_2228,In_2060);
nor U3449 (N_3449,In_1503,In_1602);
nor U3450 (N_3450,In_2183,In_380);
nor U3451 (N_3451,In_2033,In_2832);
nand U3452 (N_3452,In_183,In_502);
nand U3453 (N_3453,In_2990,In_2267);
or U3454 (N_3454,In_1181,In_175);
nor U3455 (N_3455,In_1274,In_418);
nor U3456 (N_3456,In_1355,In_1264);
and U3457 (N_3457,In_2876,In_251);
nor U3458 (N_3458,In_1527,In_861);
or U3459 (N_3459,In_2563,In_996);
or U3460 (N_3460,In_123,In_2854);
or U3461 (N_3461,In_2626,In_1936);
and U3462 (N_3462,In_2123,In_2170);
nand U3463 (N_3463,In_1928,In_1515);
nor U3464 (N_3464,In_2352,In_2626);
nor U3465 (N_3465,In_2264,In_2868);
nor U3466 (N_3466,In_2132,In_492);
nand U3467 (N_3467,In_1243,In_896);
nor U3468 (N_3468,In_2902,In_1612);
nand U3469 (N_3469,In_379,In_2);
and U3470 (N_3470,In_2067,In_1982);
nand U3471 (N_3471,In_2738,In_2362);
nor U3472 (N_3472,In_621,In_60);
nor U3473 (N_3473,In_1008,In_936);
or U3474 (N_3474,In_2769,In_2222);
and U3475 (N_3475,In_552,In_233);
and U3476 (N_3476,In_2983,In_1248);
nand U3477 (N_3477,In_2546,In_783);
nand U3478 (N_3478,In_717,In_1472);
xor U3479 (N_3479,In_2455,In_1754);
or U3480 (N_3480,In_433,In_1205);
nor U3481 (N_3481,In_960,In_2732);
nand U3482 (N_3482,In_1022,In_1542);
and U3483 (N_3483,In_655,In_1051);
and U3484 (N_3484,In_1756,In_1617);
nand U3485 (N_3485,In_2457,In_190);
and U3486 (N_3486,In_2245,In_2081);
or U3487 (N_3487,In_1550,In_1019);
nand U3488 (N_3488,In_624,In_978);
or U3489 (N_3489,In_100,In_1362);
and U3490 (N_3490,In_617,In_775);
xnor U3491 (N_3491,In_1598,In_641);
and U3492 (N_3492,In_2759,In_1240);
nor U3493 (N_3493,In_819,In_2263);
nand U3494 (N_3494,In_496,In_2834);
nor U3495 (N_3495,In_532,In_1057);
and U3496 (N_3496,In_2729,In_1576);
nand U3497 (N_3497,In_1865,In_1603);
nor U3498 (N_3498,In_2714,In_2195);
or U3499 (N_3499,In_2608,In_2906);
nand U3500 (N_3500,In_2812,In_1462);
nor U3501 (N_3501,In_1005,In_973);
nor U3502 (N_3502,In_2335,In_2018);
or U3503 (N_3503,In_2349,In_322);
and U3504 (N_3504,In_1218,In_2024);
or U3505 (N_3505,In_1369,In_1534);
nor U3506 (N_3506,In_2230,In_1893);
and U3507 (N_3507,In_38,In_386);
and U3508 (N_3508,In_824,In_2995);
or U3509 (N_3509,In_551,In_600);
nand U3510 (N_3510,In_1715,In_582);
or U3511 (N_3511,In_1106,In_1844);
or U3512 (N_3512,In_2357,In_1796);
nand U3513 (N_3513,In_235,In_54);
or U3514 (N_3514,In_2943,In_2892);
or U3515 (N_3515,In_384,In_403);
or U3516 (N_3516,In_2897,In_2242);
or U3517 (N_3517,In_1537,In_2908);
and U3518 (N_3518,In_672,In_1142);
and U3519 (N_3519,In_2974,In_2076);
xnor U3520 (N_3520,In_2969,In_1003);
or U3521 (N_3521,In_2004,In_1836);
or U3522 (N_3522,In_622,In_923);
and U3523 (N_3523,In_1333,In_2582);
and U3524 (N_3524,In_761,In_1468);
nand U3525 (N_3525,In_2294,In_1622);
and U3526 (N_3526,In_125,In_1843);
or U3527 (N_3527,In_975,In_83);
nor U3528 (N_3528,In_2740,In_522);
and U3529 (N_3529,In_1761,In_1735);
or U3530 (N_3530,In_973,In_2967);
and U3531 (N_3531,In_2927,In_1448);
nand U3532 (N_3532,In_903,In_1953);
nand U3533 (N_3533,In_180,In_2074);
nand U3534 (N_3534,In_2463,In_2174);
nand U3535 (N_3535,In_2332,In_2473);
nand U3536 (N_3536,In_2674,In_1228);
nor U3537 (N_3537,In_338,In_687);
nand U3538 (N_3538,In_1198,In_2671);
xnor U3539 (N_3539,In_925,In_897);
or U3540 (N_3540,In_1457,In_2293);
nor U3541 (N_3541,In_1529,In_2291);
nand U3542 (N_3542,In_2735,In_1067);
nor U3543 (N_3543,In_1481,In_1668);
nor U3544 (N_3544,In_577,In_2924);
or U3545 (N_3545,In_2510,In_2955);
nand U3546 (N_3546,In_1881,In_293);
and U3547 (N_3547,In_217,In_2073);
or U3548 (N_3548,In_1210,In_973);
and U3549 (N_3549,In_1484,In_739);
nor U3550 (N_3550,In_1379,In_1999);
or U3551 (N_3551,In_1702,In_2258);
or U3552 (N_3552,In_2754,In_103);
or U3553 (N_3553,In_2276,In_1539);
or U3554 (N_3554,In_26,In_532);
or U3555 (N_3555,In_532,In_272);
nor U3556 (N_3556,In_2321,In_582);
and U3557 (N_3557,In_1157,In_636);
nand U3558 (N_3558,In_118,In_2394);
nor U3559 (N_3559,In_1795,In_1218);
or U3560 (N_3560,In_1005,In_1354);
nor U3561 (N_3561,In_1592,In_2167);
nor U3562 (N_3562,In_2107,In_2490);
or U3563 (N_3563,In_558,In_2049);
nor U3564 (N_3564,In_2073,In_2276);
or U3565 (N_3565,In_2046,In_1995);
nand U3566 (N_3566,In_1085,In_1561);
or U3567 (N_3567,In_1473,In_1801);
nor U3568 (N_3568,In_814,In_737);
and U3569 (N_3569,In_2144,In_1176);
nand U3570 (N_3570,In_1620,In_108);
and U3571 (N_3571,In_1402,In_654);
nand U3572 (N_3572,In_2501,In_1281);
nand U3573 (N_3573,In_1899,In_973);
or U3574 (N_3574,In_1058,In_919);
or U3575 (N_3575,In_1301,In_530);
and U3576 (N_3576,In_1565,In_347);
or U3577 (N_3577,In_2465,In_2999);
nand U3578 (N_3578,In_2802,In_2041);
and U3579 (N_3579,In_436,In_424);
and U3580 (N_3580,In_237,In_518);
or U3581 (N_3581,In_1647,In_2159);
nand U3582 (N_3582,In_542,In_540);
nor U3583 (N_3583,In_2686,In_2334);
and U3584 (N_3584,In_2938,In_389);
nor U3585 (N_3585,In_2773,In_2812);
nand U3586 (N_3586,In_108,In_1495);
nor U3587 (N_3587,In_1448,In_797);
nor U3588 (N_3588,In_737,In_2710);
nand U3589 (N_3589,In_1240,In_127);
nor U3590 (N_3590,In_822,In_1850);
nand U3591 (N_3591,In_2739,In_1921);
and U3592 (N_3592,In_2174,In_1511);
nor U3593 (N_3593,In_899,In_382);
or U3594 (N_3594,In_1534,In_2892);
nand U3595 (N_3595,In_1560,In_1959);
nand U3596 (N_3596,In_647,In_1393);
nand U3597 (N_3597,In_2413,In_2142);
or U3598 (N_3598,In_1388,In_1577);
or U3599 (N_3599,In_981,In_390);
nand U3600 (N_3600,In_1353,In_1340);
nand U3601 (N_3601,In_577,In_484);
and U3602 (N_3602,In_2589,In_182);
and U3603 (N_3603,In_1355,In_1659);
and U3604 (N_3604,In_564,In_44);
and U3605 (N_3605,In_570,In_966);
nand U3606 (N_3606,In_309,In_440);
nor U3607 (N_3607,In_2807,In_2938);
nor U3608 (N_3608,In_2304,In_1776);
nand U3609 (N_3609,In_970,In_389);
or U3610 (N_3610,In_178,In_2198);
nand U3611 (N_3611,In_2471,In_2024);
or U3612 (N_3612,In_344,In_2162);
nor U3613 (N_3613,In_1811,In_130);
nand U3614 (N_3614,In_800,In_2311);
nor U3615 (N_3615,In_1592,In_2297);
or U3616 (N_3616,In_1909,In_1740);
nand U3617 (N_3617,In_35,In_1289);
and U3618 (N_3618,In_1687,In_1849);
or U3619 (N_3619,In_1081,In_1318);
nand U3620 (N_3620,In_498,In_2104);
and U3621 (N_3621,In_2996,In_2031);
nand U3622 (N_3622,In_2558,In_762);
nor U3623 (N_3623,In_6,In_1484);
and U3624 (N_3624,In_1266,In_2143);
nand U3625 (N_3625,In_2073,In_2055);
or U3626 (N_3626,In_403,In_556);
and U3627 (N_3627,In_957,In_2755);
nand U3628 (N_3628,In_2548,In_844);
nor U3629 (N_3629,In_1728,In_735);
and U3630 (N_3630,In_1097,In_2002);
nand U3631 (N_3631,In_623,In_1892);
or U3632 (N_3632,In_912,In_2360);
nand U3633 (N_3633,In_184,In_275);
nor U3634 (N_3634,In_1958,In_1345);
and U3635 (N_3635,In_2791,In_2044);
and U3636 (N_3636,In_1157,In_1910);
nand U3637 (N_3637,In_2651,In_1725);
nand U3638 (N_3638,In_1044,In_2230);
and U3639 (N_3639,In_2368,In_1062);
and U3640 (N_3640,In_1249,In_2632);
nand U3641 (N_3641,In_1025,In_1044);
and U3642 (N_3642,In_2620,In_2142);
nand U3643 (N_3643,In_437,In_1057);
or U3644 (N_3644,In_2062,In_2176);
nor U3645 (N_3645,In_1637,In_2467);
nand U3646 (N_3646,In_553,In_332);
and U3647 (N_3647,In_2300,In_2899);
nor U3648 (N_3648,In_1806,In_821);
nor U3649 (N_3649,In_2742,In_2951);
nand U3650 (N_3650,In_2581,In_1881);
nand U3651 (N_3651,In_340,In_1863);
nor U3652 (N_3652,In_1664,In_714);
or U3653 (N_3653,In_2317,In_1759);
nor U3654 (N_3654,In_1356,In_1788);
nand U3655 (N_3655,In_858,In_2832);
nor U3656 (N_3656,In_2183,In_1656);
and U3657 (N_3657,In_647,In_1152);
or U3658 (N_3658,In_1162,In_2731);
nand U3659 (N_3659,In_467,In_1569);
nor U3660 (N_3660,In_1925,In_1821);
and U3661 (N_3661,In_2304,In_1491);
xnor U3662 (N_3662,In_1465,In_1661);
xor U3663 (N_3663,In_321,In_2960);
nand U3664 (N_3664,In_2669,In_818);
nand U3665 (N_3665,In_1784,In_1082);
or U3666 (N_3666,In_2919,In_631);
and U3667 (N_3667,In_2144,In_1198);
xor U3668 (N_3668,In_2082,In_2565);
and U3669 (N_3669,In_2506,In_654);
and U3670 (N_3670,In_2880,In_846);
or U3671 (N_3671,In_1189,In_2680);
and U3672 (N_3672,In_2699,In_88);
nor U3673 (N_3673,In_1549,In_1502);
and U3674 (N_3674,In_372,In_1845);
nor U3675 (N_3675,In_1078,In_180);
and U3676 (N_3676,In_2566,In_494);
and U3677 (N_3677,In_1368,In_155);
or U3678 (N_3678,In_287,In_1275);
nand U3679 (N_3679,In_1159,In_2901);
nor U3680 (N_3680,In_2585,In_2951);
and U3681 (N_3681,In_39,In_126);
and U3682 (N_3682,In_1814,In_2459);
nor U3683 (N_3683,In_1314,In_902);
or U3684 (N_3684,In_1372,In_2267);
nand U3685 (N_3685,In_587,In_2858);
nand U3686 (N_3686,In_2120,In_1213);
or U3687 (N_3687,In_1615,In_1059);
nor U3688 (N_3688,In_2654,In_2816);
nor U3689 (N_3689,In_2175,In_1570);
nor U3690 (N_3690,In_1584,In_1721);
or U3691 (N_3691,In_2032,In_918);
or U3692 (N_3692,In_1233,In_2566);
and U3693 (N_3693,In_2976,In_1829);
nand U3694 (N_3694,In_1707,In_2461);
or U3695 (N_3695,In_537,In_273);
or U3696 (N_3696,In_1548,In_1349);
and U3697 (N_3697,In_2272,In_2166);
and U3698 (N_3698,In_158,In_162);
or U3699 (N_3699,In_1683,In_1030);
nor U3700 (N_3700,In_870,In_1306);
nor U3701 (N_3701,In_2941,In_374);
nand U3702 (N_3702,In_2395,In_339);
and U3703 (N_3703,In_1358,In_2472);
or U3704 (N_3704,In_1620,In_2246);
nor U3705 (N_3705,In_1499,In_1078);
or U3706 (N_3706,In_2718,In_2234);
nor U3707 (N_3707,In_1631,In_2943);
and U3708 (N_3708,In_2591,In_151);
or U3709 (N_3709,In_2501,In_1431);
nor U3710 (N_3710,In_2757,In_1386);
or U3711 (N_3711,In_74,In_745);
and U3712 (N_3712,In_949,In_2842);
nand U3713 (N_3713,In_2665,In_980);
nand U3714 (N_3714,In_1837,In_374);
or U3715 (N_3715,In_552,In_2031);
and U3716 (N_3716,In_2440,In_699);
and U3717 (N_3717,In_429,In_2726);
or U3718 (N_3718,In_1391,In_646);
and U3719 (N_3719,In_2893,In_1239);
nor U3720 (N_3720,In_1418,In_1171);
nand U3721 (N_3721,In_2948,In_740);
nor U3722 (N_3722,In_2458,In_703);
or U3723 (N_3723,In_1483,In_2841);
and U3724 (N_3724,In_2349,In_804);
nand U3725 (N_3725,In_2690,In_2962);
and U3726 (N_3726,In_1052,In_240);
or U3727 (N_3727,In_1396,In_1185);
and U3728 (N_3728,In_457,In_1249);
nand U3729 (N_3729,In_981,In_1391);
nand U3730 (N_3730,In_406,In_2467);
nand U3731 (N_3731,In_736,In_301);
nor U3732 (N_3732,In_2768,In_357);
and U3733 (N_3733,In_644,In_2620);
nor U3734 (N_3734,In_848,In_1757);
nor U3735 (N_3735,In_2245,In_942);
and U3736 (N_3736,In_751,In_1233);
nand U3737 (N_3737,In_2179,In_707);
and U3738 (N_3738,In_1404,In_879);
and U3739 (N_3739,In_955,In_260);
nor U3740 (N_3740,In_2066,In_996);
nand U3741 (N_3741,In_262,In_1330);
nor U3742 (N_3742,In_1502,In_1676);
nor U3743 (N_3743,In_136,In_1754);
nor U3744 (N_3744,In_368,In_1163);
or U3745 (N_3745,In_2717,In_2515);
and U3746 (N_3746,In_2897,In_2234);
nor U3747 (N_3747,In_1648,In_1154);
nor U3748 (N_3748,In_2266,In_2835);
nor U3749 (N_3749,In_2265,In_2680);
nor U3750 (N_3750,In_2432,In_1091);
and U3751 (N_3751,In_1601,In_500);
or U3752 (N_3752,In_1811,In_108);
or U3753 (N_3753,In_2227,In_2909);
nand U3754 (N_3754,In_1575,In_2028);
and U3755 (N_3755,In_383,In_2535);
nand U3756 (N_3756,In_2613,In_2799);
nand U3757 (N_3757,In_1253,In_370);
and U3758 (N_3758,In_822,In_2378);
and U3759 (N_3759,In_1544,In_736);
nand U3760 (N_3760,In_2114,In_1001);
nand U3761 (N_3761,In_1635,In_2477);
or U3762 (N_3762,In_2667,In_273);
nor U3763 (N_3763,In_785,In_1871);
nand U3764 (N_3764,In_84,In_2227);
nor U3765 (N_3765,In_824,In_1471);
nor U3766 (N_3766,In_2349,In_33);
or U3767 (N_3767,In_1233,In_755);
and U3768 (N_3768,In_154,In_439);
xor U3769 (N_3769,In_1102,In_1785);
and U3770 (N_3770,In_2452,In_972);
or U3771 (N_3771,In_97,In_36);
or U3772 (N_3772,In_1653,In_2773);
or U3773 (N_3773,In_1522,In_2761);
nand U3774 (N_3774,In_1628,In_2942);
nor U3775 (N_3775,In_862,In_453);
or U3776 (N_3776,In_1285,In_128);
and U3777 (N_3777,In_1952,In_2793);
nand U3778 (N_3778,In_884,In_2490);
nor U3779 (N_3779,In_1214,In_2617);
and U3780 (N_3780,In_2852,In_2731);
nand U3781 (N_3781,In_976,In_525);
or U3782 (N_3782,In_1648,In_2240);
nand U3783 (N_3783,In_1244,In_1694);
nand U3784 (N_3784,In_1869,In_2503);
nand U3785 (N_3785,In_1230,In_414);
or U3786 (N_3786,In_1173,In_1034);
nor U3787 (N_3787,In_2865,In_2545);
and U3788 (N_3788,In_2319,In_699);
or U3789 (N_3789,In_1698,In_478);
or U3790 (N_3790,In_2105,In_2435);
nor U3791 (N_3791,In_1329,In_1946);
nand U3792 (N_3792,In_863,In_1561);
nand U3793 (N_3793,In_569,In_2069);
or U3794 (N_3794,In_1000,In_705);
or U3795 (N_3795,In_1708,In_1268);
and U3796 (N_3796,In_2635,In_461);
nand U3797 (N_3797,In_384,In_602);
nor U3798 (N_3798,In_1486,In_1560);
nand U3799 (N_3799,In_2337,In_2943);
nor U3800 (N_3800,In_906,In_2821);
or U3801 (N_3801,In_2739,In_1988);
and U3802 (N_3802,In_2130,In_959);
nand U3803 (N_3803,In_1087,In_951);
or U3804 (N_3804,In_490,In_1861);
or U3805 (N_3805,In_2143,In_2696);
and U3806 (N_3806,In_278,In_2465);
and U3807 (N_3807,In_2313,In_1284);
and U3808 (N_3808,In_1585,In_1995);
nand U3809 (N_3809,In_146,In_1376);
or U3810 (N_3810,In_1767,In_1900);
nand U3811 (N_3811,In_144,In_2889);
and U3812 (N_3812,In_2252,In_16);
nor U3813 (N_3813,In_141,In_579);
nor U3814 (N_3814,In_431,In_888);
or U3815 (N_3815,In_581,In_1693);
or U3816 (N_3816,In_2484,In_2427);
nand U3817 (N_3817,In_1757,In_643);
and U3818 (N_3818,In_2590,In_1317);
nand U3819 (N_3819,In_817,In_2689);
or U3820 (N_3820,In_1154,In_253);
or U3821 (N_3821,In_2279,In_2869);
or U3822 (N_3822,In_2858,In_313);
nand U3823 (N_3823,In_1514,In_1519);
or U3824 (N_3824,In_841,In_73);
and U3825 (N_3825,In_246,In_546);
nor U3826 (N_3826,In_1292,In_2593);
nand U3827 (N_3827,In_2473,In_2440);
nor U3828 (N_3828,In_1476,In_2026);
nand U3829 (N_3829,In_2243,In_2045);
or U3830 (N_3830,In_1354,In_815);
xor U3831 (N_3831,In_1247,In_1971);
nand U3832 (N_3832,In_792,In_1678);
and U3833 (N_3833,In_1380,In_2131);
and U3834 (N_3834,In_2493,In_2706);
nand U3835 (N_3835,In_1545,In_1006);
and U3836 (N_3836,In_716,In_727);
nor U3837 (N_3837,In_2135,In_1320);
or U3838 (N_3838,In_1144,In_2634);
or U3839 (N_3839,In_1558,In_277);
nand U3840 (N_3840,In_909,In_2385);
nor U3841 (N_3841,In_2144,In_1113);
or U3842 (N_3842,In_2308,In_1650);
and U3843 (N_3843,In_2177,In_185);
and U3844 (N_3844,In_668,In_745);
or U3845 (N_3845,In_2002,In_114);
and U3846 (N_3846,In_2051,In_2910);
and U3847 (N_3847,In_2685,In_2213);
or U3848 (N_3848,In_496,In_2635);
nor U3849 (N_3849,In_2019,In_119);
nand U3850 (N_3850,In_68,In_2119);
nand U3851 (N_3851,In_512,In_2135);
nand U3852 (N_3852,In_2890,In_2769);
nand U3853 (N_3853,In_1147,In_661);
xnor U3854 (N_3854,In_2163,In_1645);
and U3855 (N_3855,In_78,In_1633);
nor U3856 (N_3856,In_1315,In_1451);
nor U3857 (N_3857,In_2266,In_2669);
nand U3858 (N_3858,In_1426,In_1196);
nand U3859 (N_3859,In_2471,In_1218);
or U3860 (N_3860,In_2699,In_269);
nand U3861 (N_3861,In_1802,In_1435);
nor U3862 (N_3862,In_636,In_1726);
and U3863 (N_3863,In_225,In_1790);
or U3864 (N_3864,In_2113,In_350);
nand U3865 (N_3865,In_1211,In_922);
nor U3866 (N_3866,In_1280,In_2299);
and U3867 (N_3867,In_1044,In_217);
or U3868 (N_3868,In_1378,In_1515);
and U3869 (N_3869,In_1458,In_342);
or U3870 (N_3870,In_792,In_484);
and U3871 (N_3871,In_612,In_606);
and U3872 (N_3872,In_1790,In_1441);
or U3873 (N_3873,In_2504,In_2211);
nor U3874 (N_3874,In_2714,In_35);
xnor U3875 (N_3875,In_2278,In_1069);
and U3876 (N_3876,In_679,In_835);
nand U3877 (N_3877,In_1116,In_2496);
or U3878 (N_3878,In_2863,In_1930);
and U3879 (N_3879,In_954,In_2694);
nor U3880 (N_3880,In_1026,In_2085);
nor U3881 (N_3881,In_2253,In_1927);
nand U3882 (N_3882,In_940,In_1378);
and U3883 (N_3883,In_2051,In_1550);
and U3884 (N_3884,In_361,In_711);
or U3885 (N_3885,In_1898,In_1801);
nand U3886 (N_3886,In_1007,In_356);
or U3887 (N_3887,In_952,In_2444);
nand U3888 (N_3888,In_2077,In_2360);
and U3889 (N_3889,In_2928,In_434);
nand U3890 (N_3890,In_2417,In_2639);
nor U3891 (N_3891,In_2746,In_906);
and U3892 (N_3892,In_2884,In_2235);
or U3893 (N_3893,In_2372,In_1101);
nand U3894 (N_3894,In_609,In_2134);
xnor U3895 (N_3895,In_765,In_475);
nand U3896 (N_3896,In_476,In_1558);
nor U3897 (N_3897,In_1087,In_18);
or U3898 (N_3898,In_1971,In_1354);
nand U3899 (N_3899,In_837,In_2450);
nor U3900 (N_3900,In_726,In_1783);
nand U3901 (N_3901,In_1958,In_380);
nand U3902 (N_3902,In_407,In_2049);
or U3903 (N_3903,In_61,In_2505);
xnor U3904 (N_3904,In_1621,In_1103);
and U3905 (N_3905,In_913,In_2914);
nor U3906 (N_3906,In_2197,In_1864);
or U3907 (N_3907,In_1061,In_1799);
and U3908 (N_3908,In_733,In_1095);
nor U3909 (N_3909,In_1067,In_178);
nor U3910 (N_3910,In_741,In_300);
or U3911 (N_3911,In_152,In_1494);
nand U3912 (N_3912,In_281,In_1446);
nor U3913 (N_3913,In_1723,In_189);
nor U3914 (N_3914,In_2354,In_869);
and U3915 (N_3915,In_2124,In_177);
nand U3916 (N_3916,In_147,In_1091);
and U3917 (N_3917,In_1502,In_963);
and U3918 (N_3918,In_1504,In_2563);
and U3919 (N_3919,In_2715,In_826);
and U3920 (N_3920,In_232,In_89);
nor U3921 (N_3921,In_2927,In_2404);
and U3922 (N_3922,In_2146,In_2245);
or U3923 (N_3923,In_2421,In_2212);
or U3924 (N_3924,In_709,In_2073);
nand U3925 (N_3925,In_1857,In_2094);
and U3926 (N_3926,In_2697,In_1105);
or U3927 (N_3927,In_1628,In_1545);
and U3928 (N_3928,In_193,In_1461);
nand U3929 (N_3929,In_501,In_1081);
nand U3930 (N_3930,In_99,In_1726);
and U3931 (N_3931,In_1157,In_307);
or U3932 (N_3932,In_30,In_1635);
nand U3933 (N_3933,In_2630,In_466);
or U3934 (N_3934,In_240,In_378);
or U3935 (N_3935,In_2362,In_774);
nand U3936 (N_3936,In_551,In_658);
nand U3937 (N_3937,In_2599,In_584);
nand U3938 (N_3938,In_421,In_1289);
nor U3939 (N_3939,In_2695,In_653);
and U3940 (N_3940,In_1662,In_1765);
nand U3941 (N_3941,In_880,In_351);
or U3942 (N_3942,In_2237,In_2815);
and U3943 (N_3943,In_2635,In_237);
nor U3944 (N_3944,In_2509,In_2933);
and U3945 (N_3945,In_1106,In_2314);
and U3946 (N_3946,In_425,In_2749);
and U3947 (N_3947,In_2194,In_1660);
and U3948 (N_3948,In_1186,In_865);
nand U3949 (N_3949,In_2368,In_797);
nor U3950 (N_3950,In_331,In_465);
nor U3951 (N_3951,In_1698,In_167);
or U3952 (N_3952,In_837,In_1008);
and U3953 (N_3953,In_2668,In_282);
and U3954 (N_3954,In_822,In_198);
or U3955 (N_3955,In_724,In_1416);
and U3956 (N_3956,In_740,In_2077);
and U3957 (N_3957,In_1853,In_887);
nor U3958 (N_3958,In_1269,In_449);
nor U3959 (N_3959,In_2622,In_1197);
and U3960 (N_3960,In_721,In_2875);
nor U3961 (N_3961,In_384,In_67);
nand U3962 (N_3962,In_1920,In_2487);
nor U3963 (N_3963,In_1017,In_416);
nand U3964 (N_3964,In_827,In_426);
and U3965 (N_3965,In_209,In_992);
nand U3966 (N_3966,In_1286,In_1818);
nor U3967 (N_3967,In_2151,In_2683);
nand U3968 (N_3968,In_1834,In_2986);
and U3969 (N_3969,In_2878,In_420);
nor U3970 (N_3970,In_2516,In_98);
and U3971 (N_3971,In_2574,In_1508);
nand U3972 (N_3972,In_1945,In_1450);
nand U3973 (N_3973,In_1173,In_913);
nand U3974 (N_3974,In_1431,In_2831);
nor U3975 (N_3975,In_1511,In_1343);
nor U3976 (N_3976,In_1207,In_2104);
nand U3977 (N_3977,In_1336,In_2065);
and U3978 (N_3978,In_1689,In_1268);
or U3979 (N_3979,In_2002,In_2631);
nor U3980 (N_3980,In_2359,In_2242);
or U3981 (N_3981,In_361,In_2120);
nand U3982 (N_3982,In_1210,In_1748);
nor U3983 (N_3983,In_2878,In_2853);
nor U3984 (N_3984,In_1806,In_1983);
and U3985 (N_3985,In_438,In_812);
nand U3986 (N_3986,In_2488,In_1026);
or U3987 (N_3987,In_2250,In_754);
and U3988 (N_3988,In_960,In_1022);
nand U3989 (N_3989,In_1937,In_2706);
and U3990 (N_3990,In_2582,In_2196);
nand U3991 (N_3991,In_2410,In_1554);
nand U3992 (N_3992,In_2705,In_48);
or U3993 (N_3993,In_2910,In_627);
nor U3994 (N_3994,In_931,In_2608);
or U3995 (N_3995,In_2994,In_968);
or U3996 (N_3996,In_2885,In_454);
or U3997 (N_3997,In_1207,In_533);
nor U3998 (N_3998,In_2679,In_2413);
nand U3999 (N_3999,In_1681,In_2241);
nor U4000 (N_4000,In_2705,In_1671);
nand U4001 (N_4001,In_1455,In_2422);
nor U4002 (N_4002,In_1705,In_1357);
nor U4003 (N_4003,In_2549,In_2880);
or U4004 (N_4004,In_1242,In_2222);
and U4005 (N_4005,In_1122,In_377);
nor U4006 (N_4006,In_520,In_743);
nor U4007 (N_4007,In_2275,In_532);
nor U4008 (N_4008,In_377,In_1885);
nor U4009 (N_4009,In_1134,In_1348);
nand U4010 (N_4010,In_2348,In_2301);
nor U4011 (N_4011,In_2832,In_1144);
and U4012 (N_4012,In_1785,In_2410);
nand U4013 (N_4013,In_2517,In_1043);
or U4014 (N_4014,In_1893,In_1785);
and U4015 (N_4015,In_1957,In_1211);
nor U4016 (N_4016,In_1073,In_851);
nand U4017 (N_4017,In_48,In_856);
or U4018 (N_4018,In_1381,In_1552);
and U4019 (N_4019,In_1099,In_1738);
and U4020 (N_4020,In_523,In_992);
nand U4021 (N_4021,In_615,In_226);
and U4022 (N_4022,In_1591,In_2279);
nand U4023 (N_4023,In_2066,In_2264);
or U4024 (N_4024,In_1758,In_1948);
and U4025 (N_4025,In_418,In_1648);
nor U4026 (N_4026,In_410,In_1579);
and U4027 (N_4027,In_2698,In_2431);
and U4028 (N_4028,In_213,In_2298);
or U4029 (N_4029,In_680,In_1198);
and U4030 (N_4030,In_921,In_2650);
and U4031 (N_4031,In_172,In_1036);
or U4032 (N_4032,In_2841,In_2934);
nor U4033 (N_4033,In_2014,In_2420);
nor U4034 (N_4034,In_514,In_973);
and U4035 (N_4035,In_1412,In_1233);
nand U4036 (N_4036,In_2090,In_1021);
nor U4037 (N_4037,In_1112,In_870);
nor U4038 (N_4038,In_2517,In_2623);
nand U4039 (N_4039,In_1452,In_517);
nor U4040 (N_4040,In_1790,In_151);
nand U4041 (N_4041,In_1298,In_263);
nand U4042 (N_4042,In_1864,In_2402);
nand U4043 (N_4043,In_1044,In_975);
nand U4044 (N_4044,In_1274,In_897);
and U4045 (N_4045,In_2067,In_2221);
and U4046 (N_4046,In_1059,In_1127);
nor U4047 (N_4047,In_665,In_3);
or U4048 (N_4048,In_617,In_1310);
and U4049 (N_4049,In_391,In_2222);
nand U4050 (N_4050,In_1830,In_712);
and U4051 (N_4051,In_490,In_1393);
nor U4052 (N_4052,In_165,In_1233);
nor U4053 (N_4053,In_1550,In_1572);
or U4054 (N_4054,In_1112,In_807);
or U4055 (N_4055,In_1568,In_2702);
and U4056 (N_4056,In_1551,In_2138);
or U4057 (N_4057,In_63,In_2786);
or U4058 (N_4058,In_2866,In_1253);
nor U4059 (N_4059,In_2989,In_2551);
nor U4060 (N_4060,In_1662,In_1568);
or U4061 (N_4061,In_898,In_2107);
xnor U4062 (N_4062,In_1183,In_2496);
nor U4063 (N_4063,In_2013,In_2110);
or U4064 (N_4064,In_46,In_1850);
or U4065 (N_4065,In_902,In_2813);
or U4066 (N_4066,In_659,In_794);
nor U4067 (N_4067,In_54,In_2011);
or U4068 (N_4068,In_1810,In_680);
or U4069 (N_4069,In_650,In_216);
nor U4070 (N_4070,In_344,In_2197);
nand U4071 (N_4071,In_2821,In_2281);
nor U4072 (N_4072,In_442,In_1777);
nor U4073 (N_4073,In_563,In_2946);
or U4074 (N_4074,In_1727,In_501);
nor U4075 (N_4075,In_568,In_1494);
nor U4076 (N_4076,In_2819,In_1591);
or U4077 (N_4077,In_2604,In_253);
and U4078 (N_4078,In_121,In_412);
nor U4079 (N_4079,In_776,In_2565);
or U4080 (N_4080,In_2946,In_2390);
nor U4081 (N_4081,In_797,In_1466);
and U4082 (N_4082,In_2874,In_1305);
nor U4083 (N_4083,In_1441,In_1423);
or U4084 (N_4084,In_2899,In_1249);
and U4085 (N_4085,In_2256,In_1024);
nor U4086 (N_4086,In_2755,In_2600);
nor U4087 (N_4087,In_787,In_683);
and U4088 (N_4088,In_792,In_2378);
nand U4089 (N_4089,In_500,In_1495);
nand U4090 (N_4090,In_1899,In_1825);
or U4091 (N_4091,In_2577,In_1009);
nand U4092 (N_4092,In_898,In_2838);
or U4093 (N_4093,In_1033,In_590);
or U4094 (N_4094,In_2434,In_1476);
and U4095 (N_4095,In_1448,In_2364);
or U4096 (N_4096,In_2998,In_1218);
nand U4097 (N_4097,In_2642,In_2809);
and U4098 (N_4098,In_1598,In_695);
nand U4099 (N_4099,In_2822,In_2804);
nand U4100 (N_4100,In_2003,In_155);
and U4101 (N_4101,In_2079,In_699);
nand U4102 (N_4102,In_2584,In_796);
or U4103 (N_4103,In_274,In_1597);
nor U4104 (N_4104,In_1749,In_484);
nor U4105 (N_4105,In_1444,In_1721);
or U4106 (N_4106,In_2793,In_906);
and U4107 (N_4107,In_1518,In_1978);
and U4108 (N_4108,In_1537,In_1717);
nor U4109 (N_4109,In_665,In_881);
nor U4110 (N_4110,In_2621,In_2709);
or U4111 (N_4111,In_2000,In_2931);
or U4112 (N_4112,In_2469,In_811);
or U4113 (N_4113,In_2595,In_21);
or U4114 (N_4114,In_172,In_1656);
or U4115 (N_4115,In_1186,In_2086);
and U4116 (N_4116,In_217,In_640);
nand U4117 (N_4117,In_1708,In_997);
or U4118 (N_4118,In_877,In_1053);
nor U4119 (N_4119,In_2057,In_1887);
nand U4120 (N_4120,In_2832,In_2901);
nor U4121 (N_4121,In_176,In_244);
or U4122 (N_4122,In_1279,In_267);
or U4123 (N_4123,In_205,In_1972);
nor U4124 (N_4124,In_875,In_1632);
and U4125 (N_4125,In_1147,In_2941);
nand U4126 (N_4126,In_945,In_1899);
nand U4127 (N_4127,In_795,In_210);
and U4128 (N_4128,In_120,In_2143);
nand U4129 (N_4129,In_225,In_1691);
or U4130 (N_4130,In_2607,In_2667);
nand U4131 (N_4131,In_2756,In_712);
or U4132 (N_4132,In_246,In_1598);
or U4133 (N_4133,In_2143,In_1352);
nand U4134 (N_4134,In_1216,In_260);
and U4135 (N_4135,In_1903,In_2686);
or U4136 (N_4136,In_1033,In_2369);
nand U4137 (N_4137,In_1384,In_1071);
and U4138 (N_4138,In_2293,In_651);
or U4139 (N_4139,In_1318,In_665);
or U4140 (N_4140,In_2844,In_1840);
nor U4141 (N_4141,In_2987,In_1383);
nand U4142 (N_4142,In_56,In_2487);
and U4143 (N_4143,In_2362,In_2348);
nand U4144 (N_4144,In_1095,In_76);
nor U4145 (N_4145,In_1275,In_1087);
and U4146 (N_4146,In_2754,In_1761);
or U4147 (N_4147,In_2941,In_769);
or U4148 (N_4148,In_1816,In_2930);
and U4149 (N_4149,In_429,In_2152);
nor U4150 (N_4150,In_2406,In_399);
or U4151 (N_4151,In_1723,In_1414);
nor U4152 (N_4152,In_2844,In_2458);
nand U4153 (N_4153,In_2787,In_2781);
xnor U4154 (N_4154,In_625,In_1267);
or U4155 (N_4155,In_1483,In_404);
and U4156 (N_4156,In_2628,In_215);
nand U4157 (N_4157,In_744,In_1398);
nand U4158 (N_4158,In_1057,In_868);
or U4159 (N_4159,In_1319,In_1206);
nand U4160 (N_4160,In_2632,In_2898);
and U4161 (N_4161,In_1514,In_1050);
and U4162 (N_4162,In_1508,In_1756);
or U4163 (N_4163,In_2084,In_1939);
nand U4164 (N_4164,In_1407,In_2387);
or U4165 (N_4165,In_897,In_995);
or U4166 (N_4166,In_2957,In_440);
nand U4167 (N_4167,In_462,In_2783);
nor U4168 (N_4168,In_2558,In_2900);
and U4169 (N_4169,In_132,In_150);
nand U4170 (N_4170,In_2925,In_1250);
or U4171 (N_4171,In_1280,In_2007);
nand U4172 (N_4172,In_2549,In_691);
nand U4173 (N_4173,In_744,In_1519);
or U4174 (N_4174,In_1486,In_645);
nor U4175 (N_4175,In_779,In_359);
nand U4176 (N_4176,In_81,In_1334);
nor U4177 (N_4177,In_372,In_2679);
nand U4178 (N_4178,In_232,In_480);
and U4179 (N_4179,In_2976,In_447);
nand U4180 (N_4180,In_638,In_2634);
nand U4181 (N_4181,In_1366,In_597);
nand U4182 (N_4182,In_2854,In_1954);
nand U4183 (N_4183,In_372,In_2543);
or U4184 (N_4184,In_1195,In_2245);
nand U4185 (N_4185,In_356,In_2330);
nand U4186 (N_4186,In_2723,In_25);
nor U4187 (N_4187,In_2378,In_1775);
or U4188 (N_4188,In_2058,In_2733);
nand U4189 (N_4189,In_1627,In_786);
nand U4190 (N_4190,In_2662,In_1335);
and U4191 (N_4191,In_1958,In_1517);
and U4192 (N_4192,In_186,In_2870);
nand U4193 (N_4193,In_2430,In_1471);
or U4194 (N_4194,In_1332,In_1929);
nand U4195 (N_4195,In_812,In_677);
nand U4196 (N_4196,In_1374,In_429);
nor U4197 (N_4197,In_620,In_176);
or U4198 (N_4198,In_2689,In_980);
nand U4199 (N_4199,In_718,In_1983);
nand U4200 (N_4200,In_1189,In_1516);
xor U4201 (N_4201,In_2492,In_1943);
nand U4202 (N_4202,In_857,In_1511);
nor U4203 (N_4203,In_1665,In_1709);
nor U4204 (N_4204,In_2490,In_599);
and U4205 (N_4205,In_1864,In_1852);
nand U4206 (N_4206,In_1174,In_627);
or U4207 (N_4207,In_675,In_2314);
or U4208 (N_4208,In_28,In_673);
nor U4209 (N_4209,In_2416,In_2487);
and U4210 (N_4210,In_964,In_2240);
nor U4211 (N_4211,In_7,In_2837);
nand U4212 (N_4212,In_2185,In_1155);
nand U4213 (N_4213,In_1308,In_653);
or U4214 (N_4214,In_1352,In_47);
nand U4215 (N_4215,In_891,In_1278);
nor U4216 (N_4216,In_131,In_1981);
and U4217 (N_4217,In_2603,In_87);
and U4218 (N_4218,In_212,In_2096);
nor U4219 (N_4219,In_2678,In_486);
or U4220 (N_4220,In_1750,In_1505);
nor U4221 (N_4221,In_2144,In_2328);
and U4222 (N_4222,In_2981,In_1228);
nand U4223 (N_4223,In_335,In_921);
nand U4224 (N_4224,In_2758,In_416);
nor U4225 (N_4225,In_597,In_1585);
nand U4226 (N_4226,In_2621,In_1735);
or U4227 (N_4227,In_2464,In_1861);
and U4228 (N_4228,In_108,In_855);
xnor U4229 (N_4229,In_2159,In_1433);
nor U4230 (N_4230,In_64,In_86);
or U4231 (N_4231,In_495,In_764);
nor U4232 (N_4232,In_899,In_1469);
xnor U4233 (N_4233,In_192,In_223);
nand U4234 (N_4234,In_2750,In_1721);
nor U4235 (N_4235,In_2206,In_24);
and U4236 (N_4236,In_828,In_136);
nand U4237 (N_4237,In_1541,In_1117);
nand U4238 (N_4238,In_2631,In_2950);
nor U4239 (N_4239,In_401,In_2282);
or U4240 (N_4240,In_1877,In_407);
and U4241 (N_4241,In_964,In_2673);
and U4242 (N_4242,In_79,In_362);
and U4243 (N_4243,In_1496,In_358);
nand U4244 (N_4244,In_790,In_1281);
nand U4245 (N_4245,In_168,In_1214);
nor U4246 (N_4246,In_1318,In_1325);
nor U4247 (N_4247,In_1198,In_2031);
and U4248 (N_4248,In_440,In_937);
nand U4249 (N_4249,In_102,In_2540);
nor U4250 (N_4250,In_1799,In_1422);
and U4251 (N_4251,In_2159,In_2324);
nand U4252 (N_4252,In_1840,In_2979);
or U4253 (N_4253,In_1868,In_2201);
nor U4254 (N_4254,In_798,In_1191);
and U4255 (N_4255,In_1904,In_2545);
nor U4256 (N_4256,In_2982,In_176);
and U4257 (N_4257,In_723,In_1850);
or U4258 (N_4258,In_555,In_2939);
nor U4259 (N_4259,In_2929,In_573);
nor U4260 (N_4260,In_2535,In_367);
nand U4261 (N_4261,In_2928,In_2939);
or U4262 (N_4262,In_1478,In_1452);
or U4263 (N_4263,In_2496,In_391);
nor U4264 (N_4264,In_1780,In_2894);
and U4265 (N_4265,In_2378,In_2114);
and U4266 (N_4266,In_2131,In_1939);
or U4267 (N_4267,In_1887,In_2466);
or U4268 (N_4268,In_1647,In_2027);
nor U4269 (N_4269,In_1572,In_913);
or U4270 (N_4270,In_1215,In_2209);
nand U4271 (N_4271,In_67,In_1587);
and U4272 (N_4272,In_2108,In_29);
nand U4273 (N_4273,In_2627,In_105);
nor U4274 (N_4274,In_2627,In_1870);
nand U4275 (N_4275,In_85,In_461);
and U4276 (N_4276,In_710,In_513);
xor U4277 (N_4277,In_515,In_690);
or U4278 (N_4278,In_1443,In_2351);
nor U4279 (N_4279,In_249,In_1063);
nand U4280 (N_4280,In_1391,In_1470);
or U4281 (N_4281,In_1373,In_1990);
and U4282 (N_4282,In_2993,In_1218);
nor U4283 (N_4283,In_2929,In_2405);
or U4284 (N_4284,In_1285,In_2947);
nor U4285 (N_4285,In_406,In_33);
nor U4286 (N_4286,In_802,In_138);
or U4287 (N_4287,In_2607,In_2597);
nor U4288 (N_4288,In_751,In_1353);
or U4289 (N_4289,In_1479,In_2850);
nor U4290 (N_4290,In_963,In_2228);
and U4291 (N_4291,In_1292,In_483);
or U4292 (N_4292,In_2383,In_2218);
or U4293 (N_4293,In_201,In_2710);
or U4294 (N_4294,In_733,In_656);
nor U4295 (N_4295,In_1964,In_279);
or U4296 (N_4296,In_2563,In_2175);
or U4297 (N_4297,In_2767,In_1024);
nand U4298 (N_4298,In_1456,In_802);
nor U4299 (N_4299,In_293,In_277);
nor U4300 (N_4300,In_2611,In_2714);
nor U4301 (N_4301,In_2386,In_437);
nand U4302 (N_4302,In_1757,In_256);
and U4303 (N_4303,In_599,In_1795);
nor U4304 (N_4304,In_385,In_2742);
or U4305 (N_4305,In_2417,In_1121);
nor U4306 (N_4306,In_2723,In_345);
nand U4307 (N_4307,In_522,In_2985);
and U4308 (N_4308,In_159,In_2416);
nor U4309 (N_4309,In_2308,In_1913);
nand U4310 (N_4310,In_836,In_1237);
and U4311 (N_4311,In_1824,In_81);
nand U4312 (N_4312,In_2692,In_1279);
or U4313 (N_4313,In_1636,In_2625);
and U4314 (N_4314,In_529,In_1140);
or U4315 (N_4315,In_1631,In_1);
xor U4316 (N_4316,In_292,In_282);
or U4317 (N_4317,In_2231,In_2644);
or U4318 (N_4318,In_2238,In_170);
nor U4319 (N_4319,In_2804,In_1812);
nor U4320 (N_4320,In_2664,In_2961);
xor U4321 (N_4321,In_2057,In_1897);
or U4322 (N_4322,In_1240,In_800);
and U4323 (N_4323,In_1357,In_1689);
or U4324 (N_4324,In_1809,In_867);
or U4325 (N_4325,In_286,In_2401);
and U4326 (N_4326,In_1965,In_2414);
nor U4327 (N_4327,In_1255,In_2263);
and U4328 (N_4328,In_1174,In_1690);
nand U4329 (N_4329,In_2923,In_1023);
and U4330 (N_4330,In_1026,In_1371);
nand U4331 (N_4331,In_1547,In_866);
and U4332 (N_4332,In_151,In_664);
nand U4333 (N_4333,In_2655,In_1182);
nand U4334 (N_4334,In_44,In_481);
and U4335 (N_4335,In_2121,In_538);
and U4336 (N_4336,In_2970,In_1605);
xnor U4337 (N_4337,In_2676,In_1209);
and U4338 (N_4338,In_816,In_2312);
or U4339 (N_4339,In_1799,In_1744);
or U4340 (N_4340,In_1555,In_829);
nor U4341 (N_4341,In_1955,In_2898);
nand U4342 (N_4342,In_932,In_573);
nand U4343 (N_4343,In_2103,In_226);
and U4344 (N_4344,In_2831,In_1788);
and U4345 (N_4345,In_1657,In_488);
and U4346 (N_4346,In_2908,In_2653);
nand U4347 (N_4347,In_920,In_1592);
and U4348 (N_4348,In_1039,In_1576);
and U4349 (N_4349,In_602,In_658);
and U4350 (N_4350,In_1266,In_2916);
nor U4351 (N_4351,In_2719,In_1787);
nor U4352 (N_4352,In_1115,In_238);
or U4353 (N_4353,In_954,In_1122);
or U4354 (N_4354,In_2991,In_1434);
nor U4355 (N_4355,In_2528,In_2517);
nand U4356 (N_4356,In_431,In_1981);
or U4357 (N_4357,In_2724,In_461);
nand U4358 (N_4358,In_2375,In_506);
xor U4359 (N_4359,In_149,In_2677);
nand U4360 (N_4360,In_1682,In_1572);
or U4361 (N_4361,In_1760,In_98);
nor U4362 (N_4362,In_2620,In_2717);
or U4363 (N_4363,In_3,In_971);
nor U4364 (N_4364,In_2158,In_2979);
nor U4365 (N_4365,In_1847,In_2741);
and U4366 (N_4366,In_1677,In_979);
nor U4367 (N_4367,In_541,In_1066);
or U4368 (N_4368,In_816,In_2847);
nor U4369 (N_4369,In_2395,In_1195);
and U4370 (N_4370,In_2248,In_624);
nand U4371 (N_4371,In_2985,In_1581);
and U4372 (N_4372,In_959,In_2839);
nand U4373 (N_4373,In_1372,In_462);
nor U4374 (N_4374,In_2645,In_8);
and U4375 (N_4375,In_325,In_767);
and U4376 (N_4376,In_527,In_1748);
and U4377 (N_4377,In_1646,In_1650);
and U4378 (N_4378,In_1484,In_2906);
nand U4379 (N_4379,In_1913,In_2354);
nand U4380 (N_4380,In_1867,In_1956);
or U4381 (N_4381,In_2561,In_2374);
and U4382 (N_4382,In_2256,In_2864);
nand U4383 (N_4383,In_2291,In_1535);
or U4384 (N_4384,In_2007,In_135);
nor U4385 (N_4385,In_2714,In_2104);
or U4386 (N_4386,In_108,In_2110);
nand U4387 (N_4387,In_1113,In_793);
nor U4388 (N_4388,In_138,In_1852);
and U4389 (N_4389,In_2610,In_1416);
or U4390 (N_4390,In_2091,In_1362);
and U4391 (N_4391,In_835,In_2715);
and U4392 (N_4392,In_2656,In_334);
nand U4393 (N_4393,In_2489,In_768);
or U4394 (N_4394,In_2127,In_208);
and U4395 (N_4395,In_923,In_1658);
nand U4396 (N_4396,In_868,In_909);
or U4397 (N_4397,In_212,In_2221);
or U4398 (N_4398,In_2210,In_2321);
nand U4399 (N_4399,In_2299,In_310);
nor U4400 (N_4400,In_1350,In_1638);
nand U4401 (N_4401,In_382,In_176);
or U4402 (N_4402,In_717,In_664);
and U4403 (N_4403,In_2037,In_1788);
nor U4404 (N_4404,In_1420,In_1075);
or U4405 (N_4405,In_1510,In_513);
nand U4406 (N_4406,In_40,In_2532);
nand U4407 (N_4407,In_1503,In_2253);
nand U4408 (N_4408,In_2518,In_13);
or U4409 (N_4409,In_214,In_2189);
and U4410 (N_4410,In_399,In_266);
nor U4411 (N_4411,In_717,In_966);
nor U4412 (N_4412,In_2901,In_1490);
and U4413 (N_4413,In_420,In_2672);
nand U4414 (N_4414,In_1566,In_2455);
and U4415 (N_4415,In_393,In_1405);
and U4416 (N_4416,In_2143,In_36);
nor U4417 (N_4417,In_143,In_25);
or U4418 (N_4418,In_2621,In_2770);
nor U4419 (N_4419,In_2562,In_2634);
nand U4420 (N_4420,In_1521,In_791);
or U4421 (N_4421,In_2066,In_2061);
nor U4422 (N_4422,In_1719,In_1496);
or U4423 (N_4423,In_2497,In_543);
nor U4424 (N_4424,In_466,In_897);
nor U4425 (N_4425,In_2488,In_1824);
nor U4426 (N_4426,In_2425,In_1533);
nand U4427 (N_4427,In_776,In_1967);
nor U4428 (N_4428,In_1866,In_2697);
or U4429 (N_4429,In_423,In_1160);
and U4430 (N_4430,In_926,In_1818);
nand U4431 (N_4431,In_2129,In_2065);
nand U4432 (N_4432,In_1197,In_1274);
nand U4433 (N_4433,In_727,In_2300);
or U4434 (N_4434,In_1586,In_202);
and U4435 (N_4435,In_132,In_858);
and U4436 (N_4436,In_1399,In_2046);
and U4437 (N_4437,In_1362,In_2788);
nor U4438 (N_4438,In_753,In_879);
nor U4439 (N_4439,In_580,In_1910);
and U4440 (N_4440,In_79,In_2041);
nor U4441 (N_4441,In_1200,In_1551);
nand U4442 (N_4442,In_409,In_175);
nor U4443 (N_4443,In_1147,In_2988);
nand U4444 (N_4444,In_392,In_1339);
nand U4445 (N_4445,In_1082,In_1707);
nor U4446 (N_4446,In_1536,In_75);
nand U4447 (N_4447,In_2808,In_922);
or U4448 (N_4448,In_745,In_2364);
or U4449 (N_4449,In_2452,In_1090);
and U4450 (N_4450,In_2807,In_2328);
and U4451 (N_4451,In_1161,In_1271);
nor U4452 (N_4452,In_436,In_1149);
xor U4453 (N_4453,In_469,In_1189);
and U4454 (N_4454,In_1606,In_482);
or U4455 (N_4455,In_2573,In_1803);
nor U4456 (N_4456,In_54,In_1222);
or U4457 (N_4457,In_491,In_1228);
or U4458 (N_4458,In_2386,In_2276);
and U4459 (N_4459,In_2774,In_2708);
nand U4460 (N_4460,In_2446,In_2957);
or U4461 (N_4461,In_2501,In_1028);
nand U4462 (N_4462,In_578,In_179);
xnor U4463 (N_4463,In_726,In_2981);
or U4464 (N_4464,In_2387,In_2237);
or U4465 (N_4465,In_2178,In_579);
nand U4466 (N_4466,In_1319,In_239);
and U4467 (N_4467,In_2681,In_2309);
nor U4468 (N_4468,In_1985,In_2382);
and U4469 (N_4469,In_2146,In_2206);
nand U4470 (N_4470,In_2873,In_2968);
or U4471 (N_4471,In_1328,In_2440);
nor U4472 (N_4472,In_662,In_2436);
and U4473 (N_4473,In_1640,In_1029);
or U4474 (N_4474,In_2513,In_1837);
nand U4475 (N_4475,In_2717,In_1033);
and U4476 (N_4476,In_556,In_1749);
nand U4477 (N_4477,In_2772,In_1100);
nand U4478 (N_4478,In_2533,In_486);
or U4479 (N_4479,In_1541,In_2453);
and U4480 (N_4480,In_186,In_1069);
and U4481 (N_4481,In_237,In_2209);
or U4482 (N_4482,In_1824,In_2230);
nor U4483 (N_4483,In_833,In_2527);
and U4484 (N_4484,In_2409,In_897);
and U4485 (N_4485,In_1338,In_1291);
nand U4486 (N_4486,In_1276,In_1572);
nor U4487 (N_4487,In_845,In_65);
or U4488 (N_4488,In_1776,In_120);
nor U4489 (N_4489,In_707,In_1145);
and U4490 (N_4490,In_1856,In_1980);
nand U4491 (N_4491,In_267,In_2740);
nor U4492 (N_4492,In_1904,In_282);
nor U4493 (N_4493,In_328,In_46);
and U4494 (N_4494,In_778,In_1456);
or U4495 (N_4495,In_684,In_1907);
and U4496 (N_4496,In_1921,In_1923);
nor U4497 (N_4497,In_2830,In_1998);
and U4498 (N_4498,In_2133,In_1747);
nor U4499 (N_4499,In_2700,In_2268);
or U4500 (N_4500,In_787,In_300);
and U4501 (N_4501,In_929,In_2309);
nor U4502 (N_4502,In_107,In_179);
or U4503 (N_4503,In_2781,In_2135);
nand U4504 (N_4504,In_1892,In_2338);
nor U4505 (N_4505,In_400,In_1881);
or U4506 (N_4506,In_398,In_2062);
or U4507 (N_4507,In_798,In_1439);
nor U4508 (N_4508,In_803,In_1463);
or U4509 (N_4509,In_2443,In_2609);
nand U4510 (N_4510,In_1522,In_2328);
and U4511 (N_4511,In_415,In_23);
nand U4512 (N_4512,In_2053,In_2913);
nor U4513 (N_4513,In_1918,In_1456);
and U4514 (N_4514,In_2285,In_2923);
nand U4515 (N_4515,In_867,In_2710);
or U4516 (N_4516,In_1657,In_2380);
and U4517 (N_4517,In_136,In_186);
nand U4518 (N_4518,In_2163,In_142);
or U4519 (N_4519,In_1717,In_1627);
nand U4520 (N_4520,In_2945,In_1398);
nand U4521 (N_4521,In_268,In_1233);
nand U4522 (N_4522,In_557,In_2948);
or U4523 (N_4523,In_590,In_486);
or U4524 (N_4524,In_1184,In_1976);
and U4525 (N_4525,In_2790,In_611);
and U4526 (N_4526,In_494,In_146);
nor U4527 (N_4527,In_1027,In_2735);
nor U4528 (N_4528,In_615,In_1891);
nand U4529 (N_4529,In_2473,In_1792);
nand U4530 (N_4530,In_16,In_1366);
or U4531 (N_4531,In_1955,In_1507);
nand U4532 (N_4532,In_1327,In_1024);
or U4533 (N_4533,In_655,In_2466);
and U4534 (N_4534,In_1634,In_813);
and U4535 (N_4535,In_987,In_507);
nand U4536 (N_4536,In_2523,In_1749);
or U4537 (N_4537,In_2141,In_234);
nand U4538 (N_4538,In_2064,In_768);
nand U4539 (N_4539,In_2260,In_890);
and U4540 (N_4540,In_2202,In_780);
nor U4541 (N_4541,In_421,In_2853);
or U4542 (N_4542,In_122,In_821);
nor U4543 (N_4543,In_1151,In_2193);
and U4544 (N_4544,In_1424,In_74);
and U4545 (N_4545,In_658,In_2562);
or U4546 (N_4546,In_636,In_2334);
or U4547 (N_4547,In_2062,In_2874);
nor U4548 (N_4548,In_378,In_2287);
nand U4549 (N_4549,In_2622,In_1546);
nand U4550 (N_4550,In_1601,In_1876);
nor U4551 (N_4551,In_123,In_1652);
nand U4552 (N_4552,In_2521,In_1794);
nor U4553 (N_4553,In_1237,In_238);
and U4554 (N_4554,In_711,In_2014);
nand U4555 (N_4555,In_2660,In_146);
or U4556 (N_4556,In_2037,In_2076);
and U4557 (N_4557,In_2532,In_1990);
nand U4558 (N_4558,In_1677,In_1656);
nor U4559 (N_4559,In_2986,In_525);
nand U4560 (N_4560,In_841,In_2145);
nand U4561 (N_4561,In_1393,In_2106);
or U4562 (N_4562,In_2319,In_402);
and U4563 (N_4563,In_1284,In_1826);
nand U4564 (N_4564,In_866,In_1473);
xnor U4565 (N_4565,In_1752,In_671);
nand U4566 (N_4566,In_61,In_519);
or U4567 (N_4567,In_2133,In_1802);
nand U4568 (N_4568,In_2599,In_549);
and U4569 (N_4569,In_2862,In_63);
and U4570 (N_4570,In_2603,In_2552);
or U4571 (N_4571,In_2497,In_1178);
nor U4572 (N_4572,In_1347,In_871);
nor U4573 (N_4573,In_2129,In_1766);
nand U4574 (N_4574,In_1173,In_1604);
or U4575 (N_4575,In_1085,In_2800);
and U4576 (N_4576,In_1293,In_2433);
or U4577 (N_4577,In_1077,In_1982);
nor U4578 (N_4578,In_524,In_2368);
or U4579 (N_4579,In_1276,In_1665);
and U4580 (N_4580,In_2313,In_1652);
nand U4581 (N_4581,In_1472,In_2340);
and U4582 (N_4582,In_1525,In_2508);
or U4583 (N_4583,In_2151,In_1405);
nand U4584 (N_4584,In_88,In_1293);
or U4585 (N_4585,In_738,In_893);
nand U4586 (N_4586,In_1745,In_2396);
or U4587 (N_4587,In_1095,In_207);
nand U4588 (N_4588,In_865,In_759);
xnor U4589 (N_4589,In_1853,In_1729);
nand U4590 (N_4590,In_1096,In_2160);
xor U4591 (N_4591,In_1251,In_1520);
nand U4592 (N_4592,In_969,In_1534);
nand U4593 (N_4593,In_2731,In_2549);
nand U4594 (N_4594,In_1615,In_2258);
nor U4595 (N_4595,In_2527,In_1653);
and U4596 (N_4596,In_668,In_233);
nor U4597 (N_4597,In_930,In_1392);
and U4598 (N_4598,In_85,In_2041);
nand U4599 (N_4599,In_1441,In_1561);
and U4600 (N_4600,In_2361,In_1849);
or U4601 (N_4601,In_2547,In_1984);
and U4602 (N_4602,In_2621,In_1559);
nand U4603 (N_4603,In_2642,In_1602);
and U4604 (N_4604,In_856,In_770);
and U4605 (N_4605,In_1630,In_1306);
nor U4606 (N_4606,In_542,In_106);
nand U4607 (N_4607,In_2883,In_2976);
or U4608 (N_4608,In_2556,In_2070);
and U4609 (N_4609,In_93,In_2574);
nand U4610 (N_4610,In_1635,In_2850);
and U4611 (N_4611,In_2482,In_1491);
nor U4612 (N_4612,In_924,In_443);
nor U4613 (N_4613,In_2467,In_313);
nor U4614 (N_4614,In_2998,In_1112);
nor U4615 (N_4615,In_1451,In_586);
nor U4616 (N_4616,In_930,In_199);
and U4617 (N_4617,In_2497,In_1244);
nor U4618 (N_4618,In_2117,In_408);
nand U4619 (N_4619,In_2302,In_1143);
nand U4620 (N_4620,In_667,In_1660);
nor U4621 (N_4621,In_607,In_1912);
or U4622 (N_4622,In_527,In_952);
or U4623 (N_4623,In_1517,In_1872);
nor U4624 (N_4624,In_2397,In_2070);
and U4625 (N_4625,In_2945,In_175);
or U4626 (N_4626,In_2815,In_2890);
nor U4627 (N_4627,In_1570,In_301);
nand U4628 (N_4628,In_91,In_2958);
nor U4629 (N_4629,In_1946,In_835);
and U4630 (N_4630,In_1939,In_2644);
nand U4631 (N_4631,In_941,In_2680);
nor U4632 (N_4632,In_2734,In_2203);
nand U4633 (N_4633,In_2695,In_1941);
nor U4634 (N_4634,In_2242,In_2520);
nor U4635 (N_4635,In_1461,In_1533);
or U4636 (N_4636,In_2194,In_2808);
or U4637 (N_4637,In_1667,In_104);
and U4638 (N_4638,In_1898,In_848);
and U4639 (N_4639,In_2038,In_1103);
and U4640 (N_4640,In_920,In_1823);
or U4641 (N_4641,In_1317,In_2253);
and U4642 (N_4642,In_28,In_1702);
and U4643 (N_4643,In_671,In_1928);
nand U4644 (N_4644,In_1994,In_1262);
nor U4645 (N_4645,In_1697,In_906);
or U4646 (N_4646,In_1078,In_1435);
and U4647 (N_4647,In_1552,In_664);
and U4648 (N_4648,In_2050,In_1833);
or U4649 (N_4649,In_1932,In_2304);
nor U4650 (N_4650,In_2875,In_2460);
nor U4651 (N_4651,In_2978,In_1147);
or U4652 (N_4652,In_1045,In_375);
nor U4653 (N_4653,In_2923,In_1982);
and U4654 (N_4654,In_1695,In_1215);
or U4655 (N_4655,In_1383,In_647);
or U4656 (N_4656,In_1092,In_1152);
nand U4657 (N_4657,In_2651,In_2471);
or U4658 (N_4658,In_1541,In_1745);
and U4659 (N_4659,In_659,In_2946);
or U4660 (N_4660,In_1813,In_1432);
nor U4661 (N_4661,In_1352,In_1654);
or U4662 (N_4662,In_1514,In_1522);
nand U4663 (N_4663,In_185,In_487);
or U4664 (N_4664,In_134,In_1108);
nand U4665 (N_4665,In_2740,In_1076);
and U4666 (N_4666,In_2311,In_2469);
nor U4667 (N_4667,In_1820,In_2900);
nand U4668 (N_4668,In_2939,In_2305);
nand U4669 (N_4669,In_2337,In_430);
nand U4670 (N_4670,In_1484,In_822);
or U4671 (N_4671,In_2787,In_371);
nand U4672 (N_4672,In_1126,In_739);
nor U4673 (N_4673,In_1861,In_890);
xor U4674 (N_4674,In_1559,In_1709);
and U4675 (N_4675,In_772,In_1111);
or U4676 (N_4676,In_789,In_2184);
or U4677 (N_4677,In_2205,In_1514);
nor U4678 (N_4678,In_1958,In_2071);
nor U4679 (N_4679,In_1377,In_1941);
nand U4680 (N_4680,In_1939,In_2469);
nor U4681 (N_4681,In_2270,In_189);
nand U4682 (N_4682,In_2250,In_2840);
nor U4683 (N_4683,In_1380,In_1738);
nand U4684 (N_4684,In_1805,In_1042);
or U4685 (N_4685,In_2172,In_2341);
and U4686 (N_4686,In_270,In_2118);
or U4687 (N_4687,In_951,In_1251);
or U4688 (N_4688,In_1286,In_2263);
or U4689 (N_4689,In_2552,In_2786);
or U4690 (N_4690,In_2534,In_2633);
or U4691 (N_4691,In_229,In_2458);
or U4692 (N_4692,In_334,In_1643);
nor U4693 (N_4693,In_1156,In_32);
and U4694 (N_4694,In_1382,In_2690);
nand U4695 (N_4695,In_1948,In_1443);
or U4696 (N_4696,In_782,In_248);
nand U4697 (N_4697,In_1419,In_789);
nand U4698 (N_4698,In_2457,In_2859);
nand U4699 (N_4699,In_455,In_2411);
nand U4700 (N_4700,In_2782,In_929);
nand U4701 (N_4701,In_1291,In_1049);
nor U4702 (N_4702,In_1176,In_1149);
and U4703 (N_4703,In_2911,In_2248);
or U4704 (N_4704,In_1907,In_383);
nand U4705 (N_4705,In_1075,In_669);
nor U4706 (N_4706,In_1235,In_2807);
and U4707 (N_4707,In_683,In_1557);
nor U4708 (N_4708,In_1013,In_1425);
nand U4709 (N_4709,In_693,In_1248);
nand U4710 (N_4710,In_2084,In_1592);
nand U4711 (N_4711,In_867,In_72);
and U4712 (N_4712,In_898,In_2762);
nor U4713 (N_4713,In_1911,In_861);
nand U4714 (N_4714,In_486,In_965);
or U4715 (N_4715,In_303,In_2069);
and U4716 (N_4716,In_2856,In_1288);
nand U4717 (N_4717,In_2875,In_2554);
nor U4718 (N_4718,In_2302,In_154);
or U4719 (N_4719,In_341,In_831);
or U4720 (N_4720,In_1608,In_231);
nor U4721 (N_4721,In_2168,In_2666);
and U4722 (N_4722,In_2594,In_1052);
and U4723 (N_4723,In_830,In_2864);
and U4724 (N_4724,In_1758,In_1533);
and U4725 (N_4725,In_1969,In_421);
nand U4726 (N_4726,In_824,In_2173);
nand U4727 (N_4727,In_80,In_2106);
nand U4728 (N_4728,In_1775,In_1544);
nor U4729 (N_4729,In_924,In_979);
nand U4730 (N_4730,In_1216,In_738);
nand U4731 (N_4731,In_440,In_2230);
and U4732 (N_4732,In_1078,In_1907);
nor U4733 (N_4733,In_416,In_813);
nor U4734 (N_4734,In_2358,In_2381);
nand U4735 (N_4735,In_1813,In_2933);
nand U4736 (N_4736,In_2901,In_886);
or U4737 (N_4737,In_1480,In_1389);
nand U4738 (N_4738,In_1872,In_2593);
nand U4739 (N_4739,In_2280,In_2538);
nand U4740 (N_4740,In_2635,In_1098);
nor U4741 (N_4741,In_1881,In_79);
and U4742 (N_4742,In_445,In_2781);
nand U4743 (N_4743,In_2005,In_1597);
nor U4744 (N_4744,In_1767,In_398);
and U4745 (N_4745,In_2000,In_840);
nand U4746 (N_4746,In_1210,In_467);
nor U4747 (N_4747,In_423,In_2884);
and U4748 (N_4748,In_2369,In_1315);
xnor U4749 (N_4749,In_2352,In_2024);
and U4750 (N_4750,In_1698,In_1582);
nor U4751 (N_4751,In_871,In_1536);
nor U4752 (N_4752,In_1679,In_126);
and U4753 (N_4753,In_1992,In_1341);
or U4754 (N_4754,In_2406,In_459);
nand U4755 (N_4755,In_1434,In_1651);
and U4756 (N_4756,In_1582,In_2997);
nor U4757 (N_4757,In_2935,In_606);
and U4758 (N_4758,In_866,In_1022);
nor U4759 (N_4759,In_497,In_1958);
nor U4760 (N_4760,In_1257,In_2694);
and U4761 (N_4761,In_1144,In_1151);
nor U4762 (N_4762,In_2084,In_1466);
nor U4763 (N_4763,In_983,In_899);
nor U4764 (N_4764,In_2765,In_2887);
nand U4765 (N_4765,In_455,In_1073);
and U4766 (N_4766,In_298,In_87);
and U4767 (N_4767,In_2877,In_2341);
nand U4768 (N_4768,In_2275,In_1466);
and U4769 (N_4769,In_2502,In_1021);
nand U4770 (N_4770,In_2779,In_1206);
or U4771 (N_4771,In_1412,In_1696);
nor U4772 (N_4772,In_886,In_411);
nor U4773 (N_4773,In_1797,In_1132);
xor U4774 (N_4774,In_697,In_1429);
nor U4775 (N_4775,In_814,In_2243);
nand U4776 (N_4776,In_2145,In_1361);
and U4777 (N_4777,In_1254,In_409);
or U4778 (N_4778,In_703,In_520);
and U4779 (N_4779,In_1051,In_1149);
nor U4780 (N_4780,In_1751,In_1636);
xor U4781 (N_4781,In_1836,In_1111);
nand U4782 (N_4782,In_2220,In_1064);
and U4783 (N_4783,In_493,In_1621);
and U4784 (N_4784,In_1390,In_957);
nor U4785 (N_4785,In_538,In_588);
nor U4786 (N_4786,In_218,In_638);
and U4787 (N_4787,In_1234,In_2438);
nand U4788 (N_4788,In_1062,In_1001);
and U4789 (N_4789,In_1564,In_2327);
nand U4790 (N_4790,In_831,In_751);
nor U4791 (N_4791,In_1236,In_2639);
nand U4792 (N_4792,In_2414,In_2732);
nor U4793 (N_4793,In_761,In_1925);
nor U4794 (N_4794,In_969,In_1033);
and U4795 (N_4795,In_2679,In_1932);
or U4796 (N_4796,In_1514,In_2541);
or U4797 (N_4797,In_2824,In_1249);
and U4798 (N_4798,In_1822,In_908);
nand U4799 (N_4799,In_1330,In_1764);
or U4800 (N_4800,In_40,In_2953);
nor U4801 (N_4801,In_897,In_1800);
nor U4802 (N_4802,In_2499,In_2262);
and U4803 (N_4803,In_426,In_157);
or U4804 (N_4804,In_1112,In_618);
nor U4805 (N_4805,In_2401,In_2596);
nand U4806 (N_4806,In_2310,In_1130);
and U4807 (N_4807,In_1057,In_1849);
xnor U4808 (N_4808,In_812,In_2009);
nor U4809 (N_4809,In_1654,In_1802);
and U4810 (N_4810,In_1914,In_1977);
or U4811 (N_4811,In_1877,In_325);
nor U4812 (N_4812,In_1106,In_592);
or U4813 (N_4813,In_2241,In_1982);
or U4814 (N_4814,In_809,In_1815);
nand U4815 (N_4815,In_274,In_818);
nand U4816 (N_4816,In_2689,In_1444);
or U4817 (N_4817,In_307,In_1745);
or U4818 (N_4818,In_714,In_653);
nor U4819 (N_4819,In_614,In_1699);
or U4820 (N_4820,In_1372,In_858);
and U4821 (N_4821,In_946,In_1238);
and U4822 (N_4822,In_1087,In_672);
nor U4823 (N_4823,In_368,In_188);
or U4824 (N_4824,In_2440,In_2214);
nor U4825 (N_4825,In_1977,In_933);
xor U4826 (N_4826,In_1905,In_938);
and U4827 (N_4827,In_2868,In_706);
and U4828 (N_4828,In_749,In_2128);
nand U4829 (N_4829,In_2135,In_2022);
nor U4830 (N_4830,In_2797,In_1130);
nand U4831 (N_4831,In_45,In_1400);
nand U4832 (N_4832,In_1598,In_1624);
nand U4833 (N_4833,In_1977,In_1709);
nor U4834 (N_4834,In_1485,In_2804);
or U4835 (N_4835,In_498,In_1059);
nor U4836 (N_4836,In_2291,In_2009);
nor U4837 (N_4837,In_2204,In_16);
nor U4838 (N_4838,In_648,In_1847);
nor U4839 (N_4839,In_1995,In_609);
nor U4840 (N_4840,In_1492,In_925);
nor U4841 (N_4841,In_2020,In_567);
xnor U4842 (N_4842,In_1917,In_1669);
and U4843 (N_4843,In_11,In_1611);
nor U4844 (N_4844,In_2472,In_341);
or U4845 (N_4845,In_2733,In_1825);
nand U4846 (N_4846,In_2708,In_1800);
or U4847 (N_4847,In_2167,In_855);
and U4848 (N_4848,In_400,In_518);
or U4849 (N_4849,In_2635,In_1949);
and U4850 (N_4850,In_2807,In_2919);
or U4851 (N_4851,In_506,In_2075);
nor U4852 (N_4852,In_1432,In_1802);
nand U4853 (N_4853,In_285,In_537);
or U4854 (N_4854,In_1779,In_208);
nand U4855 (N_4855,In_2867,In_485);
and U4856 (N_4856,In_1266,In_86);
nor U4857 (N_4857,In_797,In_473);
and U4858 (N_4858,In_1195,In_1624);
and U4859 (N_4859,In_1013,In_1169);
or U4860 (N_4860,In_1487,In_2507);
or U4861 (N_4861,In_1474,In_2681);
nand U4862 (N_4862,In_425,In_683);
and U4863 (N_4863,In_1897,In_118);
nor U4864 (N_4864,In_101,In_2042);
nor U4865 (N_4865,In_1153,In_154);
xnor U4866 (N_4866,In_73,In_1513);
and U4867 (N_4867,In_2767,In_1286);
and U4868 (N_4868,In_2502,In_1309);
nor U4869 (N_4869,In_78,In_426);
and U4870 (N_4870,In_850,In_1988);
or U4871 (N_4871,In_1097,In_2427);
nand U4872 (N_4872,In_2371,In_1493);
and U4873 (N_4873,In_2179,In_1704);
nor U4874 (N_4874,In_1416,In_871);
and U4875 (N_4875,In_1726,In_385);
nor U4876 (N_4876,In_989,In_1708);
or U4877 (N_4877,In_557,In_780);
or U4878 (N_4878,In_1000,In_1573);
nor U4879 (N_4879,In_613,In_698);
nand U4880 (N_4880,In_756,In_55);
nand U4881 (N_4881,In_268,In_2470);
nand U4882 (N_4882,In_1823,In_1358);
and U4883 (N_4883,In_1299,In_2107);
or U4884 (N_4884,In_77,In_525);
nand U4885 (N_4885,In_1725,In_160);
nand U4886 (N_4886,In_1421,In_1082);
nand U4887 (N_4887,In_1595,In_2246);
nand U4888 (N_4888,In_1590,In_1013);
nor U4889 (N_4889,In_2465,In_1547);
nor U4890 (N_4890,In_1191,In_1501);
nand U4891 (N_4891,In_1446,In_1523);
nand U4892 (N_4892,In_2907,In_972);
or U4893 (N_4893,In_2287,In_125);
nand U4894 (N_4894,In_597,In_966);
nor U4895 (N_4895,In_627,In_1504);
nand U4896 (N_4896,In_2383,In_783);
or U4897 (N_4897,In_1110,In_1458);
nor U4898 (N_4898,In_447,In_1416);
nand U4899 (N_4899,In_1476,In_392);
and U4900 (N_4900,In_1187,In_72);
nand U4901 (N_4901,In_1204,In_2521);
and U4902 (N_4902,In_1445,In_1374);
or U4903 (N_4903,In_591,In_1131);
nor U4904 (N_4904,In_2894,In_1225);
nand U4905 (N_4905,In_2457,In_1867);
and U4906 (N_4906,In_1686,In_555);
and U4907 (N_4907,In_821,In_139);
nor U4908 (N_4908,In_928,In_2528);
and U4909 (N_4909,In_600,In_2237);
and U4910 (N_4910,In_1529,In_2892);
nand U4911 (N_4911,In_2055,In_1608);
nand U4912 (N_4912,In_1729,In_1499);
nor U4913 (N_4913,In_333,In_877);
and U4914 (N_4914,In_1978,In_1953);
and U4915 (N_4915,In_2774,In_2439);
nor U4916 (N_4916,In_2539,In_2172);
and U4917 (N_4917,In_373,In_2671);
nand U4918 (N_4918,In_2786,In_2892);
or U4919 (N_4919,In_1986,In_382);
or U4920 (N_4920,In_1204,In_1555);
and U4921 (N_4921,In_1709,In_1992);
and U4922 (N_4922,In_1275,In_667);
nand U4923 (N_4923,In_1212,In_110);
or U4924 (N_4924,In_2369,In_769);
or U4925 (N_4925,In_1881,In_1600);
nor U4926 (N_4926,In_977,In_1650);
nand U4927 (N_4927,In_2294,In_2199);
nor U4928 (N_4928,In_842,In_2551);
nor U4929 (N_4929,In_1697,In_2307);
and U4930 (N_4930,In_2563,In_1038);
nor U4931 (N_4931,In_2784,In_404);
nand U4932 (N_4932,In_2587,In_802);
or U4933 (N_4933,In_985,In_1865);
nor U4934 (N_4934,In_71,In_1057);
nor U4935 (N_4935,In_2972,In_2364);
nor U4936 (N_4936,In_2984,In_2304);
or U4937 (N_4937,In_269,In_1163);
or U4938 (N_4938,In_159,In_29);
or U4939 (N_4939,In_2277,In_1759);
nor U4940 (N_4940,In_2893,In_979);
or U4941 (N_4941,In_2640,In_2223);
nand U4942 (N_4942,In_2305,In_1291);
and U4943 (N_4943,In_2485,In_370);
nand U4944 (N_4944,In_1587,In_2362);
nor U4945 (N_4945,In_2953,In_219);
xnor U4946 (N_4946,In_15,In_2059);
nor U4947 (N_4947,In_146,In_827);
and U4948 (N_4948,In_92,In_1075);
nor U4949 (N_4949,In_474,In_2406);
or U4950 (N_4950,In_1920,In_1829);
and U4951 (N_4951,In_1443,In_619);
xnor U4952 (N_4952,In_2911,In_976);
nor U4953 (N_4953,In_1507,In_982);
nand U4954 (N_4954,In_2771,In_2424);
or U4955 (N_4955,In_2995,In_2958);
or U4956 (N_4956,In_950,In_1511);
and U4957 (N_4957,In_75,In_2607);
and U4958 (N_4958,In_862,In_2427);
and U4959 (N_4959,In_1468,In_1711);
nor U4960 (N_4960,In_2472,In_1996);
nor U4961 (N_4961,In_2154,In_2613);
nand U4962 (N_4962,In_2963,In_2345);
nor U4963 (N_4963,In_397,In_401);
nor U4964 (N_4964,In_1874,In_2767);
nor U4965 (N_4965,In_2209,In_66);
or U4966 (N_4966,In_1139,In_2186);
nand U4967 (N_4967,In_740,In_860);
nor U4968 (N_4968,In_334,In_1448);
and U4969 (N_4969,In_2636,In_1307);
and U4970 (N_4970,In_782,In_1626);
and U4971 (N_4971,In_2373,In_1833);
nor U4972 (N_4972,In_1664,In_2781);
and U4973 (N_4973,In_1166,In_2297);
nor U4974 (N_4974,In_947,In_2239);
or U4975 (N_4975,In_822,In_2685);
xnor U4976 (N_4976,In_92,In_1813);
or U4977 (N_4977,In_2428,In_850);
and U4978 (N_4978,In_447,In_49);
nor U4979 (N_4979,In_2338,In_101);
or U4980 (N_4980,In_685,In_1097);
or U4981 (N_4981,In_867,In_579);
or U4982 (N_4982,In_2472,In_1485);
and U4983 (N_4983,In_20,In_1224);
nand U4984 (N_4984,In_1901,In_2017);
and U4985 (N_4985,In_1879,In_2068);
and U4986 (N_4986,In_2338,In_1649);
or U4987 (N_4987,In_278,In_1713);
and U4988 (N_4988,In_2772,In_2538);
and U4989 (N_4989,In_2452,In_1702);
or U4990 (N_4990,In_1569,In_1890);
or U4991 (N_4991,In_1699,In_2250);
xor U4992 (N_4992,In_1024,In_1731);
nor U4993 (N_4993,In_2013,In_2566);
and U4994 (N_4994,In_310,In_16);
nor U4995 (N_4995,In_2487,In_1163);
nand U4996 (N_4996,In_1698,In_1705);
or U4997 (N_4997,In_968,In_2726);
and U4998 (N_4998,In_1989,In_1775);
and U4999 (N_4999,In_2151,In_2573);
or U5000 (N_5000,N_3471,N_113);
nor U5001 (N_5001,N_2922,N_2887);
nand U5002 (N_5002,N_799,N_1556);
and U5003 (N_5003,N_3751,N_1144);
nand U5004 (N_5004,N_308,N_1984);
nand U5005 (N_5005,N_2645,N_4698);
nand U5006 (N_5006,N_3431,N_4134);
or U5007 (N_5007,N_887,N_392);
nor U5008 (N_5008,N_1772,N_3227);
nor U5009 (N_5009,N_374,N_2754);
nor U5010 (N_5010,N_2807,N_219);
nor U5011 (N_5011,N_3953,N_1006);
and U5012 (N_5012,N_661,N_2818);
or U5013 (N_5013,N_1744,N_3806);
xor U5014 (N_5014,N_1221,N_2988);
and U5015 (N_5015,N_4822,N_4977);
nor U5016 (N_5016,N_3414,N_1753);
nand U5017 (N_5017,N_633,N_3821);
and U5018 (N_5018,N_1362,N_3469);
or U5019 (N_5019,N_4974,N_51);
nand U5020 (N_5020,N_341,N_3704);
xnor U5021 (N_5021,N_4548,N_994);
nor U5022 (N_5022,N_2871,N_4087);
or U5023 (N_5023,N_3863,N_3797);
nor U5024 (N_5024,N_4445,N_2749);
nand U5025 (N_5025,N_475,N_2723);
nor U5026 (N_5026,N_4888,N_2911);
nor U5027 (N_5027,N_553,N_3947);
and U5028 (N_5028,N_4036,N_2272);
and U5029 (N_5029,N_1651,N_1113);
and U5030 (N_5030,N_686,N_3317);
and U5031 (N_5031,N_5,N_4879);
nand U5032 (N_5032,N_4662,N_3658);
nor U5033 (N_5033,N_3932,N_769);
nand U5034 (N_5034,N_2255,N_3478);
nand U5035 (N_5035,N_2928,N_3544);
or U5036 (N_5036,N_1077,N_3439);
nand U5037 (N_5037,N_330,N_3045);
xor U5038 (N_5038,N_3609,N_34);
nor U5039 (N_5039,N_2934,N_3692);
nand U5040 (N_5040,N_3060,N_3182);
nor U5041 (N_5041,N_4002,N_1389);
nand U5042 (N_5042,N_1852,N_613);
and U5043 (N_5043,N_1882,N_4075);
and U5044 (N_5044,N_4522,N_4613);
nor U5045 (N_5045,N_3400,N_508);
nand U5046 (N_5046,N_1840,N_1616);
and U5047 (N_5047,N_61,N_2487);
nor U5048 (N_5048,N_433,N_956);
or U5049 (N_5049,N_1581,N_1180);
or U5050 (N_5050,N_1212,N_623);
nor U5051 (N_5051,N_1741,N_1769);
nor U5052 (N_5052,N_455,N_3167);
or U5053 (N_5053,N_3738,N_3162);
and U5054 (N_5054,N_2417,N_1631);
nor U5055 (N_5055,N_368,N_3383);
nor U5056 (N_5056,N_3950,N_151);
or U5057 (N_5057,N_1103,N_1764);
nor U5058 (N_5058,N_2616,N_2416);
nand U5059 (N_5059,N_4792,N_532);
nor U5060 (N_5060,N_1355,N_3436);
and U5061 (N_5061,N_3380,N_667);
or U5062 (N_5062,N_3417,N_596);
and U5063 (N_5063,N_4389,N_2232);
nor U5064 (N_5064,N_4606,N_2410);
or U5065 (N_5065,N_2989,N_807);
and U5066 (N_5066,N_1097,N_1543);
or U5067 (N_5067,N_1023,N_4279);
nand U5068 (N_5068,N_4324,N_4925);
nand U5069 (N_5069,N_2980,N_3659);
nand U5070 (N_5070,N_399,N_4432);
or U5071 (N_5071,N_2197,N_2549);
or U5072 (N_5072,N_2111,N_321);
nand U5073 (N_5073,N_831,N_65);
nor U5074 (N_5074,N_3171,N_4494);
nor U5075 (N_5075,N_1228,N_2027);
nand U5076 (N_5076,N_1846,N_2896);
and U5077 (N_5077,N_871,N_1032);
nor U5078 (N_5078,N_4488,N_2314);
and U5079 (N_5079,N_2174,N_1229);
nor U5080 (N_5080,N_4346,N_2265);
and U5081 (N_5081,N_4292,N_3335);
xor U5082 (N_5082,N_2656,N_4198);
nor U5083 (N_5083,N_3212,N_4310);
or U5084 (N_5084,N_3194,N_3986);
xor U5085 (N_5085,N_411,N_1609);
and U5086 (N_5086,N_4111,N_2644);
nor U5087 (N_5087,N_485,N_2681);
nor U5088 (N_5088,N_1266,N_2923);
and U5089 (N_5089,N_4405,N_3141);
or U5090 (N_5090,N_4618,N_4766);
or U5091 (N_5091,N_645,N_940);
or U5092 (N_5092,N_3865,N_766);
and U5093 (N_5093,N_3581,N_1201);
nor U5094 (N_5094,N_2610,N_3290);
and U5095 (N_5095,N_1509,N_3463);
and U5096 (N_5096,N_3628,N_179);
or U5097 (N_5097,N_4490,N_1739);
nand U5098 (N_5098,N_4506,N_131);
nand U5099 (N_5099,N_3621,N_3473);
nor U5100 (N_5100,N_4776,N_753);
nand U5101 (N_5101,N_2028,N_2356);
and U5102 (N_5102,N_3745,N_3418);
and U5103 (N_5103,N_2408,N_3457);
and U5104 (N_5104,N_2112,N_881);
or U5105 (N_5105,N_13,N_4765);
or U5106 (N_5106,N_3352,N_2971);
nand U5107 (N_5107,N_2118,N_3152);
or U5108 (N_5108,N_4362,N_4916);
nor U5109 (N_5109,N_4273,N_1811);
and U5110 (N_5110,N_2413,N_1928);
nand U5111 (N_5111,N_3861,N_2336);
nand U5112 (N_5112,N_487,N_2013);
nand U5113 (N_5113,N_1994,N_1165);
and U5114 (N_5114,N_748,N_1506);
or U5115 (N_5115,N_561,N_1937);
nor U5116 (N_5116,N_4746,N_1956);
and U5117 (N_5117,N_3358,N_1761);
or U5118 (N_5118,N_4993,N_3511);
and U5119 (N_5119,N_1197,N_1752);
nand U5120 (N_5120,N_3228,N_339);
nor U5121 (N_5121,N_4205,N_544);
nand U5122 (N_5122,N_4825,N_878);
or U5123 (N_5123,N_2173,N_3901);
and U5124 (N_5124,N_3730,N_1474);
nand U5125 (N_5125,N_3618,N_1563);
nor U5126 (N_5126,N_1511,N_194);
nand U5127 (N_5127,N_3769,N_3148);
nor U5128 (N_5128,N_2469,N_4338);
or U5129 (N_5129,N_4539,N_583);
nand U5130 (N_5130,N_1710,N_1002);
nand U5131 (N_5131,N_3173,N_1749);
or U5132 (N_5132,N_707,N_555);
and U5133 (N_5133,N_4054,N_3153);
or U5134 (N_5134,N_3623,N_3928);
nor U5135 (N_5135,N_2148,N_873);
or U5136 (N_5136,N_1379,N_554);
nand U5137 (N_5137,N_1569,N_3568);
nor U5138 (N_5138,N_4067,N_70);
nand U5139 (N_5139,N_593,N_3438);
and U5140 (N_5140,N_1294,N_3266);
nor U5141 (N_5141,N_2052,N_134);
nor U5142 (N_5142,N_393,N_215);
or U5143 (N_5143,N_1137,N_971);
or U5144 (N_5144,N_4039,N_3886);
and U5145 (N_5145,N_1162,N_2855);
nor U5146 (N_5146,N_246,N_284);
and U5147 (N_5147,N_3739,N_1155);
or U5148 (N_5148,N_582,N_506);
nand U5149 (N_5149,N_1341,N_88);
nand U5150 (N_5150,N_4838,N_1650);
nand U5151 (N_5151,N_3512,N_1558);
nand U5152 (N_5152,N_3441,N_2169);
nor U5153 (N_5153,N_813,N_2322);
and U5154 (N_5154,N_2637,N_3295);
nor U5155 (N_5155,N_4452,N_1958);
and U5156 (N_5156,N_1330,N_3563);
nor U5157 (N_5157,N_2386,N_2977);
nor U5158 (N_5158,N_1570,N_663);
and U5159 (N_5159,N_1408,N_3864);
or U5160 (N_5160,N_4693,N_493);
nand U5161 (N_5161,N_4085,N_4008);
nor U5162 (N_5162,N_3343,N_3852);
or U5163 (N_5163,N_2390,N_2668);
nor U5164 (N_5164,N_1013,N_754);
and U5165 (N_5165,N_4632,N_4677);
or U5166 (N_5166,N_3482,N_2757);
nand U5167 (N_5167,N_298,N_3231);
and U5168 (N_5168,N_4774,N_3550);
nand U5169 (N_5169,N_4403,N_4917);
or U5170 (N_5170,N_4031,N_3775);
or U5171 (N_5171,N_2725,N_4569);
and U5172 (N_5172,N_4588,N_4713);
and U5173 (N_5173,N_840,N_1678);
nand U5174 (N_5174,N_1635,N_2569);
nand U5175 (N_5175,N_2770,N_300);
nand U5176 (N_5176,N_4985,N_4946);
nor U5177 (N_5177,N_1135,N_1272);
and U5178 (N_5178,N_4026,N_4453);
or U5179 (N_5179,N_517,N_477);
and U5180 (N_5180,N_2245,N_3236);
and U5181 (N_5181,N_2850,N_189);
or U5182 (N_5182,N_3750,N_1005);
nand U5183 (N_5183,N_597,N_981);
or U5184 (N_5184,N_3364,N_2976);
or U5185 (N_5185,N_4108,N_802);
or U5186 (N_5186,N_1093,N_240);
or U5187 (N_5187,N_446,N_3934);
or U5188 (N_5188,N_49,N_4733);
nor U5189 (N_5189,N_3712,N_2638);
nor U5190 (N_5190,N_1323,N_2744);
nand U5191 (N_5191,N_1542,N_4233);
nor U5192 (N_5192,N_1458,N_1274);
or U5193 (N_5193,N_2552,N_1056);
nor U5194 (N_5194,N_2722,N_4411);
nor U5195 (N_5195,N_458,N_3034);
nor U5196 (N_5196,N_3732,N_4410);
nand U5197 (N_5197,N_3063,N_4631);
or U5198 (N_5198,N_4248,N_1510);
nand U5199 (N_5199,N_1345,N_4671);
nand U5200 (N_5200,N_1564,N_1530);
or U5201 (N_5201,N_3201,N_4501);
and U5202 (N_5202,N_1911,N_698);
nand U5203 (N_5203,N_3940,N_1694);
nor U5204 (N_5204,N_1528,N_573);
nand U5205 (N_5205,N_237,N_1433);
nor U5206 (N_5206,N_2325,N_2539);
and U5207 (N_5207,N_932,N_1724);
and U5208 (N_5208,N_4999,N_4096);
and U5209 (N_5209,N_3240,N_1876);
nor U5210 (N_5210,N_262,N_2223);
or U5211 (N_5211,N_3718,N_2662);
or U5212 (N_5212,N_3577,N_1173);
nor U5213 (N_5213,N_2432,N_2987);
nand U5214 (N_5214,N_3019,N_3238);
nor U5215 (N_5215,N_4546,N_4424);
and U5216 (N_5216,N_4858,N_1311);
nand U5217 (N_5217,N_3580,N_2158);
or U5218 (N_5218,N_3232,N_816);
nand U5219 (N_5219,N_1169,N_733);
nor U5220 (N_5220,N_3790,N_1803);
and U5221 (N_5221,N_647,N_941);
and U5222 (N_5222,N_3432,N_2563);
nor U5223 (N_5223,N_87,N_2983);
and U5224 (N_5224,N_849,N_4296);
or U5225 (N_5225,N_4830,N_25);
or U5226 (N_5226,N_92,N_4619);
or U5227 (N_5227,N_3257,N_4213);
nor U5228 (N_5228,N_2742,N_3694);
nor U5229 (N_5229,N_3341,N_1046);
or U5230 (N_5230,N_352,N_514);
nor U5231 (N_5231,N_3858,N_2259);
nor U5232 (N_5232,N_4747,N_2992);
and U5233 (N_5233,N_4605,N_3768);
nand U5234 (N_5234,N_3848,N_4016);
and U5235 (N_5235,N_2186,N_2331);
and U5236 (N_5236,N_1053,N_4431);
and U5237 (N_5237,N_1520,N_4633);
nand U5238 (N_5238,N_3758,N_1168);
nor U5239 (N_5239,N_2229,N_1125);
nand U5240 (N_5240,N_2535,N_1797);
nand U5241 (N_5241,N_2915,N_960);
and U5242 (N_5242,N_270,N_6);
nand U5243 (N_5243,N_217,N_901);
nor U5244 (N_5244,N_3582,N_4552);
nor U5245 (N_5245,N_4795,N_2738);
and U5246 (N_5246,N_4065,N_4103);
nor U5247 (N_5247,N_1954,N_1017);
nand U5248 (N_5248,N_518,N_502);
and U5249 (N_5249,N_2652,N_775);
or U5250 (N_5250,N_3005,N_3393);
and U5251 (N_5251,N_3936,N_90);
or U5252 (N_5252,N_157,N_1337);
nor U5253 (N_5253,N_4758,N_3389);
nor U5254 (N_5254,N_4926,N_2583);
nand U5255 (N_5255,N_2809,N_1210);
nand U5256 (N_5256,N_2709,N_2454);
or U5257 (N_5257,N_4586,N_2448);
and U5258 (N_5258,N_1880,N_4268);
nand U5259 (N_5259,N_1469,N_1845);
or U5260 (N_5260,N_3595,N_2058);
or U5261 (N_5261,N_4590,N_3048);
and U5262 (N_5262,N_1282,N_171);
nor U5263 (N_5263,N_1720,N_2603);
and U5264 (N_5264,N_1964,N_4291);
nand U5265 (N_5265,N_4479,N_2654);
and U5266 (N_5266,N_2659,N_4629);
or U5267 (N_5267,N_4173,N_1603);
nand U5268 (N_5268,N_2401,N_3449);
or U5269 (N_5269,N_291,N_4033);
and U5270 (N_5270,N_132,N_2753);
and U5271 (N_5271,N_4148,N_1472);
nor U5272 (N_5272,N_423,N_2760);
nor U5273 (N_5273,N_2385,N_3668);
nand U5274 (N_5274,N_3320,N_2528);
or U5275 (N_5275,N_3873,N_1717);
or U5276 (N_5276,N_695,N_1050);
or U5277 (N_5277,N_907,N_2370);
nor U5278 (N_5278,N_4832,N_3620);
nor U5279 (N_5279,N_377,N_2511);
nor U5280 (N_5280,N_3476,N_2927);
nand U5281 (N_5281,N_636,N_1574);
or U5282 (N_5282,N_1677,N_144);
and U5283 (N_5283,N_4601,N_1837);
nor U5284 (N_5284,N_1821,N_2721);
nand U5285 (N_5285,N_2363,N_566);
nor U5286 (N_5286,N_187,N_2578);
nor U5287 (N_5287,N_2237,N_4647);
nand U5288 (N_5288,N_1889,N_3924);
xor U5289 (N_5289,N_2402,N_495);
nand U5290 (N_5290,N_1213,N_3448);
nand U5291 (N_5291,N_142,N_4630);
nand U5292 (N_5292,N_811,N_806);
xnor U5293 (N_5293,N_2618,N_1532);
nand U5294 (N_5294,N_2999,N_2559);
or U5295 (N_5295,N_2764,N_2005);
and U5296 (N_5296,N_965,N_4611);
or U5297 (N_5297,N_1926,N_513);
nand U5298 (N_5298,N_2040,N_2864);
and U5299 (N_5299,N_912,N_617);
nor U5300 (N_5300,N_82,N_4669);
and U5301 (N_5301,N_4721,N_504);
and U5302 (N_5302,N_4901,N_2920);
or U5303 (N_5303,N_2772,N_417);
or U5304 (N_5304,N_1305,N_299);
nor U5305 (N_5305,N_3744,N_1824);
or U5306 (N_5306,N_4166,N_1263);
or U5307 (N_5307,N_4339,N_2095);
and U5308 (N_5308,N_2160,N_3402);
and U5309 (N_5309,N_2224,N_3661);
or U5310 (N_5310,N_2010,N_4518);
nand U5311 (N_5311,N_325,N_2107);
and U5312 (N_5312,N_810,N_4331);
or U5313 (N_5313,N_3079,N_1499);
nand U5314 (N_5314,N_3660,N_2425);
or U5315 (N_5315,N_955,N_3771);
nand U5316 (N_5316,N_4961,N_1969);
or U5317 (N_5317,N_39,N_3589);
or U5318 (N_5318,N_1288,N_129);
or U5319 (N_5319,N_1445,N_734);
nor U5320 (N_5320,N_2137,N_3631);
and U5321 (N_5321,N_2323,N_3382);
or U5322 (N_5322,N_854,N_1416);
nor U5323 (N_5323,N_3230,N_1854);
nand U5324 (N_5324,N_265,N_3016);
and U5325 (N_5325,N_2329,N_4853);
nor U5326 (N_5326,N_4734,N_3994);
nand U5327 (N_5327,N_2514,N_2227);
or U5328 (N_5328,N_2308,N_4060);
or U5329 (N_5329,N_3114,N_1063);
nor U5330 (N_5330,N_1191,N_4711);
nand U5331 (N_5331,N_4987,N_3566);
or U5332 (N_5332,N_4221,N_2188);
or U5333 (N_5333,N_3875,N_457);
and U5334 (N_5334,N_2817,N_4818);
nand U5335 (N_5335,N_4392,N_842);
nor U5336 (N_5336,N_4791,N_4582);
xor U5337 (N_5337,N_2601,N_4653);
nor U5338 (N_5338,N_11,N_653);
or U5339 (N_5339,N_551,N_2783);
or U5340 (N_5340,N_4914,N_4335);
nor U5341 (N_5341,N_601,N_334);
nand U5342 (N_5342,N_2661,N_1388);
nor U5343 (N_5343,N_1524,N_4425);
xnor U5344 (N_5344,N_97,N_1042);
or U5345 (N_5345,N_1951,N_84);
or U5346 (N_5346,N_1832,N_4730);
nand U5347 (N_5347,N_2214,N_3639);
or U5348 (N_5348,N_3155,N_2043);
or U5349 (N_5349,N_1273,N_2543);
or U5350 (N_5350,N_1205,N_4312);
nand U5351 (N_5351,N_1881,N_4402);
nand U5352 (N_5352,N_1547,N_2919);
nor U5353 (N_5353,N_3849,N_997);
nor U5354 (N_5354,N_486,N_4604);
nand U5355 (N_5355,N_1190,N_1942);
and U5356 (N_5356,N_3465,N_700);
and U5357 (N_5357,N_2253,N_3951);
or U5358 (N_5358,N_3426,N_1602);
nand U5359 (N_5359,N_0,N_3138);
nor U5360 (N_5360,N_1498,N_2330);
nor U5361 (N_5361,N_2883,N_440);
nand U5362 (N_5362,N_4862,N_1645);
xnor U5363 (N_5363,N_470,N_4382);
or U5364 (N_5364,N_2079,N_1309);
nand U5365 (N_5365,N_3267,N_3921);
and U5366 (N_5366,N_4160,N_4602);
nor U5367 (N_5367,N_4640,N_4478);
or U5368 (N_5368,N_1242,N_3381);
nand U5369 (N_5369,N_1935,N_3018);
and U5370 (N_5370,N_4919,N_4531);
and U5371 (N_5371,N_4367,N_3397);
nand U5372 (N_5372,N_4695,N_4442);
nor U5373 (N_5373,N_1733,N_787);
or U5374 (N_5374,N_4882,N_2714);
or U5375 (N_5375,N_1027,N_3565);
nor U5376 (N_5376,N_1598,N_3347);
or U5377 (N_5377,N_3052,N_1187);
and U5378 (N_5378,N_4361,N_3995);
nor U5379 (N_5379,N_1922,N_4448);
and U5380 (N_5380,N_3029,N_1058);
and U5381 (N_5381,N_953,N_2996);
nand U5382 (N_5382,N_426,N_3579);
nand U5383 (N_5383,N_533,N_4089);
nand U5384 (N_5384,N_2975,N_4827);
or U5385 (N_5385,N_3386,N_148);
nor U5386 (N_5386,N_1421,N_4023);
nor U5387 (N_5387,N_1727,N_1507);
nand U5388 (N_5388,N_4011,N_2083);
nor U5389 (N_5389,N_3273,N_1949);
xor U5390 (N_5390,N_1658,N_139);
and U5391 (N_5391,N_4145,N_681);
and U5392 (N_5392,N_3679,N_2476);
or U5393 (N_5393,N_1847,N_2490);
nor U5394 (N_5394,N_3773,N_3388);
nand U5395 (N_5395,N_1784,N_4028);
or U5396 (N_5396,N_2282,N_2641);
nor U5397 (N_5397,N_851,N_843);
nand U5398 (N_5398,N_3355,N_762);
or U5399 (N_5399,N_80,N_560);
and U5400 (N_5400,N_407,N_2985);
or U5401 (N_5401,N_1116,N_678);
or U5402 (N_5402,N_1249,N_1833);
or U5403 (N_5403,N_1062,N_2504);
nand U5404 (N_5404,N_4610,N_516);
nor U5405 (N_5405,N_1166,N_2679);
nand U5406 (N_5406,N_177,N_2249);
or U5407 (N_5407,N_3390,N_3825);
and U5408 (N_5408,N_2834,N_2865);
nor U5409 (N_5409,N_1095,N_4068);
and U5410 (N_5410,N_208,N_3051);
nand U5411 (N_5411,N_136,N_163);
nor U5412 (N_5412,N_895,N_3695);
and U5413 (N_5413,N_3464,N_4270);
and U5414 (N_5414,N_3766,N_4568);
or U5415 (N_5415,N_4971,N_315);
or U5416 (N_5416,N_3487,N_2542);
nand U5417 (N_5417,N_401,N_292);
nor U5418 (N_5418,N_2993,N_4199);
and U5419 (N_5419,N_4664,N_3866);
and U5420 (N_5420,N_1427,N_4193);
and U5421 (N_5421,N_4401,N_982);
or U5422 (N_5422,N_846,N_4885);
or U5423 (N_5423,N_1009,N_4941);
nand U5424 (N_5424,N_540,N_3637);
or U5425 (N_5425,N_791,N_2824);
nor U5426 (N_5426,N_1703,N_375);
and U5427 (N_5427,N_1684,N_2051);
nand U5428 (N_5428,N_4377,N_3387);
nand U5429 (N_5429,N_478,N_3968);
and U5430 (N_5430,N_225,N_4197);
and U5431 (N_5431,N_1227,N_4482);
nor U5432 (N_5432,N_2859,N_3998);
nand U5433 (N_5433,N_1292,N_3818);
or U5434 (N_5434,N_2577,N_2619);
nor U5435 (N_5435,N_1214,N_4172);
and U5436 (N_5436,N_992,N_4235);
or U5437 (N_5437,N_3578,N_3413);
or U5438 (N_5438,N_2289,N_2593);
or U5439 (N_5439,N_1156,N_4871);
and U5440 (N_5440,N_4264,N_574);
and U5441 (N_5441,N_1394,N_3095);
nand U5442 (N_5442,N_2130,N_931);
nand U5443 (N_5443,N_4238,N_4020);
nand U5444 (N_5444,N_1189,N_4051);
and U5445 (N_5445,N_2302,N_4041);
nor U5446 (N_5446,N_1217,N_987);
and U5447 (N_5447,N_3931,N_2565);
nand U5448 (N_5448,N_3604,N_3147);
nor U5449 (N_5449,N_3635,N_1484);
or U5450 (N_5450,N_4934,N_1517);
nor U5451 (N_5451,N_2545,N_2254);
nor U5452 (N_5452,N_4826,N_3237);
or U5453 (N_5453,N_2660,N_1026);
or U5454 (N_5454,N_1008,N_2405);
nor U5455 (N_5455,N_926,N_723);
or U5456 (N_5456,N_4689,N_4790);
nor U5457 (N_5457,N_3027,N_3779);
and U5458 (N_5458,N_1959,N_3453);
and U5459 (N_5459,N_2632,N_1149);
or U5460 (N_5460,N_2801,N_213);
and U5461 (N_5461,N_3247,N_640);
and U5462 (N_5462,N_3530,N_903);
or U5463 (N_5463,N_4404,N_4299);
nor U5464 (N_5464,N_4315,N_2030);
xor U5465 (N_5465,N_2665,N_883);
nor U5466 (N_5466,N_1962,N_2422);
or U5467 (N_5467,N_1885,N_2019);
nor U5468 (N_5468,N_2394,N_2306);
nor U5469 (N_5469,N_602,N_2324);
nor U5470 (N_5470,N_3896,N_3493);
and U5471 (N_5471,N_2343,N_1486);
and U5472 (N_5472,N_2586,N_1407);
nand U5473 (N_5473,N_1578,N_2775);
nand U5474 (N_5474,N_1184,N_4994);
and U5475 (N_5475,N_4712,N_2344);
and U5476 (N_5476,N_379,N_185);
and U5477 (N_5477,N_2544,N_3788);
nand U5478 (N_5478,N_1634,N_1986);
and U5479 (N_5479,N_1848,N_1216);
nand U5480 (N_5480,N_1434,N_1568);
nand U5481 (N_5481,N_4716,N_1841);
or U5482 (N_5482,N_2066,N_3084);
and U5483 (N_5483,N_3172,N_1024);
nor U5484 (N_5484,N_1451,N_1731);
nand U5485 (N_5485,N_2149,N_2573);
or U5486 (N_5486,N_4256,N_4742);
nand U5487 (N_5487,N_1734,N_4966);
nand U5488 (N_5488,N_4509,N_3020);
and U5489 (N_5489,N_3937,N_2268);
and U5490 (N_5490,N_3624,N_3834);
or U5491 (N_5491,N_3612,N_2113);
and U5492 (N_5492,N_2575,N_3442);
nand U5493 (N_5493,N_3075,N_4210);
and U5494 (N_5494,N_1237,N_1614);
or U5495 (N_5495,N_2252,N_3759);
or U5496 (N_5496,N_3456,N_911);
or U5497 (N_5497,N_4617,N_803);
or U5498 (N_5498,N_4709,N_4697);
nor U5499 (N_5499,N_1610,N_4848);
or U5500 (N_5500,N_2202,N_3916);
nor U5501 (N_5501,N_3702,N_3686);
or U5502 (N_5502,N_863,N_3696);
or U5503 (N_5503,N_3502,N_1932);
nand U5504 (N_5504,N_1646,N_1145);
nor U5505 (N_5505,N_3408,N_2806);
and U5506 (N_5506,N_790,N_4038);
nor U5507 (N_5507,N_3481,N_4313);
and U5508 (N_5508,N_1182,N_3619);
or U5509 (N_5509,N_2065,N_4540);
nor U5510 (N_5510,N_59,N_1898);
or U5511 (N_5511,N_3165,N_1877);
and U5512 (N_5512,N_1334,N_1419);
and U5513 (N_5513,N_957,N_3124);
and U5514 (N_5514,N_4355,N_1508);
nor U5515 (N_5515,N_2326,N_3601);
or U5516 (N_5516,N_4151,N_4787);
nand U5517 (N_5517,N_3351,N_1112);
and U5518 (N_5518,N_2328,N_4187);
and U5519 (N_5519,N_4870,N_2068);
nor U5520 (N_5520,N_557,N_1409);
nand U5521 (N_5521,N_336,N_3708);
and U5522 (N_5522,N_2024,N_897);
or U5523 (N_5523,N_4722,N_3688);
nand U5524 (N_5524,N_2566,N_4708);
and U5525 (N_5525,N_4573,N_968);
nor U5526 (N_5526,N_2953,N_3908);
nand U5527 (N_5527,N_2843,N_1482);
or U5528 (N_5528,N_2063,N_3583);
nand U5529 (N_5529,N_1701,N_3282);
nand U5530 (N_5530,N_329,N_474);
nand U5531 (N_5531,N_744,N_1015);
or U5532 (N_5532,N_4053,N_660);
and U5533 (N_5533,N_963,N_1522);
nand U5534 (N_5534,N_2978,N_1295);
or U5535 (N_5535,N_234,N_4559);
nor U5536 (N_5536,N_2167,N_1891);
nand U5537 (N_5537,N_2768,N_4168);
or U5538 (N_5538,N_1514,N_3706);
and U5539 (N_5539,N_886,N_4793);
and U5540 (N_5540,N_824,N_1944);
or U5541 (N_5541,N_1034,N_755);
and U5542 (N_5542,N_4088,N_4308);
nand U5543 (N_5543,N_2203,N_739);
nand U5544 (N_5544,N_4353,N_2415);
and U5545 (N_5545,N_4665,N_679);
and U5546 (N_5546,N_2269,N_2582);
nand U5547 (N_5547,N_3,N_3683);
nand U5548 (N_5548,N_2060,N_2550);
nor U5549 (N_5549,N_162,N_945);
and U5550 (N_5550,N_218,N_1296);
or U5551 (N_5551,N_2631,N_4284);
nand U5552 (N_5552,N_4883,N_1018);
nor U5553 (N_5553,N_2342,N_1813);
and U5554 (N_5554,N_1719,N_2091);
and U5555 (N_5555,N_2524,N_91);
nand U5556 (N_5556,N_258,N_3359);
or U5557 (N_5557,N_1400,N_4984);
or U5558 (N_5558,N_4182,N_2092);
nor U5559 (N_5559,N_4816,N_3137);
xnor U5560 (N_5560,N_4077,N_1106);
nor U5561 (N_5561,N_4904,N_2478);
and U5562 (N_5562,N_2685,N_2481);
or U5563 (N_5563,N_1086,N_4202);
nor U5564 (N_5564,N_721,N_2451);
or U5565 (N_5565,N_1108,N_4578);
or U5566 (N_5566,N_4288,N_2621);
nor U5567 (N_5567,N_3178,N_1085);
and U5568 (N_5568,N_4345,N_2875);
nand U5569 (N_5569,N_3203,N_1192);
nor U5570 (N_5570,N_605,N_3633);
and U5571 (N_5571,N_2860,N_3607);
and U5572 (N_5572,N_2284,N_2574);
and U5573 (N_5573,N_4439,N_2743);
or U5574 (N_5574,N_937,N_4340);
nor U5575 (N_5575,N_3764,N_2138);
and U5576 (N_5576,N_364,N_3354);
or U5577 (N_5577,N_1792,N_4359);
or U5578 (N_5578,N_4413,N_2888);
nand U5579 (N_5579,N_4139,N_3851);
or U5580 (N_5580,N_924,N_2151);
and U5581 (N_5581,N_765,N_4474);
nand U5582 (N_5582,N_1397,N_2041);
nand U5583 (N_5583,N_3353,N_2280);
nor U5584 (N_5584,N_3562,N_355);
nor U5585 (N_5585,N_1254,N_4368);
nand U5586 (N_5586,N_480,N_2810);
or U5587 (N_5587,N_3100,N_3000);
nand U5588 (N_5588,N_2187,N_718);
or U5589 (N_5589,N_2436,N_4880);
nand U5590 (N_5590,N_2502,N_3008);
nand U5591 (N_5591,N_3707,N_115);
and U5592 (N_5592,N_670,N_2702);
and U5593 (N_5593,N_2628,N_4833);
or U5594 (N_5594,N_4622,N_1780);
xor U5595 (N_5595,N_4374,N_2781);
or U5596 (N_5596,N_1315,N_111);
nor U5597 (N_5597,N_4995,N_4222);
and U5598 (N_5598,N_3551,N_3017);
and U5599 (N_5599,N_951,N_4678);
nor U5600 (N_5600,N_1136,N_2930);
nor U5601 (N_5601,N_1834,N_4010);
and U5602 (N_5602,N_122,N_1915);
nor U5603 (N_5603,N_4086,N_200);
nand U5604 (N_5604,N_4098,N_3765);
and U5605 (N_5605,N_858,N_3844);
nand U5606 (N_5606,N_2921,N_4846);
and U5607 (N_5607,N_4956,N_4246);
nor U5608 (N_5608,N_2751,N_2391);
xor U5609 (N_5609,N_3556,N_4450);
nor U5610 (N_5610,N_1453,N_3762);
nand U5611 (N_5611,N_4484,N_736);
and U5612 (N_5612,N_3570,N_2874);
nor U5613 (N_5613,N_644,N_4052);
nor U5614 (N_5614,N_1328,N_212);
nand U5615 (N_5615,N_3475,N_1467);
and U5616 (N_5616,N_3823,N_1100);
and U5617 (N_5617,N_844,N_2192);
and U5618 (N_5618,N_993,N_4543);
and U5619 (N_5619,N_288,N_2366);
and U5620 (N_5620,N_2036,N_3820);
and U5621 (N_5621,N_4529,N_3677);
nand U5622 (N_5622,N_915,N_247);
nand U5623 (N_5623,N_4266,N_402);
and U5624 (N_5624,N_2791,N_668);
nor U5625 (N_5625,N_4682,N_4864);
and U5626 (N_5626,N_1704,N_3539);
nor U5627 (N_5627,N_2142,N_3776);
nor U5628 (N_5628,N_1698,N_847);
nand U5629 (N_5629,N_2498,N_1975);
or U5630 (N_5630,N_1456,N_826);
nor U5631 (N_5631,N_2995,N_1934);
or U5632 (N_5632,N_1748,N_3085);
nand U5633 (N_5633,N_4656,N_4924);
or U5634 (N_5634,N_1000,N_4133);
or U5635 (N_5635,N_2313,N_1857);
nand U5636 (N_5636,N_2305,N_4657);
or U5637 (N_5637,N_793,N_1625);
nand U5638 (N_5638,N_46,N_1504);
or U5639 (N_5639,N_1391,N_2033);
nand U5640 (N_5640,N_1529,N_4125);
and U5641 (N_5641,N_3042,N_3433);
or U5642 (N_5642,N_2968,N_950);
and U5643 (N_5643,N_1683,N_4867);
nand U5644 (N_5644,N_1488,N_1978);
nand U5645 (N_5645,N_3109,N_81);
nor U5646 (N_5646,N_4627,N_2439);
or U5647 (N_5647,N_4706,N_3028);
and U5648 (N_5648,N_2933,N_361);
xor U5649 (N_5649,N_2763,N_3547);
or U5650 (N_5650,N_1033,N_666);
and U5651 (N_5651,N_439,N_1897);
and U5652 (N_5652,N_4206,N_4527);
and U5653 (N_5653,N_2758,N_2945);
or U5654 (N_5654,N_152,N_4255);
nor U5655 (N_5655,N_386,N_2720);
and U5656 (N_5656,N_1540,N_4165);
and U5657 (N_5657,N_4978,N_3139);
or U5658 (N_5658,N_2053,N_4524);
nor U5659 (N_5659,N_2312,N_722);
and U5660 (N_5660,N_3316,N_4936);
and U5661 (N_5661,N_4217,N_121);
nand U5662 (N_5662,N_1552,N_3786);
or U5663 (N_5663,N_4550,N_453);
or U5664 (N_5664,N_1723,N_3300);
nor U5665 (N_5665,N_3061,N_720);
or U5666 (N_5666,N_2939,N_1953);
nor U5667 (N_5667,N_449,N_1548);
and U5668 (N_5668,N_1707,N_4045);
or U5669 (N_5669,N_1437,N_45);
and U5670 (N_5670,N_1587,N_3549);
or U5671 (N_5671,N_1550,N_1464);
nor U5672 (N_5672,N_3719,N_3122);
nor U5673 (N_5673,N_3149,N_4492);
or U5674 (N_5674,N_2195,N_335);
nor U5675 (N_5675,N_3218,N_3368);
or U5676 (N_5676,N_4112,N_899);
and U5677 (N_5677,N_2471,N_4763);
and U5678 (N_5678,N_1340,N_1527);
nand U5679 (N_5679,N_2465,N_468);
or U5680 (N_5680,N_3699,N_4583);
or U5681 (N_5681,N_2713,N_1431);
and U5682 (N_5682,N_2275,N_3342);
or U5683 (N_5683,N_760,N_2020);
and U5684 (N_5684,N_1064,N_1204);
and U5685 (N_5685,N_2548,N_4819);
and U5686 (N_5686,N_4473,N_4136);
and U5687 (N_5687,N_1025,N_3690);
nor U5688 (N_5688,N_3591,N_1060);
xor U5689 (N_5689,N_1545,N_3271);
and U5690 (N_5690,N_4400,N_3336);
or U5691 (N_5691,N_558,N_2178);
nor U5692 (N_5692,N_4581,N_4660);
and U5693 (N_5693,N_4293,N_3437);
nand U5694 (N_5694,N_4979,N_4223);
xor U5695 (N_5695,N_3800,N_4072);
or U5696 (N_5696,N_526,N_1370);
or U5697 (N_5697,N_2145,N_4881);
nor U5698 (N_5698,N_301,N_4937);
nor U5699 (N_5699,N_1745,N_2581);
nor U5700 (N_5700,N_3461,N_4130);
and U5701 (N_5701,N_3902,N_4218);
nand U5702 (N_5702,N_3312,N_1479);
nand U5703 (N_5703,N_1124,N_1549);
nor U5704 (N_5704,N_3314,N_4426);
or U5705 (N_5705,N_2081,N_268);
and U5706 (N_5706,N_4754,N_777);
and U5707 (N_5707,N_444,N_1048);
nand U5708 (N_5708,N_3422,N_1485);
nand U5709 (N_5709,N_3332,N_3292);
and U5710 (N_5710,N_1406,N_1059);
or U5711 (N_5711,N_1615,N_1220);
or U5712 (N_5712,N_3647,N_853);
and U5713 (N_5713,N_2979,N_1890);
or U5714 (N_5714,N_2537,N_4334);
or U5715 (N_5715,N_984,N_3987);
and U5716 (N_5716,N_2827,N_1314);
or U5717 (N_5717,N_1285,N_3385);
nand U5718 (N_5718,N_884,N_357);
nor U5719 (N_5719,N_4813,N_2453);
nand U5720 (N_5720,N_3898,N_48);
and U5721 (N_5721,N_4078,N_4342);
nand U5722 (N_5722,N_2338,N_178);
and U5723 (N_5723,N_4634,N_559);
nand U5724 (N_5724,N_3564,N_2411);
and U5725 (N_5725,N_995,N_4037);
nand U5726 (N_5726,N_4156,N_3962);
nor U5727 (N_5727,N_2935,N_4421);
nor U5728 (N_5728,N_3653,N_834);
or U5729 (N_5729,N_2840,N_2078);
nor U5730 (N_5730,N_1102,N_1712);
or U5731 (N_5731,N_1566,N_2890);
or U5732 (N_5732,N_2147,N_1147);
nor U5733 (N_5733,N_1157,N_3662);
nand U5734 (N_5734,N_2916,N_4262);
nand U5735 (N_5735,N_3545,N_2734);
nor U5736 (N_5736,N_3614,N_1491);
and U5737 (N_5737,N_376,N_1061);
xnor U5738 (N_5738,N_1332,N_2477);
or U5739 (N_5739,N_192,N_3626);
nand U5740 (N_5740,N_652,N_1721);
and U5741 (N_5741,N_1644,N_3958);
or U5742 (N_5742,N_1791,N_3836);
nor U5743 (N_5743,N_1230,N_310);
and U5744 (N_5744,N_4675,N_1259);
nor U5745 (N_5745,N_4106,N_2963);
and U5746 (N_5746,N_3829,N_1240);
and U5747 (N_5747,N_1763,N_1682);
nand U5748 (N_5748,N_4574,N_2794);
and U5749 (N_5749,N_1084,N_935);
nor U5750 (N_5750,N_4872,N_3957);
and U5751 (N_5751,N_890,N_2318);
or U5752 (N_5752,N_1830,N_3313);
or U5753 (N_5753,N_221,N_2505);
or U5754 (N_5754,N_2771,N_1265);
or U5755 (N_5755,N_1836,N_1174);
nor U5756 (N_5756,N_3443,N_1668);
or U5757 (N_5757,N_629,N_2728);
and U5758 (N_5758,N_3590,N_348);
or U5759 (N_5759,N_4686,N_1535);
nand U5760 (N_5760,N_4241,N_1659);
or U5761 (N_5761,N_2348,N_898);
nor U5762 (N_5762,N_3177,N_4175);
and U5763 (N_5763,N_3792,N_713);
nand U5764 (N_5764,N_4207,N_1041);
and U5765 (N_5765,N_4080,N_1577);
or U5766 (N_5766,N_1247,N_1781);
nand U5767 (N_5767,N_1773,N_175);
and U5768 (N_5768,N_1133,N_1359);
nand U5769 (N_5769,N_2708,N_241);
or U5770 (N_5770,N_409,N_1661);
and U5771 (N_5771,N_2389,N_4623);
and U5772 (N_5772,N_4366,N_21);
and U5773 (N_5773,N_3573,N_1215);
or U5774 (N_5774,N_4153,N_1835);
nor U5775 (N_5775,N_4415,N_2349);
nand U5776 (N_5776,N_2054,N_4061);
nand U5777 (N_5777,N_1996,N_3859);
or U5778 (N_5778,N_2590,N_4276);
and U5779 (N_5779,N_2102,N_2123);
nor U5780 (N_5780,N_3537,N_2031);
or U5781 (N_5781,N_1271,N_1118);
or U5782 (N_5782,N_75,N_2808);
nand U5783 (N_5783,N_3588,N_4957);
nor U5784 (N_5784,N_2608,N_2423);
nand U5785 (N_5785,N_4648,N_4321);
or U5786 (N_5786,N_998,N_2089);
nor U5787 (N_5787,N_697,N_4965);
nor U5788 (N_5788,N_1995,N_2561);
nand U5789 (N_5789,N_4070,N_2096);
nor U5790 (N_5790,N_3070,N_3979);
nor U5791 (N_5791,N_1680,N_572);
or U5792 (N_5792,N_93,N_1126);
and U5793 (N_5793,N_2756,N_1963);
nand U5794 (N_5794,N_2869,N_2070);
nor U5795 (N_5795,N_2218,N_3770);
or U5796 (N_5796,N_4247,N_2727);
or U5797 (N_5797,N_3001,N_4564);
nor U5798 (N_5798,N_801,N_798);
or U5799 (N_5799,N_2951,N_944);
and U5800 (N_5800,N_2235,N_2438);
or U5801 (N_5801,N_2290,N_731);
nor U5802 (N_5802,N_2952,N_3362);
or U5803 (N_5803,N_27,N_277);
nand U5804 (N_5804,N_2483,N_79);
nand U5805 (N_5805,N_782,N_530);
nand U5806 (N_5806,N_4354,N_918);
and U5807 (N_5807,N_820,N_4056);
or U5808 (N_5808,N_2146,N_4607);
and U5809 (N_5809,N_729,N_930);
nor U5810 (N_5810,N_2004,N_64);
nor U5811 (N_5811,N_3129,N_2597);
or U5812 (N_5812,N_1936,N_3816);
nor U5813 (N_5813,N_3254,N_2194);
nor U5814 (N_5814,N_460,N_4696);
nand U5815 (N_5815,N_2541,N_651);
or U5816 (N_5816,N_4316,N_2540);
nand U5817 (N_5817,N_3276,N_1239);
and U5818 (N_5818,N_4385,N_2690);
and U5819 (N_5819,N_4122,N_4062);
or U5820 (N_5820,N_1620,N_2909);
nand U5821 (N_5821,N_4298,N_267);
and U5822 (N_5822,N_2165,N_3243);
nor U5823 (N_5823,N_3856,N_571);
or U5824 (N_5824,N_4161,N_689);
and U5825 (N_5825,N_15,N_2376);
nor U5826 (N_5826,N_4903,N_4063);
nand U5827 (N_5827,N_2166,N_1559);
and U5828 (N_5828,N_4280,N_2018);
and U5829 (N_5829,N_599,N_3123);
nand U5830 (N_5830,N_4652,N_4032);
or U5831 (N_5831,N_356,N_4817);
nor U5832 (N_5832,N_4587,N_2277);
nor U5833 (N_5833,N_4234,N_4170);
or U5834 (N_5834,N_549,N_3506);
nand U5835 (N_5835,N_3778,N_4225);
nand U5836 (N_5836,N_1800,N_4521);
nand U5837 (N_5837,N_4422,N_4673);
nor U5838 (N_5838,N_4082,N_3757);
or U5839 (N_5839,N_1494,N_3508);
nor U5840 (N_5840,N_675,N_1003);
nand U5841 (N_5841,N_4449,N_2307);
nand U5842 (N_5842,N_4272,N_4158);
nand U5843 (N_5843,N_664,N_274);
or U5844 (N_5844,N_3101,N_2627);
xnor U5845 (N_5845,N_875,N_3107);
or U5846 (N_5846,N_1575,N_3561);
or U5847 (N_5847,N_4644,N_959);
nor U5848 (N_5848,N_161,N_1250);
and U5849 (N_5849,N_164,N_3166);
and U5850 (N_5850,N_2959,N_2828);
or U5851 (N_5851,N_3015,N_2682);
nor U5852 (N_5852,N_3777,N_4074);
or U5853 (N_5853,N_4676,N_275);
nor U5854 (N_5854,N_818,N_983);
and U5855 (N_5855,N_211,N_2319);
nor U5856 (N_5856,N_2732,N_1052);
xnor U5857 (N_5857,N_4828,N_2620);
or U5858 (N_5858,N_2399,N_1902);
or U5859 (N_5859,N_3248,N_3007);
nand U5860 (N_5860,N_442,N_4875);
nand U5861 (N_5861,N_4309,N_263);
nor U5862 (N_5862,N_2761,N_3412);
or U5863 (N_5863,N_4866,N_3056);
or U5864 (N_5864,N_1691,N_1805);
and U5865 (N_5865,N_2966,N_4897);
nor U5866 (N_5866,N_1399,N_1049);
nand U5867 (N_5867,N_552,N_4503);
and U5868 (N_5868,N_425,N_2364);
or U5869 (N_5869,N_4290,N_1977);
nand U5870 (N_5870,N_186,N_1842);
nand U5871 (N_5871,N_1354,N_4014);
or U5872 (N_5872,N_1455,N_4616);
or U5873 (N_5873,N_1667,N_4534);
nor U5874 (N_5874,N_740,N_1853);
and U5875 (N_5875,N_3135,N_4731);
nand U5876 (N_5876,N_2823,N_2829);
nor U5877 (N_5877,N_536,N_1709);
or U5878 (N_5878,N_3260,N_642);
and U5879 (N_5879,N_3747,N_3925);
nand U5880 (N_5880,N_384,N_2271);
nor U5881 (N_5881,N_4779,N_3784);
and U5882 (N_5882,N_3741,N_112);
nor U5883 (N_5883,N_3787,N_2404);
nand U5884 (N_5884,N_1945,N_1560);
and U5885 (N_5885,N_1148,N_3186);
and U5886 (N_5886,N_1883,N_366);
and U5887 (N_5887,N_2361,N_548);
nand U5888 (N_5888,N_4183,N_4661);
nor U5889 (N_5889,N_2175,N_3083);
nor U5890 (N_5890,N_2599,N_3241);
or U5891 (N_5891,N_1087,N_2705);
nor U5892 (N_5892,N_382,N_2379);
or U5893 (N_5893,N_3526,N_4576);
nor U5894 (N_5894,N_662,N_50);
nor U5895 (N_5895,N_1648,N_1579);
or U5896 (N_5896,N_419,N_4443);
nand U5897 (N_5897,N_388,N_779);
nand U5898 (N_5898,N_2105,N_3108);
or U5899 (N_5899,N_3440,N_1774);
nor U5900 (N_5900,N_3735,N_343);
or U5901 (N_5901,N_373,N_4105);
nor U5902 (N_5902,N_3468,N_311);
nand U5903 (N_5903,N_1177,N_1737);
nor U5904 (N_5904,N_3872,N_764);
and U5905 (N_5905,N_830,N_632);
and U5906 (N_5906,N_1806,N_4737);
and U5907 (N_5907,N_1139,N_3103);
nand U5908 (N_5908,N_1856,N_2144);
and U5909 (N_5909,N_3656,N_3080);
or U5910 (N_5910,N_2881,N_1380);
or U5911 (N_5911,N_2558,N_4873);
or U5912 (N_5912,N_3946,N_1637);
or U5913 (N_5913,N_805,N_1302);
nor U5914 (N_5914,N_2739,N_2633);
and U5915 (N_5915,N_519,N_2510);
nor U5916 (N_5916,N_3480,N_1132);
nor U5917 (N_5917,N_4719,N_4102);
nor U5918 (N_5918,N_4477,N_3646);
nand U5919 (N_5919,N_4399,N_2547);
nor U5920 (N_5920,N_2870,N_4249);
nor U5921 (N_5921,N_2787,N_3729);
nor U5922 (N_5922,N_1900,N_4381);
or U5923 (N_5923,N_703,N_3833);
nand U5924 (N_5924,N_3239,N_484);
and U5925 (N_5925,N_2820,N_600);
or U5926 (N_5926,N_3091,N_2119);
and U5927 (N_5927,N_3040,N_463);
nand U5928 (N_5928,N_4959,N_4044);
and U5929 (N_5929,N_7,N_2796);
or U5930 (N_5930,N_2206,N_2672);
nand U5931 (N_5931,N_4184,N_2181);
and U5932 (N_5932,N_4406,N_3006);
nor U5933 (N_5933,N_2087,N_1129);
or U5934 (N_5934,N_1236,N_2814);
and U5935 (N_5935,N_1590,N_4928);
and U5936 (N_5936,N_3244,N_1708);
nor U5937 (N_5937,N_2233,N_3323);
nor U5938 (N_5938,N_2917,N_3516);
nor U5939 (N_5939,N_3705,N_3132);
or U5940 (N_5940,N_4837,N_2152);
nand U5941 (N_5941,N_362,N_305);
xnor U5942 (N_5942,N_434,N_1293);
and U5943 (N_5943,N_489,N_1804);
or U5944 (N_5944,N_4736,N_2647);
nand U5945 (N_5945,N_3529,N_16);
and U5946 (N_5946,N_2830,N_22);
or U5947 (N_5947,N_3809,N_73);
or U5948 (N_5948,N_2256,N_3199);
or U5949 (N_5949,N_4525,N_4275);
or U5950 (N_5950,N_1462,N_443);
nand U5951 (N_5951,N_2086,N_1454);
and U5952 (N_5952,N_4829,N_4058);
or U5953 (N_5953,N_1153,N_3941);
nor U5954 (N_5954,N_3268,N_1044);
nand U5955 (N_5955,N_4336,N_3483);
and U5956 (N_5956,N_916,N_1662);
nor U5957 (N_5957,N_4304,N_606);
or U5958 (N_5958,N_2956,N_3616);
nand U5959 (N_5959,N_3961,N_4147);
or U5960 (N_5960,N_584,N_1154);
or U5961 (N_5961,N_2045,N_1904);
and U5962 (N_5962,N_1663,N_9);
or U5963 (N_5963,N_2833,N_3479);
nor U5964 (N_5964,N_1127,N_207);
nand U5965 (N_5965,N_578,N_620);
nor U5966 (N_5966,N_1690,N_673);
nand U5967 (N_5967,N_656,N_226);
nand U5968 (N_5968,N_3592,N_2914);
nand U5969 (N_5969,N_2397,N_4455);
nor U5970 (N_5970,N_2287,N_4417);
and U5971 (N_5971,N_973,N_2071);
or U5972 (N_5972,N_4949,N_3161);
and U5973 (N_5973,N_322,N_3086);
nor U5974 (N_5974,N_1855,N_2635);
and U5975 (N_5975,N_3310,N_3654);
and U5976 (N_5976,N_4040,N_4267);
nor U5977 (N_5977,N_1808,N_523);
and U5978 (N_5978,N_2150,N_4005);
nand U5979 (N_5979,N_1075,N_3031);
and U5980 (N_5980,N_4744,N_4042);
or U5981 (N_5981,N_3032,N_2606);
nor U5982 (N_5982,N_2367,N_3112);
nand U5983 (N_5983,N_1788,N_3068);
or U5984 (N_5984,N_1457,N_2273);
and U5985 (N_5985,N_3334,N_4227);
or U5986 (N_5986,N_3840,N_2655);
nor U5987 (N_5987,N_693,N_2320);
nand U5988 (N_5988,N_3283,N_1582);
nor U5989 (N_5989,N_104,N_4973);
nor U5990 (N_5990,N_4915,N_52);
nand U5991 (N_5991,N_2879,N_1028);
and U5992 (N_5992,N_3496,N_1393);
nor U5993 (N_5993,N_4912,N_2050);
nor U5994 (N_5994,N_1611,N_2697);
and U5995 (N_5995,N_1278,N_1864);
and U5996 (N_5996,N_2346,N_4363);
nor U5997 (N_5997,N_2244,N_3974);
or U5998 (N_5998,N_2526,N_1142);
nand U5999 (N_5999,N_756,N_269);
nand U6000 (N_6000,N_4505,N_2372);
and U6001 (N_6001,N_4498,N_1352);
nor U6002 (N_6002,N_2258,N_4236);
nor U6003 (N_6003,N_3500,N_4143);
nor U6004 (N_6004,N_2491,N_4991);
or U6005 (N_6005,N_2960,N_1251);
or U6006 (N_6006,N_466,N_4502);
nor U6007 (N_6007,N_934,N_2037);
and U6008 (N_6008,N_3291,N_1202);
and U6009 (N_6009,N_4300,N_545);
or U6010 (N_6010,N_4514,N_245);
and U6011 (N_6011,N_2164,N_1768);
nor U6012 (N_6012,N_2509,N_256);
or U6013 (N_6013,N_2495,N_874);
nand U6014 (N_6014,N_2309,N_4009);
nor U6015 (N_6015,N_3363,N_2447);
or U6016 (N_6016,N_3430,N_4178);
or U6017 (N_6017,N_4918,N_2986);
nand U6018 (N_6018,N_1561,N_1622);
and U6019 (N_6019,N_1789,N_2424);
and U6020 (N_6020,N_1178,N_3090);
nand U6021 (N_6021,N_1526,N_2689);
nor U6022 (N_6022,N_4287,N_3256);
and U6023 (N_6023,N_328,N_3299);
nor U6024 (N_6024,N_2099,N_4759);
nand U6025 (N_6025,N_146,N_4831);
xnor U6026 (N_6026,N_2589,N_1398);
nor U6027 (N_6027,N_2059,N_4185);
nor U6028 (N_6028,N_96,N_76);
nor U6029 (N_6029,N_893,N_3415);
nand U6030 (N_6030,N_2241,N_1869);
and U6031 (N_6031,N_817,N_3611);
nand U6032 (N_6032,N_2600,N_1492);
nor U6033 (N_6033,N_861,N_4433);
nand U6034 (N_6034,N_1038,N_889);
nor U6035 (N_6035,N_2962,N_2669);
nand U6036 (N_6036,N_2811,N_286);
nand U6037 (N_6037,N_3877,N_2893);
and U6038 (N_6038,N_1320,N_815);
nand U6039 (N_6039,N_1312,N_155);
and U6040 (N_6040,N_784,N_1476);
or U6041 (N_6041,N_3013,N_3760);
and U6042 (N_6042,N_4908,N_2199);
nand U6043 (N_6043,N_4209,N_2387);
nor U6044 (N_6044,N_2981,N_2716);
or U6045 (N_6045,N_2857,N_2516);
and U6046 (N_6046,N_3094,N_3867);
and U6047 (N_6047,N_949,N_4093);
nor U6048 (N_6048,N_1537,N_3366);
and U6049 (N_6049,N_562,N_2846);
and U6050 (N_6050,N_32,N_2612);
or U6051 (N_6051,N_3948,N_1786);
or U6052 (N_6052,N_1478,N_639);
nor U6053 (N_6053,N_2849,N_4735);
or U6054 (N_6054,N_223,N_2316);
nor U6055 (N_6055,N_2341,N_1179);
or U6056 (N_6056,N_3715,N_4157);
and U6057 (N_6057,N_972,N_1892);
or U6058 (N_6058,N_3205,N_2211);
nand U6059 (N_6059,N_4702,N_3226);
or U6060 (N_6060,N_3521,N_4379);
nand U6061 (N_6061,N_4729,N_708);
xnor U6062 (N_6062,N_712,N_4896);
or U6063 (N_6063,N_4840,N_2064);
or U6064 (N_6064,N_4666,N_3772);
or U6065 (N_6065,N_4751,N_2294);
nand U6066 (N_6066,N_3587,N_3264);
xnor U6067 (N_6067,N_527,N_4947);
or U6068 (N_6068,N_4626,N_243);
and U6069 (N_6069,N_4192,N_564);
nor U6070 (N_6070,N_494,N_74);
or U6071 (N_6071,N_1758,N_44);
nand U6072 (N_6072,N_3074,N_2907);
nor U6073 (N_6073,N_2240,N_3113);
or U6074 (N_6074,N_3805,N_904);
and U6075 (N_6075,N_2444,N_2609);
nor U6076 (N_6076,N_349,N_3392);
and U6077 (N_6077,N_1927,N_2642);
nand U6078 (N_6078,N_383,N_3272);
nand U6079 (N_6079,N_118,N_556);
and U6080 (N_6080,N_4913,N_3509);
or U6081 (N_6081,N_1261,N_309);
xor U6082 (N_6082,N_732,N_4109);
nor U6083 (N_6083,N_528,N_1410);
nand U6084 (N_6084,N_2286,N_4773);
and U6085 (N_6085,N_4114,N_880);
nand U6086 (N_6086,N_209,N_3082);
or U6087 (N_6087,N_165,N_2762);
or U6088 (N_6088,N_503,N_588);
and U6089 (N_6089,N_3535,N_1505);
nand U6090 (N_6090,N_1909,N_1525);
nand U6091 (N_6091,N_4710,N_4935);
or U6092 (N_6092,N_3548,N_4116);
and U6093 (N_6093,N_450,N_4092);
or U6094 (N_6094,N_643,N_1920);
nand U6095 (N_6095,N_976,N_4899);
or U6096 (N_6096,N_2692,N_3634);
xnor U6097 (N_6097,N_2412,N_467);
or U6098 (N_6098,N_257,N_1500);
and U6099 (N_6099,N_1071,N_71);
or U6100 (N_6100,N_4584,N_1425);
or U6101 (N_6101,N_3955,N_3296);
nand U6102 (N_6102,N_2468,N_4128);
or U6103 (N_6103,N_4463,N_2153);
or U6104 (N_6104,N_3929,N_507);
nor U6105 (N_6105,N_4615,N_2676);
nand U6106 (N_6106,N_2257,N_534);
or U6107 (N_6107,N_4750,N_4743);
or U6108 (N_6108,N_2437,N_2551);
or U6109 (N_6109,N_537,N_2795);
or U6110 (N_6110,N_1096,N_4491);
and U6111 (N_6111,N_1825,N_1130);
and U6112 (N_6112,N_622,N_4012);
and U6113 (N_6113,N_4739,N_3002);
nand U6114 (N_6114,N_1029,N_372);
or U6115 (N_6115,N_3281,N_4504);
nor U6116 (N_6116,N_4547,N_1207);
nor U6117 (N_6117,N_26,N_2997);
nor U6118 (N_6118,N_3938,N_702);
or U6119 (N_6119,N_3189,N_4418);
xor U6120 (N_6120,N_3275,N_4948);
nor U6121 (N_6121,N_1591,N_1381);
nor U6122 (N_6122,N_1326,N_4567);
nor U6123 (N_6123,N_1895,N_795);
nand U6124 (N_6124,N_2075,N_3909);
or U6125 (N_6125,N_1687,N_63);
or U6126 (N_6126,N_879,N_2899);
or U6127 (N_6127,N_2098,N_1300);
and U6128 (N_6128,N_1057,N_1497);
or U6129 (N_6129,N_4674,N_2176);
or U6130 (N_6130,N_3846,N_2982);
or U6131 (N_6131,N_4663,N_4841);
and U6132 (N_6132,N_3984,N_2388);
nor U6133 (N_6133,N_2501,N_631);
nand U6134 (N_6134,N_4511,N_3492);
nand U6135 (N_6135,N_2025,N_2127);
and U6136 (N_6136,N_4358,N_1333);
and U6137 (N_6137,N_3118,N_4317);
nor U6138 (N_6138,N_1626,N_414);
or U6139 (N_6139,N_1348,N_1585);
and U6140 (N_6140,N_4728,N_2464);
and U6141 (N_6141,N_690,N_2624);
and U6142 (N_6142,N_1159,N_4944);
nor U6143 (N_6143,N_1612,N_3340);
nand U6144 (N_6144,N_1538,N_4059);
and U6145 (N_6145,N_2473,N_3126);
nor U6146 (N_6146,N_159,N_1743);
or U6147 (N_6147,N_1055,N_2460);
nor U6148 (N_6148,N_3345,N_210);
or U6149 (N_6149,N_2878,N_3552);
and U6150 (N_6150,N_4163,N_3339);
and U6151 (N_6151,N_2276,N_3233);
nor U6152 (N_6152,N_1368,N_1653);
and U6153 (N_6153,N_3522,N_716);
nand U6154 (N_6154,N_2443,N_4064);
nor U6155 (N_6155,N_3761,N_3360);
and U6156 (N_6156,N_4154,N_4326);
nand U6157 (N_6157,N_1997,N_4952);
or U6158 (N_6158,N_4186,N_3837);
nor U6159 (N_6159,N_3196,N_459);
or U6160 (N_6160,N_2403,N_324);
nor U6161 (N_6161,N_2434,N_4258);
nor U6162 (N_6162,N_3265,N_1823);
and U6163 (N_6163,N_1218,N_928);
nor U6164 (N_6164,N_2002,N_4887);
and U6165 (N_6165,N_1696,N_2538);
or U6166 (N_6166,N_280,N_222);
and U6167 (N_6167,N_3462,N_3721);
nor U6168 (N_6168,N_289,N_1321);
nor U6169 (N_6169,N_1941,N_1751);
and U6170 (N_6170,N_1489,N_2450);
and U6171 (N_6171,N_3850,N_2623);
or U6172 (N_6172,N_1031,N_1107);
nor U6173 (N_6173,N_4000,N_2517);
or U6174 (N_6174,N_1423,N_317);
or U6175 (N_6175,N_1198,N_2393);
xnor U6176 (N_6176,N_872,N_436);
or U6177 (N_6177,N_1349,N_4785);
or U6178 (N_6178,N_261,N_1641);
nand U6179 (N_6179,N_3606,N_3554);
or U6180 (N_6180,N_2885,N_822);
and U6181 (N_6181,N_1122,N_447);
or U6182 (N_6182,N_3289,N_1594);
nor U6183 (N_6183,N_3855,N_3211);
xor U6184 (N_6184,N_3713,N_2457);
nand U6185 (N_6185,N_4337,N_1436);
nand U6186 (N_6186,N_2924,N_2858);
and U6187 (N_6187,N_649,N_2836);
nor U6188 (N_6188,N_1843,N_612);
and U6189 (N_6189,N_1809,N_2901);
or U6190 (N_6190,N_172,N_283);
and U6191 (N_6191,N_3815,N_894);
nand U6192 (N_6192,N_825,N_4986);
nand U6193 (N_6193,N_2532,N_354);
and U6194 (N_6194,N_3252,N_4119);
and U6195 (N_6195,N_1262,N_833);
and U6196 (N_6196,N_4815,N_917);
nor U6197 (N_6197,N_85,N_4253);
nor U6198 (N_6198,N_2567,N_1067);
nor U6199 (N_6199,N_4423,N_1310);
and U6200 (N_6200,N_3728,N_4967);
or U6201 (N_6201,N_2463,N_4169);
and U6202 (N_6202,N_421,N_2522);
or U6203 (N_6203,N_2587,N_979);
nor U6204 (N_6204,N_100,N_1385);
nand U6205 (N_6205,N_4195,N_405);
nor U6206 (N_6206,N_725,N_1970);
nand U6207 (N_6207,N_1729,N_3140);
nor U6208 (N_6208,N_757,N_3644);
or U6209 (N_6209,N_3089,N_870);
nand U6210 (N_6210,N_188,N_429);
or U6211 (N_6211,N_2994,N_2910);
xnor U6212 (N_6212,N_285,N_688);
nor U6213 (N_6213,N_3804,N_40);
and U6214 (N_6214,N_2201,N_4437);
and U6215 (N_6215,N_4493,N_4212);
and U6216 (N_6216,N_471,N_2634);
nor U6217 (N_6217,N_1851,N_2384);
nand U6218 (N_6218,N_2124,N_2533);
nor U6219 (N_6219,N_4101,N_1346);
nor U6220 (N_6220,N_1450,N_2523);
nand U6221 (N_6221,N_2014,N_3907);
nor U6222 (N_6222,N_4760,N_391);
nand U6223 (N_6223,N_2750,N_8);
nor U6224 (N_6224,N_3214,N_952);
nand U6225 (N_6225,N_2159,N_3049);
nor U6226 (N_6226,N_2168,N_191);
nand U6227 (N_6227,N_4460,N_687);
or U6228 (N_6228,N_344,N_3125);
and U6229 (N_6229,N_4485,N_1839);
nor U6230 (N_6230,N_2359,N_4167);
and U6231 (N_6231,N_4895,N_1007);
nand U6232 (N_6232,N_4802,N_1722);
or U6233 (N_6233,N_3743,N_1181);
and U6234 (N_6234,N_3318,N_1374);
and U6235 (N_6235,N_1787,N_1099);
or U6236 (N_6236,N_3882,N_3742);
and U6237 (N_6237,N_2782,N_986);
or U6238 (N_6238,N_2696,N_2117);
nand U6239 (N_6239,N_4768,N_117);
or U6240 (N_6240,N_4910,N_509);
nor U6241 (N_6241,N_966,N_4783);
and U6242 (N_6242,N_3229,N_2270);
nand U6243 (N_6243,N_619,N_2777);
and U6244 (N_6244,N_4228,N_3076);
and U6245 (N_6245,N_3262,N_746);
nor U6246 (N_6246,N_905,N_3640);
nor U6247 (N_6247,N_3810,N_169);
nor U6248 (N_6248,N_1232,N_1982);
xnor U6249 (N_6249,N_3525,N_295);
and U6250 (N_6250,N_4252,N_3405);
and U6251 (N_6251,N_4692,N_1878);
nand U6252 (N_6252,N_359,N_3012);
nand U6253 (N_6253,N_4645,N_2877);
or U6254 (N_6254,N_3763,N_1430);
or U6255 (N_6255,N_914,N_437);
and U6256 (N_6256,N_306,N_1253);
and U6257 (N_6257,N_1608,N_342);
and U6258 (N_6258,N_4905,N_327);
or U6259 (N_6259,N_867,N_3030);
and U6260 (N_6260,N_35,N_2847);
nand U6261 (N_6261,N_3371,N_1004);
nand U6262 (N_6262,N_2780,N_2062);
and U6263 (N_6263,N_684,N_4229);
nor U6264 (N_6264,N_745,N_1688);
nor U6265 (N_6265,N_2157,N_3681);
or U6266 (N_6266,N_181,N_2482);
or U6267 (N_6267,N_124,N_4555);
or U6268 (N_6268,N_4282,N_3328);
nor U6269 (N_6269,N_1676,N_1140);
and U6270 (N_6270,N_4135,N_4892);
and U6271 (N_6271,N_4740,N_1382);
nor U6272 (N_6272,N_2613,N_3159);
nand U6273 (N_6273,N_4717,N_2180);
nand U6274 (N_6274,N_4794,N_3674);
nor U6275 (N_6275,N_1358,N_978);
and U6276 (N_6276,N_1628,N_1471);
nand U6277 (N_6277,N_1801,N_1010);
nand U6278 (N_6278,N_2873,N_479);
nor U6279 (N_6279,N_714,N_4372);
nand U6280 (N_6280,N_4565,N_2221);
and U6281 (N_6281,N_2420,N_1411);
nor U6282 (N_6282,N_259,N_3667);
nand U6283 (N_6283,N_2042,N_2339);
nand U6284 (N_6284,N_3963,N_589);
nand U6285 (N_6285,N_848,N_3446);
or U6286 (N_6286,N_3322,N_381);
and U6287 (N_6287,N_778,N_1331);
nor U6288 (N_6288,N_2485,N_3454);
or U6289 (N_6289,N_183,N_36);
nand U6290 (N_6290,N_2964,N_2602);
and U6291 (N_6291,N_2701,N_2056);
or U6292 (N_6292,N_3329,N_3010);
or U6293 (N_6293,N_4771,N_2630);
and U6294 (N_6294,N_2184,N_4683);
or U6295 (N_6295,N_2260,N_2266);
or U6296 (N_6296,N_4950,N_1674);
xor U6297 (N_6297,N_29,N_4784);
and U6298 (N_6298,N_370,N_3507);
or U6299 (N_6299,N_3369,N_214);
and U6300 (N_6300,N_2706,N_254);
nand U6301 (N_6301,N_83,N_3274);
nand U6302 (N_6302,N_539,N_616);
nor U6303 (N_6303,N_2382,N_2622);
nand U6304 (N_6304,N_1447,N_427);
or U6305 (N_6305,N_1725,N_3584);
nor U6306 (N_6306,N_2207,N_948);
and U6307 (N_6307,N_1599,N_1089);
and U6308 (N_6308,N_2351,N_3830);
and U6309 (N_6309,N_1817,N_2267);
nand U6310 (N_6310,N_2496,N_3638);
or U6311 (N_6311,N_709,N_1158);
and U6312 (N_6312,N_1669,N_4015);
or U6313 (N_6313,N_2500,N_2317);
nor U6314 (N_6314,N_970,N_404);
nand U6315 (N_6315,N_838,N_4668);
nand U6316 (N_6316,N_855,N_590);
nand U6317 (N_6317,N_1583,N_3204);
nand U6318 (N_6318,N_2718,N_127);
nand U6319 (N_6319,N_1917,N_4461);
nand U6320 (N_6320,N_2653,N_318);
nor U6321 (N_6321,N_3207,N_1670);
nand U6322 (N_6322,N_126,N_615);
nand U6323 (N_6323,N_353,N_1887);
nand U6324 (N_6324,N_705,N_3338);
or U6325 (N_6325,N_3059,N_3671);
and U6326 (N_6326,N_2217,N_1121);
or U6327 (N_6327,N_638,N_67);
or U6328 (N_6328,N_1111,N_3960);
nand U6329 (N_6329,N_2392,N_3365);
and U6330 (N_6330,N_1879,N_1588);
nor U6331 (N_6331,N_2442,N_3145);
nand U6332 (N_6332,N_2462,N_1016);
and U6333 (N_6333,N_3714,N_1810);
and U6334 (N_6334,N_1619,N_4375);
or U6335 (N_6335,N_464,N_130);
or U6336 (N_6336,N_2456,N_4240);
nand U6337 (N_6337,N_28,N_706);
and U6338 (N_6338,N_1424,N_2407);
nand U6339 (N_6339,N_1054,N_2886);
nor U6340 (N_6340,N_2904,N_4224);
nor U6341 (N_6341,N_313,N_3206);
and U6342 (N_6342,N_1020,N_4715);
or U6343 (N_6343,N_3081,N_3991);
and U6344 (N_6344,N_4099,N_2375);
nor U6345 (N_6345,N_701,N_3811);
and U6346 (N_6346,N_1656,N_4594);
or U6347 (N_6347,N_2334,N_882);
nand U6348 (N_6348,N_141,N_1655);
and U6349 (N_6349,N_608,N_3541);
nand U6350 (N_6350,N_2198,N_4876);
or U6351 (N_6351,N_273,N_1633);
or U6352 (N_6352,N_2512,N_1606);
nor U6353 (N_6353,N_4084,N_3105);
nor U6354 (N_6354,N_4481,N_184);
nor U6355 (N_6355,N_2189,N_2576);
nor U6356 (N_6356,N_3857,N_4489);
or U6357 (N_6357,N_3879,N_2704);
or U6358 (N_6358,N_4329,N_3297);
or U6359 (N_6359,N_1593,N_2683);
xnor U6360 (N_6360,N_735,N_1387);
and U6361 (N_6361,N_3472,N_4242);
or U6362 (N_6362,N_4980,N_1985);
nand U6363 (N_6363,N_4561,N_990);
or U6364 (N_6364,N_524,N_752);
and U6365 (N_6365,N_2055,N_4861);
or U6366 (N_6366,N_4976,N_3900);
nand U6367 (N_6367,N_4960,N_54);
and U6368 (N_6368,N_3785,N_72);
and U6369 (N_6369,N_515,N_672);
and U6370 (N_6370,N_2354,N_1245);
or U6371 (N_6371,N_108,N_1794);
or U6372 (N_6372,N_618,N_4796);
or U6373 (N_6373,N_230,N_3831);
or U6374 (N_6374,N_4811,N_4155);
and U6375 (N_6375,N_1347,N_4050);
nor U6376 (N_6376,N_1449,N_4412);
nand U6377 (N_6377,N_3367,N_4395);
or U6378 (N_6378,N_1463,N_3524);
or U6379 (N_6379,N_1750,N_829);
and U6380 (N_6380,N_2580,N_2737);
and U6381 (N_6381,N_3807,N_1584);
nor U6382 (N_6382,N_4302,N_4277);
or U6383 (N_6383,N_3429,N_726);
nor U6384 (N_6384,N_430,N_4003);
or U6385 (N_6385,N_4761,N_1924);
nand U6386 (N_6386,N_2250,N_1930);
or U6387 (N_6387,N_2077,N_1255);
or U6388 (N_6388,N_3324,N_4958);
or U6389 (N_6389,N_4328,N_2731);
nor U6390 (N_6390,N_2046,N_287);
or U6391 (N_6391,N_1831,N_2554);
and U6392 (N_6392,N_1521,N_3357);
nor U6393 (N_6393,N_4138,N_4126);
and U6394 (N_6394,N_2965,N_4672);
nor U6395 (N_6395,N_4369,N_68);
nand U6396 (N_6396,N_4076,N_1793);
nand U6397 (N_6397,N_2029,N_730);
nor U6398 (N_6398,N_2970,N_4968);
or U6399 (N_6399,N_3813,N_4589);
nand U6400 (N_6400,N_3720,N_2335);
nor U6401 (N_6401,N_3791,N_1316);
or U6402 (N_6402,N_1554,N_1849);
nand U6403 (N_6403,N_3567,N_823);
nor U6404 (N_6404,N_1652,N_2729);
nor U6405 (N_6405,N_3072,N_2205);
or U6406 (N_6406,N_4579,N_751);
nor U6407 (N_6407,N_389,N_2649);
nand U6408 (N_6408,N_2688,N_1700);
and U6409 (N_6409,N_491,N_278);
nand U6410 (N_6410,N_3234,N_145);
nand U6411 (N_6411,N_1629,N_614);
nand U6412 (N_6412,N_4047,N_2990);
or U6413 (N_6413,N_2856,N_3269);
nand U6414 (N_6414,N_2433,N_2057);
nor U6415 (N_6415,N_919,N_4554);
and U6416 (N_6416,N_511,N_1442);
and U6417 (N_6417,N_1979,N_4603);
or U6418 (N_6418,N_3625,N_2852);
or U6419 (N_6419,N_1110,N_4962);
nor U6420 (N_6420,N_2082,N_3880);
nor U6421 (N_6421,N_2837,N_1795);
or U6422 (N_6422,N_4430,N_98);
nor U6423 (N_6423,N_2925,N_3009);
and U6424 (N_6424,N_4305,N_3143);
and U6425 (N_6425,N_3666,N_2506);
and U6426 (N_6426,N_1120,N_3435);
nand U6427 (N_6427,N_2374,N_416);
nand U6428 (N_6428,N_1304,N_3942);
and U6429 (N_6429,N_1943,N_1534);
nor U6430 (N_6430,N_4004,N_3795);
nor U6431 (N_6431,N_4289,N_1654);
and U6432 (N_6432,N_3691,N_461);
nand U6433 (N_6433,N_4597,N_3569);
nor U6434 (N_6434,N_3740,N_1414);
or U6435 (N_6435,N_1039,N_2333);
nor U6436 (N_6436,N_1893,N_4614);
nor U6437 (N_6437,N_4254,N_4953);
nand U6438 (N_6438,N_2730,N_1167);
nand U6439 (N_6439,N_3799,N_4860);
and U6440 (N_6440,N_1440,N_1546);
or U6441 (N_6441,N_4680,N_3379);
or U6442 (N_6442,N_4100,N_2162);
nand U6443 (N_6443,N_3505,N_3997);
or U6444 (N_6444,N_248,N_546);
nor U6445 (N_6445,N_4943,N_4714);
or U6446 (N_6446,N_3202,N_2274);
and U6447 (N_6447,N_1765,N_350);
nand U6448 (N_6448,N_282,N_102);
nand U6449 (N_6449,N_1531,N_4469);
and U6450 (N_6450,N_78,N_4595);
or U6451 (N_6451,N_1536,N_481);
and U6452 (N_6452,N_412,N_1268);
and U6453 (N_6453,N_2115,N_2264);
nor U6454 (N_6454,N_1931,N_3116);
or U6455 (N_6455,N_4834,N_3983);
or U6456 (N_6456,N_962,N_1475);
nand U6457 (N_6457,N_2472,N_2663);
or U6458 (N_6458,N_4226,N_1673);
and U6459 (N_6459,N_4146,N_767);
and U6460 (N_6460,N_3752,N_41);
nor U6461 (N_6461,N_2719,N_3737);
and U6462 (N_6462,N_2831,N_2936);
nor U6463 (N_6463,N_3484,N_4931);
and U6464 (N_6464,N_3796,N_432);
nand U6465 (N_6465,N_4095,N_4177);
or U6466 (N_6466,N_1477,N_1490);
nand U6467 (N_6467,N_1916,N_1976);
nand U6468 (N_6468,N_4073,N_60);
nor U6469 (N_6469,N_2755,N_1413);
nor U6470 (N_6470,N_1519,N_4859);
nor U6471 (N_6471,N_4516,N_680);
or U6472 (N_6472,N_3146,N_2161);
or U6473 (N_6473,N_3037,N_3399);
or U6474 (N_6474,N_398,N_3246);
nand U6475 (N_6475,N_2769,N_3597);
or U6476 (N_6476,N_1874,N_1091);
nand U6477 (N_6477,N_4356,N_1947);
nand U6478 (N_6478,N_490,N_2228);
nor U6479 (N_6479,N_410,N_522);
nor U6480 (N_6480,N_1383,N_3585);
nand U6481 (N_6481,N_105,N_3046);
nand U6482 (N_6482,N_835,N_800);
or U6483 (N_6483,N_1518,N_3774);
or U6484 (N_6484,N_1384,N_520);
and U6485 (N_6485,N_4149,N_12);
nor U6486 (N_6486,N_3327,N_3649);
or U6487 (N_6487,N_1051,N_3519);
nor U6488 (N_6488,N_2640,N_4371);
nand U6489 (N_6489,N_3213,N_1870);
nand U6490 (N_6490,N_2210,N_1980);
nor U6491 (N_6491,N_2657,N_4535);
nand U6492 (N_6492,N_4532,N_2585);
xor U6493 (N_6493,N_1992,N_2984);
and U6494 (N_6494,N_4013,N_3188);
nor U6495 (N_6495,N_1905,N_1280);
nor U6496 (N_6496,N_3972,N_4164);
and U6497 (N_6497,N_759,N_2125);
xnor U6498 (N_6498,N_4639,N_3675);
nand U6499 (N_6499,N_1114,N_3154);
nand U6500 (N_6500,N_4140,N_985);
xor U6501 (N_6501,N_3175,N_2116);
or U6502 (N_6502,N_3893,N_2154);
and U6503 (N_6503,N_333,N_3999);
and U6504 (N_6504,N_2301,N_3098);
nor U6505 (N_6505,N_1802,N_789);
or U6506 (N_6506,N_3306,N_819);
nor U6507 (N_6507,N_1618,N_2571);
or U6508 (N_6508,N_3294,N_3444);
and U6509 (N_6509,N_365,N_2895);
or U6510 (N_6510,N_1866,N_1875);
nand U6511 (N_6511,N_3026,N_451);
nand U6512 (N_6512,N_1613,N_4933);
nor U6513 (N_6513,N_717,N_2712);
or U6514 (N_6514,N_2378,N_396);
nor U6515 (N_6515,N_4319,N_3843);
or U6516 (N_6516,N_190,N_3557);
and U6517 (N_6517,N_1859,N_17);
and U6518 (N_6518,N_4907,N_1865);
nor U6519 (N_6519,N_2278,N_1141);
or U6520 (N_6520,N_4407,N_1209);
nor U6521 (N_6521,N_2825,N_2671);
nor U6522 (N_6522,N_1601,N_2848);
nor U6523 (N_6523,N_4278,N_1291);
xor U6524 (N_6524,N_2044,N_2114);
nor U6525 (N_6525,N_1257,N_1200);
nand U6526 (N_6526,N_1324,N_4593);
nor U6527 (N_6527,N_569,N_1697);
nand U6528 (N_6528,N_4347,N_3670);
and U6529 (N_6529,N_435,N_4451);
nand U6530 (N_6530,N_2838,N_1035);
nand U6531 (N_6531,N_603,N_2303);
nor U6532 (N_6532,N_4243,N_1037);
nand U6533 (N_6533,N_174,N_724);
nor U6534 (N_6534,N_3455,N_1906);
nand U6535 (N_6535,N_3973,N_1435);
and U6536 (N_6536,N_3518,N_2698);
or U6537 (N_6537,N_2236,N_3990);
and U6538 (N_6538,N_1643,N_2797);
or U6539 (N_6539,N_4344,N_2553);
or U6540 (N_6540,N_1666,N_3280);
xnor U6541 (N_6541,N_62,N_2126);
nand U6542 (N_6542,N_4373,N_3927);
nor U6543 (N_6543,N_1736,N_2646);
nor U6544 (N_6544,N_2067,N_2466);
or U6545 (N_6545,N_2868,N_3935);
nor U6546 (N_6546,N_1993,N_4612);
and U6547 (N_6547,N_3102,N_3553);
nand U6548 (N_6548,N_4387,N_2441);
and U6549 (N_6549,N_2710,N_168);
or U6550 (N_6550,N_2400,N_497);
and U6551 (N_6551,N_4303,N_2288);
or U6552 (N_6552,N_850,N_1699);
or U6553 (N_6553,N_3321,N_3754);
nand U6554 (N_6554,N_4127,N_4725);
nor U6555 (N_6555,N_2488,N_922);
and U6556 (N_6556,N_1850,N_3277);
and U6557 (N_6557,N_1533,N_1128);
and U6558 (N_6558,N_2212,N_180);
nand U6559 (N_6559,N_1150,N_4757);
nor U6560 (N_6560,N_1098,N_2786);
or U6561 (N_6561,N_1367,N_2804);
nand U6562 (N_6562,N_2789,N_2897);
nor U6563 (N_6563,N_676,N_4591);
nand U6564 (N_6564,N_2380,N_4416);
or U6565 (N_6565,N_3285,N_2943);
nand U6566 (N_6566,N_1186,N_2262);
nor U6567 (N_6567,N_1448,N_2231);
or U6568 (N_6568,N_1283,N_4132);
or U6569 (N_6569,N_3899,N_1194);
and U6570 (N_6570,N_2048,N_3136);
and U6571 (N_6571,N_400,N_747);
nor U6572 (N_6572,N_4295,N_3887);
or U6573 (N_6573,N_4508,N_4332);
or U6574 (N_6574,N_1319,N_3407);
and U6575 (N_6575,N_711,N_3447);
nor U6576 (N_6576,N_428,N_3144);
and U6577 (N_6577,N_3096,N_1735);
nor U6578 (N_6578,N_260,N_4393);
nand U6579 (N_6579,N_2418,N_4069);
nand U6580 (N_6580,N_1277,N_4486);
and U6581 (N_6581,N_3157,N_1553);
nor U6582 (N_6582,N_4856,N_567);
or U6583 (N_6583,N_3378,N_770);
nor U6584 (N_6584,N_2835,N_3933);
and U6585 (N_6585,N_2991,N_630);
or U6586 (N_6586,N_4738,N_2570);
nand U6587 (N_6587,N_1377,N_154);
nand U6588 (N_6588,N_3970,N_3755);
nor U6589 (N_6589,N_1513,N_3460);
and U6590 (N_6590,N_2219,N_2736);
and U6591 (N_6591,N_1047,N_473);
or U6592 (N_6592,N_3424,N_2110);
nor U6593 (N_6593,N_856,N_2854);
nand U6594 (N_6594,N_913,N_109);
or U6595 (N_6595,N_3073,N_648);
nand U6596 (N_6596,N_2248,N_4438);
and U6597 (N_6597,N_1344,N_776);
nor U6598 (N_6598,N_337,N_2475);
nor U6599 (N_6599,N_3425,N_3905);
or U6600 (N_6600,N_2213,N_345);
or U6601 (N_6601,N_2643,N_4955);
or U6602 (N_6602,N_550,N_2950);
and U6603 (N_6603,N_1428,N_1777);
nand U6604 (N_6604,N_1726,N_591);
nand U6605 (N_6605,N_4600,N_836);
or U6606 (N_6606,N_1175,N_182);
and U6607 (N_6607,N_4851,N_4189);
xnor U6608 (N_6608,N_3041,N_323);
nand U6609 (N_6609,N_4699,N_3722);
nor U6610 (N_6610,N_4681,N_4396);
or U6611 (N_6611,N_3419,N_1088);
or U6612 (N_6612,N_4580,N_1350);
and U6613 (N_6613,N_20,N_3903);
nor U6614 (N_6614,N_2826,N_2355);
nand U6615 (N_6615,N_251,N_3558);
and U6616 (N_6616,N_2365,N_4231);
and U6617 (N_6617,N_2861,N_3608);
and U6618 (N_6618,N_587,N_2607);
nor U6619 (N_6619,N_2841,N_3894);
or U6620 (N_6620,N_4360,N_3881);
nor U6621 (N_6621,N_2155,N_1718);
nor U6622 (N_6622,N_4144,N_173);
or U6623 (N_6623,N_3717,N_1640);
and U6624 (N_6624,N_1373,N_2594);
nand U6625 (N_6625,N_2428,N_2358);
nor U6626 (N_6626,N_4932,N_3959);
and U6627 (N_6627,N_4902,N_3976);
nor U6628 (N_6628,N_1967,N_2340);
or U6629 (N_6629,N_1647,N_2695);
nor U6630 (N_6630,N_4998,N_2409);
or U6631 (N_6631,N_2562,N_1185);
nor U6632 (N_6632,N_4563,N_4115);
and U6633 (N_6633,N_2677,N_3711);
or U6634 (N_6634,N_3923,N_2973);
and U6635 (N_6635,N_4562,N_4857);
and U6636 (N_6636,N_1671,N_1405);
or U6637 (N_6637,N_580,N_4376);
nand U6638 (N_6638,N_1925,N_4495);
or U6639 (N_6639,N_1919,N_1076);
and U6640 (N_6640,N_3605,N_657);
or U6641 (N_6641,N_3969,N_991);
nor U6642 (N_6642,N_3630,N_3450);
or U6643 (N_6643,N_3058,N_1313);
and U6644 (N_6644,N_1818,N_2673);
nor U6645 (N_6645,N_3195,N_3065);
or U6646 (N_6646,N_3014,N_4357);
nor U6647 (N_6647,N_3225,N_2300);
or U6648 (N_6648,N_2614,N_2200);
nor U6649 (N_6649,N_4655,N_2947);
and U6650 (N_6650,N_3598,N_4239);
and U6651 (N_6651,N_4487,N_3874);
or U6652 (N_6652,N_193,N_4462);
and U6653 (N_6653,N_33,N_2776);
and U6654 (N_6654,N_3615,N_2226);
or U6655 (N_6655,N_1770,N_4781);
nor U6656 (N_6656,N_4476,N_2972);
nand U6657 (N_6657,N_3527,N_30);
or U6658 (N_6658,N_773,N_3576);
or U6659 (N_6659,N_4598,N_106);
or U6660 (N_6660,N_3121,N_1012);
nor U6661 (N_6661,N_2905,N_3641);
and U6662 (N_6662,N_4764,N_1083);
or U6663 (N_6663,N_3533,N_3470);
nor U6664 (N_6664,N_3025,N_4429);
and U6665 (N_6665,N_592,N_4874);
or U6666 (N_6666,N_4996,N_4724);
nor U6667 (N_6667,N_2298,N_780);
or U6668 (N_6668,N_4365,N_1747);
or U6669 (N_6669,N_3977,N_2190);
or U6670 (N_6670,N_4927,N_4118);
nor U6671 (N_6671,N_909,N_1816);
or U6672 (N_6672,N_788,N_2711);
or U6673 (N_6673,N_4330,N_1466);
and U6674 (N_6674,N_4842,N_4767);
nand U6675 (N_6675,N_19,N_2435);
nor U6676 (N_6676,N_4419,N_4071);
or U6677 (N_6677,N_4196,N_1329);
nand U6678 (N_6678,N_3192,N_3531);
nand U6679 (N_6679,N_2080,N_1503);
nand U6680 (N_6680,N_3176,N_2955);
nand U6681 (N_6681,N_3803,N_659);
nor U6682 (N_6682,N_1807,N_2039);
nor U6683 (N_6683,N_3687,N_2759);
or U6684 (N_6684,N_55,N_3538);
nand U6685 (N_6685,N_281,N_4575);
nand U6686 (N_6686,N_3725,N_1422);
nand U6687 (N_6687,N_4570,N_2774);
or U6688 (N_6688,N_2461,N_808);
nor U6689 (N_6689,N_4352,N_3523);
nand U6690 (N_6690,N_4348,N_4592);
or U6691 (N_6691,N_2377,N_110);
and U6692 (N_6692,N_314,N_3571);
and U6693 (N_6693,N_2350,N_4162);
nand U6694 (N_6694,N_3870,N_646);
or U6695 (N_6695,N_3697,N_1740);
nand U6696 (N_6696,N_2310,N_2845);
nand U6697 (N_6697,N_2822,N_1828);
and U6698 (N_6698,N_2735,N_3817);
nor U6699 (N_6699,N_975,N_2555);
and U6700 (N_6700,N_2139,N_1040);
nand U6701 (N_6701,N_4409,N_4775);
or U6702 (N_6702,N_4120,N_1686);
nor U6703 (N_6703,N_1950,N_814);
nand U6704 (N_6704,N_2686,N_4970);
and U6705 (N_6705,N_4467,N_2156);
nor U6706 (N_6706,N_170,N_2012);
nand U6707 (N_6707,N_4782,N_3685);
and U6708 (N_6708,N_1914,N_3684);
and U6709 (N_6709,N_4378,N_3043);
nor U6710 (N_6710,N_1117,N_4251);
xnor U6711 (N_6711,N_397,N_1439);
and U6712 (N_6712,N_158,N_1078);
and U6713 (N_6713,N_859,N_1119);
nor U6714 (N_6714,N_395,N_3510);
and U6715 (N_6715,N_989,N_2596);
nand U6716 (N_6716,N_38,N_832);
nand U6717 (N_6717,N_3546,N_4131);
xor U6718 (N_6718,N_1327,N_1913);
nor U6719 (N_6719,N_906,N_3895);
nor U6720 (N_6720,N_3215,N_4852);
nor U6721 (N_6721,N_3445,N_576);
xor U6722 (N_6722,N_3602,N_1308);
nor U6723 (N_6723,N_1814,N_2747);
and U6724 (N_6724,N_3305,N_422);
and U6725 (N_6725,N_3884,N_1957);
nor U6726 (N_6726,N_2693,N_4824);
or U6727 (N_6727,N_3610,N_3798);
nor U6728 (N_6728,N_1081,N_4325);
or U6729 (N_6729,N_4259,N_1767);
or U6730 (N_6730,N_3209,N_683);
xnor U6731 (N_6731,N_4638,N_1146);
and U6732 (N_6732,N_1929,N_1565);
and U6733 (N_6733,N_737,N_4691);
or U6734 (N_6734,N_4975,N_2431);
and U6735 (N_6735,N_4384,N_4799);
nor U6736 (N_6736,N_1246,N_3680);
and U6737 (N_6737,N_4609,N_1516);
or U6738 (N_6738,N_1757,N_938);
nand U6739 (N_6739,N_143,N_3992);
nand U6740 (N_6740,N_1627,N_14);
nand U6741 (N_6741,N_4318,N_3594);
and U6742 (N_6742,N_954,N_2748);
nand U6743 (N_6743,N_929,N_866);
and U6744 (N_6744,N_229,N_3698);
and U6745 (N_6745,N_1746,N_4596);
nor U6746 (N_6746,N_483,N_4886);
nand U6747 (N_6747,N_3115,N_167);
nand U6748 (N_6748,N_3106,N_3749);
or U6749 (N_6749,N_326,N_4777);
and U6750 (N_6750,N_1894,N_2398);
nand U6751 (N_6751,N_4922,N_1286);
nand U6752 (N_6752,N_3528,N_3731);
nand U6753 (N_6753,N_2345,N_4786);
or U6754 (N_6754,N_1206,N_4806);
and U6755 (N_6755,N_2177,N_1555);
and U6756 (N_6756,N_4458,N_2536);
nor U6757 (N_6757,N_4294,N_3926);
and U6758 (N_6758,N_3930,N_796);
nand U6759 (N_6759,N_501,N_3709);
and U6760 (N_6760,N_4519,N_3279);
nand U6761 (N_6761,N_3642,N_1101);
or U6762 (N_6762,N_4201,N_2816);
or U6763 (N_6763,N_4283,N_1396);
or U6764 (N_6764,N_3251,N_3794);
or U6765 (N_6765,N_3542,N_2479);
nand U6766 (N_6766,N_2006,N_4850);
nor U6767 (N_6767,N_581,N_4457);
nor U6768 (N_6768,N_3917,N_2076);
and U6769 (N_6769,N_3655,N_10);
and U6770 (N_6770,N_4772,N_3689);
and U6771 (N_6771,N_4898,N_1991);
nand U6772 (N_6772,N_3191,N_2521);
nand U6773 (N_6773,N_2072,N_2866);
nor U6774 (N_6774,N_2773,N_2969);
nand U6775 (N_6775,N_3301,N_2183);
or U6776 (N_6776,N_3036,N_2948);
and U6777 (N_6777,N_107,N_1515);
nand U6778 (N_6778,N_1779,N_360);
nor U6779 (N_6779,N_3099,N_1473);
nand U6780 (N_6780,N_3586,N_885);
or U6781 (N_6781,N_2440,N_4454);
nor U6782 (N_6782,N_4496,N_3534);
nor U6783 (N_6783,N_809,N_3497);
nand U6784 (N_6784,N_1940,N_95);
and U6785 (N_6785,N_2520,N_2368);
nor U6786 (N_6786,N_3964,N_2352);
nand U6787 (N_6787,N_1080,N_3420);
nand U6788 (N_6788,N_974,N_1260);
and U6789 (N_6789,N_4625,N_1702);
and U6790 (N_6790,N_2022,N_1946);
nor U6791 (N_6791,N_2940,N_4322);
or U6792 (N_6792,N_1460,N_2459);
nand U6793 (N_6793,N_2015,N_1461);
and U6794 (N_6794,N_2595,N_266);
and U6795 (N_6795,N_3617,N_1998);
and U6796 (N_6796,N_1783,N_1501);
nand U6797 (N_6797,N_1426,N_595);
and U6798 (N_6798,N_1105,N_4208);
nand U6799 (N_6799,N_2658,N_4533);
nor U6800 (N_6800,N_413,N_3451);
or U6801 (N_6801,N_2093,N_694);
nor U6802 (N_6802,N_4814,N_253);
nor U6803 (N_6803,N_1432,N_1713);
nand U6804 (N_6804,N_4220,N_3780);
nand U6805 (N_6805,N_3672,N_4809);
nand U6806 (N_6806,N_4920,N_2853);
or U6807 (N_6807,N_525,N_4805);
or U6808 (N_6808,N_1495,N_2369);
nor U6809 (N_6809,N_4599,N_2120);
nor U6810 (N_6810,N_4964,N_896);
nor U6811 (N_6811,N_2016,N_4553);
nor U6812 (N_6812,N_996,N_786);
or U6813 (N_6813,N_2193,N_271);
or U6814 (N_6814,N_4281,N_942);
and U6815 (N_6815,N_1073,N_1123);
nor U6816 (N_6816,N_363,N_199);
or U6817 (N_6817,N_216,N_3985);
and U6818 (N_6818,N_1989,N_3404);
nor U6819 (N_6819,N_332,N_24);
nand U6820 (N_6820,N_2136,N_3966);
nor U6821 (N_6821,N_2132,N_2035);
nor U6822 (N_6822,N_1248,N_1657);
or U6823 (N_6823,N_2839,N_4137);
nor U6824 (N_6824,N_977,N_3949);
or U6825 (N_6825,N_671,N_1014);
and U6826 (N_6826,N_2073,N_4869);
and U6827 (N_6827,N_2957,N_2104);
and U6828 (N_6828,N_2844,N_4141);
or U6829 (N_6829,N_1065,N_4174);
nand U6830 (N_6830,N_575,N_1235);
nor U6831 (N_6831,N_3120,N_1420);
and U6832 (N_6832,N_3467,N_4909);
and U6833 (N_6833,N_3746,N_579);
nand U6834 (N_6834,N_611,N_3868);
and U6835 (N_6835,N_1711,N_3914);
nand U6836 (N_6836,N_2106,N_220);
nor U6837 (N_6837,N_4938,N_946);
nor U6838 (N_6838,N_2912,N_641);
or U6839 (N_6839,N_2958,N_4798);
nand U6840 (N_6840,N_3996,N_869);
nand U6841 (N_6841,N_2813,N_892);
or U6842 (N_6842,N_4083,N_1544);
nor U6843 (N_6843,N_2503,N_3971);
nor U6844 (N_6844,N_89,N_845);
or U6845 (N_6845,N_290,N_3224);
nand U6846 (N_6846,N_1386,N_1523);
nand U6847 (N_6847,N_424,N_1353);
or U6848 (N_6848,N_227,N_3980);
and U6849 (N_6849,N_4019,N_2513);
or U6850 (N_6850,N_18,N_140);
or U6851 (N_6851,N_3255,N_293);
and U6852 (N_6852,N_547,N_2296);
nand U6853 (N_6853,N_3736,N_4541);
nor U6854 (N_6854,N_865,N_2572);
or U6855 (N_6855,N_3242,N_927);
nor U6856 (N_6856,N_2851,N_123);
nand U6857 (N_6857,N_1604,N_958);
nor U6858 (N_6858,N_4500,N_2974);
or U6859 (N_6859,N_2321,N_4285);
nand U6860 (N_6860,N_923,N_2579);
nand U6861 (N_6861,N_156,N_3871);
nand U6862 (N_6862,N_2788,N_4558);
nand U6863 (N_6863,N_316,N_1143);
nand U6864 (N_6864,N_320,N_2557);
nor U6865 (N_6865,N_4755,N_2222);
or U6866 (N_6866,N_568,N_1858);
nand U6867 (N_6867,N_1567,N_3142);
nor U6868 (N_6868,N_2251,N_1325);
nand U6869 (N_6869,N_4939,N_728);
nor U6870 (N_6870,N_176,N_1109);
or U6871 (N_6871,N_4398,N_1298);
and U6872 (N_6872,N_1693,N_609);
nand U6873 (N_6873,N_4651,N_1364);
nor U6874 (N_6874,N_2285,N_2034);
and U6875 (N_6875,N_4447,N_1557);
or U6876 (N_6876,N_3197,N_1444);
nor U6877 (N_6877,N_1224,N_2812);
or U6878 (N_6878,N_2000,N_3693);
and U6879 (N_6879,N_3814,N_403);
nor U6880 (N_6880,N_4808,N_4440);
and U6881 (N_6881,N_704,N_2455);
nand U6882 (N_6882,N_598,N_4800);
or U6883 (N_6883,N_3303,N_2626);
or U6884 (N_6884,N_1968,N_2021);
nor U6885 (N_6885,N_1592,N_3190);
xor U6886 (N_6886,N_1796,N_4203);
nand U6887 (N_6887,N_445,N_4245);
or U6888 (N_6888,N_2239,N_4989);
or U6889 (N_6889,N_2592,N_2929);
nor U6890 (N_6890,N_1714,N_936);
nor U6891 (N_6891,N_4214,N_4441);
and U6892 (N_6892,N_4556,N_3629);
and U6893 (N_6893,N_2884,N_4244);
and U6894 (N_6894,N_1438,N_1161);
nand U6895 (N_6895,N_2752,N_4049);
nor U6896 (N_6896,N_3024,N_1072);
and U6897 (N_6897,N_3286,N_3733);
or U6898 (N_6898,N_57,N_3827);
or U6899 (N_6899,N_3488,N_4821);
nand U6900 (N_6900,N_3110,N_2101);
nand U6901 (N_6901,N_4435,N_2246);
nand U6902 (N_6902,N_4057,N_621);
nand U6903 (N_6903,N_4320,N_743);
nor U6904 (N_6904,N_4216,N_4810);
and U6905 (N_6905,N_2530,N_4314);
and U6906 (N_6906,N_1468,N_2699);
nand U6907 (N_6907,N_1441,N_1339);
xor U6908 (N_6908,N_1208,N_135);
nand U6909 (N_6909,N_2918,N_3897);
nand U6910 (N_6910,N_3288,N_699);
nand U6911 (N_6911,N_2049,N_1241);
or U6912 (N_6912,N_2196,N_2908);
and U6913 (N_6913,N_4456,N_2799);
nor U6914 (N_6914,N_1573,N_4480);
and U6915 (N_6915,N_3050,N_4812);
nand U6916 (N_6916,N_3657,N_3406);
nand U6917 (N_6917,N_120,N_4219);
or U6918 (N_6918,N_3828,N_4844);
or U6919 (N_6919,N_1183,N_3434);
nand U6920 (N_6920,N_761,N_828);
or U6921 (N_6921,N_2023,N_860);
nor U6922 (N_6922,N_4349,N_3038);
or U6923 (N_6923,N_1988,N_2785);
nor U6924 (N_6924,N_4906,N_4152);
or U6925 (N_6925,N_2238,N_500);
nand U6926 (N_6926,N_2103,N_2172);
and U6927 (N_6927,N_2961,N_203);
and U6928 (N_6928,N_4351,N_4530);
or U6929 (N_6929,N_3307,N_1595);
or U6930 (N_6930,N_3004,N_2133);
nor U6931 (N_6931,N_3703,N_3767);
nor U6932 (N_6932,N_4408,N_4200);
nor U6933 (N_6933,N_367,N_586);
or U6934 (N_6934,N_1730,N_346);
nand U6935 (N_6935,N_1001,N_2862);
nor U6936 (N_6936,N_3374,N_2291);
or U6937 (N_6937,N_1011,N_3304);
nor U6938 (N_6938,N_1219,N_1974);
or U6939 (N_6939,N_4055,N_1);
or U6940 (N_6940,N_2100,N_1252);
nand U6941 (N_6941,N_1649,N_727);
or U6942 (N_6942,N_390,N_2694);
or U6943 (N_6943,N_925,N_4117);
nor U6944 (N_6944,N_2458,N_1138);
and U6945 (N_6945,N_2360,N_772);
nor U6946 (N_6946,N_2191,N_3727);
or U6947 (N_6947,N_4628,N_4171);
and U6948 (N_6948,N_2792,N_3047);
or U6949 (N_6949,N_2667,N_2793);
nand U6950 (N_6950,N_804,N_469);
nand U6951 (N_6951,N_4194,N_4969);
nor U6952 (N_6952,N_4459,N_1299);
or U6953 (N_6953,N_2518,N_3064);
nand U6954 (N_6954,N_4464,N_420);
and U6955 (N_6955,N_4515,N_4865);
nor U6956 (N_6956,N_3184,N_1021);
or U6957 (N_6957,N_1131,N_4820);
nor U6958 (N_6958,N_4930,N_2163);
nand U6959 (N_6959,N_4528,N_1244);
nand U6960 (N_6960,N_4835,N_4778);
and U6961 (N_6961,N_4472,N_4386);
and U6962 (N_6962,N_1539,N_4954);
nand U6963 (N_6963,N_3845,N_43);
nor U6964 (N_6964,N_4963,N_3756);
and U6965 (N_6965,N_3054,N_2546);
nor U6966 (N_6966,N_2942,N_2131);
nand U6967 (N_6967,N_3885,N_4261);
nor U6968 (N_6968,N_719,N_3235);
and U6969 (N_6969,N_4517,N_3326);
and U6970 (N_6970,N_1082,N_1306);
or U6971 (N_6971,N_4707,N_964);
nor U6972 (N_6972,N_1738,N_1907);
nand U6973 (N_6973,N_1589,N_1621);
nand U6974 (N_6974,N_4027,N_2664);
and U6975 (N_6975,N_4726,N_774);
and U6976 (N_6976,N_4510,N_1868);
or U6977 (N_6977,N_2421,N_3978);
nand U6978 (N_6978,N_1999,N_531);
nand U6979 (N_6979,N_2534,N_3600);
or U6980 (N_6980,N_2767,N_3860);
nor U6981 (N_6981,N_2204,N_4263);
nor U6982 (N_6982,N_3298,N_1303);
nand U6983 (N_6983,N_988,N_482);
or U6984 (N_6984,N_2519,N_1403);
or U6985 (N_6985,N_2591,N_3372);
and U6986 (N_6986,N_2419,N_3370);
xnor U6987 (N_6987,N_4679,N_4659);
and U6988 (N_6988,N_742,N_1715);
nand U6989 (N_6989,N_4048,N_2182);
nand U6990 (N_6990,N_4104,N_3593);
or U6991 (N_6991,N_2395,N_2938);
and U6992 (N_6992,N_4684,N_738);
nor U6993 (N_6993,N_1226,N_3663);
nand U6994 (N_6994,N_2032,N_3824);
or U6995 (N_6995,N_431,N_2515);
nand U6996 (N_6996,N_1888,N_3869);
nand U6997 (N_6997,N_2605,N_3676);
or U6998 (N_6998,N_4380,N_4884);
and U6999 (N_6999,N_1921,N_369);
nand U7000 (N_7000,N_1290,N_2678);
or U7001 (N_7001,N_1572,N_1318);
and U7002 (N_7002,N_3835,N_23);
nor U7003 (N_7003,N_4434,N_1196);
or U7004 (N_7004,N_4643,N_1395);
and U7005 (N_7005,N_2900,N_3918);
or U7006 (N_7006,N_3466,N_4839);
or U7007 (N_7007,N_1443,N_1338);
and U7008 (N_7008,N_3847,N_535);
or U7009 (N_7009,N_2017,N_2648);
nor U7010 (N_7010,N_2467,N_4364);
and U7011 (N_7011,N_201,N_2452);
or U7012 (N_7012,N_4343,N_3168);
nand U7013 (N_7013,N_1446,N_2892);
or U7014 (N_7014,N_4507,N_2903);
or U7015 (N_7015,N_3185,N_69);
or U7016 (N_7016,N_235,N_650);
nor U7017 (N_7017,N_3293,N_2135);
and U7018 (N_7018,N_1269,N_3981);
nand U7019 (N_7019,N_4311,N_4649);
nor U7020 (N_7020,N_3514,N_1480);
nand U7021 (N_7021,N_3575,N_3504);
or U7022 (N_7022,N_3128,N_2357);
or U7023 (N_7023,N_116,N_4414);
and U7024 (N_7024,N_2508,N_4566);
and U7025 (N_7025,N_4520,N_1030);
or U7026 (N_7026,N_4769,N_2819);
or U7027 (N_7027,N_340,N_304);
or U7028 (N_7028,N_99,N_1861);
and U7029 (N_7029,N_4420,N_538);
and U7030 (N_7030,N_4297,N_655);
nor U7031 (N_7031,N_1483,N_4843);
nand U7032 (N_7032,N_1225,N_2954);
nor U7033 (N_7033,N_1910,N_1541);
and U7034 (N_7034,N_4877,N_3801);
nor U7035 (N_7035,N_448,N_3396);
nand U7036 (N_7036,N_2598,N_3789);
and U7037 (N_7037,N_4690,N_2474);
nand U7038 (N_7038,N_841,N_4536);
or U7039 (N_7039,N_665,N_3333);
nand U7040 (N_7040,N_1679,N_3819);
nand U7041 (N_7041,N_2141,N_3543);
or U7042 (N_7042,N_771,N_1623);
nand U7043 (N_7043,N_2832,N_1418);
and U7044 (N_7044,N_1716,N_3193);
or U7045 (N_7045,N_634,N_3179);
and U7046 (N_7046,N_452,N_4091);
nor U7047 (N_7047,N_1871,N_3423);
nand U7048 (N_7048,N_236,N_1983);
or U7049 (N_7049,N_4741,N_521);
and U7050 (N_7050,N_4286,N_876);
nand U7051 (N_7051,N_4179,N_2332);
nand U7052 (N_7052,N_1972,N_3574);
or U7053 (N_7053,N_3555,N_394);
and U7054 (N_7054,N_1276,N_812);
and U7055 (N_7055,N_47,N_3498);
nand U7056 (N_7056,N_347,N_3346);
nor U7057 (N_7057,N_4250,N_1624);
or U7058 (N_7058,N_943,N_2741);
nor U7059 (N_7059,N_1923,N_3133);
and U7060 (N_7060,N_4545,N_763);
nand U7061 (N_7061,N_2011,N_3913);
or U7062 (N_7062,N_691,N_2651);
or U7063 (N_7063,N_1366,N_637);
nand U7064 (N_7064,N_2373,N_1238);
nand U7065 (N_7065,N_3022,N_31);
nor U7066 (N_7066,N_1074,N_205);
and U7067 (N_7067,N_1785,N_768);
nand U7068 (N_7068,N_4940,N_2507);
or U7069 (N_7069,N_1365,N_3067);
or U7070 (N_7070,N_1371,N_1695);
and U7071 (N_7071,N_3650,N_2492);
or U7072 (N_7072,N_1908,N_505);
nor U7073 (N_7073,N_125,N_3944);
and U7074 (N_7074,N_4097,N_2283);
nand U7075 (N_7075,N_3160,N_3716);
nor U7076 (N_7076,N_1642,N_4854);
nand U7077 (N_7077,N_3223,N_4732);
or U7078 (N_7078,N_153,N_228);
and U7079 (N_7079,N_1417,N_2446);
or U7080 (N_7080,N_3922,N_1732);
nand U7081 (N_7081,N_2292,N_3920);
or U7082 (N_7082,N_999,N_3208);
nand U7083 (N_7083,N_4204,N_4513);
nor U7084 (N_7084,N_58,N_1392);
nor U7085 (N_7085,N_2122,N_1607);
nor U7086 (N_7086,N_1317,N_3409);
and U7087 (N_7087,N_4121,N_2007);
nand U7088 (N_7088,N_947,N_3348);
nand U7089 (N_7089,N_150,N_4470);
nor U7090 (N_7090,N_4006,N_276);
nand U7091 (N_7091,N_4526,N_2209);
and U7092 (N_7092,N_3350,N_1465);
and U7093 (N_7093,N_541,N_2008);
or U7094 (N_7094,N_4181,N_3536);
nor U7095 (N_7095,N_933,N_3559);
or U7096 (N_7096,N_4142,N_2381);
nor U7097 (N_7097,N_1844,N_331);
nor U7098 (N_7098,N_3428,N_3130);
nor U7099 (N_7099,N_3643,N_2353);
nand U7100 (N_7100,N_4066,N_2842);
or U7101 (N_7101,N_1289,N_4836);
and U7102 (N_7102,N_4891,N_961);
and U7103 (N_7103,N_137,N_476);
and U7104 (N_7104,N_4667,N_1759);
nand U7105 (N_7105,N_2815,N_1164);
nor U7106 (N_7106,N_3952,N_4911);
or U7107 (N_7107,N_1766,N_312);
nand U7108 (N_7108,N_1638,N_877);
nand U7109 (N_7109,N_3183,N_1195);
and U7110 (N_7110,N_888,N_1873);
and U7111 (N_7111,N_160,N_1043);
nand U7112 (N_7112,N_1948,N_2216);
nand U7113 (N_7113,N_4544,N_1952);
nand U7114 (N_7114,N_3912,N_1571);
and U7115 (N_7115,N_1756,N_2001);
and U7116 (N_7116,N_3151,N_4271);
nor U7117 (N_7117,N_2926,N_750);
nand U7118 (N_7118,N_4090,N_2998);
and U7119 (N_7119,N_224,N_2880);
nor U7120 (N_7120,N_2625,N_2315);
nand U7121 (N_7121,N_1322,N_4900);
nor U7122 (N_7122,N_862,N_2666);
and U7123 (N_7123,N_2556,N_4752);
and U7124 (N_7124,N_1301,N_4557);
nor U7125 (N_7125,N_4333,N_3245);
and U7126 (N_7126,N_1258,N_1094);
and U7127 (N_7127,N_2568,N_2779);
nor U7128 (N_7128,N_3967,N_272);
nand U7129 (N_7129,N_4538,N_4191);
and U7130 (N_7130,N_1493,N_3401);
and U7131 (N_7131,N_1822,N_2311);
or U7132 (N_7132,N_4701,N_3131);
and U7133 (N_7133,N_3416,N_1079);
nor U7134 (N_7134,N_2717,N_4446);
nor U7135 (N_7135,N_3200,N_4444);
nor U7136 (N_7136,N_1336,N_1576);
or U7137 (N_7137,N_53,N_3939);
nor U7138 (N_7138,N_488,N_1279);
or U7139 (N_7139,N_1762,N_297);
nand U7140 (N_7140,N_607,N_3163);
nor U7141 (N_7141,N_380,N_1728);
nand U7142 (N_7142,N_1452,N_239);
and U7143 (N_7143,N_3309,N_42);
and U7144 (N_7144,N_821,N_1378);
nand U7145 (N_7145,N_2470,N_577);
or U7146 (N_7146,N_4301,N_3375);
or U7147 (N_7147,N_3975,N_4123);
and U7148 (N_7148,N_2499,N_3069);
or U7149 (N_7149,N_624,N_2406);
nor U7150 (N_7150,N_3258,N_4350);
and U7151 (N_7151,N_2636,N_3532);
and U7152 (N_7152,N_4046,N_3253);
nand U7153 (N_7153,N_715,N_2684);
or U7154 (N_7154,N_4921,N_2784);
and U7155 (N_7155,N_696,N_147);
and U7156 (N_7156,N_4427,N_1090);
or U7157 (N_7157,N_1066,N_3033);
nand U7158 (N_7158,N_3284,N_1152);
and U7159 (N_7159,N_1234,N_279);
nand U7160 (N_7160,N_839,N_1459);
and U7161 (N_7161,N_1689,N_4025);
nand U7162 (N_7162,N_3311,N_1487);
and U7163 (N_7163,N_1351,N_2185);
or U7164 (N_7164,N_3039,N_498);
or U7165 (N_7165,N_4436,N_1223);
and U7166 (N_7166,N_741,N_3910);
and U7167 (N_7167,N_2941,N_252);
nand U7168 (N_7168,N_542,N_3403);
xor U7169 (N_7169,N_1231,N_3700);
and U7170 (N_7170,N_692,N_3181);
and U7171 (N_7171,N_2821,N_921);
nand U7172 (N_7172,N_1151,N_4770);
and U7173 (N_7173,N_1675,N_1551);
or U7174 (N_7174,N_3726,N_3652);
and U7175 (N_7175,N_785,N_2026);
nand U7176 (N_7176,N_3988,N_202);
nand U7177 (N_7177,N_3376,N_2584);
nand U7178 (N_7178,N_4230,N_1754);
or U7179 (N_7179,N_3915,N_4391);
and U7180 (N_7180,N_3485,N_3724);
nand U7181 (N_7181,N_4549,N_2746);
nor U7182 (N_7182,N_939,N_1685);
or U7183 (N_7183,N_3491,N_1971);
nor U7184 (N_7184,N_1343,N_2109);
and U7185 (N_7185,N_3560,N_2898);
nor U7186 (N_7186,N_4756,N_2383);
nand U7187 (N_7187,N_1199,N_3883);
nand U7188 (N_7188,N_2946,N_2715);
and U7189 (N_7189,N_4030,N_86);
nand U7190 (N_7190,N_2525,N_1605);
nor U7191 (N_7191,N_4560,N_4465);
and U7192 (N_7192,N_2629,N_2872);
nand U7193 (N_7193,N_3053,N_2670);
nor U7194 (N_7194,N_4571,N_2805);
and U7195 (N_7195,N_2493,N_2766);
and U7196 (N_7196,N_1470,N_4180);
and U7197 (N_7197,N_454,N_2937);
or U7198 (N_7198,N_1826,N_2038);
nor U7199 (N_7199,N_3119,N_233);
and U7200 (N_7200,N_2494,N_4523);
or U7201 (N_7201,N_94,N_685);
and U7202 (N_7202,N_101,N_1172);
nand U7203 (N_7203,N_232,N_3673);
and U7204 (N_7204,N_4497,N_1966);
nor U7205 (N_7205,N_4468,N_2009);
nand U7206 (N_7206,N_2121,N_2560);
and U7207 (N_7207,N_1838,N_3513);
nand U7208 (N_7208,N_4893,N_1884);
nand U7209 (N_7209,N_4024,N_1896);
xor U7210 (N_7210,N_1775,N_2362);
nor U7211 (N_7211,N_338,N_2489);
and U7212 (N_7212,N_3421,N_3945);
nand U7213 (N_7213,N_3344,N_1275);
nand U7214 (N_7214,N_2617,N_4237);
and U7215 (N_7215,N_3044,N_3219);
nand U7216 (N_7216,N_4749,N_565);
xor U7217 (N_7217,N_1660,N_626);
nand U7218 (N_7218,N_3331,N_2097);
and U7219 (N_7219,N_1901,N_2304);
nand U7220 (N_7220,N_3956,N_4878);
or U7221 (N_7221,N_980,N_3603);
and U7222 (N_7222,N_4397,N_1069);
or U7223 (N_7223,N_462,N_654);
and U7224 (N_7224,N_4257,N_1203);
and U7225 (N_7225,N_1630,N_3648);
and U7226 (N_7226,N_635,N_4685);
nor U7227 (N_7227,N_3156,N_625);
nand U7228 (N_7228,N_4620,N_4428);
or U7229 (N_7229,N_3411,N_3832);
and U7230 (N_7230,N_1193,N_255);
or U7231 (N_7231,N_1933,N_2327);
or U7232 (N_7232,N_4801,N_3377);
and U7233 (N_7233,N_4894,N_1281);
and U7234 (N_7234,N_4700,N_1092);
nand U7235 (N_7235,N_1163,N_4269);
and U7236 (N_7236,N_3891,N_797);
nor U7237 (N_7237,N_570,N_3495);
or U7238 (N_7238,N_2215,N_3217);
or U7239 (N_7239,N_2088,N_4658);
nor U7240 (N_7240,N_4537,N_3499);
and U7241 (N_7241,N_3259,N_710);
nand U7242 (N_7242,N_1863,N_3373);
nand U7243 (N_7243,N_3093,N_2700);
or U7244 (N_7244,N_406,N_77);
and U7245 (N_7245,N_1115,N_2949);
or U7246 (N_7246,N_792,N_1022);
or U7247 (N_7247,N_627,N_1401);
and U7248 (N_7248,N_4635,N_4997);
nor U7249 (N_7249,N_2803,N_2615);
nor U7250 (N_7250,N_4215,N_1918);
and U7251 (N_7251,N_3854,N_2932);
and U7252 (N_7252,N_2863,N_1284);
and U7253 (N_7253,N_2279,N_472);
or U7254 (N_7254,N_3077,N_2604);
nand U7255 (N_7255,N_1267,N_4390);
or U7256 (N_7256,N_3104,N_2371);
and U7257 (N_7257,N_3515,N_2295);
and U7258 (N_7258,N_103,N_1664);
and U7259 (N_7259,N_3842,N_3216);
nand U7260 (N_7260,N_1562,N_1170);
and U7261 (N_7261,N_4823,N_1404);
or U7262 (N_7262,N_2588,N_3812);
nor U7263 (N_7263,N_499,N_2687);
nor U7264 (N_7264,N_837,N_2680);
and U7265 (N_7265,N_1361,N_4471);
nor U7266 (N_7266,N_3278,N_1264);
or U7267 (N_7267,N_3486,N_4176);
or U7268 (N_7268,N_3221,N_3889);
nand U7269 (N_7269,N_1134,N_231);
or U7270 (N_7270,N_3839,N_2778);
nand U7271 (N_7271,N_3263,N_3302);
nand U7272 (N_7272,N_1307,N_2263);
nand U7273 (N_7273,N_4992,N_3664);
nor U7274 (N_7274,N_4124,N_1070);
nand U7275 (N_7275,N_1356,N_510);
and U7276 (N_7276,N_857,N_1342);
nor U7277 (N_7277,N_852,N_1580);
nor U7278 (N_7278,N_4654,N_1771);
or U7279 (N_7279,N_4035,N_303);
nor U7280 (N_7280,N_1243,N_4720);
nor U7281 (N_7281,N_4370,N_1639);
and U7282 (N_7282,N_4341,N_4753);
or U7283 (N_7283,N_378,N_4990);
nor U7284 (N_7284,N_1776,N_3087);
nand U7285 (N_7285,N_2430,N_1068);
nand U7286 (N_7286,N_244,N_910);
or U7287 (N_7287,N_2480,N_3220);
or U7288 (N_7288,N_3169,N_1357);
and U7289 (N_7289,N_3210,N_1104);
or U7290 (N_7290,N_2230,N_3782);
or U7291 (N_7291,N_119,N_418);
nor U7292 (N_7292,N_4688,N_3890);
and U7293 (N_7293,N_1335,N_3723);
and U7294 (N_7294,N_794,N_385);
nor U7295 (N_7295,N_1706,N_492);
nor U7296 (N_7296,N_3349,N_2906);
or U7297 (N_7297,N_1960,N_4942);
nor U7298 (N_7298,N_4670,N_2047);
and U7299 (N_7299,N_238,N_512);
nor U7300 (N_7300,N_585,N_4789);
nand U7301 (N_7301,N_3066,N_4762);
nor U7302 (N_7302,N_149,N_920);
nor U7303 (N_7303,N_4017,N_2299);
nand U7304 (N_7304,N_1376,N_3035);
and U7305 (N_7305,N_3748,N_2967);
and U7306 (N_7306,N_4079,N_3088);
nand U7307 (N_7307,N_3198,N_3489);
and U7308 (N_7308,N_441,N_1860);
nand U7309 (N_7309,N_529,N_1705);
xnor U7310 (N_7310,N_2867,N_3356);
nand U7311 (N_7311,N_2445,N_1829);
or U7312 (N_7312,N_3710,N_1965);
nand U7313 (N_7313,N_3682,N_1987);
nor U7314 (N_7314,N_1372,N_2798);
and U7315 (N_7315,N_1160,N_1955);
or U7316 (N_7316,N_4951,N_4001);
or U7317 (N_7317,N_2085,N_2611);
nand U7318 (N_7318,N_4260,N_3622);
nor U7319 (N_7319,N_3781,N_3097);
nand U7320 (N_7320,N_2143,N_543);
nand U7321 (N_7321,N_4081,N_3394);
nand U7322 (N_7322,N_4982,N_2242);
and U7323 (N_7323,N_371,N_3287);
nor U7324 (N_7324,N_2337,N_2765);
nor U7325 (N_7325,N_4022,N_3982);
nand U7326 (N_7326,N_1375,N_2170);
or U7327 (N_7327,N_1402,N_3651);
or U7328 (N_7328,N_3474,N_1390);
and U7329 (N_7329,N_3337,N_3180);
nand U7330 (N_7330,N_1512,N_3627);
or U7331 (N_7331,N_1415,N_4029);
nor U7332 (N_7332,N_2140,N_3645);
or U7333 (N_7333,N_1681,N_1938);
or U7334 (N_7334,N_610,N_2003);
or U7335 (N_7335,N_1045,N_1815);
nor U7336 (N_7336,N_1799,N_3261);
nor U7337 (N_7337,N_3906,N_3753);
nand U7338 (N_7338,N_4475,N_2733);
nand U7339 (N_7339,N_4094,N_749);
nand U7340 (N_7340,N_2069,N_3919);
and U7341 (N_7341,N_900,N_4983);
or U7342 (N_7342,N_2234,N_3134);
nand U7343 (N_7343,N_1597,N_3062);
or U7344 (N_7344,N_2902,N_827);
or U7345 (N_7345,N_864,N_604);
nor U7346 (N_7346,N_1036,N_242);
nand U7347 (N_7347,N_4845,N_4190);
nor U7348 (N_7348,N_496,N_2281);
or U7349 (N_7349,N_4043,N_1429);
xor U7350 (N_7350,N_3078,N_2220);
nor U7351 (N_7351,N_902,N_4981);
nor U7352 (N_7352,N_2347,N_1812);
and U7353 (N_7353,N_4542,N_1760);
and U7354 (N_7354,N_4804,N_4107);
or U7355 (N_7355,N_4624,N_1990);
nand U7356 (N_7356,N_4972,N_1270);
and U7357 (N_7357,N_3150,N_3701);
nor U7358 (N_7358,N_250,N_3427);
or U7359 (N_7359,N_2484,N_3862);
nor U7360 (N_7360,N_3222,N_3111);
and U7361 (N_7361,N_1778,N_3250);
and U7362 (N_7362,N_2790,N_4704);
nand U7363 (N_7363,N_4807,N_2674);
nand U7364 (N_7364,N_195,N_3853);
or U7365 (N_7365,N_4483,N_4642);
or U7366 (N_7366,N_2802,N_2889);
nand U7367 (N_7367,N_1502,N_4705);
nand U7368 (N_7368,N_3572,N_3398);
nand U7369 (N_7369,N_868,N_3632);
nand U7370 (N_7370,N_908,N_2931);
and U7371 (N_7371,N_4551,N_3315);
nor U7372 (N_7372,N_1586,N_4232);
nor U7373 (N_7373,N_2084,N_4274);
nand U7374 (N_7374,N_3826,N_1496);
nor U7375 (N_7375,N_1798,N_2208);
nor U7376 (N_7376,N_2882,N_4110);
or U7377 (N_7377,N_3170,N_196);
nor U7378 (N_7378,N_3838,N_4847);
nor U7379 (N_7379,N_674,N_3459);
and U7380 (N_7380,N_4923,N_1782);
and U7381 (N_7381,N_3055,N_197);
nor U7382 (N_7382,N_3503,N_3993);
nor U7383 (N_7383,N_594,N_4868);
xnor U7384 (N_7384,N_1360,N_4307);
or U7385 (N_7385,N_3904,N_4650);
nand U7386 (N_7386,N_4797,N_4585);
nand U7387 (N_7387,N_3678,N_2497);
nand U7388 (N_7388,N_2396,N_2429);
or U7389 (N_7389,N_4007,N_3734);
nand U7390 (N_7390,N_2426,N_3023);
nor U7391 (N_7391,N_2090,N_4499);
and U7392 (N_7392,N_114,N_1171);
nand U7393 (N_7393,N_4694,N_4512);
nor U7394 (N_7394,N_3395,N_2261);
nor U7395 (N_7395,N_4021,N_1961);
nand U7396 (N_7396,N_4855,N_2094);
or U7397 (N_7397,N_387,N_3127);
nor U7398 (N_7398,N_4150,N_4388);
nand U7399 (N_7399,N_2129,N_2913);
and U7400 (N_7400,N_319,N_1632);
and U7401 (N_7401,N_3249,N_465);
nand U7402 (N_7402,N_658,N_3822);
or U7403 (N_7403,N_4803,N_4748);
or U7404 (N_7404,N_1820,N_2414);
or U7405 (N_7405,N_1287,N_3517);
nand U7406 (N_7406,N_2944,N_2108);
nor U7407 (N_7407,N_1672,N_2293);
and U7408 (N_7408,N_2427,N_3613);
nor U7409 (N_7409,N_1790,N_1481);
nor U7410 (N_7410,N_4889,N_4129);
nand U7411 (N_7411,N_2691,N_4718);
nand U7412 (N_7412,N_1973,N_1867);
nand U7413 (N_7413,N_2745,N_2650);
or U7414 (N_7414,N_1256,N_3458);
nand U7415 (N_7415,N_3117,N_3669);
or U7416 (N_7416,N_3808,N_56);
or U7417 (N_7417,N_3003,N_4687);
or U7418 (N_7418,N_4466,N_2074);
and U7419 (N_7419,N_2894,N_3490);
or U7420 (N_7420,N_3477,N_3384);
and U7421 (N_7421,N_3319,N_2891);
nand U7422 (N_7422,N_1222,N_783);
nor U7423 (N_7423,N_3520,N_4723);
and U7424 (N_7424,N_2724,N_1019);
and U7425 (N_7425,N_969,N_967);
nor U7426 (N_7426,N_3892,N_3802);
and U7427 (N_7427,N_1899,N_1369);
or U7428 (N_7428,N_3636,N_3391);
and U7429 (N_7429,N_2247,N_4572);
nand U7430 (N_7430,N_4788,N_4929);
nand U7431 (N_7431,N_4,N_66);
nand U7432 (N_7432,N_294,N_2179);
nor U7433 (N_7433,N_3876,N_4383);
nor U7434 (N_7434,N_4159,N_1363);
nand U7435 (N_7435,N_198,N_3325);
and U7436 (N_7436,N_4265,N_4637);
nor U7437 (N_7437,N_133,N_3174);
or U7438 (N_7438,N_2449,N_1819);
nor U7439 (N_7439,N_1886,N_1912);
or U7440 (N_7440,N_128,N_3965);
nor U7441 (N_7441,N_4727,N_4636);
nor U7442 (N_7442,N_37,N_358);
or U7443 (N_7443,N_206,N_3596);
nor U7444 (N_7444,N_3954,N_1636);
or U7445 (N_7445,N_3410,N_1827);
or U7446 (N_7446,N_2134,N_3092);
nor U7447 (N_7447,N_204,N_2639);
nand U7448 (N_7448,N_4945,N_4780);
and U7449 (N_7449,N_3841,N_408);
nand U7450 (N_7450,N_3057,N_3494);
and U7451 (N_7451,N_415,N_2529);
nor U7452 (N_7452,N_4745,N_3011);
and U7453 (N_7453,N_438,N_2527);
or U7454 (N_7454,N_3164,N_4394);
nand U7455 (N_7455,N_891,N_4018);
or U7456 (N_7456,N_138,N_2225);
nand U7457 (N_7457,N_2,N_3021);
nor U7458 (N_7458,N_166,N_2876);
nand U7459 (N_7459,N_1297,N_4211);
nand U7460 (N_7460,N_4327,N_4641);
and U7461 (N_7461,N_2675,N_1617);
nand U7462 (N_7462,N_2726,N_4863);
and U7463 (N_7463,N_4988,N_4890);
or U7464 (N_7464,N_758,N_1412);
xor U7465 (N_7465,N_456,N_1903);
and U7466 (N_7466,N_1692,N_2703);
nor U7467 (N_7467,N_4577,N_3330);
nor U7468 (N_7468,N_2243,N_563);
nor U7469 (N_7469,N_4646,N_264);
nor U7470 (N_7470,N_3943,N_2297);
nor U7471 (N_7471,N_1742,N_2707);
nor U7472 (N_7472,N_3501,N_3361);
nand U7473 (N_7473,N_3665,N_2171);
nand U7474 (N_7474,N_3911,N_682);
nor U7475 (N_7475,N_1862,N_2061);
nand U7476 (N_7476,N_3158,N_4188);
or U7477 (N_7477,N_3878,N_249);
and U7478 (N_7478,N_4306,N_3308);
or U7479 (N_7479,N_1211,N_4621);
or U7480 (N_7480,N_307,N_4703);
nand U7481 (N_7481,N_781,N_3270);
nand U7482 (N_7482,N_2531,N_4608);
and U7483 (N_7483,N_677,N_1665);
and U7484 (N_7484,N_3071,N_4849);
nor U7485 (N_7485,N_2740,N_1981);
or U7486 (N_7486,N_1872,N_3452);
and U7487 (N_7487,N_1176,N_351);
and U7488 (N_7488,N_3540,N_3888);
nor U7489 (N_7489,N_296,N_3599);
or U7490 (N_7490,N_2564,N_2486);
nor U7491 (N_7491,N_1188,N_4113);
and U7492 (N_7492,N_1233,N_628);
and U7493 (N_7493,N_1755,N_2128);
nand U7494 (N_7494,N_3793,N_3989);
nand U7495 (N_7495,N_4323,N_1939);
nor U7496 (N_7496,N_3783,N_1596);
and U7497 (N_7497,N_1600,N_3187);
nand U7498 (N_7498,N_302,N_669);
nor U7499 (N_7499,N_2800,N_4034);
nand U7500 (N_7500,N_3571,N_4195);
nor U7501 (N_7501,N_2566,N_1399);
or U7502 (N_7502,N_3599,N_4919);
nand U7503 (N_7503,N_517,N_4527);
and U7504 (N_7504,N_1767,N_2796);
and U7505 (N_7505,N_221,N_4593);
nand U7506 (N_7506,N_4923,N_210);
or U7507 (N_7507,N_3566,N_4380);
or U7508 (N_7508,N_2925,N_417);
and U7509 (N_7509,N_3596,N_3507);
nand U7510 (N_7510,N_884,N_1060);
nor U7511 (N_7511,N_894,N_4710);
nand U7512 (N_7512,N_299,N_609);
or U7513 (N_7513,N_4931,N_3742);
or U7514 (N_7514,N_3607,N_1782);
or U7515 (N_7515,N_4625,N_2651);
and U7516 (N_7516,N_55,N_3493);
or U7517 (N_7517,N_2735,N_3881);
nand U7518 (N_7518,N_353,N_3919);
nand U7519 (N_7519,N_405,N_4318);
nor U7520 (N_7520,N_1839,N_3378);
nor U7521 (N_7521,N_4710,N_2540);
and U7522 (N_7522,N_1773,N_4717);
nand U7523 (N_7523,N_581,N_2873);
or U7524 (N_7524,N_4330,N_1926);
or U7525 (N_7525,N_718,N_4573);
and U7526 (N_7526,N_2784,N_1996);
nor U7527 (N_7527,N_4281,N_1617);
nand U7528 (N_7528,N_2285,N_3208);
nand U7529 (N_7529,N_571,N_1121);
nor U7530 (N_7530,N_4043,N_891);
nor U7531 (N_7531,N_2458,N_2216);
or U7532 (N_7532,N_468,N_3930);
nor U7533 (N_7533,N_1393,N_3127);
and U7534 (N_7534,N_3234,N_549);
or U7535 (N_7535,N_281,N_4392);
and U7536 (N_7536,N_70,N_1961);
nor U7537 (N_7537,N_3757,N_231);
nor U7538 (N_7538,N_3458,N_1975);
nand U7539 (N_7539,N_2899,N_2389);
nor U7540 (N_7540,N_694,N_164);
nand U7541 (N_7541,N_3416,N_625);
nand U7542 (N_7542,N_666,N_216);
and U7543 (N_7543,N_832,N_1120);
nand U7544 (N_7544,N_4301,N_1323);
nand U7545 (N_7545,N_3515,N_3612);
and U7546 (N_7546,N_3972,N_4198);
xor U7547 (N_7547,N_164,N_3088);
or U7548 (N_7548,N_2378,N_3094);
and U7549 (N_7549,N_3774,N_2438);
nor U7550 (N_7550,N_2530,N_1795);
nor U7551 (N_7551,N_2157,N_2120);
or U7552 (N_7552,N_2022,N_4603);
nor U7553 (N_7553,N_2452,N_2411);
nand U7554 (N_7554,N_3738,N_22);
nand U7555 (N_7555,N_3214,N_1031);
nand U7556 (N_7556,N_602,N_3252);
or U7557 (N_7557,N_3508,N_4515);
or U7558 (N_7558,N_1140,N_4747);
nand U7559 (N_7559,N_2563,N_3854);
nand U7560 (N_7560,N_1320,N_4900);
nor U7561 (N_7561,N_834,N_2808);
nand U7562 (N_7562,N_3177,N_4587);
and U7563 (N_7563,N_1426,N_1427);
nor U7564 (N_7564,N_3766,N_3835);
or U7565 (N_7565,N_2949,N_1652);
nand U7566 (N_7566,N_4938,N_3585);
nor U7567 (N_7567,N_1182,N_4236);
nor U7568 (N_7568,N_4305,N_4224);
nor U7569 (N_7569,N_1030,N_161);
and U7570 (N_7570,N_1459,N_1955);
nor U7571 (N_7571,N_4492,N_4723);
or U7572 (N_7572,N_898,N_2670);
and U7573 (N_7573,N_1032,N_1603);
nor U7574 (N_7574,N_2489,N_4795);
nand U7575 (N_7575,N_434,N_1515);
nor U7576 (N_7576,N_3547,N_2265);
or U7577 (N_7577,N_2183,N_2780);
and U7578 (N_7578,N_2498,N_237);
or U7579 (N_7579,N_4313,N_2748);
nand U7580 (N_7580,N_1292,N_2076);
or U7581 (N_7581,N_275,N_2055);
and U7582 (N_7582,N_4586,N_4489);
nor U7583 (N_7583,N_2706,N_3947);
and U7584 (N_7584,N_607,N_2288);
or U7585 (N_7585,N_1102,N_3706);
nand U7586 (N_7586,N_4701,N_1896);
or U7587 (N_7587,N_1141,N_1467);
nand U7588 (N_7588,N_1437,N_1480);
or U7589 (N_7589,N_1125,N_1959);
or U7590 (N_7590,N_208,N_451);
nand U7591 (N_7591,N_4953,N_120);
nand U7592 (N_7592,N_1631,N_2889);
nor U7593 (N_7593,N_1772,N_1089);
and U7594 (N_7594,N_1810,N_4157);
and U7595 (N_7595,N_4542,N_2909);
nand U7596 (N_7596,N_1050,N_4260);
nand U7597 (N_7597,N_2758,N_2453);
xor U7598 (N_7598,N_1473,N_4251);
or U7599 (N_7599,N_3494,N_952);
nand U7600 (N_7600,N_3403,N_4962);
or U7601 (N_7601,N_1438,N_3182);
and U7602 (N_7602,N_1341,N_355);
or U7603 (N_7603,N_4815,N_4192);
nand U7604 (N_7604,N_2507,N_4519);
and U7605 (N_7605,N_1211,N_4733);
or U7606 (N_7606,N_4032,N_2340);
xor U7607 (N_7607,N_3725,N_3954);
nand U7608 (N_7608,N_3844,N_1732);
nand U7609 (N_7609,N_1086,N_2337);
and U7610 (N_7610,N_4814,N_3754);
nor U7611 (N_7611,N_1714,N_4777);
or U7612 (N_7612,N_4817,N_3776);
and U7613 (N_7613,N_3329,N_2398);
nand U7614 (N_7614,N_1989,N_4990);
nand U7615 (N_7615,N_1232,N_2895);
nand U7616 (N_7616,N_1213,N_1272);
and U7617 (N_7617,N_3774,N_4655);
nand U7618 (N_7618,N_1528,N_4035);
nand U7619 (N_7619,N_2577,N_3049);
nand U7620 (N_7620,N_463,N_2966);
nor U7621 (N_7621,N_2235,N_3346);
or U7622 (N_7622,N_4898,N_999);
and U7623 (N_7623,N_672,N_2262);
and U7624 (N_7624,N_3856,N_456);
and U7625 (N_7625,N_3801,N_4148);
nand U7626 (N_7626,N_4038,N_2559);
nor U7627 (N_7627,N_2269,N_3021);
nor U7628 (N_7628,N_4465,N_283);
or U7629 (N_7629,N_3938,N_2882);
nor U7630 (N_7630,N_2812,N_4004);
or U7631 (N_7631,N_2769,N_380);
nand U7632 (N_7632,N_690,N_4700);
nand U7633 (N_7633,N_4656,N_4914);
or U7634 (N_7634,N_2499,N_837);
nand U7635 (N_7635,N_1366,N_2543);
or U7636 (N_7636,N_375,N_4562);
nor U7637 (N_7637,N_3121,N_2645);
or U7638 (N_7638,N_4480,N_1476);
nor U7639 (N_7639,N_4197,N_1692);
nand U7640 (N_7640,N_4691,N_116);
nand U7641 (N_7641,N_3350,N_4587);
nand U7642 (N_7642,N_163,N_3043);
nor U7643 (N_7643,N_4538,N_273);
nor U7644 (N_7644,N_1498,N_2893);
nor U7645 (N_7645,N_2092,N_1565);
or U7646 (N_7646,N_2978,N_4976);
or U7647 (N_7647,N_2898,N_1159);
and U7648 (N_7648,N_1315,N_4289);
nand U7649 (N_7649,N_1244,N_4355);
nor U7650 (N_7650,N_1922,N_3916);
and U7651 (N_7651,N_4407,N_1515);
nor U7652 (N_7652,N_1628,N_1010);
nor U7653 (N_7653,N_551,N_3779);
and U7654 (N_7654,N_1011,N_3945);
nand U7655 (N_7655,N_1890,N_4597);
and U7656 (N_7656,N_4924,N_2542);
and U7657 (N_7657,N_2249,N_2939);
and U7658 (N_7658,N_2014,N_3869);
nand U7659 (N_7659,N_879,N_3304);
or U7660 (N_7660,N_4889,N_3944);
nor U7661 (N_7661,N_3264,N_3532);
nand U7662 (N_7662,N_3121,N_2904);
nand U7663 (N_7663,N_671,N_4975);
or U7664 (N_7664,N_3173,N_1278);
nand U7665 (N_7665,N_3466,N_3279);
or U7666 (N_7666,N_2578,N_2730);
and U7667 (N_7667,N_3914,N_3683);
and U7668 (N_7668,N_4039,N_1743);
and U7669 (N_7669,N_3119,N_3859);
and U7670 (N_7670,N_2340,N_1630);
or U7671 (N_7671,N_4249,N_1776);
and U7672 (N_7672,N_192,N_1732);
nand U7673 (N_7673,N_2527,N_366);
or U7674 (N_7674,N_1406,N_4631);
and U7675 (N_7675,N_310,N_4923);
or U7676 (N_7676,N_3737,N_1800);
and U7677 (N_7677,N_1533,N_1117);
and U7678 (N_7678,N_3456,N_1165);
nand U7679 (N_7679,N_4543,N_622);
or U7680 (N_7680,N_3507,N_2342);
nand U7681 (N_7681,N_2773,N_2250);
nor U7682 (N_7682,N_2613,N_1038);
and U7683 (N_7683,N_4617,N_3819);
or U7684 (N_7684,N_487,N_2705);
or U7685 (N_7685,N_3753,N_1865);
or U7686 (N_7686,N_2666,N_1896);
nor U7687 (N_7687,N_3672,N_4423);
or U7688 (N_7688,N_45,N_994);
or U7689 (N_7689,N_1971,N_633);
and U7690 (N_7690,N_3462,N_2875);
and U7691 (N_7691,N_410,N_1031);
and U7692 (N_7692,N_179,N_2537);
nor U7693 (N_7693,N_2825,N_2819);
nand U7694 (N_7694,N_1478,N_3013);
nor U7695 (N_7695,N_3693,N_4752);
or U7696 (N_7696,N_4822,N_2889);
or U7697 (N_7697,N_2118,N_1773);
or U7698 (N_7698,N_1204,N_4727);
or U7699 (N_7699,N_1027,N_317);
nand U7700 (N_7700,N_2470,N_4297);
or U7701 (N_7701,N_851,N_2947);
nand U7702 (N_7702,N_4268,N_4041);
nand U7703 (N_7703,N_3076,N_1313);
nor U7704 (N_7704,N_3827,N_3121);
nand U7705 (N_7705,N_1103,N_82);
and U7706 (N_7706,N_2712,N_4535);
and U7707 (N_7707,N_2403,N_4434);
nor U7708 (N_7708,N_4367,N_1623);
and U7709 (N_7709,N_3789,N_4990);
and U7710 (N_7710,N_1376,N_3539);
and U7711 (N_7711,N_129,N_4760);
xor U7712 (N_7712,N_2231,N_1699);
nand U7713 (N_7713,N_3981,N_431);
nor U7714 (N_7714,N_1031,N_3801);
and U7715 (N_7715,N_3534,N_4287);
nor U7716 (N_7716,N_561,N_4569);
and U7717 (N_7717,N_1421,N_3023);
nand U7718 (N_7718,N_1289,N_4483);
nor U7719 (N_7719,N_3104,N_419);
or U7720 (N_7720,N_3020,N_710);
nor U7721 (N_7721,N_2374,N_2349);
and U7722 (N_7722,N_1201,N_1779);
or U7723 (N_7723,N_3843,N_306);
nor U7724 (N_7724,N_687,N_446);
nor U7725 (N_7725,N_3558,N_1739);
nand U7726 (N_7726,N_3081,N_1246);
and U7727 (N_7727,N_834,N_3352);
xnor U7728 (N_7728,N_3418,N_3347);
nor U7729 (N_7729,N_973,N_3910);
nor U7730 (N_7730,N_1532,N_352);
and U7731 (N_7731,N_3491,N_4395);
xor U7732 (N_7732,N_3876,N_4995);
nand U7733 (N_7733,N_2091,N_2350);
or U7734 (N_7734,N_4013,N_2);
nand U7735 (N_7735,N_2234,N_1916);
nand U7736 (N_7736,N_3716,N_4338);
nor U7737 (N_7737,N_3647,N_1317);
and U7738 (N_7738,N_1317,N_3741);
nand U7739 (N_7739,N_1165,N_4356);
and U7740 (N_7740,N_4204,N_1413);
nand U7741 (N_7741,N_2260,N_3568);
nand U7742 (N_7742,N_709,N_1752);
and U7743 (N_7743,N_2339,N_429);
and U7744 (N_7744,N_1522,N_2659);
or U7745 (N_7745,N_49,N_1341);
or U7746 (N_7746,N_1442,N_1166);
nor U7747 (N_7747,N_826,N_2186);
nor U7748 (N_7748,N_1076,N_3133);
nor U7749 (N_7749,N_1058,N_2720);
nand U7750 (N_7750,N_1283,N_1175);
or U7751 (N_7751,N_146,N_344);
and U7752 (N_7752,N_4075,N_1443);
and U7753 (N_7753,N_4532,N_1334);
nand U7754 (N_7754,N_1318,N_827);
nand U7755 (N_7755,N_592,N_2210);
nor U7756 (N_7756,N_2291,N_3892);
or U7757 (N_7757,N_757,N_129);
and U7758 (N_7758,N_1254,N_1663);
nor U7759 (N_7759,N_1045,N_4544);
nand U7760 (N_7760,N_3647,N_4439);
and U7761 (N_7761,N_4153,N_1048);
or U7762 (N_7762,N_2829,N_3139);
and U7763 (N_7763,N_2405,N_4196);
and U7764 (N_7764,N_4175,N_473);
nand U7765 (N_7765,N_1625,N_4970);
nand U7766 (N_7766,N_4335,N_3165);
and U7767 (N_7767,N_2212,N_4688);
nor U7768 (N_7768,N_3984,N_1764);
nand U7769 (N_7769,N_4605,N_1055);
or U7770 (N_7770,N_550,N_3190);
nor U7771 (N_7771,N_4426,N_2286);
nand U7772 (N_7772,N_3570,N_4162);
nand U7773 (N_7773,N_4824,N_1136);
or U7774 (N_7774,N_4527,N_1253);
nor U7775 (N_7775,N_1837,N_1167);
and U7776 (N_7776,N_760,N_1256);
nor U7777 (N_7777,N_3356,N_3247);
or U7778 (N_7778,N_665,N_688);
or U7779 (N_7779,N_4532,N_2664);
and U7780 (N_7780,N_3258,N_2488);
nor U7781 (N_7781,N_3727,N_2570);
nor U7782 (N_7782,N_2781,N_3767);
xnor U7783 (N_7783,N_154,N_469);
or U7784 (N_7784,N_2760,N_2980);
nand U7785 (N_7785,N_2309,N_3928);
or U7786 (N_7786,N_4896,N_98);
nor U7787 (N_7787,N_2346,N_1578);
nor U7788 (N_7788,N_2063,N_3772);
nand U7789 (N_7789,N_3673,N_314);
or U7790 (N_7790,N_3080,N_3056);
and U7791 (N_7791,N_2180,N_1660);
and U7792 (N_7792,N_1925,N_3083);
nor U7793 (N_7793,N_2060,N_265);
nand U7794 (N_7794,N_4929,N_863);
nor U7795 (N_7795,N_1257,N_840);
or U7796 (N_7796,N_3,N_2261);
nand U7797 (N_7797,N_3673,N_1268);
or U7798 (N_7798,N_1120,N_1806);
nand U7799 (N_7799,N_4847,N_1230);
nor U7800 (N_7800,N_3509,N_4605);
or U7801 (N_7801,N_1851,N_4631);
nor U7802 (N_7802,N_2428,N_957);
nor U7803 (N_7803,N_4360,N_1070);
and U7804 (N_7804,N_3971,N_4692);
nor U7805 (N_7805,N_3111,N_721);
or U7806 (N_7806,N_2153,N_3664);
nor U7807 (N_7807,N_1445,N_3162);
nor U7808 (N_7808,N_2500,N_3377);
and U7809 (N_7809,N_2600,N_3280);
nand U7810 (N_7810,N_1265,N_2907);
and U7811 (N_7811,N_2641,N_4754);
and U7812 (N_7812,N_2548,N_3954);
nand U7813 (N_7813,N_440,N_2859);
nor U7814 (N_7814,N_2508,N_3948);
nand U7815 (N_7815,N_767,N_4369);
xnor U7816 (N_7816,N_3653,N_2257);
and U7817 (N_7817,N_2403,N_3249);
nor U7818 (N_7818,N_965,N_3279);
nand U7819 (N_7819,N_3048,N_371);
or U7820 (N_7820,N_4873,N_1339);
and U7821 (N_7821,N_4323,N_4546);
nand U7822 (N_7822,N_1454,N_848);
or U7823 (N_7823,N_603,N_2142);
nor U7824 (N_7824,N_471,N_920);
nor U7825 (N_7825,N_1267,N_1039);
and U7826 (N_7826,N_4304,N_3277);
nor U7827 (N_7827,N_473,N_2279);
or U7828 (N_7828,N_3585,N_1901);
nand U7829 (N_7829,N_2177,N_3008);
nor U7830 (N_7830,N_1334,N_4062);
or U7831 (N_7831,N_3059,N_4154);
or U7832 (N_7832,N_80,N_1546);
or U7833 (N_7833,N_2514,N_2255);
nand U7834 (N_7834,N_1010,N_4908);
nand U7835 (N_7835,N_2990,N_1422);
nor U7836 (N_7836,N_2795,N_1949);
nand U7837 (N_7837,N_2037,N_4448);
and U7838 (N_7838,N_366,N_3979);
nand U7839 (N_7839,N_1405,N_2767);
nand U7840 (N_7840,N_1852,N_2677);
or U7841 (N_7841,N_1619,N_2438);
or U7842 (N_7842,N_302,N_3093);
and U7843 (N_7843,N_3422,N_4102);
nor U7844 (N_7844,N_3462,N_2090);
and U7845 (N_7845,N_866,N_1174);
nand U7846 (N_7846,N_1205,N_2052);
nand U7847 (N_7847,N_4660,N_478);
nor U7848 (N_7848,N_593,N_1753);
nand U7849 (N_7849,N_2851,N_4413);
nor U7850 (N_7850,N_3382,N_3059);
nand U7851 (N_7851,N_4154,N_2219);
nor U7852 (N_7852,N_1185,N_1912);
or U7853 (N_7853,N_508,N_3360);
or U7854 (N_7854,N_2205,N_2537);
xnor U7855 (N_7855,N_4258,N_2781);
and U7856 (N_7856,N_915,N_689);
or U7857 (N_7857,N_164,N_1553);
nor U7858 (N_7858,N_4828,N_1920);
and U7859 (N_7859,N_4481,N_1931);
nand U7860 (N_7860,N_756,N_1422);
nor U7861 (N_7861,N_1829,N_2637);
nor U7862 (N_7862,N_4073,N_2959);
nor U7863 (N_7863,N_3789,N_1203);
or U7864 (N_7864,N_645,N_4980);
or U7865 (N_7865,N_2919,N_3748);
nand U7866 (N_7866,N_3026,N_2425);
nand U7867 (N_7867,N_2641,N_3975);
and U7868 (N_7868,N_934,N_3339);
nor U7869 (N_7869,N_4563,N_603);
or U7870 (N_7870,N_354,N_3801);
nor U7871 (N_7871,N_406,N_1886);
nor U7872 (N_7872,N_870,N_4583);
or U7873 (N_7873,N_680,N_3974);
or U7874 (N_7874,N_3251,N_1240);
nand U7875 (N_7875,N_2500,N_3222);
nor U7876 (N_7876,N_1332,N_3598);
and U7877 (N_7877,N_3833,N_3611);
nor U7878 (N_7878,N_4628,N_1522);
or U7879 (N_7879,N_3424,N_3284);
nor U7880 (N_7880,N_4212,N_3765);
and U7881 (N_7881,N_744,N_4774);
nor U7882 (N_7882,N_3521,N_3108);
xor U7883 (N_7883,N_13,N_2194);
nor U7884 (N_7884,N_1170,N_4043);
nor U7885 (N_7885,N_2791,N_4925);
nor U7886 (N_7886,N_1055,N_1474);
nand U7887 (N_7887,N_688,N_1950);
and U7888 (N_7888,N_3727,N_3204);
nor U7889 (N_7889,N_1663,N_1690);
nor U7890 (N_7890,N_77,N_1688);
or U7891 (N_7891,N_2986,N_4117);
nor U7892 (N_7892,N_3573,N_697);
nand U7893 (N_7893,N_2929,N_3647);
nand U7894 (N_7894,N_4856,N_1021);
nand U7895 (N_7895,N_1972,N_4732);
nor U7896 (N_7896,N_2958,N_3869);
or U7897 (N_7897,N_3589,N_3953);
and U7898 (N_7898,N_4453,N_1872);
and U7899 (N_7899,N_864,N_4886);
and U7900 (N_7900,N_3018,N_716);
nor U7901 (N_7901,N_661,N_1638);
and U7902 (N_7902,N_914,N_4920);
and U7903 (N_7903,N_4721,N_1042);
nor U7904 (N_7904,N_1851,N_4248);
nand U7905 (N_7905,N_1939,N_2357);
or U7906 (N_7906,N_4964,N_632);
nand U7907 (N_7907,N_4725,N_1624);
and U7908 (N_7908,N_3305,N_2339);
nor U7909 (N_7909,N_3912,N_4398);
nand U7910 (N_7910,N_1915,N_1858);
nor U7911 (N_7911,N_3403,N_4146);
nor U7912 (N_7912,N_2230,N_461);
and U7913 (N_7913,N_4362,N_4023);
and U7914 (N_7914,N_1291,N_1518);
and U7915 (N_7915,N_461,N_573);
or U7916 (N_7916,N_2216,N_1566);
or U7917 (N_7917,N_961,N_3606);
nor U7918 (N_7918,N_42,N_3248);
nor U7919 (N_7919,N_3572,N_4429);
and U7920 (N_7920,N_1554,N_1176);
nand U7921 (N_7921,N_3203,N_1214);
or U7922 (N_7922,N_1597,N_1967);
or U7923 (N_7923,N_2199,N_4612);
or U7924 (N_7924,N_4154,N_1018);
nor U7925 (N_7925,N_1,N_1454);
and U7926 (N_7926,N_3349,N_4053);
nand U7927 (N_7927,N_2602,N_1080);
nand U7928 (N_7928,N_4967,N_4620);
and U7929 (N_7929,N_4987,N_4186);
or U7930 (N_7930,N_3237,N_3235);
nand U7931 (N_7931,N_2004,N_4709);
nor U7932 (N_7932,N_3564,N_2224);
and U7933 (N_7933,N_594,N_1040);
nor U7934 (N_7934,N_2138,N_328);
nor U7935 (N_7935,N_3456,N_1675);
and U7936 (N_7936,N_4162,N_4295);
nand U7937 (N_7937,N_1298,N_3075);
or U7938 (N_7938,N_309,N_4489);
nand U7939 (N_7939,N_2868,N_3766);
or U7940 (N_7940,N_2625,N_40);
nand U7941 (N_7941,N_1952,N_687);
or U7942 (N_7942,N_4836,N_1022);
and U7943 (N_7943,N_3011,N_1348);
nor U7944 (N_7944,N_518,N_262);
and U7945 (N_7945,N_2951,N_4624);
nand U7946 (N_7946,N_2732,N_3169);
nor U7947 (N_7947,N_1197,N_2931);
nand U7948 (N_7948,N_2380,N_2926);
nor U7949 (N_7949,N_208,N_2898);
or U7950 (N_7950,N_136,N_4027);
and U7951 (N_7951,N_865,N_2439);
and U7952 (N_7952,N_1062,N_741);
nand U7953 (N_7953,N_3994,N_1374);
nand U7954 (N_7954,N_1117,N_727);
nand U7955 (N_7955,N_2135,N_2146);
nor U7956 (N_7956,N_458,N_1626);
or U7957 (N_7957,N_4993,N_3907);
xnor U7958 (N_7958,N_3442,N_2900);
or U7959 (N_7959,N_2085,N_348);
nand U7960 (N_7960,N_3174,N_1464);
nand U7961 (N_7961,N_1760,N_2864);
and U7962 (N_7962,N_1446,N_4799);
or U7963 (N_7963,N_2440,N_321);
nand U7964 (N_7964,N_3231,N_1885);
nand U7965 (N_7965,N_4535,N_2662);
nand U7966 (N_7966,N_2318,N_301);
or U7967 (N_7967,N_271,N_4813);
nor U7968 (N_7968,N_1801,N_4523);
nor U7969 (N_7969,N_1458,N_275);
nand U7970 (N_7970,N_1463,N_3487);
nand U7971 (N_7971,N_3255,N_3942);
nor U7972 (N_7972,N_2462,N_1303);
nor U7973 (N_7973,N_4476,N_1442);
or U7974 (N_7974,N_1106,N_3241);
or U7975 (N_7975,N_3964,N_4340);
nor U7976 (N_7976,N_2986,N_2612);
nor U7977 (N_7977,N_2913,N_3723);
or U7978 (N_7978,N_4877,N_3811);
or U7979 (N_7979,N_2095,N_4553);
and U7980 (N_7980,N_208,N_1578);
and U7981 (N_7981,N_515,N_488);
nor U7982 (N_7982,N_326,N_798);
and U7983 (N_7983,N_1637,N_3600);
and U7984 (N_7984,N_1105,N_1113);
or U7985 (N_7985,N_3383,N_1159);
or U7986 (N_7986,N_3344,N_1651);
nand U7987 (N_7987,N_1623,N_554);
nor U7988 (N_7988,N_3704,N_4081);
nand U7989 (N_7989,N_425,N_2079);
nand U7990 (N_7990,N_3201,N_1877);
xor U7991 (N_7991,N_3654,N_4478);
nor U7992 (N_7992,N_1518,N_3365);
nand U7993 (N_7993,N_2708,N_2080);
nand U7994 (N_7994,N_2910,N_2683);
nor U7995 (N_7995,N_1462,N_3619);
and U7996 (N_7996,N_4081,N_1117);
xnor U7997 (N_7997,N_1766,N_2839);
and U7998 (N_7998,N_1302,N_4914);
nor U7999 (N_7999,N_2874,N_1908);
or U8000 (N_8000,N_4257,N_3877);
nor U8001 (N_8001,N_1792,N_2980);
and U8002 (N_8002,N_4756,N_1320);
nand U8003 (N_8003,N_3602,N_4537);
or U8004 (N_8004,N_3024,N_4828);
nand U8005 (N_8005,N_608,N_306);
and U8006 (N_8006,N_2398,N_3475);
nand U8007 (N_8007,N_3956,N_1755);
or U8008 (N_8008,N_2574,N_2014);
nand U8009 (N_8009,N_936,N_2774);
nor U8010 (N_8010,N_3641,N_818);
nand U8011 (N_8011,N_525,N_2739);
and U8012 (N_8012,N_4367,N_1775);
and U8013 (N_8013,N_4582,N_3987);
nor U8014 (N_8014,N_2139,N_4299);
nor U8015 (N_8015,N_519,N_1545);
nor U8016 (N_8016,N_4200,N_1456);
nor U8017 (N_8017,N_3667,N_3796);
nand U8018 (N_8018,N_1566,N_4793);
nand U8019 (N_8019,N_1079,N_4374);
nand U8020 (N_8020,N_4235,N_194);
nand U8021 (N_8021,N_3722,N_610);
nand U8022 (N_8022,N_1790,N_4960);
and U8023 (N_8023,N_2768,N_4472);
or U8024 (N_8024,N_2085,N_4300);
and U8025 (N_8025,N_2436,N_2871);
nand U8026 (N_8026,N_1203,N_3854);
or U8027 (N_8027,N_2534,N_2990);
or U8028 (N_8028,N_1486,N_3552);
and U8029 (N_8029,N_3225,N_1315);
nor U8030 (N_8030,N_4438,N_731);
nor U8031 (N_8031,N_4958,N_2212);
nand U8032 (N_8032,N_2160,N_2700);
nand U8033 (N_8033,N_3598,N_3574);
and U8034 (N_8034,N_4372,N_4298);
or U8035 (N_8035,N_442,N_1337);
nand U8036 (N_8036,N_1660,N_3239);
or U8037 (N_8037,N_1789,N_1405);
or U8038 (N_8038,N_2954,N_3431);
and U8039 (N_8039,N_1536,N_1812);
nand U8040 (N_8040,N_2167,N_46);
nand U8041 (N_8041,N_1480,N_1554);
nand U8042 (N_8042,N_1103,N_3317);
or U8043 (N_8043,N_4579,N_2372);
and U8044 (N_8044,N_2330,N_418);
and U8045 (N_8045,N_2512,N_4900);
or U8046 (N_8046,N_1276,N_3858);
nand U8047 (N_8047,N_1061,N_4676);
and U8048 (N_8048,N_2091,N_4070);
nand U8049 (N_8049,N_3886,N_4193);
nand U8050 (N_8050,N_962,N_4245);
nor U8051 (N_8051,N_1269,N_1362);
nand U8052 (N_8052,N_3276,N_362);
nor U8053 (N_8053,N_2689,N_3945);
nor U8054 (N_8054,N_1926,N_2729);
and U8055 (N_8055,N_1061,N_995);
nand U8056 (N_8056,N_3381,N_4979);
nand U8057 (N_8057,N_4083,N_3835);
and U8058 (N_8058,N_2051,N_739);
nand U8059 (N_8059,N_3509,N_2629);
nand U8060 (N_8060,N_1327,N_3941);
or U8061 (N_8061,N_3315,N_4728);
and U8062 (N_8062,N_3412,N_3637);
and U8063 (N_8063,N_2303,N_975);
or U8064 (N_8064,N_2246,N_4401);
or U8065 (N_8065,N_1974,N_90);
nor U8066 (N_8066,N_2557,N_4120);
nand U8067 (N_8067,N_1837,N_3207);
or U8068 (N_8068,N_3432,N_104);
or U8069 (N_8069,N_1448,N_2930);
nor U8070 (N_8070,N_282,N_573);
nor U8071 (N_8071,N_2659,N_2291);
nand U8072 (N_8072,N_79,N_111);
nand U8073 (N_8073,N_2282,N_1018);
nand U8074 (N_8074,N_1119,N_2616);
nand U8075 (N_8075,N_88,N_481);
nand U8076 (N_8076,N_2121,N_3889);
nand U8077 (N_8077,N_844,N_1270);
nor U8078 (N_8078,N_3723,N_2308);
nor U8079 (N_8079,N_1509,N_1290);
and U8080 (N_8080,N_1105,N_1396);
nor U8081 (N_8081,N_3496,N_2098);
and U8082 (N_8082,N_232,N_3666);
or U8083 (N_8083,N_3519,N_3755);
nor U8084 (N_8084,N_4655,N_3416);
nor U8085 (N_8085,N_2061,N_2301);
nand U8086 (N_8086,N_356,N_2529);
nor U8087 (N_8087,N_3858,N_4184);
or U8088 (N_8088,N_2230,N_2719);
nor U8089 (N_8089,N_726,N_1911);
nor U8090 (N_8090,N_148,N_301);
nor U8091 (N_8091,N_2257,N_4583);
and U8092 (N_8092,N_1575,N_4003);
nor U8093 (N_8093,N_4911,N_36);
nand U8094 (N_8094,N_3237,N_4065);
or U8095 (N_8095,N_940,N_4585);
nand U8096 (N_8096,N_2463,N_1462);
and U8097 (N_8097,N_4475,N_2410);
nor U8098 (N_8098,N_4907,N_3694);
or U8099 (N_8099,N_1505,N_2063);
and U8100 (N_8100,N_2701,N_3081);
nor U8101 (N_8101,N_2614,N_935);
nor U8102 (N_8102,N_2332,N_1887);
nand U8103 (N_8103,N_3285,N_4108);
and U8104 (N_8104,N_424,N_229);
and U8105 (N_8105,N_279,N_500);
nand U8106 (N_8106,N_2981,N_1964);
nor U8107 (N_8107,N_132,N_135);
and U8108 (N_8108,N_154,N_4567);
nor U8109 (N_8109,N_1281,N_4686);
or U8110 (N_8110,N_2271,N_1630);
nand U8111 (N_8111,N_4211,N_2803);
nor U8112 (N_8112,N_4426,N_2534);
or U8113 (N_8113,N_2463,N_1300);
nand U8114 (N_8114,N_3498,N_2906);
nand U8115 (N_8115,N_1395,N_2777);
and U8116 (N_8116,N_829,N_1502);
or U8117 (N_8117,N_3132,N_246);
or U8118 (N_8118,N_4616,N_3926);
or U8119 (N_8119,N_4440,N_1572);
nor U8120 (N_8120,N_1777,N_4912);
or U8121 (N_8121,N_4910,N_546);
or U8122 (N_8122,N_3589,N_4982);
or U8123 (N_8123,N_2294,N_257);
and U8124 (N_8124,N_1652,N_2023);
nor U8125 (N_8125,N_1550,N_4630);
nor U8126 (N_8126,N_887,N_2851);
or U8127 (N_8127,N_3597,N_4572);
and U8128 (N_8128,N_1305,N_472);
nor U8129 (N_8129,N_3932,N_3827);
and U8130 (N_8130,N_32,N_857);
and U8131 (N_8131,N_937,N_3616);
nor U8132 (N_8132,N_120,N_3344);
nand U8133 (N_8133,N_4339,N_1557);
and U8134 (N_8134,N_1674,N_4800);
or U8135 (N_8135,N_1554,N_1460);
nand U8136 (N_8136,N_300,N_4128);
nand U8137 (N_8137,N_1933,N_496);
or U8138 (N_8138,N_2760,N_2425);
and U8139 (N_8139,N_2596,N_4358);
and U8140 (N_8140,N_4092,N_1793);
or U8141 (N_8141,N_2802,N_1219);
and U8142 (N_8142,N_4463,N_2062);
nor U8143 (N_8143,N_1696,N_1453);
nand U8144 (N_8144,N_712,N_4864);
nand U8145 (N_8145,N_2311,N_4579);
nand U8146 (N_8146,N_769,N_2900);
nand U8147 (N_8147,N_3344,N_1099);
nand U8148 (N_8148,N_1357,N_3783);
or U8149 (N_8149,N_4139,N_1686);
and U8150 (N_8150,N_3806,N_1094);
nand U8151 (N_8151,N_1380,N_2943);
xor U8152 (N_8152,N_3869,N_3022);
nand U8153 (N_8153,N_3627,N_3);
nand U8154 (N_8154,N_1938,N_4567);
nor U8155 (N_8155,N_384,N_2254);
nand U8156 (N_8156,N_1622,N_4770);
nor U8157 (N_8157,N_4619,N_4310);
nand U8158 (N_8158,N_3008,N_973);
nand U8159 (N_8159,N_63,N_1293);
or U8160 (N_8160,N_3821,N_896);
and U8161 (N_8161,N_602,N_1211);
and U8162 (N_8162,N_1587,N_2111);
nand U8163 (N_8163,N_1984,N_42);
nor U8164 (N_8164,N_520,N_4247);
and U8165 (N_8165,N_4504,N_3421);
nand U8166 (N_8166,N_981,N_2084);
nor U8167 (N_8167,N_2715,N_4855);
and U8168 (N_8168,N_2795,N_600);
nand U8169 (N_8169,N_3985,N_2275);
nand U8170 (N_8170,N_741,N_1128);
or U8171 (N_8171,N_4974,N_1995);
nor U8172 (N_8172,N_2749,N_4101);
nand U8173 (N_8173,N_4366,N_3525);
and U8174 (N_8174,N_7,N_38);
and U8175 (N_8175,N_4349,N_4417);
nand U8176 (N_8176,N_1884,N_1757);
or U8177 (N_8177,N_3453,N_2108);
and U8178 (N_8178,N_2627,N_1306);
nand U8179 (N_8179,N_3676,N_3027);
nand U8180 (N_8180,N_3467,N_3748);
and U8181 (N_8181,N_1805,N_2128);
or U8182 (N_8182,N_1286,N_843);
and U8183 (N_8183,N_35,N_1418);
nor U8184 (N_8184,N_998,N_4979);
nand U8185 (N_8185,N_4808,N_4303);
or U8186 (N_8186,N_4320,N_3390);
nor U8187 (N_8187,N_1866,N_2432);
nor U8188 (N_8188,N_3279,N_1554);
or U8189 (N_8189,N_1767,N_2549);
nor U8190 (N_8190,N_1050,N_1109);
nor U8191 (N_8191,N_4821,N_1017);
or U8192 (N_8192,N_4190,N_4170);
nor U8193 (N_8193,N_4921,N_3227);
nor U8194 (N_8194,N_2472,N_1138);
or U8195 (N_8195,N_1411,N_1258);
or U8196 (N_8196,N_2220,N_2720);
and U8197 (N_8197,N_4869,N_2808);
nand U8198 (N_8198,N_3363,N_762);
or U8199 (N_8199,N_2098,N_1774);
and U8200 (N_8200,N_3077,N_3155);
nand U8201 (N_8201,N_2667,N_1494);
nor U8202 (N_8202,N_1456,N_3216);
or U8203 (N_8203,N_51,N_2188);
or U8204 (N_8204,N_3959,N_1819);
or U8205 (N_8205,N_4577,N_1242);
nor U8206 (N_8206,N_4205,N_569);
and U8207 (N_8207,N_605,N_3756);
and U8208 (N_8208,N_3342,N_2328);
or U8209 (N_8209,N_3761,N_1553);
and U8210 (N_8210,N_3768,N_3830);
and U8211 (N_8211,N_2622,N_3525);
nand U8212 (N_8212,N_2630,N_1278);
nand U8213 (N_8213,N_766,N_1821);
or U8214 (N_8214,N_2575,N_1304);
nand U8215 (N_8215,N_4325,N_4797);
nor U8216 (N_8216,N_4236,N_1407);
or U8217 (N_8217,N_4613,N_2177);
or U8218 (N_8218,N_1525,N_2755);
nand U8219 (N_8219,N_8,N_563);
or U8220 (N_8220,N_1317,N_1319);
nand U8221 (N_8221,N_2293,N_2955);
and U8222 (N_8222,N_4714,N_1887);
and U8223 (N_8223,N_4582,N_1981);
and U8224 (N_8224,N_379,N_1586);
and U8225 (N_8225,N_2838,N_1542);
or U8226 (N_8226,N_1469,N_3850);
and U8227 (N_8227,N_2838,N_3760);
nand U8228 (N_8228,N_1932,N_570);
nand U8229 (N_8229,N_4277,N_950);
nor U8230 (N_8230,N_597,N_1756);
nand U8231 (N_8231,N_3555,N_2273);
and U8232 (N_8232,N_2386,N_1592);
nand U8233 (N_8233,N_2063,N_223);
and U8234 (N_8234,N_2629,N_3427);
nand U8235 (N_8235,N_892,N_4642);
nand U8236 (N_8236,N_4131,N_4610);
nor U8237 (N_8237,N_133,N_144);
or U8238 (N_8238,N_923,N_3994);
nand U8239 (N_8239,N_1344,N_2542);
nand U8240 (N_8240,N_2641,N_340);
or U8241 (N_8241,N_579,N_3269);
and U8242 (N_8242,N_292,N_4851);
and U8243 (N_8243,N_2588,N_4394);
or U8244 (N_8244,N_2785,N_285);
nand U8245 (N_8245,N_1323,N_2236);
or U8246 (N_8246,N_3332,N_762);
nand U8247 (N_8247,N_3597,N_4229);
nand U8248 (N_8248,N_4886,N_4350);
and U8249 (N_8249,N_1863,N_4622);
nand U8250 (N_8250,N_4349,N_1355);
and U8251 (N_8251,N_4897,N_1723);
nor U8252 (N_8252,N_4079,N_2418);
or U8253 (N_8253,N_2214,N_1940);
nor U8254 (N_8254,N_4266,N_4094);
or U8255 (N_8255,N_2716,N_892);
nor U8256 (N_8256,N_4684,N_2685);
and U8257 (N_8257,N_2738,N_1373);
and U8258 (N_8258,N_2063,N_3105);
nor U8259 (N_8259,N_1222,N_1538);
nand U8260 (N_8260,N_434,N_3039);
or U8261 (N_8261,N_2753,N_2831);
or U8262 (N_8262,N_3148,N_3754);
or U8263 (N_8263,N_2812,N_555);
and U8264 (N_8264,N_3940,N_2793);
nand U8265 (N_8265,N_1504,N_1460);
or U8266 (N_8266,N_1884,N_4847);
nand U8267 (N_8267,N_4979,N_2968);
or U8268 (N_8268,N_3023,N_2528);
or U8269 (N_8269,N_4821,N_1639);
nor U8270 (N_8270,N_2068,N_49);
nand U8271 (N_8271,N_4212,N_4877);
nor U8272 (N_8272,N_939,N_2873);
or U8273 (N_8273,N_4895,N_3356);
and U8274 (N_8274,N_3215,N_322);
nor U8275 (N_8275,N_384,N_2392);
and U8276 (N_8276,N_4582,N_1545);
nor U8277 (N_8277,N_3824,N_2883);
nor U8278 (N_8278,N_324,N_4108);
or U8279 (N_8279,N_2153,N_1136);
nand U8280 (N_8280,N_1242,N_697);
nor U8281 (N_8281,N_3526,N_3867);
nand U8282 (N_8282,N_1067,N_2450);
nand U8283 (N_8283,N_2470,N_3474);
or U8284 (N_8284,N_2612,N_4484);
nor U8285 (N_8285,N_4330,N_4308);
and U8286 (N_8286,N_3571,N_4352);
nor U8287 (N_8287,N_535,N_4118);
nor U8288 (N_8288,N_181,N_2896);
nor U8289 (N_8289,N_4308,N_400);
nand U8290 (N_8290,N_2580,N_2088);
nor U8291 (N_8291,N_947,N_1174);
nor U8292 (N_8292,N_1569,N_895);
and U8293 (N_8293,N_923,N_4441);
nor U8294 (N_8294,N_4269,N_3071);
nand U8295 (N_8295,N_2577,N_2670);
nand U8296 (N_8296,N_3147,N_555);
or U8297 (N_8297,N_1563,N_4655);
and U8298 (N_8298,N_225,N_4542);
or U8299 (N_8299,N_3501,N_2540);
nand U8300 (N_8300,N_1151,N_427);
and U8301 (N_8301,N_986,N_4256);
nand U8302 (N_8302,N_335,N_405);
and U8303 (N_8303,N_3271,N_3664);
nand U8304 (N_8304,N_3622,N_4897);
nand U8305 (N_8305,N_4682,N_3967);
nor U8306 (N_8306,N_467,N_3646);
nand U8307 (N_8307,N_1514,N_2973);
and U8308 (N_8308,N_341,N_4038);
or U8309 (N_8309,N_1840,N_3017);
xor U8310 (N_8310,N_3626,N_3096);
nor U8311 (N_8311,N_998,N_3833);
or U8312 (N_8312,N_568,N_2985);
or U8313 (N_8313,N_3057,N_856);
nand U8314 (N_8314,N_3619,N_2523);
nand U8315 (N_8315,N_3075,N_3149);
nor U8316 (N_8316,N_1370,N_4584);
and U8317 (N_8317,N_1023,N_1901);
or U8318 (N_8318,N_2685,N_548);
nand U8319 (N_8319,N_1604,N_4069);
nor U8320 (N_8320,N_83,N_3575);
nand U8321 (N_8321,N_1305,N_2272);
or U8322 (N_8322,N_750,N_3410);
and U8323 (N_8323,N_3746,N_1723);
nand U8324 (N_8324,N_1755,N_554);
nor U8325 (N_8325,N_909,N_1588);
and U8326 (N_8326,N_1388,N_4973);
nand U8327 (N_8327,N_4085,N_2257);
or U8328 (N_8328,N_456,N_1586);
or U8329 (N_8329,N_2208,N_235);
or U8330 (N_8330,N_3685,N_3611);
or U8331 (N_8331,N_2062,N_2038);
nand U8332 (N_8332,N_1769,N_3913);
nand U8333 (N_8333,N_4817,N_148);
nor U8334 (N_8334,N_3273,N_1125);
nand U8335 (N_8335,N_3031,N_3101);
or U8336 (N_8336,N_3762,N_2301);
nand U8337 (N_8337,N_1533,N_4310);
nor U8338 (N_8338,N_2700,N_92);
nor U8339 (N_8339,N_3944,N_14);
nand U8340 (N_8340,N_3049,N_895);
nand U8341 (N_8341,N_1249,N_2807);
or U8342 (N_8342,N_4919,N_1735);
or U8343 (N_8343,N_458,N_77);
and U8344 (N_8344,N_4954,N_2926);
or U8345 (N_8345,N_2225,N_1117);
nand U8346 (N_8346,N_1745,N_4151);
nand U8347 (N_8347,N_2039,N_4397);
and U8348 (N_8348,N_4127,N_274);
nand U8349 (N_8349,N_2651,N_4712);
or U8350 (N_8350,N_3484,N_3534);
or U8351 (N_8351,N_2568,N_2900);
and U8352 (N_8352,N_2363,N_146);
or U8353 (N_8353,N_1397,N_4123);
nand U8354 (N_8354,N_3103,N_761);
and U8355 (N_8355,N_4973,N_4975);
or U8356 (N_8356,N_2536,N_2657);
and U8357 (N_8357,N_764,N_3838);
nor U8358 (N_8358,N_3506,N_266);
or U8359 (N_8359,N_2300,N_2353);
and U8360 (N_8360,N_4099,N_2448);
and U8361 (N_8361,N_1581,N_1189);
nor U8362 (N_8362,N_4691,N_4110);
or U8363 (N_8363,N_3876,N_4376);
nor U8364 (N_8364,N_4979,N_3633);
and U8365 (N_8365,N_4662,N_3827);
or U8366 (N_8366,N_2320,N_2216);
nor U8367 (N_8367,N_1311,N_4740);
and U8368 (N_8368,N_3192,N_1882);
nand U8369 (N_8369,N_4209,N_1429);
or U8370 (N_8370,N_4581,N_1581);
nand U8371 (N_8371,N_663,N_1662);
nor U8372 (N_8372,N_296,N_3980);
nor U8373 (N_8373,N_3160,N_285);
and U8374 (N_8374,N_130,N_2594);
nor U8375 (N_8375,N_1880,N_505);
nor U8376 (N_8376,N_2597,N_805);
nand U8377 (N_8377,N_872,N_4524);
or U8378 (N_8378,N_2596,N_1027);
nand U8379 (N_8379,N_831,N_1327);
or U8380 (N_8380,N_1883,N_4951);
or U8381 (N_8381,N_3566,N_4289);
nor U8382 (N_8382,N_3818,N_4973);
or U8383 (N_8383,N_1479,N_2727);
or U8384 (N_8384,N_2363,N_2490);
or U8385 (N_8385,N_2530,N_4289);
and U8386 (N_8386,N_2534,N_2491);
or U8387 (N_8387,N_3572,N_4683);
and U8388 (N_8388,N_798,N_225);
nand U8389 (N_8389,N_4861,N_3497);
or U8390 (N_8390,N_2799,N_1341);
nand U8391 (N_8391,N_3184,N_363);
nor U8392 (N_8392,N_4726,N_4274);
nor U8393 (N_8393,N_3215,N_2977);
or U8394 (N_8394,N_3759,N_328);
and U8395 (N_8395,N_4449,N_3701);
xnor U8396 (N_8396,N_646,N_57);
nand U8397 (N_8397,N_3399,N_567);
nor U8398 (N_8398,N_2880,N_2916);
xnor U8399 (N_8399,N_3671,N_3309);
and U8400 (N_8400,N_989,N_2150);
nand U8401 (N_8401,N_1077,N_4873);
or U8402 (N_8402,N_2687,N_3153);
nor U8403 (N_8403,N_680,N_2242);
or U8404 (N_8404,N_3641,N_4388);
or U8405 (N_8405,N_4357,N_2264);
or U8406 (N_8406,N_4062,N_2906);
nand U8407 (N_8407,N_4794,N_1884);
or U8408 (N_8408,N_2063,N_2658);
or U8409 (N_8409,N_3263,N_2781);
nor U8410 (N_8410,N_2627,N_1119);
nor U8411 (N_8411,N_126,N_2224);
or U8412 (N_8412,N_1465,N_4877);
or U8413 (N_8413,N_4000,N_3926);
nor U8414 (N_8414,N_1153,N_441);
nor U8415 (N_8415,N_4730,N_2387);
nor U8416 (N_8416,N_3393,N_983);
and U8417 (N_8417,N_2505,N_1213);
nand U8418 (N_8418,N_3731,N_290);
nand U8419 (N_8419,N_4091,N_1829);
nand U8420 (N_8420,N_3416,N_2849);
nor U8421 (N_8421,N_4432,N_2298);
and U8422 (N_8422,N_2533,N_1028);
nand U8423 (N_8423,N_723,N_3490);
and U8424 (N_8424,N_1403,N_2051);
nor U8425 (N_8425,N_3863,N_1167);
nand U8426 (N_8426,N_3774,N_3353);
and U8427 (N_8427,N_3226,N_3640);
nand U8428 (N_8428,N_2551,N_4046);
or U8429 (N_8429,N_3294,N_3342);
and U8430 (N_8430,N_817,N_3602);
nand U8431 (N_8431,N_978,N_1500);
nor U8432 (N_8432,N_1713,N_1728);
nor U8433 (N_8433,N_2410,N_1512);
nor U8434 (N_8434,N_761,N_1995);
nor U8435 (N_8435,N_3071,N_4343);
nand U8436 (N_8436,N_4622,N_4766);
nor U8437 (N_8437,N_3286,N_1999);
and U8438 (N_8438,N_4215,N_1208);
and U8439 (N_8439,N_4313,N_3738);
and U8440 (N_8440,N_101,N_2432);
nor U8441 (N_8441,N_4495,N_4054);
and U8442 (N_8442,N_3390,N_2524);
nor U8443 (N_8443,N_4133,N_1798);
or U8444 (N_8444,N_827,N_1280);
or U8445 (N_8445,N_2070,N_4677);
and U8446 (N_8446,N_3768,N_3444);
nand U8447 (N_8447,N_2306,N_3502);
and U8448 (N_8448,N_3580,N_1376);
nor U8449 (N_8449,N_871,N_1208);
nand U8450 (N_8450,N_2564,N_3219);
nand U8451 (N_8451,N_4010,N_3411);
and U8452 (N_8452,N_681,N_378);
nor U8453 (N_8453,N_4033,N_3486);
nor U8454 (N_8454,N_2466,N_4458);
nand U8455 (N_8455,N_1198,N_1597);
nor U8456 (N_8456,N_3374,N_3543);
nor U8457 (N_8457,N_1476,N_4523);
or U8458 (N_8458,N_2739,N_3546);
nor U8459 (N_8459,N_4917,N_718);
and U8460 (N_8460,N_3907,N_1826);
nor U8461 (N_8461,N_3727,N_3236);
and U8462 (N_8462,N_4588,N_1554);
or U8463 (N_8463,N_3946,N_2186);
nand U8464 (N_8464,N_4883,N_3539);
nor U8465 (N_8465,N_408,N_270);
nand U8466 (N_8466,N_2893,N_1547);
or U8467 (N_8467,N_2409,N_4673);
and U8468 (N_8468,N_2110,N_4017);
nor U8469 (N_8469,N_3359,N_3810);
nor U8470 (N_8470,N_4923,N_4989);
and U8471 (N_8471,N_3537,N_4448);
nor U8472 (N_8472,N_4446,N_885);
nor U8473 (N_8473,N_802,N_2639);
nand U8474 (N_8474,N_4621,N_4111);
and U8475 (N_8475,N_4250,N_444);
nor U8476 (N_8476,N_4310,N_274);
and U8477 (N_8477,N_1401,N_1782);
nor U8478 (N_8478,N_1641,N_4269);
nor U8479 (N_8479,N_4497,N_1532);
nor U8480 (N_8480,N_4936,N_2544);
nor U8481 (N_8481,N_2017,N_4605);
and U8482 (N_8482,N_4078,N_1622);
and U8483 (N_8483,N_4247,N_4801);
nand U8484 (N_8484,N_613,N_331);
or U8485 (N_8485,N_3060,N_3269);
or U8486 (N_8486,N_3728,N_3678);
nand U8487 (N_8487,N_2977,N_2527);
nor U8488 (N_8488,N_4823,N_48);
nand U8489 (N_8489,N_781,N_2436);
and U8490 (N_8490,N_3933,N_2600);
nor U8491 (N_8491,N_2959,N_2236);
nand U8492 (N_8492,N_3033,N_3531);
nor U8493 (N_8493,N_3886,N_1123);
nand U8494 (N_8494,N_834,N_2652);
or U8495 (N_8495,N_4118,N_2930);
and U8496 (N_8496,N_4635,N_4028);
nor U8497 (N_8497,N_140,N_2588);
nand U8498 (N_8498,N_3203,N_4586);
or U8499 (N_8499,N_3933,N_3528);
or U8500 (N_8500,N_2160,N_4244);
nand U8501 (N_8501,N_3796,N_599);
xor U8502 (N_8502,N_2364,N_2888);
or U8503 (N_8503,N_1780,N_4506);
or U8504 (N_8504,N_2139,N_3310);
nand U8505 (N_8505,N_2082,N_1619);
nand U8506 (N_8506,N_682,N_3280);
nand U8507 (N_8507,N_3505,N_4227);
and U8508 (N_8508,N_2950,N_4746);
nand U8509 (N_8509,N_2398,N_4982);
nand U8510 (N_8510,N_2315,N_1673);
nor U8511 (N_8511,N_1494,N_2027);
nor U8512 (N_8512,N_615,N_3576);
or U8513 (N_8513,N_354,N_745);
or U8514 (N_8514,N_2064,N_1820);
and U8515 (N_8515,N_1655,N_3363);
and U8516 (N_8516,N_734,N_3375);
nor U8517 (N_8517,N_2421,N_4468);
nand U8518 (N_8518,N_95,N_3427);
or U8519 (N_8519,N_219,N_729);
nor U8520 (N_8520,N_1850,N_4095);
nand U8521 (N_8521,N_2277,N_1403);
nand U8522 (N_8522,N_1257,N_1214);
and U8523 (N_8523,N_2729,N_3029);
or U8524 (N_8524,N_2804,N_4111);
nand U8525 (N_8525,N_4705,N_1472);
or U8526 (N_8526,N_2651,N_936);
and U8527 (N_8527,N_190,N_1488);
or U8528 (N_8528,N_2139,N_2416);
nand U8529 (N_8529,N_4068,N_3532);
nand U8530 (N_8530,N_4731,N_2544);
and U8531 (N_8531,N_3137,N_2270);
nor U8532 (N_8532,N_2057,N_4158);
nor U8533 (N_8533,N_2851,N_3617);
and U8534 (N_8534,N_4383,N_3792);
nor U8535 (N_8535,N_3103,N_207);
nand U8536 (N_8536,N_2010,N_3949);
and U8537 (N_8537,N_894,N_2631);
nor U8538 (N_8538,N_3935,N_3988);
and U8539 (N_8539,N_808,N_3957);
nand U8540 (N_8540,N_4835,N_1766);
or U8541 (N_8541,N_4570,N_4029);
or U8542 (N_8542,N_4410,N_4632);
nand U8543 (N_8543,N_3465,N_971);
nor U8544 (N_8544,N_2340,N_1129);
nand U8545 (N_8545,N_483,N_1057);
and U8546 (N_8546,N_4228,N_3489);
nand U8547 (N_8547,N_752,N_990);
or U8548 (N_8548,N_586,N_835);
nor U8549 (N_8549,N_270,N_62);
nor U8550 (N_8550,N_196,N_4437);
nand U8551 (N_8551,N_1348,N_4632);
or U8552 (N_8552,N_3877,N_2532);
or U8553 (N_8553,N_1343,N_2409);
nor U8554 (N_8554,N_3828,N_399);
nor U8555 (N_8555,N_2230,N_4903);
nor U8556 (N_8556,N_209,N_3580);
nor U8557 (N_8557,N_4900,N_4597);
and U8558 (N_8558,N_387,N_3690);
nor U8559 (N_8559,N_2283,N_3405);
nor U8560 (N_8560,N_936,N_3052);
nor U8561 (N_8561,N_851,N_1402);
or U8562 (N_8562,N_2333,N_3196);
and U8563 (N_8563,N_180,N_410);
nor U8564 (N_8564,N_1356,N_392);
nand U8565 (N_8565,N_2678,N_2652);
or U8566 (N_8566,N_3887,N_2311);
or U8567 (N_8567,N_3183,N_4150);
nand U8568 (N_8568,N_4702,N_3790);
nor U8569 (N_8569,N_3814,N_1675);
nand U8570 (N_8570,N_2850,N_2601);
or U8571 (N_8571,N_61,N_3005);
and U8572 (N_8572,N_1158,N_544);
nand U8573 (N_8573,N_1516,N_3811);
and U8574 (N_8574,N_3061,N_4571);
nand U8575 (N_8575,N_2314,N_672);
or U8576 (N_8576,N_1024,N_1549);
or U8577 (N_8577,N_2622,N_4703);
nor U8578 (N_8578,N_3204,N_338);
nand U8579 (N_8579,N_858,N_2753);
and U8580 (N_8580,N_49,N_4631);
nand U8581 (N_8581,N_939,N_1309);
and U8582 (N_8582,N_88,N_4024);
and U8583 (N_8583,N_2893,N_2957);
nand U8584 (N_8584,N_1246,N_178);
nor U8585 (N_8585,N_3995,N_3832);
nand U8586 (N_8586,N_2357,N_2520);
nand U8587 (N_8587,N_2098,N_2357);
or U8588 (N_8588,N_2229,N_2242);
nor U8589 (N_8589,N_4033,N_1118);
and U8590 (N_8590,N_1911,N_1689);
or U8591 (N_8591,N_52,N_1866);
nor U8592 (N_8592,N_4467,N_2182);
nor U8593 (N_8593,N_1711,N_4845);
nand U8594 (N_8594,N_1358,N_549);
nor U8595 (N_8595,N_3143,N_510);
or U8596 (N_8596,N_3710,N_4371);
nor U8597 (N_8597,N_17,N_2679);
or U8598 (N_8598,N_3209,N_2445);
or U8599 (N_8599,N_1454,N_4966);
and U8600 (N_8600,N_2973,N_2787);
and U8601 (N_8601,N_4839,N_3168);
and U8602 (N_8602,N_3915,N_3255);
and U8603 (N_8603,N_4721,N_2087);
or U8604 (N_8604,N_2159,N_1421);
nand U8605 (N_8605,N_4134,N_1909);
or U8606 (N_8606,N_3282,N_4751);
or U8607 (N_8607,N_2922,N_1289);
and U8608 (N_8608,N_303,N_2665);
or U8609 (N_8609,N_2483,N_2864);
or U8610 (N_8610,N_4599,N_3083);
and U8611 (N_8611,N_4111,N_2851);
nor U8612 (N_8612,N_4155,N_1229);
or U8613 (N_8613,N_3104,N_4038);
and U8614 (N_8614,N_2686,N_2581);
or U8615 (N_8615,N_1749,N_3971);
nand U8616 (N_8616,N_906,N_3011);
nand U8617 (N_8617,N_558,N_1551);
nor U8618 (N_8618,N_2987,N_304);
or U8619 (N_8619,N_2791,N_975);
nand U8620 (N_8620,N_3047,N_3670);
or U8621 (N_8621,N_3529,N_1537);
or U8622 (N_8622,N_2419,N_1276);
and U8623 (N_8623,N_1219,N_2037);
nor U8624 (N_8624,N_2922,N_2228);
and U8625 (N_8625,N_2729,N_3334);
or U8626 (N_8626,N_3171,N_2365);
or U8627 (N_8627,N_3076,N_997);
and U8628 (N_8628,N_2003,N_3224);
and U8629 (N_8629,N_1836,N_3908);
nand U8630 (N_8630,N_1226,N_4789);
nand U8631 (N_8631,N_432,N_2740);
or U8632 (N_8632,N_3754,N_4008);
and U8633 (N_8633,N_1402,N_654);
or U8634 (N_8634,N_4178,N_3477);
and U8635 (N_8635,N_1762,N_1454);
nand U8636 (N_8636,N_4425,N_217);
nand U8637 (N_8637,N_273,N_3841);
or U8638 (N_8638,N_4993,N_2249);
or U8639 (N_8639,N_500,N_1857);
nand U8640 (N_8640,N_1001,N_363);
or U8641 (N_8641,N_450,N_434);
and U8642 (N_8642,N_1315,N_508);
and U8643 (N_8643,N_1390,N_4696);
or U8644 (N_8644,N_3897,N_2701);
nor U8645 (N_8645,N_3483,N_3403);
and U8646 (N_8646,N_498,N_1638);
nor U8647 (N_8647,N_4456,N_818);
nor U8648 (N_8648,N_3547,N_736);
nor U8649 (N_8649,N_1539,N_2605);
or U8650 (N_8650,N_3060,N_773);
nand U8651 (N_8651,N_3724,N_4881);
nor U8652 (N_8652,N_286,N_1483);
nand U8653 (N_8653,N_2839,N_436);
nand U8654 (N_8654,N_2207,N_3740);
nor U8655 (N_8655,N_591,N_2945);
nand U8656 (N_8656,N_1588,N_3073);
and U8657 (N_8657,N_4994,N_1718);
and U8658 (N_8658,N_3679,N_4030);
and U8659 (N_8659,N_2152,N_3750);
or U8660 (N_8660,N_4511,N_732);
or U8661 (N_8661,N_674,N_2608);
nand U8662 (N_8662,N_410,N_2907);
nand U8663 (N_8663,N_2049,N_4081);
and U8664 (N_8664,N_273,N_3915);
or U8665 (N_8665,N_3876,N_4577);
nor U8666 (N_8666,N_3593,N_808);
and U8667 (N_8667,N_1242,N_1599);
nor U8668 (N_8668,N_4892,N_1082);
nand U8669 (N_8669,N_764,N_3256);
and U8670 (N_8670,N_1284,N_3990);
or U8671 (N_8671,N_1709,N_965);
nand U8672 (N_8672,N_1833,N_4831);
nor U8673 (N_8673,N_2818,N_3071);
or U8674 (N_8674,N_1303,N_1345);
nor U8675 (N_8675,N_4247,N_1369);
nand U8676 (N_8676,N_1268,N_141);
nand U8677 (N_8677,N_3138,N_4964);
nand U8678 (N_8678,N_2975,N_3486);
and U8679 (N_8679,N_3262,N_980);
and U8680 (N_8680,N_1489,N_4251);
or U8681 (N_8681,N_130,N_4777);
and U8682 (N_8682,N_737,N_4056);
nand U8683 (N_8683,N_246,N_2670);
or U8684 (N_8684,N_3229,N_1630);
nand U8685 (N_8685,N_4922,N_1801);
nor U8686 (N_8686,N_1138,N_3703);
nand U8687 (N_8687,N_3212,N_2034);
or U8688 (N_8688,N_4648,N_1297);
nor U8689 (N_8689,N_2899,N_805);
and U8690 (N_8690,N_2501,N_741);
or U8691 (N_8691,N_687,N_1599);
and U8692 (N_8692,N_710,N_1861);
or U8693 (N_8693,N_4884,N_1471);
or U8694 (N_8694,N_4200,N_2739);
nand U8695 (N_8695,N_2556,N_1597);
nor U8696 (N_8696,N_229,N_4874);
nor U8697 (N_8697,N_3774,N_3857);
nand U8698 (N_8698,N_1874,N_2927);
nor U8699 (N_8699,N_3119,N_4720);
nor U8700 (N_8700,N_3799,N_3221);
nand U8701 (N_8701,N_3977,N_2552);
and U8702 (N_8702,N_4290,N_3360);
nor U8703 (N_8703,N_4787,N_2870);
nand U8704 (N_8704,N_2473,N_2948);
and U8705 (N_8705,N_2296,N_1275);
nand U8706 (N_8706,N_2523,N_156);
and U8707 (N_8707,N_3214,N_1621);
and U8708 (N_8708,N_4701,N_3531);
and U8709 (N_8709,N_2267,N_199);
and U8710 (N_8710,N_4940,N_1901);
nor U8711 (N_8711,N_1576,N_2992);
nor U8712 (N_8712,N_2330,N_712);
and U8713 (N_8713,N_3734,N_1997);
nor U8714 (N_8714,N_2003,N_2611);
nor U8715 (N_8715,N_4303,N_1809);
nor U8716 (N_8716,N_269,N_4280);
or U8717 (N_8717,N_4540,N_1490);
nand U8718 (N_8718,N_627,N_754);
or U8719 (N_8719,N_4493,N_3320);
or U8720 (N_8720,N_4603,N_4763);
xor U8721 (N_8721,N_751,N_1835);
or U8722 (N_8722,N_3301,N_2160);
nor U8723 (N_8723,N_1465,N_4096);
and U8724 (N_8724,N_763,N_1987);
and U8725 (N_8725,N_4711,N_4497);
and U8726 (N_8726,N_2195,N_2978);
nand U8727 (N_8727,N_3860,N_4641);
nor U8728 (N_8728,N_3421,N_2797);
or U8729 (N_8729,N_4233,N_922);
and U8730 (N_8730,N_2748,N_1169);
and U8731 (N_8731,N_2363,N_2999);
nand U8732 (N_8732,N_1852,N_4115);
xnor U8733 (N_8733,N_4522,N_1292);
or U8734 (N_8734,N_1547,N_1209);
or U8735 (N_8735,N_3468,N_824);
nor U8736 (N_8736,N_1197,N_4458);
nand U8737 (N_8737,N_2163,N_459);
and U8738 (N_8738,N_2492,N_2408);
or U8739 (N_8739,N_559,N_803);
and U8740 (N_8740,N_1183,N_2164);
and U8741 (N_8741,N_4357,N_4891);
and U8742 (N_8742,N_246,N_786);
nor U8743 (N_8743,N_4151,N_970);
nand U8744 (N_8744,N_3111,N_3724);
nand U8745 (N_8745,N_560,N_3944);
nand U8746 (N_8746,N_247,N_1692);
nand U8747 (N_8747,N_285,N_3074);
or U8748 (N_8748,N_3864,N_1644);
or U8749 (N_8749,N_4174,N_60);
or U8750 (N_8750,N_1396,N_3557);
or U8751 (N_8751,N_4826,N_4997);
and U8752 (N_8752,N_2805,N_903);
or U8753 (N_8753,N_767,N_908);
nor U8754 (N_8754,N_4902,N_1909);
nor U8755 (N_8755,N_3587,N_4952);
and U8756 (N_8756,N_3591,N_1853);
nand U8757 (N_8757,N_991,N_2787);
and U8758 (N_8758,N_2406,N_267);
nor U8759 (N_8759,N_2236,N_3727);
nor U8760 (N_8760,N_4679,N_518);
or U8761 (N_8761,N_2559,N_1480);
or U8762 (N_8762,N_3087,N_3453);
nor U8763 (N_8763,N_707,N_1518);
and U8764 (N_8764,N_682,N_650);
nor U8765 (N_8765,N_4232,N_4209);
and U8766 (N_8766,N_3369,N_2871);
or U8767 (N_8767,N_4033,N_847);
nor U8768 (N_8768,N_204,N_2088);
or U8769 (N_8769,N_660,N_3736);
and U8770 (N_8770,N_2266,N_3304);
or U8771 (N_8771,N_3780,N_664);
and U8772 (N_8772,N_2609,N_4699);
and U8773 (N_8773,N_1917,N_3524);
and U8774 (N_8774,N_767,N_2475);
or U8775 (N_8775,N_1044,N_4922);
nor U8776 (N_8776,N_4988,N_4511);
and U8777 (N_8777,N_2941,N_4612);
nand U8778 (N_8778,N_4853,N_2460);
and U8779 (N_8779,N_4570,N_2546);
xnor U8780 (N_8780,N_852,N_4135);
or U8781 (N_8781,N_753,N_908);
or U8782 (N_8782,N_2003,N_1713);
nor U8783 (N_8783,N_1783,N_770);
and U8784 (N_8784,N_4728,N_1806);
or U8785 (N_8785,N_4396,N_3468);
and U8786 (N_8786,N_1109,N_4377);
and U8787 (N_8787,N_4173,N_1063);
nor U8788 (N_8788,N_462,N_4062);
xnor U8789 (N_8789,N_330,N_2429);
nand U8790 (N_8790,N_1216,N_2558);
or U8791 (N_8791,N_3933,N_2020);
nand U8792 (N_8792,N_144,N_3461);
or U8793 (N_8793,N_1358,N_843);
nor U8794 (N_8794,N_2314,N_3612);
or U8795 (N_8795,N_3247,N_3690);
xnor U8796 (N_8796,N_324,N_602);
or U8797 (N_8797,N_4023,N_3839);
xor U8798 (N_8798,N_1544,N_296);
and U8799 (N_8799,N_4928,N_4090);
nor U8800 (N_8800,N_417,N_2868);
or U8801 (N_8801,N_1827,N_537);
nor U8802 (N_8802,N_1759,N_1525);
nor U8803 (N_8803,N_290,N_842);
nand U8804 (N_8804,N_1796,N_4715);
and U8805 (N_8805,N_3518,N_1403);
nand U8806 (N_8806,N_316,N_3269);
and U8807 (N_8807,N_3732,N_2099);
or U8808 (N_8808,N_3441,N_552);
and U8809 (N_8809,N_1189,N_2614);
and U8810 (N_8810,N_2914,N_1473);
nand U8811 (N_8811,N_1659,N_767);
or U8812 (N_8812,N_3469,N_4064);
nor U8813 (N_8813,N_981,N_2432);
nor U8814 (N_8814,N_3036,N_2965);
nand U8815 (N_8815,N_2124,N_2108);
and U8816 (N_8816,N_4759,N_3993);
nand U8817 (N_8817,N_2666,N_4195);
nor U8818 (N_8818,N_199,N_652);
nor U8819 (N_8819,N_906,N_648);
or U8820 (N_8820,N_4690,N_836);
nand U8821 (N_8821,N_3490,N_3523);
nor U8822 (N_8822,N_4661,N_2791);
and U8823 (N_8823,N_217,N_2973);
nand U8824 (N_8824,N_3765,N_2586);
nand U8825 (N_8825,N_3042,N_2194);
nand U8826 (N_8826,N_721,N_3440);
or U8827 (N_8827,N_1633,N_1520);
nand U8828 (N_8828,N_647,N_542);
nand U8829 (N_8829,N_664,N_3647);
nor U8830 (N_8830,N_3847,N_1466);
and U8831 (N_8831,N_4109,N_1927);
and U8832 (N_8832,N_1916,N_4132);
or U8833 (N_8833,N_3549,N_4644);
nand U8834 (N_8834,N_4151,N_2759);
nor U8835 (N_8835,N_758,N_2396);
and U8836 (N_8836,N_3258,N_2256);
and U8837 (N_8837,N_4367,N_215);
or U8838 (N_8838,N_1073,N_1060);
and U8839 (N_8839,N_2512,N_3638);
nor U8840 (N_8840,N_3702,N_3829);
and U8841 (N_8841,N_160,N_3585);
nand U8842 (N_8842,N_411,N_3239);
or U8843 (N_8843,N_139,N_1368);
nand U8844 (N_8844,N_384,N_938);
and U8845 (N_8845,N_3164,N_249);
nor U8846 (N_8846,N_1982,N_4954);
or U8847 (N_8847,N_1393,N_2148);
and U8848 (N_8848,N_2573,N_335);
and U8849 (N_8849,N_1103,N_828);
or U8850 (N_8850,N_4574,N_536);
and U8851 (N_8851,N_1319,N_4236);
and U8852 (N_8852,N_2087,N_3306);
or U8853 (N_8853,N_46,N_210);
nor U8854 (N_8854,N_4953,N_810);
or U8855 (N_8855,N_4287,N_2552);
or U8856 (N_8856,N_3093,N_600);
and U8857 (N_8857,N_2364,N_3684);
and U8858 (N_8858,N_0,N_3725);
or U8859 (N_8859,N_1411,N_2708);
nor U8860 (N_8860,N_508,N_4567);
nand U8861 (N_8861,N_1839,N_2161);
and U8862 (N_8862,N_186,N_3355);
or U8863 (N_8863,N_1014,N_2593);
nor U8864 (N_8864,N_604,N_4445);
nor U8865 (N_8865,N_1619,N_4372);
or U8866 (N_8866,N_3105,N_3730);
and U8867 (N_8867,N_692,N_3999);
nand U8868 (N_8868,N_4559,N_3276);
and U8869 (N_8869,N_806,N_4907);
or U8870 (N_8870,N_602,N_1245);
and U8871 (N_8871,N_1041,N_119);
and U8872 (N_8872,N_4164,N_792);
nor U8873 (N_8873,N_1141,N_360);
nor U8874 (N_8874,N_4163,N_2755);
and U8875 (N_8875,N_4474,N_2927);
nand U8876 (N_8876,N_4910,N_3810);
or U8877 (N_8877,N_2628,N_3050);
nand U8878 (N_8878,N_854,N_2335);
nand U8879 (N_8879,N_4431,N_4160);
nor U8880 (N_8880,N_3828,N_4423);
and U8881 (N_8881,N_3608,N_2002);
nand U8882 (N_8882,N_1761,N_2004);
and U8883 (N_8883,N_1840,N_2393);
nand U8884 (N_8884,N_1913,N_2186);
nand U8885 (N_8885,N_1374,N_1564);
nand U8886 (N_8886,N_4129,N_1481);
nand U8887 (N_8887,N_2133,N_3047);
nand U8888 (N_8888,N_1601,N_1550);
and U8889 (N_8889,N_1782,N_4970);
and U8890 (N_8890,N_288,N_2988);
nor U8891 (N_8891,N_1708,N_4206);
and U8892 (N_8892,N_3640,N_2642);
and U8893 (N_8893,N_1018,N_4251);
or U8894 (N_8894,N_4410,N_1258);
nand U8895 (N_8895,N_3497,N_824);
nor U8896 (N_8896,N_4927,N_1623);
and U8897 (N_8897,N_4597,N_1060);
nand U8898 (N_8898,N_3774,N_2755);
nor U8899 (N_8899,N_4790,N_2856);
nand U8900 (N_8900,N_4528,N_4870);
and U8901 (N_8901,N_1079,N_3697);
and U8902 (N_8902,N_3673,N_1545);
or U8903 (N_8903,N_2021,N_4611);
and U8904 (N_8904,N_290,N_3752);
and U8905 (N_8905,N_4167,N_986);
nand U8906 (N_8906,N_1608,N_4563);
and U8907 (N_8907,N_3460,N_1065);
nand U8908 (N_8908,N_942,N_2244);
and U8909 (N_8909,N_757,N_2799);
nand U8910 (N_8910,N_702,N_1209);
nor U8911 (N_8911,N_3064,N_4575);
nand U8912 (N_8912,N_1414,N_4117);
and U8913 (N_8913,N_1450,N_4452);
and U8914 (N_8914,N_4372,N_4396);
nor U8915 (N_8915,N_22,N_3360);
and U8916 (N_8916,N_660,N_1167);
nand U8917 (N_8917,N_329,N_3561);
or U8918 (N_8918,N_2233,N_774);
or U8919 (N_8919,N_4621,N_1991);
nand U8920 (N_8920,N_4650,N_3868);
or U8921 (N_8921,N_2338,N_3447);
and U8922 (N_8922,N_82,N_72);
and U8923 (N_8923,N_2478,N_991);
nand U8924 (N_8924,N_3403,N_424);
nor U8925 (N_8925,N_4353,N_3936);
nand U8926 (N_8926,N_4359,N_4740);
nor U8927 (N_8927,N_3067,N_2055);
or U8928 (N_8928,N_4544,N_3637);
nor U8929 (N_8929,N_2815,N_4581);
and U8930 (N_8930,N_2205,N_3192);
and U8931 (N_8931,N_815,N_2883);
xor U8932 (N_8932,N_2115,N_4848);
nor U8933 (N_8933,N_1856,N_1871);
nand U8934 (N_8934,N_745,N_2975);
nor U8935 (N_8935,N_4563,N_3689);
or U8936 (N_8936,N_4459,N_3165);
and U8937 (N_8937,N_392,N_958);
nand U8938 (N_8938,N_454,N_3401);
nand U8939 (N_8939,N_3616,N_4899);
or U8940 (N_8940,N_4083,N_196);
nor U8941 (N_8941,N_1250,N_3055);
or U8942 (N_8942,N_2549,N_3480);
nor U8943 (N_8943,N_3093,N_2268);
nand U8944 (N_8944,N_2062,N_3934);
nand U8945 (N_8945,N_1360,N_3390);
and U8946 (N_8946,N_3869,N_2448);
nor U8947 (N_8947,N_1370,N_955);
and U8948 (N_8948,N_2245,N_629);
and U8949 (N_8949,N_3677,N_1948);
or U8950 (N_8950,N_286,N_182);
nand U8951 (N_8951,N_4493,N_1203);
or U8952 (N_8952,N_3736,N_2595);
and U8953 (N_8953,N_3490,N_1298);
nor U8954 (N_8954,N_2851,N_1303);
or U8955 (N_8955,N_1068,N_3217);
xnor U8956 (N_8956,N_4062,N_3260);
and U8957 (N_8957,N_3237,N_3162);
and U8958 (N_8958,N_2885,N_2366);
and U8959 (N_8959,N_2265,N_3533);
nand U8960 (N_8960,N_2488,N_1243);
nor U8961 (N_8961,N_4561,N_2305);
nand U8962 (N_8962,N_4804,N_1777);
nor U8963 (N_8963,N_839,N_987);
nand U8964 (N_8964,N_3927,N_3356);
nor U8965 (N_8965,N_4341,N_3974);
nor U8966 (N_8966,N_3817,N_3161);
nand U8967 (N_8967,N_3118,N_750);
and U8968 (N_8968,N_2056,N_3826);
and U8969 (N_8969,N_2055,N_2169);
or U8970 (N_8970,N_4814,N_549);
and U8971 (N_8971,N_3893,N_4868);
and U8972 (N_8972,N_3099,N_1130);
nand U8973 (N_8973,N_370,N_4643);
nand U8974 (N_8974,N_1311,N_3392);
and U8975 (N_8975,N_2998,N_653);
and U8976 (N_8976,N_3653,N_4333);
or U8977 (N_8977,N_1203,N_3805);
xor U8978 (N_8978,N_3094,N_446);
nand U8979 (N_8979,N_1583,N_3056);
nand U8980 (N_8980,N_3518,N_4120);
nand U8981 (N_8981,N_1653,N_1767);
nor U8982 (N_8982,N_2594,N_4875);
or U8983 (N_8983,N_3620,N_2202);
and U8984 (N_8984,N_3983,N_651);
or U8985 (N_8985,N_4273,N_1022);
or U8986 (N_8986,N_1388,N_4621);
nand U8987 (N_8987,N_136,N_4972);
nor U8988 (N_8988,N_3557,N_3019);
nand U8989 (N_8989,N_2653,N_3089);
or U8990 (N_8990,N_385,N_1401);
or U8991 (N_8991,N_407,N_3261);
and U8992 (N_8992,N_4467,N_2812);
nor U8993 (N_8993,N_3099,N_2025);
nor U8994 (N_8994,N_4089,N_918);
or U8995 (N_8995,N_2950,N_3532);
nor U8996 (N_8996,N_3040,N_941);
and U8997 (N_8997,N_4983,N_3816);
and U8998 (N_8998,N_310,N_2661);
nor U8999 (N_8999,N_2313,N_2060);
or U9000 (N_9000,N_3775,N_179);
nand U9001 (N_9001,N_3639,N_3903);
and U9002 (N_9002,N_3996,N_230);
nor U9003 (N_9003,N_2534,N_2209);
and U9004 (N_9004,N_2396,N_4490);
and U9005 (N_9005,N_265,N_4738);
and U9006 (N_9006,N_870,N_2197);
and U9007 (N_9007,N_3381,N_818);
and U9008 (N_9008,N_1276,N_4629);
or U9009 (N_9009,N_4577,N_1041);
or U9010 (N_9010,N_2276,N_4787);
and U9011 (N_9011,N_1073,N_341);
and U9012 (N_9012,N_4418,N_4369);
or U9013 (N_9013,N_615,N_2457);
nand U9014 (N_9014,N_132,N_4663);
and U9015 (N_9015,N_4377,N_1037);
nor U9016 (N_9016,N_1580,N_4022);
or U9017 (N_9017,N_3894,N_1154);
or U9018 (N_9018,N_52,N_1428);
and U9019 (N_9019,N_2711,N_4839);
nor U9020 (N_9020,N_4697,N_2376);
and U9021 (N_9021,N_4751,N_3512);
and U9022 (N_9022,N_2681,N_4313);
or U9023 (N_9023,N_383,N_229);
and U9024 (N_9024,N_17,N_4190);
and U9025 (N_9025,N_2580,N_3162);
or U9026 (N_9026,N_2873,N_1424);
nand U9027 (N_9027,N_646,N_4054);
or U9028 (N_9028,N_3151,N_3323);
or U9029 (N_9029,N_471,N_3029);
nand U9030 (N_9030,N_2443,N_1196);
xor U9031 (N_9031,N_1764,N_3443);
and U9032 (N_9032,N_1426,N_2672);
nand U9033 (N_9033,N_1143,N_765);
nor U9034 (N_9034,N_4492,N_4445);
nor U9035 (N_9035,N_2911,N_531);
or U9036 (N_9036,N_698,N_1055);
nand U9037 (N_9037,N_65,N_1210);
nand U9038 (N_9038,N_293,N_633);
nand U9039 (N_9039,N_3411,N_2724);
and U9040 (N_9040,N_4880,N_1330);
or U9041 (N_9041,N_4443,N_4875);
and U9042 (N_9042,N_648,N_2260);
and U9043 (N_9043,N_309,N_952);
and U9044 (N_9044,N_2146,N_2011);
nor U9045 (N_9045,N_117,N_155);
and U9046 (N_9046,N_4212,N_1086);
nor U9047 (N_9047,N_2133,N_4895);
nor U9048 (N_9048,N_1659,N_640);
xnor U9049 (N_9049,N_3526,N_3625);
and U9050 (N_9050,N_4240,N_677);
nand U9051 (N_9051,N_974,N_284);
or U9052 (N_9052,N_4124,N_987);
nor U9053 (N_9053,N_569,N_118);
nor U9054 (N_9054,N_252,N_4266);
and U9055 (N_9055,N_3838,N_4955);
nor U9056 (N_9056,N_2664,N_1962);
nor U9057 (N_9057,N_2585,N_572);
and U9058 (N_9058,N_67,N_1222);
nor U9059 (N_9059,N_887,N_75);
and U9060 (N_9060,N_4671,N_4185);
or U9061 (N_9061,N_2012,N_4176);
or U9062 (N_9062,N_4123,N_207);
nor U9063 (N_9063,N_1241,N_4932);
nor U9064 (N_9064,N_3177,N_4306);
nor U9065 (N_9065,N_2671,N_3882);
and U9066 (N_9066,N_2911,N_4586);
and U9067 (N_9067,N_2121,N_2267);
nand U9068 (N_9068,N_1333,N_792);
and U9069 (N_9069,N_1541,N_488);
nor U9070 (N_9070,N_2440,N_4767);
or U9071 (N_9071,N_3590,N_1696);
nor U9072 (N_9072,N_3824,N_2615);
or U9073 (N_9073,N_3889,N_4145);
or U9074 (N_9074,N_1989,N_1037);
and U9075 (N_9075,N_3305,N_3703);
nand U9076 (N_9076,N_4345,N_3203);
and U9077 (N_9077,N_2762,N_2299);
nor U9078 (N_9078,N_384,N_2681);
and U9079 (N_9079,N_295,N_345);
nand U9080 (N_9080,N_4217,N_4194);
nand U9081 (N_9081,N_1485,N_1457);
and U9082 (N_9082,N_2739,N_3478);
and U9083 (N_9083,N_3725,N_2776);
nand U9084 (N_9084,N_641,N_1970);
or U9085 (N_9085,N_4877,N_976);
and U9086 (N_9086,N_3468,N_2365);
nand U9087 (N_9087,N_3802,N_1192);
nand U9088 (N_9088,N_2115,N_4156);
nand U9089 (N_9089,N_233,N_1444);
and U9090 (N_9090,N_3071,N_4162);
or U9091 (N_9091,N_4737,N_2444);
and U9092 (N_9092,N_2831,N_3);
or U9093 (N_9093,N_1589,N_3680);
and U9094 (N_9094,N_379,N_4027);
or U9095 (N_9095,N_2303,N_2842);
nand U9096 (N_9096,N_2756,N_3108);
or U9097 (N_9097,N_4946,N_2055);
nand U9098 (N_9098,N_612,N_3451);
and U9099 (N_9099,N_875,N_2668);
nor U9100 (N_9100,N_866,N_4253);
or U9101 (N_9101,N_29,N_1974);
and U9102 (N_9102,N_2426,N_4029);
nor U9103 (N_9103,N_3172,N_1825);
and U9104 (N_9104,N_3947,N_1191);
or U9105 (N_9105,N_1381,N_2);
and U9106 (N_9106,N_4106,N_372);
or U9107 (N_9107,N_4025,N_1647);
and U9108 (N_9108,N_1058,N_3971);
nor U9109 (N_9109,N_3002,N_717);
nand U9110 (N_9110,N_4181,N_5);
nor U9111 (N_9111,N_841,N_283);
nand U9112 (N_9112,N_610,N_3663);
or U9113 (N_9113,N_2737,N_4354);
nand U9114 (N_9114,N_2966,N_2123);
nor U9115 (N_9115,N_1638,N_3681);
or U9116 (N_9116,N_4143,N_370);
nand U9117 (N_9117,N_345,N_1175);
and U9118 (N_9118,N_995,N_380);
nand U9119 (N_9119,N_4812,N_1090);
nor U9120 (N_9120,N_2499,N_2355);
nand U9121 (N_9121,N_1962,N_2003);
nor U9122 (N_9122,N_1928,N_2709);
or U9123 (N_9123,N_417,N_1642);
nor U9124 (N_9124,N_2745,N_2845);
or U9125 (N_9125,N_1869,N_1526);
nor U9126 (N_9126,N_2608,N_2037);
nor U9127 (N_9127,N_2388,N_3686);
nand U9128 (N_9128,N_2344,N_4881);
or U9129 (N_9129,N_4653,N_1059);
or U9130 (N_9130,N_1477,N_1918);
xnor U9131 (N_9131,N_2943,N_1648);
nor U9132 (N_9132,N_1287,N_1581);
nor U9133 (N_9133,N_3637,N_4765);
or U9134 (N_9134,N_600,N_3675);
and U9135 (N_9135,N_1165,N_1044);
nand U9136 (N_9136,N_4893,N_2794);
and U9137 (N_9137,N_709,N_4107);
or U9138 (N_9138,N_1182,N_4527);
and U9139 (N_9139,N_3195,N_4591);
nor U9140 (N_9140,N_2940,N_2711);
or U9141 (N_9141,N_4004,N_2006);
nand U9142 (N_9142,N_4821,N_4073);
xor U9143 (N_9143,N_1278,N_2353);
nor U9144 (N_9144,N_2194,N_353);
and U9145 (N_9145,N_4641,N_1378);
or U9146 (N_9146,N_1662,N_4826);
and U9147 (N_9147,N_1883,N_2779);
nor U9148 (N_9148,N_2534,N_3292);
and U9149 (N_9149,N_4899,N_3200);
nand U9150 (N_9150,N_392,N_1076);
or U9151 (N_9151,N_668,N_4028);
nand U9152 (N_9152,N_1022,N_2580);
and U9153 (N_9153,N_722,N_515);
and U9154 (N_9154,N_4946,N_3918);
or U9155 (N_9155,N_303,N_1319);
and U9156 (N_9156,N_2845,N_4917);
or U9157 (N_9157,N_524,N_2334);
nand U9158 (N_9158,N_4755,N_851);
nor U9159 (N_9159,N_4826,N_3824);
or U9160 (N_9160,N_4497,N_2831);
and U9161 (N_9161,N_2573,N_341);
xor U9162 (N_9162,N_2489,N_2018);
nor U9163 (N_9163,N_2935,N_4034);
nor U9164 (N_9164,N_3649,N_3981);
or U9165 (N_9165,N_3845,N_101);
nor U9166 (N_9166,N_1374,N_2016);
or U9167 (N_9167,N_3743,N_2665);
nand U9168 (N_9168,N_1454,N_2996);
or U9169 (N_9169,N_2715,N_1201);
and U9170 (N_9170,N_3983,N_3404);
or U9171 (N_9171,N_187,N_1788);
and U9172 (N_9172,N_3425,N_2861);
nand U9173 (N_9173,N_2469,N_1540);
nor U9174 (N_9174,N_2664,N_768);
and U9175 (N_9175,N_4386,N_4219);
or U9176 (N_9176,N_4033,N_2884);
or U9177 (N_9177,N_2041,N_3025);
nor U9178 (N_9178,N_2936,N_3314);
or U9179 (N_9179,N_2583,N_2142);
nand U9180 (N_9180,N_1736,N_3868);
and U9181 (N_9181,N_1470,N_3609);
nand U9182 (N_9182,N_911,N_1103);
nor U9183 (N_9183,N_3149,N_4001);
and U9184 (N_9184,N_352,N_2492);
or U9185 (N_9185,N_1594,N_1138);
and U9186 (N_9186,N_1675,N_4203);
nor U9187 (N_9187,N_1396,N_2080);
or U9188 (N_9188,N_1695,N_582);
and U9189 (N_9189,N_2804,N_641);
or U9190 (N_9190,N_4196,N_4017);
or U9191 (N_9191,N_1780,N_4599);
and U9192 (N_9192,N_4220,N_2024);
and U9193 (N_9193,N_4810,N_3261);
or U9194 (N_9194,N_3059,N_1604);
and U9195 (N_9195,N_4843,N_1246);
or U9196 (N_9196,N_1243,N_2855);
and U9197 (N_9197,N_1989,N_1739);
nor U9198 (N_9198,N_3142,N_3878);
or U9199 (N_9199,N_3574,N_82);
nand U9200 (N_9200,N_45,N_408);
or U9201 (N_9201,N_3648,N_4801);
nor U9202 (N_9202,N_31,N_4929);
nor U9203 (N_9203,N_4736,N_4778);
nor U9204 (N_9204,N_2799,N_1494);
or U9205 (N_9205,N_897,N_4936);
nand U9206 (N_9206,N_4189,N_4085);
or U9207 (N_9207,N_1020,N_4424);
nand U9208 (N_9208,N_4399,N_4427);
nand U9209 (N_9209,N_2277,N_4559);
nand U9210 (N_9210,N_1926,N_4524);
or U9211 (N_9211,N_1057,N_671);
nand U9212 (N_9212,N_251,N_953);
and U9213 (N_9213,N_1183,N_1574);
xor U9214 (N_9214,N_4531,N_4468);
nand U9215 (N_9215,N_594,N_29);
nand U9216 (N_9216,N_533,N_2690);
nand U9217 (N_9217,N_2299,N_4571);
nand U9218 (N_9218,N_3692,N_1026);
or U9219 (N_9219,N_2124,N_1912);
nand U9220 (N_9220,N_3048,N_2371);
nand U9221 (N_9221,N_586,N_22);
nand U9222 (N_9222,N_4851,N_3494);
nor U9223 (N_9223,N_1856,N_4426);
nand U9224 (N_9224,N_202,N_1297);
nand U9225 (N_9225,N_1166,N_1208);
nand U9226 (N_9226,N_617,N_4531);
or U9227 (N_9227,N_3256,N_1042);
or U9228 (N_9228,N_1247,N_2779);
nor U9229 (N_9229,N_2844,N_2848);
nand U9230 (N_9230,N_154,N_3229);
or U9231 (N_9231,N_271,N_630);
nand U9232 (N_9232,N_3561,N_3953);
or U9233 (N_9233,N_671,N_3114);
or U9234 (N_9234,N_3011,N_4916);
and U9235 (N_9235,N_517,N_3402);
or U9236 (N_9236,N_1529,N_744);
and U9237 (N_9237,N_3652,N_2008);
nand U9238 (N_9238,N_283,N_3494);
nand U9239 (N_9239,N_4400,N_3187);
nor U9240 (N_9240,N_792,N_2759);
or U9241 (N_9241,N_578,N_3896);
xnor U9242 (N_9242,N_4426,N_1239);
nand U9243 (N_9243,N_2972,N_4602);
nor U9244 (N_9244,N_2889,N_4305);
or U9245 (N_9245,N_1157,N_2452);
and U9246 (N_9246,N_559,N_194);
nor U9247 (N_9247,N_2382,N_1707);
nor U9248 (N_9248,N_949,N_2800);
nand U9249 (N_9249,N_2985,N_1813);
nor U9250 (N_9250,N_1216,N_1508);
or U9251 (N_9251,N_88,N_1296);
nand U9252 (N_9252,N_1022,N_2503);
or U9253 (N_9253,N_4389,N_2584);
and U9254 (N_9254,N_2490,N_3740);
nand U9255 (N_9255,N_471,N_1636);
and U9256 (N_9256,N_2258,N_4713);
nor U9257 (N_9257,N_1430,N_2340);
nor U9258 (N_9258,N_2040,N_2446);
or U9259 (N_9259,N_3983,N_4511);
nand U9260 (N_9260,N_948,N_935);
nand U9261 (N_9261,N_4473,N_2663);
or U9262 (N_9262,N_2600,N_4696);
nand U9263 (N_9263,N_4424,N_312);
or U9264 (N_9264,N_1464,N_2494);
and U9265 (N_9265,N_4601,N_245);
nor U9266 (N_9266,N_3313,N_4341);
and U9267 (N_9267,N_4286,N_3702);
or U9268 (N_9268,N_1081,N_4260);
or U9269 (N_9269,N_4577,N_1458);
nor U9270 (N_9270,N_2813,N_4090);
nand U9271 (N_9271,N_3173,N_1584);
and U9272 (N_9272,N_4515,N_496);
and U9273 (N_9273,N_815,N_4885);
nand U9274 (N_9274,N_145,N_3298);
nor U9275 (N_9275,N_2257,N_325);
nand U9276 (N_9276,N_3746,N_4748);
or U9277 (N_9277,N_3987,N_4921);
and U9278 (N_9278,N_1111,N_1070);
or U9279 (N_9279,N_332,N_1107);
and U9280 (N_9280,N_898,N_578);
and U9281 (N_9281,N_1174,N_3871);
nor U9282 (N_9282,N_45,N_1913);
nor U9283 (N_9283,N_2234,N_1174);
nor U9284 (N_9284,N_2521,N_449);
nor U9285 (N_9285,N_1405,N_616);
nor U9286 (N_9286,N_2844,N_2042);
nor U9287 (N_9287,N_4901,N_2789);
nand U9288 (N_9288,N_3898,N_3692);
or U9289 (N_9289,N_831,N_3689);
nor U9290 (N_9290,N_574,N_1881);
or U9291 (N_9291,N_4450,N_4999);
or U9292 (N_9292,N_3518,N_864);
nand U9293 (N_9293,N_499,N_4962);
and U9294 (N_9294,N_2354,N_2268);
nor U9295 (N_9295,N_2508,N_3018);
or U9296 (N_9296,N_4920,N_3903);
or U9297 (N_9297,N_3909,N_2978);
nor U9298 (N_9298,N_677,N_1350);
or U9299 (N_9299,N_1112,N_2408);
and U9300 (N_9300,N_4144,N_3662);
nand U9301 (N_9301,N_4607,N_4323);
and U9302 (N_9302,N_2992,N_4527);
or U9303 (N_9303,N_129,N_3908);
or U9304 (N_9304,N_4878,N_2624);
nand U9305 (N_9305,N_3601,N_4056);
or U9306 (N_9306,N_3766,N_3669);
nor U9307 (N_9307,N_3757,N_3849);
nor U9308 (N_9308,N_2919,N_4703);
nor U9309 (N_9309,N_3685,N_580);
xor U9310 (N_9310,N_1933,N_3782);
and U9311 (N_9311,N_1298,N_1788);
and U9312 (N_9312,N_1036,N_4152);
nor U9313 (N_9313,N_4258,N_2571);
and U9314 (N_9314,N_3988,N_2895);
and U9315 (N_9315,N_1311,N_4126);
or U9316 (N_9316,N_3427,N_22);
nand U9317 (N_9317,N_4118,N_2951);
or U9318 (N_9318,N_2669,N_403);
nand U9319 (N_9319,N_2326,N_1682);
nor U9320 (N_9320,N_3468,N_1293);
nand U9321 (N_9321,N_539,N_3397);
nand U9322 (N_9322,N_2273,N_4121);
and U9323 (N_9323,N_148,N_3053);
nand U9324 (N_9324,N_1904,N_1821);
nand U9325 (N_9325,N_2278,N_3188);
nor U9326 (N_9326,N_4953,N_3018);
or U9327 (N_9327,N_4792,N_1467);
nor U9328 (N_9328,N_3654,N_4024);
nand U9329 (N_9329,N_3938,N_951);
and U9330 (N_9330,N_4189,N_3340);
or U9331 (N_9331,N_2324,N_2585);
or U9332 (N_9332,N_770,N_2615);
and U9333 (N_9333,N_2862,N_1460);
nor U9334 (N_9334,N_1886,N_656);
or U9335 (N_9335,N_4027,N_4711);
and U9336 (N_9336,N_2578,N_4845);
nand U9337 (N_9337,N_2176,N_2162);
or U9338 (N_9338,N_3022,N_3946);
nor U9339 (N_9339,N_4892,N_2576);
nor U9340 (N_9340,N_4461,N_4663);
and U9341 (N_9341,N_2818,N_2507);
and U9342 (N_9342,N_919,N_4432);
and U9343 (N_9343,N_2295,N_4918);
and U9344 (N_9344,N_2097,N_2426);
xor U9345 (N_9345,N_2648,N_2850);
or U9346 (N_9346,N_2000,N_924);
nor U9347 (N_9347,N_3541,N_1010);
nor U9348 (N_9348,N_4045,N_3006);
nand U9349 (N_9349,N_3539,N_3680);
nand U9350 (N_9350,N_1130,N_1323);
or U9351 (N_9351,N_2417,N_3870);
nand U9352 (N_9352,N_4318,N_3590);
and U9353 (N_9353,N_3637,N_868);
nor U9354 (N_9354,N_4214,N_3019);
nor U9355 (N_9355,N_3318,N_4176);
nor U9356 (N_9356,N_2018,N_81);
nand U9357 (N_9357,N_1454,N_3119);
or U9358 (N_9358,N_1539,N_280);
or U9359 (N_9359,N_2615,N_739);
or U9360 (N_9360,N_4376,N_3320);
nor U9361 (N_9361,N_2621,N_1743);
or U9362 (N_9362,N_2620,N_1686);
or U9363 (N_9363,N_1084,N_2023);
and U9364 (N_9364,N_4733,N_4172);
nand U9365 (N_9365,N_1688,N_96);
nand U9366 (N_9366,N_1834,N_3988);
or U9367 (N_9367,N_1267,N_844);
and U9368 (N_9368,N_2564,N_39);
and U9369 (N_9369,N_4409,N_2093);
or U9370 (N_9370,N_1902,N_2134);
nor U9371 (N_9371,N_2919,N_3689);
nor U9372 (N_9372,N_3250,N_3619);
or U9373 (N_9373,N_2049,N_3146);
nand U9374 (N_9374,N_463,N_2343);
or U9375 (N_9375,N_4801,N_2968);
nor U9376 (N_9376,N_1846,N_3983);
or U9377 (N_9377,N_3167,N_4802);
or U9378 (N_9378,N_373,N_4786);
nand U9379 (N_9379,N_1998,N_4432);
or U9380 (N_9380,N_3332,N_3562);
or U9381 (N_9381,N_498,N_4261);
nor U9382 (N_9382,N_1131,N_921);
nor U9383 (N_9383,N_1517,N_45);
nand U9384 (N_9384,N_355,N_650);
nand U9385 (N_9385,N_1568,N_462);
or U9386 (N_9386,N_4717,N_3158);
nor U9387 (N_9387,N_1842,N_2958);
nor U9388 (N_9388,N_2823,N_1070);
nor U9389 (N_9389,N_4878,N_241);
or U9390 (N_9390,N_2185,N_4791);
and U9391 (N_9391,N_1117,N_1650);
or U9392 (N_9392,N_754,N_566);
or U9393 (N_9393,N_2989,N_3793);
or U9394 (N_9394,N_1588,N_4507);
or U9395 (N_9395,N_2183,N_117);
xor U9396 (N_9396,N_2510,N_4538);
and U9397 (N_9397,N_2370,N_4419);
and U9398 (N_9398,N_1157,N_4057);
and U9399 (N_9399,N_1105,N_4153);
and U9400 (N_9400,N_3648,N_3924);
and U9401 (N_9401,N_2692,N_1093);
and U9402 (N_9402,N_3041,N_601);
nand U9403 (N_9403,N_878,N_215);
nor U9404 (N_9404,N_2137,N_1121);
and U9405 (N_9405,N_736,N_3019);
or U9406 (N_9406,N_371,N_3982);
nand U9407 (N_9407,N_3997,N_1831);
and U9408 (N_9408,N_552,N_4560);
nand U9409 (N_9409,N_3946,N_2313);
nand U9410 (N_9410,N_3917,N_1025);
nor U9411 (N_9411,N_4052,N_4999);
nand U9412 (N_9412,N_202,N_388);
or U9413 (N_9413,N_435,N_2658);
or U9414 (N_9414,N_535,N_3543);
nor U9415 (N_9415,N_3046,N_3031);
nand U9416 (N_9416,N_2224,N_168);
xnor U9417 (N_9417,N_1520,N_479);
and U9418 (N_9418,N_3542,N_2071);
nor U9419 (N_9419,N_1372,N_1375);
and U9420 (N_9420,N_4999,N_2957);
and U9421 (N_9421,N_3058,N_1581);
and U9422 (N_9422,N_890,N_2733);
and U9423 (N_9423,N_2387,N_4844);
or U9424 (N_9424,N_308,N_3516);
or U9425 (N_9425,N_1803,N_1533);
nor U9426 (N_9426,N_4172,N_918);
or U9427 (N_9427,N_3256,N_4846);
nand U9428 (N_9428,N_1122,N_472);
nand U9429 (N_9429,N_4009,N_1532);
nor U9430 (N_9430,N_4172,N_5);
and U9431 (N_9431,N_1217,N_3128);
nand U9432 (N_9432,N_1816,N_2861);
xnor U9433 (N_9433,N_1936,N_907);
nand U9434 (N_9434,N_948,N_1693);
and U9435 (N_9435,N_753,N_938);
nand U9436 (N_9436,N_2345,N_468);
nand U9437 (N_9437,N_1594,N_1515);
and U9438 (N_9438,N_3630,N_4449);
nor U9439 (N_9439,N_3236,N_3483);
nor U9440 (N_9440,N_1320,N_4472);
nor U9441 (N_9441,N_120,N_743);
or U9442 (N_9442,N_2929,N_1369);
nor U9443 (N_9443,N_2194,N_1382);
or U9444 (N_9444,N_3850,N_2732);
or U9445 (N_9445,N_3916,N_102);
nor U9446 (N_9446,N_1416,N_1299);
nor U9447 (N_9447,N_2597,N_819);
or U9448 (N_9448,N_2268,N_3630);
nand U9449 (N_9449,N_1896,N_1284);
and U9450 (N_9450,N_4401,N_633);
and U9451 (N_9451,N_3168,N_1447);
or U9452 (N_9452,N_2981,N_171);
or U9453 (N_9453,N_1512,N_1965);
nor U9454 (N_9454,N_1405,N_3180);
nor U9455 (N_9455,N_1285,N_3677);
nand U9456 (N_9456,N_1777,N_4075);
nand U9457 (N_9457,N_4187,N_1487);
nor U9458 (N_9458,N_4525,N_3024);
nor U9459 (N_9459,N_4635,N_3471);
or U9460 (N_9460,N_1782,N_2008);
or U9461 (N_9461,N_4030,N_1824);
and U9462 (N_9462,N_1243,N_2287);
nor U9463 (N_9463,N_197,N_4630);
nand U9464 (N_9464,N_2864,N_1489);
and U9465 (N_9465,N_4158,N_98);
or U9466 (N_9466,N_4801,N_904);
or U9467 (N_9467,N_390,N_3174);
nor U9468 (N_9468,N_2176,N_325);
and U9469 (N_9469,N_3946,N_3966);
or U9470 (N_9470,N_3881,N_1838);
nor U9471 (N_9471,N_2288,N_388);
and U9472 (N_9472,N_2732,N_4293);
nand U9473 (N_9473,N_3136,N_1817);
nand U9474 (N_9474,N_1655,N_3435);
nor U9475 (N_9475,N_3115,N_3866);
and U9476 (N_9476,N_301,N_1241);
or U9477 (N_9477,N_3243,N_4233);
or U9478 (N_9478,N_3231,N_4832);
and U9479 (N_9479,N_1763,N_3567);
and U9480 (N_9480,N_34,N_4682);
or U9481 (N_9481,N_3717,N_1956);
or U9482 (N_9482,N_1096,N_4458);
or U9483 (N_9483,N_4892,N_3370);
or U9484 (N_9484,N_3431,N_1554);
nor U9485 (N_9485,N_1153,N_3718);
nor U9486 (N_9486,N_1801,N_1626);
and U9487 (N_9487,N_1068,N_886);
or U9488 (N_9488,N_581,N_243);
nor U9489 (N_9489,N_4716,N_699);
and U9490 (N_9490,N_2508,N_246);
or U9491 (N_9491,N_1690,N_1191);
or U9492 (N_9492,N_601,N_1348);
nand U9493 (N_9493,N_2187,N_2638);
and U9494 (N_9494,N_3849,N_387);
nor U9495 (N_9495,N_1778,N_1312);
and U9496 (N_9496,N_2894,N_1023);
or U9497 (N_9497,N_1640,N_1424);
or U9498 (N_9498,N_1505,N_2797);
nor U9499 (N_9499,N_2631,N_4366);
nand U9500 (N_9500,N_2240,N_2093);
nor U9501 (N_9501,N_4681,N_223);
nand U9502 (N_9502,N_1472,N_2023);
nand U9503 (N_9503,N_4090,N_3349);
and U9504 (N_9504,N_2840,N_2744);
nor U9505 (N_9505,N_1919,N_748);
nor U9506 (N_9506,N_4616,N_1609);
xor U9507 (N_9507,N_2654,N_3294);
and U9508 (N_9508,N_4803,N_866);
nand U9509 (N_9509,N_3147,N_3844);
or U9510 (N_9510,N_2844,N_255);
nor U9511 (N_9511,N_2094,N_2265);
or U9512 (N_9512,N_2132,N_3602);
nor U9513 (N_9513,N_1159,N_4829);
nor U9514 (N_9514,N_3347,N_3931);
and U9515 (N_9515,N_2057,N_4461);
or U9516 (N_9516,N_387,N_3237);
or U9517 (N_9517,N_268,N_567);
nor U9518 (N_9518,N_500,N_1687);
and U9519 (N_9519,N_1288,N_4685);
nor U9520 (N_9520,N_2192,N_1115);
nor U9521 (N_9521,N_2687,N_876);
and U9522 (N_9522,N_4541,N_2524);
or U9523 (N_9523,N_2522,N_1328);
nand U9524 (N_9524,N_1076,N_549);
nand U9525 (N_9525,N_2704,N_4565);
xor U9526 (N_9526,N_3578,N_4402);
nand U9527 (N_9527,N_196,N_3800);
nand U9528 (N_9528,N_3934,N_2371);
and U9529 (N_9529,N_584,N_3172);
or U9530 (N_9530,N_4071,N_3926);
nand U9531 (N_9531,N_4405,N_1281);
and U9532 (N_9532,N_3779,N_4881);
nor U9533 (N_9533,N_999,N_4789);
or U9534 (N_9534,N_3859,N_4056);
nand U9535 (N_9535,N_4621,N_4942);
nor U9536 (N_9536,N_985,N_2868);
or U9537 (N_9537,N_3863,N_3325);
nand U9538 (N_9538,N_159,N_2862);
nand U9539 (N_9539,N_478,N_306);
and U9540 (N_9540,N_4488,N_1523);
or U9541 (N_9541,N_1882,N_524);
nor U9542 (N_9542,N_714,N_2108);
nand U9543 (N_9543,N_1046,N_2545);
nor U9544 (N_9544,N_4247,N_2636);
and U9545 (N_9545,N_3041,N_274);
nand U9546 (N_9546,N_3413,N_476);
nand U9547 (N_9547,N_3580,N_4565);
and U9548 (N_9548,N_167,N_4373);
nand U9549 (N_9549,N_1014,N_76);
and U9550 (N_9550,N_3409,N_3576);
or U9551 (N_9551,N_4236,N_188);
nand U9552 (N_9552,N_3652,N_4172);
or U9553 (N_9553,N_3687,N_4735);
and U9554 (N_9554,N_3687,N_3476);
nand U9555 (N_9555,N_2169,N_1571);
or U9556 (N_9556,N_3069,N_1682);
and U9557 (N_9557,N_2451,N_3201);
and U9558 (N_9558,N_308,N_2372);
nand U9559 (N_9559,N_3291,N_767);
and U9560 (N_9560,N_3,N_1016);
nor U9561 (N_9561,N_647,N_2581);
nor U9562 (N_9562,N_4917,N_3387);
nor U9563 (N_9563,N_2586,N_3036);
and U9564 (N_9564,N_1690,N_1818);
and U9565 (N_9565,N_1257,N_1953);
nor U9566 (N_9566,N_117,N_564);
or U9567 (N_9567,N_3342,N_354);
and U9568 (N_9568,N_539,N_1400);
nand U9569 (N_9569,N_2010,N_228);
and U9570 (N_9570,N_3383,N_4033);
nor U9571 (N_9571,N_1436,N_1363);
and U9572 (N_9572,N_3903,N_3362);
and U9573 (N_9573,N_4743,N_340);
nor U9574 (N_9574,N_2147,N_19);
nand U9575 (N_9575,N_882,N_4017);
or U9576 (N_9576,N_3773,N_623);
and U9577 (N_9577,N_3666,N_3921);
nand U9578 (N_9578,N_3277,N_1151);
nor U9579 (N_9579,N_1670,N_4930);
or U9580 (N_9580,N_3944,N_33);
and U9581 (N_9581,N_202,N_2754);
nor U9582 (N_9582,N_319,N_2927);
and U9583 (N_9583,N_4803,N_1043);
nor U9584 (N_9584,N_695,N_4367);
or U9585 (N_9585,N_4023,N_1007);
nor U9586 (N_9586,N_2671,N_2787);
nand U9587 (N_9587,N_904,N_2869);
nor U9588 (N_9588,N_2362,N_4944);
and U9589 (N_9589,N_4520,N_54);
and U9590 (N_9590,N_4929,N_436);
or U9591 (N_9591,N_2576,N_233);
or U9592 (N_9592,N_4357,N_315);
nand U9593 (N_9593,N_4589,N_1936);
or U9594 (N_9594,N_4721,N_3626);
or U9595 (N_9595,N_2468,N_2311);
nand U9596 (N_9596,N_1844,N_1534);
nor U9597 (N_9597,N_4951,N_1581);
or U9598 (N_9598,N_4072,N_312);
nor U9599 (N_9599,N_4206,N_3651);
or U9600 (N_9600,N_923,N_2447);
nand U9601 (N_9601,N_3290,N_1591);
nand U9602 (N_9602,N_2066,N_2411);
or U9603 (N_9603,N_2908,N_4449);
or U9604 (N_9604,N_2984,N_3149);
and U9605 (N_9605,N_170,N_728);
nand U9606 (N_9606,N_4969,N_139);
and U9607 (N_9607,N_1976,N_3760);
nor U9608 (N_9608,N_1741,N_3818);
nand U9609 (N_9609,N_4764,N_745);
nand U9610 (N_9610,N_1289,N_2101);
and U9611 (N_9611,N_2088,N_274);
nand U9612 (N_9612,N_4311,N_127);
or U9613 (N_9613,N_3843,N_770);
and U9614 (N_9614,N_4101,N_194);
or U9615 (N_9615,N_4938,N_4266);
nand U9616 (N_9616,N_4253,N_1566);
nand U9617 (N_9617,N_1047,N_3501);
and U9618 (N_9618,N_504,N_3053);
nand U9619 (N_9619,N_2054,N_277);
nor U9620 (N_9620,N_3724,N_129);
nand U9621 (N_9621,N_3887,N_1233);
nand U9622 (N_9622,N_505,N_4354);
nor U9623 (N_9623,N_2112,N_3741);
nor U9624 (N_9624,N_4620,N_804);
and U9625 (N_9625,N_4149,N_1581);
or U9626 (N_9626,N_3138,N_4155);
nand U9627 (N_9627,N_1568,N_3186);
nor U9628 (N_9628,N_3210,N_971);
nor U9629 (N_9629,N_819,N_1861);
or U9630 (N_9630,N_2715,N_1056);
or U9631 (N_9631,N_1352,N_4424);
or U9632 (N_9632,N_1518,N_2432);
nor U9633 (N_9633,N_856,N_4713);
nor U9634 (N_9634,N_3302,N_1707);
nand U9635 (N_9635,N_721,N_2985);
and U9636 (N_9636,N_249,N_257);
nor U9637 (N_9637,N_3551,N_3328);
or U9638 (N_9638,N_4486,N_2860);
or U9639 (N_9639,N_2415,N_2186);
nor U9640 (N_9640,N_2339,N_173);
nand U9641 (N_9641,N_701,N_3317);
nand U9642 (N_9642,N_172,N_1231);
nor U9643 (N_9643,N_1217,N_4687);
or U9644 (N_9644,N_1518,N_0);
or U9645 (N_9645,N_4752,N_4195);
and U9646 (N_9646,N_4518,N_4424);
or U9647 (N_9647,N_815,N_4644);
or U9648 (N_9648,N_4747,N_1851);
nand U9649 (N_9649,N_2318,N_1314);
or U9650 (N_9650,N_622,N_1106);
nand U9651 (N_9651,N_1723,N_1335);
nand U9652 (N_9652,N_1062,N_4693);
nand U9653 (N_9653,N_681,N_3482);
nor U9654 (N_9654,N_297,N_3613);
or U9655 (N_9655,N_2488,N_772);
nor U9656 (N_9656,N_1399,N_1566);
nor U9657 (N_9657,N_1414,N_720);
nor U9658 (N_9658,N_691,N_4519);
and U9659 (N_9659,N_3068,N_419);
nor U9660 (N_9660,N_3703,N_4829);
or U9661 (N_9661,N_134,N_1091);
nand U9662 (N_9662,N_504,N_1849);
and U9663 (N_9663,N_4166,N_4896);
nor U9664 (N_9664,N_1001,N_2828);
and U9665 (N_9665,N_1604,N_94);
and U9666 (N_9666,N_1708,N_3482);
nor U9667 (N_9667,N_1649,N_4003);
or U9668 (N_9668,N_674,N_2454);
and U9669 (N_9669,N_1315,N_2294);
and U9670 (N_9670,N_3048,N_65);
nand U9671 (N_9671,N_2807,N_1191);
nand U9672 (N_9672,N_3975,N_468);
and U9673 (N_9673,N_3109,N_580);
and U9674 (N_9674,N_3769,N_4835);
nor U9675 (N_9675,N_9,N_1660);
and U9676 (N_9676,N_4260,N_2933);
nand U9677 (N_9677,N_2357,N_478);
or U9678 (N_9678,N_1459,N_3772);
nand U9679 (N_9679,N_3067,N_1207);
nand U9680 (N_9680,N_2178,N_2733);
or U9681 (N_9681,N_702,N_4105);
nor U9682 (N_9682,N_2305,N_4327);
or U9683 (N_9683,N_4760,N_4706);
nor U9684 (N_9684,N_978,N_2060);
nor U9685 (N_9685,N_4701,N_3682);
or U9686 (N_9686,N_309,N_3177);
nand U9687 (N_9687,N_2798,N_1309);
nor U9688 (N_9688,N_2504,N_4930);
and U9689 (N_9689,N_1702,N_1288);
nand U9690 (N_9690,N_1912,N_4103);
nor U9691 (N_9691,N_2908,N_627);
and U9692 (N_9692,N_2991,N_240);
nand U9693 (N_9693,N_1315,N_4026);
and U9694 (N_9694,N_3220,N_652);
or U9695 (N_9695,N_859,N_4326);
nand U9696 (N_9696,N_2210,N_1380);
nand U9697 (N_9697,N_4072,N_3320);
nor U9698 (N_9698,N_3653,N_3983);
nand U9699 (N_9699,N_744,N_1392);
nand U9700 (N_9700,N_67,N_3768);
nand U9701 (N_9701,N_2943,N_2437);
or U9702 (N_9702,N_3260,N_4295);
nand U9703 (N_9703,N_4827,N_934);
nor U9704 (N_9704,N_2656,N_3420);
and U9705 (N_9705,N_275,N_2755);
nand U9706 (N_9706,N_4471,N_4226);
and U9707 (N_9707,N_1849,N_97);
or U9708 (N_9708,N_2029,N_4321);
nand U9709 (N_9709,N_1799,N_3620);
nor U9710 (N_9710,N_3304,N_1052);
and U9711 (N_9711,N_2550,N_3237);
or U9712 (N_9712,N_1154,N_2216);
nand U9713 (N_9713,N_1469,N_473);
nand U9714 (N_9714,N_4084,N_1590);
or U9715 (N_9715,N_2402,N_2613);
nand U9716 (N_9716,N_2909,N_1509);
and U9717 (N_9717,N_863,N_3251);
and U9718 (N_9718,N_4689,N_2772);
nand U9719 (N_9719,N_1761,N_3020);
nand U9720 (N_9720,N_1208,N_1266);
nor U9721 (N_9721,N_3391,N_3696);
nand U9722 (N_9722,N_2301,N_1581);
and U9723 (N_9723,N_3145,N_3496);
and U9724 (N_9724,N_4080,N_4564);
nor U9725 (N_9725,N_3544,N_3493);
or U9726 (N_9726,N_4585,N_3300);
or U9727 (N_9727,N_4338,N_1890);
or U9728 (N_9728,N_1230,N_4638);
nand U9729 (N_9729,N_2125,N_2697);
nand U9730 (N_9730,N_1579,N_3037);
and U9731 (N_9731,N_2181,N_3141);
or U9732 (N_9732,N_686,N_4164);
nand U9733 (N_9733,N_4979,N_4327);
or U9734 (N_9734,N_545,N_3696);
and U9735 (N_9735,N_4628,N_4056);
or U9736 (N_9736,N_605,N_3929);
nor U9737 (N_9737,N_1929,N_2300);
nor U9738 (N_9738,N_4922,N_425);
nor U9739 (N_9739,N_1249,N_2091);
and U9740 (N_9740,N_40,N_2802);
and U9741 (N_9741,N_969,N_1615);
nand U9742 (N_9742,N_3792,N_975);
nand U9743 (N_9743,N_2229,N_4966);
nor U9744 (N_9744,N_4559,N_4953);
nor U9745 (N_9745,N_3436,N_1957);
and U9746 (N_9746,N_3846,N_1187);
nand U9747 (N_9747,N_1523,N_1407);
nor U9748 (N_9748,N_3988,N_1595);
and U9749 (N_9749,N_1762,N_910);
nand U9750 (N_9750,N_3567,N_4070);
nor U9751 (N_9751,N_1150,N_4356);
nor U9752 (N_9752,N_1277,N_4196);
or U9753 (N_9753,N_3645,N_3707);
or U9754 (N_9754,N_3011,N_1433);
nor U9755 (N_9755,N_3658,N_4063);
nor U9756 (N_9756,N_3899,N_2990);
and U9757 (N_9757,N_2241,N_2661);
nor U9758 (N_9758,N_819,N_193);
and U9759 (N_9759,N_3891,N_1600);
or U9760 (N_9760,N_2722,N_1530);
nand U9761 (N_9761,N_2816,N_4148);
and U9762 (N_9762,N_2719,N_947);
nor U9763 (N_9763,N_4071,N_4218);
nor U9764 (N_9764,N_1179,N_390);
and U9765 (N_9765,N_3982,N_142);
nor U9766 (N_9766,N_215,N_46);
nor U9767 (N_9767,N_1751,N_4535);
or U9768 (N_9768,N_4868,N_2127);
or U9769 (N_9769,N_1210,N_1256);
and U9770 (N_9770,N_4760,N_2209);
nand U9771 (N_9771,N_158,N_4369);
or U9772 (N_9772,N_1972,N_2812);
or U9773 (N_9773,N_4091,N_2329);
nand U9774 (N_9774,N_2059,N_890);
nor U9775 (N_9775,N_386,N_4112);
and U9776 (N_9776,N_4010,N_1299);
and U9777 (N_9777,N_3676,N_3929);
nand U9778 (N_9778,N_2833,N_422);
and U9779 (N_9779,N_63,N_4716);
and U9780 (N_9780,N_1464,N_4566);
and U9781 (N_9781,N_218,N_708);
nor U9782 (N_9782,N_3049,N_3656);
nor U9783 (N_9783,N_3773,N_1262);
nor U9784 (N_9784,N_3776,N_1093);
or U9785 (N_9785,N_4431,N_4227);
nor U9786 (N_9786,N_359,N_1852);
and U9787 (N_9787,N_1577,N_4422);
and U9788 (N_9788,N_2820,N_3787);
nor U9789 (N_9789,N_2945,N_612);
nor U9790 (N_9790,N_597,N_3929);
and U9791 (N_9791,N_2849,N_2033);
nand U9792 (N_9792,N_1998,N_2332);
or U9793 (N_9793,N_2490,N_3161);
or U9794 (N_9794,N_203,N_4977);
or U9795 (N_9795,N_3570,N_2449);
nand U9796 (N_9796,N_1244,N_4564);
nor U9797 (N_9797,N_696,N_4745);
nand U9798 (N_9798,N_2860,N_78);
nand U9799 (N_9799,N_2647,N_2147);
and U9800 (N_9800,N_4948,N_2009);
and U9801 (N_9801,N_4137,N_2454);
nand U9802 (N_9802,N_1587,N_2372);
or U9803 (N_9803,N_2096,N_3045);
nor U9804 (N_9804,N_1710,N_52);
or U9805 (N_9805,N_3926,N_2216);
or U9806 (N_9806,N_4150,N_241);
or U9807 (N_9807,N_1414,N_3491);
and U9808 (N_9808,N_1555,N_3306);
nand U9809 (N_9809,N_4181,N_3904);
and U9810 (N_9810,N_3438,N_4087);
nor U9811 (N_9811,N_1816,N_4282);
and U9812 (N_9812,N_1031,N_2181);
and U9813 (N_9813,N_3965,N_40);
nor U9814 (N_9814,N_675,N_2865);
nor U9815 (N_9815,N_1413,N_4192);
or U9816 (N_9816,N_874,N_690);
nand U9817 (N_9817,N_933,N_1294);
nor U9818 (N_9818,N_483,N_1840);
nand U9819 (N_9819,N_1184,N_1141);
xor U9820 (N_9820,N_1227,N_4541);
and U9821 (N_9821,N_1223,N_170);
nand U9822 (N_9822,N_1013,N_3621);
and U9823 (N_9823,N_2878,N_4714);
and U9824 (N_9824,N_4081,N_2612);
or U9825 (N_9825,N_4823,N_4208);
nor U9826 (N_9826,N_872,N_3722);
or U9827 (N_9827,N_2559,N_3821);
nor U9828 (N_9828,N_3942,N_4447);
or U9829 (N_9829,N_4214,N_1726);
or U9830 (N_9830,N_3866,N_2726);
nand U9831 (N_9831,N_1062,N_1973);
or U9832 (N_9832,N_3384,N_1941);
and U9833 (N_9833,N_3172,N_449);
nor U9834 (N_9834,N_1080,N_152);
and U9835 (N_9835,N_1164,N_1367);
and U9836 (N_9836,N_2943,N_4748);
nor U9837 (N_9837,N_2395,N_3590);
or U9838 (N_9838,N_419,N_2740);
and U9839 (N_9839,N_343,N_4614);
nand U9840 (N_9840,N_1475,N_4752);
nand U9841 (N_9841,N_3694,N_2108);
nor U9842 (N_9842,N_4384,N_3921);
nor U9843 (N_9843,N_665,N_525);
or U9844 (N_9844,N_4790,N_2931);
or U9845 (N_9845,N_3285,N_937);
or U9846 (N_9846,N_3423,N_4670);
or U9847 (N_9847,N_1773,N_3312);
nor U9848 (N_9848,N_2344,N_4254);
nand U9849 (N_9849,N_1846,N_3428);
nor U9850 (N_9850,N_3272,N_3676);
nor U9851 (N_9851,N_2253,N_4426);
or U9852 (N_9852,N_2317,N_1957);
and U9853 (N_9853,N_4063,N_647);
and U9854 (N_9854,N_1612,N_1606);
or U9855 (N_9855,N_2638,N_1048);
or U9856 (N_9856,N_3598,N_1200);
nand U9857 (N_9857,N_428,N_1035);
or U9858 (N_9858,N_307,N_783);
and U9859 (N_9859,N_4364,N_1226);
nand U9860 (N_9860,N_3079,N_3325);
and U9861 (N_9861,N_4423,N_2599);
nor U9862 (N_9862,N_4932,N_4242);
or U9863 (N_9863,N_3105,N_2834);
nand U9864 (N_9864,N_4872,N_4832);
nor U9865 (N_9865,N_3182,N_773);
or U9866 (N_9866,N_2375,N_1368);
nor U9867 (N_9867,N_287,N_2773);
nand U9868 (N_9868,N_1093,N_4598);
or U9869 (N_9869,N_493,N_235);
nand U9870 (N_9870,N_4105,N_2158);
and U9871 (N_9871,N_1866,N_3403);
nor U9872 (N_9872,N_4194,N_3192);
nor U9873 (N_9873,N_12,N_3528);
and U9874 (N_9874,N_444,N_4511);
or U9875 (N_9875,N_37,N_4347);
nand U9876 (N_9876,N_256,N_3768);
and U9877 (N_9877,N_2878,N_4098);
and U9878 (N_9878,N_245,N_3455);
nand U9879 (N_9879,N_3894,N_4302);
or U9880 (N_9880,N_1781,N_927);
and U9881 (N_9881,N_2258,N_2706);
and U9882 (N_9882,N_1683,N_2357);
nand U9883 (N_9883,N_2326,N_995);
or U9884 (N_9884,N_1185,N_3478);
nor U9885 (N_9885,N_81,N_2338);
or U9886 (N_9886,N_2465,N_2615);
nand U9887 (N_9887,N_4167,N_1017);
or U9888 (N_9888,N_979,N_3570);
and U9889 (N_9889,N_4879,N_407);
and U9890 (N_9890,N_3245,N_2927);
or U9891 (N_9891,N_1481,N_2936);
nand U9892 (N_9892,N_1234,N_4027);
or U9893 (N_9893,N_196,N_4511);
and U9894 (N_9894,N_2351,N_4030);
nor U9895 (N_9895,N_3000,N_2915);
nor U9896 (N_9896,N_575,N_1182);
and U9897 (N_9897,N_3578,N_1789);
nand U9898 (N_9898,N_382,N_1426);
and U9899 (N_9899,N_1118,N_1414);
or U9900 (N_9900,N_1588,N_2013);
or U9901 (N_9901,N_2903,N_2805);
and U9902 (N_9902,N_475,N_1325);
or U9903 (N_9903,N_2765,N_1452);
or U9904 (N_9904,N_299,N_589);
nand U9905 (N_9905,N_1042,N_2852);
nand U9906 (N_9906,N_3309,N_3630);
nand U9907 (N_9907,N_2951,N_2725);
or U9908 (N_9908,N_3727,N_2023);
nand U9909 (N_9909,N_2858,N_1720);
or U9910 (N_9910,N_1514,N_2213);
and U9911 (N_9911,N_2934,N_2269);
or U9912 (N_9912,N_4620,N_4636);
nand U9913 (N_9913,N_2787,N_2922);
and U9914 (N_9914,N_2824,N_1143);
nor U9915 (N_9915,N_925,N_4695);
nor U9916 (N_9916,N_3283,N_2562);
or U9917 (N_9917,N_2713,N_2764);
or U9918 (N_9918,N_2545,N_550);
or U9919 (N_9919,N_4363,N_2767);
or U9920 (N_9920,N_4481,N_3041);
and U9921 (N_9921,N_3211,N_4752);
nor U9922 (N_9922,N_1835,N_2554);
and U9923 (N_9923,N_3727,N_1518);
nor U9924 (N_9924,N_2787,N_480);
xnor U9925 (N_9925,N_4109,N_4528);
and U9926 (N_9926,N_2033,N_2678);
nor U9927 (N_9927,N_9,N_3509);
or U9928 (N_9928,N_4605,N_872);
or U9929 (N_9929,N_3972,N_968);
and U9930 (N_9930,N_515,N_4266);
or U9931 (N_9931,N_776,N_968);
or U9932 (N_9932,N_1018,N_731);
nor U9933 (N_9933,N_3571,N_2221);
nor U9934 (N_9934,N_268,N_4635);
nand U9935 (N_9935,N_3044,N_1954);
and U9936 (N_9936,N_4250,N_725);
nor U9937 (N_9937,N_3205,N_191);
or U9938 (N_9938,N_27,N_3588);
and U9939 (N_9939,N_2515,N_993);
and U9940 (N_9940,N_3131,N_3099);
and U9941 (N_9941,N_2672,N_2804);
nand U9942 (N_9942,N_4114,N_4404);
nand U9943 (N_9943,N_841,N_3982);
and U9944 (N_9944,N_1293,N_811);
nand U9945 (N_9945,N_4164,N_2547);
or U9946 (N_9946,N_2608,N_781);
and U9947 (N_9947,N_134,N_3320);
nor U9948 (N_9948,N_3820,N_1357);
and U9949 (N_9949,N_4740,N_2765);
or U9950 (N_9950,N_4456,N_413);
nand U9951 (N_9951,N_1978,N_2114);
nand U9952 (N_9952,N_4565,N_4246);
or U9953 (N_9953,N_3312,N_4421);
and U9954 (N_9954,N_577,N_1565);
nand U9955 (N_9955,N_1932,N_924);
nand U9956 (N_9956,N_840,N_3832);
nand U9957 (N_9957,N_1891,N_2363);
nor U9958 (N_9958,N_802,N_1674);
nand U9959 (N_9959,N_3079,N_2087);
and U9960 (N_9960,N_1710,N_4679);
and U9961 (N_9961,N_1555,N_1024);
or U9962 (N_9962,N_2745,N_4917);
or U9963 (N_9963,N_1430,N_418);
or U9964 (N_9964,N_1691,N_4624);
nand U9965 (N_9965,N_1,N_4482);
or U9966 (N_9966,N_289,N_3888);
or U9967 (N_9967,N_4021,N_1751);
nand U9968 (N_9968,N_3081,N_3992);
nor U9969 (N_9969,N_451,N_645);
nor U9970 (N_9970,N_2631,N_925);
nand U9971 (N_9971,N_2019,N_3593);
nand U9972 (N_9972,N_2392,N_3465);
xor U9973 (N_9973,N_459,N_491);
or U9974 (N_9974,N_3010,N_1911);
nor U9975 (N_9975,N_3944,N_3669);
nor U9976 (N_9976,N_2804,N_947);
nand U9977 (N_9977,N_938,N_2467);
nand U9978 (N_9978,N_1224,N_1542);
nor U9979 (N_9979,N_932,N_4781);
nand U9980 (N_9980,N_935,N_3729);
and U9981 (N_9981,N_1748,N_2201);
and U9982 (N_9982,N_2848,N_1686);
or U9983 (N_9983,N_3430,N_1293);
and U9984 (N_9984,N_505,N_4921);
nand U9985 (N_9985,N_4006,N_4199);
or U9986 (N_9986,N_1139,N_3395);
and U9987 (N_9987,N_1683,N_660);
nor U9988 (N_9988,N_3546,N_173);
nand U9989 (N_9989,N_2573,N_3889);
nand U9990 (N_9990,N_813,N_722);
nor U9991 (N_9991,N_3459,N_306);
nor U9992 (N_9992,N_1592,N_3426);
nand U9993 (N_9993,N_4130,N_2895);
or U9994 (N_9994,N_3521,N_3883);
nand U9995 (N_9995,N_2518,N_3322);
nand U9996 (N_9996,N_1096,N_1655);
or U9997 (N_9997,N_802,N_1591);
or U9998 (N_9998,N_1788,N_2635);
and U9999 (N_9999,N_2245,N_1621);
nor U10000 (N_10000,N_5556,N_9269);
and U10001 (N_10001,N_6046,N_6061);
nand U10002 (N_10002,N_6440,N_8607);
nand U10003 (N_10003,N_7797,N_6762);
nand U10004 (N_10004,N_8506,N_7180);
nand U10005 (N_10005,N_5674,N_7382);
and U10006 (N_10006,N_6935,N_8274);
nand U10007 (N_10007,N_9218,N_8981);
nor U10008 (N_10008,N_5699,N_6251);
and U10009 (N_10009,N_8832,N_5055);
nor U10010 (N_10010,N_7102,N_6719);
and U10011 (N_10011,N_6337,N_6274);
nor U10012 (N_10012,N_5973,N_9879);
nor U10013 (N_10013,N_8386,N_8530);
nor U10014 (N_10014,N_5801,N_5914);
nor U10015 (N_10015,N_7188,N_9579);
and U10016 (N_10016,N_8139,N_9621);
and U10017 (N_10017,N_5080,N_8884);
or U10018 (N_10018,N_7848,N_5191);
or U10019 (N_10019,N_5423,N_6032);
or U10020 (N_10020,N_5348,N_8923);
nor U10021 (N_10021,N_8562,N_9843);
nor U10022 (N_10022,N_8264,N_5396);
nor U10023 (N_10023,N_7458,N_7865);
nor U10024 (N_10024,N_6887,N_6107);
or U10025 (N_10025,N_7498,N_6172);
or U10026 (N_10026,N_8907,N_6280);
nor U10027 (N_10027,N_7740,N_7289);
nor U10028 (N_10028,N_9671,N_9943);
nor U10029 (N_10029,N_6875,N_8622);
nand U10030 (N_10030,N_8691,N_8427);
nor U10031 (N_10031,N_7245,N_7192);
or U10032 (N_10032,N_6739,N_6850);
nand U10033 (N_10033,N_5573,N_7973);
or U10034 (N_10034,N_7697,N_5721);
or U10035 (N_10035,N_9990,N_5135);
nand U10036 (N_10036,N_8171,N_6276);
and U10037 (N_10037,N_8715,N_9503);
nor U10038 (N_10038,N_5074,N_8678);
and U10039 (N_10039,N_5300,N_6306);
nand U10040 (N_10040,N_6245,N_9106);
nor U10041 (N_10041,N_8507,N_7581);
xnor U10042 (N_10042,N_7648,N_9273);
and U10043 (N_10043,N_9558,N_7216);
nor U10044 (N_10044,N_7628,N_5966);
nand U10045 (N_10045,N_5990,N_5864);
nor U10046 (N_10046,N_8540,N_5944);
nor U10047 (N_10047,N_7704,N_6416);
and U10048 (N_10048,N_9900,N_7656);
or U10049 (N_10049,N_6959,N_6231);
and U10050 (N_10050,N_8410,N_7995);
or U10051 (N_10051,N_8569,N_5459);
or U10052 (N_10052,N_7197,N_7889);
and U10053 (N_10053,N_9117,N_8974);
and U10054 (N_10054,N_6065,N_8773);
or U10055 (N_10055,N_7957,N_5697);
or U10056 (N_10056,N_5856,N_5620);
and U10057 (N_10057,N_8007,N_5871);
or U10058 (N_10058,N_6104,N_6545);
or U10059 (N_10059,N_9324,N_5068);
nand U10060 (N_10060,N_6173,N_7271);
and U10061 (N_10061,N_8851,N_6674);
and U10062 (N_10062,N_6813,N_7376);
nand U10063 (N_10063,N_7940,N_5416);
and U10064 (N_10064,N_8781,N_6248);
xor U10065 (N_10065,N_9901,N_7443);
or U10066 (N_10066,N_5660,N_7110);
nand U10067 (N_10067,N_8722,N_9052);
nor U10068 (N_10068,N_9443,N_7675);
or U10069 (N_10069,N_8253,N_7478);
or U10070 (N_10070,N_7296,N_5849);
and U10071 (N_10071,N_8709,N_6476);
nand U10072 (N_10072,N_6543,N_5593);
or U10073 (N_10073,N_6267,N_9340);
nor U10074 (N_10074,N_8431,N_8434);
xnor U10075 (N_10075,N_9794,N_9693);
and U10076 (N_10076,N_9413,N_6659);
or U10077 (N_10077,N_6426,N_9213);
and U10078 (N_10078,N_7378,N_7115);
or U10079 (N_10079,N_9424,N_7379);
and U10080 (N_10080,N_6080,N_9742);
nand U10081 (N_10081,N_7856,N_8278);
nand U10082 (N_10082,N_9044,N_7613);
nand U10083 (N_10083,N_6782,N_8340);
and U10084 (N_10084,N_7472,N_8319);
nand U10085 (N_10085,N_5291,N_5271);
and U10086 (N_10086,N_6682,N_6871);
nand U10087 (N_10087,N_9246,N_7429);
or U10088 (N_10088,N_7442,N_9423);
or U10089 (N_10089,N_6301,N_8873);
nand U10090 (N_10090,N_5527,N_9686);
nand U10091 (N_10091,N_9205,N_7061);
nand U10092 (N_10092,N_5298,N_6976);
nand U10093 (N_10093,N_6646,N_5277);
or U10094 (N_10094,N_5269,N_7359);
nor U10095 (N_10095,N_8254,N_5198);
nor U10096 (N_10096,N_9487,N_7732);
nand U10097 (N_10097,N_5469,N_9612);
or U10098 (N_10098,N_7263,N_8233);
nor U10099 (N_10099,N_6376,N_6811);
and U10100 (N_10100,N_5181,N_7918);
nor U10101 (N_10101,N_6077,N_6825);
and U10102 (N_10102,N_6213,N_8449);
nor U10103 (N_10103,N_5126,N_7905);
and U10104 (N_10104,N_9958,N_8774);
nor U10105 (N_10105,N_6764,N_8684);
or U10106 (N_10106,N_6743,N_5779);
nand U10107 (N_10107,N_6592,N_9851);
nand U10108 (N_10108,N_8675,N_9823);
or U10109 (N_10109,N_9048,N_9922);
nor U10110 (N_10110,N_6244,N_5663);
or U10111 (N_10111,N_7034,N_5369);
or U10112 (N_10112,N_6505,N_6638);
or U10113 (N_10113,N_5683,N_5006);
xor U10114 (N_10114,N_8658,N_5650);
and U10115 (N_10115,N_6473,N_7850);
nand U10116 (N_10116,N_5767,N_7333);
nand U10117 (N_10117,N_5594,N_7300);
nor U10118 (N_10118,N_5463,N_8797);
nand U10119 (N_10119,N_7570,N_7463);
nor U10120 (N_10120,N_5398,N_6726);
or U10121 (N_10121,N_7313,N_9198);
and U10122 (N_10122,N_8258,N_9908);
nand U10123 (N_10123,N_6938,N_7605);
and U10124 (N_10124,N_7974,N_8719);
and U10125 (N_10125,N_9972,N_6379);
nor U10126 (N_10126,N_9695,N_7608);
and U10127 (N_10127,N_6017,N_9880);
and U10128 (N_10128,N_8854,N_7982);
nand U10129 (N_10129,N_9435,N_6330);
or U10130 (N_10130,N_9708,N_6135);
or U10131 (N_10131,N_8296,N_6933);
nand U10132 (N_10132,N_9475,N_9027);
nor U10133 (N_10133,N_6981,N_5066);
nand U10134 (N_10134,N_9685,N_5471);
nand U10135 (N_10135,N_8619,N_8966);
nand U10136 (N_10136,N_9296,N_9867);
and U10137 (N_10137,N_7899,N_8766);
nor U10138 (N_10138,N_7710,N_9422);
or U10139 (N_10139,N_6859,N_7031);
and U10140 (N_10140,N_5585,N_7065);
or U10141 (N_10141,N_6684,N_5429);
or U10142 (N_10142,N_7037,N_7189);
nand U10143 (N_10143,N_5301,N_5977);
nand U10144 (N_10144,N_7389,N_8770);
or U10145 (N_10145,N_7947,N_8631);
and U10146 (N_10146,N_9986,N_8163);
or U10147 (N_10147,N_6314,N_6413);
and U10148 (N_10148,N_5497,N_7018);
and U10149 (N_10149,N_5168,N_8747);
nand U10150 (N_10150,N_9690,N_9816);
nand U10151 (N_10151,N_6908,N_6730);
nand U10152 (N_10152,N_7421,N_7325);
nand U10153 (N_10153,N_7992,N_5102);
and U10154 (N_10154,N_5377,N_7803);
and U10155 (N_10155,N_6751,N_9022);
or U10156 (N_10156,N_5393,N_7235);
or U10157 (N_10157,N_7910,N_9400);
or U10158 (N_10158,N_5194,N_5252);
or U10159 (N_10159,N_5983,N_9862);
or U10160 (N_10160,N_7521,N_9008);
nor U10161 (N_10161,N_7209,N_6150);
or U10162 (N_10162,N_9601,N_8858);
or U10163 (N_10163,N_6857,N_6230);
or U10164 (N_10164,N_8105,N_6686);
and U10165 (N_10165,N_8201,N_7044);
and U10166 (N_10166,N_9751,N_8841);
nor U10167 (N_10167,N_6309,N_5776);
nor U10168 (N_10168,N_6845,N_8457);
nor U10169 (N_10169,N_6613,N_9093);
nand U10170 (N_10170,N_6395,N_7367);
nand U10171 (N_10171,N_6443,N_6121);
nand U10172 (N_10172,N_8503,N_7738);
nand U10173 (N_10173,N_7595,N_5725);
nand U10174 (N_10174,N_7911,N_7211);
nand U10175 (N_10175,N_8203,N_6237);
nor U10176 (N_10176,N_8051,N_5927);
or U10177 (N_10177,N_6964,N_6161);
nor U10178 (N_10178,N_6670,N_6088);
and U10179 (N_10179,N_6785,N_8000);
and U10180 (N_10180,N_7532,N_6289);
and U10181 (N_10181,N_8932,N_8943);
or U10182 (N_10182,N_7920,N_5486);
nor U10183 (N_10183,N_9959,N_7248);
and U10184 (N_10184,N_6576,N_7097);
nand U10185 (N_10185,N_8284,N_9185);
and U10186 (N_10186,N_8630,N_9745);
nor U10187 (N_10187,N_5996,N_9945);
nand U10188 (N_10188,N_6369,N_5127);
or U10189 (N_10189,N_7924,N_5138);
nand U10190 (N_10190,N_8725,N_5691);
and U10191 (N_10191,N_7322,N_8147);
or U10192 (N_10192,N_9419,N_9462);
nand U10193 (N_10193,N_9358,N_7691);
or U10194 (N_10194,N_9268,N_6969);
and U10195 (N_10195,N_6240,N_5610);
or U10196 (N_10196,N_7474,N_9910);
nor U10197 (N_10197,N_8070,N_8897);
or U10198 (N_10198,N_9602,N_7128);
nand U10199 (N_10199,N_5521,N_9049);
nand U10200 (N_10200,N_9872,N_7091);
nand U10201 (N_10201,N_9662,N_7822);
or U10202 (N_10202,N_8094,N_5360);
or U10203 (N_10203,N_6821,N_6480);
nor U10204 (N_10204,N_7900,N_9500);
and U10205 (N_10205,N_7806,N_7591);
and U10206 (N_10206,N_6953,N_6790);
and U10207 (N_10207,N_6787,N_7393);
nor U10208 (N_10208,N_6937,N_9798);
and U10209 (N_10209,N_5645,N_5617);
nor U10210 (N_10210,N_9599,N_8086);
and U10211 (N_10211,N_6112,N_9194);
or U10212 (N_10212,N_7304,N_5531);
and U10213 (N_10213,N_5861,N_6948);
nand U10214 (N_10214,N_6652,N_6699);
nand U10215 (N_10215,N_5468,N_8523);
nand U10216 (N_10216,N_9878,N_8361);
nand U10217 (N_10217,N_7385,N_6770);
nor U10218 (N_10218,N_9129,N_7154);
nand U10219 (N_10219,N_6936,N_8515);
and U10220 (N_10220,N_6508,N_6129);
nor U10221 (N_10221,N_8522,N_9277);
nand U10222 (N_10222,N_8305,N_8988);
or U10223 (N_10223,N_7721,N_8793);
or U10224 (N_10224,N_9970,N_8124);
xnor U10225 (N_10225,N_6013,N_5355);
nand U10226 (N_10226,N_7970,N_7129);
and U10227 (N_10227,N_5110,N_8487);
and U10228 (N_10228,N_6057,N_8968);
and U10229 (N_10229,N_9494,N_6671);
or U10230 (N_10230,N_6229,N_5481);
or U10231 (N_10231,N_9393,N_6865);
and U10232 (N_10232,N_9221,N_7459);
or U10233 (N_10233,N_8938,N_7702);
nand U10234 (N_10234,N_9086,N_7694);
or U10235 (N_10235,N_5107,N_8387);
and U10236 (N_10236,N_5710,N_6383);
or U10237 (N_10237,N_6106,N_8601);
nor U10238 (N_10238,N_6010,N_5233);
and U10239 (N_10239,N_9013,N_5251);
nor U10240 (N_10240,N_8557,N_5470);
or U10241 (N_10241,N_5129,N_7662);
and U10242 (N_10242,N_7347,N_7764);
and U10243 (N_10243,N_6449,N_5222);
nor U10244 (N_10244,N_7058,N_7890);
nor U10245 (N_10245,N_9676,N_5104);
or U10246 (N_10246,N_8223,N_8861);
and U10247 (N_10247,N_5430,N_7301);
nor U10248 (N_10248,N_7767,N_9156);
nor U10249 (N_10249,N_5606,N_9075);
and U10250 (N_10250,N_5276,N_5790);
or U10251 (N_10251,N_6621,N_5193);
and U10252 (N_10252,N_8128,N_8760);
nand U10253 (N_10253,N_6678,N_7706);
and U10254 (N_10254,N_7559,N_6510);
nor U10255 (N_10255,N_5064,N_9190);
nor U10256 (N_10256,N_7722,N_7433);
nor U10257 (N_10257,N_5751,N_5955);
nand U10258 (N_10258,N_7334,N_7564);
and U10259 (N_10259,N_9598,N_8888);
or U10260 (N_10260,N_5530,N_5759);
or U10261 (N_10261,N_6370,N_7863);
and U10262 (N_10262,N_8418,N_9800);
nor U10263 (N_10263,N_9699,N_8597);
nor U10264 (N_10264,N_5239,N_9021);
and U10265 (N_10265,N_7201,N_9425);
or U10266 (N_10266,N_5073,N_8865);
and U10267 (N_10267,N_9208,N_9811);
and U10268 (N_10268,N_7161,N_9035);
and U10269 (N_10269,N_6446,N_8823);
and U10270 (N_10270,N_8686,N_5265);
nor U10271 (N_10271,N_9337,N_7109);
and U10272 (N_10272,N_5343,N_5908);
nand U10273 (N_10273,N_6332,N_5451);
or U10274 (N_10274,N_6818,N_9460);
and U10275 (N_10275,N_9804,N_8038);
and U10276 (N_10276,N_9292,N_9622);
nand U10277 (N_10277,N_8043,N_7365);
nand U10278 (N_10278,N_8137,N_6523);
and U10279 (N_10279,N_7361,N_6290);
nor U10280 (N_10280,N_6663,N_6047);
nand U10281 (N_10281,N_8210,N_5506);
or U10282 (N_10282,N_9114,N_9272);
and U10283 (N_10283,N_8756,N_7090);
nor U10284 (N_10284,N_5382,N_6374);
and U10285 (N_10285,N_7466,N_8959);
nand U10286 (N_10286,N_9531,N_9232);
and U10287 (N_10287,N_7555,N_5563);
and U10288 (N_10288,N_6950,N_9128);
nor U10289 (N_10289,N_8009,N_7768);
and U10290 (N_10290,N_9749,N_5304);
and U10291 (N_10291,N_5515,N_7545);
nor U10292 (N_10292,N_8947,N_8176);
nor U10293 (N_10293,N_6734,N_9130);
nor U10294 (N_10294,N_5465,N_5859);
or U10295 (N_10295,N_8422,N_7386);
and U10296 (N_10296,N_8821,N_8558);
and U10297 (N_10297,N_8555,N_6873);
nor U10298 (N_10298,N_5088,N_9654);
or U10299 (N_10299,N_9728,N_9061);
nor U10300 (N_10300,N_8824,N_6500);
nand U10301 (N_10301,N_6792,N_7026);
nor U10302 (N_10302,N_5101,N_8961);
and U10303 (N_10303,N_7494,N_6673);
nand U10304 (N_10304,N_7993,N_6533);
and U10305 (N_10305,N_5789,N_5568);
or U10306 (N_10306,N_8628,N_6463);
nor U10307 (N_10307,N_7885,N_5324);
or U10308 (N_10308,N_8552,N_6534);
nand U10309 (N_10309,N_5597,N_5082);
nor U10310 (N_10310,N_7649,N_8097);
nand U10311 (N_10311,N_9165,N_8430);
nor U10312 (N_10312,N_6468,N_9980);
or U10313 (N_10313,N_5796,N_7544);
nor U10314 (N_10314,N_8735,N_9000);
nand U10315 (N_10315,N_7875,N_6602);
and U10316 (N_10316,N_7309,N_7823);
nor U10317 (N_10317,N_6136,N_6362);
nand U10318 (N_10318,N_8759,N_7030);
and U10319 (N_10319,N_7854,N_9316);
nand U10320 (N_10320,N_7846,N_6212);
and U10321 (N_10321,N_5115,N_9866);
nand U10322 (N_10322,N_9732,N_5510);
and U10323 (N_10323,N_7081,N_6412);
nand U10324 (N_10324,N_6171,N_8906);
nand U10325 (N_10325,N_6155,N_5445);
nand U10326 (N_10326,N_9665,N_9037);
and U10327 (N_10327,N_7944,N_6322);
nor U10328 (N_10328,N_8772,N_8882);
nor U10329 (N_10329,N_6893,N_8291);
nand U10330 (N_10330,N_9588,N_8717);
and U10331 (N_10331,N_7895,N_5120);
xor U10332 (N_10332,N_6909,N_9444);
or U10333 (N_10333,N_7236,N_7210);
nor U10334 (N_10334,N_7549,N_6585);
and U10335 (N_10335,N_7931,N_7709);
or U10336 (N_10336,N_5844,N_5030);
and U10337 (N_10337,N_5057,N_8615);
nor U10338 (N_10338,N_6551,N_7729);
or U10339 (N_10339,N_5351,N_9678);
nor U10340 (N_10340,N_6823,N_8050);
nand U10341 (N_10341,N_7476,N_7047);
and U10342 (N_10342,N_5187,N_6093);
nor U10343 (N_10343,N_7265,N_5009);
nand U10344 (N_10344,N_9445,N_5547);
and U10345 (N_10345,N_6722,N_7832);
nand U10346 (N_10346,N_7703,N_8189);
or U10347 (N_10347,N_7215,N_5083);
and U10348 (N_10348,N_8579,N_5043);
and U10349 (N_10349,N_8461,N_8435);
and U10350 (N_10350,N_7810,N_5241);
xor U10351 (N_10351,N_8462,N_8328);
nor U10352 (N_10352,N_8196,N_5098);
or U10353 (N_10353,N_8842,N_8857);
and U10354 (N_10354,N_7111,N_9585);
and U10355 (N_10355,N_6997,N_9528);
or U10356 (N_10356,N_5449,N_7571);
nand U10357 (N_10357,N_8092,N_6250);
or U10358 (N_10358,N_6725,N_5903);
nand U10359 (N_10359,N_7191,N_7513);
nand U10360 (N_10360,N_6986,N_8269);
nand U10361 (N_10361,N_5877,N_9987);
or U10362 (N_10362,N_8004,N_8183);
and U10363 (N_10363,N_9799,N_5791);
nand U10364 (N_10364,N_9092,N_5456);
and U10365 (N_10365,N_6907,N_9944);
and U10366 (N_10366,N_8334,N_9160);
nand U10367 (N_10367,N_7624,N_8993);
nand U10368 (N_10368,N_7232,N_7711);
and U10369 (N_10369,N_9836,N_7755);
nor U10370 (N_10370,N_5605,N_5338);
and U10371 (N_10371,N_7609,N_7253);
or U10372 (N_10372,N_9385,N_6353);
or U10373 (N_10373,N_8478,N_6524);
and U10374 (N_10374,N_9111,N_5945);
and U10375 (N_10375,N_7765,N_5015);
nand U10376 (N_10376,N_5132,N_8452);
or U10377 (N_10377,N_8384,N_5569);
nand U10378 (N_10378,N_6452,N_6339);
or U10379 (N_10379,N_7566,N_9507);
nor U10380 (N_10380,N_6174,N_5152);
nand U10381 (N_10381,N_5406,N_6819);
nand U10382 (N_10382,N_8395,N_5409);
nor U10383 (N_10383,N_8153,N_7627);
nand U10384 (N_10384,N_7772,N_7486);
nor U10385 (N_10385,N_9465,N_5285);
and U10386 (N_10386,N_9930,N_6731);
nor U10387 (N_10387,N_6254,N_6874);
and U10388 (N_10388,N_7408,N_6522);
nand U10389 (N_10389,N_8811,N_8718);
or U10390 (N_10390,N_7354,N_9279);
or U10391 (N_10391,N_8589,N_6114);
or U10392 (N_10392,N_7139,N_7845);
nand U10393 (N_10393,N_6848,N_6115);
and U10394 (N_10394,N_5330,N_6016);
nand U10395 (N_10395,N_7160,N_9633);
nand U10396 (N_10396,N_8099,N_8860);
nand U10397 (N_10397,N_7348,N_8761);
or U10398 (N_10398,N_7901,N_5166);
or U10399 (N_10399,N_6268,N_9429);
nor U10400 (N_10400,N_5170,N_7470);
nand U10401 (N_10401,N_5346,N_8531);
nand U10402 (N_10402,N_7418,N_5923);
nand U10403 (N_10403,N_9555,N_6196);
or U10404 (N_10404,N_7923,N_9143);
or U10405 (N_10405,N_7269,N_8185);
nand U10406 (N_10406,N_9782,N_9321);
or U10407 (N_10407,N_7985,N_5206);
nor U10408 (N_10408,N_5078,N_8133);
or U10409 (N_10409,N_5418,N_9125);
nand U10410 (N_10410,N_6170,N_8875);
nand U10411 (N_10411,N_6528,N_7377);
nor U10412 (N_10412,N_5525,N_8621);
nor U10413 (N_10413,N_8587,N_8985);
and U10414 (N_10414,N_6842,N_8880);
and U10415 (N_10415,N_9939,N_7606);
and U10416 (N_10416,N_9565,N_5780);
nand U10417 (N_10417,N_5412,N_7661);
and U10418 (N_10418,N_9136,N_9216);
nand U10419 (N_10419,N_8707,N_9062);
nor U10420 (N_10420,N_6342,N_8481);
or U10421 (N_10421,N_6712,N_8998);
or U10422 (N_10422,N_6949,N_9711);
nor U10423 (N_10423,N_8162,N_7069);
nand U10424 (N_10424,N_6750,N_6346);
or U10425 (N_10425,N_8843,N_5705);
and U10426 (N_10426,N_6629,N_7186);
or U10427 (N_10427,N_5947,N_9498);
nand U10428 (N_10428,N_5069,N_5119);
nand U10429 (N_10429,N_5242,N_5722);
nor U10430 (N_10430,N_6559,N_6128);
or U10431 (N_10431,N_6134,N_7336);
nand U10432 (N_10432,N_9834,N_7909);
nand U10433 (N_10433,N_9744,N_9511);
nor U10434 (N_10434,N_6656,N_5503);
and U10435 (N_10435,N_9164,N_7956);
or U10436 (N_10436,N_9110,N_8277);
nand U10437 (N_10437,N_9295,N_9572);
or U10438 (N_10438,N_9078,N_6263);
xnor U10439 (N_10439,N_6068,N_7381);
or U10440 (N_10440,N_8467,N_6679);
and U10441 (N_10441,N_9530,N_8568);
and U10442 (N_10442,N_6096,N_7113);
nor U10443 (N_10443,N_8376,N_6367);
and U10444 (N_10444,N_9542,N_6816);
nand U10445 (N_10445,N_5906,N_9440);
and U10446 (N_10446,N_8787,N_7835);
or U10447 (N_10447,N_8828,N_9384);
or U10448 (N_10448,N_7552,N_6978);
and U10449 (N_10449,N_7739,N_6292);
nor U10450 (N_10450,N_8316,N_5411);
or U10451 (N_10451,N_5623,N_6485);
or U10452 (N_10452,N_9717,N_5148);
or U10453 (N_10453,N_8280,N_7237);
and U10454 (N_10454,N_7456,N_5245);
nand U10455 (N_10455,N_5283,N_8117);
or U10456 (N_10456,N_8542,N_8309);
or U10457 (N_10457,N_7094,N_6064);
or U10458 (N_10458,N_5898,N_8089);
and U10459 (N_10459,N_8371,N_9477);
or U10460 (N_10460,N_6403,N_9963);
nor U10461 (N_10461,N_7556,N_9640);
nor U10462 (N_10462,N_5608,N_5477);
or U10463 (N_10463,N_8475,N_9339);
and U10464 (N_10464,N_9858,N_7883);
or U10465 (N_10465,N_9071,N_9434);
nor U10466 (N_10466,N_6275,N_7482);
nand U10467 (N_10467,N_5060,N_8406);
nor U10468 (N_10468,N_9981,N_5384);
nor U10469 (N_10469,N_9016,N_5799);
nand U10470 (N_10470,N_5428,N_5777);
nand U10471 (N_10471,N_5146,N_6898);
nor U10472 (N_10472,N_6020,N_6755);
or U10473 (N_10473,N_6490,N_8742);
xor U10474 (N_10474,N_7092,N_9937);
and U10475 (N_10475,N_9535,N_7104);
and U10476 (N_10476,N_8207,N_5022);
nor U10477 (N_10477,N_7131,N_9195);
and U10478 (N_10478,N_9919,N_6633);
or U10479 (N_10479,N_9303,N_9705);
or U10480 (N_10480,N_8012,N_5008);
nand U10481 (N_10481,N_5176,N_9574);
or U10482 (N_10482,N_7255,N_8739);
or U10483 (N_10483,N_7267,N_6051);
and U10484 (N_10484,N_8152,N_8211);
nand U10485 (N_10485,N_9036,N_7604);
or U10486 (N_10486,N_9797,N_5425);
nor U10487 (N_10487,N_8640,N_8287);
and U10488 (N_10488,N_8915,N_7434);
and U10489 (N_10489,N_5352,N_8335);
or U10490 (N_10490,N_7533,N_9673);
nand U10491 (N_10491,N_6145,N_9084);
nor U10492 (N_10492,N_8146,N_9390);
or U10493 (N_10493,N_5524,N_7541);
nor U10494 (N_10494,N_9825,N_5546);
nor U10495 (N_10495,N_9853,N_5708);
and U10496 (N_10496,N_6558,N_5259);
and U10497 (N_10497,N_6757,N_8202);
or U10498 (N_10498,N_9895,N_6573);
nor U10499 (N_10499,N_8927,N_8792);
nor U10500 (N_10500,N_5720,N_5231);
or U10501 (N_10501,N_5733,N_8818);
and U10502 (N_10502,N_6914,N_5336);
or U10503 (N_10503,N_8486,N_8807);
xnor U10504 (N_10504,N_8169,N_6272);
nor U10505 (N_10505,N_9145,N_5354);
nor U10506 (N_10506,N_5444,N_5543);
xnor U10507 (N_10507,N_7960,N_5960);
nor U10508 (N_10508,N_5118,N_5192);
or U10509 (N_10509,N_8257,N_7127);
and U10510 (N_10510,N_7343,N_7335);
nor U10511 (N_10511,N_9014,N_8268);
and U10512 (N_10512,N_8967,N_5667);
nor U10513 (N_10513,N_9010,N_5240);
nor U10514 (N_10514,N_8876,N_9039);
or U10515 (N_10515,N_7063,N_9214);
or U10516 (N_10516,N_9831,N_6273);
nor U10517 (N_10517,N_6747,N_7499);
or U10518 (N_10518,N_5440,N_8941);
nor U10519 (N_10519,N_9418,N_9967);
or U10520 (N_10520,N_7099,N_5337);
nor U10521 (N_10521,N_8281,N_9283);
nand U10522 (N_10522,N_7495,N_6258);
and U10523 (N_10523,N_7022,N_6404);
or U10524 (N_10524,N_8276,N_7419);
and U10525 (N_10525,N_9200,N_8065);
nor U10526 (N_10526,N_7020,N_8156);
nand U10527 (N_10527,N_6716,N_8177);
nand U10528 (N_10528,N_8919,N_5402);
nor U10529 (N_10529,N_9824,N_7813);
nor U10530 (N_10530,N_5890,N_7542);
or U10531 (N_10531,N_8513,N_9677);
and U10532 (N_10532,N_8213,N_8389);
or U10533 (N_10533,N_6360,N_8563);
or U10534 (N_10534,N_7103,N_7546);
nand U10535 (N_10535,N_8931,N_9940);
or U10536 (N_10536,N_6456,N_7670);
and U10537 (N_10537,N_5928,N_8986);
nor U10538 (N_10538,N_5494,N_8380);
nand U10539 (N_10539,N_7280,N_6595);
nor U10540 (N_10540,N_9138,N_9567);
nand U10541 (N_10541,N_8238,N_7002);
or U10542 (N_10542,N_7747,N_6736);
and U10543 (N_10543,N_5392,N_7954);
nor U10544 (N_10544,N_7651,N_6605);
or U10545 (N_10545,N_9456,N_8846);
nor U10546 (N_10546,N_6915,N_7838);
and U10547 (N_10547,N_6192,N_5495);
and U10548 (N_10548,N_7547,N_8535);
nand U10549 (N_10549,N_5238,N_5975);
and U10550 (N_10550,N_5034,N_6767);
and U10551 (N_10551,N_9480,N_7718);
nor U10552 (N_10552,N_5860,N_8492);
nand U10553 (N_10553,N_9256,N_6407);
and U10554 (N_10554,N_6516,N_7519);
and U10555 (N_10555,N_7975,N_8491);
or U10556 (N_10556,N_5504,N_6351);
nand U10557 (N_10557,N_7321,N_6433);
and U10558 (N_10558,N_7312,N_9561);
and U10559 (N_10559,N_9822,N_8816);
or U10560 (N_10560,N_5290,N_5509);
nor U10561 (N_10561,N_7086,N_5208);
nor U10562 (N_10562,N_9864,N_5358);
nand U10563 (N_10563,N_7610,N_5851);
and U10564 (N_10564,N_5934,N_6085);
nor U10565 (N_10565,N_8062,N_5436);
and U10566 (N_10566,N_7288,N_6888);
and U10567 (N_10567,N_8444,N_7614);
nor U10568 (N_10568,N_6372,N_7511);
nand U10569 (N_10569,N_6968,N_9857);
and U10570 (N_10570,N_5072,N_7855);
or U10571 (N_10571,N_5334,N_9573);
or U10572 (N_10572,N_8005,N_5825);
and U10573 (N_10573,N_7870,N_8063);
or U10574 (N_10574,N_9399,N_5619);
nor U10575 (N_10575,N_8733,N_6913);
nand U10576 (N_10576,N_5281,N_6582);
and U10577 (N_10577,N_9226,N_5937);
and U10578 (N_10578,N_9302,N_8639);
and U10579 (N_10579,N_8834,N_6749);
nand U10580 (N_10580,N_9336,N_7228);
or U10581 (N_10581,N_9847,N_5824);
and U10582 (N_10582,N_9204,N_9239);
nor U10583 (N_10583,N_9826,N_9540);
or U10584 (N_10584,N_9684,N_5637);
and U10585 (N_10585,N_8235,N_9038);
or U10586 (N_10586,N_5802,N_9554);
and U10587 (N_10587,N_5103,N_6927);
nor U10588 (N_10588,N_5076,N_8485);
or U10589 (N_10589,N_6664,N_9330);
or U10590 (N_10590,N_5554,N_8353);
nor U10591 (N_10591,N_7064,N_8071);
or U10592 (N_10592,N_5682,N_8289);
nand U10593 (N_10593,N_9458,N_7229);
or U10594 (N_10594,N_7504,N_6998);
nor U10595 (N_10595,N_5413,N_9361);
or U10596 (N_10596,N_8886,N_9263);
nor U10597 (N_10597,N_7233,N_6846);
or U10598 (N_10598,N_9848,N_8637);
and U10599 (N_10599,N_7514,N_7200);
nand U10600 (N_10600,N_6220,N_7256);
nor U10601 (N_10601,N_7388,N_8076);
or U10602 (N_10602,N_6704,N_6036);
nor U10603 (N_10603,N_7036,N_6878);
or U10604 (N_10604,N_9485,N_6650);
and U10605 (N_10605,N_8785,N_6014);
xor U10606 (N_10606,N_9903,N_6181);
and U10607 (N_10607,N_6054,N_9806);
nand U10608 (N_10608,N_8646,N_7185);
or U10609 (N_10609,N_5748,N_5838);
and U10610 (N_10610,N_8890,N_8412);
or U10611 (N_10611,N_5086,N_8690);
nand U10612 (N_10612,N_8645,N_5302);
nor U10613 (N_10613,N_5113,N_6814);
nand U10614 (N_10614,N_7249,N_7349);
and U10615 (N_10615,N_5564,N_8158);
nor U10616 (N_10616,N_8660,N_6184);
nand U10617 (N_10617,N_7217,N_5004);
nor U10618 (N_10618,N_6738,N_7809);
nor U10619 (N_10619,N_8664,N_6518);
and U10620 (N_10620,N_7584,N_5327);
or U10621 (N_10621,N_5757,N_9366);
nor U10622 (N_10622,N_5917,N_9133);
and U10623 (N_10623,N_8838,N_8783);
and U10624 (N_10624,N_6539,N_9647);
and U10625 (N_10625,N_8574,N_7879);
or U10626 (N_10626,N_8891,N_9270);
nand U10627 (N_10627,N_5863,N_7006);
nand U10628 (N_10628,N_9754,N_8671);
nor U10629 (N_10629,N_7222,N_5311);
nand U10630 (N_10630,N_8963,N_6729);
nor U10631 (N_10631,N_8578,N_6098);
and U10632 (N_10632,N_9615,N_5046);
and U10633 (N_10633,N_9913,N_7946);
nand U10634 (N_10634,N_9680,N_6885);
or U10635 (N_10635,N_5702,N_9317);
and U10636 (N_10636,N_8543,N_6579);
nand U10637 (N_10637,N_8229,N_6023);
xnor U10638 (N_10638,N_6622,N_6100);
xor U10639 (N_10639,N_9447,N_9529);
nor U10640 (N_10640,N_7029,N_8442);
nor U10641 (N_10641,N_7087,N_9070);
nand U10642 (N_10642,N_8079,N_7942);
and U10643 (N_10643,N_6234,N_6393);
or U10644 (N_10644,N_5600,N_7719);
and U10645 (N_10645,N_7672,N_5771);
nor U10646 (N_10646,N_6753,N_7560);
nand U10647 (N_10647,N_7744,N_5654);
and U10648 (N_10648,N_7676,N_8383);
nand U10649 (N_10649,N_6975,N_5735);
nand U10650 (N_10650,N_5028,N_7663);
nand U10651 (N_10651,N_6955,N_8681);
and U10652 (N_10652,N_5822,N_9112);
nor U10653 (N_10653,N_7150,N_7133);
nor U10654 (N_10654,N_5764,N_8553);
or U10655 (N_10655,N_8697,N_9610);
nor U10656 (N_10656,N_7019,N_5993);
or U10657 (N_10657,N_5523,N_7475);
nand U10658 (N_10658,N_6578,N_5099);
and U10659 (N_10659,N_7578,N_5747);
nor U10660 (N_10660,N_7828,N_7903);
or U10661 (N_10661,N_9545,N_8323);
nor U10662 (N_10662,N_6099,N_7460);
and U10663 (N_10663,N_5769,N_8357);
xnor U10664 (N_10664,N_9163,N_7921);
or U10665 (N_10665,N_7851,N_9620);
and U10666 (N_10666,N_9609,N_6000);
and U10667 (N_10667,N_9403,N_6189);
nor U10668 (N_10668,N_8360,N_9884);
nand U10669 (N_10669,N_8632,N_6343);
or U10670 (N_10670,N_5133,N_9469);
or U10671 (N_10671,N_6916,N_7652);
nand U10672 (N_10672,N_7778,N_6496);
nor U10673 (N_10673,N_6478,N_5368);
nor U10674 (N_10674,N_6930,N_7683);
nand U10675 (N_10675,N_7598,N_5685);
nor U10676 (N_10676,N_6723,N_5453);
and U10677 (N_10677,N_5091,N_5414);
or U10678 (N_10678,N_5387,N_7306);
or U10679 (N_10679,N_9298,N_8040);
or U10680 (N_10680,N_6182,N_7949);
or U10681 (N_10681,N_8822,N_9603);
or U10682 (N_10682,N_6987,N_5105);
nor U10683 (N_10683,N_9357,N_6567);
nor U10684 (N_10684,N_9553,N_7685);
nand U10685 (N_10685,N_5033,N_9600);
and U10686 (N_10686,N_5447,N_6774);
or U10687 (N_10687,N_6198,N_8155);
or U10688 (N_10688,N_6203,N_5026);
or U10689 (N_10689,N_6146,N_7290);
or U10690 (N_10690,N_6527,N_5116);
nand U10691 (N_10691,N_9248,N_7461);
nor U10692 (N_10692,N_7487,N_8075);
or U10693 (N_10693,N_9551,N_7980);
nand U10694 (N_10694,N_7659,N_5968);
nor U10695 (N_10695,N_5084,N_6667);
nor U10696 (N_10696,N_9450,N_7345);
and U10697 (N_10697,N_8374,N_7785);
nor U10698 (N_10698,N_6952,N_8710);
and U10699 (N_10699,N_7144,N_7713);
or U10700 (N_10700,N_6474,N_8980);
nand U10701 (N_10701,N_8413,N_8356);
or U10702 (N_10702,N_9034,N_9722);
and U10703 (N_10703,N_7407,N_7820);
and U10704 (N_10704,N_8529,N_8061);
or U10705 (N_10705,N_6201,N_6619);
nand U10706 (N_10706,N_7773,N_6019);
nor U10707 (N_10707,N_8325,N_9490);
or U10708 (N_10708,N_8626,N_5052);
nand U10709 (N_10709,N_7100,N_6027);
nor U10710 (N_10710,N_7252,N_6772);
or U10711 (N_10711,N_6498,N_5612);
and U10712 (N_10712,N_9368,N_6502);
and U10713 (N_10713,N_6078,N_9351);
or U10714 (N_10714,N_8566,N_7314);
nor U10715 (N_10715,N_9294,N_6167);
nor U10716 (N_10716,N_6070,N_6598);
nand U10717 (N_10717,N_9829,N_8179);
or U10718 (N_10718,N_7868,N_9849);
or U10719 (N_10719,N_8167,N_7902);
or U10720 (N_10720,N_8157,N_7638);
or U10721 (N_10721,N_5805,N_5604);
nor U10722 (N_10722,N_8674,N_8330);
or U10723 (N_10723,N_9018,N_8649);
or U10724 (N_10724,N_5400,N_7368);
and U10725 (N_10725,N_7490,N_7815);
nor U10726 (N_10726,N_6479,N_5627);
nor U10727 (N_10727,N_8460,N_8836);
or U10728 (N_10728,N_7688,N_7134);
or U10729 (N_10729,N_7095,N_5312);
nand U10730 (N_10730,N_9063,N_8206);
and U10731 (N_10731,N_7563,N_9406);
nand U10732 (N_10732,N_6012,N_6381);
nand U10733 (N_10733,N_8957,N_8161);
nand U10734 (N_10734,N_8192,N_6428);
and U10735 (N_10735,N_8627,N_8910);
or U10736 (N_10736,N_9516,N_8477);
and U10737 (N_10737,N_6356,N_9859);
and U10738 (N_10738,N_7291,N_7330);
nand U10739 (N_10739,N_9242,N_6294);
nor U10740 (N_10740,N_6455,N_5599);
or U10741 (N_10741,N_6238,N_7213);
nand U10742 (N_10742,N_5437,N_7413);
nand U10743 (N_10743,N_5359,N_5865);
nor U10744 (N_10744,N_7225,N_9066);
nor U10745 (N_10745,N_9791,N_9360);
and U10746 (N_10746,N_7266,N_8394);
or U10747 (N_10747,N_9736,N_9240);
nand U10748 (N_10748,N_9257,N_5403);
and U10749 (N_10749,N_9787,N_6205);
and U10750 (N_10750,N_7793,N_9707);
and U10751 (N_10751,N_5474,N_5813);
nor U10752 (N_10752,N_7853,N_7760);
or U10753 (N_10753,N_5042,N_5012);
nand U10754 (N_10754,N_6302,N_6321);
nor U10755 (N_10755,N_7423,N_6840);
nand U10756 (N_10756,N_7175,N_9841);
or U10757 (N_10757,N_7350,N_8113);
or U10758 (N_10758,N_8221,N_9306);
and U10759 (N_10759,N_9278,N_6109);
nor U10760 (N_10760,N_8728,N_8165);
nand U10761 (N_10761,N_5742,N_5707);
or U10762 (N_10762,N_7025,N_5629);
and U10763 (N_10763,N_7976,N_5526);
nand U10764 (N_10764,N_7357,N_5763);
or U10765 (N_10765,N_9712,N_8738);
or U10766 (N_10766,N_9838,N_8720);
or U10767 (N_10767,N_8576,N_8170);
nor U10768 (N_10768,N_5885,N_9028);
nand U10769 (N_10769,N_9581,N_6784);
nor U10770 (N_10770,N_5581,N_5306);
nor U10771 (N_10771,N_7548,N_7374);
and U10772 (N_10772,N_7664,N_8236);
nand U10773 (N_10773,N_7893,N_5701);
nand U10774 (N_10774,N_5331,N_7807);
nor U10775 (N_10775,N_7181,N_6958);
or U10776 (N_10776,N_9793,N_9372);
or U10777 (N_10777,N_8241,N_5961);
nor U10778 (N_10778,N_7963,N_7427);
nor U10779 (N_10779,N_9889,N_5125);
or U10780 (N_10780,N_6758,N_7311);
and U10781 (N_10781,N_9057,N_6076);
or U10782 (N_10782,N_8453,N_9319);
nand U10783 (N_10783,N_5153,N_5997);
or U10784 (N_10784,N_7402,N_9342);
and U10785 (N_10785,N_6417,N_8944);
or U10786 (N_10786,N_9023,N_9902);
and U10787 (N_10787,N_5112,N_5092);
nand U10788 (N_10788,N_5434,N_8666);
and U10789 (N_10789,N_8519,N_5770);
nand U10790 (N_10790,N_8614,N_9367);
nor U10791 (N_10791,N_7705,N_8539);
nor U10792 (N_10792,N_7062,N_8482);
nor U10793 (N_10793,N_9761,N_9819);
and U10794 (N_10794,N_6385,N_7394);
nand U10795 (N_10795,N_7587,N_5940);
nor U10796 (N_10796,N_9152,N_9168);
nand U10797 (N_10797,N_5219,N_8642);
nor U10798 (N_10798,N_5752,N_6003);
and U10799 (N_10799,N_8073,N_6537);
nand U10800 (N_10800,N_7169,N_7015);
and U10801 (N_10801,N_5226,N_9446);
nor U10802 (N_10802,N_5848,N_8749);
and U10803 (N_10803,N_6359,N_7754);
and U10804 (N_10804,N_6943,N_8301);
or U10805 (N_10805,N_8423,N_8303);
or U10806 (N_10806,N_6015,N_8712);
or U10807 (N_10807,N_9898,N_9166);
and U10808 (N_10808,N_7583,N_9437);
and U10809 (N_10809,N_6226,N_9225);
and U10810 (N_10810,N_8734,N_5150);
and U10811 (N_10811,N_5561,N_6609);
or U10812 (N_10812,N_6041,N_8653);
or U10813 (N_10813,N_8310,N_7116);
nand U10814 (N_10814,N_6043,N_7916);
nor U10815 (N_10815,N_8337,N_8782);
and U10816 (N_10816,N_7791,N_8517);
nand U10817 (N_10817,N_7998,N_8730);
and U10818 (N_10818,N_9484,N_5988);
or U10819 (N_10819,N_8724,N_7358);
nand U10820 (N_10820,N_7000,N_9335);
nor U10821 (N_10821,N_5766,N_7106);
nand U10822 (N_10822,N_8527,N_7007);
and U10823 (N_10823,N_5549,N_8127);
nand U10824 (N_10824,N_6741,N_9897);
nand U10825 (N_10825,N_7529,N_8682);
and U10826 (N_10826,N_6541,N_6560);
nor U10827 (N_10827,N_6756,N_5924);
and U10828 (N_10828,N_6328,N_9888);
nor U10829 (N_10829,N_9224,N_9772);
nor U10830 (N_10830,N_6861,N_9481);
and U10831 (N_10831,N_7305,N_9548);
or U10832 (N_10832,N_8017,N_5688);
or U10833 (N_10833,N_5478,N_9291);
or U10834 (N_10834,N_5555,N_7303);
xnor U10835 (N_10835,N_9549,N_7634);
nor U10836 (N_10836,N_6960,N_8688);
or U10837 (N_10837,N_8087,N_6891);
nand U10838 (N_10838,N_8228,N_9290);
and U10839 (N_10839,N_8143,N_9814);
nand U10840 (N_10840,N_5981,N_7568);
nand U10841 (N_10841,N_8871,N_6901);
nand U10842 (N_10842,N_6239,N_8283);
nand U10843 (N_10843,N_8575,N_7392);
or U10844 (N_10844,N_5893,N_6457);
nand U10845 (N_10845,N_6961,N_5999);
and U10846 (N_10846,N_7138,N_9534);
nor U10847 (N_10847,N_7405,N_5641);
xnor U10848 (N_10848,N_5160,N_7052);
nand U10849 (N_10849,N_9096,N_6336);
nor U10850 (N_10850,N_9969,N_8218);
nand U10851 (N_10851,N_9318,N_7727);
nand U10852 (N_10852,N_8794,N_7827);
nand U10853 (N_10853,N_9759,N_8757);
or U10854 (N_10854,N_8784,N_6809);
and U10855 (N_10855,N_7576,N_8365);
nor U10856 (N_10856,N_7395,N_9636);
or U10857 (N_10857,N_5558,N_8020);
nor U10858 (N_10858,N_5755,N_6617);
nand U10859 (N_10859,N_9628,N_5212);
and U10860 (N_10860,N_8641,N_8900);
nor U10861 (N_10861,N_7517,N_7431);
nor U10862 (N_10862,N_5728,N_7049);
and U10863 (N_10863,N_7712,N_5000);
nor U10864 (N_10864,N_9597,N_9228);
xor U10865 (N_10865,N_5874,N_8916);
nor U10866 (N_10866,N_5686,N_5340);
nand U10867 (N_10867,N_5698,N_6236);
nor U10868 (N_10868,N_9098,N_9352);
nor U10869 (N_10869,N_7426,N_8024);
and U10870 (N_10870,N_7452,N_8594);
or U10871 (N_10871,N_5694,N_5536);
nor U10872 (N_10872,N_9774,N_5854);
or U10873 (N_10873,N_8536,N_7390);
and U10874 (N_10874,N_7462,N_6329);
nand U10875 (N_10875,N_8788,N_6791);
nor U10876 (N_10876,N_7798,N_9323);
nor U10877 (N_10877,N_7176,N_9409);
nor U10878 (N_10878,N_5492,N_7156);
nor U10879 (N_10879,N_6928,N_5552);
or U10880 (N_10880,N_7616,N_5491);
nor U10881 (N_10881,N_8878,N_8329);
nor U10882 (N_10882,N_7699,N_5220);
or U10883 (N_10883,N_8085,N_5875);
and U10884 (N_10884,N_8288,N_8741);
nor U10885 (N_10885,N_5054,N_5432);
nand U10886 (N_10886,N_9807,N_8965);
nor U10887 (N_10887,N_9132,N_5891);
xnor U10888 (N_10888,N_9890,N_9155);
nor U10889 (N_10889,N_9449,N_9150);
or U10890 (N_10890,N_5778,N_5765);
and U10891 (N_10891,N_9436,N_6980);
and U10892 (N_10892,N_5284,N_6879);
or U10893 (N_10893,N_5321,N_5476);
and U10894 (N_10894,N_9584,N_7001);
or U10895 (N_10895,N_6575,N_8991);
nor U10896 (N_10896,N_5575,N_8343);
and U10897 (N_10897,N_6442,N_7515);
nand U10898 (N_10898,N_8266,N_8037);
nand U10899 (N_10899,N_6834,N_6470);
nor U10900 (N_10900,N_7234,N_6087);
or U10901 (N_10901,N_8883,N_6116);
nor U10902 (N_10902,N_9203,N_5274);
or U10903 (N_10903,N_6951,N_6929);
or U10904 (N_10904,N_6165,N_8046);
nand U10905 (N_10905,N_9047,N_7320);
or U10906 (N_10906,N_5464,N_9504);
and U10907 (N_10907,N_9674,N_9381);
nor U10908 (N_10908,N_6977,N_6810);
or U10909 (N_10909,N_6125,N_9730);
and U10910 (N_10910,N_7422,N_7666);
or U10911 (N_10911,N_6450,N_6265);
or U10912 (N_10912,N_9979,N_8359);
or U10913 (N_10913,N_8399,N_8190);
and U10914 (N_10914,N_6399,N_6683);
nor U10915 (N_10915,N_5114,N_5901);
nor U10916 (N_10916,N_7677,N_9669);
nor U10917 (N_10917,N_8154,N_5255);
nand U10918 (N_10918,N_7859,N_9559);
nor U10919 (N_10919,N_5915,N_5024);
nor U10920 (N_10920,N_6042,N_9766);
nand U10921 (N_10921,N_7043,N_7708);
nand U10922 (N_10922,N_5389,N_8969);
nand U10923 (N_10923,N_7400,N_8514);
or U10924 (N_10924,N_7945,N_6319);
nand U10925 (N_10925,N_5535,N_5473);
and U10926 (N_10926,N_6906,N_9438);
and U10927 (N_10927,N_9350,N_5642);
xnor U10928 (N_10928,N_7554,N_5932);
or U10929 (N_10929,N_6503,N_5933);
nand U10930 (N_10930,N_6858,N_8680);
nor U10931 (N_10931,N_8617,N_5579);
nor U10932 (N_10932,N_9891,N_9151);
nor U10933 (N_10933,N_6357,N_8771);
and U10934 (N_10934,N_5909,N_5140);
nand U10935 (N_10935,N_8402,N_8746);
nor U10936 (N_10936,N_6548,N_7804);
and U10937 (N_10937,N_5740,N_5806);
and U10938 (N_10938,N_7004,N_8072);
or U10939 (N_10939,N_5002,N_5189);
and U10940 (N_10940,N_9689,N_8499);
nor U10941 (N_10941,N_9430,N_8972);
or U10942 (N_10942,N_5957,N_6831);
and U10943 (N_10943,N_8837,N_6347);
nand U10944 (N_10944,N_8994,N_8804);
or U10945 (N_10945,N_9334,N_9905);
and U10946 (N_10946,N_5852,N_9805);
nor U10947 (N_10947,N_6348,N_9353);
and U10948 (N_10948,N_6187,N_8148);
and U10949 (N_10949,N_7951,N_5196);
nand U10950 (N_10950,N_8249,N_5718);
nor U10951 (N_10951,N_7227,N_7936);
and U10952 (N_10952,N_9161,N_5053);
or U10953 (N_10953,N_9080,N_7406);
or U10954 (N_10954,N_5315,N_6974);
nand U10955 (N_10955,N_7146,N_5310);
nor U10956 (N_10956,N_6807,N_6702);
or U10957 (N_10957,N_8001,N_5895);
and U10958 (N_10958,N_7728,N_5616);
nand U10959 (N_10959,N_5567,N_9120);
nand U10960 (N_10960,N_5056,N_5134);
and U10961 (N_10961,N_6631,N_7650);
and U10962 (N_10962,N_9582,N_7684);
and U10963 (N_10963,N_5768,N_7059);
and U10964 (N_10964,N_5808,N_9193);
or U10965 (N_10965,N_8740,N_5965);
and U10966 (N_10966,N_9637,N_5706);
and U10967 (N_10967,N_8827,N_5842);
nand U10968 (N_10968,N_8852,N_5540);
or U10969 (N_10969,N_6763,N_8436);
or U10970 (N_10970,N_8752,N_5040);
nand U10971 (N_10971,N_6151,N_9614);
nand U10972 (N_10972,N_8704,N_5149);
nand U10973 (N_10973,N_7978,N_6271);
nor U10974 (N_10974,N_6363,N_9991);
or U10975 (N_10975,N_7857,N_9105);
and U10976 (N_10976,N_6430,N_9017);
nand U10977 (N_10977,N_9941,N_7908);
nor U10978 (N_10978,N_9953,N_9513);
nor U10979 (N_10979,N_8973,N_5136);
and U10980 (N_10980,N_5803,N_9015);
or U10981 (N_10981,N_9266,N_8438);
nor U10982 (N_10982,N_6031,N_9099);
and U10983 (N_10983,N_8194,N_8348);
nor U10984 (N_10984,N_6458,N_5576);
nor U10985 (N_10985,N_6299,N_8795);
nand U10986 (N_10986,N_7137,N_5010);
or U10987 (N_10987,N_9192,N_6746);
nor U10988 (N_10988,N_5417,N_8262);
xor U10989 (N_10989,N_9904,N_8670);
and U10990 (N_10990,N_7259,N_6312);
and U10991 (N_10991,N_9012,N_6985);
or U10992 (N_10992,N_9315,N_7881);
and U10993 (N_10993,N_7750,N_6111);
or U10994 (N_10994,N_5077,N_5894);
and U10995 (N_10995,N_9726,N_6493);
and U10996 (N_10996,N_8066,N_8088);
nand U10997 (N_10997,N_5391,N_8894);
and U10998 (N_10998,N_6513,N_5551);
nor U10999 (N_10999,N_7543,N_9113);
and U11000 (N_11000,N_7847,N_7636);
nor U11001 (N_11001,N_6554,N_6038);
and U11002 (N_11002,N_5237,N_7603);
nand U11003 (N_11003,N_9102,N_5570);
and U11004 (N_11004,N_6300,N_5374);
nand U11005 (N_11005,N_6860,N_9255);
or U11006 (N_11006,N_7796,N_9282);
nor U11007 (N_11007,N_6798,N_9002);
nand U11008 (N_11008,N_8022,N_7525);
nor U11009 (N_11009,N_8166,N_8470);
and U11010 (N_11010,N_6044,N_6597);
or U11011 (N_11011,N_6880,N_6983);
nand U11012 (N_11012,N_6995,N_8098);
or U11013 (N_11013,N_9348,N_7964);
nand U11014 (N_11014,N_7988,N_9996);
nand U11015 (N_11015,N_7276,N_6776);
nand U11016 (N_11016,N_5858,N_6401);
nor U11017 (N_11017,N_6657,N_8318);
nand U11018 (N_11018,N_7024,N_5836);
nor U11019 (N_11019,N_8528,N_5630);
or U11020 (N_11020,N_5364,N_6624);
and U11021 (N_11021,N_5332,N_9267);
and U11022 (N_11022,N_9648,N_6669);
and U11023 (N_11023,N_7887,N_5972);
and U11024 (N_11024,N_7489,N_5659);
nand U11025 (N_11025,N_5935,N_8572);
or U11026 (N_11026,N_7079,N_7928);
xor U11027 (N_11027,N_5184,N_8501);
and U11028 (N_11028,N_8654,N_8789);
nand U11029 (N_11029,N_9116,N_9382);
and U11030 (N_11030,N_8036,N_7351);
nand U11031 (N_11031,N_6469,N_9064);
nand U11032 (N_11032,N_7873,N_8936);
or U11033 (N_11033,N_9174,N_7308);
nand U11034 (N_11034,N_5815,N_8469);
or U11035 (N_11035,N_6962,N_5866);
or U11036 (N_11036,N_9899,N_9954);
or U11037 (N_11037,N_9104,N_6611);
or U11038 (N_11038,N_8554,N_6530);
nor U11039 (N_11039,N_8300,N_6410);
or U11040 (N_11040,N_9177,N_7535);
and U11041 (N_11041,N_8659,N_5793);
nand U11042 (N_11042,N_7182,N_9591);
and U11043 (N_11043,N_6481,N_8116);
nor U11044 (N_11044,N_9144,N_7869);
nor U11045 (N_11045,N_6033,N_6285);
or U11046 (N_11046,N_7724,N_9731);
nand U11047 (N_11047,N_6317,N_5011);
nor U11048 (N_11048,N_9779,N_7415);
nand U11049 (N_11049,N_6235,N_7929);
nor U11050 (N_11050,N_6439,N_5305);
nand U11051 (N_11051,N_5075,N_6323);
or U11052 (N_11052,N_6886,N_8132);
nand U11053 (N_11053,N_6852,N_8777);
and U11054 (N_11054,N_8977,N_9896);
or U11055 (N_11055,N_6462,N_8342);
and U11056 (N_11056,N_8693,N_8358);
nor U11057 (N_11057,N_9073,N_7257);
nand U11058 (N_11058,N_5565,N_7319);
or U11059 (N_11059,N_7310,N_5736);
nand U11060 (N_11060,N_5726,N_5541);
nand U11061 (N_11061,N_6291,N_5820);
nand U11062 (N_11062,N_8059,N_5595);
nor U11063 (N_11063,N_7621,N_5716);
or U11064 (N_11064,N_9734,N_8997);
nand U11065 (N_11065,N_5978,N_5316);
nor U11066 (N_11066,N_8096,N_6375);
nor U11067 (N_11067,N_9842,N_8160);
nor U11068 (N_11068,N_8778,N_9617);
or U11069 (N_11069,N_8149,N_7105);
and U11070 (N_11070,N_9428,N_9079);
nand U11071 (N_11071,N_8953,N_7867);
nand U11072 (N_11072,N_9389,N_5256);
nand U11073 (N_11073,N_5508,N_9672);
nand U11074 (N_11074,N_5724,N_7324);
or U11075 (N_11075,N_9875,N_8216);
nand U11076 (N_11076,N_5936,N_9363);
or U11077 (N_11077,N_8379,N_9499);
nor U11078 (N_11078,N_6824,N_8853);
nor U11079 (N_11079,N_9589,N_7934);
nand U11080 (N_11080,N_9948,N_5544);
nand U11081 (N_11081,N_8351,N_9427);
nand U11082 (N_11082,N_5518,N_6666);
nor U11083 (N_11083,N_8984,N_8178);
nand U11084 (N_11084,N_9586,N_7328);
and U11085 (N_11085,N_8045,N_9929);
and U11086 (N_11086,N_6642,N_7907);
nor U11087 (N_11087,N_9191,N_6318);
nand U11088 (N_11088,N_9649,N_8810);
and U11089 (N_11089,N_5013,N_7371);
and U11090 (N_11090,N_5625,N_7632);
xnor U11091 (N_11091,N_9817,N_7927);
xor U11092 (N_11092,N_9522,N_5263);
or U11093 (N_11093,N_7411,N_8556);
or U11094 (N_11094,N_7078,N_6277);
and U11095 (N_11095,N_9696,N_6881);
nand U11096 (N_11096,N_5282,N_5234);
or U11097 (N_11097,N_7042,N_8306);
nand U11098 (N_11098,N_5931,N_5693);
nand U11099 (N_11099,N_5275,N_7293);
or U11100 (N_11100,N_8247,N_5520);
nor U11101 (N_11101,N_7170,N_8848);
and U11102 (N_11102,N_6789,N_6984);
nand U11103 (N_11103,N_6142,N_5458);
or U11104 (N_11104,N_9746,N_8002);
nor U11105 (N_11105,N_5876,N_6668);
nor U11106 (N_11106,N_9416,N_6195);
or U11107 (N_11107,N_6604,N_6862);
or U11108 (N_11108,N_8921,N_6035);
and U11109 (N_11109,N_8222,N_7488);
nand U11110 (N_11110,N_9375,N_8400);
and U11111 (N_11111,N_9041,N_5534);
and U11112 (N_11112,N_9650,N_9727);
nand U11113 (N_11113,N_9383,N_8011);
nand U11114 (N_11114,N_7720,N_8468);
or U11115 (N_11115,N_7569,N_9845);
or U11116 (N_11116,N_9916,N_8102);
or U11117 (N_11117,N_8251,N_8409);
or U11118 (N_11118,N_8864,N_5097);
nand U11119 (N_11119,N_9300,N_6759);
or U11120 (N_11120,N_5872,N_9792);
nor U11121 (N_11121,N_7646,N_5622);
or U11122 (N_11122,N_8570,N_7484);
nand U11123 (N_11123,N_9569,N_5826);
nand U11124 (N_11124,N_6471,N_7226);
nand U11125 (N_11125,N_7033,N_9915);
nand U11126 (N_11126,N_8084,N_8559);
nor U11127 (N_11127,N_7601,N_7919);
nor U11128 (N_11128,N_8541,N_9118);
nor U11129 (N_11129,N_5270,N_6697);
and U11130 (N_11130,N_6315,N_9220);
nand U11131 (N_11131,N_8567,N_8432);
nor U11132 (N_11132,N_8498,N_9127);
or U11133 (N_11133,N_6942,N_6495);
nor U11134 (N_11134,N_5571,N_5603);
nor U11135 (N_11135,N_8256,N_9984);
or U11136 (N_11136,N_9040,N_9396);
nand U11137 (N_11137,N_9169,N_7884);
or U11138 (N_11138,N_9844,N_7506);
nand U11139 (N_11139,N_7886,N_7251);
and U11140 (N_11140,N_5225,N_7445);
and U11141 (N_11141,N_7858,N_6324);
nand U11142 (N_11142,N_8495,N_8123);
nor U11143 (N_11143,N_5807,N_6847);
or U11144 (N_11144,N_9452,N_6529);
and U11145 (N_11145,N_5087,N_7585);
or U11146 (N_11146,N_5788,N_9961);
or U11147 (N_11147,N_7190,N_8373);
nand U11148 (N_11148,N_8844,N_6806);
nand U11149 (N_11149,N_9882,N_9223);
nand U11150 (N_11150,N_7896,N_5059);
and U11151 (N_11151,N_8215,N_8516);
and U11152 (N_11152,N_6593,N_9638);
nor U11153 (N_11153,N_6760,N_5236);
or U11154 (N_11154,N_5781,N_9245);
nor U11155 (N_11155,N_9183,N_8913);
or U11156 (N_11156,N_9083,N_9209);
nor U11157 (N_11157,N_9189,N_6056);
and U11158 (N_11158,N_8708,N_7876);
nand U11159 (N_11159,N_9411,N_6732);
xor U11160 (N_11160,N_9635,N_6639);
and U11161 (N_11161,N_8100,N_5185);
or U11162 (N_11162,N_8025,N_5756);
and U11163 (N_11163,N_5512,N_9471);
and U11164 (N_11164,N_9158,N_9785);
nor U11165 (N_11165,N_5985,N_6022);
nor U11166 (N_11166,N_7925,N_8590);
nand U11167 (N_11167,N_8455,N_8488);
nor U11168 (N_11168,N_6419,N_5483);
nor U11169 (N_11169,N_7505,N_9928);
nor U11170 (N_11170,N_6437,N_7327);
nand U11171 (N_11171,N_5804,N_5643);
nand U11172 (N_11172,N_6690,N_7250);
nor U11173 (N_11173,N_6021,N_6841);
or U11174 (N_11174,N_9332,N_9763);
and U11175 (N_11175,N_6103,N_5408);
or U11176 (N_11176,N_6127,N_9691);
nand U11177 (N_11177,N_5839,N_5475);
nand U11178 (N_11178,N_9918,N_8464);
nor U11179 (N_11179,N_6133,N_8583);
nor U11180 (N_11180,N_7667,N_9395);
and U11181 (N_11181,N_9489,N_5609);
nand U11182 (N_11182,N_8479,N_7961);
and U11183 (N_11183,N_6429,N_9483);
nand U11184 (N_11184,N_9713,N_8912);
nor U11185 (N_11185,N_7451,N_5715);
and U11186 (N_11186,N_6775,N_6820);
or U11187 (N_11187,N_6341,N_5958);
and U11188 (N_11188,N_5634,N_5900);
and U11189 (N_11189,N_5461,N_8706);
nor U11190 (N_11190,N_7551,N_8987);
and U11191 (N_11191,N_6123,N_5232);
nor U11192 (N_11192,N_6939,N_5018);
nand U11193 (N_11193,N_8407,N_5713);
xnor U11194 (N_11194,N_5253,N_7780);
or U11195 (N_11195,N_5167,N_5472);
and U11196 (N_11196,N_6255,N_8893);
or U11197 (N_11197,N_8885,N_6241);
or U11198 (N_11198,N_6414,N_6910);
nor U11199 (N_11199,N_7539,N_9215);
or U11200 (N_11200,N_9329,N_6562);
or U11201 (N_11201,N_8172,N_7787);
nor U11202 (N_11202,N_9739,N_7573);
and U11203 (N_11203,N_9861,N_6616);
nor U11204 (N_11204,N_8364,N_9783);
nor U11205 (N_11205,N_9123,N_7752);
nor U11206 (N_11206,N_7468,N_9846);
xor U11207 (N_11207,N_8392,N_5326);
and U11208 (N_11208,N_8537,N_6298);
and U11209 (N_11209,N_5810,N_9656);
and U11210 (N_11210,N_5749,N_9314);
and U11211 (N_11211,N_9076,N_7481);
or U11212 (N_11212,N_9706,N_8297);
nor U11213 (N_11213,N_6144,N_8126);
or U11214 (N_11214,N_6499,N_9201);
or U11215 (N_11215,N_9401,N_6577);
nand U11216 (N_11216,N_9188,N_9757);
nor U11217 (N_11217,N_7991,N_6900);
and U11218 (N_11218,N_9408,N_6921);
nand U11219 (N_11219,N_7246,N_9577);
or U11220 (N_11220,N_7085,N_9470);
nor U11221 (N_11221,N_6623,N_6991);
or U11222 (N_11222,N_5714,N_8052);
and U11223 (N_11223,N_6836,N_8829);
nand U11224 (N_11224,N_7048,N_8344);
nor U11225 (N_11225,N_8199,N_8497);
nand U11226 (N_11226,N_5653,N_8956);
or U11227 (N_11227,N_5921,N_8799);
nand U11228 (N_11228,N_5727,N_7816);
nor U11229 (N_11229,N_9697,N_5881);
nor U11230 (N_11230,N_6086,N_6610);
or U11231 (N_11231,N_8421,N_8078);
or U11232 (N_11232,N_7114,N_8625);
xnor U11233 (N_11233,N_7979,N_6090);
and U11234 (N_11234,N_8393,N_5250);
and U11235 (N_11235,N_9249,N_7307);
nand U11236 (N_11236,N_5574,N_9293);
and U11237 (N_11237,N_9107,N_7369);
nor U11238 (N_11238,N_7733,N_6694);
or U11239 (N_11239,N_9923,N_8960);
and U11240 (N_11240,N_7695,N_8687);
nand U11241 (N_11241,N_6795,N_8616);
nor U11242 (N_11242,N_7597,N_8090);
nand U11243 (N_11243,N_7120,N_8091);
nand U11244 (N_11244,N_9238,N_9645);
and U11245 (N_11245,N_6331,N_8368);
or U11246 (N_11246,N_6973,N_9328);
and U11247 (N_11247,N_5498,N_6069);
nor U11248 (N_11248,N_9251,N_7112);
or U11249 (N_11249,N_7698,N_9894);
nor U11250 (N_11250,N_5636,N_5488);
nor U11251 (N_11251,N_6583,N_7938);
nand U11252 (N_11252,N_7508,N_9262);
and U11253 (N_11253,N_7003,N_9681);
nor U11254 (N_11254,N_5442,N_5247);
nor U11255 (N_11255,N_7412,N_8754);
nor U11256 (N_11256,N_5289,N_6094);
and U11257 (N_11257,N_8835,N_9643);
nor U11258 (N_11258,N_9512,N_9510);
or U11259 (N_11259,N_7119,N_6208);
and U11260 (N_11260,N_7326,N_5845);
and U11261 (N_11261,N_5823,N_6920);
and U11262 (N_11262,N_5156,N_9619);
or U11263 (N_11263,N_8474,N_9921);
nor U11264 (N_11264,N_8839,N_8729);
nor U11265 (N_11265,N_6771,N_6696);
nand U11266 (N_11266,N_5157,N_7844);
or U11267 (N_11267,N_8548,N_8652);
nand U11268 (N_11268,N_8768,N_5335);
and U11269 (N_11269,N_8168,N_9914);
nand U11270 (N_11270,N_5415,N_8911);
or U11271 (N_11271,N_6695,N_8378);
nor U11272 (N_11272,N_6868,N_7602);
and U11273 (N_11273,N_6641,N_5926);
xnor U11274 (N_11274,N_6926,N_8242);
and U11275 (N_11275,N_9659,N_8714);
and U11276 (N_11276,N_6438,N_7199);
or U11277 (N_11277,N_5438,N_7177);
nor U11278 (N_11278,N_7012,N_9252);
or U11279 (N_11279,N_8275,N_5969);
nor U11280 (N_11280,N_7204,N_6672);
or U11281 (N_11281,N_5689,N_9557);
or U11282 (N_11282,N_6130,N_5837);
nand U11283 (N_11283,N_6486,N_8175);
or U11284 (N_11284,N_6802,N_9304);
and U11285 (N_11285,N_8948,N_7912);
or U11286 (N_11286,N_8564,N_6647);
or U11287 (N_11287,N_6521,N_8008);
xor U11288 (N_11288,N_9241,N_8580);
nor U11289 (N_11289,N_8122,N_7842);
and U11290 (N_11290,N_5760,N_5424);
nor U11291 (N_11291,N_5218,N_9976);
and U11292 (N_11292,N_6895,N_6919);
nand U11293 (N_11293,N_7736,N_9258);
or U11294 (N_11294,N_7136,N_6059);
or U11295 (N_11295,N_9873,N_7414);
and U11296 (N_11296,N_9058,N_6625);
nor U11297 (N_11297,N_5467,N_8585);
nand U11298 (N_11298,N_5675,N_6454);
and U11299 (N_11299,N_9042,N_6599);
nor U11300 (N_11300,N_7781,N_6822);
nor U11301 (N_11301,N_5712,N_8198);
nor U11302 (N_11302,N_9146,N_5904);
or U11303 (N_11303,N_8863,N_7157);
or U11304 (N_11304,N_7008,N_9931);
nand U11305 (N_11305,N_8355,N_7152);
and U11306 (N_11306,N_5821,N_6637);
nor U11307 (N_11307,N_6607,N_9613);
nand U11308 (N_11308,N_6266,N_7107);
or U11309 (N_11309,N_9082,N_9473);
nand U11310 (N_11310,N_7509,N_9032);
and U11311 (N_11311,N_5318,N_7510);
and U11312 (N_11312,N_8044,N_9421);
or U11313 (N_11313,N_7612,N_8618);
and U11314 (N_11314,N_7469,N_6944);
or U11315 (N_11315,N_5047,N_5294);
nand U11316 (N_11316,N_6089,N_9735);
nand U11317 (N_11317,N_9738,N_9233);
or U11318 (N_11318,N_5383,N_5147);
or U11319 (N_11319,N_8292,N_6194);
nor U11320 (N_11320,N_5652,N_5970);
nor U11321 (N_11321,N_8217,N_9995);
nand U11322 (N_11322,N_6311,N_9951);
nor U11323 (N_11323,N_8141,N_8989);
nand U11324 (N_11324,N_7726,N_5362);
nand U11325 (N_11325,N_5287,N_6709);
and U11326 (N_11326,N_8006,N_9886);
nor U11327 (N_11327,N_8366,N_5907);
nand U11328 (N_11328,N_9325,N_5216);
or U11329 (N_11329,N_5372,N_8667);
nor U11330 (N_11330,N_9432,N_5454);
nor U11331 (N_11331,N_8502,N_9005);
nand U11332 (N_11332,N_8896,N_7986);
nand U11333 (N_11333,N_9758,N_6733);
nand U11334 (N_11334,N_6724,N_6008);
nor U11335 (N_11335,N_9397,N_9808);
and U11336 (N_11336,N_7497,N_7208);
nor U11337 (N_11337,N_8565,N_5980);
and U11338 (N_11338,N_6340,N_8401);
or U11339 (N_11339,N_8473,N_8525);
nor U11340 (N_11340,N_7520,N_8225);
or U11341 (N_11341,N_6854,N_6296);
and U11342 (N_11342,N_8111,N_6095);
nand U11343 (N_11343,N_9583,N_7286);
or U11344 (N_11344,N_7068,N_7496);
and U11345 (N_11345,N_7035,N_5342);
nor U11346 (N_11346,N_7792,N_7642);
nor U11347 (N_11347,N_7438,N_7770);
and U11348 (N_11348,N_6387,N_9605);
and U11349 (N_11349,N_5179,N_9056);
nand U11350 (N_11350,N_7843,N_6282);
nor U11351 (N_11351,N_5325,N_7071);
or U11352 (N_11352,N_6648,N_7799);
nor U11353 (N_11353,N_6432,N_6752);
and U11354 (N_11354,N_5485,N_9652);
nor U11355 (N_11355,N_6092,N_6970);
nor U11356 (N_11356,N_5696,N_6902);
nand U11357 (N_11357,N_7013,N_9721);
or U11358 (N_11358,N_9250,N_7617);
and U11359 (N_11359,N_7387,N_8352);
nor U11360 (N_11360,N_7619,N_7424);
nor U11361 (N_11361,N_5719,N_5350);
and U11362 (N_11362,N_9243,N_9374);
or U11363 (N_11363,N_7756,N_6918);
and U11364 (N_11364,N_7040,N_6632);
xnor U11365 (N_11365,N_5188,N_6982);
nor U11366 (N_11366,N_8700,N_6148);
nand U11367 (N_11367,N_5918,N_9417);
nor U11368 (N_11368,N_6803,N_6143);
nand U11369 (N_11369,N_7247,N_7473);
or U11370 (N_11370,N_6420,N_8809);
nor U11371 (N_11371,N_8053,N_8814);
nor U11372 (N_11372,N_6400,N_6817);
nor U11373 (N_11373,N_8129,N_9701);
nor U11374 (N_11374,N_6110,N_9176);
nor U11375 (N_11375,N_6188,N_5347);
nor U11376 (N_11376,N_8840,N_6382);
nor U11377 (N_11377,N_5158,N_7981);
nor U11378 (N_11378,N_7027,N_6252);
nor U11379 (N_11379,N_9518,N_7862);
nor U11380 (N_11380,N_6796,N_7840);
and U11381 (N_11381,N_9946,N_8509);
or U11382 (N_11382,N_9501,N_5979);
nand U11383 (N_11383,N_6507,N_5021);
xor U11384 (N_11384,N_7550,N_5831);
nand U11385 (N_11385,N_6675,N_7155);
or U11386 (N_11386,N_5835,N_5723);
and U11387 (N_11387,N_5754,N_7344);
or U11388 (N_11388,N_8187,N_7660);
or U11389 (N_11389,N_7852,N_6620);
or U11390 (N_11390,N_8833,N_6305);
nand U11391 (N_11391,N_7759,N_6692);
nor U11392 (N_11392,N_7171,N_9632);
nor U11393 (N_11393,N_7500,N_8743);
nand U11394 (N_11394,N_8060,N_7260);
or U11395 (N_11395,N_6139,N_7240);
nand U11396 (N_11396,N_7825,N_6924);
or U11397 (N_11397,N_8058,N_8293);
nand U11398 (N_11398,N_9179,N_8074);
and U11399 (N_11399,N_7352,N_8304);
and U11400 (N_11400,N_5121,N_5500);
nand U11401 (N_11401,N_9644,N_8909);
xnor U11402 (N_11402,N_5214,N_8573);
nor U11403 (N_11403,N_5868,N_8634);
xnor U11404 (N_11404,N_6199,N_7404);
and U11405 (N_11405,N_8950,N_5457);
and U11406 (N_11406,N_9629,N_9431);
nand U11407 (N_11407,N_7375,N_9781);
nor U11408 (N_11408,N_8765,N_9222);
and U11409 (N_11409,N_9521,N_9495);
nand U11410 (N_11410,N_5580,N_6717);
and U11411 (N_11411,N_8665,N_5976);
and U11412 (N_11412,N_9871,N_5186);
or U11413 (N_11413,N_7457,N_7122);
nand U11414 (N_11414,N_5772,N_9702);
and U11415 (N_11415,N_6422,N_9926);
xnor U11416 (N_11416,N_6075,N_9911);
nand U11417 (N_11417,N_6867,N_8949);
nand U11418 (N_11418,N_9308,N_5490);
or U11419 (N_11419,N_5879,N_9704);
nand U11420 (N_11420,N_9840,N_9275);
xor U11421 (N_11421,N_9960,N_6618);
nand U11422 (N_11422,N_6279,N_5067);
or U11423 (N_11423,N_6176,N_6264);
or U11424 (N_11424,N_6833,N_5048);
nand U11425 (N_11425,N_5626,N_5094);
nand U11426 (N_11426,N_9276,N_6037);
and U11427 (N_11427,N_5745,N_9818);
nand U11428 (N_11428,N_8958,N_6402);
and U11429 (N_11429,N_7446,N_9720);
nand U11430 (N_11430,N_6688,N_8879);
nand U11431 (N_11431,N_6215,N_7962);
or U11432 (N_11432,N_9802,N_9322);
or U11433 (N_11433,N_6445,N_8955);
and U11434 (N_11434,N_6154,N_7958);
and U11435 (N_11435,N_8801,N_6581);
and U11436 (N_11436,N_8510,N_8862);
nand U11437 (N_11437,N_9170,N_8307);
nand U11438 (N_11438,N_8996,N_8874);
nor U11439 (N_11439,N_5586,N_5419);
nand U11440 (N_11440,N_6138,N_6872);
nor U11441 (N_11441,N_6028,N_6295);
nor U11442 (N_11442,N_9046,N_9331);
or U11443 (N_11443,N_8982,N_5124);
nand U11444 (N_11444,N_9387,N_9343);
and U11445 (N_11445,N_7915,N_8048);
or U11446 (N_11446,N_6221,N_7645);
or U11447 (N_11447,N_8655,N_9594);
nand U11448 (N_11448,N_9765,N_5853);
nand U11449 (N_11449,N_5533,N_9694);
nor U11450 (N_11450,N_5299,N_8181);
nand U11451 (N_11451,N_5514,N_5032);
or U11452 (N_11452,N_5517,N_7653);
or U11453 (N_11453,N_8895,N_9139);
nand U11454 (N_11454,N_8889,N_6166);
and U11455 (N_11455,N_8581,N_9349);
and U11456 (N_11456,N_9124,N_7080);
nand U11457 (N_11457,N_8290,N_5079);
nand U11458 (N_11458,N_5162,N_6491);
nor U11459 (N_11459,N_7501,N_8067);
nor U11460 (N_11460,N_5982,N_5435);
nor U11461 (N_11461,N_5583,N_7906);
nor U11462 (N_11462,N_8302,N_6897);
or U11463 (N_11463,N_5591,N_5410);
or U11464 (N_11464,N_6594,N_7527);
nand U11465 (N_11465,N_6338,N_7596);
or U11466 (N_11466,N_5655,N_7477);
nor U11467 (N_11467,N_6304,N_7801);
or U11468 (N_11468,N_8922,N_7669);
or U11469 (N_11469,N_8971,N_8745);
or U11470 (N_11470,N_6568,N_9463);
nand U11471 (N_11471,N_8101,N_5215);
xor U11472 (N_11472,N_9973,N_9122);
nand U11473 (N_11473,N_7955,N_5371);
nand U11474 (N_11474,N_6197,N_9870);
nand U11475 (N_11475,N_9344,N_6856);
and U11476 (N_11476,N_5711,N_5482);
and U11477 (N_11477,N_6781,N_9741);
and U11478 (N_11478,N_9497,N_7074);
and U11479 (N_11479,N_6434,N_5613);
xor U11480 (N_11480,N_7874,N_9966);
nand U11481 (N_11481,N_6335,N_9657);
nor U11482 (N_11482,N_7939,N_6654);
or U11483 (N_11483,N_9982,N_9997);
or U11484 (N_11484,N_6464,N_6084);
or U11485 (N_11485,N_6676,N_8935);
nor U11486 (N_11486,N_8695,N_9089);
nor U11487 (N_11487,N_9595,N_5224);
nor U11488 (N_11488,N_7270,N_5249);
or U11489 (N_11489,N_6864,N_8520);
or U11490 (N_11490,N_7149,N_7644);
nand U11491 (N_11491,N_8702,N_7416);
and U11492 (N_11492,N_9679,N_6349);
and U11493 (N_11493,N_6925,N_5938);
and U11494 (N_11494,N_9947,N_6520);
nand U11495 (N_11495,N_5085,N_6561);
nand U11496 (N_11496,N_6892,N_9538);
or U11497 (N_11497,N_5948,N_7965);
and U11498 (N_11498,N_7196,N_6740);
nor U11499 (N_11499,N_8926,N_7172);
or U11500 (N_11500,N_9378,N_6884);
nand U11501 (N_11501,N_5319,N_5058);
and U11502 (N_11502,N_7600,N_6354);
nor U11503 (N_11503,N_8534,N_8428);
or U11504 (N_11504,N_9925,N_7761);
nor U11505 (N_11505,N_9433,N_7341);
nor U11506 (N_11506,N_6636,N_9777);
or U11507 (N_11507,N_9892,N_7221);
nand U11508 (N_11508,N_9182,N_7641);
nor U11509 (N_11509,N_9934,N_9526);
nor U11510 (N_11510,N_8465,N_5952);
or U11511 (N_11511,N_9885,N_7817);
nand U11512 (N_11512,N_9253,N_9687);
nor U11513 (N_11513,N_6904,N_5553);
or U11514 (N_11514,N_8933,N_7696);
or U11515 (N_11515,N_8267,N_9747);
or U11516 (N_11516,N_8138,N_8114);
nor U11517 (N_11517,N_5884,N_7372);
and U11518 (N_11518,N_7864,N_6773);
nand U11519 (N_11519,N_5050,N_6896);
and U11520 (N_11520,N_8673,N_9134);
and U11521 (N_11521,N_7599,N_5111);
or U11522 (N_11522,N_9004,N_9033);
and U11523 (N_11523,N_9030,N_7284);
nor U11524 (N_11524,N_5731,N_6711);
nor U11525 (N_11525,N_8285,N_5666);
nand U11526 (N_11526,N_5738,N_5782);
nand U11527 (N_11527,N_8226,N_6526);
and U11528 (N_11528,N_5014,N_6160);
and U11529 (N_11529,N_6001,N_5991);
nand U11530 (N_11530,N_8142,N_5031);
nand U11531 (N_11531,N_8231,N_5783);
or U11532 (N_11532,N_5093,N_8314);
and U11533 (N_11533,N_5260,N_7950);
or U11534 (N_11534,N_6742,N_5592);
or U11535 (N_11535,N_8815,N_6844);
nor U11536 (N_11536,N_8881,N_6805);
and U11537 (N_11537,N_6801,N_6555);
or U11538 (N_11538,N_8259,N_8604);
nor U11539 (N_11539,N_5373,N_5598);
or U11540 (N_11540,N_7315,N_7841);
nand U11541 (N_11541,N_9006,N_9461);
or U11542 (N_11542,N_5615,N_6050);
and U11543 (N_11543,N_8298,N_9924);
nand U11544 (N_11544,N_8995,N_8560);
and U11545 (N_11545,N_7355,N_6316);
or U11546 (N_11546,N_6627,N_6040);
and U11547 (N_11547,N_7984,N_5462);
and U11548 (N_11548,N_6797,N_6228);
xnor U11549 (N_11549,N_8414,N_9142);
and U11550 (N_11550,N_5061,N_9616);
nor U11551 (N_11551,N_7430,N_8662);
nor U11552 (N_11552,N_7639,N_6905);
or U11553 (N_11553,N_8870,N_5669);
and U11554 (N_11554,N_7789,N_7829);
or U11555 (N_11555,N_5178,N_8311);
or U11556 (N_11556,N_6680,N_7631);
or U11557 (N_11557,N_6249,N_8021);
or U11558 (N_11558,N_6649,N_5925);
nand U11559 (N_11559,N_7751,N_8027);
or U11560 (N_11560,N_5687,N_5089);
or U11561 (N_11561,N_7657,N_9626);
or U11562 (N_11562,N_9627,N_9964);
nor U11563 (N_11563,N_5690,N_5911);
or U11564 (N_11564,N_6119,N_5100);
or U11565 (N_11565,N_7483,N_7005);
nand U11566 (N_11566,N_5381,N_9868);
and U11567 (N_11567,N_9103,N_7179);
nor U11568 (N_11568,N_8107,N_6512);
and U11569 (N_11569,N_9570,N_6934);
or U11570 (N_11570,N_6839,N_5264);
nor U11571 (N_11571,N_5460,N_6153);
and U11572 (N_11572,N_9426,N_8856);
nor U11573 (N_11573,N_7615,N_8015);
nand U11574 (N_11574,N_8610,N_7239);
and U11575 (N_11575,N_7287,N_7162);
xor U11576 (N_11576,N_7243,N_6152);
nor U11577 (N_11577,N_7538,N_9618);
and U11578 (N_11578,N_5217,N_5339);
or U11579 (N_11579,N_8014,N_7409);
nor U11580 (N_11580,N_7580,N_7611);
nor U11581 (N_11581,N_5550,N_6278);
and U11582 (N_11582,N_9893,N_7742);
nor U11583 (N_11583,N_6829,N_6186);
nor U11584 (N_11584,N_8214,N_5286);
nor U11585 (N_11585,N_8830,N_7126);
nor U11586 (N_11586,N_6735,N_8694);
and U11587 (N_11587,N_7140,N_6783);
nand U11588 (N_11588,N_7588,N_9297);
nor U11589 (N_11589,N_9575,N_7268);
nor U11590 (N_11590,N_5001,N_6661);
nor U11591 (N_11591,N_9091,N_9479);
or U11592 (N_11592,N_8620,N_9286);
and U11593 (N_11593,N_8592,N_8270);
nand U11594 (N_11594,N_8047,N_9710);
or U11595 (N_11595,N_8446,N_5202);
and U11596 (N_11596,N_5971,N_7428);
and U11597 (N_11597,N_9700,N_7999);
nor U11598 (N_11598,N_7124,N_7299);
or U11599 (N_11599,N_5328,N_7178);
or U11600 (N_11600,N_9341,N_7658);
nor U11601 (N_11601,N_6766,N_5049);
nand U11602 (N_11602,N_5664,N_6687);
nor U11603 (N_11603,N_6204,N_9532);
and U11604 (N_11604,N_9743,N_9874);
nand U11605 (N_11605,N_8463,N_7045);
nand U11606 (N_11606,N_7295,N_9956);
nand U11607 (N_11607,N_9833,N_9280);
or U11608 (N_11608,N_6917,N_5920);
nor U11609 (N_11609,N_5293,N_9472);
or U11610 (N_11610,N_9608,N_5678);
nand U11611 (N_11611,N_9955,N_7735);
and U11612 (N_11612,N_7996,N_6207);
or U11613 (N_11613,N_8648,N_9488);
nor U11614 (N_11614,N_5841,N_7277);
nor U11615 (N_11615,N_5390,N_7821);
and U11616 (N_11616,N_7435,N_6219);
or U11617 (N_11617,N_8767,N_6993);
and U11618 (N_11618,N_6519,N_8197);
nor U11619 (N_11619,N_8925,N_9854);
nand U11620 (N_11620,N_5679,N_7278);
nor U11621 (N_11621,N_5070,N_7959);
nor U11622 (N_11622,N_8679,N_9661);
or U11623 (N_11623,N_8701,N_5800);
and U11624 (N_11624,N_5939,N_9971);
and U11625 (N_11625,N_8408,N_9624);
nor U11626 (N_11626,N_7647,N_6972);
or U11627 (N_11627,N_7364,N_5775);
nor U11628 (N_11628,N_7917,N_9153);
or U11629 (N_11629,N_6941,N_5631);
nand U11630 (N_11630,N_5677,N_5794);
nand U11631 (N_11631,N_5878,N_8952);
nor U11632 (N_11632,N_8892,N_5818);
nand U11633 (N_11633,N_9466,N_7776);
or U11634 (N_11634,N_7281,N_7076);
nand U11635 (N_11635,N_8458,N_5537);
or U11636 (N_11636,N_7121,N_5361);
or U11637 (N_11637,N_7332,N_5899);
and U11638 (N_11638,N_5366,N_6388);
nand U11639 (N_11639,N_9985,N_6855);
nand U11640 (N_11640,N_5267,N_8898);
or U11641 (N_11641,N_6178,N_5175);
nand U11642 (N_11642,N_8454,N_8140);
or U11643 (N_11643,N_9420,N_6843);
or U11644 (N_11644,N_6708,N_7914);
and U11645 (N_11645,N_9442,N_9883);
or U11646 (N_11646,N_6460,N_7522);
nor U11647 (N_11647,N_9839,N_5375);
and U11648 (N_11648,N_8456,N_8396);
nand U11649 (N_11649,N_9520,N_9069);
or U11650 (N_11650,N_9448,N_8812);
or U11651 (N_11651,N_7794,N_5817);
nor U11652 (N_11652,N_6705,N_8790);
or U11653 (N_11653,N_6963,N_8983);
and U11654 (N_11654,N_8538,N_9514);
and U11655 (N_11655,N_5183,N_9942);
nor U11656 (N_11656,N_5388,N_7158);
nand U11657 (N_11657,N_6488,N_8448);
nand U11658 (N_11658,N_5607,N_8439);
nand U11659 (N_11659,N_5207,N_8584);
and U11660 (N_11660,N_8119,N_5341);
nor U11661 (N_11661,N_8650,N_6108);
nand U11662 (N_11662,N_6405,N_8990);
and U11663 (N_11663,N_8918,N_9024);
nand U11664 (N_11664,N_5873,N_9468);
nor U11665 (N_11665,N_6071,N_6540);
nor U11666 (N_11666,N_7282,N_8248);
nor U11667 (N_11667,N_6326,N_8633);
nand U11668 (N_11668,N_6007,N_8736);
xor U11669 (N_11669,N_5386,N_8110);
and U11670 (N_11670,N_9906,N_6156);
nand U11671 (N_11671,N_6477,N_7937);
nand U11672 (N_11672,N_8546,N_8698);
nand U11673 (N_11673,N_8347,N_7492);
or U11674 (N_11674,N_6378,N_5280);
nand U11675 (N_11675,N_8683,N_6451);
nand U11676 (N_11676,N_7725,N_8561);
nand U11677 (N_11677,N_7839,N_9327);
or U11678 (N_11678,N_5323,N_9506);
nor U11679 (N_11679,N_9566,N_7618);
and U11680 (N_11680,N_9492,N_9231);
or U11681 (N_11681,N_7671,N_9312);
nand U11682 (N_11682,N_7758,N_9932);
and U11683 (N_11683,N_6310,N_6572);
or U11684 (N_11684,N_9933,N_8613);
or U11685 (N_11685,N_7440,N_7643);
or U11686 (N_11686,N_8964,N_6355);
nand U11687 (N_11687,N_7060,N_8945);
xor U11688 (N_11688,N_6391,N_6371);
nor U11689 (N_11689,N_5367,N_5953);
nand U11690 (N_11690,N_9404,N_5589);
and U11691 (N_11691,N_5394,N_9952);
nand U11692 (N_11692,N_7096,N_5171);
and U11693 (N_11693,N_7860,N_9237);
nand U11694 (N_11694,N_8643,N_6398);
nor U11695 (N_11695,N_7039,N_9527);
or U11696 (N_11696,N_9978,N_8093);
or U11697 (N_11697,N_7741,N_6660);
and U11698 (N_11698,N_9815,N_5896);
or U11699 (N_11699,N_6214,N_5131);
or U11700 (N_11700,N_6899,N_9196);
or U11701 (N_11701,N_5762,N_7668);
and U11702 (N_11702,N_9265,N_8472);
and U11703 (N_11703,N_6163,N_9786);
nand U11704 (N_11704,N_5106,N_8689);
and U11705 (N_11705,N_6126,N_9568);
or U11706 (N_11706,N_7717,N_5357);
nand U11707 (N_11707,N_9658,N_8349);
nor U11708 (N_11708,N_8243,N_8611);
and U11709 (N_11709,N_8273,N_7774);
nor U11710 (N_11710,N_6536,N_9576);
or U11711 (N_11711,N_6966,N_8975);
nor U11712 (N_11712,N_9762,N_8588);
or U11713 (N_11713,N_5704,N_7279);
xor U11714 (N_11714,N_6466,N_8381);
nand U11715 (N_11715,N_6297,N_6058);
or U11716 (N_11716,N_9388,N_7441);
nand U11717 (N_11717,N_7145,N_6352);
and U11718 (N_11718,N_5279,N_9641);
nand U11719 (N_11719,N_5025,N_6588);
nor U11720 (N_11720,N_6447,N_8869);
nor U11721 (N_11721,N_6270,N_6903);
nor U11722 (N_11722,N_8866,N_9974);
nand U11723 (N_11723,N_6563,N_6063);
or U11724 (N_11724,N_5798,N_5204);
nor U11725 (N_11725,N_5984,N_9370);
nand U11726 (N_11726,N_7871,N_9776);
or U11727 (N_11727,N_8635,N_5143);
or U11728 (N_11728,N_5880,N_7935);
or U11729 (N_11729,N_7164,N_5322);
nand U11730 (N_11730,N_7837,N_9230);
nand U11731 (N_11731,N_5673,N_8970);
nor U11732 (N_11732,N_9051,N_9486);
nor U11733 (N_11733,N_7524,N_6325);
or U11734 (N_11734,N_5511,N_6768);
or U11735 (N_11735,N_5487,N_6074);
nand U11736 (N_11736,N_7363,N_6644);
nor U11737 (N_11737,N_8134,N_5023);
and U11738 (N_11738,N_9667,N_5892);
nand U11739 (N_11739,N_7757,N_8385);
nand U11740 (N_11740,N_6922,N_8265);
nand U11741 (N_11741,N_6004,N_6113);
or U11742 (N_11742,N_8391,N_6564);
nor U11743 (N_11743,N_7302,N_9740);
and U11744 (N_11744,N_8859,N_9796);
or U11745 (N_11745,N_7183,N_5272);
and U11746 (N_11746,N_6535,N_5577);
xnor U11747 (N_11747,N_9311,N_6168);
or U11748 (N_11748,N_9140,N_9949);
and U11749 (N_11749,N_6384,N_6971);
nor U11750 (N_11750,N_6786,N_6700);
and U11751 (N_11751,N_5532,N_8350);
and U11752 (N_11752,N_7218,N_9869);
or U11753 (N_11753,N_5223,N_7790);
nor U11754 (N_11754,N_6614,N_5632);
and U11755 (N_11755,N_9181,N_5039);
or U11756 (N_11756,N_9509,N_8419);
and U11757 (N_11757,N_9229,N_8602);
or U11758 (N_11758,N_9175,N_6283);
xnor U11759 (N_11759,N_6425,N_7159);
or U11760 (N_11760,N_8159,N_5173);
nand U11761 (N_11761,N_6701,N_9376);
or U11762 (N_11762,N_9968,N_9718);
or U11763 (N_11763,N_7151,N_8606);
nor U11764 (N_11764,N_8763,N_8013);
nor U11765 (N_11765,N_9053,N_7084);
and U11766 (N_11766,N_9975,N_9453);
and U11767 (N_11767,N_9131,N_9950);
nor U11768 (N_11768,N_7399,N_9289);
or U11769 (N_11769,N_5122,N_9197);
or U11770 (N_11770,N_5035,N_8039);
nand U11771 (N_11771,N_9556,N_6147);
nor U11772 (N_11772,N_8758,N_8205);
and U11773 (N_11773,N_8753,N_7932);
nand U11774 (N_11774,N_5670,N_6467);
nand U11775 (N_11775,N_9988,N_6368);
nor U11776 (N_11776,N_7678,N_5258);
or U11777 (N_11777,N_8624,N_7880);
nand U11778 (N_11778,N_7977,N_8219);
nor U11779 (N_11779,N_8294,N_7707);
nor U11780 (N_11780,N_9563,N_5230);
nand U11781 (N_11781,N_8164,N_6217);
and U11782 (N_11782,N_5638,N_6655);
and U11783 (N_11783,N_7674,N_8375);
or U11784 (N_11784,N_8320,N_8550);
nor U11785 (N_11785,N_6615,N_5095);
and U11786 (N_11786,N_9750,N_9359);
or U11787 (N_11787,N_5195,N_8532);
xor U11788 (N_11788,N_5519,N_5433);
or U11789 (N_11789,N_8440,N_8081);
nand U11790 (N_11790,N_7242,N_8459);
or U11791 (N_11791,N_9415,N_6851);
or U11792 (N_11792,N_9977,N_6990);
nor U11793 (N_11793,N_5787,N_6140);
or U11794 (N_11794,N_7941,N_6081);
nand U11795 (N_11795,N_8723,N_7023);
nand U11796 (N_11796,N_7479,N_7193);
and U11797 (N_11797,N_9087,N_8322);
nor U11798 (N_11798,N_7485,N_9379);
nand U11799 (N_11799,N_7969,N_8976);
nor U11800 (N_11800,N_8295,N_8151);
or U11801 (N_11801,N_5784,N_5809);
or U11802 (N_11802,N_6710,N_6253);
or U11803 (N_11803,N_5295,N_6137);
and U11804 (N_11804,N_7990,N_9770);
and U11805 (N_11805,N_9493,N_8657);
nor U11806 (N_11806,N_7050,N_5210);
nor U11807 (N_11807,N_5177,N_7093);
nor U11808 (N_11808,N_8240,N_9876);
nand U11809 (N_11809,N_6122,N_9788);
and U11810 (N_11810,N_8034,N_9025);
nand U11811 (N_11811,N_8644,N_8608);
xnor U11812 (N_11812,N_7782,N_7410);
or U11813 (N_11813,N_6380,N_6737);
nor U11814 (N_11814,N_8951,N_9126);
or U11815 (N_11815,N_6589,N_7360);
nand U11816 (N_11816,N_5741,N_5967);
and U11817 (N_11817,N_9803,N_7082);
and U11818 (N_11818,N_5450,N_7454);
or U11819 (N_11819,N_5213,N_6164);
nand U11820 (N_11820,N_6484,N_7802);
or U11821 (N_11821,N_8605,N_7021);
nor U11822 (N_11822,N_9009,N_8028);
and U11823 (N_11823,N_8035,N_5647);
and U11824 (N_11824,N_9301,N_5516);
nand U11825 (N_11825,N_5180,N_8825);
nand U11826 (N_11826,N_9755,N_5501);
nand U11827 (N_11827,N_8136,N_6837);
nor U11828 (N_11828,N_7088,N_8928);
nor U11829 (N_11829,N_7346,N_9285);
nor U11830 (N_11830,N_6052,N_6957);
nor U11831 (N_11831,N_8791,N_6608);
and U11832 (N_11832,N_6628,N_7238);
nand U11833 (N_11833,N_8914,N_5943);
and U11834 (N_11834,N_8370,N_9402);
nand U11835 (N_11835,N_8808,N_6281);
or U11836 (N_11836,N_6177,N_7055);
nand U11837 (N_11837,N_7338,N_6288);
or U11838 (N_11838,N_6053,N_9983);
nor U11839 (N_11839,N_8341,N_8692);
or U11840 (N_11840,N_7261,N_5036);
or U11841 (N_11841,N_9171,N_5658);
nand U11842 (N_11842,N_5203,N_6327);
or U11843 (N_11843,N_9723,N_6141);
and U11844 (N_11844,N_6225,N_5439);
nor U11845 (N_11845,N_9999,N_9095);
nand U11846 (N_11846,N_9345,N_6345);
or U11847 (N_11847,N_6547,N_7878);
nor U11848 (N_11848,N_6665,N_8204);
or U11849 (N_11849,N_8424,N_6532);
and U11850 (N_11850,N_7331,N_9211);
xnor U11851 (N_11851,N_6097,N_5421);
nand U11852 (N_11852,N_5618,N_5887);
or U11853 (N_11853,N_5426,N_7814);
or U11854 (N_11854,N_9752,N_7384);
nor U11855 (N_11855,N_8239,N_6083);
and U11856 (N_11856,N_7493,N_9398);
and U11857 (N_11857,N_7654,N_9663);
or U11858 (N_11858,N_5930,N_6482);
or U11859 (N_11859,N_8954,N_5427);
nand U11860 (N_11860,N_7948,N_6693);
nor U11861 (N_11861,N_5646,N_6048);
nand U11862 (N_11862,N_9623,N_7894);
nor U11863 (N_11863,N_6005,N_6487);
or U11864 (N_11864,N_6863,N_7997);
xor U11865 (N_11865,N_8324,N_8521);
and U11866 (N_11866,N_5941,N_6465);
xnor U11867 (N_11867,N_7275,N_7194);
or U11868 (N_11868,N_9920,N_8064);
nand U11869 (N_11869,N_9611,N_9860);
or U11870 (N_11870,N_5949,N_9210);
nor U11871 (N_11871,N_9059,N_5758);
and U11872 (N_11872,N_7046,N_9137);
nand U11873 (N_11873,N_5016,N_5974);
and U11874 (N_11874,N_7540,N_9380);
nor U11875 (N_11875,N_8451,N_5420);
and U11876 (N_11876,N_6049,N_8480);
or U11877 (N_11877,N_5397,N_5559);
nor U11878 (N_11878,N_8339,N_7067);
nor U11879 (N_11879,N_5329,N_8817);
nor U11880 (N_11880,N_9692,N_7530);
and U11881 (N_11881,N_8593,N_7679);
or U11882 (N_11882,N_6911,N_5992);
xnor U11883 (N_11883,N_6427,N_7117);
nor U11884 (N_11884,N_5986,N_5379);
and U11885 (N_11885,N_7523,N_6931);
nand U11886 (N_11886,N_8080,N_8109);
or U11887 (N_11887,N_9184,N_7198);
and U11888 (N_11888,N_8466,N_9219);
nor U11889 (N_11889,N_9454,N_5163);
nor U11890 (N_11890,N_8363,N_7766);
and U11891 (N_11891,N_7383,N_9072);
and U11892 (N_11892,N_9274,N_6546);
xnor U11893 (N_11893,N_8321,N_6124);
nand U11894 (N_11894,N_6590,N_9756);
or U11895 (N_11895,N_7966,N_7952);
nor U11896 (N_11896,N_6091,N_7397);
nor U11897 (N_11897,N_9227,N_7373);
nand U11898 (N_11898,N_9604,N_8272);
or U11899 (N_11899,N_6101,N_8180);
nand U11900 (N_11900,N_9560,N_8716);
and U11901 (N_11901,N_5812,N_8077);
nor U11902 (N_11902,N_6193,N_5902);
or U11903 (N_11903,N_8069,N_7142);
and U11904 (N_11904,N_5422,N_6553);
or U11905 (N_11905,N_6698,N_6511);
nor U11906 (N_11906,N_5404,N_9482);
or U11907 (N_11907,N_6828,N_5635);
nor U11908 (N_11908,N_6877,N_7665);
nand U11909 (N_11909,N_8490,N_7051);
and U11910 (N_11910,N_7231,N_9639);
and U11911 (N_11911,N_5096,N_6992);
and U11912 (N_11912,N_7800,N_5850);
or U11913 (N_11913,N_5538,N_9646);
nor U11914 (N_11914,N_6396,N_8877);
nor U11915 (N_11915,N_5228,N_8286);
nand U11916 (N_11916,N_6556,N_7403);
and U11917 (N_11917,N_6566,N_9957);
nand U11918 (N_11918,N_9355,N_8903);
or U11919 (N_11919,N_7148,N_6574);
nor U11920 (N_11920,N_9264,N_6689);
or U11921 (N_11921,N_8651,N_5278);
or U11922 (N_11922,N_7398,N_6361);
or U11923 (N_11923,N_5484,N_7153);
and U11924 (N_11924,N_7453,N_7586);
nor U11925 (N_11925,N_7834,N_5027);
and U11926 (N_11926,N_5661,N_6210);
or U11927 (N_11927,N_5761,N_7503);
nand U11928 (N_11928,N_7748,N_7028);
nor U11929 (N_11929,N_9698,N_9199);
nor U11930 (N_11930,N_5345,N_6313);
or U11931 (N_11931,N_9007,N_9373);
or U11932 (N_11932,N_9141,N_9055);
nor U11933 (N_11933,N_6149,N_8696);
nor U11934 (N_11934,N_9474,N_5959);
nand U11935 (N_11935,N_5130,N_6453);
and U11936 (N_11936,N_9536,N_8118);
nand U11937 (N_11937,N_6232,N_5963);
and U11938 (N_11938,N_9026,N_5846);
nor U11939 (N_11939,N_8599,N_9180);
nor U11940 (N_11940,N_6778,N_6408);
nand U11941 (N_11941,N_8103,N_9827);
nand U11942 (N_11942,N_7053,N_5700);
or U11943 (N_11943,N_7737,N_5950);
nand U11944 (N_11944,N_6131,N_9003);
nand U11945 (N_11945,N_9235,N_7701);
nor U11946 (N_11946,N_6557,N_9668);
or U11947 (N_11947,N_6515,N_8191);
and U11948 (N_11948,N_7165,N_7089);
or U11949 (N_11949,N_8332,N_5123);
nor U11950 (N_11950,N_8867,N_9459);
nor U11951 (N_11951,N_8338,N_7318);
nand U11952 (N_11952,N_7655,N_8260);
and U11953 (N_11953,N_9365,N_5588);
nand U11954 (N_11954,N_6286,N_5505);
or U11955 (N_11955,N_5190,N_6827);
nor U11956 (N_11956,N_6956,N_5221);
nand U11957 (N_11957,N_8372,N_5888);
or U11958 (N_11958,N_5662,N_8403);
xnor U11959 (N_11959,N_9909,N_6261);
nor U11960 (N_11960,N_6509,N_7339);
nor U11961 (N_11961,N_7830,N_9912);
nand U11962 (N_11962,N_8315,N_9455);
and U11963 (N_11963,N_8713,N_6159);
and U11964 (N_11964,N_6923,N_8623);
and U11965 (N_11965,N_8232,N_7016);
or U11966 (N_11966,N_8336,N_6996);
nor U11967 (N_11967,N_7471,N_8905);
or U11968 (N_11968,N_9207,N_6718);
and U11969 (N_11969,N_8377,N_8445);
and U11970 (N_11970,N_6549,N_6826);
nand U11971 (N_11971,N_9202,N_7425);
or U11972 (N_11972,N_9546,N_7882);
or U11973 (N_11973,N_9236,N_8769);
nand U11974 (N_11974,N_7743,N_5703);
nor U11975 (N_11975,N_8145,N_5942);
nand U11976 (N_11976,N_5870,N_8571);
or U11977 (N_11977,N_9719,N_7716);
or U11978 (N_11978,N_6262,N_7913);
nor U11979 (N_11979,N_8112,N_6542);
and U11980 (N_11980,N_6591,N_7010);
and U11981 (N_11981,N_6815,N_6243);
and U11982 (N_11982,N_6364,N_8125);
or U11983 (N_11983,N_6550,N_7417);
nor U11984 (N_11984,N_6406,N_9050);
or U11985 (N_11985,N_7715,N_8508);
and U11986 (N_11986,N_5349,N_6497);
and U11987 (N_11987,N_6185,N_9863);
nand U11988 (N_11988,N_8484,N_8411);
or U11989 (N_11989,N_5657,N_9784);
nand U11990 (N_11990,N_8212,N_5292);
and U11991 (N_11991,N_8279,N_5814);
nand U11992 (N_11992,N_8727,N_8227);
and U11993 (N_11993,N_7777,N_9515);
nand U11994 (N_11994,N_6788,N_8261);
nand U11995 (N_11995,N_7575,N_8748);
and U11996 (N_11996,N_7135,N_5448);
nand U11997 (N_11997,N_8930,N_6073);
xor U11998 (N_11998,N_7565,N_7891);
nand U11999 (N_11999,N_8115,N_9552);
and U12000 (N_12000,N_8547,N_7987);
nor U12001 (N_12001,N_6183,N_7967);
or U12002 (N_12002,N_6677,N_6055);
nor U12003 (N_12003,N_8685,N_5797);
and U12004 (N_12004,N_5489,N_9587);
or U12005 (N_12005,N_6227,N_7380);
and U12006 (N_12006,N_5493,N_8312);
nand U12007 (N_12007,N_6006,N_7640);
or U12008 (N_12008,N_6777,N_8030);
nand U12009 (N_12009,N_5496,N_7805);
nor U12010 (N_12010,N_9149,N_6603);
nor U12011 (N_12011,N_6707,N_6011);
or U12012 (N_12012,N_7017,N_5913);
or U12013 (N_12013,N_7836,N_6691);
or U12014 (N_12014,N_7241,N_9917);
and U12015 (N_12015,N_5407,N_6303);
nand U12016 (N_12016,N_5954,N_7689);
or U12017 (N_12017,N_5684,N_6211);
nand U12018 (N_12018,N_5912,N_8762);
nor U12019 (N_12019,N_9760,N_9045);
nand U12020 (N_12020,N_6640,N_9392);
and U12021 (N_12021,N_9675,N_7223);
nand U12022 (N_12022,N_7769,N_5065);
and U12023 (N_12023,N_6293,N_6067);
or U12024 (N_12024,N_8234,N_8669);
xor U12025 (N_12025,N_6804,N_7173);
and U12026 (N_12026,N_9414,N_8780);
nor U12027 (N_12027,N_6912,N_7507);
nand U12028 (N_12028,N_9346,N_5431);
or U12029 (N_12029,N_6870,N_7254);
nor U12030 (N_12030,N_5254,N_6989);
nor U12031 (N_12031,N_9307,N_9935);
nor U12032 (N_12032,N_6191,N_7730);
and U12033 (N_12033,N_8420,N_8367);
and U12034 (N_12034,N_9992,N_6946);
nand U12035 (N_12035,N_8899,N_5528);
nor U12036 (N_12036,N_8656,N_7926);
or U12037 (N_12037,N_8676,N_5548);
nand U12038 (N_12038,N_6223,N_5303);
and U12039 (N_12039,N_6890,N_6876);
nor U12040 (N_12040,N_7686,N_6869);
nand U12041 (N_12041,N_6169,N_7448);
nor U12042 (N_12042,N_8397,N_6685);
and U12043 (N_12043,N_6853,N_5019);
or U12044 (N_12044,N_8942,N_6259);
nand U12045 (N_12045,N_5951,N_7401);
or U12046 (N_12046,N_9764,N_7212);
and U12047 (N_12047,N_7057,N_6780);
nor U12048 (N_12048,N_6118,N_8668);
nor U12049 (N_12049,N_7298,N_9550);
nand U12050 (N_12050,N_8042,N_9651);
and U12051 (N_12051,N_6308,N_9703);
or U12052 (N_12052,N_7784,N_9244);
or U12053 (N_12053,N_7083,N_8494);
and U12054 (N_12054,N_5785,N_6034);
nand U12055 (N_12055,N_9670,N_9313);
nor U12056 (N_12056,N_9247,N_8744);
and U12057 (N_12057,N_5889,N_5401);
or U12058 (N_12058,N_7824,N_8415);
nand U12059 (N_12059,N_8826,N_8255);
nor U12060 (N_12060,N_7285,N_5307);
nor U12061 (N_12061,N_7983,N_5681);
and U12062 (N_12062,N_9147,N_6492);
nand U12063 (N_12063,N_8803,N_6745);
nor U12064 (N_12064,N_8582,N_6377);
or U12065 (N_12065,N_9809,N_7123);
or U12066 (N_12066,N_6344,N_9688);
nor U12067 (N_12067,N_9135,N_7897);
and U12068 (N_12068,N_6389,N_9391);
nor U12069 (N_12069,N_8902,N_6024);
or U12070 (N_12070,N_9377,N_6082);
or U12071 (N_12071,N_9347,N_5695);
and U12072 (N_12072,N_6945,N_7077);
and U12073 (N_12073,N_9178,N_7582);
or U12074 (N_12074,N_6517,N_9801);
and U12075 (N_12075,N_8831,N_6552);
nand U12076 (N_12076,N_5502,N_6584);
nor U12077 (N_12077,N_7826,N_7141);
or U12078 (N_12078,N_9060,N_7526);
nor U12079 (N_12079,N_8224,N_7272);
nand U12080 (N_12080,N_6421,N_5139);
and U12081 (N_12081,N_6662,N_7516);
or U12082 (N_12082,N_8398,N_8849);
nor U12083 (N_12083,N_9154,N_5946);
nand U12084 (N_12084,N_5692,N_8326);
or U12085 (N_12085,N_8416,N_6988);
and U12086 (N_12086,N_9261,N_6162);
nor U12087 (N_12087,N_9356,N_8282);
and U12088 (N_12088,N_6158,N_9094);
nor U12089 (N_12089,N_6334,N_8999);
and U12090 (N_12090,N_9533,N_9148);
or U12091 (N_12091,N_7723,N_9938);
nand U12092 (N_12092,N_7589,N_6392);
nand U12093 (N_12093,N_9525,N_6260);
and U12094 (N_12094,N_9714,N_8244);
nor U12095 (N_12095,N_9865,N_7163);
nand U12096 (N_12096,N_8703,N_6651);
nand U12097 (N_12097,N_7783,N_5266);
nand U12098 (N_12098,N_5443,N_7118);
or U12099 (N_12099,N_8779,N_7888);
nor U12100 (N_12100,N_7130,N_9019);
nor U12101 (N_12101,N_9281,N_9769);
nor U12102 (N_12102,N_7594,N_5041);
or U12103 (N_12103,N_5211,N_7633);
and U12104 (N_12104,N_7283,N_6744);
xor U12105 (N_12105,N_5587,N_8220);
and U12106 (N_12106,N_9369,N_8433);
and U12107 (N_12107,N_5446,N_8016);
nor U12108 (N_12108,N_7866,N_6883);
and U12109 (N_12109,N_8962,N_7512);
nand U12110 (N_12110,N_8437,N_5737);
nor U12111 (N_12111,N_5452,N_7014);
or U12112 (N_12112,N_8737,N_9907);
nand U12113 (N_12113,N_6793,N_7680);
nand U12114 (N_12114,N_9607,N_6441);
nor U12115 (N_12115,N_8104,N_8595);
and U12116 (N_12116,N_8082,N_7745);
nor U12117 (N_12117,N_7635,N_6570);
nand U12118 (N_12118,N_7625,N_9767);
and U12119 (N_12119,N_5989,N_5562);
nand U12120 (N_12120,N_8450,N_9547);
nand U12121 (N_12121,N_8802,N_8018);
or U12122 (N_12122,N_5601,N_9810);
nand U12123 (N_12123,N_9653,N_7258);
nand U12124 (N_12124,N_5235,N_9828);
nand U12125 (N_12125,N_7994,N_9085);
nand U12126 (N_12126,N_5867,N_9881);
nand U12127 (N_12127,N_5109,N_5161);
and U12128 (N_12128,N_8083,N_8647);
or U12129 (N_12129,N_5309,N_8500);
nor U12130 (N_12130,N_6643,N_5855);
or U12131 (N_12131,N_9464,N_7771);
nor U12132 (N_12132,N_6157,N_9299);
and U12133 (N_12133,N_9097,N_7779);
and U12134 (N_12134,N_6501,N_7317);
and U12135 (N_12135,N_9729,N_6418);
xor U12136 (N_12136,N_9631,N_7623);
nand U12137 (N_12137,N_6373,N_7174);
nor U12138 (N_12138,N_8144,N_8150);
nor U12139 (N_12139,N_9994,N_5840);
nor U12140 (N_12140,N_8049,N_5639);
xor U12141 (N_12141,N_6514,N_9043);
nor U12142 (N_12142,N_9284,N_9543);
nor U12143 (N_12143,N_9119,N_6967);
or U12144 (N_12144,N_5308,N_6247);
and U12145 (N_12145,N_8182,N_9716);
or U12146 (N_12146,N_5145,N_7812);
nor U12147 (N_12147,N_8245,N_5910);
nand U12148 (N_12148,N_6242,N_6461);
xor U12149 (N_12149,N_6612,N_5744);
or U12150 (N_12150,N_5229,N_5774);
or U12151 (N_12151,N_9715,N_9725);
nand U12152 (N_12152,N_9778,N_9157);
and U12153 (N_12153,N_6009,N_7449);
or U12154 (N_12154,N_5003,N_5169);
and U12155 (N_12155,N_7056,N_7108);
nor U12156 (N_12156,N_6102,N_5051);
xnor U12157 (N_12157,N_9590,N_8195);
nand U12158 (N_12158,N_6390,N_9562);
nand U12159 (N_12159,N_7788,N_8252);
or U12160 (N_12160,N_9206,N_6320);
and U12161 (N_12161,N_5709,N_9748);
nor U12162 (N_12162,N_8031,N_7692);
or U12163 (N_12163,N_5037,N_6287);
nand U12164 (N_12164,N_9031,N_8820);
nand U12165 (N_12165,N_8805,N_6794);
nand U12166 (N_12166,N_9081,N_8908);
or U12167 (N_12167,N_9537,N_7184);
nand U12168 (N_12168,N_7620,N_5380);
and U12169 (N_12169,N_6630,N_8544);
and U12170 (N_12170,N_5455,N_5020);
nor U12171 (N_12171,N_5833,N_8920);
or U12172 (N_12172,N_5353,N_8524);
xor U12173 (N_12173,N_9642,N_6018);
nor U12174 (N_12174,N_6026,N_6066);
xor U12175 (N_12175,N_8600,N_6720);
and U12176 (N_12176,N_8354,N_5399);
and U12177 (N_12177,N_5590,N_5090);
nand U12178 (N_12178,N_9505,N_8056);
nor U12179 (N_12179,N_5017,N_6030);
nor U12180 (N_12180,N_9101,N_5811);
and U12181 (N_12181,N_7849,N_9386);
nor U12182 (N_12182,N_7011,N_8992);
or U12183 (N_12183,N_5614,N_5261);
or U12184 (N_12184,N_7294,N_7577);
and U12185 (N_12185,N_9020,N_6994);
or U12186 (N_12186,N_7749,N_8526);
or U12187 (N_12187,N_5827,N_5199);
or U12188 (N_12188,N_7562,N_9625);
and U12189 (N_12189,N_8271,N_7070);
and U12190 (N_12190,N_5038,N_9394);
or U12191 (N_12191,N_5296,N_5743);
nor U12192 (N_12192,N_9508,N_8346);
nor U12193 (N_12193,N_6489,N_5734);
nor U12194 (N_12194,N_5830,N_5395);
or U12195 (N_12195,N_6246,N_6079);
nand U12196 (N_12196,N_6544,N_9167);
nand U12197 (N_12197,N_9457,N_8441);
nand U12198 (N_12198,N_7195,N_6713);
and U12199 (N_12199,N_6029,N_5651);
nand U12200 (N_12200,N_6645,N_8250);
nor U12201 (N_12201,N_5370,N_6269);
and U12202 (N_12202,N_8019,N_9519);
nor U12203 (N_12203,N_8471,N_8591);
nor U12204 (N_12204,N_7455,N_5499);
and U12205 (N_12205,N_7444,N_7262);
nor U12206 (N_12206,N_8904,N_5137);
nor U12207 (N_12207,N_5819,N_9821);
nand U12208 (N_12208,N_6284,N_5154);
nor U12209 (N_12209,N_7244,N_8313);
nor U12210 (N_12210,N_6626,N_7439);
and U12211 (N_12211,N_9775,N_9271);
and U12212 (N_12212,N_5739,N_8186);
and U12213 (N_12213,N_9524,N_9067);
or U12214 (N_12214,N_8672,N_7831);
nand U12215 (N_12215,N_6444,N_6606);
nor U12216 (N_12216,N_9832,N_6531);
or U12217 (N_12217,N_5648,N_6838);
and U12218 (N_12218,N_8699,N_8549);
or U12219 (N_12219,N_9371,N_5987);
or U12220 (N_12220,N_8929,N_8755);
nor U12221 (N_12221,N_9088,N_5172);
nand U12222 (N_12222,N_5886,N_7682);
and U12223 (N_12223,N_7592,N_7622);
or U12224 (N_12224,N_6779,N_7531);
or U12225 (N_12225,N_6703,N_7342);
and U12226 (N_12226,N_8404,N_6206);
nand U12227 (N_12227,N_8946,N_6423);
xor U12228 (N_12228,N_8847,N_5071);
and U12229 (N_12229,N_7567,N_8263);
nand U12230 (N_12230,N_8940,N_8545);
or U12231 (N_12231,N_8382,N_5246);
nor U12232 (N_12232,N_8800,N_9259);
or U12233 (N_12233,N_8055,N_7219);
or U12234 (N_12234,N_6190,N_9288);
or U12235 (N_12235,N_6721,N_6475);
nand U12236 (N_12236,N_5144,N_7098);
and U12237 (N_12237,N_9634,N_8845);
nor U12238 (N_12238,N_5746,N_7391);
nand U12239 (N_12239,N_5572,N_9539);
nand U12240 (N_12240,N_8504,N_5479);
and U12241 (N_12241,N_5676,N_5244);
nor U12242 (N_12242,N_7353,N_5962);
nor U12243 (N_12243,N_9517,N_8751);
or U12244 (N_12244,N_8057,N_5197);
and U12245 (N_12245,N_7971,N_6569);
nor U12246 (N_12246,N_5209,N_6224);
nand U12247 (N_12247,N_6117,N_7356);
nor U12248 (N_12248,N_5151,N_6748);
or U12249 (N_12249,N_6866,N_7593);
nor U12250 (N_12250,N_8032,N_5640);
nand U12251 (N_12251,N_8638,N_5680);
or U12252 (N_12252,N_7220,N_5142);
or U12253 (N_12253,N_7329,N_6999);
nand U12254 (N_12254,N_8705,N_5621);
or U12255 (N_12255,N_7892,N_7637);
nand U12256 (N_12256,N_8193,N_7230);
nand U12257 (N_12257,N_8551,N_8237);
nor U12258 (N_12258,N_7147,N_9310);
or U12259 (N_12259,N_7420,N_5832);
xnor U12260 (N_12260,N_6506,N_7274);
and U12261 (N_12261,N_9451,N_5566);
and U12262 (N_12262,N_6596,N_7502);
or U12263 (N_12263,N_5582,N_8230);
or U12264 (N_12264,N_6397,N_7292);
or U12265 (N_12265,N_6800,N_5611);
xnor U12266 (N_12266,N_8496,N_7075);
or U12267 (N_12267,N_9441,N_8184);
nor U12268 (N_12268,N_9109,N_8505);
nand U12269 (N_12269,N_9660,N_7491);
nand U12270 (N_12270,N_7607,N_9159);
nor U12271 (N_12271,N_5182,N_8246);
nor U12272 (N_12272,N_5480,N_7972);
nand U12273 (N_12273,N_9287,N_9927);
or U12274 (N_12274,N_8208,N_9596);
or U12275 (N_12275,N_6350,N_8003);
nor U12276 (N_12276,N_6202,N_6765);
nor U12277 (N_12277,N_7205,N_5005);
nor U12278 (N_12278,N_7447,N_6411);
nor U12279 (N_12279,N_9571,N_9989);
or U12280 (N_12280,N_8405,N_5786);
nand U12281 (N_12281,N_7786,N_5649);
nor U12282 (N_12282,N_9172,N_5539);
nand U12283 (N_12283,N_8489,N_9309);
nor U12284 (N_12284,N_7922,N_8776);
nor U12285 (N_12285,N_5919,N_9121);
nand U12286 (N_12286,N_8131,N_7072);
or U12287 (N_12287,N_9068,N_7989);
nor U12288 (N_12288,N_7101,N_9753);
nand U12289 (N_12289,N_6808,N_6635);
nor U12290 (N_12290,N_6706,N_9364);
nand U12291 (N_12291,N_7214,N_9115);
nand U12292 (N_12292,N_9965,N_7630);
nor U12293 (N_12293,N_9683,N_7943);
nor U12294 (N_12294,N_5029,N_9491);
or U12295 (N_12295,N_9173,N_5273);
or U12296 (N_12296,N_9254,N_6728);
and U12297 (N_12297,N_8924,N_7224);
nand U12298 (N_12298,N_8533,N_7370);
nor U12299 (N_12299,N_7362,N_8978);
or U12300 (N_12300,N_8299,N_7032);
and U12301 (N_12301,N_7968,N_7528);
nand U12302 (N_12302,N_5560,N_6222);
or U12303 (N_12303,N_8786,N_9108);
nor U12304 (N_12304,N_6039,N_5507);
nor U12305 (N_12305,N_6200,N_9606);
nand U12306 (N_12306,N_5376,N_7819);
or U12307 (N_12307,N_5644,N_6218);
and U12308 (N_12308,N_8200,N_7536);
nor U12309 (N_12309,N_7207,N_6947);
nand U12310 (N_12310,N_7450,N_5297);
or U12311 (N_12311,N_8026,N_9564);
nor U12312 (N_12312,N_5141,N_8388);
or U12313 (N_12313,N_8518,N_5730);
xor U12314 (N_12314,N_5201,N_5317);
nand U12315 (N_12315,N_8188,N_8476);
nand U12316 (N_12316,N_6882,N_5671);
and U12317 (N_12317,N_9724,N_6653);
nor U12318 (N_12318,N_5314,N_5063);
or U12319 (N_12319,N_7557,N_5356);
nand U12320 (N_12320,N_8033,N_5108);
nor U12321 (N_12321,N_8173,N_9090);
nor U12322 (N_12322,N_8939,N_9217);
or U12323 (N_12323,N_5816,N_9887);
nor U12324 (N_12324,N_6601,N_9795);
nand U12325 (N_12325,N_6580,N_8010);
nor U12326 (N_12326,N_5843,N_5378);
nor U12327 (N_12327,N_8121,N_5405);
and U12328 (N_12328,N_9771,N_6179);
nand U12329 (N_12329,N_6835,N_8417);
nand U12330 (N_12330,N_7572,N_9011);
nor U12331 (N_12331,N_8711,N_5155);
nor U12332 (N_12332,N_9338,N_8721);
nand U12333 (N_12333,N_5262,N_5044);
nor U12334 (N_12334,N_5243,N_8095);
and U12335 (N_12335,N_9580,N_6727);
nand U12336 (N_12336,N_7432,N_5717);
nor U12337 (N_12337,N_7054,N_9812);
or U12338 (N_12338,N_6681,N_8429);
and U12339 (N_12339,N_5750,N_7700);
or U12340 (N_12340,N_9162,N_9709);
nor U12341 (N_12341,N_6072,N_6525);
and U12342 (N_12342,N_8345,N_8209);
nand U12343 (N_12343,N_9768,N_8068);
nand U12344 (N_12344,N_8029,N_5320);
and U12345 (N_12345,N_9733,N_9476);
and U12346 (N_12346,N_5205,N_8390);
or U12347 (N_12347,N_5007,N_7933);
or U12348 (N_12348,N_5288,N_6025);
or U12349 (N_12349,N_7833,N_8331);
xnor U12350 (N_12350,N_9578,N_5165);
and U12351 (N_12351,N_9655,N_5994);
nand U12352 (N_12352,N_5897,N_9789);
nand U12353 (N_12353,N_8609,N_7753);
nand U12354 (N_12354,N_5732,N_7168);
and U12355 (N_12355,N_9001,N_6233);
nor U12356 (N_12356,N_7746,N_6209);
and U12357 (N_12357,N_6415,N_6386);
nand U12358 (N_12358,N_9305,N_5656);
nor U12359 (N_12359,N_7626,N_8174);
or U12360 (N_12360,N_8120,N_9439);
nand U12361 (N_12361,N_9074,N_7467);
nor U12362 (N_12362,N_9478,N_6366);
nand U12363 (N_12363,N_9412,N_6889);
or U12364 (N_12364,N_5795,N_6045);
and U12365 (N_12365,N_8775,N_8327);
nor U12366 (N_12366,N_9856,N_7316);
nand U12367 (N_12367,N_8483,N_6132);
or U12368 (N_12368,N_8872,N_6333);
and U12369 (N_12369,N_9502,N_8887);
nor U12370 (N_12370,N_8362,N_8596);
and U12371 (N_12371,N_6634,N_6409);
or U12372 (N_12372,N_5672,N_8813);
nand U12373 (N_12373,N_8612,N_9855);
and U12374 (N_12374,N_6849,N_7534);
nand U12375 (N_12375,N_5542,N_9666);
and U12376 (N_12376,N_5248,N_6932);
and U12377 (N_12377,N_9065,N_7811);
nand U12378 (N_12378,N_5385,N_7872);
or U12379 (N_12379,N_7687,N_5829);
nor U12380 (N_12380,N_5164,N_8447);
or U12381 (N_12381,N_5522,N_6600);
nor U12382 (N_12382,N_6431,N_9820);
and U12383 (N_12383,N_7861,N_9773);
or U12384 (N_12384,N_7038,N_5956);
and U12385 (N_12385,N_8726,N_7818);
nand U12386 (N_12386,N_5227,N_8577);
nand U12387 (N_12387,N_7681,N_7590);
or U12388 (N_12388,N_9362,N_7009);
or U12389 (N_12389,N_5557,N_9998);
nand U12390 (N_12390,N_8511,N_5862);
and U12391 (N_12391,N_9029,N_8443);
nor U12392 (N_12392,N_9186,N_8054);
nor U12393 (N_12393,N_5081,N_8732);
and U12394 (N_12394,N_9837,N_9852);
and U12395 (N_12395,N_5441,N_8512);
nor U12396 (N_12396,N_6799,N_5633);
and U12397 (N_12397,N_7297,N_9260);
or U12398 (N_12398,N_9054,N_6586);
and U12399 (N_12399,N_5159,N_6769);
nand U12400 (N_12400,N_7898,N_5964);
and U12401 (N_12401,N_8426,N_9962);
nor U12402 (N_12402,N_5905,N_6060);
nor U12403 (N_12403,N_6436,N_7264);
nor U12404 (N_12404,N_7558,N_8937);
nor U12405 (N_12405,N_5174,N_7206);
nand U12406 (N_12406,N_8023,N_8850);
or U12407 (N_12407,N_5668,N_6120);
or U12408 (N_12408,N_9877,N_7166);
nor U12409 (N_12409,N_5313,N_7579);
nor U12410 (N_12410,N_9077,N_8855);
xnor U12411 (N_12411,N_7203,N_6483);
nand U12412 (N_12412,N_9790,N_9326);
nor U12413 (N_12413,N_5045,N_8135);
nand U12414 (N_12414,N_6504,N_6658);
nand U12415 (N_12415,N_8108,N_9993);
and U12416 (N_12416,N_8317,N_6257);
nor U12417 (N_12417,N_8750,N_9407);
or U12418 (N_12418,N_6754,N_6894);
nor U12419 (N_12419,N_9813,N_5753);
nor U12420 (N_12420,N_6307,N_5529);
nor U12421 (N_12421,N_7167,N_5929);
or U12422 (N_12422,N_6494,N_8369);
nand U12423 (N_12423,N_6832,N_9544);
nor U12424 (N_12424,N_8917,N_5578);
nand U12425 (N_12425,N_5257,N_6940);
nand U12426 (N_12426,N_5729,N_8901);
and U12427 (N_12427,N_6394,N_6105);
xor U12428 (N_12428,N_8493,N_5847);
nand U12429 (N_12429,N_6256,N_7795);
nor U12430 (N_12430,N_7561,N_7731);
and U12431 (N_12431,N_8868,N_9541);
nor U12432 (N_12432,N_8106,N_6715);
or U12433 (N_12433,N_8731,N_8798);
or U12434 (N_12434,N_9234,N_5062);
and U12435 (N_12435,N_6565,N_9100);
or U12436 (N_12436,N_8598,N_5792);
or U12437 (N_12437,N_8636,N_5333);
and U12438 (N_12438,N_7877,N_7537);
nor U12439 (N_12439,N_8425,N_5628);
nand U12440 (N_12440,N_6175,N_8934);
or U12441 (N_12441,N_8629,N_7125);
or U12442 (N_12442,N_5665,N_8819);
and U12443 (N_12443,N_9320,N_9593);
or U12444 (N_12444,N_6979,N_6587);
nor U12445 (N_12445,N_9592,N_7693);
and U12446 (N_12446,N_7340,N_7480);
or U12447 (N_12447,N_7066,N_6538);
nand U12448 (N_12448,N_8806,N_7518);
and U12449 (N_12449,N_5545,N_7187);
or U12450 (N_12450,N_5117,N_7904);
or U12451 (N_12451,N_6472,N_5995);
or U12452 (N_12452,N_8677,N_8663);
nand U12453 (N_12453,N_7132,N_9830);
or U12454 (N_12454,N_6365,N_9780);
nand U12455 (N_12455,N_5268,N_8661);
or U12456 (N_12456,N_6002,N_6448);
nand U12457 (N_12457,N_9212,N_6965);
and U12458 (N_12458,N_8796,N_6424);
and U12459 (N_12459,N_5128,N_7762);
and U12460 (N_12460,N_7273,N_8979);
nand U12461 (N_12461,N_7073,N_5584);
nor U12462 (N_12462,N_6954,N_7436);
and U12463 (N_12463,N_9664,N_6571);
or U12464 (N_12464,N_7366,N_5596);
and U12465 (N_12465,N_8586,N_6180);
nor U12466 (N_12466,N_7337,N_5466);
or U12467 (N_12467,N_7775,N_9405);
and U12468 (N_12468,N_9630,N_5998);
nor U12469 (N_12469,N_7464,N_7574);
nand U12470 (N_12470,N_6761,N_5773);
nor U12471 (N_12471,N_5922,N_5916);
and U12472 (N_12472,N_7202,N_8041);
or U12473 (N_12473,N_5834,N_9496);
nand U12474 (N_12474,N_7143,N_5363);
nand U12475 (N_12475,N_9850,N_6062);
and U12476 (N_12476,N_7714,N_9187);
nand U12477 (N_12477,N_6714,N_8603);
nand U12478 (N_12478,N_7323,N_9333);
and U12479 (N_12479,N_5828,N_5365);
or U12480 (N_12480,N_5200,N_8333);
nor U12481 (N_12481,N_5344,N_7465);
nor U12482 (N_12482,N_7690,N_7763);
and U12483 (N_12483,N_9410,N_7437);
or U12484 (N_12484,N_9523,N_7808);
or U12485 (N_12485,N_5857,N_9936);
nand U12486 (N_12486,N_8308,N_5869);
nand U12487 (N_12487,N_5602,N_6812);
and U12488 (N_12488,N_7953,N_7629);
and U12489 (N_12489,N_5883,N_6216);
nand U12490 (N_12490,N_8764,N_7673);
nand U12491 (N_12491,N_9682,N_6358);
nor U12492 (N_12492,N_9354,N_5513);
nand U12493 (N_12493,N_7734,N_8130);
nand U12494 (N_12494,N_7396,N_6435);
nor U12495 (N_12495,N_9737,N_9835);
or U12496 (N_12496,N_6830,N_5882);
or U12497 (N_12497,N_9467,N_5624);
nand U12498 (N_12498,N_7553,N_7041);
and U12499 (N_12499,N_7930,N_6459);
and U12500 (N_12500,N_5440,N_8904);
and U12501 (N_12501,N_7242,N_8029);
and U12502 (N_12502,N_8124,N_9939);
and U12503 (N_12503,N_9712,N_5229);
nor U12504 (N_12504,N_6076,N_6322);
or U12505 (N_12505,N_7158,N_5992);
and U12506 (N_12506,N_9366,N_9571);
or U12507 (N_12507,N_6720,N_6191);
nor U12508 (N_12508,N_9980,N_8988);
nand U12509 (N_12509,N_5983,N_9121);
nand U12510 (N_12510,N_7524,N_9992);
nand U12511 (N_12511,N_6541,N_5516);
and U12512 (N_12512,N_8075,N_6840);
nand U12513 (N_12513,N_6272,N_6237);
nor U12514 (N_12514,N_9659,N_5234);
and U12515 (N_12515,N_6820,N_7948);
nor U12516 (N_12516,N_8608,N_7621);
or U12517 (N_12517,N_7220,N_6664);
nor U12518 (N_12518,N_7714,N_9975);
or U12519 (N_12519,N_7270,N_5488);
or U12520 (N_12520,N_8970,N_6872);
nand U12521 (N_12521,N_9418,N_6510);
nor U12522 (N_12522,N_5497,N_7456);
and U12523 (N_12523,N_6182,N_7984);
nor U12524 (N_12524,N_7979,N_9551);
or U12525 (N_12525,N_7817,N_6853);
and U12526 (N_12526,N_5929,N_9908);
and U12527 (N_12527,N_7016,N_9371);
nor U12528 (N_12528,N_6209,N_8423);
nor U12529 (N_12529,N_7585,N_8137);
and U12530 (N_12530,N_6254,N_6753);
nand U12531 (N_12531,N_5763,N_6441);
nand U12532 (N_12532,N_9934,N_9286);
and U12533 (N_12533,N_5686,N_5200);
and U12534 (N_12534,N_9449,N_5882);
nor U12535 (N_12535,N_8511,N_6687);
nor U12536 (N_12536,N_9704,N_6524);
or U12537 (N_12537,N_9892,N_5012);
nand U12538 (N_12538,N_7662,N_6283);
or U12539 (N_12539,N_8256,N_8497);
and U12540 (N_12540,N_9642,N_8292);
xor U12541 (N_12541,N_6483,N_5036);
nor U12542 (N_12542,N_5306,N_8340);
nor U12543 (N_12543,N_7131,N_8208);
nand U12544 (N_12544,N_8386,N_9805);
or U12545 (N_12545,N_9763,N_7922);
nor U12546 (N_12546,N_9531,N_5308);
or U12547 (N_12547,N_7150,N_6085);
nand U12548 (N_12548,N_6528,N_7503);
and U12549 (N_12549,N_7080,N_7858);
nor U12550 (N_12550,N_8845,N_6076);
nand U12551 (N_12551,N_6751,N_5502);
nor U12552 (N_12552,N_6887,N_7950);
nor U12553 (N_12553,N_9434,N_6020);
and U12554 (N_12554,N_5856,N_5861);
or U12555 (N_12555,N_5022,N_7684);
nor U12556 (N_12556,N_5087,N_8324);
and U12557 (N_12557,N_6071,N_9472);
nor U12558 (N_12558,N_7845,N_9697);
and U12559 (N_12559,N_9981,N_5660);
nor U12560 (N_12560,N_5252,N_6208);
or U12561 (N_12561,N_7846,N_9703);
or U12562 (N_12562,N_8047,N_7481);
nor U12563 (N_12563,N_9290,N_9824);
or U12564 (N_12564,N_6218,N_5502);
nor U12565 (N_12565,N_9060,N_9105);
and U12566 (N_12566,N_7744,N_7290);
nor U12567 (N_12567,N_9886,N_6531);
and U12568 (N_12568,N_5607,N_6455);
and U12569 (N_12569,N_5175,N_9857);
or U12570 (N_12570,N_8261,N_9837);
nand U12571 (N_12571,N_7299,N_6037);
or U12572 (N_12572,N_6279,N_9115);
and U12573 (N_12573,N_9589,N_6977);
or U12574 (N_12574,N_8258,N_5791);
and U12575 (N_12575,N_8695,N_8991);
and U12576 (N_12576,N_6360,N_7677);
nor U12577 (N_12577,N_8206,N_9413);
or U12578 (N_12578,N_5876,N_8215);
or U12579 (N_12579,N_8241,N_5437);
nand U12580 (N_12580,N_5276,N_8274);
nor U12581 (N_12581,N_9161,N_8194);
nand U12582 (N_12582,N_9326,N_8444);
nor U12583 (N_12583,N_6719,N_6025);
nand U12584 (N_12584,N_9368,N_6311);
or U12585 (N_12585,N_6996,N_8498);
or U12586 (N_12586,N_5446,N_8314);
and U12587 (N_12587,N_8276,N_8482);
nor U12588 (N_12588,N_7127,N_5064);
and U12589 (N_12589,N_5676,N_7019);
nand U12590 (N_12590,N_6483,N_9013);
nand U12591 (N_12591,N_7782,N_6630);
and U12592 (N_12592,N_7195,N_5955);
or U12593 (N_12593,N_9901,N_8332);
nand U12594 (N_12594,N_8953,N_7127);
nor U12595 (N_12595,N_8160,N_7858);
and U12596 (N_12596,N_6101,N_7433);
and U12597 (N_12597,N_7306,N_7175);
nand U12598 (N_12598,N_6113,N_8486);
nor U12599 (N_12599,N_5646,N_9501);
and U12600 (N_12600,N_8805,N_7146);
and U12601 (N_12601,N_6850,N_6480);
or U12602 (N_12602,N_9721,N_5070);
nand U12603 (N_12603,N_5605,N_8375);
or U12604 (N_12604,N_5068,N_9825);
nand U12605 (N_12605,N_8908,N_6391);
nand U12606 (N_12606,N_9474,N_9489);
and U12607 (N_12607,N_8009,N_9042);
and U12608 (N_12608,N_5115,N_9508);
and U12609 (N_12609,N_5021,N_8549);
nor U12610 (N_12610,N_5737,N_6436);
and U12611 (N_12611,N_5415,N_9356);
and U12612 (N_12612,N_8065,N_9957);
and U12613 (N_12613,N_7932,N_9908);
xnor U12614 (N_12614,N_7652,N_8513);
nor U12615 (N_12615,N_5023,N_5057);
and U12616 (N_12616,N_5809,N_5922);
nand U12617 (N_12617,N_6587,N_7235);
nor U12618 (N_12618,N_5668,N_5496);
and U12619 (N_12619,N_9467,N_9776);
xor U12620 (N_12620,N_6660,N_9741);
and U12621 (N_12621,N_6382,N_5278);
or U12622 (N_12622,N_6412,N_8429);
or U12623 (N_12623,N_7271,N_7024);
nor U12624 (N_12624,N_5045,N_7730);
nand U12625 (N_12625,N_6363,N_7557);
or U12626 (N_12626,N_7895,N_6308);
and U12627 (N_12627,N_9148,N_5448);
nor U12628 (N_12628,N_7264,N_8900);
nand U12629 (N_12629,N_6494,N_6609);
nand U12630 (N_12630,N_6698,N_8999);
nand U12631 (N_12631,N_8028,N_5145);
nand U12632 (N_12632,N_6272,N_9312);
or U12633 (N_12633,N_8644,N_9460);
nand U12634 (N_12634,N_6986,N_8756);
or U12635 (N_12635,N_6916,N_5244);
nand U12636 (N_12636,N_6551,N_8874);
or U12637 (N_12637,N_6301,N_9279);
and U12638 (N_12638,N_6646,N_7153);
and U12639 (N_12639,N_5996,N_5752);
or U12640 (N_12640,N_6725,N_5340);
or U12641 (N_12641,N_8650,N_7044);
nand U12642 (N_12642,N_5261,N_7599);
nand U12643 (N_12643,N_6268,N_8765);
nor U12644 (N_12644,N_5093,N_8854);
nand U12645 (N_12645,N_8604,N_7914);
or U12646 (N_12646,N_8606,N_5143);
or U12647 (N_12647,N_6716,N_5873);
or U12648 (N_12648,N_7416,N_7445);
nand U12649 (N_12649,N_9091,N_8520);
nor U12650 (N_12650,N_9151,N_5772);
nand U12651 (N_12651,N_8338,N_6284);
and U12652 (N_12652,N_7446,N_5894);
or U12653 (N_12653,N_9547,N_9555);
nor U12654 (N_12654,N_5314,N_8197);
nand U12655 (N_12655,N_5377,N_5953);
nor U12656 (N_12656,N_7380,N_7323);
and U12657 (N_12657,N_9578,N_6188);
and U12658 (N_12658,N_9369,N_9048);
nand U12659 (N_12659,N_6256,N_5156);
or U12660 (N_12660,N_9467,N_6958);
and U12661 (N_12661,N_9851,N_7585);
or U12662 (N_12662,N_9846,N_9058);
or U12663 (N_12663,N_9908,N_7812);
or U12664 (N_12664,N_5018,N_7766);
and U12665 (N_12665,N_9505,N_7531);
nor U12666 (N_12666,N_9018,N_5778);
and U12667 (N_12667,N_8377,N_9531);
or U12668 (N_12668,N_7250,N_9850);
or U12669 (N_12669,N_9646,N_7534);
nor U12670 (N_12670,N_9962,N_6074);
and U12671 (N_12671,N_8827,N_5418);
and U12672 (N_12672,N_5970,N_7620);
and U12673 (N_12673,N_6018,N_5456);
nand U12674 (N_12674,N_7693,N_5430);
and U12675 (N_12675,N_6237,N_7667);
nand U12676 (N_12676,N_9321,N_8314);
or U12677 (N_12677,N_5181,N_8444);
and U12678 (N_12678,N_8881,N_9330);
nor U12679 (N_12679,N_7917,N_8929);
or U12680 (N_12680,N_5656,N_8075);
and U12681 (N_12681,N_6472,N_9045);
nor U12682 (N_12682,N_7476,N_9688);
nor U12683 (N_12683,N_9009,N_8367);
or U12684 (N_12684,N_8654,N_8003);
or U12685 (N_12685,N_8093,N_5887);
nor U12686 (N_12686,N_7863,N_8530);
nand U12687 (N_12687,N_6928,N_6313);
nor U12688 (N_12688,N_8307,N_6664);
nand U12689 (N_12689,N_6614,N_6420);
nor U12690 (N_12690,N_7049,N_6478);
nor U12691 (N_12691,N_6633,N_5733);
and U12692 (N_12692,N_8105,N_6949);
nand U12693 (N_12693,N_7216,N_9855);
and U12694 (N_12694,N_9068,N_8070);
or U12695 (N_12695,N_5464,N_7044);
nand U12696 (N_12696,N_8848,N_8659);
nor U12697 (N_12697,N_5721,N_9464);
or U12698 (N_12698,N_9866,N_5666);
and U12699 (N_12699,N_8456,N_5831);
or U12700 (N_12700,N_7264,N_6243);
or U12701 (N_12701,N_6398,N_6093);
nor U12702 (N_12702,N_6888,N_5851);
nand U12703 (N_12703,N_7163,N_9787);
nand U12704 (N_12704,N_8127,N_9981);
and U12705 (N_12705,N_7777,N_9765);
or U12706 (N_12706,N_9732,N_5940);
or U12707 (N_12707,N_5233,N_9055);
and U12708 (N_12708,N_7555,N_9411);
and U12709 (N_12709,N_7621,N_6726);
nor U12710 (N_12710,N_9398,N_6388);
nor U12711 (N_12711,N_6784,N_7152);
nor U12712 (N_12712,N_8061,N_7705);
nor U12713 (N_12713,N_8822,N_8792);
nand U12714 (N_12714,N_8763,N_8059);
nand U12715 (N_12715,N_5038,N_7752);
or U12716 (N_12716,N_7969,N_8188);
nor U12717 (N_12717,N_7775,N_9499);
nor U12718 (N_12718,N_5040,N_8043);
nand U12719 (N_12719,N_9178,N_7999);
nor U12720 (N_12720,N_7663,N_9391);
nand U12721 (N_12721,N_6410,N_6833);
nand U12722 (N_12722,N_5564,N_7740);
or U12723 (N_12723,N_5426,N_7769);
nor U12724 (N_12724,N_7507,N_5775);
and U12725 (N_12725,N_6776,N_8677);
or U12726 (N_12726,N_6917,N_6836);
or U12727 (N_12727,N_9545,N_9450);
nand U12728 (N_12728,N_7992,N_7977);
or U12729 (N_12729,N_7625,N_9036);
nor U12730 (N_12730,N_7763,N_6465);
and U12731 (N_12731,N_9290,N_8614);
nand U12732 (N_12732,N_5657,N_5750);
nor U12733 (N_12733,N_7730,N_8319);
nand U12734 (N_12734,N_6660,N_8305);
nor U12735 (N_12735,N_9807,N_5128);
xor U12736 (N_12736,N_8334,N_7448);
nor U12737 (N_12737,N_7869,N_5094);
nor U12738 (N_12738,N_5742,N_9940);
and U12739 (N_12739,N_7614,N_9558);
or U12740 (N_12740,N_9123,N_7901);
and U12741 (N_12741,N_6483,N_5495);
nand U12742 (N_12742,N_6560,N_5324);
or U12743 (N_12743,N_9699,N_7892);
nand U12744 (N_12744,N_5557,N_9282);
and U12745 (N_12745,N_7804,N_8388);
or U12746 (N_12746,N_9563,N_6474);
and U12747 (N_12747,N_9682,N_9271);
or U12748 (N_12748,N_8411,N_6022);
or U12749 (N_12749,N_5554,N_9384);
nor U12750 (N_12750,N_6059,N_6441);
or U12751 (N_12751,N_5717,N_9651);
nor U12752 (N_12752,N_9128,N_8504);
nor U12753 (N_12753,N_9770,N_8886);
nor U12754 (N_12754,N_9219,N_5892);
and U12755 (N_12755,N_8156,N_7982);
nor U12756 (N_12756,N_7641,N_5907);
and U12757 (N_12757,N_7512,N_6565);
nand U12758 (N_12758,N_8143,N_7249);
and U12759 (N_12759,N_7052,N_5651);
nor U12760 (N_12760,N_8955,N_8611);
or U12761 (N_12761,N_6843,N_7939);
nor U12762 (N_12762,N_9815,N_9833);
and U12763 (N_12763,N_7665,N_8087);
and U12764 (N_12764,N_8948,N_9056);
and U12765 (N_12765,N_8224,N_6449);
or U12766 (N_12766,N_9194,N_7043);
nor U12767 (N_12767,N_7526,N_6826);
nand U12768 (N_12768,N_9181,N_6400);
or U12769 (N_12769,N_8214,N_7238);
or U12770 (N_12770,N_5788,N_6828);
nor U12771 (N_12771,N_7423,N_8389);
nand U12772 (N_12772,N_6010,N_9374);
or U12773 (N_12773,N_5562,N_8458);
xnor U12774 (N_12774,N_6111,N_8336);
nand U12775 (N_12775,N_5187,N_7752);
nor U12776 (N_12776,N_7340,N_9493);
and U12777 (N_12777,N_6149,N_6585);
and U12778 (N_12778,N_6337,N_8359);
nand U12779 (N_12779,N_7812,N_8931);
and U12780 (N_12780,N_9168,N_9284);
and U12781 (N_12781,N_8070,N_6478);
nor U12782 (N_12782,N_9443,N_9759);
xor U12783 (N_12783,N_9634,N_7574);
and U12784 (N_12784,N_6526,N_9181);
nor U12785 (N_12785,N_6981,N_7328);
nor U12786 (N_12786,N_8326,N_6185);
or U12787 (N_12787,N_8286,N_8458);
and U12788 (N_12788,N_5847,N_7523);
and U12789 (N_12789,N_5251,N_5871);
nand U12790 (N_12790,N_8955,N_9647);
nand U12791 (N_12791,N_7795,N_5084);
or U12792 (N_12792,N_5669,N_9715);
and U12793 (N_12793,N_6923,N_7587);
or U12794 (N_12794,N_7812,N_7917);
nor U12795 (N_12795,N_9764,N_9506);
and U12796 (N_12796,N_5211,N_8173);
nor U12797 (N_12797,N_7861,N_9571);
or U12798 (N_12798,N_6026,N_5215);
nand U12799 (N_12799,N_8731,N_8919);
and U12800 (N_12800,N_8560,N_5759);
or U12801 (N_12801,N_7350,N_7459);
nand U12802 (N_12802,N_5178,N_5750);
nor U12803 (N_12803,N_8372,N_8872);
nor U12804 (N_12804,N_8976,N_8665);
or U12805 (N_12805,N_8488,N_6802);
and U12806 (N_12806,N_7332,N_6026);
and U12807 (N_12807,N_6783,N_5137);
xnor U12808 (N_12808,N_6766,N_8696);
and U12809 (N_12809,N_8084,N_6435);
or U12810 (N_12810,N_9745,N_6606);
nor U12811 (N_12811,N_5495,N_5421);
nand U12812 (N_12812,N_9114,N_9647);
nor U12813 (N_12813,N_9094,N_7256);
nand U12814 (N_12814,N_9416,N_8434);
nand U12815 (N_12815,N_8123,N_7774);
nor U12816 (N_12816,N_8895,N_8447);
nor U12817 (N_12817,N_5395,N_8194);
nand U12818 (N_12818,N_7377,N_5042);
nor U12819 (N_12819,N_6452,N_5980);
nor U12820 (N_12820,N_5666,N_5116);
nor U12821 (N_12821,N_9292,N_6797);
nand U12822 (N_12822,N_7816,N_8091);
nor U12823 (N_12823,N_5450,N_7868);
or U12824 (N_12824,N_7034,N_9352);
or U12825 (N_12825,N_8761,N_9161);
and U12826 (N_12826,N_9189,N_8623);
nor U12827 (N_12827,N_7388,N_8693);
nand U12828 (N_12828,N_7335,N_9422);
or U12829 (N_12829,N_7816,N_7886);
and U12830 (N_12830,N_8448,N_9877);
nor U12831 (N_12831,N_6614,N_7824);
nor U12832 (N_12832,N_8887,N_8804);
and U12833 (N_12833,N_6250,N_9428);
and U12834 (N_12834,N_7510,N_9639);
nor U12835 (N_12835,N_6901,N_5778);
nand U12836 (N_12836,N_9640,N_7407);
or U12837 (N_12837,N_5004,N_7984);
nand U12838 (N_12838,N_5376,N_6637);
xor U12839 (N_12839,N_6938,N_6046);
and U12840 (N_12840,N_8486,N_6806);
and U12841 (N_12841,N_9948,N_7024);
nor U12842 (N_12842,N_7408,N_8008);
or U12843 (N_12843,N_7850,N_7461);
nand U12844 (N_12844,N_9752,N_8971);
and U12845 (N_12845,N_8082,N_6827);
or U12846 (N_12846,N_9433,N_6420);
or U12847 (N_12847,N_5661,N_7907);
nor U12848 (N_12848,N_5931,N_9149);
nor U12849 (N_12849,N_6368,N_9715);
nand U12850 (N_12850,N_8029,N_8728);
nor U12851 (N_12851,N_7177,N_5218);
nand U12852 (N_12852,N_6855,N_6556);
nor U12853 (N_12853,N_9964,N_8615);
nand U12854 (N_12854,N_8912,N_9021);
nand U12855 (N_12855,N_5869,N_7890);
nand U12856 (N_12856,N_6694,N_6828);
nor U12857 (N_12857,N_8692,N_9852);
and U12858 (N_12858,N_6564,N_6096);
and U12859 (N_12859,N_6554,N_7686);
or U12860 (N_12860,N_9230,N_8081);
and U12861 (N_12861,N_5887,N_5493);
and U12862 (N_12862,N_9515,N_7899);
nor U12863 (N_12863,N_8950,N_9619);
xor U12864 (N_12864,N_8091,N_7455);
or U12865 (N_12865,N_6378,N_6650);
nor U12866 (N_12866,N_9539,N_7401);
and U12867 (N_12867,N_8405,N_9257);
nand U12868 (N_12868,N_7688,N_8745);
nor U12869 (N_12869,N_5408,N_5587);
nor U12870 (N_12870,N_8483,N_7319);
or U12871 (N_12871,N_8270,N_9139);
nor U12872 (N_12872,N_7740,N_6498);
and U12873 (N_12873,N_5742,N_8696);
nand U12874 (N_12874,N_6823,N_8482);
nor U12875 (N_12875,N_8007,N_6390);
and U12876 (N_12876,N_9189,N_8882);
or U12877 (N_12877,N_8889,N_5043);
and U12878 (N_12878,N_8332,N_6267);
or U12879 (N_12879,N_7714,N_7008);
nor U12880 (N_12880,N_7681,N_7557);
and U12881 (N_12881,N_6507,N_7825);
nor U12882 (N_12882,N_7236,N_8515);
nand U12883 (N_12883,N_7274,N_8927);
and U12884 (N_12884,N_9827,N_5159);
or U12885 (N_12885,N_7512,N_7854);
and U12886 (N_12886,N_8948,N_6139);
nor U12887 (N_12887,N_9891,N_9617);
and U12888 (N_12888,N_9434,N_7502);
nor U12889 (N_12889,N_8462,N_7229);
nand U12890 (N_12890,N_9441,N_6240);
or U12891 (N_12891,N_8602,N_6490);
nor U12892 (N_12892,N_9079,N_8679);
nor U12893 (N_12893,N_6524,N_5063);
or U12894 (N_12894,N_5116,N_8806);
or U12895 (N_12895,N_7795,N_7543);
nor U12896 (N_12896,N_5994,N_5604);
nand U12897 (N_12897,N_7118,N_7238);
and U12898 (N_12898,N_7138,N_7688);
and U12899 (N_12899,N_9867,N_8225);
nor U12900 (N_12900,N_9403,N_6322);
nor U12901 (N_12901,N_6305,N_8676);
or U12902 (N_12902,N_5601,N_7146);
nand U12903 (N_12903,N_9919,N_9250);
nor U12904 (N_12904,N_9388,N_8443);
or U12905 (N_12905,N_5409,N_6203);
and U12906 (N_12906,N_9143,N_9984);
nand U12907 (N_12907,N_7724,N_8143);
and U12908 (N_12908,N_5636,N_8137);
nor U12909 (N_12909,N_9892,N_7955);
nand U12910 (N_12910,N_6330,N_5685);
and U12911 (N_12911,N_8430,N_9635);
or U12912 (N_12912,N_5029,N_5543);
nor U12913 (N_12913,N_6855,N_6365);
and U12914 (N_12914,N_9537,N_7203);
nor U12915 (N_12915,N_9864,N_6248);
and U12916 (N_12916,N_8153,N_8935);
or U12917 (N_12917,N_9065,N_7255);
and U12918 (N_12918,N_5031,N_5796);
or U12919 (N_12919,N_8636,N_8453);
nor U12920 (N_12920,N_6359,N_8254);
or U12921 (N_12921,N_8694,N_8890);
and U12922 (N_12922,N_6722,N_7268);
or U12923 (N_12923,N_8171,N_9221);
nor U12924 (N_12924,N_9333,N_9700);
and U12925 (N_12925,N_7825,N_8872);
nor U12926 (N_12926,N_8537,N_6906);
and U12927 (N_12927,N_8892,N_5908);
nor U12928 (N_12928,N_9733,N_6748);
nand U12929 (N_12929,N_9223,N_8190);
or U12930 (N_12930,N_5149,N_6344);
and U12931 (N_12931,N_9009,N_8307);
nand U12932 (N_12932,N_7965,N_8950);
and U12933 (N_12933,N_5380,N_7382);
nor U12934 (N_12934,N_6311,N_9362);
or U12935 (N_12935,N_9456,N_7089);
nor U12936 (N_12936,N_5141,N_9287);
xor U12937 (N_12937,N_8192,N_5409);
or U12938 (N_12938,N_5795,N_9981);
nor U12939 (N_12939,N_5801,N_8520);
nand U12940 (N_12940,N_9491,N_6734);
nand U12941 (N_12941,N_7620,N_5448);
or U12942 (N_12942,N_9100,N_6059);
or U12943 (N_12943,N_5848,N_9114);
and U12944 (N_12944,N_9765,N_6450);
or U12945 (N_12945,N_8786,N_9636);
nor U12946 (N_12946,N_5478,N_5722);
or U12947 (N_12947,N_5825,N_7273);
nor U12948 (N_12948,N_6938,N_7678);
or U12949 (N_12949,N_9900,N_6120);
or U12950 (N_12950,N_5059,N_7861);
or U12951 (N_12951,N_7285,N_6250);
or U12952 (N_12952,N_5626,N_9327);
and U12953 (N_12953,N_9325,N_9365);
nor U12954 (N_12954,N_6783,N_8198);
and U12955 (N_12955,N_5175,N_8819);
or U12956 (N_12956,N_8704,N_5349);
nand U12957 (N_12957,N_8281,N_9350);
nor U12958 (N_12958,N_5026,N_8907);
nand U12959 (N_12959,N_7118,N_8130);
and U12960 (N_12960,N_6824,N_8605);
nor U12961 (N_12961,N_8228,N_8317);
or U12962 (N_12962,N_6551,N_8525);
nand U12963 (N_12963,N_5245,N_7361);
nand U12964 (N_12964,N_6920,N_6624);
nor U12965 (N_12965,N_7234,N_5217);
nor U12966 (N_12966,N_5967,N_6468);
or U12967 (N_12967,N_5004,N_6661);
and U12968 (N_12968,N_7667,N_6577);
and U12969 (N_12969,N_5729,N_7957);
and U12970 (N_12970,N_7121,N_8643);
or U12971 (N_12971,N_8695,N_9999);
or U12972 (N_12972,N_9933,N_6145);
or U12973 (N_12973,N_8074,N_5832);
nor U12974 (N_12974,N_5796,N_7111);
or U12975 (N_12975,N_9919,N_5972);
nand U12976 (N_12976,N_9110,N_6806);
nand U12977 (N_12977,N_6636,N_8764);
nand U12978 (N_12978,N_8704,N_9174);
nand U12979 (N_12979,N_9363,N_7751);
and U12980 (N_12980,N_5153,N_8891);
or U12981 (N_12981,N_5258,N_6272);
or U12982 (N_12982,N_5472,N_5032);
nand U12983 (N_12983,N_6549,N_9821);
nand U12984 (N_12984,N_6733,N_5363);
xnor U12985 (N_12985,N_7543,N_6659);
nand U12986 (N_12986,N_6117,N_5992);
nand U12987 (N_12987,N_9818,N_7809);
nor U12988 (N_12988,N_9051,N_5614);
nand U12989 (N_12989,N_6252,N_9602);
or U12990 (N_12990,N_6035,N_9596);
xor U12991 (N_12991,N_5360,N_7879);
nor U12992 (N_12992,N_5214,N_7686);
or U12993 (N_12993,N_8823,N_9253);
nand U12994 (N_12994,N_6424,N_9164);
and U12995 (N_12995,N_9811,N_8205);
and U12996 (N_12996,N_7019,N_9484);
nand U12997 (N_12997,N_7686,N_8254);
and U12998 (N_12998,N_6171,N_5465);
nor U12999 (N_12999,N_5100,N_7106);
nand U13000 (N_13000,N_7465,N_9143);
and U13001 (N_13001,N_8062,N_5362);
or U13002 (N_13002,N_9233,N_6600);
nor U13003 (N_13003,N_7589,N_7409);
nand U13004 (N_13004,N_7154,N_6622);
or U13005 (N_13005,N_9397,N_9015);
nand U13006 (N_13006,N_6926,N_5178);
and U13007 (N_13007,N_7812,N_8660);
nand U13008 (N_13008,N_8759,N_9182);
and U13009 (N_13009,N_9102,N_5647);
or U13010 (N_13010,N_7899,N_8074);
and U13011 (N_13011,N_8176,N_8771);
nand U13012 (N_13012,N_9493,N_9393);
or U13013 (N_13013,N_6876,N_7564);
and U13014 (N_13014,N_5117,N_7096);
or U13015 (N_13015,N_7066,N_5098);
nand U13016 (N_13016,N_5005,N_8812);
and U13017 (N_13017,N_8947,N_9168);
or U13018 (N_13018,N_6135,N_5164);
and U13019 (N_13019,N_8413,N_5681);
nor U13020 (N_13020,N_6879,N_5338);
or U13021 (N_13021,N_7751,N_9940);
or U13022 (N_13022,N_8575,N_8417);
nor U13023 (N_13023,N_5174,N_7494);
nor U13024 (N_13024,N_8974,N_8488);
nor U13025 (N_13025,N_8194,N_7593);
and U13026 (N_13026,N_6850,N_7972);
nor U13027 (N_13027,N_5194,N_9333);
nor U13028 (N_13028,N_7786,N_6879);
or U13029 (N_13029,N_8726,N_6285);
nand U13030 (N_13030,N_7988,N_8984);
nand U13031 (N_13031,N_9849,N_6807);
and U13032 (N_13032,N_6722,N_7808);
and U13033 (N_13033,N_8676,N_7184);
nor U13034 (N_13034,N_9046,N_9701);
nor U13035 (N_13035,N_8225,N_9779);
or U13036 (N_13036,N_9382,N_5112);
and U13037 (N_13037,N_7508,N_9264);
or U13038 (N_13038,N_9702,N_6756);
nor U13039 (N_13039,N_8554,N_6526);
or U13040 (N_13040,N_9589,N_5204);
nand U13041 (N_13041,N_9210,N_5806);
nor U13042 (N_13042,N_6505,N_9008);
nand U13043 (N_13043,N_7048,N_7933);
nor U13044 (N_13044,N_5706,N_7366);
or U13045 (N_13045,N_8694,N_9231);
nor U13046 (N_13046,N_8595,N_8349);
and U13047 (N_13047,N_9034,N_7829);
xnor U13048 (N_13048,N_7623,N_8043);
or U13049 (N_13049,N_5058,N_8386);
nand U13050 (N_13050,N_6284,N_8751);
or U13051 (N_13051,N_6744,N_8714);
nand U13052 (N_13052,N_7951,N_5749);
nor U13053 (N_13053,N_6730,N_7525);
or U13054 (N_13054,N_7948,N_5951);
nand U13055 (N_13055,N_8502,N_6284);
and U13056 (N_13056,N_7863,N_8365);
or U13057 (N_13057,N_6717,N_5974);
or U13058 (N_13058,N_5808,N_8084);
nand U13059 (N_13059,N_5353,N_5052);
and U13060 (N_13060,N_5280,N_6588);
and U13061 (N_13061,N_5975,N_6115);
and U13062 (N_13062,N_9120,N_8016);
nor U13063 (N_13063,N_7311,N_9116);
nand U13064 (N_13064,N_9779,N_9954);
nand U13065 (N_13065,N_7491,N_5554);
and U13066 (N_13066,N_5205,N_5719);
nand U13067 (N_13067,N_7733,N_6727);
nor U13068 (N_13068,N_5842,N_6357);
nand U13069 (N_13069,N_7324,N_8055);
and U13070 (N_13070,N_5722,N_8515);
nor U13071 (N_13071,N_9346,N_5855);
nor U13072 (N_13072,N_7533,N_5007);
nor U13073 (N_13073,N_7701,N_5294);
and U13074 (N_13074,N_6044,N_8929);
or U13075 (N_13075,N_6084,N_8252);
and U13076 (N_13076,N_7259,N_5074);
and U13077 (N_13077,N_7950,N_6679);
nand U13078 (N_13078,N_5753,N_8981);
xor U13079 (N_13079,N_8286,N_6153);
nor U13080 (N_13080,N_5668,N_8877);
or U13081 (N_13081,N_9525,N_8871);
nor U13082 (N_13082,N_6605,N_5660);
and U13083 (N_13083,N_6075,N_8091);
and U13084 (N_13084,N_5948,N_5988);
and U13085 (N_13085,N_6245,N_7943);
nor U13086 (N_13086,N_8351,N_7568);
nand U13087 (N_13087,N_7844,N_9923);
and U13088 (N_13088,N_7337,N_9412);
or U13089 (N_13089,N_8828,N_6622);
or U13090 (N_13090,N_9693,N_6869);
and U13091 (N_13091,N_5699,N_9644);
nor U13092 (N_13092,N_9368,N_6155);
nand U13093 (N_13093,N_9054,N_9773);
and U13094 (N_13094,N_6763,N_8359);
nand U13095 (N_13095,N_6339,N_8664);
nor U13096 (N_13096,N_6673,N_6596);
or U13097 (N_13097,N_8446,N_8058);
and U13098 (N_13098,N_7545,N_8014);
and U13099 (N_13099,N_6699,N_8051);
or U13100 (N_13100,N_6051,N_9527);
or U13101 (N_13101,N_9875,N_8457);
nor U13102 (N_13102,N_7168,N_5977);
and U13103 (N_13103,N_6199,N_8544);
nor U13104 (N_13104,N_8059,N_6892);
nor U13105 (N_13105,N_9521,N_8693);
or U13106 (N_13106,N_8649,N_6800);
or U13107 (N_13107,N_8479,N_5721);
or U13108 (N_13108,N_5175,N_8997);
xor U13109 (N_13109,N_8538,N_5219);
or U13110 (N_13110,N_5363,N_7959);
and U13111 (N_13111,N_5287,N_5171);
and U13112 (N_13112,N_5739,N_6359);
and U13113 (N_13113,N_9798,N_6929);
or U13114 (N_13114,N_7621,N_8334);
nand U13115 (N_13115,N_6358,N_5746);
nor U13116 (N_13116,N_8005,N_7512);
xnor U13117 (N_13117,N_9003,N_9043);
nor U13118 (N_13118,N_7608,N_8110);
nor U13119 (N_13119,N_9793,N_6532);
or U13120 (N_13120,N_5056,N_5810);
nor U13121 (N_13121,N_6111,N_8587);
nor U13122 (N_13122,N_8026,N_8676);
nor U13123 (N_13123,N_9387,N_5549);
and U13124 (N_13124,N_5916,N_9969);
and U13125 (N_13125,N_6192,N_5680);
nand U13126 (N_13126,N_7294,N_9105);
nor U13127 (N_13127,N_9684,N_8596);
nor U13128 (N_13128,N_6511,N_6911);
or U13129 (N_13129,N_8006,N_7001);
or U13130 (N_13130,N_8135,N_8831);
or U13131 (N_13131,N_9307,N_5116);
and U13132 (N_13132,N_7613,N_6717);
or U13133 (N_13133,N_6435,N_8195);
nand U13134 (N_13134,N_6555,N_7090);
and U13135 (N_13135,N_5599,N_5918);
nand U13136 (N_13136,N_8884,N_8644);
and U13137 (N_13137,N_8157,N_8524);
and U13138 (N_13138,N_9972,N_8556);
and U13139 (N_13139,N_5535,N_6609);
and U13140 (N_13140,N_5790,N_5853);
nor U13141 (N_13141,N_7126,N_8855);
or U13142 (N_13142,N_6270,N_6511);
nand U13143 (N_13143,N_7063,N_7318);
nor U13144 (N_13144,N_6312,N_7087);
or U13145 (N_13145,N_6060,N_9412);
or U13146 (N_13146,N_6125,N_8393);
and U13147 (N_13147,N_7916,N_5738);
or U13148 (N_13148,N_8755,N_8422);
or U13149 (N_13149,N_9546,N_6917);
or U13150 (N_13150,N_6250,N_5567);
and U13151 (N_13151,N_9629,N_8367);
nand U13152 (N_13152,N_6036,N_8186);
and U13153 (N_13153,N_7397,N_8286);
or U13154 (N_13154,N_6716,N_8873);
or U13155 (N_13155,N_6057,N_9342);
nor U13156 (N_13156,N_9296,N_9397);
or U13157 (N_13157,N_6948,N_9105);
and U13158 (N_13158,N_8318,N_8029);
nor U13159 (N_13159,N_6947,N_5190);
or U13160 (N_13160,N_8722,N_8737);
and U13161 (N_13161,N_9284,N_6261);
nand U13162 (N_13162,N_7749,N_9572);
or U13163 (N_13163,N_9143,N_9788);
or U13164 (N_13164,N_9307,N_9952);
and U13165 (N_13165,N_8431,N_8931);
and U13166 (N_13166,N_9183,N_6027);
nand U13167 (N_13167,N_7960,N_8594);
nor U13168 (N_13168,N_8317,N_8176);
nor U13169 (N_13169,N_7939,N_5314);
and U13170 (N_13170,N_6210,N_8582);
nor U13171 (N_13171,N_6582,N_5481);
nand U13172 (N_13172,N_7245,N_6292);
or U13173 (N_13173,N_6575,N_8814);
nor U13174 (N_13174,N_8214,N_7831);
nand U13175 (N_13175,N_9302,N_8025);
nand U13176 (N_13176,N_5338,N_6302);
and U13177 (N_13177,N_7876,N_6981);
and U13178 (N_13178,N_8511,N_6131);
and U13179 (N_13179,N_7315,N_8633);
nor U13180 (N_13180,N_5253,N_6848);
and U13181 (N_13181,N_7177,N_5907);
nand U13182 (N_13182,N_8878,N_5765);
and U13183 (N_13183,N_9044,N_6063);
or U13184 (N_13184,N_5907,N_9402);
and U13185 (N_13185,N_9825,N_6218);
or U13186 (N_13186,N_9588,N_5257);
nand U13187 (N_13187,N_6050,N_5303);
nand U13188 (N_13188,N_5960,N_6847);
and U13189 (N_13189,N_7423,N_7801);
or U13190 (N_13190,N_8079,N_5891);
or U13191 (N_13191,N_6159,N_9572);
nand U13192 (N_13192,N_7950,N_8456);
or U13193 (N_13193,N_6629,N_9945);
nand U13194 (N_13194,N_6013,N_6712);
nand U13195 (N_13195,N_6098,N_6312);
or U13196 (N_13196,N_6282,N_5884);
and U13197 (N_13197,N_5148,N_6763);
nor U13198 (N_13198,N_5858,N_6441);
nor U13199 (N_13199,N_8424,N_9796);
and U13200 (N_13200,N_7415,N_5098);
nor U13201 (N_13201,N_7814,N_9712);
and U13202 (N_13202,N_8439,N_9415);
nand U13203 (N_13203,N_7998,N_8672);
and U13204 (N_13204,N_9895,N_5143);
nand U13205 (N_13205,N_9415,N_8844);
nand U13206 (N_13206,N_6130,N_6597);
and U13207 (N_13207,N_5323,N_6592);
nor U13208 (N_13208,N_8130,N_8903);
nand U13209 (N_13209,N_7846,N_9983);
and U13210 (N_13210,N_9488,N_5519);
and U13211 (N_13211,N_7603,N_6105);
or U13212 (N_13212,N_5890,N_9380);
and U13213 (N_13213,N_6570,N_8613);
or U13214 (N_13214,N_6087,N_8751);
or U13215 (N_13215,N_9512,N_8765);
nor U13216 (N_13216,N_5317,N_9676);
and U13217 (N_13217,N_7970,N_5537);
nand U13218 (N_13218,N_8371,N_9253);
nor U13219 (N_13219,N_6097,N_9899);
nor U13220 (N_13220,N_9901,N_7465);
or U13221 (N_13221,N_5752,N_9891);
nand U13222 (N_13222,N_8889,N_6605);
nand U13223 (N_13223,N_9715,N_5505);
or U13224 (N_13224,N_6270,N_8124);
nand U13225 (N_13225,N_8151,N_5467);
nand U13226 (N_13226,N_6862,N_8674);
or U13227 (N_13227,N_8270,N_8700);
nand U13228 (N_13228,N_6752,N_8371);
nor U13229 (N_13229,N_6852,N_8342);
or U13230 (N_13230,N_7071,N_5455);
or U13231 (N_13231,N_9505,N_9662);
or U13232 (N_13232,N_5171,N_7545);
nor U13233 (N_13233,N_9899,N_6187);
nand U13234 (N_13234,N_6009,N_8295);
or U13235 (N_13235,N_6027,N_7769);
or U13236 (N_13236,N_8628,N_5350);
nand U13237 (N_13237,N_6370,N_6719);
nor U13238 (N_13238,N_6128,N_8555);
nor U13239 (N_13239,N_7015,N_5877);
or U13240 (N_13240,N_7054,N_9972);
nand U13241 (N_13241,N_6034,N_9045);
nand U13242 (N_13242,N_5107,N_9833);
and U13243 (N_13243,N_9882,N_7815);
nor U13244 (N_13244,N_7399,N_9942);
and U13245 (N_13245,N_8678,N_8839);
and U13246 (N_13246,N_9608,N_5816);
and U13247 (N_13247,N_6459,N_9422);
nand U13248 (N_13248,N_9685,N_6735);
or U13249 (N_13249,N_6843,N_6008);
nand U13250 (N_13250,N_5763,N_6910);
nand U13251 (N_13251,N_8614,N_5323);
and U13252 (N_13252,N_5303,N_6668);
nor U13253 (N_13253,N_6275,N_8773);
nand U13254 (N_13254,N_6598,N_7142);
nor U13255 (N_13255,N_7045,N_7039);
nor U13256 (N_13256,N_6435,N_7276);
or U13257 (N_13257,N_6289,N_5265);
or U13258 (N_13258,N_7877,N_6877);
or U13259 (N_13259,N_9031,N_8674);
nor U13260 (N_13260,N_5835,N_9874);
or U13261 (N_13261,N_5558,N_8843);
nand U13262 (N_13262,N_7672,N_6237);
nand U13263 (N_13263,N_9450,N_8044);
or U13264 (N_13264,N_8283,N_6617);
nor U13265 (N_13265,N_8500,N_9043);
and U13266 (N_13266,N_9835,N_5774);
or U13267 (N_13267,N_9837,N_9939);
nor U13268 (N_13268,N_5714,N_7044);
or U13269 (N_13269,N_6287,N_6995);
or U13270 (N_13270,N_9202,N_7502);
xor U13271 (N_13271,N_6358,N_6733);
or U13272 (N_13272,N_8325,N_5740);
nand U13273 (N_13273,N_6299,N_9397);
or U13274 (N_13274,N_8107,N_9748);
or U13275 (N_13275,N_9461,N_9545);
and U13276 (N_13276,N_9758,N_6019);
nand U13277 (N_13277,N_9860,N_5674);
and U13278 (N_13278,N_9644,N_5503);
nand U13279 (N_13279,N_5579,N_8040);
and U13280 (N_13280,N_5385,N_9237);
or U13281 (N_13281,N_8435,N_8400);
and U13282 (N_13282,N_7776,N_8927);
nand U13283 (N_13283,N_5083,N_9525);
or U13284 (N_13284,N_5383,N_6658);
nor U13285 (N_13285,N_9790,N_9906);
nor U13286 (N_13286,N_8209,N_5328);
nand U13287 (N_13287,N_6024,N_9900);
or U13288 (N_13288,N_9985,N_5334);
or U13289 (N_13289,N_5302,N_6466);
or U13290 (N_13290,N_9750,N_6826);
nor U13291 (N_13291,N_7625,N_6180);
or U13292 (N_13292,N_5527,N_5419);
nand U13293 (N_13293,N_5043,N_9163);
nand U13294 (N_13294,N_7014,N_5950);
or U13295 (N_13295,N_5405,N_5181);
nand U13296 (N_13296,N_5970,N_9030);
nor U13297 (N_13297,N_6879,N_6182);
or U13298 (N_13298,N_6361,N_8651);
or U13299 (N_13299,N_7117,N_6726);
nor U13300 (N_13300,N_8603,N_9822);
nor U13301 (N_13301,N_5975,N_5323);
nor U13302 (N_13302,N_7929,N_6517);
nor U13303 (N_13303,N_8057,N_8353);
and U13304 (N_13304,N_5205,N_5136);
nand U13305 (N_13305,N_6921,N_6082);
and U13306 (N_13306,N_7764,N_8614);
and U13307 (N_13307,N_5002,N_8796);
nand U13308 (N_13308,N_5310,N_6204);
or U13309 (N_13309,N_7818,N_8522);
or U13310 (N_13310,N_8827,N_5077);
or U13311 (N_13311,N_6570,N_9902);
or U13312 (N_13312,N_8964,N_6244);
nand U13313 (N_13313,N_5879,N_7485);
nor U13314 (N_13314,N_5501,N_6387);
or U13315 (N_13315,N_5242,N_9910);
or U13316 (N_13316,N_8606,N_9923);
nand U13317 (N_13317,N_9902,N_7922);
nand U13318 (N_13318,N_8273,N_8699);
and U13319 (N_13319,N_7614,N_5046);
and U13320 (N_13320,N_5270,N_9557);
or U13321 (N_13321,N_8482,N_6562);
nor U13322 (N_13322,N_8138,N_8310);
and U13323 (N_13323,N_5333,N_8864);
nand U13324 (N_13324,N_6620,N_5575);
nand U13325 (N_13325,N_9035,N_8577);
and U13326 (N_13326,N_8830,N_8640);
nor U13327 (N_13327,N_6104,N_7649);
nor U13328 (N_13328,N_6452,N_8985);
nand U13329 (N_13329,N_9315,N_9010);
nor U13330 (N_13330,N_8765,N_8086);
nand U13331 (N_13331,N_6103,N_6663);
or U13332 (N_13332,N_8943,N_7713);
or U13333 (N_13333,N_5999,N_9377);
and U13334 (N_13334,N_8487,N_7460);
or U13335 (N_13335,N_6414,N_6095);
nor U13336 (N_13336,N_9576,N_6174);
nor U13337 (N_13337,N_5247,N_7847);
nand U13338 (N_13338,N_6350,N_9222);
nor U13339 (N_13339,N_7836,N_7982);
nand U13340 (N_13340,N_6796,N_9584);
and U13341 (N_13341,N_6069,N_6062);
nand U13342 (N_13342,N_6789,N_5402);
and U13343 (N_13343,N_6710,N_9876);
nor U13344 (N_13344,N_6487,N_8258);
nor U13345 (N_13345,N_6258,N_5118);
nand U13346 (N_13346,N_7007,N_8481);
or U13347 (N_13347,N_6357,N_9608);
nor U13348 (N_13348,N_7234,N_9377);
nand U13349 (N_13349,N_9502,N_9997);
and U13350 (N_13350,N_7486,N_9407);
or U13351 (N_13351,N_5918,N_5075);
and U13352 (N_13352,N_8855,N_8533);
and U13353 (N_13353,N_6208,N_6344);
and U13354 (N_13354,N_7130,N_5647);
nor U13355 (N_13355,N_7564,N_7455);
or U13356 (N_13356,N_6234,N_9130);
nand U13357 (N_13357,N_7121,N_6541);
nor U13358 (N_13358,N_8031,N_8479);
and U13359 (N_13359,N_9206,N_5282);
nor U13360 (N_13360,N_5615,N_7578);
nor U13361 (N_13361,N_7128,N_8940);
or U13362 (N_13362,N_8081,N_7666);
nand U13363 (N_13363,N_9889,N_6298);
and U13364 (N_13364,N_5676,N_5718);
nor U13365 (N_13365,N_7635,N_6645);
or U13366 (N_13366,N_6404,N_6642);
nor U13367 (N_13367,N_6296,N_8805);
nand U13368 (N_13368,N_7230,N_8930);
nor U13369 (N_13369,N_7126,N_8493);
nand U13370 (N_13370,N_8517,N_9594);
and U13371 (N_13371,N_9444,N_8201);
or U13372 (N_13372,N_9546,N_8109);
and U13373 (N_13373,N_5841,N_5047);
and U13374 (N_13374,N_6404,N_5012);
and U13375 (N_13375,N_8376,N_8064);
nand U13376 (N_13376,N_6218,N_6860);
nor U13377 (N_13377,N_7166,N_6719);
or U13378 (N_13378,N_5642,N_8064);
or U13379 (N_13379,N_9324,N_5327);
nor U13380 (N_13380,N_6624,N_5661);
and U13381 (N_13381,N_7705,N_5379);
nor U13382 (N_13382,N_6185,N_8708);
nor U13383 (N_13383,N_5711,N_9532);
nand U13384 (N_13384,N_6333,N_6188);
and U13385 (N_13385,N_6613,N_9160);
and U13386 (N_13386,N_9918,N_6124);
nor U13387 (N_13387,N_7858,N_5349);
nor U13388 (N_13388,N_8722,N_9228);
nor U13389 (N_13389,N_6781,N_7781);
or U13390 (N_13390,N_6595,N_6378);
nor U13391 (N_13391,N_5414,N_8390);
nand U13392 (N_13392,N_6957,N_7964);
nand U13393 (N_13393,N_5247,N_8594);
and U13394 (N_13394,N_5098,N_7596);
and U13395 (N_13395,N_9618,N_7050);
nor U13396 (N_13396,N_6710,N_7104);
or U13397 (N_13397,N_7917,N_7286);
xor U13398 (N_13398,N_6079,N_7086);
nand U13399 (N_13399,N_7621,N_9412);
nor U13400 (N_13400,N_9301,N_9337);
or U13401 (N_13401,N_6032,N_7499);
and U13402 (N_13402,N_6782,N_8034);
or U13403 (N_13403,N_9101,N_9737);
or U13404 (N_13404,N_6495,N_7699);
or U13405 (N_13405,N_7796,N_6140);
or U13406 (N_13406,N_5600,N_6642);
nor U13407 (N_13407,N_7357,N_6178);
nor U13408 (N_13408,N_9936,N_8739);
nor U13409 (N_13409,N_9060,N_5201);
and U13410 (N_13410,N_7540,N_9410);
or U13411 (N_13411,N_8136,N_7546);
xor U13412 (N_13412,N_7236,N_5406);
nor U13413 (N_13413,N_8417,N_9166);
nand U13414 (N_13414,N_7189,N_7979);
and U13415 (N_13415,N_8208,N_8316);
nor U13416 (N_13416,N_7436,N_5504);
or U13417 (N_13417,N_6975,N_6063);
nand U13418 (N_13418,N_8265,N_9713);
nand U13419 (N_13419,N_9323,N_9379);
or U13420 (N_13420,N_6681,N_9943);
and U13421 (N_13421,N_5461,N_8233);
or U13422 (N_13422,N_5847,N_6260);
or U13423 (N_13423,N_7705,N_8171);
nand U13424 (N_13424,N_5702,N_8699);
or U13425 (N_13425,N_7926,N_7260);
nor U13426 (N_13426,N_7294,N_6967);
and U13427 (N_13427,N_8627,N_5268);
or U13428 (N_13428,N_6094,N_9608);
nand U13429 (N_13429,N_9027,N_5168);
or U13430 (N_13430,N_5255,N_7697);
or U13431 (N_13431,N_7654,N_6632);
nand U13432 (N_13432,N_5495,N_5557);
and U13433 (N_13433,N_5551,N_8235);
nor U13434 (N_13434,N_6131,N_6171);
nand U13435 (N_13435,N_6201,N_6842);
nor U13436 (N_13436,N_5898,N_6244);
and U13437 (N_13437,N_5692,N_8872);
nand U13438 (N_13438,N_7165,N_6678);
nand U13439 (N_13439,N_8364,N_5959);
nor U13440 (N_13440,N_5679,N_5407);
and U13441 (N_13441,N_5690,N_8303);
and U13442 (N_13442,N_7552,N_7930);
or U13443 (N_13443,N_9337,N_6046);
and U13444 (N_13444,N_9741,N_6830);
nand U13445 (N_13445,N_5891,N_6347);
nand U13446 (N_13446,N_6980,N_6503);
nand U13447 (N_13447,N_6740,N_7524);
nand U13448 (N_13448,N_5404,N_7140);
xnor U13449 (N_13449,N_5271,N_9964);
or U13450 (N_13450,N_9138,N_6032);
and U13451 (N_13451,N_9349,N_5593);
nor U13452 (N_13452,N_5374,N_5934);
nand U13453 (N_13453,N_7211,N_7853);
nand U13454 (N_13454,N_9013,N_9365);
nand U13455 (N_13455,N_9379,N_9733);
and U13456 (N_13456,N_6995,N_7947);
and U13457 (N_13457,N_8077,N_6025);
and U13458 (N_13458,N_8058,N_5019);
or U13459 (N_13459,N_7032,N_8429);
and U13460 (N_13460,N_9989,N_7303);
nor U13461 (N_13461,N_8704,N_6960);
nor U13462 (N_13462,N_6697,N_9198);
nand U13463 (N_13463,N_7843,N_9329);
and U13464 (N_13464,N_7749,N_9059);
and U13465 (N_13465,N_7755,N_6018);
nand U13466 (N_13466,N_9240,N_8324);
or U13467 (N_13467,N_7255,N_5917);
and U13468 (N_13468,N_6120,N_8115);
nand U13469 (N_13469,N_8206,N_9777);
nand U13470 (N_13470,N_8888,N_7424);
xor U13471 (N_13471,N_6925,N_9048);
xor U13472 (N_13472,N_8156,N_9227);
and U13473 (N_13473,N_8991,N_5847);
and U13474 (N_13474,N_8758,N_7961);
or U13475 (N_13475,N_5334,N_9685);
nor U13476 (N_13476,N_8172,N_9058);
and U13477 (N_13477,N_5973,N_6887);
nand U13478 (N_13478,N_5203,N_5837);
and U13479 (N_13479,N_9972,N_9683);
or U13480 (N_13480,N_6569,N_9049);
and U13481 (N_13481,N_8294,N_6329);
nand U13482 (N_13482,N_7821,N_5769);
nor U13483 (N_13483,N_9337,N_9625);
nand U13484 (N_13484,N_9924,N_8245);
and U13485 (N_13485,N_5304,N_8617);
nand U13486 (N_13486,N_5915,N_8269);
nor U13487 (N_13487,N_8606,N_9911);
nor U13488 (N_13488,N_5024,N_6336);
or U13489 (N_13489,N_8652,N_5417);
or U13490 (N_13490,N_6630,N_6869);
nor U13491 (N_13491,N_5320,N_6928);
nand U13492 (N_13492,N_5756,N_9117);
nand U13493 (N_13493,N_9226,N_6434);
or U13494 (N_13494,N_8965,N_7452);
and U13495 (N_13495,N_9784,N_5591);
and U13496 (N_13496,N_9393,N_8164);
or U13497 (N_13497,N_7575,N_9735);
nor U13498 (N_13498,N_8135,N_7675);
nor U13499 (N_13499,N_5490,N_7621);
and U13500 (N_13500,N_8938,N_5676);
or U13501 (N_13501,N_7177,N_6537);
and U13502 (N_13502,N_8439,N_6403);
and U13503 (N_13503,N_8614,N_6218);
and U13504 (N_13504,N_9970,N_5394);
nor U13505 (N_13505,N_6884,N_9724);
xnor U13506 (N_13506,N_7187,N_7113);
nor U13507 (N_13507,N_8731,N_6881);
or U13508 (N_13508,N_6455,N_6519);
or U13509 (N_13509,N_6832,N_5938);
and U13510 (N_13510,N_6386,N_7341);
nand U13511 (N_13511,N_5713,N_8747);
and U13512 (N_13512,N_5280,N_8542);
nand U13513 (N_13513,N_7336,N_9091);
or U13514 (N_13514,N_6367,N_7713);
or U13515 (N_13515,N_7612,N_7579);
or U13516 (N_13516,N_8545,N_5625);
or U13517 (N_13517,N_8660,N_9803);
nand U13518 (N_13518,N_6171,N_6863);
nand U13519 (N_13519,N_5150,N_9558);
and U13520 (N_13520,N_6414,N_7952);
and U13521 (N_13521,N_9861,N_8044);
or U13522 (N_13522,N_9216,N_8646);
nor U13523 (N_13523,N_7380,N_8783);
nand U13524 (N_13524,N_6031,N_5295);
nor U13525 (N_13525,N_8973,N_8228);
nor U13526 (N_13526,N_8279,N_7533);
nand U13527 (N_13527,N_6681,N_5493);
nor U13528 (N_13528,N_8956,N_9463);
or U13529 (N_13529,N_6191,N_5735);
and U13530 (N_13530,N_6684,N_7390);
nand U13531 (N_13531,N_5126,N_5650);
nand U13532 (N_13532,N_7888,N_9761);
or U13533 (N_13533,N_6577,N_6654);
or U13534 (N_13534,N_8838,N_7427);
nand U13535 (N_13535,N_7323,N_6280);
nor U13536 (N_13536,N_9257,N_9003);
or U13537 (N_13537,N_7595,N_7717);
and U13538 (N_13538,N_5140,N_5960);
nor U13539 (N_13539,N_6972,N_5606);
nor U13540 (N_13540,N_7755,N_8853);
nand U13541 (N_13541,N_6218,N_7077);
or U13542 (N_13542,N_7425,N_9036);
or U13543 (N_13543,N_7425,N_9700);
and U13544 (N_13544,N_8740,N_7802);
or U13545 (N_13545,N_6151,N_8730);
nand U13546 (N_13546,N_5937,N_6865);
and U13547 (N_13547,N_6604,N_9997);
or U13548 (N_13548,N_7370,N_7270);
and U13549 (N_13549,N_6335,N_8496);
and U13550 (N_13550,N_9358,N_5909);
or U13551 (N_13551,N_6315,N_6263);
and U13552 (N_13552,N_8360,N_6725);
xor U13553 (N_13553,N_6376,N_7668);
nor U13554 (N_13554,N_6048,N_7620);
nand U13555 (N_13555,N_7471,N_7498);
nand U13556 (N_13556,N_9814,N_5081);
nand U13557 (N_13557,N_5671,N_9013);
nor U13558 (N_13558,N_5569,N_5510);
and U13559 (N_13559,N_8775,N_7486);
or U13560 (N_13560,N_9889,N_7677);
nand U13561 (N_13561,N_9396,N_5164);
and U13562 (N_13562,N_9954,N_5160);
and U13563 (N_13563,N_6855,N_6067);
or U13564 (N_13564,N_9135,N_6464);
or U13565 (N_13565,N_9243,N_7202);
or U13566 (N_13566,N_9231,N_8255);
nor U13567 (N_13567,N_6255,N_9003);
nand U13568 (N_13568,N_6171,N_6187);
nand U13569 (N_13569,N_9280,N_8499);
or U13570 (N_13570,N_6385,N_5810);
or U13571 (N_13571,N_8615,N_5056);
or U13572 (N_13572,N_7905,N_9037);
nand U13573 (N_13573,N_7689,N_5260);
and U13574 (N_13574,N_8781,N_5686);
and U13575 (N_13575,N_5625,N_7051);
and U13576 (N_13576,N_9771,N_8115);
and U13577 (N_13577,N_5761,N_8479);
nand U13578 (N_13578,N_7046,N_9671);
nand U13579 (N_13579,N_6501,N_6024);
nand U13580 (N_13580,N_8074,N_7955);
nand U13581 (N_13581,N_9677,N_8465);
and U13582 (N_13582,N_7978,N_7812);
or U13583 (N_13583,N_6888,N_9197);
nand U13584 (N_13584,N_9291,N_9481);
or U13585 (N_13585,N_6277,N_8304);
and U13586 (N_13586,N_6975,N_8602);
nor U13587 (N_13587,N_7883,N_6542);
nand U13588 (N_13588,N_9826,N_7442);
and U13589 (N_13589,N_7059,N_9600);
nor U13590 (N_13590,N_5274,N_5980);
nor U13591 (N_13591,N_7703,N_7142);
or U13592 (N_13592,N_8284,N_8242);
and U13593 (N_13593,N_8055,N_5010);
nor U13594 (N_13594,N_9066,N_5446);
nor U13595 (N_13595,N_8531,N_7233);
nor U13596 (N_13596,N_7896,N_6719);
and U13597 (N_13597,N_9127,N_6787);
or U13598 (N_13598,N_7731,N_9835);
or U13599 (N_13599,N_8648,N_8676);
nand U13600 (N_13600,N_7326,N_9036);
nor U13601 (N_13601,N_5023,N_7428);
nor U13602 (N_13602,N_8870,N_6885);
and U13603 (N_13603,N_5661,N_9255);
nand U13604 (N_13604,N_5684,N_8413);
nand U13605 (N_13605,N_6709,N_8426);
nand U13606 (N_13606,N_5986,N_7402);
nor U13607 (N_13607,N_5381,N_5864);
and U13608 (N_13608,N_9856,N_7620);
nor U13609 (N_13609,N_6181,N_8433);
nand U13610 (N_13610,N_7120,N_5752);
nand U13611 (N_13611,N_8815,N_7218);
and U13612 (N_13612,N_8583,N_6141);
and U13613 (N_13613,N_8963,N_5511);
nor U13614 (N_13614,N_5162,N_6687);
nand U13615 (N_13615,N_6197,N_6761);
nand U13616 (N_13616,N_5498,N_7049);
nand U13617 (N_13617,N_8727,N_7842);
nor U13618 (N_13618,N_5194,N_6533);
and U13619 (N_13619,N_8978,N_8995);
or U13620 (N_13620,N_6896,N_8943);
or U13621 (N_13621,N_5895,N_7986);
or U13622 (N_13622,N_7957,N_5531);
nor U13623 (N_13623,N_7936,N_9886);
and U13624 (N_13624,N_7112,N_8970);
nor U13625 (N_13625,N_7064,N_9119);
and U13626 (N_13626,N_6206,N_8817);
nand U13627 (N_13627,N_9233,N_6387);
and U13628 (N_13628,N_9332,N_9822);
nand U13629 (N_13629,N_7372,N_5111);
or U13630 (N_13630,N_5874,N_8175);
and U13631 (N_13631,N_8525,N_7588);
nor U13632 (N_13632,N_9459,N_5012);
and U13633 (N_13633,N_9091,N_9655);
nand U13634 (N_13634,N_5336,N_9400);
or U13635 (N_13635,N_6760,N_5076);
nand U13636 (N_13636,N_9511,N_8666);
nor U13637 (N_13637,N_8084,N_7832);
or U13638 (N_13638,N_7072,N_8260);
nand U13639 (N_13639,N_7738,N_8414);
nor U13640 (N_13640,N_8144,N_5753);
nand U13641 (N_13641,N_6184,N_5883);
and U13642 (N_13642,N_8238,N_8602);
nand U13643 (N_13643,N_9882,N_6505);
or U13644 (N_13644,N_6419,N_7411);
nand U13645 (N_13645,N_9922,N_9081);
and U13646 (N_13646,N_9918,N_7394);
nand U13647 (N_13647,N_8157,N_7968);
and U13648 (N_13648,N_8526,N_7447);
nand U13649 (N_13649,N_9365,N_7215);
and U13650 (N_13650,N_5349,N_8518);
nand U13651 (N_13651,N_9443,N_8737);
nand U13652 (N_13652,N_9796,N_9756);
or U13653 (N_13653,N_8494,N_5398);
or U13654 (N_13654,N_6122,N_5638);
nand U13655 (N_13655,N_9454,N_7001);
nor U13656 (N_13656,N_5051,N_8417);
nor U13657 (N_13657,N_9554,N_6405);
nor U13658 (N_13658,N_6737,N_7625);
or U13659 (N_13659,N_8907,N_8583);
and U13660 (N_13660,N_8520,N_6640);
nor U13661 (N_13661,N_7001,N_5101);
and U13662 (N_13662,N_5699,N_6991);
nor U13663 (N_13663,N_6098,N_5731);
nand U13664 (N_13664,N_8059,N_5705);
or U13665 (N_13665,N_8906,N_7490);
or U13666 (N_13666,N_6667,N_5288);
nand U13667 (N_13667,N_9641,N_5314);
or U13668 (N_13668,N_7534,N_5234);
nand U13669 (N_13669,N_6442,N_8594);
nand U13670 (N_13670,N_6631,N_5660);
nor U13671 (N_13671,N_6597,N_9061);
nand U13672 (N_13672,N_5324,N_7246);
nand U13673 (N_13673,N_8802,N_9963);
nor U13674 (N_13674,N_7714,N_6272);
xnor U13675 (N_13675,N_7809,N_8816);
nor U13676 (N_13676,N_7538,N_8674);
or U13677 (N_13677,N_6089,N_5857);
nand U13678 (N_13678,N_5878,N_7892);
nor U13679 (N_13679,N_7799,N_6485);
or U13680 (N_13680,N_7543,N_6398);
and U13681 (N_13681,N_8702,N_8374);
or U13682 (N_13682,N_9834,N_5721);
or U13683 (N_13683,N_8278,N_6577);
nand U13684 (N_13684,N_8264,N_8796);
and U13685 (N_13685,N_8203,N_7608);
nand U13686 (N_13686,N_9433,N_7082);
or U13687 (N_13687,N_7147,N_9472);
or U13688 (N_13688,N_5120,N_8079);
nor U13689 (N_13689,N_8849,N_5924);
or U13690 (N_13690,N_7283,N_9699);
or U13691 (N_13691,N_5093,N_5561);
nand U13692 (N_13692,N_7794,N_6538);
nand U13693 (N_13693,N_8851,N_6077);
or U13694 (N_13694,N_9428,N_6274);
and U13695 (N_13695,N_9143,N_6774);
or U13696 (N_13696,N_7102,N_9920);
or U13697 (N_13697,N_5718,N_8012);
or U13698 (N_13698,N_8012,N_7608);
and U13699 (N_13699,N_6375,N_8596);
and U13700 (N_13700,N_8059,N_8863);
nor U13701 (N_13701,N_6050,N_7333);
or U13702 (N_13702,N_8059,N_8570);
nor U13703 (N_13703,N_5347,N_7942);
nand U13704 (N_13704,N_7259,N_7150);
or U13705 (N_13705,N_8305,N_8924);
nand U13706 (N_13706,N_5271,N_7786);
and U13707 (N_13707,N_9120,N_7198);
or U13708 (N_13708,N_5670,N_7962);
nor U13709 (N_13709,N_9945,N_9168);
nand U13710 (N_13710,N_6212,N_7368);
or U13711 (N_13711,N_6491,N_8774);
or U13712 (N_13712,N_6327,N_9340);
nor U13713 (N_13713,N_5797,N_6735);
and U13714 (N_13714,N_6911,N_7743);
and U13715 (N_13715,N_5084,N_5810);
and U13716 (N_13716,N_6144,N_6130);
nor U13717 (N_13717,N_7290,N_5177);
nand U13718 (N_13718,N_5403,N_8471);
nand U13719 (N_13719,N_6237,N_7997);
nor U13720 (N_13720,N_8442,N_9505);
nand U13721 (N_13721,N_7812,N_5246);
and U13722 (N_13722,N_8652,N_8658);
and U13723 (N_13723,N_5813,N_9288);
or U13724 (N_13724,N_6214,N_9387);
nor U13725 (N_13725,N_9486,N_5287);
nor U13726 (N_13726,N_6111,N_7327);
nor U13727 (N_13727,N_9756,N_7604);
or U13728 (N_13728,N_6270,N_6279);
nand U13729 (N_13729,N_5940,N_6493);
nor U13730 (N_13730,N_6759,N_9377);
and U13731 (N_13731,N_9871,N_6951);
nand U13732 (N_13732,N_6729,N_6057);
nand U13733 (N_13733,N_5930,N_6914);
nor U13734 (N_13734,N_6615,N_5406);
and U13735 (N_13735,N_9075,N_6482);
and U13736 (N_13736,N_6962,N_5634);
nand U13737 (N_13737,N_8521,N_6103);
and U13738 (N_13738,N_5010,N_5178);
nand U13739 (N_13739,N_7281,N_7130);
nor U13740 (N_13740,N_6601,N_5457);
or U13741 (N_13741,N_5005,N_6513);
or U13742 (N_13742,N_7716,N_7486);
or U13743 (N_13743,N_9907,N_7897);
nand U13744 (N_13744,N_8306,N_6692);
nor U13745 (N_13745,N_7909,N_9145);
nor U13746 (N_13746,N_9285,N_7854);
nor U13747 (N_13747,N_8895,N_5329);
nand U13748 (N_13748,N_6385,N_6997);
and U13749 (N_13749,N_6040,N_6983);
and U13750 (N_13750,N_7042,N_7129);
or U13751 (N_13751,N_7580,N_9304);
or U13752 (N_13752,N_5049,N_9108);
and U13753 (N_13753,N_7988,N_6610);
nand U13754 (N_13754,N_6435,N_5869);
or U13755 (N_13755,N_6416,N_7557);
nor U13756 (N_13756,N_6739,N_7260);
and U13757 (N_13757,N_8188,N_9686);
and U13758 (N_13758,N_6939,N_7068);
nand U13759 (N_13759,N_7051,N_6777);
and U13760 (N_13760,N_6252,N_8610);
nor U13761 (N_13761,N_9741,N_6188);
nand U13762 (N_13762,N_6006,N_7351);
or U13763 (N_13763,N_6212,N_8230);
nor U13764 (N_13764,N_9760,N_5136);
nor U13765 (N_13765,N_6440,N_7124);
and U13766 (N_13766,N_8021,N_9248);
or U13767 (N_13767,N_7642,N_6332);
nor U13768 (N_13768,N_6339,N_8246);
and U13769 (N_13769,N_7130,N_8806);
or U13770 (N_13770,N_5733,N_8376);
and U13771 (N_13771,N_8338,N_8459);
or U13772 (N_13772,N_5009,N_8258);
or U13773 (N_13773,N_6097,N_7569);
and U13774 (N_13774,N_8943,N_5433);
or U13775 (N_13775,N_9508,N_8771);
nand U13776 (N_13776,N_7286,N_8457);
or U13777 (N_13777,N_9456,N_6972);
nand U13778 (N_13778,N_5598,N_7670);
nand U13779 (N_13779,N_8729,N_6219);
nand U13780 (N_13780,N_5896,N_8941);
and U13781 (N_13781,N_5788,N_7625);
xor U13782 (N_13782,N_6879,N_8124);
nand U13783 (N_13783,N_6873,N_6187);
and U13784 (N_13784,N_7039,N_5199);
nand U13785 (N_13785,N_8857,N_5596);
nand U13786 (N_13786,N_9243,N_8957);
nand U13787 (N_13787,N_9683,N_8893);
or U13788 (N_13788,N_5703,N_9641);
and U13789 (N_13789,N_7659,N_5176);
or U13790 (N_13790,N_6724,N_9853);
nor U13791 (N_13791,N_7598,N_9574);
nor U13792 (N_13792,N_6797,N_7085);
nand U13793 (N_13793,N_5485,N_8847);
or U13794 (N_13794,N_6942,N_7451);
nand U13795 (N_13795,N_6321,N_7909);
nor U13796 (N_13796,N_8537,N_8776);
or U13797 (N_13797,N_6426,N_9212);
or U13798 (N_13798,N_7586,N_5423);
and U13799 (N_13799,N_9652,N_5931);
nand U13800 (N_13800,N_9924,N_8363);
nand U13801 (N_13801,N_7701,N_7111);
nand U13802 (N_13802,N_9840,N_8857);
nor U13803 (N_13803,N_5431,N_6939);
or U13804 (N_13804,N_5520,N_6574);
nor U13805 (N_13805,N_7802,N_5331);
nor U13806 (N_13806,N_7743,N_8973);
and U13807 (N_13807,N_9382,N_8160);
nand U13808 (N_13808,N_8207,N_7212);
and U13809 (N_13809,N_5168,N_7087);
or U13810 (N_13810,N_7379,N_5621);
or U13811 (N_13811,N_9076,N_6505);
or U13812 (N_13812,N_5901,N_9092);
nand U13813 (N_13813,N_7223,N_7714);
nand U13814 (N_13814,N_9128,N_9536);
and U13815 (N_13815,N_6444,N_7190);
nand U13816 (N_13816,N_7486,N_8089);
nor U13817 (N_13817,N_5041,N_5529);
nand U13818 (N_13818,N_7630,N_9336);
and U13819 (N_13819,N_5396,N_5576);
nand U13820 (N_13820,N_6849,N_9614);
nor U13821 (N_13821,N_6792,N_6442);
nand U13822 (N_13822,N_5843,N_5213);
or U13823 (N_13823,N_7382,N_9532);
nand U13824 (N_13824,N_6015,N_7405);
nand U13825 (N_13825,N_8913,N_8633);
and U13826 (N_13826,N_5532,N_7365);
and U13827 (N_13827,N_8292,N_8205);
and U13828 (N_13828,N_6489,N_7165);
nor U13829 (N_13829,N_8931,N_7562);
or U13830 (N_13830,N_7436,N_9648);
nor U13831 (N_13831,N_9565,N_5827);
nand U13832 (N_13832,N_6933,N_5258);
or U13833 (N_13833,N_8700,N_5052);
or U13834 (N_13834,N_6856,N_9826);
and U13835 (N_13835,N_9772,N_9180);
nor U13836 (N_13836,N_8557,N_9641);
and U13837 (N_13837,N_9612,N_7466);
or U13838 (N_13838,N_6764,N_5521);
nor U13839 (N_13839,N_7065,N_7417);
nand U13840 (N_13840,N_5227,N_6622);
or U13841 (N_13841,N_8702,N_9432);
and U13842 (N_13842,N_7740,N_9451);
and U13843 (N_13843,N_7914,N_5152);
or U13844 (N_13844,N_8359,N_6197);
and U13845 (N_13845,N_8257,N_8092);
nand U13846 (N_13846,N_8035,N_7774);
or U13847 (N_13847,N_8321,N_5281);
or U13848 (N_13848,N_5003,N_7990);
nand U13849 (N_13849,N_9896,N_8830);
or U13850 (N_13850,N_8348,N_7391);
or U13851 (N_13851,N_5118,N_5826);
or U13852 (N_13852,N_7764,N_6506);
and U13853 (N_13853,N_6512,N_8534);
and U13854 (N_13854,N_8976,N_5801);
nor U13855 (N_13855,N_9895,N_8711);
nand U13856 (N_13856,N_8847,N_8019);
or U13857 (N_13857,N_7455,N_9269);
nand U13858 (N_13858,N_8552,N_7182);
nand U13859 (N_13859,N_8877,N_6420);
or U13860 (N_13860,N_7819,N_6928);
and U13861 (N_13861,N_9005,N_8152);
nor U13862 (N_13862,N_7749,N_5224);
nor U13863 (N_13863,N_7472,N_5158);
nand U13864 (N_13864,N_6823,N_9476);
and U13865 (N_13865,N_9489,N_5552);
nand U13866 (N_13866,N_6379,N_7647);
nor U13867 (N_13867,N_9331,N_7708);
nand U13868 (N_13868,N_8917,N_9197);
nand U13869 (N_13869,N_6765,N_8127);
nor U13870 (N_13870,N_6758,N_8514);
or U13871 (N_13871,N_6194,N_7860);
nor U13872 (N_13872,N_9227,N_9426);
and U13873 (N_13873,N_6158,N_7032);
nor U13874 (N_13874,N_8846,N_7996);
nor U13875 (N_13875,N_7354,N_5827);
or U13876 (N_13876,N_5496,N_8193);
and U13877 (N_13877,N_5462,N_5849);
or U13878 (N_13878,N_7200,N_6062);
and U13879 (N_13879,N_8141,N_8564);
and U13880 (N_13880,N_7084,N_5018);
nor U13881 (N_13881,N_8915,N_5201);
nor U13882 (N_13882,N_7757,N_8990);
and U13883 (N_13883,N_9303,N_7561);
nand U13884 (N_13884,N_9420,N_5243);
or U13885 (N_13885,N_8015,N_7739);
or U13886 (N_13886,N_5735,N_6285);
nor U13887 (N_13887,N_8138,N_7404);
nand U13888 (N_13888,N_9816,N_9942);
or U13889 (N_13889,N_6956,N_9967);
nand U13890 (N_13890,N_8761,N_6597);
nand U13891 (N_13891,N_6200,N_8266);
nand U13892 (N_13892,N_6739,N_6111);
nand U13893 (N_13893,N_7933,N_6307);
nand U13894 (N_13894,N_7159,N_5675);
nand U13895 (N_13895,N_9015,N_5331);
nand U13896 (N_13896,N_9084,N_8362);
and U13897 (N_13897,N_9564,N_9524);
or U13898 (N_13898,N_6245,N_9914);
nand U13899 (N_13899,N_8354,N_5301);
or U13900 (N_13900,N_9177,N_9540);
and U13901 (N_13901,N_9070,N_9773);
nor U13902 (N_13902,N_8397,N_6838);
or U13903 (N_13903,N_9625,N_7486);
nor U13904 (N_13904,N_9987,N_7020);
or U13905 (N_13905,N_7923,N_8638);
nand U13906 (N_13906,N_6407,N_6664);
nand U13907 (N_13907,N_9139,N_6818);
and U13908 (N_13908,N_8970,N_8287);
nor U13909 (N_13909,N_8456,N_7582);
or U13910 (N_13910,N_7458,N_6808);
or U13911 (N_13911,N_8787,N_8452);
nor U13912 (N_13912,N_7932,N_9782);
or U13913 (N_13913,N_6962,N_7899);
or U13914 (N_13914,N_6555,N_5457);
nand U13915 (N_13915,N_9921,N_8908);
nand U13916 (N_13916,N_9936,N_5816);
nand U13917 (N_13917,N_9202,N_7460);
or U13918 (N_13918,N_9004,N_7626);
nand U13919 (N_13919,N_8973,N_7575);
nor U13920 (N_13920,N_6173,N_5731);
nor U13921 (N_13921,N_8375,N_5317);
or U13922 (N_13922,N_7487,N_6555);
and U13923 (N_13923,N_8832,N_7062);
nand U13924 (N_13924,N_6378,N_7762);
or U13925 (N_13925,N_9739,N_6753);
or U13926 (N_13926,N_7165,N_5969);
nand U13927 (N_13927,N_8668,N_9087);
nor U13928 (N_13928,N_9180,N_9711);
nor U13929 (N_13929,N_5088,N_6668);
and U13930 (N_13930,N_8638,N_8209);
and U13931 (N_13931,N_6577,N_7935);
nand U13932 (N_13932,N_8766,N_8551);
or U13933 (N_13933,N_9166,N_5163);
nor U13934 (N_13934,N_5129,N_7030);
and U13935 (N_13935,N_7390,N_6625);
or U13936 (N_13936,N_8224,N_6000);
and U13937 (N_13937,N_5017,N_8098);
nor U13938 (N_13938,N_9088,N_8525);
and U13939 (N_13939,N_7446,N_7062);
nand U13940 (N_13940,N_9009,N_9399);
or U13941 (N_13941,N_5885,N_5839);
or U13942 (N_13942,N_8315,N_7242);
nand U13943 (N_13943,N_9956,N_6695);
and U13944 (N_13944,N_7779,N_6087);
nand U13945 (N_13945,N_5781,N_8676);
nor U13946 (N_13946,N_9174,N_9228);
nand U13947 (N_13947,N_8167,N_5783);
nor U13948 (N_13948,N_6401,N_9284);
and U13949 (N_13949,N_9136,N_6631);
and U13950 (N_13950,N_8026,N_8239);
or U13951 (N_13951,N_6937,N_7252);
and U13952 (N_13952,N_8210,N_8989);
xnor U13953 (N_13953,N_8912,N_7079);
nor U13954 (N_13954,N_7999,N_8551);
nand U13955 (N_13955,N_5517,N_7674);
and U13956 (N_13956,N_5016,N_8429);
or U13957 (N_13957,N_9204,N_5563);
or U13958 (N_13958,N_7731,N_5508);
nor U13959 (N_13959,N_9510,N_7946);
nor U13960 (N_13960,N_8696,N_5773);
nor U13961 (N_13961,N_9027,N_6737);
nor U13962 (N_13962,N_9260,N_5566);
or U13963 (N_13963,N_8405,N_5791);
and U13964 (N_13964,N_6020,N_5908);
nor U13965 (N_13965,N_7130,N_5672);
and U13966 (N_13966,N_7756,N_6280);
or U13967 (N_13967,N_7925,N_9397);
and U13968 (N_13968,N_6237,N_8424);
or U13969 (N_13969,N_8997,N_7345);
xor U13970 (N_13970,N_6183,N_7644);
or U13971 (N_13971,N_5479,N_5150);
nor U13972 (N_13972,N_8511,N_6307);
nand U13973 (N_13973,N_6373,N_9756);
nand U13974 (N_13974,N_7003,N_7267);
nor U13975 (N_13975,N_8701,N_7695);
and U13976 (N_13976,N_9917,N_6186);
nand U13977 (N_13977,N_6270,N_7225);
nor U13978 (N_13978,N_8667,N_5873);
and U13979 (N_13979,N_8057,N_5271);
nor U13980 (N_13980,N_6577,N_5270);
nor U13981 (N_13981,N_5252,N_5225);
nand U13982 (N_13982,N_5670,N_8095);
nand U13983 (N_13983,N_8038,N_7885);
or U13984 (N_13984,N_7599,N_7122);
and U13985 (N_13985,N_7701,N_7831);
nand U13986 (N_13986,N_6112,N_6708);
and U13987 (N_13987,N_6006,N_9820);
or U13988 (N_13988,N_5230,N_9632);
and U13989 (N_13989,N_7368,N_5224);
nor U13990 (N_13990,N_8986,N_7364);
nor U13991 (N_13991,N_9031,N_7884);
or U13992 (N_13992,N_5937,N_8514);
or U13993 (N_13993,N_5836,N_7171);
nand U13994 (N_13994,N_6943,N_6007);
or U13995 (N_13995,N_5594,N_7798);
or U13996 (N_13996,N_5164,N_9401);
or U13997 (N_13997,N_7896,N_8169);
and U13998 (N_13998,N_7392,N_5475);
nor U13999 (N_13999,N_6877,N_9089);
nor U14000 (N_14000,N_5486,N_9864);
nand U14001 (N_14001,N_7974,N_9909);
nor U14002 (N_14002,N_8874,N_7133);
nor U14003 (N_14003,N_8821,N_7531);
xor U14004 (N_14004,N_9424,N_6597);
nand U14005 (N_14005,N_9187,N_8641);
or U14006 (N_14006,N_8088,N_9265);
nor U14007 (N_14007,N_7655,N_6913);
and U14008 (N_14008,N_6565,N_9828);
nand U14009 (N_14009,N_6396,N_5186);
nor U14010 (N_14010,N_6994,N_7149);
and U14011 (N_14011,N_7393,N_5606);
and U14012 (N_14012,N_9875,N_5929);
nor U14013 (N_14013,N_6814,N_8234);
or U14014 (N_14014,N_6283,N_6323);
or U14015 (N_14015,N_7706,N_5852);
and U14016 (N_14016,N_6072,N_6440);
nor U14017 (N_14017,N_6411,N_6854);
or U14018 (N_14018,N_9175,N_6045);
or U14019 (N_14019,N_7347,N_8861);
and U14020 (N_14020,N_6391,N_8689);
nand U14021 (N_14021,N_5868,N_6198);
nand U14022 (N_14022,N_9127,N_9128);
or U14023 (N_14023,N_9832,N_7735);
and U14024 (N_14024,N_8808,N_8564);
or U14025 (N_14025,N_9285,N_6342);
nor U14026 (N_14026,N_6690,N_5218);
nor U14027 (N_14027,N_8959,N_6782);
or U14028 (N_14028,N_6553,N_9760);
or U14029 (N_14029,N_9269,N_7595);
and U14030 (N_14030,N_9657,N_5198);
nand U14031 (N_14031,N_9842,N_5831);
and U14032 (N_14032,N_9394,N_6732);
or U14033 (N_14033,N_7449,N_8222);
or U14034 (N_14034,N_6272,N_5298);
nor U14035 (N_14035,N_8746,N_8274);
nand U14036 (N_14036,N_7431,N_5831);
or U14037 (N_14037,N_7339,N_7194);
nand U14038 (N_14038,N_6320,N_5441);
nor U14039 (N_14039,N_6051,N_6488);
nand U14040 (N_14040,N_6927,N_5106);
xor U14041 (N_14041,N_6629,N_6350);
or U14042 (N_14042,N_8579,N_6133);
and U14043 (N_14043,N_6349,N_9895);
or U14044 (N_14044,N_9749,N_5153);
and U14045 (N_14045,N_5060,N_7012);
nand U14046 (N_14046,N_5346,N_6884);
nand U14047 (N_14047,N_7798,N_5364);
and U14048 (N_14048,N_6640,N_9146);
and U14049 (N_14049,N_8481,N_7814);
nor U14050 (N_14050,N_8905,N_6933);
nor U14051 (N_14051,N_8350,N_6342);
or U14052 (N_14052,N_8065,N_8015);
xor U14053 (N_14053,N_6205,N_8313);
nand U14054 (N_14054,N_6854,N_6155);
nand U14055 (N_14055,N_7852,N_8161);
and U14056 (N_14056,N_6852,N_5075);
nand U14057 (N_14057,N_6747,N_5587);
nor U14058 (N_14058,N_6290,N_7589);
or U14059 (N_14059,N_9902,N_8736);
and U14060 (N_14060,N_9995,N_6311);
and U14061 (N_14061,N_8653,N_7761);
and U14062 (N_14062,N_7845,N_6584);
and U14063 (N_14063,N_6769,N_7226);
nand U14064 (N_14064,N_8202,N_9257);
nand U14065 (N_14065,N_7686,N_7859);
and U14066 (N_14066,N_6813,N_6619);
or U14067 (N_14067,N_7387,N_9328);
nand U14068 (N_14068,N_8448,N_9273);
and U14069 (N_14069,N_9674,N_7896);
and U14070 (N_14070,N_8355,N_7103);
nor U14071 (N_14071,N_5870,N_6726);
nor U14072 (N_14072,N_8470,N_7454);
and U14073 (N_14073,N_6281,N_9320);
nand U14074 (N_14074,N_9294,N_9142);
nor U14075 (N_14075,N_7963,N_8027);
or U14076 (N_14076,N_9499,N_9065);
nand U14077 (N_14077,N_9482,N_7024);
nand U14078 (N_14078,N_8469,N_7219);
and U14079 (N_14079,N_7768,N_9909);
or U14080 (N_14080,N_5606,N_6673);
nand U14081 (N_14081,N_6050,N_7589);
nor U14082 (N_14082,N_8394,N_6817);
and U14083 (N_14083,N_8223,N_5395);
nand U14084 (N_14084,N_8016,N_9214);
nand U14085 (N_14085,N_6940,N_9428);
nor U14086 (N_14086,N_9201,N_6746);
nand U14087 (N_14087,N_7743,N_5541);
nor U14088 (N_14088,N_9775,N_6559);
and U14089 (N_14089,N_9291,N_7466);
or U14090 (N_14090,N_8996,N_6553);
nor U14091 (N_14091,N_8213,N_8080);
nor U14092 (N_14092,N_5275,N_9140);
nor U14093 (N_14093,N_7141,N_5053);
and U14094 (N_14094,N_5284,N_7488);
and U14095 (N_14095,N_7091,N_7394);
and U14096 (N_14096,N_7429,N_6725);
and U14097 (N_14097,N_5006,N_7399);
nand U14098 (N_14098,N_8139,N_6977);
nand U14099 (N_14099,N_5776,N_6228);
or U14100 (N_14100,N_5045,N_9007);
nor U14101 (N_14101,N_6287,N_8630);
or U14102 (N_14102,N_5596,N_9536);
nor U14103 (N_14103,N_8556,N_8671);
and U14104 (N_14104,N_7551,N_5300);
or U14105 (N_14105,N_5579,N_7659);
and U14106 (N_14106,N_9229,N_6144);
and U14107 (N_14107,N_6982,N_5085);
nor U14108 (N_14108,N_7087,N_6856);
nand U14109 (N_14109,N_6076,N_5603);
or U14110 (N_14110,N_8891,N_5343);
or U14111 (N_14111,N_6991,N_7757);
or U14112 (N_14112,N_5423,N_5955);
nand U14113 (N_14113,N_9830,N_9667);
nor U14114 (N_14114,N_6583,N_6522);
nand U14115 (N_14115,N_9433,N_6851);
nor U14116 (N_14116,N_9385,N_9862);
nand U14117 (N_14117,N_5882,N_9188);
nand U14118 (N_14118,N_9133,N_9530);
nor U14119 (N_14119,N_8312,N_5723);
and U14120 (N_14120,N_6965,N_7995);
and U14121 (N_14121,N_8090,N_5392);
nand U14122 (N_14122,N_7475,N_8303);
nor U14123 (N_14123,N_8579,N_9163);
and U14124 (N_14124,N_5504,N_7782);
or U14125 (N_14125,N_7993,N_5587);
and U14126 (N_14126,N_5606,N_5164);
or U14127 (N_14127,N_7023,N_6451);
nand U14128 (N_14128,N_8744,N_9352);
and U14129 (N_14129,N_9588,N_8693);
or U14130 (N_14130,N_6162,N_6094);
and U14131 (N_14131,N_9705,N_8821);
or U14132 (N_14132,N_5126,N_8378);
and U14133 (N_14133,N_5511,N_6241);
nand U14134 (N_14134,N_5508,N_8505);
nand U14135 (N_14135,N_6654,N_5427);
nand U14136 (N_14136,N_8448,N_9055);
and U14137 (N_14137,N_9546,N_9559);
and U14138 (N_14138,N_6744,N_8941);
nand U14139 (N_14139,N_8094,N_6266);
nor U14140 (N_14140,N_8178,N_9665);
nor U14141 (N_14141,N_7798,N_5979);
nand U14142 (N_14142,N_7315,N_5235);
nor U14143 (N_14143,N_8311,N_5155);
or U14144 (N_14144,N_8524,N_7395);
nand U14145 (N_14145,N_5640,N_9783);
and U14146 (N_14146,N_9840,N_9454);
and U14147 (N_14147,N_6247,N_5087);
or U14148 (N_14148,N_8336,N_8435);
or U14149 (N_14149,N_5456,N_9465);
nand U14150 (N_14150,N_8118,N_9491);
or U14151 (N_14151,N_8248,N_9613);
nand U14152 (N_14152,N_7335,N_6086);
or U14153 (N_14153,N_8832,N_6639);
and U14154 (N_14154,N_8612,N_5383);
and U14155 (N_14155,N_5548,N_6409);
nand U14156 (N_14156,N_8904,N_7441);
nand U14157 (N_14157,N_5653,N_5619);
nand U14158 (N_14158,N_9307,N_7374);
nor U14159 (N_14159,N_5266,N_9215);
nand U14160 (N_14160,N_8785,N_6579);
or U14161 (N_14161,N_8405,N_6703);
and U14162 (N_14162,N_5765,N_7647);
nor U14163 (N_14163,N_8270,N_6611);
or U14164 (N_14164,N_9556,N_7707);
and U14165 (N_14165,N_7365,N_9206);
nor U14166 (N_14166,N_7381,N_7939);
nand U14167 (N_14167,N_7898,N_7700);
and U14168 (N_14168,N_6979,N_5665);
nand U14169 (N_14169,N_5381,N_8016);
and U14170 (N_14170,N_6086,N_8455);
or U14171 (N_14171,N_9044,N_7655);
nor U14172 (N_14172,N_8353,N_7352);
nand U14173 (N_14173,N_6084,N_5960);
and U14174 (N_14174,N_9063,N_7248);
and U14175 (N_14175,N_7909,N_6229);
or U14176 (N_14176,N_8260,N_6123);
nand U14177 (N_14177,N_6249,N_8182);
nand U14178 (N_14178,N_6358,N_6888);
and U14179 (N_14179,N_7202,N_8098);
or U14180 (N_14180,N_6825,N_8250);
and U14181 (N_14181,N_7161,N_7859);
nand U14182 (N_14182,N_7940,N_9135);
and U14183 (N_14183,N_8009,N_6494);
nand U14184 (N_14184,N_8550,N_5164);
nor U14185 (N_14185,N_9964,N_9407);
or U14186 (N_14186,N_5729,N_7574);
or U14187 (N_14187,N_5736,N_9149);
and U14188 (N_14188,N_5432,N_8024);
nor U14189 (N_14189,N_8675,N_6217);
or U14190 (N_14190,N_9488,N_5525);
nand U14191 (N_14191,N_9633,N_6587);
or U14192 (N_14192,N_6469,N_5924);
or U14193 (N_14193,N_7295,N_7422);
or U14194 (N_14194,N_8316,N_8210);
and U14195 (N_14195,N_8771,N_6122);
or U14196 (N_14196,N_8513,N_6777);
or U14197 (N_14197,N_5536,N_9938);
and U14198 (N_14198,N_8562,N_8097);
nor U14199 (N_14199,N_7081,N_6750);
or U14200 (N_14200,N_6855,N_6998);
nor U14201 (N_14201,N_5373,N_7927);
nor U14202 (N_14202,N_9872,N_7490);
nand U14203 (N_14203,N_6616,N_6513);
nand U14204 (N_14204,N_5462,N_8646);
nand U14205 (N_14205,N_7734,N_6962);
and U14206 (N_14206,N_7054,N_7533);
nand U14207 (N_14207,N_8917,N_8654);
or U14208 (N_14208,N_6124,N_5402);
nand U14209 (N_14209,N_5609,N_5039);
nor U14210 (N_14210,N_8859,N_5628);
nand U14211 (N_14211,N_8141,N_7412);
or U14212 (N_14212,N_9505,N_7097);
or U14213 (N_14213,N_6924,N_6530);
xor U14214 (N_14214,N_8383,N_6632);
nor U14215 (N_14215,N_8176,N_5455);
or U14216 (N_14216,N_8286,N_7458);
nand U14217 (N_14217,N_7503,N_9896);
and U14218 (N_14218,N_7287,N_6196);
and U14219 (N_14219,N_5552,N_6726);
or U14220 (N_14220,N_5193,N_8452);
nor U14221 (N_14221,N_8195,N_5762);
or U14222 (N_14222,N_5086,N_9985);
or U14223 (N_14223,N_9308,N_6480);
nor U14224 (N_14224,N_7901,N_6818);
nor U14225 (N_14225,N_5674,N_5870);
nand U14226 (N_14226,N_6866,N_5475);
or U14227 (N_14227,N_5187,N_5580);
nor U14228 (N_14228,N_5174,N_9699);
and U14229 (N_14229,N_5175,N_9847);
or U14230 (N_14230,N_5090,N_8430);
and U14231 (N_14231,N_5443,N_9612);
and U14232 (N_14232,N_7037,N_7647);
nand U14233 (N_14233,N_8128,N_6390);
nand U14234 (N_14234,N_7236,N_9465);
or U14235 (N_14235,N_8477,N_6856);
and U14236 (N_14236,N_9921,N_6980);
nor U14237 (N_14237,N_7817,N_5755);
nor U14238 (N_14238,N_8524,N_7820);
nand U14239 (N_14239,N_9676,N_8069);
and U14240 (N_14240,N_5981,N_6475);
and U14241 (N_14241,N_8051,N_6254);
nand U14242 (N_14242,N_5930,N_7468);
or U14243 (N_14243,N_8184,N_5732);
or U14244 (N_14244,N_6682,N_5764);
nor U14245 (N_14245,N_7371,N_7272);
nand U14246 (N_14246,N_6025,N_5028);
or U14247 (N_14247,N_6671,N_8528);
and U14248 (N_14248,N_6740,N_9951);
nor U14249 (N_14249,N_9642,N_9781);
nand U14250 (N_14250,N_5967,N_9852);
and U14251 (N_14251,N_8490,N_8245);
nand U14252 (N_14252,N_8067,N_9030);
nor U14253 (N_14253,N_8029,N_9747);
or U14254 (N_14254,N_9973,N_6673);
nand U14255 (N_14255,N_6971,N_9061);
or U14256 (N_14256,N_5175,N_8604);
nand U14257 (N_14257,N_7493,N_9607);
nand U14258 (N_14258,N_8211,N_6770);
nand U14259 (N_14259,N_5375,N_9025);
and U14260 (N_14260,N_6328,N_7895);
or U14261 (N_14261,N_6868,N_7625);
and U14262 (N_14262,N_5354,N_8646);
or U14263 (N_14263,N_7473,N_6710);
nand U14264 (N_14264,N_8945,N_5484);
nand U14265 (N_14265,N_6959,N_7558);
or U14266 (N_14266,N_5738,N_7983);
and U14267 (N_14267,N_6141,N_6747);
or U14268 (N_14268,N_6812,N_9697);
nor U14269 (N_14269,N_8488,N_8055);
nor U14270 (N_14270,N_9640,N_7021);
or U14271 (N_14271,N_9860,N_9916);
nand U14272 (N_14272,N_9184,N_7930);
and U14273 (N_14273,N_8433,N_6430);
and U14274 (N_14274,N_9228,N_5663);
and U14275 (N_14275,N_9249,N_9200);
or U14276 (N_14276,N_7231,N_5587);
nand U14277 (N_14277,N_7610,N_6445);
and U14278 (N_14278,N_7300,N_7177);
or U14279 (N_14279,N_9391,N_5128);
and U14280 (N_14280,N_8558,N_8448);
and U14281 (N_14281,N_8451,N_9977);
and U14282 (N_14282,N_9389,N_8698);
xor U14283 (N_14283,N_5678,N_8336);
nor U14284 (N_14284,N_8543,N_8077);
nand U14285 (N_14285,N_5390,N_8636);
nor U14286 (N_14286,N_7515,N_9284);
nor U14287 (N_14287,N_9358,N_6166);
nor U14288 (N_14288,N_7095,N_7150);
nor U14289 (N_14289,N_9161,N_7065);
xor U14290 (N_14290,N_5519,N_7276);
nand U14291 (N_14291,N_6325,N_8789);
and U14292 (N_14292,N_8846,N_5858);
and U14293 (N_14293,N_6215,N_8212);
and U14294 (N_14294,N_6350,N_5063);
or U14295 (N_14295,N_6117,N_8243);
and U14296 (N_14296,N_7016,N_6894);
nand U14297 (N_14297,N_5515,N_6422);
or U14298 (N_14298,N_7254,N_8348);
and U14299 (N_14299,N_6620,N_6438);
and U14300 (N_14300,N_7531,N_5755);
nor U14301 (N_14301,N_9983,N_5930);
nand U14302 (N_14302,N_5350,N_6763);
nand U14303 (N_14303,N_8318,N_6454);
or U14304 (N_14304,N_5718,N_8524);
and U14305 (N_14305,N_8520,N_8299);
nand U14306 (N_14306,N_9295,N_7351);
or U14307 (N_14307,N_9922,N_7080);
nand U14308 (N_14308,N_5380,N_8868);
or U14309 (N_14309,N_5864,N_8106);
xnor U14310 (N_14310,N_9803,N_8757);
and U14311 (N_14311,N_5652,N_7494);
and U14312 (N_14312,N_6022,N_5915);
nor U14313 (N_14313,N_5186,N_8653);
nand U14314 (N_14314,N_9731,N_7752);
or U14315 (N_14315,N_9086,N_8888);
nor U14316 (N_14316,N_8359,N_8317);
nand U14317 (N_14317,N_6361,N_7104);
nand U14318 (N_14318,N_6200,N_5812);
nor U14319 (N_14319,N_6689,N_7727);
and U14320 (N_14320,N_7105,N_8194);
nand U14321 (N_14321,N_8840,N_5776);
nand U14322 (N_14322,N_8656,N_9284);
and U14323 (N_14323,N_5080,N_5425);
nand U14324 (N_14324,N_5029,N_9292);
or U14325 (N_14325,N_8297,N_9643);
or U14326 (N_14326,N_9251,N_6494);
nand U14327 (N_14327,N_8279,N_6497);
nand U14328 (N_14328,N_6102,N_8228);
nand U14329 (N_14329,N_8348,N_7607);
or U14330 (N_14330,N_5790,N_7997);
nand U14331 (N_14331,N_6987,N_6087);
nor U14332 (N_14332,N_8135,N_6367);
nor U14333 (N_14333,N_9555,N_6945);
and U14334 (N_14334,N_7548,N_5917);
or U14335 (N_14335,N_9591,N_6987);
and U14336 (N_14336,N_9682,N_8735);
nand U14337 (N_14337,N_9231,N_9269);
xor U14338 (N_14338,N_7748,N_8385);
or U14339 (N_14339,N_8756,N_8744);
or U14340 (N_14340,N_5191,N_5158);
or U14341 (N_14341,N_5381,N_6950);
nand U14342 (N_14342,N_7511,N_6429);
and U14343 (N_14343,N_9027,N_7325);
nor U14344 (N_14344,N_8089,N_7628);
nor U14345 (N_14345,N_6117,N_9040);
nor U14346 (N_14346,N_7852,N_6413);
or U14347 (N_14347,N_9240,N_7263);
or U14348 (N_14348,N_7363,N_8679);
nand U14349 (N_14349,N_5198,N_7417);
nor U14350 (N_14350,N_9859,N_6093);
and U14351 (N_14351,N_9841,N_5965);
or U14352 (N_14352,N_5874,N_8889);
nand U14353 (N_14353,N_7378,N_7298);
and U14354 (N_14354,N_8351,N_8676);
nor U14355 (N_14355,N_6107,N_9737);
or U14356 (N_14356,N_5545,N_9618);
or U14357 (N_14357,N_9965,N_6473);
or U14358 (N_14358,N_6416,N_6324);
nor U14359 (N_14359,N_7124,N_5881);
and U14360 (N_14360,N_6693,N_6197);
or U14361 (N_14361,N_5589,N_6640);
nand U14362 (N_14362,N_5085,N_7919);
or U14363 (N_14363,N_9815,N_6239);
and U14364 (N_14364,N_7492,N_6144);
and U14365 (N_14365,N_8601,N_8365);
nand U14366 (N_14366,N_7074,N_6488);
nand U14367 (N_14367,N_6072,N_8919);
nand U14368 (N_14368,N_6166,N_6100);
or U14369 (N_14369,N_9259,N_7116);
and U14370 (N_14370,N_6331,N_9319);
or U14371 (N_14371,N_9039,N_5136);
nand U14372 (N_14372,N_6361,N_9682);
or U14373 (N_14373,N_6755,N_7275);
or U14374 (N_14374,N_7149,N_8318);
nor U14375 (N_14375,N_5704,N_5257);
and U14376 (N_14376,N_6929,N_8083);
and U14377 (N_14377,N_5153,N_7166);
nor U14378 (N_14378,N_8284,N_8293);
nand U14379 (N_14379,N_9212,N_7622);
nand U14380 (N_14380,N_8866,N_9526);
nand U14381 (N_14381,N_9063,N_8433);
and U14382 (N_14382,N_9098,N_8181);
or U14383 (N_14383,N_9650,N_8000);
or U14384 (N_14384,N_8301,N_5954);
nor U14385 (N_14385,N_9295,N_7756);
nand U14386 (N_14386,N_9981,N_9576);
or U14387 (N_14387,N_8493,N_9573);
nor U14388 (N_14388,N_7456,N_6039);
nor U14389 (N_14389,N_6369,N_6869);
nand U14390 (N_14390,N_9829,N_9436);
or U14391 (N_14391,N_7297,N_9286);
nor U14392 (N_14392,N_8043,N_6335);
nand U14393 (N_14393,N_7150,N_7764);
or U14394 (N_14394,N_7059,N_5008);
nand U14395 (N_14395,N_9165,N_9808);
nor U14396 (N_14396,N_7113,N_9167);
or U14397 (N_14397,N_5737,N_8604);
nor U14398 (N_14398,N_5979,N_5708);
or U14399 (N_14399,N_8483,N_7095);
nor U14400 (N_14400,N_8615,N_9863);
or U14401 (N_14401,N_8170,N_9871);
and U14402 (N_14402,N_6342,N_8629);
or U14403 (N_14403,N_5248,N_7032);
and U14404 (N_14404,N_7765,N_7884);
nand U14405 (N_14405,N_6943,N_8725);
and U14406 (N_14406,N_5561,N_7695);
nor U14407 (N_14407,N_8656,N_5586);
or U14408 (N_14408,N_5079,N_8925);
xor U14409 (N_14409,N_5232,N_8320);
or U14410 (N_14410,N_7388,N_6154);
or U14411 (N_14411,N_8942,N_8759);
nand U14412 (N_14412,N_7813,N_5600);
and U14413 (N_14413,N_7451,N_8522);
or U14414 (N_14414,N_6942,N_8148);
or U14415 (N_14415,N_5648,N_5730);
nor U14416 (N_14416,N_9491,N_6639);
and U14417 (N_14417,N_6173,N_8560);
and U14418 (N_14418,N_6426,N_8719);
and U14419 (N_14419,N_6555,N_5025);
or U14420 (N_14420,N_5960,N_7143);
or U14421 (N_14421,N_8244,N_5063);
nor U14422 (N_14422,N_8466,N_8247);
or U14423 (N_14423,N_9356,N_8069);
nor U14424 (N_14424,N_5071,N_8207);
nor U14425 (N_14425,N_9865,N_5750);
nor U14426 (N_14426,N_7113,N_6197);
or U14427 (N_14427,N_6542,N_7060);
or U14428 (N_14428,N_7746,N_5633);
and U14429 (N_14429,N_9103,N_8856);
and U14430 (N_14430,N_8227,N_7559);
nor U14431 (N_14431,N_7519,N_5129);
and U14432 (N_14432,N_5238,N_7802);
or U14433 (N_14433,N_6310,N_8120);
or U14434 (N_14434,N_5614,N_6996);
nand U14435 (N_14435,N_8631,N_5041);
or U14436 (N_14436,N_9606,N_8310);
nor U14437 (N_14437,N_6776,N_7328);
nor U14438 (N_14438,N_9922,N_5190);
nand U14439 (N_14439,N_7672,N_7801);
and U14440 (N_14440,N_8865,N_7142);
nor U14441 (N_14441,N_7492,N_5889);
and U14442 (N_14442,N_9997,N_8578);
nand U14443 (N_14443,N_7317,N_7961);
and U14444 (N_14444,N_8669,N_6244);
nand U14445 (N_14445,N_7944,N_5289);
and U14446 (N_14446,N_9661,N_8298);
and U14447 (N_14447,N_7911,N_7552);
nand U14448 (N_14448,N_7480,N_5796);
nand U14449 (N_14449,N_8298,N_8804);
or U14450 (N_14450,N_5324,N_5921);
nand U14451 (N_14451,N_5891,N_7041);
nand U14452 (N_14452,N_9135,N_5643);
nand U14453 (N_14453,N_5755,N_7502);
or U14454 (N_14454,N_8688,N_6853);
or U14455 (N_14455,N_9786,N_8109);
or U14456 (N_14456,N_9129,N_7644);
xnor U14457 (N_14457,N_9269,N_8424);
nand U14458 (N_14458,N_8584,N_6848);
and U14459 (N_14459,N_9286,N_6813);
or U14460 (N_14460,N_6927,N_9707);
nor U14461 (N_14461,N_7289,N_7362);
nor U14462 (N_14462,N_6627,N_5710);
and U14463 (N_14463,N_5264,N_6300);
nor U14464 (N_14464,N_9407,N_5038);
or U14465 (N_14465,N_5890,N_5586);
and U14466 (N_14466,N_8434,N_8871);
nand U14467 (N_14467,N_7304,N_6297);
nor U14468 (N_14468,N_6954,N_6024);
or U14469 (N_14469,N_9222,N_5486);
nand U14470 (N_14470,N_6087,N_6887);
and U14471 (N_14471,N_5306,N_6475);
nand U14472 (N_14472,N_5944,N_7389);
nor U14473 (N_14473,N_5446,N_7682);
and U14474 (N_14474,N_8869,N_8002);
nand U14475 (N_14475,N_8530,N_8873);
nand U14476 (N_14476,N_7378,N_9703);
nand U14477 (N_14477,N_9562,N_7713);
nand U14478 (N_14478,N_6413,N_7392);
or U14479 (N_14479,N_6909,N_9646);
nand U14480 (N_14480,N_7783,N_7901);
nor U14481 (N_14481,N_9920,N_6281);
nand U14482 (N_14482,N_7253,N_6444);
nand U14483 (N_14483,N_8230,N_6724);
and U14484 (N_14484,N_9679,N_9713);
xor U14485 (N_14485,N_5613,N_8768);
or U14486 (N_14486,N_9150,N_9491);
or U14487 (N_14487,N_6332,N_8520);
or U14488 (N_14488,N_7209,N_5352);
nand U14489 (N_14489,N_8724,N_5289);
and U14490 (N_14490,N_7957,N_9210);
nand U14491 (N_14491,N_7858,N_5814);
or U14492 (N_14492,N_9200,N_7888);
nand U14493 (N_14493,N_6720,N_9280);
nor U14494 (N_14494,N_9251,N_7665);
nor U14495 (N_14495,N_7731,N_5277);
and U14496 (N_14496,N_5841,N_6564);
or U14497 (N_14497,N_7218,N_9618);
nor U14498 (N_14498,N_6917,N_8917);
xor U14499 (N_14499,N_9963,N_7700);
nor U14500 (N_14500,N_9196,N_6860);
nand U14501 (N_14501,N_6102,N_6595);
and U14502 (N_14502,N_9290,N_5475);
nor U14503 (N_14503,N_7040,N_7888);
nor U14504 (N_14504,N_5881,N_6538);
nand U14505 (N_14505,N_9149,N_7429);
nand U14506 (N_14506,N_7735,N_6436);
or U14507 (N_14507,N_9129,N_9356);
nor U14508 (N_14508,N_6771,N_5881);
and U14509 (N_14509,N_8521,N_6937);
or U14510 (N_14510,N_9802,N_8420);
or U14511 (N_14511,N_9027,N_9325);
nand U14512 (N_14512,N_6002,N_5574);
nor U14513 (N_14513,N_5651,N_5981);
nand U14514 (N_14514,N_6117,N_5036);
nor U14515 (N_14515,N_9305,N_7442);
and U14516 (N_14516,N_6109,N_5611);
nor U14517 (N_14517,N_6253,N_8416);
and U14518 (N_14518,N_9032,N_9822);
nor U14519 (N_14519,N_5578,N_9933);
and U14520 (N_14520,N_6947,N_6317);
or U14521 (N_14521,N_5143,N_8758);
or U14522 (N_14522,N_5429,N_6501);
and U14523 (N_14523,N_6020,N_9756);
or U14524 (N_14524,N_5840,N_8902);
or U14525 (N_14525,N_8348,N_6560);
nand U14526 (N_14526,N_6428,N_6574);
nand U14527 (N_14527,N_8814,N_7842);
and U14528 (N_14528,N_6290,N_9632);
and U14529 (N_14529,N_9223,N_9235);
or U14530 (N_14530,N_7702,N_5710);
and U14531 (N_14531,N_9061,N_7083);
nor U14532 (N_14532,N_8640,N_9364);
nor U14533 (N_14533,N_8911,N_5843);
nor U14534 (N_14534,N_7585,N_7344);
or U14535 (N_14535,N_7961,N_8691);
and U14536 (N_14536,N_9010,N_8775);
and U14537 (N_14537,N_5829,N_6927);
nor U14538 (N_14538,N_7846,N_5710);
and U14539 (N_14539,N_6325,N_5091);
and U14540 (N_14540,N_7759,N_9102);
and U14541 (N_14541,N_9744,N_8764);
nor U14542 (N_14542,N_8094,N_7097);
and U14543 (N_14543,N_7133,N_9434);
xnor U14544 (N_14544,N_7745,N_9357);
nor U14545 (N_14545,N_5169,N_5815);
or U14546 (N_14546,N_6763,N_5873);
nand U14547 (N_14547,N_7422,N_8408);
or U14548 (N_14548,N_6953,N_9178);
nand U14549 (N_14549,N_5963,N_8435);
nand U14550 (N_14550,N_9761,N_7442);
and U14551 (N_14551,N_8558,N_6313);
nor U14552 (N_14552,N_6286,N_8882);
nor U14553 (N_14553,N_8292,N_8192);
or U14554 (N_14554,N_7546,N_9336);
or U14555 (N_14555,N_7284,N_6138);
nor U14556 (N_14556,N_9150,N_9973);
and U14557 (N_14557,N_7143,N_9940);
nor U14558 (N_14558,N_6270,N_8242);
and U14559 (N_14559,N_9504,N_5348);
nor U14560 (N_14560,N_5928,N_8348);
or U14561 (N_14561,N_9642,N_8064);
or U14562 (N_14562,N_8198,N_8362);
nand U14563 (N_14563,N_6406,N_5708);
and U14564 (N_14564,N_7291,N_7421);
nor U14565 (N_14565,N_9615,N_7104);
or U14566 (N_14566,N_5156,N_6966);
and U14567 (N_14567,N_9089,N_8693);
nand U14568 (N_14568,N_7975,N_9344);
or U14569 (N_14569,N_9009,N_7051);
or U14570 (N_14570,N_8078,N_8410);
nor U14571 (N_14571,N_6717,N_7072);
nor U14572 (N_14572,N_5190,N_9015);
nor U14573 (N_14573,N_9842,N_8045);
and U14574 (N_14574,N_5588,N_7000);
and U14575 (N_14575,N_6974,N_7845);
xor U14576 (N_14576,N_7569,N_6307);
and U14577 (N_14577,N_9467,N_8153);
nand U14578 (N_14578,N_6465,N_9089);
nor U14579 (N_14579,N_9152,N_5086);
nor U14580 (N_14580,N_7612,N_7512);
nor U14581 (N_14581,N_7231,N_6535);
and U14582 (N_14582,N_6552,N_9697);
nand U14583 (N_14583,N_5003,N_6162);
or U14584 (N_14584,N_5211,N_5780);
or U14585 (N_14585,N_7693,N_9574);
nand U14586 (N_14586,N_6657,N_6662);
nand U14587 (N_14587,N_9387,N_5897);
or U14588 (N_14588,N_9076,N_7372);
nor U14589 (N_14589,N_9762,N_5561);
xor U14590 (N_14590,N_6559,N_7053);
and U14591 (N_14591,N_6993,N_7611);
nor U14592 (N_14592,N_8145,N_5753);
and U14593 (N_14593,N_6905,N_9409);
nor U14594 (N_14594,N_9035,N_8988);
nand U14595 (N_14595,N_9763,N_7874);
and U14596 (N_14596,N_6987,N_7694);
nor U14597 (N_14597,N_6020,N_8447);
and U14598 (N_14598,N_8040,N_6246);
and U14599 (N_14599,N_9328,N_6762);
nand U14600 (N_14600,N_5240,N_6443);
nand U14601 (N_14601,N_5016,N_8969);
nor U14602 (N_14602,N_7133,N_7054);
nor U14603 (N_14603,N_5410,N_8021);
nand U14604 (N_14604,N_7449,N_5952);
and U14605 (N_14605,N_7420,N_6467);
and U14606 (N_14606,N_7067,N_8844);
xor U14607 (N_14607,N_9665,N_9354);
and U14608 (N_14608,N_7206,N_9320);
nor U14609 (N_14609,N_7779,N_6775);
and U14610 (N_14610,N_5164,N_5523);
nand U14611 (N_14611,N_5627,N_6907);
nand U14612 (N_14612,N_7448,N_5323);
nand U14613 (N_14613,N_7689,N_6991);
or U14614 (N_14614,N_7522,N_5653);
nor U14615 (N_14615,N_9116,N_9059);
or U14616 (N_14616,N_9403,N_5670);
nor U14617 (N_14617,N_5367,N_7049);
nand U14618 (N_14618,N_6185,N_6227);
or U14619 (N_14619,N_7731,N_6611);
nor U14620 (N_14620,N_6509,N_7204);
xor U14621 (N_14621,N_7211,N_9748);
nand U14622 (N_14622,N_9429,N_6035);
and U14623 (N_14623,N_9591,N_7899);
and U14624 (N_14624,N_7229,N_6650);
nand U14625 (N_14625,N_8107,N_7165);
and U14626 (N_14626,N_7133,N_9531);
nand U14627 (N_14627,N_8127,N_8936);
or U14628 (N_14628,N_7420,N_7917);
and U14629 (N_14629,N_9780,N_7413);
nor U14630 (N_14630,N_7476,N_5862);
nor U14631 (N_14631,N_6933,N_6180);
or U14632 (N_14632,N_6398,N_6367);
nand U14633 (N_14633,N_6598,N_5267);
or U14634 (N_14634,N_6328,N_6198);
and U14635 (N_14635,N_7112,N_6863);
and U14636 (N_14636,N_7467,N_6666);
nor U14637 (N_14637,N_7506,N_5217);
or U14638 (N_14638,N_9605,N_7696);
nand U14639 (N_14639,N_7833,N_7982);
nor U14640 (N_14640,N_5531,N_5154);
or U14641 (N_14641,N_6096,N_9062);
nor U14642 (N_14642,N_6416,N_8730);
and U14643 (N_14643,N_7577,N_6994);
and U14644 (N_14644,N_9992,N_5781);
and U14645 (N_14645,N_6999,N_7289);
nand U14646 (N_14646,N_6861,N_8978);
nand U14647 (N_14647,N_6640,N_9296);
and U14648 (N_14648,N_9792,N_9892);
or U14649 (N_14649,N_7763,N_8107);
nor U14650 (N_14650,N_7652,N_6316);
nor U14651 (N_14651,N_7506,N_8578);
nand U14652 (N_14652,N_7601,N_8577);
nand U14653 (N_14653,N_6349,N_5916);
nor U14654 (N_14654,N_9912,N_5115);
or U14655 (N_14655,N_7451,N_7942);
nand U14656 (N_14656,N_7026,N_6056);
or U14657 (N_14657,N_9011,N_8208);
nand U14658 (N_14658,N_6476,N_7095);
nor U14659 (N_14659,N_9017,N_5492);
xor U14660 (N_14660,N_8323,N_5949);
nor U14661 (N_14661,N_8661,N_7420);
nand U14662 (N_14662,N_8929,N_8053);
and U14663 (N_14663,N_5999,N_8917);
nand U14664 (N_14664,N_7173,N_9094);
and U14665 (N_14665,N_8606,N_8908);
nand U14666 (N_14666,N_5138,N_9159);
nor U14667 (N_14667,N_5691,N_7327);
nor U14668 (N_14668,N_8017,N_5752);
nor U14669 (N_14669,N_9248,N_6242);
or U14670 (N_14670,N_9621,N_6265);
and U14671 (N_14671,N_9988,N_8786);
and U14672 (N_14672,N_9179,N_8554);
nor U14673 (N_14673,N_6549,N_9482);
nand U14674 (N_14674,N_8488,N_8908);
nor U14675 (N_14675,N_8055,N_5896);
nand U14676 (N_14676,N_9896,N_8615);
and U14677 (N_14677,N_5788,N_5711);
or U14678 (N_14678,N_9669,N_7286);
nand U14679 (N_14679,N_7935,N_8860);
or U14680 (N_14680,N_7826,N_6023);
nor U14681 (N_14681,N_5348,N_6339);
nor U14682 (N_14682,N_7017,N_6017);
or U14683 (N_14683,N_5756,N_8023);
nand U14684 (N_14684,N_5803,N_9458);
and U14685 (N_14685,N_5949,N_6821);
nor U14686 (N_14686,N_9418,N_8611);
or U14687 (N_14687,N_7113,N_5432);
or U14688 (N_14688,N_9283,N_9019);
nand U14689 (N_14689,N_6976,N_9925);
nor U14690 (N_14690,N_7617,N_6930);
and U14691 (N_14691,N_6383,N_5191);
nand U14692 (N_14692,N_5349,N_8883);
xnor U14693 (N_14693,N_6785,N_7622);
nor U14694 (N_14694,N_8320,N_8272);
nor U14695 (N_14695,N_8317,N_8967);
nand U14696 (N_14696,N_7721,N_8976);
or U14697 (N_14697,N_6659,N_9639);
nor U14698 (N_14698,N_7789,N_7864);
or U14699 (N_14699,N_5724,N_6503);
nand U14700 (N_14700,N_8666,N_8722);
nand U14701 (N_14701,N_8000,N_9367);
or U14702 (N_14702,N_9876,N_8050);
and U14703 (N_14703,N_8722,N_8574);
nor U14704 (N_14704,N_5434,N_6326);
or U14705 (N_14705,N_6729,N_8313);
or U14706 (N_14706,N_6240,N_7513);
nor U14707 (N_14707,N_9708,N_7534);
nor U14708 (N_14708,N_9310,N_8846);
nor U14709 (N_14709,N_7392,N_9273);
and U14710 (N_14710,N_7284,N_9336);
nand U14711 (N_14711,N_9689,N_5163);
nor U14712 (N_14712,N_6230,N_9973);
or U14713 (N_14713,N_6957,N_7082);
nand U14714 (N_14714,N_8267,N_9277);
nor U14715 (N_14715,N_9966,N_8315);
or U14716 (N_14716,N_9768,N_6496);
nor U14717 (N_14717,N_7148,N_7371);
nand U14718 (N_14718,N_5120,N_7417);
nand U14719 (N_14719,N_5157,N_6616);
nor U14720 (N_14720,N_8101,N_6520);
nor U14721 (N_14721,N_9447,N_7667);
nor U14722 (N_14722,N_6625,N_6684);
and U14723 (N_14723,N_6879,N_7351);
nand U14724 (N_14724,N_6407,N_9691);
nor U14725 (N_14725,N_8820,N_7819);
nor U14726 (N_14726,N_8583,N_8807);
nand U14727 (N_14727,N_5263,N_8837);
and U14728 (N_14728,N_8332,N_7940);
and U14729 (N_14729,N_9782,N_5067);
nor U14730 (N_14730,N_5268,N_7185);
or U14731 (N_14731,N_8325,N_5734);
or U14732 (N_14732,N_8027,N_7243);
nand U14733 (N_14733,N_7971,N_6897);
and U14734 (N_14734,N_7804,N_5161);
nand U14735 (N_14735,N_6760,N_7649);
nand U14736 (N_14736,N_8934,N_8807);
nand U14737 (N_14737,N_5357,N_5746);
nor U14738 (N_14738,N_9433,N_9171);
nand U14739 (N_14739,N_8566,N_5467);
nor U14740 (N_14740,N_6958,N_8346);
nand U14741 (N_14741,N_6124,N_9152);
nor U14742 (N_14742,N_5838,N_6655);
nor U14743 (N_14743,N_5239,N_8454);
and U14744 (N_14744,N_7056,N_7538);
nor U14745 (N_14745,N_9513,N_8227);
nor U14746 (N_14746,N_7598,N_9537);
nor U14747 (N_14747,N_7360,N_9171);
and U14748 (N_14748,N_8830,N_6281);
and U14749 (N_14749,N_8062,N_9774);
or U14750 (N_14750,N_8895,N_6037);
or U14751 (N_14751,N_6610,N_5935);
and U14752 (N_14752,N_5623,N_5587);
and U14753 (N_14753,N_7628,N_6211);
and U14754 (N_14754,N_9757,N_9787);
and U14755 (N_14755,N_9499,N_6818);
nor U14756 (N_14756,N_9331,N_9764);
nor U14757 (N_14757,N_5298,N_9726);
nand U14758 (N_14758,N_8671,N_7259);
or U14759 (N_14759,N_9391,N_6844);
or U14760 (N_14760,N_8893,N_9520);
or U14761 (N_14761,N_6849,N_8457);
and U14762 (N_14762,N_8617,N_5322);
or U14763 (N_14763,N_7497,N_5443);
nor U14764 (N_14764,N_8679,N_7155);
and U14765 (N_14765,N_7492,N_7467);
or U14766 (N_14766,N_5035,N_6554);
or U14767 (N_14767,N_7066,N_7584);
and U14768 (N_14768,N_5826,N_6036);
or U14769 (N_14769,N_6286,N_6498);
nor U14770 (N_14770,N_5363,N_8087);
nor U14771 (N_14771,N_5571,N_6731);
and U14772 (N_14772,N_9357,N_8596);
nand U14773 (N_14773,N_7180,N_7703);
and U14774 (N_14774,N_6139,N_9519);
nor U14775 (N_14775,N_9050,N_8323);
nand U14776 (N_14776,N_6227,N_8952);
and U14777 (N_14777,N_8948,N_5777);
and U14778 (N_14778,N_7817,N_6200);
and U14779 (N_14779,N_6568,N_9516);
nor U14780 (N_14780,N_7130,N_9085);
nor U14781 (N_14781,N_8819,N_8078);
nand U14782 (N_14782,N_6179,N_9498);
and U14783 (N_14783,N_5410,N_7292);
nand U14784 (N_14784,N_6041,N_9644);
or U14785 (N_14785,N_7608,N_8512);
or U14786 (N_14786,N_5321,N_9867);
and U14787 (N_14787,N_9951,N_9388);
nor U14788 (N_14788,N_6617,N_9910);
nand U14789 (N_14789,N_8507,N_9810);
nand U14790 (N_14790,N_5478,N_8121);
or U14791 (N_14791,N_5815,N_6837);
nand U14792 (N_14792,N_9302,N_6034);
nand U14793 (N_14793,N_8442,N_6961);
or U14794 (N_14794,N_8414,N_8659);
nand U14795 (N_14795,N_8349,N_7695);
or U14796 (N_14796,N_8784,N_8631);
or U14797 (N_14797,N_6335,N_7301);
nand U14798 (N_14798,N_5053,N_5249);
nand U14799 (N_14799,N_9425,N_7571);
nand U14800 (N_14800,N_7936,N_6455);
or U14801 (N_14801,N_5240,N_7019);
or U14802 (N_14802,N_7623,N_8011);
nor U14803 (N_14803,N_8539,N_9183);
and U14804 (N_14804,N_8101,N_5072);
nand U14805 (N_14805,N_5830,N_9943);
nor U14806 (N_14806,N_5131,N_8876);
nor U14807 (N_14807,N_5357,N_6498);
or U14808 (N_14808,N_6029,N_7788);
nor U14809 (N_14809,N_5800,N_9694);
and U14810 (N_14810,N_7668,N_5433);
or U14811 (N_14811,N_8812,N_9502);
and U14812 (N_14812,N_9665,N_5511);
or U14813 (N_14813,N_9680,N_5560);
or U14814 (N_14814,N_5195,N_7752);
nand U14815 (N_14815,N_6510,N_5856);
or U14816 (N_14816,N_5297,N_6854);
nor U14817 (N_14817,N_8261,N_5361);
nor U14818 (N_14818,N_5330,N_8963);
or U14819 (N_14819,N_6798,N_9162);
nor U14820 (N_14820,N_7139,N_5524);
nor U14821 (N_14821,N_6407,N_9725);
or U14822 (N_14822,N_8496,N_7838);
nor U14823 (N_14823,N_7894,N_5904);
or U14824 (N_14824,N_7821,N_5740);
or U14825 (N_14825,N_6245,N_8133);
and U14826 (N_14826,N_6192,N_6400);
and U14827 (N_14827,N_6695,N_5663);
or U14828 (N_14828,N_6236,N_5374);
nor U14829 (N_14829,N_6699,N_7472);
and U14830 (N_14830,N_5814,N_5317);
nand U14831 (N_14831,N_6786,N_6240);
nor U14832 (N_14832,N_6248,N_9231);
or U14833 (N_14833,N_6764,N_8253);
and U14834 (N_14834,N_9507,N_7820);
nand U14835 (N_14835,N_5348,N_9082);
nor U14836 (N_14836,N_9598,N_9857);
or U14837 (N_14837,N_7675,N_5700);
and U14838 (N_14838,N_6894,N_7892);
or U14839 (N_14839,N_5462,N_8369);
nor U14840 (N_14840,N_7037,N_7568);
or U14841 (N_14841,N_6721,N_5693);
and U14842 (N_14842,N_9911,N_7683);
nor U14843 (N_14843,N_9708,N_8033);
nor U14844 (N_14844,N_6736,N_6126);
nand U14845 (N_14845,N_9947,N_9622);
nand U14846 (N_14846,N_8619,N_7397);
nand U14847 (N_14847,N_7015,N_6415);
nor U14848 (N_14848,N_7220,N_6413);
nand U14849 (N_14849,N_9353,N_9461);
nand U14850 (N_14850,N_5936,N_9805);
nand U14851 (N_14851,N_7599,N_9602);
or U14852 (N_14852,N_9048,N_9197);
and U14853 (N_14853,N_6201,N_7812);
or U14854 (N_14854,N_8116,N_8442);
or U14855 (N_14855,N_7315,N_6756);
and U14856 (N_14856,N_7064,N_8009);
nor U14857 (N_14857,N_7367,N_6423);
or U14858 (N_14858,N_6098,N_8904);
and U14859 (N_14859,N_9708,N_7750);
or U14860 (N_14860,N_8850,N_5906);
or U14861 (N_14861,N_8383,N_7344);
nor U14862 (N_14862,N_7820,N_5167);
and U14863 (N_14863,N_7292,N_6659);
and U14864 (N_14864,N_7745,N_9087);
or U14865 (N_14865,N_5199,N_5249);
nor U14866 (N_14866,N_8804,N_9335);
nor U14867 (N_14867,N_9364,N_9122);
nor U14868 (N_14868,N_9691,N_6278);
and U14869 (N_14869,N_7929,N_9890);
or U14870 (N_14870,N_5940,N_6983);
nand U14871 (N_14871,N_8788,N_6074);
xnor U14872 (N_14872,N_9460,N_8493);
nor U14873 (N_14873,N_9041,N_7944);
and U14874 (N_14874,N_7281,N_6476);
or U14875 (N_14875,N_7185,N_9826);
and U14876 (N_14876,N_9517,N_8029);
or U14877 (N_14877,N_8867,N_9854);
nand U14878 (N_14878,N_9257,N_9406);
or U14879 (N_14879,N_6385,N_5443);
nor U14880 (N_14880,N_6003,N_5594);
nor U14881 (N_14881,N_6959,N_8274);
and U14882 (N_14882,N_8140,N_8292);
and U14883 (N_14883,N_6819,N_8674);
or U14884 (N_14884,N_7438,N_7673);
or U14885 (N_14885,N_8306,N_7977);
nor U14886 (N_14886,N_9753,N_6657);
nand U14887 (N_14887,N_8008,N_8420);
nor U14888 (N_14888,N_7908,N_6156);
nor U14889 (N_14889,N_7027,N_7065);
nor U14890 (N_14890,N_7340,N_5865);
nand U14891 (N_14891,N_5755,N_9552);
or U14892 (N_14892,N_7767,N_8162);
nor U14893 (N_14893,N_9557,N_8959);
nand U14894 (N_14894,N_7580,N_5005);
nand U14895 (N_14895,N_7884,N_6083);
nor U14896 (N_14896,N_7259,N_8257);
nor U14897 (N_14897,N_6431,N_7557);
nor U14898 (N_14898,N_7865,N_9885);
nor U14899 (N_14899,N_7795,N_5377);
nor U14900 (N_14900,N_9457,N_9355);
and U14901 (N_14901,N_7142,N_9550);
nor U14902 (N_14902,N_5942,N_9965);
nand U14903 (N_14903,N_9628,N_6771);
nor U14904 (N_14904,N_8635,N_8457);
or U14905 (N_14905,N_7393,N_5601);
nand U14906 (N_14906,N_8156,N_8010);
nor U14907 (N_14907,N_9000,N_6356);
nand U14908 (N_14908,N_9220,N_8313);
nand U14909 (N_14909,N_6784,N_9665);
nor U14910 (N_14910,N_9974,N_8287);
or U14911 (N_14911,N_9782,N_5229);
or U14912 (N_14912,N_5274,N_6846);
and U14913 (N_14913,N_7834,N_8021);
or U14914 (N_14914,N_7782,N_7280);
or U14915 (N_14915,N_9250,N_7297);
or U14916 (N_14916,N_6720,N_7089);
nor U14917 (N_14917,N_5929,N_8167);
and U14918 (N_14918,N_5227,N_6602);
nor U14919 (N_14919,N_8632,N_6684);
nand U14920 (N_14920,N_7114,N_8464);
and U14921 (N_14921,N_5105,N_6828);
or U14922 (N_14922,N_5648,N_6706);
nand U14923 (N_14923,N_5383,N_5043);
or U14924 (N_14924,N_7184,N_7785);
nand U14925 (N_14925,N_5593,N_8382);
or U14926 (N_14926,N_9815,N_9505);
nor U14927 (N_14927,N_9787,N_8219);
nand U14928 (N_14928,N_5047,N_8971);
or U14929 (N_14929,N_6274,N_6300);
nor U14930 (N_14930,N_5939,N_5458);
nor U14931 (N_14931,N_8990,N_9332);
nand U14932 (N_14932,N_6993,N_5859);
or U14933 (N_14933,N_7970,N_5219);
nor U14934 (N_14934,N_8773,N_7354);
nand U14935 (N_14935,N_6102,N_7102);
or U14936 (N_14936,N_6814,N_8948);
nor U14937 (N_14937,N_6386,N_9522);
nor U14938 (N_14938,N_5346,N_9998);
or U14939 (N_14939,N_7715,N_7401);
or U14940 (N_14940,N_9551,N_8806);
and U14941 (N_14941,N_8155,N_8545);
nor U14942 (N_14942,N_8663,N_6145);
or U14943 (N_14943,N_8091,N_8434);
nand U14944 (N_14944,N_7077,N_9630);
or U14945 (N_14945,N_8355,N_7075);
nor U14946 (N_14946,N_8579,N_9140);
nor U14947 (N_14947,N_8795,N_6686);
or U14948 (N_14948,N_7801,N_5946);
nand U14949 (N_14949,N_5417,N_5348);
nand U14950 (N_14950,N_6672,N_9601);
or U14951 (N_14951,N_7517,N_5176);
nor U14952 (N_14952,N_8530,N_9097);
or U14953 (N_14953,N_9585,N_9400);
or U14954 (N_14954,N_7215,N_6908);
or U14955 (N_14955,N_8249,N_6443);
or U14956 (N_14956,N_7878,N_5900);
or U14957 (N_14957,N_8194,N_5741);
nand U14958 (N_14958,N_8812,N_7186);
nand U14959 (N_14959,N_9371,N_5249);
and U14960 (N_14960,N_7649,N_6271);
nor U14961 (N_14961,N_6289,N_8943);
or U14962 (N_14962,N_8031,N_7732);
and U14963 (N_14963,N_7008,N_8831);
nand U14964 (N_14964,N_7955,N_8780);
nor U14965 (N_14965,N_7244,N_7423);
and U14966 (N_14966,N_6931,N_8553);
or U14967 (N_14967,N_7591,N_5572);
nand U14968 (N_14968,N_5716,N_7012);
nor U14969 (N_14969,N_8230,N_8996);
nand U14970 (N_14970,N_6458,N_5834);
nand U14971 (N_14971,N_9203,N_8325);
nand U14972 (N_14972,N_7023,N_9459);
and U14973 (N_14973,N_8786,N_6909);
and U14974 (N_14974,N_6908,N_7097);
nor U14975 (N_14975,N_5473,N_7338);
xnor U14976 (N_14976,N_6253,N_6670);
and U14977 (N_14977,N_7081,N_9299);
nand U14978 (N_14978,N_9011,N_5633);
and U14979 (N_14979,N_9756,N_8825);
or U14980 (N_14980,N_9520,N_9175);
or U14981 (N_14981,N_5833,N_8929);
or U14982 (N_14982,N_6298,N_6433);
nand U14983 (N_14983,N_6724,N_6352);
nor U14984 (N_14984,N_5198,N_7730);
or U14985 (N_14985,N_8826,N_7842);
nor U14986 (N_14986,N_9126,N_9281);
and U14987 (N_14987,N_5804,N_9402);
or U14988 (N_14988,N_7931,N_5805);
nand U14989 (N_14989,N_9104,N_5192);
nand U14990 (N_14990,N_5894,N_7894);
or U14991 (N_14991,N_7343,N_7011);
nand U14992 (N_14992,N_8625,N_5347);
and U14993 (N_14993,N_8505,N_7173);
nor U14994 (N_14994,N_5810,N_8753);
or U14995 (N_14995,N_7019,N_8984);
or U14996 (N_14996,N_9550,N_6267);
and U14997 (N_14997,N_9289,N_7114);
nand U14998 (N_14998,N_8615,N_6710);
nand U14999 (N_14999,N_6966,N_6794);
nor U15000 (N_15000,N_10808,N_14379);
nand U15001 (N_15001,N_12635,N_11442);
nor U15002 (N_15002,N_11476,N_13508);
nand U15003 (N_15003,N_11112,N_13371);
nor U15004 (N_15004,N_11861,N_12935);
and U15005 (N_15005,N_13080,N_11863);
and U15006 (N_15006,N_10990,N_10747);
and U15007 (N_15007,N_14053,N_14477);
nor U15008 (N_15008,N_14141,N_12077);
nor U15009 (N_15009,N_11032,N_10198);
nand U15010 (N_15010,N_10149,N_11837);
or U15011 (N_15011,N_12158,N_12697);
nand U15012 (N_15012,N_12460,N_14295);
or U15013 (N_15013,N_13214,N_12989);
and U15014 (N_15014,N_14862,N_12601);
and U15015 (N_15015,N_13399,N_10493);
nor U15016 (N_15016,N_12062,N_12627);
and U15017 (N_15017,N_11995,N_13370);
xnor U15018 (N_15018,N_10051,N_12821);
nor U15019 (N_15019,N_11139,N_12897);
nor U15020 (N_15020,N_12625,N_13088);
or U15021 (N_15021,N_14592,N_14464);
nand U15022 (N_15022,N_10937,N_13547);
nor U15023 (N_15023,N_14750,N_14072);
and U15024 (N_15024,N_11297,N_10619);
nand U15025 (N_15025,N_11952,N_13453);
and U15026 (N_15026,N_14349,N_14480);
and U15027 (N_15027,N_11488,N_13792);
nand U15028 (N_15028,N_11343,N_11178);
and U15029 (N_15029,N_10509,N_13386);
or U15030 (N_15030,N_13879,N_13805);
xor U15031 (N_15031,N_13362,N_10642);
nor U15032 (N_15032,N_13662,N_10878);
nand U15033 (N_15033,N_14010,N_12513);
and U15034 (N_15034,N_11936,N_11512);
or U15035 (N_15035,N_13537,N_11968);
nor U15036 (N_15036,N_10162,N_14932);
and U15037 (N_15037,N_11843,N_14763);
and U15038 (N_15038,N_12688,N_13069);
or U15039 (N_15039,N_12547,N_14009);
or U15040 (N_15040,N_11081,N_13378);
nor U15041 (N_15041,N_12856,N_12857);
or U15042 (N_15042,N_14908,N_12340);
or U15043 (N_15043,N_14043,N_12745);
and U15044 (N_15044,N_13440,N_11966);
and U15045 (N_15045,N_14935,N_12047);
and U15046 (N_15046,N_14805,N_14201);
or U15047 (N_15047,N_10068,N_13498);
nand U15048 (N_15048,N_12562,N_10394);
or U15049 (N_15049,N_11043,N_12503);
or U15050 (N_15050,N_10185,N_11485);
or U15051 (N_15051,N_13005,N_13142);
and U15052 (N_15052,N_11576,N_13583);
nand U15053 (N_15053,N_10161,N_13392);
nor U15054 (N_15054,N_11593,N_11201);
and U15055 (N_15055,N_11963,N_14425);
nor U15056 (N_15056,N_10345,N_13111);
nand U15057 (N_15057,N_13947,N_10825);
nor U15058 (N_15058,N_11132,N_14760);
or U15059 (N_15059,N_13319,N_11867);
nor U15060 (N_15060,N_12822,N_12032);
and U15061 (N_15061,N_14291,N_14687);
nand U15062 (N_15062,N_11763,N_11188);
and U15063 (N_15063,N_10041,N_10268);
nand U15064 (N_15064,N_12643,N_10508);
nor U15065 (N_15065,N_13798,N_13235);
and U15066 (N_15066,N_11959,N_11249);
or U15067 (N_15067,N_12235,N_14775);
or U15068 (N_15068,N_11571,N_13604);
nand U15069 (N_15069,N_10171,N_10823);
and U15070 (N_15070,N_14797,N_13169);
or U15071 (N_15071,N_14699,N_12452);
and U15072 (N_15072,N_14368,N_12837);
nand U15073 (N_15073,N_11379,N_14086);
nand U15074 (N_15074,N_10444,N_14710);
nor U15075 (N_15075,N_10404,N_11236);
or U15076 (N_15076,N_11886,N_11631);
nor U15077 (N_15077,N_11222,N_14910);
and U15078 (N_15078,N_14114,N_10675);
and U15079 (N_15079,N_12286,N_14757);
or U15080 (N_15080,N_14815,N_12828);
or U15081 (N_15081,N_13841,N_11753);
nand U15082 (N_15082,N_13667,N_12679);
and U15083 (N_15083,N_12248,N_13634);
and U15084 (N_15084,N_14284,N_13196);
or U15085 (N_15085,N_14494,N_13172);
nand U15086 (N_15086,N_10361,N_13028);
nand U15087 (N_15087,N_13382,N_13497);
nand U15088 (N_15088,N_11326,N_14411);
and U15089 (N_15089,N_12663,N_14023);
and U15090 (N_15090,N_11701,N_12882);
nand U15091 (N_15091,N_10193,N_14279);
or U15092 (N_15092,N_14694,N_11432);
nand U15093 (N_15093,N_11725,N_12031);
and U15094 (N_15094,N_12401,N_10869);
and U15095 (N_15095,N_10028,N_13874);
or U15096 (N_15096,N_14709,N_13670);
and U15097 (N_15097,N_12303,N_11662);
nand U15098 (N_15098,N_11786,N_10058);
nor U15099 (N_15099,N_11879,N_11862);
nand U15100 (N_15100,N_10875,N_13188);
nand U15101 (N_15101,N_14383,N_13231);
and U15102 (N_15102,N_14904,N_11412);
or U15103 (N_15103,N_12693,N_11819);
and U15104 (N_15104,N_10608,N_11364);
nor U15105 (N_15105,N_11623,N_14752);
nand U15106 (N_15106,N_14591,N_12993);
nand U15107 (N_15107,N_12858,N_12937);
nor U15108 (N_15108,N_10606,N_12215);
or U15109 (N_15109,N_11667,N_12398);
and U15110 (N_15110,N_13760,N_11308);
nand U15111 (N_15111,N_14593,N_10164);
or U15112 (N_15112,N_14623,N_10874);
nor U15113 (N_15113,N_14215,N_13285);
nor U15114 (N_15114,N_14437,N_10527);
and U15115 (N_15115,N_10353,N_14265);
and U15116 (N_15116,N_12768,N_11594);
xor U15117 (N_15117,N_12468,N_10661);
nand U15118 (N_15118,N_13513,N_13819);
and U15119 (N_15119,N_14831,N_11301);
or U15120 (N_15120,N_13344,N_10632);
nor U15121 (N_15121,N_12556,N_11979);
and U15122 (N_15122,N_13922,N_10671);
nor U15123 (N_15123,N_11305,N_13121);
and U15124 (N_15124,N_14223,N_12023);
nand U15125 (N_15125,N_14803,N_11806);
nand U15126 (N_15126,N_12408,N_13936);
nand U15127 (N_15127,N_11760,N_13778);
nand U15128 (N_15128,N_14817,N_12714);
and U15129 (N_15129,N_13683,N_12021);
nor U15130 (N_15130,N_12859,N_12879);
or U15131 (N_15131,N_13430,N_11585);
nand U15132 (N_15132,N_12400,N_10759);
and U15133 (N_15133,N_13212,N_11816);
nand U15134 (N_15134,N_12881,N_13522);
nor U15135 (N_15135,N_13108,N_14917);
or U15136 (N_15136,N_13131,N_12593);
nor U15137 (N_15137,N_10548,N_14030);
or U15138 (N_15138,N_12252,N_11820);
or U15139 (N_15139,N_11542,N_12181);
nor U15140 (N_15140,N_10749,N_13691);
and U15141 (N_15141,N_14941,N_13518);
nand U15142 (N_15142,N_11764,N_12082);
nor U15143 (N_15143,N_14345,N_10475);
nand U15144 (N_15144,N_14766,N_11254);
and U15145 (N_15145,N_12998,N_11513);
or U15146 (N_15146,N_14886,N_11358);
nand U15147 (N_15147,N_12591,N_11164);
nand U15148 (N_15148,N_10641,N_13967);
nor U15149 (N_15149,N_11983,N_13999);
nand U15150 (N_15150,N_14585,N_14548);
nand U15151 (N_15151,N_14317,N_10796);
nand U15152 (N_15152,N_11591,N_11160);
nor U15153 (N_15153,N_10303,N_12916);
nor U15154 (N_15154,N_14997,N_11857);
or U15155 (N_15155,N_10929,N_14181);
nor U15156 (N_15156,N_14981,N_11565);
nor U15157 (N_15157,N_10334,N_11864);
and U15158 (N_15158,N_10428,N_13880);
nor U15159 (N_15159,N_14896,N_10775);
or U15160 (N_15160,N_10063,N_11238);
nand U15161 (N_15161,N_11729,N_14088);
nor U15162 (N_15162,N_11940,N_12033);
nand U15163 (N_15163,N_10147,N_14404);
nand U15164 (N_15164,N_13727,N_14857);
nor U15165 (N_15165,N_10468,N_12182);
and U15166 (N_15166,N_12175,N_12670);
xnor U15167 (N_15167,N_14033,N_14951);
or U15168 (N_15168,N_13367,N_11618);
nand U15169 (N_15169,N_10811,N_11179);
or U15170 (N_15170,N_14270,N_14370);
nand U15171 (N_15171,N_14157,N_11289);
nand U15172 (N_15172,N_11429,N_13376);
nand U15173 (N_15173,N_13867,N_11762);
nand U15174 (N_15174,N_10052,N_10265);
nor U15175 (N_15175,N_12131,N_13763);
or U15176 (N_15176,N_12708,N_14773);
and U15177 (N_15177,N_13588,N_13032);
nor U15178 (N_15178,N_14628,N_12926);
and U15179 (N_15179,N_10994,N_11775);
nand U15180 (N_15180,N_12150,N_14583);
nand U15181 (N_15181,N_14060,N_14034);
nand U15182 (N_15182,N_10190,N_11997);
nand U15183 (N_15183,N_13755,N_11135);
nand U15184 (N_15184,N_10368,N_14983);
nor U15185 (N_15185,N_13355,N_10628);
or U15186 (N_15186,N_13656,N_10914);
nand U15187 (N_15187,N_13448,N_11166);
nor U15188 (N_15188,N_10492,N_10941);
xor U15189 (N_15189,N_14662,N_10554);
nand U15190 (N_15190,N_13152,N_10383);
nor U15191 (N_15191,N_11814,N_13322);
nand U15192 (N_15192,N_10377,N_11812);
nand U15193 (N_15193,N_14745,N_13192);
and U15194 (N_15194,N_13380,N_13254);
and U15195 (N_15195,N_12491,N_13642);
nand U15196 (N_15196,N_12242,N_12793);
nor U15197 (N_15197,N_13988,N_12519);
or U15198 (N_15198,N_14216,N_12843);
nor U15199 (N_15199,N_10340,N_13165);
or U15200 (N_15200,N_10278,N_11070);
nor U15201 (N_15201,N_13669,N_13881);
or U15202 (N_15202,N_13109,N_11477);
and U15203 (N_15203,N_12093,N_12337);
and U15204 (N_15204,N_12344,N_10782);
and U15205 (N_15205,N_13351,N_11713);
nor U15206 (N_15206,N_14439,N_10395);
and U15207 (N_15207,N_10230,N_13470);
or U15208 (N_15208,N_13789,N_14285);
nand U15209 (N_15209,N_14684,N_11443);
or U15210 (N_15210,N_13707,N_10788);
and U15211 (N_15211,N_11770,N_14144);
or U15212 (N_15212,N_10460,N_11727);
nor U15213 (N_15213,N_13124,N_10216);
and U15214 (N_15214,N_10537,N_12001);
nor U15215 (N_15215,N_10237,N_14465);
nand U15216 (N_15216,N_10301,N_14565);
nand U15217 (N_15217,N_10648,N_13290);
and U15218 (N_15218,N_13052,N_10656);
and U15219 (N_15219,N_10282,N_14203);
or U15220 (N_15220,N_12335,N_11791);
nor U15221 (N_15221,N_12944,N_12059);
xnor U15222 (N_15222,N_13671,N_11445);
nor U15223 (N_15223,N_14726,N_10089);
nand U15224 (N_15224,N_11214,N_13284);
or U15225 (N_15225,N_14994,N_14047);
or U15226 (N_15226,N_12063,N_14354);
nand U15227 (N_15227,N_13815,N_11163);
or U15228 (N_15228,N_11597,N_10911);
and U15229 (N_15229,N_13694,N_10705);
and U15230 (N_15230,N_13216,N_13586);
and U15231 (N_15231,N_13049,N_10917);
or U15232 (N_15232,N_11507,N_13233);
nand U15233 (N_15233,N_11716,N_14723);
and U15234 (N_15234,N_13985,N_10506);
nand U15235 (N_15235,N_11502,N_12675);
or U15236 (N_15236,N_14446,N_10567);
nand U15237 (N_15237,N_11552,N_10127);
nor U15238 (N_15238,N_12192,N_14800);
and U15239 (N_15239,N_11553,N_11490);
and U15240 (N_15240,N_14827,N_12109);
or U15241 (N_15241,N_12255,N_10598);
nand U15242 (N_15242,N_11102,N_10202);
and U15243 (N_15243,N_10317,N_10812);
or U15244 (N_15244,N_11311,N_12350);
or U15245 (N_15245,N_14676,N_10450);
nand U15246 (N_15246,N_11548,N_14542);
or U15247 (N_15247,N_12734,N_14074);
nor U15248 (N_15248,N_12863,N_13971);
and U15249 (N_15249,N_10634,N_14454);
nor U15250 (N_15250,N_12883,N_13341);
or U15251 (N_15251,N_11744,N_11818);
or U15252 (N_15252,N_12939,N_10709);
and U15253 (N_15253,N_12095,N_14649);
or U15254 (N_15254,N_10943,N_13684);
or U15255 (N_15255,N_10349,N_12798);
and U15256 (N_15256,N_10693,N_13031);
and U15257 (N_15257,N_10668,N_11742);
or U15258 (N_15258,N_11221,N_10735);
and U15259 (N_15259,N_10767,N_14619);
nand U15260 (N_15260,N_11710,N_10768);
nor U15261 (N_15261,N_10088,N_12477);
nor U15262 (N_15262,N_11482,N_13208);
or U15263 (N_15263,N_11537,N_13037);
or U15264 (N_15264,N_10729,N_14422);
nor U15265 (N_15265,N_14125,N_13607);
and U15266 (N_15266,N_12359,N_13054);
nor U15267 (N_15267,N_10546,N_12207);
and U15268 (N_15268,N_10667,N_14235);
nor U15269 (N_15269,N_12665,N_11381);
nor U15270 (N_15270,N_11899,N_13421);
and U15271 (N_15271,N_12457,N_12145);
nor U15272 (N_15272,N_14283,N_14966);
and U15273 (N_15273,N_13060,N_13368);
or U15274 (N_15274,N_10575,N_12766);
nand U15275 (N_15275,N_11817,N_13123);
or U15276 (N_15276,N_14517,N_12880);
nor U15277 (N_15277,N_13477,N_14021);
nand U15278 (N_15278,N_11954,N_13925);
and U15279 (N_15279,N_13217,N_12361);
nand U15280 (N_15280,N_12819,N_12396);
nor U15281 (N_15281,N_14701,N_10133);
nand U15282 (N_15282,N_13945,N_13542);
nand U15283 (N_15283,N_12183,N_13160);
nand U15284 (N_15284,N_12247,N_12508);
nand U15285 (N_15285,N_12736,N_10163);
nand U15286 (N_15286,N_12617,N_11419);
nor U15287 (N_15287,N_12966,N_12572);
and U15288 (N_15288,N_13850,N_14423);
or U15289 (N_15289,N_14200,N_14461);
nand U15290 (N_15290,N_10044,N_10580);
nand U15291 (N_15291,N_11699,N_14609);
nor U15292 (N_15292,N_10047,N_13941);
nor U15293 (N_15293,N_13664,N_10523);
nand U15294 (N_15294,N_11156,N_14737);
and U15295 (N_15295,N_13270,N_14244);
nand U15296 (N_15296,N_14725,N_12802);
nand U15297 (N_15297,N_10605,N_12517);
nor U15298 (N_15298,N_12539,N_14778);
nand U15299 (N_15299,N_10949,N_12105);
nor U15300 (N_15300,N_11091,N_12085);
nor U15301 (N_15301,N_10474,N_10741);
and U15302 (N_15302,N_10263,N_11389);
nand U15303 (N_15303,N_12762,N_13602);
and U15304 (N_15304,N_12185,N_10889);
or U15305 (N_15305,N_13744,N_10321);
and U15306 (N_15306,N_10388,N_11397);
and U15307 (N_15307,N_11598,N_14596);
nor U15308 (N_15308,N_10098,N_13712);
and U15309 (N_15309,N_10888,N_11986);
and U15310 (N_15310,N_12487,N_14842);
nor U15311 (N_15311,N_14079,N_12614);
and U15312 (N_15312,N_11134,N_11914);
nor U15313 (N_15313,N_13565,N_14399);
or U15314 (N_15314,N_14453,N_10480);
nand U15315 (N_15315,N_13832,N_13245);
and U15316 (N_15316,N_12659,N_11588);
nand U15317 (N_15317,N_10000,N_13242);
nor U15318 (N_15318,N_14607,N_12342);
or U15319 (N_15319,N_14897,N_14485);
and U15320 (N_15320,N_10827,N_13483);
or U15321 (N_15321,N_13799,N_12003);
and U15322 (N_15322,N_13632,N_14004);
nand U15323 (N_15323,N_13749,N_13445);
nor U15324 (N_15324,N_14921,N_12414);
nor U15325 (N_15325,N_13061,N_11802);
nand U15326 (N_15326,N_14080,N_14447);
nand U15327 (N_15327,N_10046,N_11341);
and U15328 (N_15328,N_12710,N_13992);
nand U15329 (N_15329,N_10924,N_14669);
or U15330 (N_15330,N_14905,N_10625);
nor U15331 (N_15331,N_11549,N_10573);
nand U15332 (N_15332,N_14294,N_12731);
nand U15333 (N_15333,N_13576,N_14866);
nand U15334 (N_15334,N_13260,N_14729);
nand U15335 (N_15335,N_10602,N_14320);
nor U15336 (N_15336,N_14656,N_10545);
nor U15337 (N_15337,N_14540,N_12190);
and U15338 (N_15338,N_11972,N_14885);
nand U15339 (N_15339,N_14918,N_12450);
or U15340 (N_15340,N_14845,N_11480);
or U15341 (N_15341,N_10013,N_13577);
or U15342 (N_15342,N_10210,N_14873);
nor U15343 (N_15343,N_14631,N_12648);
and U15344 (N_15344,N_10950,N_12971);
and U15345 (N_15345,N_11789,N_11388);
nor U15346 (N_15346,N_12630,N_13699);
nor U15347 (N_15347,N_13311,N_14007);
nand U15348 (N_15348,N_13892,N_10389);
nor U15349 (N_15349,N_14324,N_14025);
or U15350 (N_15350,N_14850,N_12680);
nor U15351 (N_15351,N_11281,N_13743);
nand U15352 (N_15352,N_14512,N_13595);
or U15353 (N_15353,N_11253,N_13578);
nand U15354 (N_15354,N_13682,N_10452);
nor U15355 (N_15355,N_14581,N_12026);
nor U15356 (N_15356,N_11491,N_14603);
nor U15357 (N_15357,N_13891,N_13651);
and U15358 (N_15358,N_12632,N_11300);
and U15359 (N_15359,N_14924,N_14503);
nor U15360 (N_15360,N_10845,N_13237);
and U15361 (N_15361,N_13296,N_12706);
nor U15362 (N_15362,N_13346,N_14974);
and U15363 (N_15363,N_11154,N_13639);
or U15364 (N_15364,N_12232,N_13894);
nand U15365 (N_15365,N_11447,N_14559);
or U15366 (N_15366,N_13885,N_11366);
and U15367 (N_15367,N_10030,N_10274);
nand U15368 (N_15368,N_10243,N_14174);
or U15369 (N_15369,N_13998,N_12641);
or U15370 (N_15370,N_14832,N_14037);
nand U15371 (N_15371,N_13558,N_13105);
or U15372 (N_15372,N_14663,N_10835);
or U15373 (N_15373,N_13385,N_10390);
xor U15374 (N_15374,N_14696,N_13006);
nand U15375 (N_15375,N_14632,N_12057);
nor U15376 (N_15376,N_10027,N_14521);
and U15377 (N_15377,N_13675,N_13514);
nand U15378 (N_15378,N_11099,N_13143);
and U15379 (N_15379,N_12536,N_14516);
nor U15380 (N_15380,N_10771,N_14736);
and U15381 (N_15381,N_14658,N_10558);
nor U15382 (N_15382,N_13776,N_13816);
nand U15383 (N_15383,N_14054,N_11185);
nand U15384 (N_15384,N_10560,N_11088);
or U15385 (N_15385,N_11721,N_12369);
and U15386 (N_15386,N_14550,N_13249);
nand U15387 (N_15387,N_11518,N_11093);
or U15388 (N_15388,N_11145,N_13467);
nand U15389 (N_15389,N_12540,N_13638);
nand U15390 (N_15390,N_12898,N_11520);
and U15391 (N_15391,N_14195,N_11212);
nand U15392 (N_15392,N_13862,N_12574);
and U15393 (N_15393,N_10977,N_14206);
nand U15394 (N_15394,N_13929,N_13701);
and U15395 (N_15395,N_13531,N_13794);
nand U15396 (N_15396,N_10148,N_12498);
nand U15397 (N_15397,N_14865,N_13865);
and U15398 (N_15398,N_13055,N_11884);
and U15399 (N_15399,N_14947,N_13451);
nand U15400 (N_15400,N_10684,N_12418);
or U15401 (N_15401,N_12968,N_11930);
or U15402 (N_15402,N_13047,N_11055);
nor U15403 (N_15403,N_12024,N_13059);
nand U15404 (N_15404,N_11714,N_12462);
nand U15405 (N_15405,N_13661,N_12186);
nand U15406 (N_15406,N_13927,N_13584);
nor U15407 (N_15407,N_11831,N_12667);
or U15408 (N_15408,N_12522,N_10220);
nand U15409 (N_15409,N_13845,N_11604);
or U15410 (N_15410,N_10297,N_11624);
nor U15411 (N_15411,N_14878,N_12126);
nor U15412 (N_15412,N_10876,N_12723);
nand U15413 (N_15413,N_11526,N_10152);
or U15414 (N_15414,N_10685,N_12984);
nor U15415 (N_15415,N_10945,N_11411);
nor U15416 (N_15416,N_10329,N_10908);
or U15417 (N_15417,N_11916,N_13013);
nor U15418 (N_15418,N_13062,N_14535);
and U15419 (N_15419,N_11161,N_14492);
nand U15420 (N_15420,N_13875,N_14197);
or U15421 (N_15421,N_13170,N_11910);
nand U15422 (N_15422,N_13110,N_11352);
or U15423 (N_15423,N_13572,N_12410);
nand U15424 (N_15424,N_13413,N_13544);
or U15425 (N_15425,N_11039,N_12301);
and U15426 (N_15426,N_14500,N_12291);
nor U15427 (N_15427,N_11918,N_10498);
or U15428 (N_15428,N_13087,N_14705);
nor U15429 (N_15429,N_11263,N_14858);
or U15430 (N_15430,N_11931,N_14400);
nor U15431 (N_15431,N_14431,N_12445);
nand U15432 (N_15432,N_13318,N_11673);
nor U15433 (N_15433,N_13198,N_10424);
nor U15434 (N_15434,N_14618,N_14626);
or U15435 (N_15435,N_11635,N_11467);
nand U15436 (N_15436,N_11649,N_12773);
or U15437 (N_15437,N_14525,N_11656);
nor U15438 (N_15438,N_13752,N_10073);
nand U15439 (N_15439,N_11670,N_13698);
and U15440 (N_15440,N_14171,N_12046);
or U15441 (N_15441,N_11908,N_11107);
nor U15442 (N_15442,N_13851,N_13014);
and U15443 (N_15443,N_14364,N_10344);
and U15444 (N_15444,N_10092,N_10189);
or U15445 (N_15445,N_10359,N_10666);
nand U15446 (N_15446,N_10953,N_14801);
nor U15447 (N_15447,N_10337,N_14879);
and U15448 (N_15448,N_12306,N_10173);
nor U15449 (N_15449,N_14617,N_12674);
or U15450 (N_15450,N_12904,N_11345);
and U15451 (N_15451,N_13079,N_11122);
or U15452 (N_15452,N_11805,N_11310);
nand U15453 (N_15453,N_14308,N_13153);
nand U15454 (N_15454,N_12683,N_14251);
and U15455 (N_15455,N_12903,N_10553);
nor U15456 (N_15456,N_10490,N_13112);
nor U15457 (N_15457,N_13325,N_10094);
or U15458 (N_15458,N_11387,N_14682);
and U15459 (N_15459,N_10905,N_13837);
and U15460 (N_15460,N_11257,N_10556);
nor U15461 (N_15461,N_14097,N_10160);
nor U15462 (N_15462,N_14936,N_12141);
or U15463 (N_15463,N_11260,N_10240);
nand U15464 (N_15464,N_12780,N_12196);
or U15465 (N_15465,N_14315,N_13914);
or U15466 (N_15466,N_14601,N_10414);
nand U15467 (N_15467,N_14382,N_11720);
and U15468 (N_15468,N_12467,N_13419);
nor U15469 (N_15469,N_11945,N_14992);
and U15470 (N_15470,N_14706,N_14388);
nor U15471 (N_15471,N_12733,N_12165);
or U15472 (N_15472,N_10754,N_12644);
and U15473 (N_15473,N_10998,N_11004);
and U15474 (N_15474,N_13147,N_12669);
nand U15475 (N_15475,N_14481,N_11778);
and U15476 (N_15476,N_14169,N_13569);
nand U15477 (N_15477,N_13431,N_10954);
nor U15478 (N_15478,N_10902,N_14142);
xor U15479 (N_15479,N_11798,N_10138);
nor U15480 (N_15480,N_11211,N_12042);
nor U15481 (N_15481,N_11689,N_13435);
and U15482 (N_15482,N_14436,N_11357);
nor U15483 (N_15483,N_12417,N_13120);
and U15484 (N_15484,N_10588,N_13333);
or U15485 (N_15485,N_14872,N_14799);
or U15486 (N_15486,N_11275,N_14579);
or U15487 (N_15487,N_10143,N_13136);
nand U15488 (N_15488,N_13277,N_13460);
or U15489 (N_15489,N_13429,N_12698);
and U15490 (N_15490,N_14042,N_14305);
nor U15491 (N_15491,N_14300,N_14980);
nor U15492 (N_15492,N_11367,N_13406);
and U15493 (N_15493,N_14491,N_11439);
nor U15494 (N_15494,N_13986,N_14119);
nand U15495 (N_15495,N_10516,N_11461);
or U15496 (N_15496,N_12276,N_13156);
nor U15497 (N_15497,N_10140,N_13058);
or U15498 (N_15498,N_11903,N_12902);
or U15499 (N_15499,N_10422,N_14887);
nand U15500 (N_15500,N_11965,N_11306);
nor U15501 (N_15501,N_11209,N_10036);
or U15502 (N_15502,N_11640,N_10318);
and U15503 (N_15503,N_12595,N_10310);
nor U15504 (N_15504,N_14620,N_14520);
xor U15505 (N_15505,N_10100,N_11787);
nor U15506 (N_15506,N_14681,N_14061);
nor U15507 (N_15507,N_10346,N_12399);
nor U15508 (N_15508,N_12923,N_13556);
or U15509 (N_15509,N_11022,N_11730);
or U15510 (N_15510,N_10280,N_11765);
nand U15511 (N_15511,N_14022,N_13720);
nor U15512 (N_15512,N_14457,N_10895);
and U15513 (N_15513,N_14380,N_14753);
nor U15514 (N_15514,N_13745,N_12685);
nor U15515 (N_15515,N_13200,N_14435);
nor U15516 (N_15516,N_13739,N_14965);
or U15517 (N_15517,N_11922,N_13688);
or U15518 (N_15518,N_11394,N_11087);
nand U15519 (N_15519,N_11492,N_12660);
or U15520 (N_15520,N_12871,N_14989);
nor U15521 (N_15521,N_14639,N_10784);
or U15522 (N_15522,N_12015,N_11912);
and U15523 (N_15523,N_10645,N_14970);
nor U15524 (N_15524,N_12266,N_12147);
and U15525 (N_15525,N_11794,N_14526);
nor U15526 (N_15526,N_11136,N_13339);
and U15527 (N_15527,N_10514,N_11815);
or U15528 (N_15528,N_14275,N_11013);
or U15529 (N_15529,N_10300,N_12726);
and U15530 (N_15530,N_14961,N_12628);
nand U15531 (N_15531,N_11530,N_14769);
or U15532 (N_15532,N_13528,N_14959);
nand U15533 (N_15533,N_14395,N_11085);
nand U15534 (N_15534,N_11407,N_14720);
nor U15535 (N_15535,N_14780,N_13930);
nand U15536 (N_15536,N_10881,N_11804);
nand U15537 (N_15537,N_13599,N_10760);
nor U15538 (N_15538,N_14653,N_12161);
or U15539 (N_15539,N_14670,N_11127);
nand U15540 (N_15540,N_14685,N_10525);
and U15541 (N_15541,N_13501,N_11252);
and U15542 (N_15542,N_13051,N_11259);
and U15543 (N_15543,N_13177,N_11114);
nand U15544 (N_15544,N_14813,N_13877);
or U15545 (N_15545,N_14569,N_12137);
nor U15546 (N_15546,N_10139,N_12044);
nor U15547 (N_15547,N_11065,N_11534);
nor U15548 (N_15548,N_11944,N_10209);
nand U15549 (N_15549,N_11650,N_12805);
nor U15550 (N_15550,N_10438,N_12582);
or U15551 (N_15551,N_12156,N_13710);
nor U15552 (N_15552,N_11062,N_10187);
and U15553 (N_15553,N_10376,N_10702);
nand U15554 (N_15554,N_11799,N_11704);
or U15555 (N_15555,N_13256,N_11738);
and U15556 (N_15556,N_11170,N_11846);
and U15557 (N_15557,N_10180,N_13075);
or U15558 (N_15558,N_10272,N_12101);
or U15559 (N_15559,N_14227,N_13117);
nor U15560 (N_15560,N_10583,N_11000);
or U15561 (N_15561,N_12373,N_10948);
and U15562 (N_15562,N_13264,N_12209);
and U15563 (N_15563,N_11609,N_12565);
nor U15564 (N_15564,N_11978,N_12074);
nor U15565 (N_15565,N_12389,N_13887);
or U15566 (N_15566,N_12655,N_10055);
nor U15567 (N_15567,N_10004,N_14489);
nand U15568 (N_15568,N_13747,N_14237);
and U15569 (N_15569,N_12271,N_14450);
nor U15570 (N_15570,N_14589,N_11575);
nand U15571 (N_15571,N_10649,N_13861);
or U15572 (N_15572,N_10365,N_10324);
or U15573 (N_15573,N_11679,N_14167);
nor U15574 (N_15574,N_11248,N_11675);
or U15575 (N_15575,N_10257,N_11064);
or U15576 (N_15576,N_11801,N_14329);
nor U15577 (N_15577,N_11438,N_12007);
and U15578 (N_15578,N_12831,N_14571);
and U15579 (N_15579,N_11195,N_12194);
or U15580 (N_15580,N_12323,N_10797);
nand U15581 (N_15581,N_10820,N_11587);
or U15582 (N_15582,N_14825,N_11116);
and U15583 (N_15583,N_13502,N_13275);
nor U15584 (N_15584,N_14598,N_10085);
nor U15585 (N_15585,N_13077,N_11299);
and U15586 (N_15586,N_12846,N_14083);
and U15587 (N_15587,N_11887,N_13272);
or U15588 (N_15588,N_10212,N_12925);
and U15589 (N_15589,N_10522,N_12224);
nor U15590 (N_15590,N_12482,N_11406);
and U15591 (N_15591,N_14281,N_11625);
nor U15592 (N_15592,N_13488,N_10557);
nand U15593 (N_15593,N_13412,N_11705);
and U15594 (N_15594,N_13409,N_14063);
and U15595 (N_15595,N_12691,N_11052);
or U15596 (N_15596,N_10793,N_10410);
nand U15597 (N_15597,N_13981,N_10660);
and U15598 (N_15598,N_10719,N_12449);
and U15599 (N_15599,N_13955,N_12234);
nor U15600 (N_15600,N_12741,N_10012);
nor U15601 (N_15601,N_10338,N_14507);
nor U15602 (N_15602,N_10551,N_11685);
and U15603 (N_15603,N_10544,N_10507);
and U15604 (N_15604,N_10769,N_12949);
nand U15605 (N_15605,N_12484,N_11479);
and U15606 (N_15606,N_13304,N_14938);
xor U15607 (N_15607,N_13015,N_10922);
nor U15608 (N_15608,N_12758,N_12578);
nand U15609 (N_15609,N_13164,N_10067);
or U15610 (N_15610,N_14332,N_13629);
nand U15611 (N_15611,N_13906,N_14544);
xnor U15612 (N_15612,N_13826,N_12729);
and U15613 (N_15613,N_13303,N_13010);
nor U15614 (N_15614,N_13232,N_11202);
and U15615 (N_15615,N_12416,N_10232);
nor U15616 (N_15616,N_11210,N_13179);
and U15617 (N_15617,N_11386,N_13676);
nand U15618 (N_15618,N_12921,N_11947);
nor U15619 (N_15619,N_13626,N_13774);
nand U15620 (N_15620,N_13899,N_13973);
nor U15621 (N_15621,N_10963,N_11466);
and U15622 (N_15622,N_12849,N_10847);
or U15623 (N_15623,N_14335,N_12448);
or U15624 (N_15624,N_10860,N_12884);
nand U15625 (N_15625,N_13526,N_10665);
nand U15626 (N_15626,N_11766,N_14363);
or U15627 (N_15627,N_14066,N_14148);
or U15628 (N_15628,N_11527,N_12084);
nor U15629 (N_15629,N_13765,N_11615);
and U15630 (N_15630,N_14859,N_13102);
nor U15631 (N_15631,N_13631,N_12890);
nand U15632 (N_15632,N_14943,N_13974);
and U15633 (N_15633,N_11462,N_12621);
or U15634 (N_15634,N_13377,N_10503);
nand U15635 (N_15635,N_14040,N_11403);
or U15636 (N_15636,N_11589,N_12385);
nor U15637 (N_15637,N_11001,N_12208);
or U15638 (N_15638,N_14646,N_14008);
or U15639 (N_15639,N_14250,N_11143);
and U15640 (N_15640,N_12384,N_14252);
nand U15641 (N_15641,N_10206,N_10613);
or U15642 (N_15642,N_10621,N_13384);
nor U15643 (N_15643,N_11590,N_10104);
nor U15644 (N_15644,N_13189,N_11274);
or U15645 (N_15645,N_13806,N_12962);
nor U15646 (N_15646,N_11885,N_14143);
and U15647 (N_15647,N_12328,N_14101);
or U15648 (N_15648,N_11703,N_13041);
or U15649 (N_15649,N_14534,N_12761);
and U15650 (N_15650,N_12386,N_13132);
or U15651 (N_15651,N_10416,N_12511);
nand U15652 (N_15652,N_11086,N_13494);
nand U15653 (N_15653,N_13288,N_14116);
nand U15654 (N_15654,N_10217,N_10298);
nor U15655 (N_15655,N_10720,N_11504);
nand U15656 (N_15656,N_11878,N_11241);
or U15657 (N_15657,N_11418,N_14742);
nor U15658 (N_15658,N_10205,N_13298);
nor U15659 (N_15659,N_13645,N_10002);
nand U15660 (N_15660,N_13389,N_10926);
nand U15661 (N_15661,N_13085,N_11495);
or U15662 (N_15662,N_14176,N_13539);
nand U15663 (N_15663,N_14408,N_10841);
nand U15664 (N_15664,N_12825,N_11444);
or U15665 (N_15665,N_12555,N_11167);
and U15666 (N_15666,N_10113,N_10267);
nor U15667 (N_15667,N_14926,N_12133);
or U15668 (N_15668,N_14939,N_10799);
or U15669 (N_15669,N_11827,N_11307);
xnor U15670 (N_15670,N_10141,N_14056);
nor U15671 (N_15671,N_14255,N_11581);
nand U15672 (N_15672,N_11668,N_12040);
or U15673 (N_15673,N_10366,N_14180);
nand U15674 (N_15674,N_10136,N_13236);
nor U15675 (N_15675,N_10328,N_12214);
and U15676 (N_15676,N_12979,N_11928);
nand U15677 (N_15677,N_13158,N_13603);
or U15678 (N_15678,N_12587,N_11279);
xnor U15679 (N_15679,N_12702,N_12382);
or U15680 (N_15680,N_11018,N_10643);
or U15681 (N_15681,N_10574,N_10604);
or U15682 (N_15682,N_10834,N_10064);
nand U15683 (N_15683,N_13366,N_14545);
or U15684 (N_15684,N_14287,N_14090);
nand U15685 (N_15685,N_13564,N_10743);
nand U15686 (N_15686,N_14152,N_10589);
nand U15687 (N_15687,N_14712,N_13499);
and U15688 (N_15688,N_12218,N_10681);
or U15689 (N_15689,N_13019,N_12251);
and U15690 (N_15690,N_14330,N_10188);
nand U15691 (N_15691,N_12173,N_13934);
and U15692 (N_15692,N_14751,N_14254);
nand U15693 (N_15693,N_12607,N_12256);
or U15694 (N_15694,N_13324,N_11033);
nor U15695 (N_15695,N_12220,N_11010);
or U15696 (N_15696,N_12440,N_12838);
nor U15697 (N_15697,N_11830,N_11877);
nand U15698 (N_15698,N_13176,N_13306);
nand U15699 (N_15699,N_10391,N_12869);
and U15700 (N_15700,N_10077,N_11133);
or U15701 (N_15701,N_10195,N_14509);
nand U15702 (N_15702,N_10773,N_14019);
nand U15703 (N_15703,N_11375,N_10846);
nor U15704 (N_15704,N_10960,N_14155);
or U15705 (N_15705,N_12709,N_14442);
nor U15706 (N_15706,N_11459,N_13969);
or U15707 (N_15707,N_14625,N_11921);
nand U15708 (N_15708,N_12480,N_11977);
or U15709 (N_15709,N_14673,N_11839);
or U15710 (N_15710,N_14039,N_11076);
and U15711 (N_15711,N_12176,N_14272);
nand U15712 (N_15712,N_14239,N_14950);
nor U15713 (N_15713,N_13292,N_14085);
nor U15714 (N_15714,N_11034,N_13338);
nor U15715 (N_15715,N_12043,N_14969);
nor U15716 (N_15716,N_13617,N_12069);
nand U15717 (N_15717,N_12946,N_10955);
nand U15718 (N_15718,N_13797,N_12474);
nand U15719 (N_15719,N_12483,N_14533);
or U15720 (N_15720,N_12891,N_14102);
nor U15721 (N_15721,N_10145,N_10804);
nand U15722 (N_15722,N_14012,N_11608);
nand U15723 (N_15723,N_13716,N_12115);
xor U15724 (N_15724,N_12135,N_12393);
or U15725 (N_15725,N_10755,N_13379);
or U15726 (N_15726,N_10590,N_13980);
and U15727 (N_15727,N_14708,N_11613);
nand U15728 (N_15728,N_11661,N_10400);
or U15729 (N_15729,N_11123,N_10591);
nand U15730 (N_15730,N_11268,N_12728);
nand U15731 (N_15731,N_14146,N_11614);
nor U15732 (N_15732,N_14473,N_11881);
nand U15733 (N_15733,N_11292,N_10952);
and U15734 (N_15734,N_14867,N_10981);
nand U15735 (N_15735,N_10561,N_13972);
or U15736 (N_15736,N_14719,N_12633);
or U15737 (N_15737,N_13408,N_10142);
nor U15738 (N_15738,N_11246,N_10677);
nand U15739 (N_15739,N_12302,N_13255);
and U15740 (N_15740,N_11706,N_12581);
or U15741 (N_15741,N_10259,N_12681);
or U15742 (N_15742,N_11014,N_14006);
and U15743 (N_15743,N_10458,N_11821);
nor U15744 (N_15744,N_13740,N_12542);
or U15745 (N_15745,N_13195,N_13516);
or U15746 (N_15746,N_14134,N_12292);
nand U15747 (N_15747,N_12961,N_12356);
xor U15748 (N_15748,N_11929,N_11280);
and U15749 (N_15749,N_10348,N_14531);
xnor U15750 (N_15750,N_12744,N_11355);
nor U15751 (N_15751,N_10119,N_14051);
and U15752 (N_15752,N_12171,N_12735);
or U15753 (N_15753,N_14312,N_11756);
nand U15754 (N_15754,N_12022,N_12603);
nand U15755 (N_15755,N_13309,N_12584);
nand U15756 (N_15756,N_13689,N_13822);
nor U15757 (N_15757,N_10486,N_12790);
nand U15758 (N_15758,N_14633,N_13705);
and U15759 (N_15759,N_12258,N_10454);
nand U15760 (N_15760,N_10931,N_11645);
or U15761 (N_15761,N_11147,N_14661);
or U15762 (N_15762,N_13687,N_13035);
nand U15763 (N_15763,N_12223,N_14475);
or U15764 (N_15764,N_11718,N_13373);
nor U15765 (N_15765,N_10009,N_10056);
and U15766 (N_15766,N_12899,N_14229);
or U15767 (N_15767,N_13618,N_12606);
nand U15768 (N_15768,N_12975,N_10708);
nor U15769 (N_15769,N_10364,N_12279);
nand U15770 (N_15770,N_11360,N_14323);
nand U15771 (N_15771,N_11069,N_10870);
nand U15772 (N_15772,N_12743,N_11359);
or U15773 (N_15773,N_11883,N_11369);
nor U15774 (N_15774,N_10247,N_14407);
or U15775 (N_15775,N_14732,N_11012);
or U15776 (N_15776,N_10115,N_10107);
and U15777 (N_15777,N_12094,N_14547);
nand U15778 (N_15778,N_12326,N_10568);
or U15779 (N_15779,N_12605,N_13505);
or U15780 (N_15780,N_12052,N_14973);
nand U15781 (N_15781,N_13697,N_11421);
nand U15782 (N_15782,N_11636,N_14484);
or U15783 (N_15783,N_12608,N_11841);
nor U15784 (N_15784,N_13234,N_14107);
nand U15785 (N_15785,N_14115,N_11546);
nand U15786 (N_15786,N_14161,N_12870);
nand U15787 (N_15787,N_11175,N_14132);
nor U15788 (N_15788,N_13616,N_10111);
nand U15789 (N_15789,N_14151,N_10437);
or U15790 (N_15790,N_12827,N_12783);
nand U15791 (N_15791,N_12760,N_10543);
nand U15792 (N_15792,N_13621,N_13050);
and U15793 (N_15793,N_13954,N_10221);
nand U15794 (N_15794,N_14374,N_11750);
and U15795 (N_15795,N_14173,N_14744);
xnor U15796 (N_15796,N_13840,N_14029);
or U15797 (N_15797,N_10547,N_14326);
or U15798 (N_15798,N_14506,N_11540);
nand U15799 (N_15799,N_13956,N_12933);
and U15800 (N_15800,N_10821,N_13184);
nor U15801 (N_15801,N_10879,N_14645);
nor U15802 (N_15802,N_10794,N_10951);
or U15803 (N_15803,N_12797,N_13842);
and U15804 (N_15804,N_11487,N_10214);
nand U15805 (N_15805,N_11680,N_12791);
and U15806 (N_15806,N_10810,N_12647);
and U15807 (N_15807,N_11208,N_12970);
and U15808 (N_15808,N_10802,N_11989);
or U15809 (N_15809,N_13046,N_13563);
nand U15810 (N_15810,N_10001,N_14241);
and U15811 (N_15811,N_10223,N_14361);
or U15812 (N_15812,N_11550,N_10048);
or U15813 (N_15813,N_14316,N_10097);
nand U15814 (N_15814,N_11776,N_12588);
or U15815 (N_15815,N_13400,N_10144);
nor U15816 (N_15816,N_14456,N_12752);
and U15817 (N_15817,N_14105,N_12378);
or U15818 (N_15818,N_13790,N_13067);
and U15819 (N_15819,N_14964,N_12671);
nand U15820 (N_15820,N_12640,N_14510);
or U15821 (N_15821,N_10933,N_10638);
nand U15822 (N_15822,N_14523,N_10920);
nand U15823 (N_15823,N_11119,N_10550);
and U15824 (N_15824,N_14577,N_12568);
or U15825 (N_15825,N_13022,N_14433);
and U15826 (N_15826,N_14912,N_14389);
nand U15827 (N_15827,N_11859,N_14955);
nand U15828 (N_15828,N_11365,N_12456);
nand U15829 (N_15829,N_12114,N_10150);
nand U15830 (N_15830,N_11865,N_10236);
and U15831 (N_15831,N_14774,N_11073);
and U15832 (N_15832,N_14782,N_14234);
or U15833 (N_15833,N_14638,N_10351);
or U15834 (N_15834,N_13987,N_12381);
nor U15835 (N_15835,N_13374,N_10445);
or U15836 (N_15836,N_10233,N_10776);
nor U15837 (N_15837,N_12355,N_14956);
nor U15838 (N_15838,N_13876,N_10213);
or U15839 (N_15839,N_11772,N_13116);
and U15840 (N_15840,N_13082,N_12756);
or U15841 (N_15841,N_14972,N_12808);
and U15842 (N_15842,N_12473,N_10900);
or U15843 (N_15843,N_13680,N_11612);
nor U15844 (N_15844,N_11205,N_10674);
or U15845 (N_15845,N_14076,N_11866);
nor U15846 (N_15846,N_13646,N_14869);
or U15847 (N_15847,N_14342,N_12550);
nor U15848 (N_15848,N_13326,N_11067);
or U15849 (N_15849,N_11996,N_11316);
and U15850 (N_15850,N_13507,N_14331);
nor U15851 (N_15851,N_13428,N_12537);
or U15852 (N_15852,N_13735,N_12501);
or U15853 (N_15853,N_13643,N_14014);
or U15854 (N_15854,N_10315,N_11267);
and U15855 (N_15855,N_10696,N_12283);
nand U15856 (N_15856,N_12955,N_14402);
or U15857 (N_15857,N_10239,N_14414);
and U15858 (N_15858,N_11572,N_10215);
and U15859 (N_15859,N_12036,N_14003);
or U15860 (N_15860,N_11449,N_10816);
nor U15861 (N_15861,N_11448,N_12433);
nand U15862 (N_15862,N_12905,N_10283);
or U15863 (N_15863,N_10673,N_13615);
nor U15864 (N_15864,N_12820,N_11602);
and U15865 (N_15865,N_13222,N_13276);
or U15866 (N_15866,N_13628,N_10620);
nor U15867 (N_15867,N_10435,N_10584);
nand U15868 (N_15868,N_13924,N_11149);
nand U15869 (N_15869,N_10017,N_10844);
nor U15870 (N_15870,N_13771,N_13135);
and U15871 (N_15871,N_14536,N_13417);
or U15872 (N_15872,N_10360,N_11642);
or U15873 (N_15873,N_13786,N_12521);
and U15874 (N_15874,N_14153,N_13263);
nand U15875 (N_15875,N_12058,N_10039);
nand U15876 (N_15876,N_12211,N_12246);
or U15877 (N_15877,N_13253,N_10325);
nor U15878 (N_15878,N_11811,N_11247);
nor U15879 (N_15879,N_11192,N_11200);
or U15880 (N_15880,N_11567,N_13481);
nor U15881 (N_15881,N_11998,N_12221);
nand U15882 (N_15882,N_11408,N_14067);
nor U15883 (N_15883,N_11942,N_13278);
nor U15884 (N_15884,N_10789,N_12799);
or U15885 (N_15885,N_10156,N_11168);
and U15886 (N_15886,N_12078,N_11582);
and U15887 (N_15887,N_12420,N_10530);
xnor U15888 (N_15888,N_12230,N_14900);
or U15889 (N_15889,N_14898,N_13321);
nand U15890 (N_15890,N_11734,N_12512);
nor U15891 (N_15891,N_10636,N_11924);
or U15892 (N_15892,N_14605,N_14922);
nand U15893 (N_15893,N_10090,N_13336);
xnor U15894 (N_15894,N_13279,N_13099);
nor U15895 (N_15895,N_11025,N_11023);
and U15896 (N_15896,N_13757,N_11627);
nand U15897 (N_15897,N_12965,N_10883);
or U15898 (N_15898,N_11007,N_11974);
and U15899 (N_15899,N_14488,N_14448);
nor U15900 (N_15900,N_10552,N_10595);
and U15901 (N_15901,N_11888,N_10786);
nor U15902 (N_15902,N_11752,N_13259);
nor U15903 (N_15903,N_12097,N_13866);
nand U15904 (N_15904,N_10251,N_10332);
nand U15905 (N_15905,N_11327,N_12377);
nand U15906 (N_15906,N_14434,N_12510);
nor U15907 (N_15907,N_14428,N_13886);
nand U15908 (N_15908,N_14149,N_10476);
nand U15909 (N_15909,N_14674,N_10197);
or U15910 (N_15910,N_11079,N_13769);
nand U15911 (N_15911,N_12431,N_12423);
xor U15912 (N_15912,N_11113,N_12972);
or U15913 (N_15913,N_10826,N_10287);
nand U15914 (N_15914,N_14641,N_11011);
nor U15915 (N_15915,N_11676,N_14990);
or U15916 (N_15916,N_12823,N_13846);
nand U15917 (N_15917,N_11380,N_10025);
or U15918 (N_15918,N_11218,N_13641);
and U15919 (N_15919,N_11509,N_12786);
nor U15920 (N_15920,N_10930,N_14225);
nor U15921 (N_15921,N_14233,N_13240);
and U15922 (N_15922,N_12407,N_11181);
nor U15923 (N_15923,N_14791,N_14138);
nor U15924 (N_15924,N_12387,N_14392);
nor U15925 (N_15925,N_12390,N_10040);
xnor U15926 (N_15926,N_13751,N_10885);
nand U15927 (N_15927,N_14211,N_12282);
or U15928 (N_15928,N_14854,N_14189);
nand U15929 (N_15929,N_13884,N_13248);
nor U15930 (N_15930,N_10018,N_11951);
nor U15931 (N_15931,N_13057,N_10646);
nand U15932 (N_15932,N_13659,N_13197);
nand U15933 (N_15933,N_10991,N_13375);
nand U15934 (N_15934,N_12842,N_13480);
or U15935 (N_15935,N_11619,N_12268);
nand U15936 (N_15936,N_13728,N_12717);
and U15937 (N_15937,N_12615,N_11555);
and U15938 (N_15938,N_13076,N_14952);
nand U15939 (N_15939,N_10670,N_12330);
nor U15940 (N_15940,N_14159,N_12338);
and U15941 (N_15941,N_11900,N_10923);
nand U15942 (N_15942,N_11294,N_13908);
or U15943 (N_15943,N_12738,N_14416);
xnor U15944 (N_15944,N_12817,N_13779);
or U15945 (N_15945,N_12742,N_13574);
nand U15946 (N_15946,N_13246,N_11904);
and U15947 (N_15947,N_11925,N_12453);
nand U15948 (N_15948,N_11186,N_13471);
nor U15949 (N_15949,N_10170,N_10079);
nor U15950 (N_15950,N_14553,N_14210);
and U15951 (N_15951,N_12191,N_12907);
and U15952 (N_15952,N_12851,N_10698);
nor U15953 (N_15953,N_13187,N_13996);
nor U15954 (N_15954,N_12206,N_11368);
or U15955 (N_15955,N_11111,N_12244);
nor U15956 (N_15956,N_12425,N_10352);
and U15957 (N_15957,N_11536,N_10912);
nand U15958 (N_15958,N_13800,N_13397);
and U15959 (N_15959,N_10418,N_11350);
and U15960 (N_15960,N_14306,N_13299);
nand U15961 (N_15961,N_11505,N_11105);
and U15962 (N_15962,N_13446,N_14309);
or U15963 (N_15963,N_13310,N_10118);
and U15964 (N_15964,N_12217,N_14707);
and U15965 (N_15965,N_11824,N_11933);
nor U15966 (N_15966,N_13825,N_14643);
and U15967 (N_15967,N_11748,N_13950);
and U15968 (N_15968,N_10813,N_10398);
or U15969 (N_15969,N_11822,N_11829);
and U15970 (N_15970,N_14027,N_11084);
and U15971 (N_15971,N_13206,N_14137);
nand U15972 (N_15972,N_10124,N_12411);
nor U15973 (N_15973,N_12620,N_12216);
or U15974 (N_15974,N_12439,N_13395);
nand U15975 (N_15975,N_14084,N_13016);
nand U15976 (N_15976,N_14919,N_14717);
nand U15977 (N_15977,N_11251,N_11639);
and U15978 (N_15978,N_14081,N_12294);
nand U15979 (N_15979,N_10234,N_11041);
or U15980 (N_15980,N_11199,N_10227);
nor U15981 (N_15981,N_11452,N_12375);
nor U15982 (N_15982,N_12363,N_13007);
or U15983 (N_15983,N_11349,N_14957);
or U15984 (N_15984,N_11771,N_12170);
nor U15985 (N_15985,N_11810,N_11040);
nand U15986 (N_15986,N_14578,N_13893);
nor U15987 (N_15987,N_13302,N_12832);
nand U15988 (N_15988,N_12160,N_10644);
or U15989 (N_15989,N_14834,N_10520);
nor U15990 (N_15990,N_12794,N_13003);
or U15991 (N_15991,N_14182,N_14325);
xnor U15992 (N_15992,N_13597,N_14595);
nand U15993 (N_15993,N_11298,N_11060);
and U15994 (N_15994,N_13593,N_11061);
nand U15995 (N_15995,N_14561,N_11809);
nand U15996 (N_15996,N_12250,N_13931);
nand U15997 (N_15997,N_14884,N_12107);
nor U15998 (N_15998,N_14471,N_11237);
nor U15999 (N_15999,N_11063,N_10290);
and U16000 (N_16000,N_12927,N_11674);
nor U16001 (N_16001,N_14580,N_14073);
and U16002 (N_16002,N_10363,N_12986);
nand U16003 (N_16003,N_11709,N_14122);
xnor U16004 (N_16004,N_12459,N_12755);
or U16005 (N_16005,N_12331,N_12942);
nor U16006 (N_16006,N_13900,N_14563);
nor U16007 (N_16007,N_12368,N_10330);
or U16008 (N_16008,N_10481,N_11044);
nor U16009 (N_16009,N_13436,N_12152);
nand U16010 (N_16010,N_12976,N_12090);
or U16011 (N_16011,N_11266,N_13161);
nand U16012 (N_16012,N_11595,N_14011);
and U16013 (N_16013,N_13154,N_14421);
and U16014 (N_16014,N_13788,N_12120);
and U16015 (N_16015,N_10043,N_12198);
or U16016 (N_16016,N_13452,N_11440);
nor U16017 (N_16017,N_12492,N_12366);
nor U16018 (N_16018,N_14158,N_10286);
nand U16019 (N_16019,N_10730,N_11422);
nor U16020 (N_16020,N_13393,N_13753);
nand U16021 (N_16021,N_14868,N_14214);
nor U16022 (N_16022,N_10478,N_12546);
nand U16023 (N_16023,N_11906,N_13622);
nor U16024 (N_16024,N_11897,N_12960);
or U16025 (N_16025,N_12873,N_12875);
and U16026 (N_16026,N_13095,N_11969);
nand U16027 (N_16027,N_13860,N_14222);
nor U16028 (N_16028,N_11496,N_13857);
nor U16029 (N_16029,N_13959,N_10049);
or U16030 (N_16030,N_14828,N_10798);
and U16031 (N_16031,N_10350,N_10401);
and U16032 (N_16032,N_11538,N_11198);
nor U16033 (N_16033,N_13356,N_13273);
nand U16034 (N_16034,N_11950,N_13459);
nand U16035 (N_16035,N_14711,N_13512);
nor U16036 (N_16036,N_12722,N_12333);
nand U16037 (N_16037,N_12504,N_12573);
and U16038 (N_16038,N_12025,N_13686);
nor U16039 (N_16039,N_14327,N_11621);
or U16040 (N_16040,N_10652,N_10959);
nand U16041 (N_16041,N_14914,N_13612);
or U16042 (N_16042,N_14147,N_12163);
and U16043 (N_16043,N_11453,N_12656);
nand U16044 (N_16044,N_12123,N_11638);
or U16045 (N_16045,N_12360,N_11678);
nor U16046 (N_16046,N_10679,N_13719);
nand U16047 (N_16047,N_13418,N_12713);
nand U16048 (N_16048,N_11501,N_11622);
or U16049 (N_16049,N_11337,N_14218);
and U16050 (N_16050,N_13223,N_14786);
nor U16051 (N_16051,N_14381,N_12419);
nor U16052 (N_16052,N_10499,N_12796);
nand U16053 (N_16053,N_14278,N_10443);
and U16054 (N_16054,N_12269,N_11515);
and U16055 (N_16055,N_13100,N_10166);
and U16056 (N_16056,N_10707,N_10182);
or U16057 (N_16057,N_12050,N_13937);
and U16058 (N_16058,N_11228,N_12129);
or U16059 (N_16059,N_14849,N_13101);
nand U16060 (N_16060,N_13873,N_10984);
and U16061 (N_16061,N_12088,N_11543);
nor U16062 (N_16062,N_11666,N_13194);
or U16063 (N_16063,N_10578,N_10629);
xor U16064 (N_16064,N_12275,N_11681);
and U16065 (N_16065,N_11092,N_10082);
nand U16066 (N_16066,N_12394,N_13097);
nor U16067 (N_16067,N_12765,N_12297);
nand U16068 (N_16068,N_10857,N_10863);
or U16069 (N_16069,N_12840,N_13783);
nor U16070 (N_16070,N_14597,N_13449);
or U16071 (N_16071,N_10327,N_12571);
nand U16072 (N_16072,N_13345,N_10637);
or U16073 (N_16073,N_12130,N_14713);
nor U16074 (N_16074,N_10446,N_10014);
nand U16075 (N_16075,N_10687,N_13590);
and U16076 (N_16076,N_14794,N_11875);
and U16077 (N_16077,N_14846,N_12816);
nor U16078 (N_16078,N_14268,N_14654);
and U16079 (N_16079,N_12528,N_13157);
or U16080 (N_16080,N_14552,N_14458);
nand U16081 (N_16081,N_12841,N_11962);
or U16082 (N_16082,N_14731,N_14131);
nor U16083 (N_16083,N_14529,N_12388);
nor U16084 (N_16084,N_11755,N_14749);
or U16085 (N_16085,N_13407,N_10367);
and U16086 (N_16086,N_11913,N_11828);
nand U16087 (N_16087,N_13173,N_14417);
or U16088 (N_16088,N_12159,N_12830);
nor U16089 (N_16089,N_10864,N_10722);
nand U16090 (N_16090,N_11735,N_11891);
nor U16091 (N_16091,N_10582,N_12203);
nor U16092 (N_16092,N_14377,N_14636);
or U16093 (N_16093,N_11683,N_13186);
nor U16094 (N_16094,N_11570,N_10439);
nor U16095 (N_16095,N_11229,N_10249);
or U16096 (N_16096,N_13096,N_13551);
nor U16097 (N_16097,N_13935,N_10335);
or U16098 (N_16098,N_14768,N_12672);
nand U16099 (N_16099,N_11682,N_11446);
nor U16100 (N_16100,N_11939,N_13297);
and U16101 (N_16101,N_13961,N_14562);
or U16102 (N_16102,N_10928,N_10540);
nor U16103 (N_16103,N_14502,N_13141);
and U16104 (N_16104,N_10277,N_12098);
nor U16105 (N_16105,N_10686,N_14334);
or U16106 (N_16106,N_11870,N_11270);
nand U16107 (N_16107,N_11493,N_14697);
nand U16108 (N_16108,N_13878,N_12139);
or U16109 (N_16109,N_12855,N_14977);
or U16110 (N_16110,N_14172,N_12458);
nor U16111 (N_16111,N_11956,N_11457);
and U16112 (N_16112,N_11158,N_10640);
and U16113 (N_16113,N_10678,N_13949);
and U16114 (N_16114,N_13693,N_13475);
and U16115 (N_16115,N_14541,N_13957);
or U16116 (N_16116,N_10536,N_14232);
nor U16117 (N_16117,N_10910,N_12853);
and U16118 (N_16118,N_13946,N_10839);
and U16119 (N_16119,N_14419,N_10037);
or U16120 (N_16120,N_13359,N_14490);
nor U16121 (N_16121,N_10921,N_12070);
and U16122 (N_16122,N_12563,N_13305);
nand U16123 (N_16123,N_10184,N_12915);
and U16124 (N_16124,N_14771,N_14178);
or U16125 (N_16125,N_13185,N_11416);
nor U16126 (N_16126,N_11304,N_12320);
and U16127 (N_16127,N_12034,N_10615);
or U16128 (N_16128,N_10925,N_12039);
nand U16129 (N_16129,N_12824,N_14934);
nand U16130 (N_16130,N_12866,N_13951);
nor U16131 (N_16131,N_10128,N_10132);
or U16132 (N_16132,N_13209,N_10783);
and U16133 (N_16133,N_13468,N_10612);
or U16134 (N_16134,N_11410,N_13044);
nor U16135 (N_16135,N_10470,N_13482);
or U16136 (N_16136,N_13090,N_12288);
nor U16137 (N_16137,N_14629,N_12345);
nor U16138 (N_16138,N_13469,N_10891);
nor U16139 (N_16139,N_11152,N_14806);
nor U16140 (N_16140,N_10066,N_13241);
nor U16141 (N_16141,N_12138,N_11434);
or U16142 (N_16142,N_11395,N_11005);
nand U16143 (N_16143,N_12651,N_14224);
and U16144 (N_16144,N_11115,N_12490);
or U16145 (N_16145,N_12012,N_11151);
nor U16146 (N_16146,N_13423,N_11700);
or U16147 (N_16147,N_12631,N_11347);
or U16148 (N_16148,N_10614,N_12318);
nand U16149 (N_16149,N_14976,N_12002);
nand U16150 (N_16150,N_12272,N_12144);
nand U16151 (N_16151,N_14648,N_10706);
or U16152 (N_16152,N_14077,N_13939);
nand U16153 (N_16153,N_10396,N_13425);
nand U16154 (N_16154,N_12357,N_14299);
nand U16155 (N_16155,N_10626,N_12701);
and U16156 (N_16156,N_10961,N_13098);
or U16157 (N_16157,N_10918,N_14128);
and U16158 (N_16158,N_13557,N_13833);
nor U16159 (N_16159,N_14735,N_11784);
and U16160 (N_16160,N_12721,N_13864);
xnor U16161 (N_16161,N_12694,N_12711);
nor U16162 (N_16162,N_14376,N_13721);
or U16163 (N_16163,N_10765,N_13447);
or U16164 (N_16164,N_10650,N_13247);
and U16165 (N_16165,N_13540,N_10432);
or U16166 (N_16166,N_10381,N_13962);
and U16167 (N_16167,N_14044,N_12035);
or U16168 (N_16168,N_12664,N_10689);
and U16169 (N_16169,N_14260,N_11129);
nor U16170 (N_16170,N_13750,N_10822);
nand U16171 (N_16171,N_12829,N_13265);
nand U16172 (N_16172,N_14860,N_14031);
nand U16173 (N_16173,N_14657,N_12564);
nand U16174 (N_16174,N_13554,N_12515);
and U16175 (N_16175,N_14996,N_13534);
nand U16176 (N_16176,N_14387,N_10901);
nand U16177 (N_16177,N_11747,N_10733);
nand U16178 (N_16178,N_10944,N_10080);
and U16179 (N_16179,N_11454,N_13856);
nor U16180 (N_16180,N_11180,N_12687);
and U16181 (N_16181,N_10586,N_13535);
or U16182 (N_16182,N_12151,N_13692);
nor U16183 (N_16183,N_14901,N_11686);
nand U16184 (N_16184,N_11958,N_13521);
nor U16185 (N_16185,N_11287,N_13300);
or U16186 (N_16186,N_13898,N_12305);
or U16187 (N_16187,N_13608,N_12642);
and U16188 (N_16188,N_13913,N_13414);
nand U16189 (N_16189,N_12270,N_13053);
and U16190 (N_16190,N_10125,N_14373);
and U16191 (N_16191,N_12690,N_10403);
or U16192 (N_16192,N_11525,N_11599);
nand U16193 (N_16193,N_10339,N_13266);
nor U16194 (N_16194,N_10842,N_14546);
nand U16195 (N_16195,N_12391,N_12913);
nand U16196 (N_16196,N_10781,N_12014);
nor U16197 (N_16197,N_14621,N_11669);
nand U16198 (N_16198,N_14410,N_10801);
nand U16199 (N_16199,N_11800,N_10571);
and U16200 (N_16200,N_10369,N_13633);
or U16201 (N_16201,N_13848,N_11920);
nand U16202 (N_16202,N_11313,N_14193);
or U16203 (N_16203,N_10872,N_12712);
and U16204 (N_16204,N_10248,N_11003);
nand U16205 (N_16205,N_11919,N_13818);
nand U16206 (N_16206,N_13282,N_11182);
or U16207 (N_16207,N_12747,N_13545);
nor U16208 (N_16208,N_10024,N_12619);
or U16209 (N_16209,N_11869,N_13785);
or U16210 (N_16210,N_11009,N_13552);
nor U16211 (N_16211,N_14282,N_13733);
nor U16212 (N_16212,N_13654,N_11882);
and U16213 (N_16213,N_10208,N_13017);
nand U16214 (N_16214,N_12862,N_10487);
and U16215 (N_16215,N_12112,N_10072);
or U16216 (N_16216,N_14406,N_14198);
or U16217 (N_16217,N_13350,N_14610);
nor U16218 (N_16218,N_10837,N_13226);
nor U16219 (N_16219,N_11844,N_11239);
and U16220 (N_16220,N_11797,N_12586);
or U16221 (N_16221,N_14140,N_10293);
nor U16222 (N_16222,N_12526,N_14508);
and U16223 (N_16223,N_14049,N_13663);
nand U16224 (N_16224,N_10717,N_11423);
and U16225 (N_16225,N_12892,N_12777);
nand U16226 (N_16226,N_13713,N_11522);
and U16227 (N_16227,N_14984,N_11736);
and U16228 (N_16228,N_12104,N_14139);
and U16229 (N_16229,N_14930,N_11607);
and U16230 (N_16230,N_12495,N_10312);
and U16231 (N_16231,N_12383,N_14647);
or U16232 (N_16232,N_11743,N_14945);
and U16233 (N_16233,N_10007,N_12103);
nand U16234 (N_16234,N_10563,N_11498);
or U16235 (N_16235,N_12293,N_14322);
and U16236 (N_16236,N_12872,N_11901);
nand U16237 (N_16237,N_13817,N_10975);
nand U16238 (N_16238,N_14611,N_10572);
and U16239 (N_16239,N_10828,N_13709);
nor U16240 (N_16240,N_10211,N_11508);
and U16241 (N_16241,N_14336,N_11016);
and U16242 (N_16242,N_13155,N_10809);
or U16243 (N_16243,N_14652,N_10123);
and U16244 (N_16244,N_12332,N_11707);
or U16245 (N_16245,N_10840,N_14691);
and U16246 (N_16246,N_12312,N_14478);
nor U16247 (N_16247,N_12348,N_13107);
nand U16248 (N_16248,N_11402,N_14722);
nor U16249 (N_16249,N_13456,N_11250);
nor U16250 (N_16250,N_14555,N_11695);
xor U16251 (N_16251,N_10409,N_11342);
nor U16252 (N_16252,N_10299,N_10165);
or U16253 (N_16253,N_12558,N_13063);
and U16254 (N_16254,N_12557,N_13793);
and U16255 (N_16255,N_10532,N_13890);
nor U16256 (N_16256,N_11563,N_10393);
and U16257 (N_16257,N_14000,N_12922);
nand U16258 (N_16258,N_11991,N_12475);
or U16259 (N_16259,N_10313,N_10059);
and U16260 (N_16260,N_12695,N_12847);
nand U16261 (N_16261,N_12549,N_14767);
nor U16262 (N_16262,N_14343,N_12233);
nand U16263 (N_16263,N_10062,N_12704);
or U16264 (N_16264,N_14062,N_11376);
and U16265 (N_16265,N_10703,N_14788);
nand U16266 (N_16266,N_14680,N_11577);
or U16267 (N_16267,N_10831,N_11071);
nand U16268 (N_16268,N_10491,N_14409);
and U16269 (N_16269,N_12803,N_11985);
nor U16270 (N_16270,N_13491,N_11833);
nand U16271 (N_16271,N_13942,N_10824);
nor U16272 (N_16272,N_11926,N_14413);
nor U16273 (N_16273,N_13787,N_11981);
or U16274 (N_16274,N_14360,N_10500);
or U16275 (N_16275,N_14958,N_11169);
nand U16276 (N_16276,N_11561,N_14057);
nor U16277 (N_16277,N_14338,N_14864);
nand U16278 (N_16278,N_10496,N_13496);
or U16279 (N_16279,N_10633,N_12516);
or U16280 (N_16280,N_11935,N_14741);
or U16281 (N_16281,N_11644,N_11348);
nand U16282 (N_16282,N_12996,N_11894);
nor U16283 (N_16283,N_14064,N_10093);
or U16284 (N_16284,N_11293,N_11058);
and U16285 (N_16285,N_12351,N_12646);
nor U16286 (N_16286,N_13070,N_10851);
and U16287 (N_16287,N_13700,N_11037);
nor U16288 (N_16288,N_13203,N_11603);
and U16289 (N_16289,N_11189,N_13993);
or U16290 (N_16290,N_11414,N_10281);
nor U16291 (N_16291,N_13791,N_10420);
nor U16292 (N_16292,N_11967,N_12049);
or U16293 (N_16293,N_14469,N_12629);
nand U16294 (N_16294,N_11469,N_14046);
or U16295 (N_16295,N_12188,N_13600);
nand U16296 (N_16296,N_10042,N_13149);
and U16297 (N_16297,N_12204,N_13828);
nor U16298 (N_16298,N_13134,N_12100);
nor U16299 (N_16299,N_14292,N_13167);
nand U16300 (N_16300,N_12336,N_13690);
and U16301 (N_16301,N_12696,N_13672);
nand U16302 (N_16302,N_11532,N_12426);
or U16303 (N_16303,N_13093,N_14303);
nand U16304 (N_16304,N_14588,N_13308);
nor U16305 (N_16305,N_13180,N_12403);
and U16306 (N_16306,N_10459,N_14186);
and U16307 (N_16307,N_11964,N_12005);
nor U16308 (N_16308,N_10609,N_13920);
and U16309 (N_16309,N_14467,N_11845);
and U16310 (N_16310,N_12737,N_14650);
nand U16311 (N_16311,N_12245,N_13560);
and U16312 (N_16312,N_10966,N_10331);
nand U16313 (N_16313,N_14050,N_12649);
and U16314 (N_16314,N_14616,N_12739);
and U16315 (N_16315,N_10752,N_14587);
nand U16316 (N_16316,N_13433,N_10980);
or U16317 (N_16317,N_10510,N_13012);
and U16318 (N_16318,N_12974,N_14129);
and U16319 (N_16319,N_14302,N_14038);
and U16320 (N_16320,N_10246,N_12809);
and U16321 (N_16321,N_12920,N_10319);
or U16322 (N_16322,N_14819,N_14393);
and U16323 (N_16323,N_14035,N_11617);
xnor U16324 (N_16324,N_10440,N_14220);
or U16325 (N_16325,N_11332,N_14995);
nand U16326 (N_16326,N_10471,N_14441);
nor U16327 (N_16327,N_10785,N_13953);
or U16328 (N_16328,N_10387,N_13191);
nand U16329 (N_16329,N_10725,N_14202);
nand U16330 (N_16330,N_14212,N_14394);
nand U16331 (N_16331,N_11430,N_12531);
and U16332 (N_16332,N_14963,N_11272);
nor U16333 (N_16333,N_13820,N_10564);
nor U16334 (N_16334,N_11852,N_13970);
or U16335 (N_16335,N_10833,N_10442);
and U16336 (N_16336,N_10988,N_13515);
nand U16337 (N_16337,N_11559,N_11130);
nor U16338 (N_16338,N_13219,N_10426);
nand U16339 (N_16339,N_11474,N_11573);
nand U16340 (N_16340,N_14071,N_10091);
and U16341 (N_16341,N_14890,N_10680);
and U16342 (N_16342,N_12982,N_10987);
nor U16343 (N_16343,N_12570,N_10168);
nand U16344 (N_16344,N_12985,N_11460);
and U16345 (N_16345,N_14117,N_11194);
and U16346 (N_16346,N_14514,N_13283);
and U16347 (N_16347,N_12523,N_10472);
or U16348 (N_16348,N_10019,N_10275);
nand U16349 (N_16349,N_12140,N_14184);
nor U16350 (N_16350,N_10639,N_13159);
nand U16351 (N_16351,N_12602,N_10126);
and U16352 (N_16352,N_13858,N_10867);
and U16353 (N_16353,N_14055,N_13391);
or U16354 (N_16354,N_13405,N_14163);
or U16355 (N_16355,N_10074,N_12527);
nor U16356 (N_16356,N_13984,N_12839);
or U16357 (N_16357,N_11796,N_10466);
and U16358 (N_16358,N_10316,N_11244);
or U16359 (N_16359,N_11584,N_14123);
nand U16360 (N_16360,N_10070,N_11711);
and U16361 (N_16361,N_10497,N_12850);
nor U16362 (N_16362,N_14993,N_10322);
xnor U16363 (N_16363,N_10518,N_13204);
or U16364 (N_16364,N_11231,N_11340);
nor U16365 (N_16365,N_13230,N_14747);
and U16366 (N_16366,N_13314,N_11315);
nor U16367 (N_16367,N_12189,N_10803);
nor U16368 (N_16368,N_11807,N_13582);
nor U16369 (N_16369,N_12757,N_10204);
nand U16370 (N_16370,N_13213,N_10676);
or U16371 (N_16371,N_11108,N_11273);
or U16372 (N_16372,N_10790,N_10714);
or U16373 (N_16373,N_12287,N_10086);
nand U16374 (N_16374,N_14058,N_10913);
nand U16375 (N_16375,N_13580,N_12929);
or U16376 (N_16376,N_11511,N_13736);
nor U16377 (N_16377,N_12017,N_10222);
or U16378 (N_16378,N_12243,N_12936);
xnor U16379 (N_16379,N_13027,N_10271);
and U16380 (N_16380,N_13555,N_12560);
or U16381 (N_16381,N_12195,N_13589);
nor U16382 (N_16382,N_13904,N_11120);
nor U16383 (N_16383,N_14024,N_11142);
nor U16384 (N_16384,N_14369,N_14853);
or U16385 (N_16385,N_13349,N_13286);
and U16386 (N_16386,N_10362,N_12437);
nand U16387 (N_16387,N_10996,N_13034);
nand U16388 (N_16388,N_14612,N_13294);
or U16389 (N_16389,N_12684,N_12030);
nor U16390 (N_16390,N_10618,N_11314);
or U16391 (N_16391,N_11436,N_14743);
nand U16392 (N_16392,N_11450,N_12497);
nand U16393 (N_16393,N_11471,N_11941);
nor U16394 (N_16394,N_13162,N_11726);
nor U16395 (N_16395,N_14429,N_10038);
nor U16396 (N_16396,N_11605,N_13463);
or U16397 (N_16397,N_11354,N_12718);
or U16398 (N_16398,N_11566,N_11854);
and U16399 (N_16399,N_11329,N_10700);
or U16400 (N_16400,N_13824,N_10764);
or U16401 (N_16401,N_10106,N_14288);
nor U16402 (N_16402,N_11481,N_12319);
or U16403 (N_16403,N_10179,N_14156);
and U16404 (N_16404,N_11020,N_13065);
nand U16405 (N_16405,N_14693,N_12947);
and U16406 (N_16406,N_10273,N_14942);
nor U16407 (N_16407,N_10766,N_12818);
nand U16408 (N_16408,N_13888,N_13853);
xor U16409 (N_16409,N_10320,N_13801);
nor U16410 (N_16410,N_13903,N_11646);
nor U16411 (N_16411,N_12678,N_11697);
and U16412 (N_16412,N_13252,N_11148);
nor U16413 (N_16413,N_11696,N_10992);
nand U16414 (N_16414,N_14501,N_14624);
or U16415 (N_16415,N_12071,N_12089);
nor U16416 (N_16416,N_11628,N_13668);
nor U16417 (N_16417,N_12544,N_11125);
and U16418 (N_16418,N_12910,N_10135);
nand U16419 (N_16419,N_12422,N_13472);
and U16420 (N_16420,N_10427,N_12541);
nand U16421 (N_16421,N_10780,N_14651);
and U16422 (N_16422,N_10916,N_14824);
and U16423 (N_16423,N_13596,N_12096);
nand U16424 (N_16424,N_10005,N_13011);
nand U16425 (N_16425,N_12579,N_13567);
nor U16426 (N_16426,N_10154,N_14861);
or U16427 (N_16427,N_14756,N_13834);
nand U16428 (N_16428,N_12861,N_10264);
and U16429 (N_16429,N_12525,N_11873);
nor U16430 (N_16430,N_11335,N_11104);
or U16431 (N_16431,N_10479,N_12596);
nand U16432 (N_16432,N_13964,N_12201);
and U16433 (N_16433,N_12371,N_14727);
or U16434 (N_16434,N_14891,N_14933);
and U16435 (N_16435,N_11396,N_12502);
or U16436 (N_16436,N_11761,N_12956);
or U16437 (N_16437,N_12769,N_11174);
and U16438 (N_16438,N_12813,N_13912);
nor U16439 (N_16439,N_10819,N_12900);
and U16440 (N_16440,N_13221,N_10354);
or U16441 (N_16441,N_13025,N_10178);
nand U16442 (N_16442,N_13741,N_13658);
or U16443 (N_16443,N_10997,N_14844);
or U16444 (N_16444,N_10385,N_12634);
and U16445 (N_16445,N_12992,N_10976);
or U16446 (N_16446,N_12299,N_13174);
nand U16447 (N_16447,N_14975,N_12432);
nand U16448 (N_16448,N_13648,N_10623);
or U16449 (N_16449,N_11657,N_13910);
and U16450 (N_16450,N_12963,N_12894);
and U16451 (N_16451,N_11215,N_11574);
or U16452 (N_16452,N_11586,N_12124);
nand U16453 (N_16453,N_11606,N_12339);
and U16454 (N_16454,N_10174,N_13396);
nor U16455 (N_16455,N_10464,N_13625);
or U16456 (N_16456,N_12060,N_14856);
nor U16457 (N_16457,N_12810,N_11993);
nand U16458 (N_16458,N_14248,N_14160);
and U16459 (N_16459,N_12240,N_11390);
or U16460 (N_16460,N_11653,N_11988);
and U16461 (N_16461,N_11098,N_13103);
and U16462 (N_16462,N_13991,N_11533);
and U16463 (N_16463,N_13681,N_14871);
nor U16464 (N_16464,N_11330,N_10103);
and U16465 (N_16465,N_11286,N_13402);
and U16466 (N_16466,N_11860,N_11851);
or U16467 (N_16467,N_11401,N_14362);
or U16468 (N_16468,N_11106,N_12441);
nor U16469 (N_16469,N_14913,N_14367);
nand U16470 (N_16470,N_11234,N_14496);
nor U16471 (N_16471,N_12699,N_10411);
or U16472 (N_16472,N_10577,N_13968);
xnor U16473 (N_16473,N_10449,N_11562);
nor U16474 (N_16474,N_11739,N_14703);
nand U16475 (N_16475,N_14175,N_11312);
or U16476 (N_16476,N_10750,N_12259);
nand U16477 (N_16477,N_12076,N_12461);
nor U16478 (N_16478,N_13323,N_12945);
nor U16479 (N_16479,N_10715,N_14991);
nor U16480 (N_16480,N_13210,N_14604);
nand U16481 (N_16481,N_10488,N_14584);
or U16482 (N_16482,N_10818,N_10655);
or U16483 (N_16483,N_12187,N_11006);
or U16484 (N_16484,N_10850,N_11291);
or U16485 (N_16485,N_14028,N_13443);
nor U16486 (N_16486,N_14640,N_14205);
and U16487 (N_16487,N_12174,N_12436);
and U16488 (N_16488,N_14698,N_12154);
nand U16489 (N_16489,N_10146,N_12143);
nor U16490 (N_16490,N_14245,N_14314);
or U16491 (N_16491,N_13510,N_13829);
xor U16492 (N_16492,N_13810,N_12740);
nor U16493 (N_16493,N_14036,N_14276);
nand U16494 (N_16494,N_11524,N_14236);
nand U16495 (N_16495,N_12463,N_12227);
or U16496 (N_16496,N_12645,N_13328);
nor U16497 (N_16497,N_14271,N_14889);
nor U16498 (N_16498,N_14808,N_13613);
nor U16499 (N_16499,N_12054,N_12048);
nand U16500 (N_16500,N_13591,N_12008);
nor U16501 (N_16501,N_12226,N_13465);
nor U16502 (N_16502,N_11556,N_14016);
nand U16503 (N_16503,N_12724,N_14538);
and U16504 (N_16504,N_13619,N_14045);
and U16505 (N_16505,N_10669,N_10862);
and U16506 (N_16506,N_10370,N_10983);
or U16507 (N_16507,N_12213,N_12789);
and U16508 (N_16508,N_12957,N_12125);
nor U16509 (N_16509,N_14841,N_13490);
nand U16510 (N_16510,N_11849,N_13072);
and U16511 (N_16511,N_11265,N_10342);
nor U16512 (N_16512,N_10096,N_14715);
or U16513 (N_16513,N_12415,N_11708);
and U16514 (N_16514,N_10010,N_13844);
nand U16515 (N_16515,N_13269,N_14256);
and U16516 (N_16516,N_11045,N_10723);
nand U16517 (N_16517,N_14968,N_14875);
and U16518 (N_16518,N_14798,N_12455);
or U16519 (N_16519,N_12999,N_14796);
nor U16520 (N_16520,N_10859,N_14740);
nand U16521 (N_16521,N_14739,N_13033);
nand U16522 (N_16522,N_11110,N_12254);
nor U16523 (N_16523,N_13008,N_12771);
and U16524 (N_16524,N_14789,N_12000);
or U16525 (N_16525,N_12787,N_12087);
or U16526 (N_16526,N_11346,N_10191);
nor U16527 (N_16527,N_14261,N_14748);
nand U16528 (N_16528,N_14075,N_11243);
nor U16529 (N_16529,N_11781,N_13770);
nand U16530 (N_16530,N_13657,N_11463);
or U16531 (N_16531,N_10122,N_14468);
nor U16532 (N_16532,N_12264,N_14511);
nor U16533 (N_16533,N_11141,N_11544);
or U16534 (N_16534,N_12374,N_14372);
nand U16535 (N_16535,N_12434,N_14733);
or U16536 (N_16536,N_14761,N_14759);
nand U16537 (N_16537,N_13438,N_13038);
or U16538 (N_16538,N_10306,N_11890);
nand U16539 (N_16539,N_14479,N_11823);
or U16540 (N_16540,N_10624,N_11754);
and U16541 (N_16541,N_13205,N_10630);
nor U16542 (N_16542,N_13387,N_13268);
and U16543 (N_16543,N_13094,N_11258);
nand U16544 (N_16544,N_12529,N_14386);
or U16545 (N_16545,N_13715,N_11002);
nor U16546 (N_16546,N_10203,N_10186);
or U16547 (N_16547,N_10461,N_13364);
or U16548 (N_16548,N_12075,N_13836);
or U16549 (N_16549,N_11660,N_10120);
nand U16550 (N_16550,N_10177,N_11665);
nand U16551 (N_16551,N_12874,N_12720);
nor U16552 (N_16552,N_10778,N_11338);
nand U16553 (N_16553,N_13630,N_10529);
and U16554 (N_16554,N_11990,N_10936);
and U16555 (N_16555,N_11319,N_13870);
and U16556 (N_16556,N_10770,N_11317);
nand U16557 (N_16557,N_14318,N_13579);
and U16558 (N_16558,N_13614,N_14843);
and U16559 (N_16559,N_11382,N_13525);
or U16560 (N_16560,N_10517,N_11153);
and U16561 (N_16561,N_12127,N_11693);
nand U16562 (N_16562,N_14289,N_13479);
and U16563 (N_16563,N_11850,N_10374);
or U16564 (N_16564,N_12053,N_14466);
or U16565 (N_16565,N_13307,N_11664);
nand U16566 (N_16566,N_10562,N_12886);
nor U16567 (N_16567,N_11224,N_11318);
xor U16568 (N_16568,N_14902,N_10467);
nand U16569 (N_16569,N_12784,N_13566);
and U16570 (N_16570,N_10713,N_11596);
nand U16571 (N_16571,N_11424,N_14209);
and U16572 (N_16572,N_11717,N_13519);
or U16573 (N_16573,N_10172,N_11027);
nand U16574 (N_16574,N_10985,N_13024);
or U16575 (N_16575,N_12274,N_13966);
and U16576 (N_16576,N_13383,N_11255);
nor U16577 (N_16577,N_12310,N_12778);
or U16578 (N_16578,N_11564,N_14017);
or U16579 (N_16579,N_10653,N_14177);
and U16580 (N_16580,N_10357,N_10521);
nand U16581 (N_16581,N_12179,N_10159);
and U16582 (N_16582,N_11949,N_11630);
and U16583 (N_16583,N_13585,N_14954);
and U16584 (N_16584,N_11499,N_12806);
nor U16585 (N_16585,N_12716,N_14113);
nor U16586 (N_16586,N_13137,N_10865);
and U16587 (N_16587,N_10542,N_14734);
or U16588 (N_16588,N_11083,N_13895);
nand U16589 (N_16589,N_12273,N_13573);
nand U16590 (N_16590,N_10724,N_10716);
nor U16591 (N_16591,N_13202,N_14576);
xor U16592 (N_16592,N_12362,N_11220);
and U16593 (N_16593,N_13533,N_13071);
and U16594 (N_16594,N_14418,N_12987);
nor U16595 (N_16595,N_13485,N_13064);
or U16596 (N_16596,N_13289,N_12700);
and U16597 (N_16597,N_13902,N_14937);
nand U16598 (N_16598,N_12278,N_12108);
nor U16599 (N_16599,N_13262,N_13703);
nor U16600 (N_16600,N_14721,N_13002);
or U16601 (N_16601,N_11600,N_12991);
or U16602 (N_16602,N_12566,N_11353);
or U16603 (N_16603,N_11144,N_11207);
and U16604 (N_16604,N_14059,N_10581);
and U16605 (N_16605,N_11992,N_14894);
xnor U16606 (N_16606,N_12692,N_13909);
and U16607 (N_16607,N_12943,N_11339);
and U16608 (N_16608,N_10358,N_13331);
nor U16609 (N_16609,N_10695,N_13293);
nor U16610 (N_16610,N_13193,N_11641);
or U16611 (N_16611,N_10631,N_11980);
and U16612 (N_16612,N_10087,N_11101);
nor U16613 (N_16613,N_10740,N_10683);
and U16614 (N_16614,N_12835,N_13543);
or U16615 (N_16615,N_12284,N_11404);
or U16616 (N_16616,N_13838,N_14826);
nor U16617 (N_16617,N_14838,N_14755);
and U16618 (N_16618,N_14852,N_13905);
or U16619 (N_16619,N_10226,N_11692);
and U16620 (N_16620,N_14002,N_14444);
nand U16621 (N_16621,N_14679,N_14566);
or U16622 (N_16622,N_11261,N_14482);
or U16623 (N_16623,N_13780,N_14333);
nor U16624 (N_16624,N_12779,N_11616);
nor U16625 (N_16625,N_10485,N_11759);
or U16626 (N_16626,N_13138,N_11427);
or U16627 (N_16627,N_14962,N_13795);
or U16628 (N_16628,N_14483,N_12444);
or U16629 (N_16629,N_14385,N_13457);
or U16630 (N_16630,N_13347,N_14539);
nand U16631 (N_16631,N_11737,N_10569);
nand U16632 (N_16632,N_10965,N_10379);
nor U16633 (N_16633,N_12928,N_14231);
or U16634 (N_16634,N_12051,N_13224);
and U16635 (N_16635,N_11066,N_11190);
and U16636 (N_16636,N_13722,N_10276);
nand U16637 (N_16637,N_10763,N_13334);
nand U16638 (N_16638,N_13363,N_13320);
nand U16639 (N_16639,N_11171,N_11633);
and U16640 (N_16640,N_11514,N_13529);
and U16641 (N_16641,N_12479,N_12980);
nor U16642 (N_16642,N_11223,N_14883);
and U16643 (N_16643,N_10795,N_12134);
nor U16644 (N_16644,N_14923,N_14746);
or U16645 (N_16645,N_12507,N_10473);
xnor U16646 (N_16646,N_12122,N_14820);
or U16647 (N_16647,N_13390,N_12836);
and U16648 (N_16648,N_10015,N_13166);
nor U16649 (N_16649,N_10791,N_13261);
and U16650 (N_16650,N_14213,N_13581);
and U16651 (N_16651,N_11056,N_11858);
or U16652 (N_16652,N_11451,N_11651);
or U16653 (N_16653,N_12464,N_10515);
nor U16654 (N_16654,N_12983,N_12657);
or U16655 (N_16655,N_10792,N_12977);
and U16656 (N_16656,N_12748,N_14286);
and U16657 (N_16657,N_12376,N_12430);
or U16658 (N_16658,N_10032,N_13316);
and U16659 (N_16659,N_12514,N_14792);
nor U16660 (N_16660,N_12493,N_10502);
and U16661 (N_16661,N_12719,N_14204);
nor U16662 (N_16662,N_10441,N_14870);
and U16663 (N_16663,N_12309,N_14700);
nor U16664 (N_16664,N_14783,N_12552);
and U16665 (N_16665,N_13115,N_14802);
and U16666 (N_16666,N_14430,N_12466);
or U16667 (N_16667,N_13764,N_13464);
and U16668 (N_16668,N_10200,N_11500);
nor U16669 (N_16669,N_13932,N_13372);
or U16670 (N_16670,N_12594,N_14443);
nor U16671 (N_16671,N_14622,N_11187);
and U16672 (N_16672,N_14505,N_13029);
nor U16673 (N_16673,N_14199,N_10753);
nand U16674 (N_16674,N_12995,N_10528);
or U16675 (N_16675,N_10592,N_10815);
nand U16676 (N_16676,N_10417,N_14568);
nor U16677 (N_16677,N_11372,N_11370);
nand U16678 (N_16678,N_13199,N_13546);
nor U16679 (N_16679,N_14949,N_13717);
and U16680 (N_16680,N_10710,N_14518);
and U16681 (N_16681,N_10772,N_11035);
nand U16682 (N_16682,N_12346,N_11038);
and U16683 (N_16683,N_10535,N_13426);
nor U16684 (N_16684,N_14390,N_11943);
nor U16685 (N_16685,N_11672,N_10664);
nor U16686 (N_16686,N_11892,N_10576);
or U16687 (N_16687,N_10830,N_13762);
and U16688 (N_16688,N_12202,N_12064);
nand U16689 (N_16689,N_14463,N_13225);
or U16690 (N_16690,N_13923,N_12499);
and U16691 (N_16691,N_11655,N_14150);
nand U16692 (N_16692,N_11868,N_12155);
and U16693 (N_16693,N_13601,N_11975);
or U16694 (N_16694,N_10737,N_12545);
or U16695 (N_16695,N_12281,N_13849);
nand U16696 (N_16696,N_14678,N_14560);
nor U16697 (N_16697,N_12950,N_13274);
nand U16698 (N_16698,N_14269,N_14881);
or U16699 (N_16699,N_10425,N_14240);
nand U16700 (N_16700,N_14979,N_14005);
and U16701 (N_16701,N_12770,N_14925);
or U16702 (N_16702,N_11663,N_12260);
and U16703 (N_16703,N_12612,N_11690);
and U16704 (N_16704,N_12788,N_12325);
or U16705 (N_16705,N_11510,N_14384);
nand U16706 (N_16706,N_14445,N_12785);
nand U16707 (N_16707,N_10993,N_12327);
nor U16708 (N_16708,N_11790,N_11048);
nand U16709 (N_16709,N_14249,N_12715);
nand U16710 (N_16710,N_14313,N_10294);
nand U16711 (N_16711,N_14403,N_10597);
and U16712 (N_16712,N_13352,N_11497);
nand U16713 (N_16713,N_14145,N_12844);
nor U16714 (N_16714,N_11324,N_11836);
and U16715 (N_16715,N_14321,N_10382);
or U16716 (N_16716,N_13043,N_13965);
or U16717 (N_16717,N_14094,N_12707);
and U16718 (N_16718,N_12222,N_14247);
nand U16719 (N_16719,N_14020,N_10183);
nand U16720 (N_16720,N_10462,N_13759);
or U16721 (N_16721,N_12804,N_13073);
and U16722 (N_16722,N_12852,N_12654);
and U16723 (N_16723,N_14793,N_14440);
nor U16724 (N_16724,N_11230,N_13754);
nand U16725 (N_16725,N_10758,N_10787);
or U16726 (N_16726,N_11955,N_12166);
and U16727 (N_16727,N_13360,N_10101);
or U16728 (N_16728,N_11521,N_11503);
nor U16729 (N_16729,N_14513,N_10969);
and U16730 (N_16730,N_13332,N_14221);
or U16731 (N_16731,N_10896,N_11399);
nor U16732 (N_16732,N_13454,N_14290);
or U16733 (N_16733,N_11847,N_11309);
nand U16734 (N_16734,N_13990,N_12249);
or U16735 (N_16735,N_12689,N_13926);
nand U16736 (N_16736,N_14190,N_13852);
and U16737 (N_16737,N_10130,N_11030);
and U16738 (N_16738,N_12532,N_12118);
and U16739 (N_16739,N_14396,N_13636);
nor U16740 (N_16740,N_14602,N_10397);
and U16741 (N_16741,N_13704,N_12354);
and U16742 (N_16742,N_13868,N_11377);
and U16743 (N_16743,N_11068,N_13882);
nor U16744 (N_16744,N_11733,N_13814);
and U16745 (N_16745,N_11516,N_11659);
nand U16746 (N_16746,N_14351,N_11124);
nor U16747 (N_16747,N_12317,N_10886);
nor U16748 (N_16748,N_14346,N_14162);
nor U16749 (N_16749,N_10939,N_14971);
nand U16750 (N_16750,N_10489,N_10020);
or U16751 (N_16751,N_12912,N_14695);
nand U16752 (N_16752,N_12567,N_11643);
or U16753 (N_16753,N_10117,N_11741);
and U16754 (N_16754,N_11155,N_14228);
or U16755 (N_16755,N_14297,N_12280);
nand U16756 (N_16756,N_14777,N_11082);
nand U16757 (N_16757,N_10347,N_14836);
or U16758 (N_16758,N_12321,N_14188);
nand U16759 (N_16759,N_12091,N_12136);
nor U16760 (N_16760,N_13492,N_12392);
and U16761 (N_16761,N_11331,N_12767);
and U16762 (N_16762,N_11999,N_12978);
nand U16763 (N_16763,N_11441,N_12486);
and U16764 (N_16764,N_10167,N_13129);
or U16765 (N_16765,N_12146,N_13474);
or U16766 (N_16766,N_10311,N_11976);
nor U16767 (N_16767,N_11774,N_12800);
or U16768 (N_16768,N_10800,N_12061);
nor U16769 (N_16769,N_14310,N_12997);
or U16770 (N_16770,N_14718,N_12447);
and U16771 (N_16771,N_13520,N_10084);
xor U16772 (N_16772,N_10890,N_14829);
nor U16773 (N_16773,N_10745,N_14728);
or U16774 (N_16774,N_10744,N_12774);
nor U16775 (N_16775,N_10305,N_14358);
nand U16776 (N_16776,N_13175,N_14998);
nand U16777 (N_16777,N_12583,N_10434);
nand U16778 (N_16778,N_14804,N_13450);
and U16779 (N_16779,N_14724,N_13427);
nand U16780 (N_16780,N_10748,N_11957);
and U16781 (N_16781,N_13811,N_10524);
nand U16782 (N_16782,N_13623,N_10021);
and U16783 (N_16783,N_13411,N_11046);
or U16784 (N_16784,N_10269,N_10739);
nor U16785 (N_16785,N_11777,N_10616);
and U16786 (N_16786,N_10731,N_13106);
nor U16787 (N_16787,N_13835,N_12938);
nand U16788 (N_16788,N_11290,N_13504);
or U16789 (N_16789,N_10593,N_11848);
nand U16790 (N_16790,N_12028,N_14664);
xor U16791 (N_16791,N_13178,N_12404);
and U16792 (N_16792,N_12236,N_12343);
or U16793 (N_16793,N_10973,N_12367);
nor U16794 (N_16794,N_14986,N_10201);
and U16795 (N_16795,N_14341,N_13784);
and U16796 (N_16796,N_10932,N_13767);
and U16797 (N_16797,N_11529,N_12341);
xnor U16798 (N_16798,N_10611,N_10225);
nor U16799 (N_16799,N_14557,N_14839);
and U16800 (N_16800,N_13398,N_13244);
nand U16801 (N_16801,N_10947,N_13369);
nor U16802 (N_16802,N_14179,N_14880);
xnor U16803 (N_16803,N_13982,N_14911);
or U16804 (N_16804,N_11620,N_14985);
nand U16805 (N_16805,N_14135,N_11558);
nand U16806 (N_16806,N_10181,N_14582);
and U16807 (N_16807,N_13381,N_14810);
nand U16808 (N_16808,N_12893,N_14353);
and U16809 (N_16809,N_11072,N_12402);
nand U16810 (N_16810,N_14812,N_10129);
nand U16811 (N_16811,N_10761,N_12157);
nor U16812 (N_16812,N_12561,N_11333);
and U16813 (N_16813,N_12406,N_13361);
and U16814 (N_16814,N_12442,N_12682);
nor U16815 (N_16815,N_12148,N_13301);
and U16816 (N_16816,N_14776,N_10538);
or U16817 (N_16817,N_14840,N_12878);
or U16818 (N_16818,N_10942,N_11322);
nor U16819 (N_16819,N_12263,N_10108);
or U16820 (N_16820,N_13977,N_13830);
and U16821 (N_16821,N_11626,N_10940);
or U16822 (N_16822,N_11204,N_12443);
nor U16823 (N_16823,N_12754,N_11856);
nand U16824 (N_16824,N_13083,N_10814);
nand U16825 (N_16825,N_12580,N_10244);
nand U16826 (N_16826,N_10413,N_12056);
and U16827 (N_16827,N_11832,N_14426);
nor U16828 (N_16828,N_13486,N_12102);
nor U16829 (N_16829,N_11483,N_12969);
or U16830 (N_16830,N_11240,N_12010);
or U16831 (N_16831,N_12178,N_11321);
or U16832 (N_16832,N_10742,N_14328);
nor U16833 (N_16833,N_14586,N_11528);
or U16834 (N_16834,N_10022,N_14765);
or U16835 (N_16835,N_13201,N_11121);
nand U16836 (N_16836,N_13295,N_13415);
and U16837 (N_16837,N_14714,N_14931);
nor U16838 (N_16838,N_10662,N_12622);
and U16839 (N_16839,N_13571,N_10738);
nor U16840 (N_16840,N_10531,N_10974);
nor U16841 (N_16841,N_13113,N_12776);
nand U16842 (N_16842,N_14273,N_10296);
and U16843 (N_16843,N_13627,N_12592);
nor U16844 (N_16844,N_13039,N_14916);
and U16845 (N_16845,N_13001,N_12934);
nand U16846 (N_16846,N_14130,N_13357);
nand U16847 (N_16847,N_13635,N_13804);
and U16848 (N_16848,N_11579,N_14183);
nor U16849 (N_16849,N_10176,N_14876);
or U16850 (N_16850,N_10603,N_12019);
or U16851 (N_16851,N_12600,N_11031);
xor U16852 (N_16852,N_14716,N_10386);
nand U16853 (N_16853,N_13933,N_10011);
or U16854 (N_16854,N_12435,N_14554);
and U16855 (N_16855,N_10057,N_10465);
and U16856 (N_16856,N_13042,N_14630);
or U16857 (N_16857,N_10196,N_14391);
or U16858 (N_16858,N_14424,N_13462);
or U16859 (N_16859,N_12041,N_12569);
and U16860 (N_16860,N_12225,N_13056);
nor U16861 (N_16861,N_11994,N_11269);
or U16862 (N_16862,N_13807,N_11278);
and U16863 (N_16863,N_12918,N_13530);
or U16864 (N_16864,N_10534,N_12068);
xnor U16865 (N_16865,N_13126,N_14476);
nor U16866 (N_16866,N_10175,N_10378);
and U16867 (N_16867,N_14528,N_13871);
or U16868 (N_16868,N_10855,N_11629);
nand U16869 (N_16869,N_10053,N_14530);
nand U16870 (N_16870,N_12277,N_11902);
and U16871 (N_16871,N_11896,N_11580);
or U16872 (N_16872,N_14497,N_11475);
nand U16873 (N_16873,N_11420,N_10635);
or U16874 (N_16874,N_10852,N_12530);
and U16875 (N_16875,N_10477,N_12485);
nand U16876 (N_16876,N_14230,N_10341);
or U16877 (N_16877,N_13919,N_14344);
nand U16878 (N_16878,N_10285,N_13711);
and U16879 (N_16879,N_12424,N_12172);
and U16880 (N_16880,N_12638,N_11611);
and U16881 (N_16881,N_11671,N_11264);
nor U16882 (N_16882,N_14627,N_13706);
and U16883 (N_16883,N_10495,N_11934);
or U16884 (N_16884,N_12469,N_10006);
nand U16885 (N_16885,N_10979,N_13782);
nor U16886 (N_16886,N_10627,N_13227);
nor U16887 (N_16887,N_13911,N_14340);
nor U16888 (N_16888,N_12662,N_11203);
or U16889 (N_16889,N_12811,N_13495);
nand U16890 (N_16890,N_11793,N_11654);
or U16891 (N_16891,N_12686,N_12405);
nand U16892 (N_16892,N_10512,N_12029);
or U16893 (N_16893,N_10110,N_12006);
nand U16894 (N_16894,N_13280,N_11431);
nor U16895 (N_16895,N_12964,N_11417);
or U16896 (N_16896,N_14337,N_14848);
or U16897 (N_16897,N_13228,N_10279);
or U16898 (N_16898,N_13620,N_13358);
or U16899 (N_16899,N_10856,N_13181);
or U16900 (N_16900,N_10956,N_11059);
and U16901 (N_16901,N_12267,N_11323);
nor U16902 (N_16902,N_12812,N_11647);
nand U16903 (N_16903,N_10023,N_10697);
nand U16904 (N_16904,N_12751,N_13251);
and U16905 (N_16905,N_12197,N_11478);
and U16906 (N_16906,N_13074,N_11096);
or U16907 (N_16907,N_10231,N_10672);
and U16908 (N_16908,N_13182,N_11732);
or U16909 (N_16909,N_10229,N_10412);
nor U16910 (N_16910,N_11872,N_12111);
nand U16911 (N_16911,N_11923,N_11075);
nand U16912 (N_16912,N_11658,N_14307);
or U16913 (N_16913,N_11078,N_10694);
and U16914 (N_16914,N_12465,N_10601);
and U16915 (N_16915,N_14015,N_11383);
nand U16916 (N_16916,N_14187,N_11021);
and U16917 (N_16917,N_13422,N_14041);
or U16918 (N_16918,N_11425,N_13144);
or U16919 (N_16919,N_14262,N_12624);
and U16920 (N_16920,N_11320,N_11437);
nand U16921 (N_16921,N_10899,N_12590);
and U16922 (N_16922,N_10309,N_11409);
and U16923 (N_16923,N_13979,N_12867);
nand U16924 (N_16924,N_12959,N_14967);
nand U16925 (N_16925,N_11288,N_13183);
nor U16926 (N_16926,N_13592,N_10355);
nor U16927 (N_16927,N_12428,N_10323);
nor U16928 (N_16928,N_10989,N_10832);
or U16929 (N_16929,N_12438,N_11557);
nand U16930 (N_16930,N_11150,N_12315);
or U16931 (N_16931,N_13503,N_10238);
nor U16932 (N_16932,N_13674,N_11517);
nand U16933 (N_16933,N_12623,N_11911);
or U16934 (N_16934,N_13843,N_14672);
and U16935 (N_16935,N_14263,N_11276);
or U16936 (N_16936,N_14168,N_13921);
nand U16937 (N_16937,N_12575,N_11932);
nor U16938 (N_16938,N_10076,N_11688);
or U16939 (N_16939,N_14522,N_10511);
nor U16940 (N_16940,N_11569,N_13678);
or U16941 (N_16941,N_11731,N_14068);
or U16942 (N_16942,N_12618,N_10570);
nor U16943 (N_16943,N_13257,N_10071);
or U16944 (N_16944,N_12184,N_12011);
nand U16945 (N_16945,N_11719,N_11117);
and U16946 (N_16946,N_10131,N_13211);
nand U16947 (N_16947,N_10494,N_11109);
or U16948 (N_16948,N_11893,N_13640);
nand U16949 (N_16949,N_11053,N_10065);
nand U16950 (N_16950,N_12604,N_12611);
nand U16951 (N_16951,N_11361,N_11808);
nor U16952 (N_16952,N_14104,N_10829);
and U16953 (N_16953,N_13171,N_12807);
nand U16954 (N_16954,N_13738,N_14124);
nor U16955 (N_16955,N_14851,N_11426);
or U16956 (N_16956,N_12509,N_11826);
or U16957 (N_16957,N_10295,N_14551);
nor U16958 (N_16958,N_12471,N_10456);
nand U16959 (N_16959,N_13424,N_13918);
and U16960 (N_16960,N_11769,N_12168);
and U16961 (N_16961,N_12548,N_11213);
nand U16962 (N_16962,N_11984,N_14355);
nor U16963 (N_16963,N_14784,N_10853);
nand U16964 (N_16964,N_14594,N_14830);
xnor U16965 (N_16965,N_12609,N_11074);
or U16966 (N_16966,N_11568,N_14401);
or U16967 (N_16967,N_14226,N_14821);
or U16968 (N_16968,N_13725,N_10304);
nand U16969 (N_16969,N_13575,N_10915);
or U16970 (N_16970,N_10291,N_12616);
or U16971 (N_16971,N_10034,N_11384);
nand U16972 (N_16972,N_14185,N_13026);
nand U16973 (N_16973,N_13036,N_12772);
nand U16974 (N_16974,N_14899,N_14906);
nor U16975 (N_16975,N_12792,N_13000);
nand U16976 (N_16976,N_12470,N_10533);
nor U16977 (N_16977,N_14264,N_14615);
xor U16978 (N_16978,N_10927,N_12478);
nor U16979 (N_16979,N_13994,N_14196);
nand U16980 (N_16980,N_11601,N_11915);
nor U16981 (N_16981,N_14948,N_13855);
and U16982 (N_16982,N_10594,N_13168);
nor U16983 (N_16983,N_11398,N_12551);
nor U16984 (N_16984,N_12239,N_13928);
nand U16985 (N_16985,N_10199,N_12307);
or U16986 (N_16986,N_14537,N_10095);
nor U16987 (N_16987,N_13089,N_10579);
or U16988 (N_16988,N_14688,N_12257);
nor U16989 (N_16989,N_11842,N_14668);
nand U16990 (N_16990,N_14909,N_11227);
or U16991 (N_16991,N_13500,N_10399);
and U16992 (N_16992,N_10408,N_10617);
nand U16993 (N_16993,N_11531,N_10336);
or U16994 (N_16994,N_11905,N_13813);
or U16995 (N_16995,N_14026,N_11042);
nor U16996 (N_16996,N_13478,N_14754);
or U16997 (N_16997,N_12262,N_10169);
or U16998 (N_16998,N_10026,N_12013);
and U16999 (N_16999,N_10501,N_12352);
nor U17000 (N_17000,N_11245,N_10455);
or U17001 (N_17001,N_10513,N_14103);
nor U17002 (N_17002,N_10858,N_11838);
nand U17003 (N_17003,N_13401,N_12296);
nor U17004 (N_17004,N_13761,N_14420);
nand U17005 (N_17005,N_14121,N_13258);
nor U17006 (N_17006,N_10962,N_14524);
or U17007 (N_17007,N_14790,N_11216);
nor U17008 (N_17008,N_12322,N_14635);
and U17009 (N_17009,N_12038,N_12896);
or U17010 (N_17010,N_11987,N_12749);
nor U17011 (N_17011,N_14438,N_11328);
or U17012 (N_17012,N_11961,N_10762);
and U17013 (N_17013,N_13218,N_13489);
nand U17014 (N_17014,N_12364,N_13649);
nand U17015 (N_17015,N_10848,N_14359);
nand U17016 (N_17016,N_10777,N_11363);
and U17017 (N_17017,N_13916,N_10105);
or U17018 (N_17018,N_14432,N_14267);
nor U17019 (N_17019,N_12200,N_14893);
nand U17020 (N_17020,N_10659,N_11874);
nand U17021 (N_17021,N_11184,N_10333);
and U17022 (N_17022,N_13125,N_12725);
and U17023 (N_17023,N_10882,N_14207);
and U17024 (N_17024,N_13404,N_13229);
and U17025 (N_17025,N_12750,N_11813);
xnor U17026 (N_17026,N_13587,N_12919);
and U17027 (N_17027,N_11094,N_10736);
and U17028 (N_17028,N_13291,N_12045);
nor U17029 (N_17029,N_13394,N_12205);
nor U17030 (N_17030,N_11256,N_11795);
xnor U17031 (N_17031,N_10690,N_12228);
nor U17032 (N_17032,N_13938,N_10817);
or U17033 (N_17033,N_12909,N_11694);
or U17034 (N_17034,N_13695,N_11560);
xor U17035 (N_17035,N_14895,N_10008);
and U17036 (N_17036,N_10258,N_12086);
or U17037 (N_17037,N_12395,N_11176);
nand U17038 (N_17038,N_11783,N_10078);
nor U17039 (N_17039,N_14493,N_14847);
and U17040 (N_17040,N_13220,N_10270);
nand U17041 (N_17041,N_14606,N_10807);
or U17042 (N_17042,N_12833,N_10457);
nand U17043 (N_17043,N_12500,N_10289);
and U17044 (N_17044,N_10250,N_10559);
nand U17045 (N_17045,N_11047,N_14689);
or U17046 (N_17046,N_12308,N_12199);
and U17047 (N_17047,N_12083,N_11385);
or U17048 (N_17048,N_10371,N_13665);
or U17049 (N_17049,N_14837,N_14018);
nand U17050 (N_17050,N_11773,N_10029);
nor U17051 (N_17051,N_11583,N_14319);
and U17052 (N_17052,N_11026,N_14779);
nor U17053 (N_17053,N_14704,N_10407);
and U17054 (N_17054,N_12065,N_10102);
nor U17055 (N_17055,N_13839,N_14452);
or U17056 (N_17056,N_10995,N_11880);
nand U17057 (N_17057,N_11909,N_11545);
or U17058 (N_17058,N_12329,N_10429);
nand U17059 (N_17059,N_11970,N_13976);
or U17060 (N_17060,N_12380,N_11172);
nor U17061 (N_17061,N_12676,N_14472);
nand U17062 (N_17062,N_13907,N_14543);
and U17063 (N_17063,N_14069,N_12212);
and U17064 (N_17064,N_10151,N_12908);
and U17065 (N_17065,N_11371,N_12290);
and U17066 (N_17066,N_13673,N_11271);
nand U17067 (N_17067,N_14347,N_13327);
and U17068 (N_17068,N_11191,N_14833);
nand U17069 (N_17069,N_10463,N_14487);
nand U17070 (N_17070,N_14098,N_12055);
and U17071 (N_17071,N_14412,N_13487);
and U17072 (N_17072,N_13812,N_13532);
or U17073 (N_17073,N_10721,N_11126);
and U17074 (N_17074,N_14304,N_14665);
nand U17075 (N_17075,N_12732,N_12901);
nand U17076 (N_17076,N_12895,N_12520);
nand U17077 (N_17077,N_10016,N_13605);
nor U17078 (N_17078,N_11960,N_13729);
nor U17079 (N_17079,N_14978,N_11008);
and U17080 (N_17080,N_11173,N_11413);
or U17081 (N_17081,N_10075,N_10326);
nor U17082 (N_17082,N_13018,N_14133);
nor U17083 (N_17083,N_12397,N_10266);
nand U17084 (N_17084,N_11691,N_10779);
nor U17085 (N_17085,N_10854,N_12413);
xor U17086 (N_17086,N_13140,N_14671);
and U17087 (N_17087,N_14816,N_12932);
nand U17088 (N_17088,N_11840,N_13287);
and U17089 (N_17089,N_12324,N_12653);
nor U17090 (N_17090,N_12524,N_11118);
and U17091 (N_17091,N_14532,N_14089);
or U17092 (N_17092,N_11792,N_12953);
or U17093 (N_17093,N_13562,N_13139);
nor U17094 (N_17094,N_12379,N_12924);
or U17095 (N_17095,N_14106,N_12650);
nor U17096 (N_17096,N_12119,N_12781);
nor U17097 (N_17097,N_14110,N_12004);
or U17098 (N_17098,N_13808,N_11196);
nor U17099 (N_17099,N_11054,N_10732);
nor U17100 (N_17100,N_13317,N_14375);
or U17101 (N_17101,N_13609,N_14667);
nor U17102 (N_17102,N_12121,N_12951);
nor U17103 (N_17103,N_11728,N_10934);
and U17104 (N_17104,N_12472,N_12116);
nand U17105 (N_17105,N_13122,N_10081);
or U17106 (N_17106,N_14907,N_13084);
and U17107 (N_17107,N_13570,N_12295);
and U17108 (N_17108,N_14770,N_11592);
nor U17109 (N_17109,N_13731,N_12066);
nand U17110 (N_17110,N_13081,N_11472);
xor U17111 (N_17111,N_12037,N_13527);
or U17112 (N_17112,N_14126,N_13854);
and U17113 (N_17113,N_14953,N_13466);
and U17114 (N_17114,N_14772,N_13637);
and U17115 (N_17115,N_13758,N_11392);
nand U17116 (N_17116,N_14892,N_11140);
nand U17117 (N_17117,N_14929,N_12868);
or U17118 (N_17118,N_13444,N_13559);
and U17119 (N_17119,N_11746,N_10526);
nor U17120 (N_17120,N_14572,N_13068);
nor U17121 (N_17121,N_14032,N_12079);
or U17122 (N_17122,N_12153,N_13511);
or U17123 (N_17123,N_12237,N_10050);
and U17124 (N_17124,N_14570,N_11782);
nor U17125 (N_17125,N_10898,N_11325);
nand U17126 (N_17126,N_10405,N_13190);
nand U17127 (N_17127,N_10565,N_12930);
nand U17128 (N_17128,N_10970,N_14246);
and U17129 (N_17129,N_11465,N_14460);
and U17130 (N_17130,N_14462,N_12589);
nor U17131 (N_17131,N_12906,N_14099);
and U17132 (N_17132,N_10877,N_10704);
or U17133 (N_17133,N_12914,N_10069);
nor U17134 (N_17134,N_10060,N_11049);
nor U17135 (N_17135,N_11080,N_10647);
nand U17136 (N_17136,N_10207,N_12231);
nor U17137 (N_17137,N_10887,N_14164);
nand U17138 (N_17138,N_11898,N_12219);
and U17139 (N_17139,N_12169,N_13410);
or U17140 (N_17140,N_11128,N_13045);
nand U17141 (N_17141,N_14082,N_13647);
or U17142 (N_17142,N_12311,N_11684);
or U17143 (N_17143,N_11336,N_13048);
and U17144 (N_17144,N_14877,N_14499);
and U17145 (N_17145,N_11177,N_14470);
or U17146 (N_17146,N_11539,N_10307);
nand U17147 (N_17147,N_13348,N_13561);
nor U17148 (N_17148,N_12826,N_13679);
and U17149 (N_17149,N_10555,N_11578);
nor U17150 (N_17150,N_14600,N_11484);
or U17151 (N_17151,N_11788,N_13104);
xnor U17152 (N_17152,N_10946,N_13021);
nand U17153 (N_17153,N_13239,N_12229);
and U17154 (N_17154,N_11486,N_14575);
and U17155 (N_17155,N_11015,N_10599);
or U17156 (N_17156,N_10849,N_11029);
and U17157 (N_17157,N_13958,N_10431);
or U17158 (N_17158,N_10654,N_12072);
or U17159 (N_17159,N_11303,N_10109);
nor U17160 (N_17160,N_13978,N_11712);
nor U17161 (N_17161,N_14242,N_13803);
and U17162 (N_17162,N_10884,N_13536);
and U17163 (N_17163,N_13329,N_10242);
nand U17164 (N_17164,N_13883,N_14988);
and U17165 (N_17165,N_11494,N_14764);
and U17166 (N_17166,N_12494,N_13708);
nand U17167 (N_17167,N_14730,N_11095);
nor U17168 (N_17168,N_14762,N_10288);
nand U17169 (N_17169,N_10504,N_13549);
nand U17170 (N_17170,N_11489,N_14243);
nor U17171 (N_17171,N_12081,N_11785);
and U17172 (N_17172,N_13207,N_10657);
and U17173 (N_17173,N_14170,N_14785);
nand U17174 (N_17174,N_13734,N_12476);
or U17175 (N_17175,N_10566,N_13215);
nand U17176 (N_17176,N_13509,N_11146);
and U17177 (N_17177,N_14365,N_13737);
nor U17178 (N_17178,N_13548,N_12316);
and U17179 (N_17179,N_13766,N_10134);
nor U17180 (N_17180,N_10314,N_10904);
or U17181 (N_17181,N_14378,N_14915);
nor U17182 (N_17182,N_10682,N_11825);
and U17183 (N_17183,N_10999,N_10112);
nor U17184 (N_17184,N_11982,N_10607);
nor U17185 (N_17185,N_11226,N_11468);
nand U17186 (N_17186,N_11019,N_12652);
and U17187 (N_17187,N_10031,N_13742);
nor U17188 (N_17188,N_13335,N_14781);
or U17189 (N_17189,N_12911,N_10447);
or U17190 (N_17190,N_12353,N_14960);
or U17191 (N_17191,N_13133,N_10469);
nand U17192 (N_17192,N_12834,N_10688);
or U17193 (N_17193,N_12372,N_12637);
nand U17194 (N_17194,N_12876,N_10375);
nor U17195 (N_17195,N_13538,N_10871);
and U17196 (N_17196,N_11551,N_12848);
nor U17197 (N_17197,N_13458,N_11751);
nand U17198 (N_17198,N_13847,N_11855);
nor U17199 (N_17199,N_13250,N_10519);
and U17200 (N_17200,N_14855,N_11907);
nor U17201 (N_17201,N_11554,N_12553);
nor U17202 (N_17202,N_10260,N_12298);
and U17203 (N_17203,N_13773,N_11637);
or U17204 (N_17204,N_10392,N_14371);
or U17205 (N_17205,N_10701,N_13493);
nand U17206 (N_17206,N_14208,N_13119);
or U17207 (N_17207,N_14219,N_10252);
or U17208 (N_17208,N_12300,N_12981);
or U17209 (N_17209,N_10373,N_13066);
and U17210 (N_17210,N_11937,N_13541);
and U17211 (N_17211,N_11378,N_14356);
and U17212 (N_17212,N_10868,N_13653);
nand U17213 (N_17213,N_12865,N_12730);
nor U17214 (N_17214,N_10539,N_12668);
nand U17215 (N_17215,N_12099,N_11768);
nand U17216 (N_17216,N_13775,N_10600);
nand U17217 (N_17217,N_11193,N_12167);
and U17218 (N_17218,N_10433,N_10734);
nor U17219 (N_17219,N_10505,N_13150);
or U17220 (N_17220,N_13975,N_13983);
xor U17221 (N_17221,N_13823,N_13611);
nor U17222 (N_17222,N_13127,N_10255);
and U17223 (N_17223,N_12128,N_11740);
nand U17224 (N_17224,N_12889,N_11767);
nand U17225 (N_17225,N_11089,N_10253);
nor U17226 (N_17226,N_13238,N_13078);
and U17227 (N_17227,N_10356,N_14690);
nand U17228 (N_17228,N_14567,N_14944);
nor U17229 (N_17229,N_14660,N_13434);
or U17230 (N_17230,N_10806,N_12538);
and U17231 (N_17231,N_14882,N_12113);
or U17232 (N_17232,N_10549,N_10054);
nand U17233 (N_17233,N_10746,N_14556);
nand U17234 (N_17234,N_10873,N_11138);
nand U17235 (N_17235,N_13963,N_14013);
nor U17236 (N_17236,N_13118,N_13896);
and U17237 (N_17237,N_10757,N_11938);
nor U17238 (N_17238,N_10585,N_11895);
nor U17239 (N_17239,N_12815,N_14686);
nand U17240 (N_17240,N_12446,N_12887);
or U17241 (N_17241,N_14927,N_10228);
or U17242 (N_17242,N_10453,N_12162);
and U17243 (N_17243,N_12543,N_11077);
nand U17244 (N_17244,N_12533,N_13756);
and U17245 (N_17245,N_11183,N_14527);
or U17246 (N_17246,N_10157,N_14474);
and U17247 (N_17247,N_10957,N_12534);
and U17248 (N_17248,N_12488,N_14298);
or U17249 (N_17249,N_12559,N_10292);
nor U17250 (N_17250,N_12814,N_10663);
and U17251 (N_17251,N_14874,N_14065);
and U17252 (N_17252,N_12554,N_13416);
or U17253 (N_17253,N_13437,N_11876);
nor U17254 (N_17254,N_10971,N_12746);
nand U17255 (N_17255,N_12210,N_11677);
nand U17256 (N_17256,N_10284,N_13553);
xnor U17257 (N_17257,N_10892,N_12764);
nand U17258 (N_17258,N_11159,N_13655);
or U17259 (N_17259,N_11028,N_11097);
nand U17260 (N_17260,N_14127,N_12429);
nor U17261 (N_17261,N_11523,N_10448);
nand U17262 (N_17262,N_12577,N_10541);
nand U17263 (N_17263,N_14405,N_12080);
nand U17264 (N_17264,N_14987,N_11948);
and U17265 (N_17265,N_10843,N_12506);
or U17266 (N_17266,N_11036,N_13943);
nand U17267 (N_17267,N_14451,N_10972);
or U17268 (N_17268,N_14495,N_13781);
nand U17269 (N_17269,N_12285,N_10245);
or U17270 (N_17270,N_13267,N_10099);
or U17271 (N_17271,N_12877,N_13461);
and U17272 (N_17272,N_12180,N_11749);
and U17273 (N_17273,N_13476,N_12313);
nand U17274 (N_17274,N_12535,N_14558);
and U17275 (N_17275,N_12854,N_12990);
and U17276 (N_17276,N_10938,N_12238);
or U17277 (N_17277,N_14888,N_13917);
nor U17278 (N_17278,N_10894,N_14573);
nand U17279 (N_17279,N_14519,N_13863);
nand U17280 (N_17280,N_13718,N_13365);
or U17281 (N_17281,N_12673,N_14738);
nor U17282 (N_17282,N_12451,N_14940);
or U17283 (N_17283,N_10121,N_14835);
or U17284 (N_17284,N_11050,N_14092);
nor U17285 (N_17285,N_13330,N_10235);
and U17286 (N_17286,N_12967,N_12067);
and U17287 (N_17287,N_12599,N_10718);
nand U17288 (N_17288,N_10805,N_11757);
nor U17289 (N_17289,N_13685,N_13340);
nand U17290 (N_17290,N_14515,N_13915);
and U17291 (N_17291,N_11724,N_10158);
or U17292 (N_17292,N_11351,N_14814);
and U17293 (N_17293,N_14637,N_12801);
nor U17294 (N_17294,N_14415,N_13952);
nor U17295 (N_17295,N_11405,N_12948);
nand U17296 (N_17296,N_14683,N_14928);
nor U17297 (N_17297,N_12639,N_13831);
and U17298 (N_17298,N_13271,N_14311);
and U17299 (N_17299,N_14078,N_11871);
nor U17300 (N_17300,N_11356,N_12973);
or U17301 (N_17301,N_10451,N_11131);
or U17302 (N_17302,N_11541,N_12860);
nor U17303 (N_17303,N_14277,N_11197);
and U17304 (N_17304,N_13040,N_13872);
nor U17305 (N_17305,N_13403,N_12864);
nand U17306 (N_17306,N_13312,N_11219);
or U17307 (N_17307,N_12241,N_11927);
or U17308 (N_17308,N_11634,N_10114);
or U17309 (N_17309,N_14154,N_12193);
and U17310 (N_17310,N_14108,N_13772);
and U17311 (N_17311,N_13598,N_13114);
nor U17312 (N_17312,N_10699,N_10751);
nand U17313 (N_17313,N_14818,N_12677);
or U17314 (N_17314,N_11953,N_12703);
nor U17315 (N_17315,N_14266,N_10262);
nand U17316 (N_17316,N_14257,N_13337);
and U17317 (N_17317,N_10727,N_13997);
nand U17318 (N_17318,N_13660,N_13702);
or U17319 (N_17319,N_10935,N_14296);
and U17320 (N_17320,N_13748,N_13086);
and U17321 (N_17321,N_13030,N_11973);
nand U17322 (N_17322,N_13020,N_11853);
nor U17323 (N_17323,N_12092,N_12261);
nor U17324 (N_17324,N_13989,N_10919);
nor U17325 (N_17325,N_13650,N_10384);
and U17326 (N_17326,N_11834,N_10482);
nor U17327 (N_17327,N_13524,N_12289);
and U17328 (N_17328,N_14293,N_13732);
or U17329 (N_17329,N_14048,N_12016);
and U17330 (N_17330,N_14659,N_14644);
and U17331 (N_17331,N_11745,N_12009);
and U17332 (N_17332,N_13746,N_12117);
nand U17333 (N_17333,N_12658,N_10691);
or U17334 (N_17334,N_12666,N_10903);
and U17335 (N_17335,N_14692,N_10756);
nor U17336 (N_17336,N_11519,N_13281);
or U17337 (N_17337,N_10194,N_11458);
nor U17338 (N_17338,N_14348,N_12917);
nand U17339 (N_17339,N_14397,N_13145);
xnor U17340 (N_17340,N_13441,N_11277);
and U17341 (N_17341,N_10406,N_12409);
xnor U17342 (N_17342,N_13004,N_11473);
or U17343 (N_17343,N_11283,N_12489);
xnor U17344 (N_17344,N_13550,N_11435);
and U17345 (N_17345,N_12481,N_12106);
and U17346 (N_17346,N_13128,N_12626);
or U17347 (N_17347,N_14192,N_10484);
nor U17348 (N_17348,N_11057,N_12164);
nand U17349 (N_17349,N_10421,N_11780);
or U17350 (N_17350,N_10343,N_14795);
nand U17351 (N_17351,N_10218,N_10430);
nand U17352 (N_17352,N_10224,N_14677);
nor U17353 (N_17353,N_11391,N_10261);
nor U17354 (N_17354,N_11702,N_10035);
xnor U17355 (N_17355,N_13897,N_12636);
and U17356 (N_17356,N_10003,N_12132);
nor U17357 (N_17357,N_12505,N_12370);
nor U17358 (N_17358,N_11090,N_12613);
and U17359 (N_17359,N_11456,N_10254);
or U17360 (N_17360,N_11610,N_13944);
or U17361 (N_17361,N_12027,N_13506);
or U17362 (N_17362,N_12782,N_14807);
nand U17363 (N_17363,N_12365,N_12020);
nand U17364 (N_17364,N_13606,N_10986);
nor U17365 (N_17365,N_11470,N_10897);
nand U17366 (N_17366,N_14498,N_13023);
nand U17367 (N_17367,N_12412,N_14590);
or U17368 (N_17368,N_14809,N_12265);
or U17369 (N_17369,N_13517,N_10712);
or U17370 (N_17370,N_12149,N_11206);
nand U17371 (N_17371,N_13724,N_12994);
and U17372 (N_17372,N_14655,N_11428);
or U17373 (N_17373,N_13353,N_10033);
nand U17374 (N_17374,N_14120,N_13146);
or U17375 (N_17375,N_10372,N_11282);
xnor U17376 (N_17376,N_14599,N_11506);
and U17377 (N_17377,N_11917,N_14087);
or U17378 (N_17378,N_12177,N_14920);
and U17379 (N_17379,N_10861,N_11157);
or U17380 (N_17380,N_13388,N_13714);
and U17381 (N_17381,N_12314,N_10596);
nor U17382 (N_17382,N_10982,N_10423);
xnor U17383 (N_17383,N_14574,N_13726);
nand U17384 (N_17384,N_14787,N_10692);
nand U17385 (N_17385,N_10192,N_14486);
or U17386 (N_17386,N_12454,N_13677);
and U17387 (N_17387,N_13859,N_13354);
nand U17388 (N_17388,N_10308,N_10219);
nand U17389 (N_17389,N_11374,N_10045);
nor U17390 (N_17390,N_12349,N_13730);
nor U17391 (N_17391,N_12952,N_13777);
and U17392 (N_17392,N_14096,N_13666);
nor U17393 (N_17393,N_10083,N_14459);
or U17394 (N_17394,N_14946,N_14982);
nand U17395 (N_17395,N_10893,N_10380);
and U17396 (N_17396,N_14822,N_14366);
and U17397 (N_17397,N_13644,N_14166);
and U17398 (N_17398,N_13473,N_14100);
or U17399 (N_17399,N_11535,N_13484);
nor U17400 (N_17400,N_12597,N_10155);
and U17401 (N_17401,N_10967,N_14608);
and U17402 (N_17402,N_11652,N_11296);
nand U17403 (N_17403,N_13568,N_13869);
or U17404 (N_17404,N_13009,N_14352);
nand U17405 (N_17405,N_13313,N_14634);
and U17406 (N_17406,N_13091,N_10968);
and U17407 (N_17407,N_14109,N_13802);
nand U17408 (N_17408,N_11889,N_12661);
and U17409 (N_17409,N_13092,N_14564);
or U17410 (N_17410,N_13130,N_13523);
nand U17411 (N_17411,N_12795,N_12988);
nand U17412 (N_17412,N_14357,N_12763);
and U17413 (N_17413,N_10907,N_13610);
or U17414 (N_17414,N_14191,N_11344);
nand U17415 (N_17415,N_10610,N_11295);
nor U17416 (N_17416,N_13315,N_11400);
nor U17417 (N_17417,N_11648,N_14301);
or U17418 (N_17418,N_10436,N_13809);
nand U17419 (N_17419,N_13151,N_10726);
nand U17420 (N_17420,N_12253,N_11165);
and U17421 (N_17421,N_12954,N_11100);
and U17422 (N_17422,N_10415,N_14549);
and U17423 (N_17423,N_10419,N_14398);
nor U17424 (N_17424,N_14093,N_11235);
and U17425 (N_17425,N_11433,N_13889);
nor U17426 (N_17426,N_13821,N_11262);
nand U17427 (N_17427,N_10774,N_14863);
nor U17428 (N_17428,N_10906,N_10137);
and U17429 (N_17429,N_14095,N_14449);
and U17430 (N_17430,N_12304,N_12347);
and U17431 (N_17431,N_12941,N_11715);
nor U17432 (N_17432,N_11393,N_13243);
nand U17433 (N_17433,N_12940,N_13940);
and U17434 (N_17434,N_10153,N_13455);
and U17435 (N_17435,N_11217,N_12427);
or U17436 (N_17436,N_11373,N_11722);
or U17437 (N_17437,N_10866,N_14427);
and U17438 (N_17438,N_12888,N_14274);
nor U17439 (N_17439,N_14253,N_11723);
nand U17440 (N_17440,N_11137,N_14702);
nor U17441 (N_17441,N_14136,N_12358);
or U17442 (N_17442,N_11051,N_13439);
nand U17443 (N_17443,N_10964,N_13995);
or U17444 (N_17444,N_13796,N_10302);
or U17445 (N_17445,N_11225,N_11232);
nor U17446 (N_17446,N_13163,N_11687);
nor U17447 (N_17447,N_11803,N_13652);
nand U17448 (N_17448,N_13696,N_10958);
nand U17449 (N_17449,N_12576,N_10728);
or U17450 (N_17450,N_13901,N_11698);
nor U17451 (N_17451,N_13827,N_10622);
nand U17452 (N_17452,N_14999,N_12775);
nand U17453 (N_17453,N_10241,N_12610);
or U17454 (N_17454,N_11971,N_14111);
nor U17455 (N_17455,N_10978,N_14642);
nor U17456 (N_17456,N_13342,N_13420);
nand U17457 (N_17457,N_13148,N_14118);
and U17458 (N_17458,N_11415,N_14052);
nand U17459 (N_17459,N_14091,N_13442);
nor U17460 (N_17460,N_11017,N_12110);
nor U17461 (N_17461,N_10658,N_10587);
and U17462 (N_17462,N_12421,N_14217);
nor U17463 (N_17463,N_14758,N_14112);
and U17464 (N_17464,N_12845,N_14675);
nand U17465 (N_17465,N_13624,N_14613);
nor U17466 (N_17466,N_11242,N_11103);
nand U17467 (N_17467,N_12931,N_14811);
or U17468 (N_17468,N_14666,N_10483);
nand U17469 (N_17469,N_14194,N_12958);
nand U17470 (N_17470,N_10256,N_14258);
nor U17471 (N_17471,N_11162,N_14823);
or U17472 (N_17472,N_12705,N_14238);
nand U17473 (N_17473,N_12334,N_10836);
or U17474 (N_17474,N_11455,N_10061);
and U17475 (N_17475,N_12759,N_11464);
or U17476 (N_17476,N_14070,N_12518);
nand U17477 (N_17477,N_11835,N_14280);
and U17478 (N_17478,N_14614,N_14165);
or U17479 (N_17479,N_11284,N_10909);
nand U17480 (N_17480,N_12885,N_13960);
or U17481 (N_17481,N_12598,N_14339);
nor U17482 (N_17482,N_13343,N_11946);
or U17483 (N_17483,N_11758,N_13723);
or U17484 (N_17484,N_11632,N_12496);
and U17485 (N_17485,N_10711,N_10651);
or U17486 (N_17486,N_12753,N_11233);
nor U17487 (N_17487,N_11547,N_12727);
and U17488 (N_17488,N_11779,N_14903);
and U17489 (N_17489,N_11362,N_13594);
and U17490 (N_17490,N_10880,N_14455);
or U17491 (N_17491,N_12585,N_12142);
nand U17492 (N_17492,N_14350,N_13768);
and U17493 (N_17493,N_10838,N_13432);
nor U17494 (N_17494,N_13948,N_11285);
or U17495 (N_17495,N_14259,N_12018);
and U17496 (N_17496,N_10402,N_14001);
and U17497 (N_17497,N_14504,N_12073);
or U17498 (N_17498,N_10116,N_11334);
nor U17499 (N_17499,N_11024,N_11302);
and U17500 (N_17500,N_14468,N_14814);
or U17501 (N_17501,N_10894,N_14396);
and U17502 (N_17502,N_10891,N_13301);
nor U17503 (N_17503,N_13106,N_11102);
or U17504 (N_17504,N_11310,N_12584);
nor U17505 (N_17505,N_12182,N_10152);
nand U17506 (N_17506,N_11548,N_14726);
or U17507 (N_17507,N_14556,N_13364);
nand U17508 (N_17508,N_13651,N_14538);
nor U17509 (N_17509,N_14228,N_13048);
nor U17510 (N_17510,N_14035,N_10681);
xor U17511 (N_17511,N_12717,N_14836);
xor U17512 (N_17512,N_12938,N_14397);
xnor U17513 (N_17513,N_14643,N_12438);
nand U17514 (N_17514,N_14101,N_13012);
or U17515 (N_17515,N_11119,N_11895);
nand U17516 (N_17516,N_10942,N_13382);
xor U17517 (N_17517,N_10111,N_11692);
nand U17518 (N_17518,N_12106,N_11708);
nor U17519 (N_17519,N_12962,N_11847);
and U17520 (N_17520,N_10139,N_12080);
or U17521 (N_17521,N_14486,N_14152);
or U17522 (N_17522,N_11180,N_14493);
and U17523 (N_17523,N_14564,N_14720);
nor U17524 (N_17524,N_13999,N_13171);
nor U17525 (N_17525,N_10406,N_10351);
and U17526 (N_17526,N_11753,N_11267);
nor U17527 (N_17527,N_13220,N_13585);
nor U17528 (N_17528,N_14803,N_14620);
nor U17529 (N_17529,N_11937,N_10923);
and U17530 (N_17530,N_10406,N_11001);
or U17531 (N_17531,N_10004,N_11117);
nor U17532 (N_17532,N_11899,N_14188);
and U17533 (N_17533,N_12024,N_11007);
or U17534 (N_17534,N_12652,N_13386);
nand U17535 (N_17535,N_10083,N_11817);
nor U17536 (N_17536,N_13316,N_10120);
nor U17537 (N_17537,N_10707,N_13090);
nor U17538 (N_17538,N_14263,N_10626);
or U17539 (N_17539,N_13350,N_12271);
and U17540 (N_17540,N_14350,N_10282);
or U17541 (N_17541,N_14002,N_11299);
nand U17542 (N_17542,N_14093,N_11262);
nand U17543 (N_17543,N_10099,N_10859);
nor U17544 (N_17544,N_11912,N_12906);
and U17545 (N_17545,N_11054,N_14599);
or U17546 (N_17546,N_11281,N_12209);
nand U17547 (N_17547,N_14916,N_12115);
nor U17548 (N_17548,N_12839,N_13308);
nor U17549 (N_17549,N_13669,N_14342);
or U17550 (N_17550,N_12484,N_12250);
nand U17551 (N_17551,N_14236,N_12934);
and U17552 (N_17552,N_10611,N_13387);
and U17553 (N_17553,N_10333,N_14857);
or U17554 (N_17554,N_10829,N_13608);
or U17555 (N_17555,N_10468,N_14235);
and U17556 (N_17556,N_11134,N_10224);
nand U17557 (N_17557,N_10926,N_13471);
and U17558 (N_17558,N_10442,N_12386);
nor U17559 (N_17559,N_14358,N_10464);
or U17560 (N_17560,N_13904,N_11598);
nand U17561 (N_17561,N_10593,N_11347);
nand U17562 (N_17562,N_11513,N_12100);
nor U17563 (N_17563,N_11139,N_11224);
nor U17564 (N_17564,N_14809,N_11928);
and U17565 (N_17565,N_10778,N_13884);
nand U17566 (N_17566,N_10276,N_11685);
nor U17567 (N_17567,N_13127,N_12995);
nor U17568 (N_17568,N_14468,N_11352);
and U17569 (N_17569,N_12958,N_13009);
and U17570 (N_17570,N_11218,N_10806);
or U17571 (N_17571,N_14084,N_11082);
and U17572 (N_17572,N_12682,N_12336);
nor U17573 (N_17573,N_11021,N_12334);
nor U17574 (N_17574,N_12049,N_11565);
and U17575 (N_17575,N_13348,N_13217);
nand U17576 (N_17576,N_14300,N_10468);
or U17577 (N_17577,N_10990,N_10649);
and U17578 (N_17578,N_14786,N_11822);
nand U17579 (N_17579,N_13944,N_14680);
or U17580 (N_17580,N_13316,N_14755);
nand U17581 (N_17581,N_11239,N_14884);
or U17582 (N_17582,N_13620,N_13496);
nand U17583 (N_17583,N_12982,N_13516);
or U17584 (N_17584,N_14194,N_11024);
or U17585 (N_17585,N_14838,N_11245);
nand U17586 (N_17586,N_14540,N_12198);
nand U17587 (N_17587,N_13446,N_13422);
nand U17588 (N_17588,N_10557,N_11461);
and U17589 (N_17589,N_11901,N_12405);
or U17590 (N_17590,N_11016,N_11935);
nand U17591 (N_17591,N_14980,N_11414);
nand U17592 (N_17592,N_12186,N_13603);
nand U17593 (N_17593,N_10837,N_10300);
nand U17594 (N_17594,N_10705,N_12259);
nor U17595 (N_17595,N_13232,N_12717);
nor U17596 (N_17596,N_13911,N_12362);
nor U17597 (N_17597,N_14069,N_11044);
nor U17598 (N_17598,N_10834,N_14966);
or U17599 (N_17599,N_13704,N_14620);
or U17600 (N_17600,N_11910,N_14573);
nand U17601 (N_17601,N_13397,N_11019);
nand U17602 (N_17602,N_10641,N_10958);
or U17603 (N_17603,N_11457,N_12306);
nand U17604 (N_17604,N_10642,N_13214);
xor U17605 (N_17605,N_11964,N_10533);
or U17606 (N_17606,N_14318,N_12624);
nand U17607 (N_17607,N_12276,N_12715);
and U17608 (N_17608,N_10769,N_12718);
and U17609 (N_17609,N_11563,N_11480);
nor U17610 (N_17610,N_10983,N_13137);
nand U17611 (N_17611,N_12614,N_12608);
and U17612 (N_17612,N_11339,N_12933);
or U17613 (N_17613,N_14093,N_13772);
and U17614 (N_17614,N_13105,N_14929);
and U17615 (N_17615,N_13026,N_12653);
and U17616 (N_17616,N_11549,N_11293);
or U17617 (N_17617,N_13495,N_11626);
and U17618 (N_17618,N_10627,N_11821);
and U17619 (N_17619,N_14472,N_14023);
nor U17620 (N_17620,N_11525,N_13200);
or U17621 (N_17621,N_12702,N_14502);
or U17622 (N_17622,N_12567,N_14903);
and U17623 (N_17623,N_10686,N_12240);
or U17624 (N_17624,N_12308,N_14128);
and U17625 (N_17625,N_10641,N_10094);
nand U17626 (N_17626,N_13453,N_11753);
nor U17627 (N_17627,N_11212,N_12538);
or U17628 (N_17628,N_12397,N_12589);
nand U17629 (N_17629,N_12572,N_14264);
or U17630 (N_17630,N_12888,N_14741);
or U17631 (N_17631,N_13696,N_13774);
and U17632 (N_17632,N_12317,N_11243);
and U17633 (N_17633,N_14892,N_10532);
or U17634 (N_17634,N_11707,N_11482);
and U17635 (N_17635,N_11982,N_14402);
nor U17636 (N_17636,N_12965,N_11407);
nor U17637 (N_17637,N_10416,N_14655);
and U17638 (N_17638,N_10987,N_11048);
nand U17639 (N_17639,N_14280,N_12166);
nand U17640 (N_17640,N_10874,N_12433);
and U17641 (N_17641,N_10658,N_13355);
and U17642 (N_17642,N_12658,N_11420);
and U17643 (N_17643,N_13917,N_12608);
nand U17644 (N_17644,N_13807,N_11294);
nand U17645 (N_17645,N_14536,N_11563);
or U17646 (N_17646,N_13919,N_12900);
nor U17647 (N_17647,N_11046,N_14312);
and U17648 (N_17648,N_13046,N_12987);
and U17649 (N_17649,N_11611,N_14638);
or U17650 (N_17650,N_12428,N_13768);
nor U17651 (N_17651,N_13015,N_12576);
nand U17652 (N_17652,N_11361,N_11206);
nor U17653 (N_17653,N_12170,N_11288);
or U17654 (N_17654,N_13425,N_13634);
and U17655 (N_17655,N_10145,N_12076);
nand U17656 (N_17656,N_12735,N_14824);
nor U17657 (N_17657,N_10958,N_12415);
nand U17658 (N_17658,N_12771,N_11830);
nor U17659 (N_17659,N_14948,N_10139);
and U17660 (N_17660,N_10163,N_12594);
or U17661 (N_17661,N_12616,N_10977);
or U17662 (N_17662,N_11426,N_14148);
or U17663 (N_17663,N_12246,N_14790);
and U17664 (N_17664,N_12656,N_13223);
or U17665 (N_17665,N_10501,N_13496);
or U17666 (N_17666,N_13621,N_10597);
nor U17667 (N_17667,N_10098,N_11195);
and U17668 (N_17668,N_11641,N_10756);
or U17669 (N_17669,N_11357,N_11982);
nand U17670 (N_17670,N_14649,N_11848);
or U17671 (N_17671,N_11338,N_14860);
nor U17672 (N_17672,N_10801,N_11849);
or U17673 (N_17673,N_12342,N_13463);
nor U17674 (N_17674,N_13635,N_11612);
nor U17675 (N_17675,N_11192,N_10532);
and U17676 (N_17676,N_11582,N_11596);
and U17677 (N_17677,N_11762,N_11535);
nand U17678 (N_17678,N_14570,N_11182);
or U17679 (N_17679,N_10183,N_10932);
nor U17680 (N_17680,N_14472,N_11950);
or U17681 (N_17681,N_11897,N_14704);
nand U17682 (N_17682,N_11128,N_12402);
and U17683 (N_17683,N_14015,N_12976);
and U17684 (N_17684,N_10930,N_10216);
nand U17685 (N_17685,N_10977,N_10243);
nor U17686 (N_17686,N_11485,N_10514);
or U17687 (N_17687,N_12752,N_10302);
nor U17688 (N_17688,N_10567,N_14694);
and U17689 (N_17689,N_14782,N_11604);
and U17690 (N_17690,N_14672,N_13873);
or U17691 (N_17691,N_13577,N_12884);
nor U17692 (N_17692,N_14726,N_13620);
nor U17693 (N_17693,N_10067,N_11316);
or U17694 (N_17694,N_14138,N_13284);
xnor U17695 (N_17695,N_10481,N_11551);
nand U17696 (N_17696,N_13678,N_14017);
nand U17697 (N_17697,N_14018,N_14501);
nand U17698 (N_17698,N_14877,N_12510);
nand U17699 (N_17699,N_12208,N_13999);
nand U17700 (N_17700,N_14938,N_11575);
or U17701 (N_17701,N_13944,N_14724);
nor U17702 (N_17702,N_14374,N_11326);
or U17703 (N_17703,N_12488,N_11076);
and U17704 (N_17704,N_11941,N_11809);
nor U17705 (N_17705,N_13978,N_10480);
nand U17706 (N_17706,N_11077,N_14648);
nand U17707 (N_17707,N_12331,N_10509);
nor U17708 (N_17708,N_13118,N_13790);
nand U17709 (N_17709,N_14175,N_14512);
or U17710 (N_17710,N_13924,N_10691);
nand U17711 (N_17711,N_11920,N_13332);
nor U17712 (N_17712,N_10866,N_13903);
nand U17713 (N_17713,N_10853,N_12479);
nand U17714 (N_17714,N_13760,N_11473);
nor U17715 (N_17715,N_10393,N_14832);
nor U17716 (N_17716,N_11358,N_11331);
nor U17717 (N_17717,N_14383,N_14037);
or U17718 (N_17718,N_14793,N_12301);
nand U17719 (N_17719,N_13836,N_10613);
or U17720 (N_17720,N_13306,N_13758);
nand U17721 (N_17721,N_10121,N_12851);
or U17722 (N_17722,N_11112,N_14418);
or U17723 (N_17723,N_13290,N_12642);
nand U17724 (N_17724,N_10215,N_13761);
nand U17725 (N_17725,N_14826,N_13906);
nand U17726 (N_17726,N_14230,N_12893);
nor U17727 (N_17727,N_13579,N_14357);
nor U17728 (N_17728,N_12233,N_14202);
nor U17729 (N_17729,N_11526,N_13464);
or U17730 (N_17730,N_14238,N_10278);
and U17731 (N_17731,N_10723,N_11780);
and U17732 (N_17732,N_10332,N_12133);
nand U17733 (N_17733,N_11381,N_12062);
and U17734 (N_17734,N_12650,N_11633);
and U17735 (N_17735,N_12645,N_13074);
nor U17736 (N_17736,N_10879,N_10560);
or U17737 (N_17737,N_11420,N_14066);
or U17738 (N_17738,N_10145,N_12783);
nand U17739 (N_17739,N_11958,N_13049);
nand U17740 (N_17740,N_12541,N_11595);
xor U17741 (N_17741,N_14761,N_10335);
nand U17742 (N_17742,N_10958,N_10480);
nand U17743 (N_17743,N_11974,N_13439);
nor U17744 (N_17744,N_10170,N_14928);
nor U17745 (N_17745,N_10775,N_13123);
and U17746 (N_17746,N_12492,N_12195);
nor U17747 (N_17747,N_14326,N_10108);
or U17748 (N_17748,N_13428,N_13090);
or U17749 (N_17749,N_14518,N_11091);
nor U17750 (N_17750,N_12827,N_12828);
and U17751 (N_17751,N_11508,N_13366);
nand U17752 (N_17752,N_10773,N_10851);
nor U17753 (N_17753,N_13999,N_10266);
nand U17754 (N_17754,N_12305,N_14154);
nand U17755 (N_17755,N_13507,N_13715);
nor U17756 (N_17756,N_12255,N_11344);
and U17757 (N_17757,N_13687,N_13761);
nand U17758 (N_17758,N_11877,N_11246);
nand U17759 (N_17759,N_14301,N_12709);
nand U17760 (N_17760,N_10727,N_12213);
or U17761 (N_17761,N_11123,N_14448);
nor U17762 (N_17762,N_13430,N_11448);
and U17763 (N_17763,N_13094,N_13260);
nor U17764 (N_17764,N_11534,N_13919);
nand U17765 (N_17765,N_10372,N_11647);
and U17766 (N_17766,N_12541,N_10481);
and U17767 (N_17767,N_10465,N_11503);
nor U17768 (N_17768,N_14416,N_10444);
and U17769 (N_17769,N_10351,N_11347);
nor U17770 (N_17770,N_11266,N_13239);
nand U17771 (N_17771,N_11226,N_12516);
nand U17772 (N_17772,N_13092,N_11351);
and U17773 (N_17773,N_12613,N_12735);
nand U17774 (N_17774,N_13076,N_11527);
and U17775 (N_17775,N_11737,N_14225);
nand U17776 (N_17776,N_13925,N_11750);
and U17777 (N_17777,N_11730,N_14924);
or U17778 (N_17778,N_14691,N_13746);
nor U17779 (N_17779,N_10833,N_10073);
or U17780 (N_17780,N_14500,N_13437);
and U17781 (N_17781,N_11549,N_12025);
nor U17782 (N_17782,N_11314,N_12960);
xor U17783 (N_17783,N_11940,N_10193);
or U17784 (N_17784,N_11440,N_13810);
nand U17785 (N_17785,N_10993,N_11155);
nand U17786 (N_17786,N_12804,N_10700);
nand U17787 (N_17787,N_12917,N_13028);
and U17788 (N_17788,N_12895,N_13153);
nor U17789 (N_17789,N_14685,N_13415);
or U17790 (N_17790,N_12473,N_10180);
and U17791 (N_17791,N_12905,N_10166);
and U17792 (N_17792,N_12183,N_13962);
and U17793 (N_17793,N_10575,N_10856);
and U17794 (N_17794,N_13378,N_11838);
or U17795 (N_17795,N_14512,N_10304);
nand U17796 (N_17796,N_12147,N_14745);
and U17797 (N_17797,N_13403,N_13687);
and U17798 (N_17798,N_10467,N_11366);
nor U17799 (N_17799,N_14009,N_14414);
or U17800 (N_17800,N_13102,N_14191);
nor U17801 (N_17801,N_13000,N_14452);
or U17802 (N_17802,N_14706,N_14033);
nand U17803 (N_17803,N_10837,N_10853);
nand U17804 (N_17804,N_12562,N_10350);
nand U17805 (N_17805,N_10602,N_11833);
nor U17806 (N_17806,N_14541,N_13207);
nor U17807 (N_17807,N_14081,N_11124);
and U17808 (N_17808,N_12821,N_14541);
nand U17809 (N_17809,N_10702,N_12078);
nand U17810 (N_17810,N_12467,N_10721);
xor U17811 (N_17811,N_12033,N_12337);
or U17812 (N_17812,N_10336,N_12747);
and U17813 (N_17813,N_10738,N_14637);
or U17814 (N_17814,N_13649,N_14757);
and U17815 (N_17815,N_13013,N_11830);
or U17816 (N_17816,N_10032,N_12044);
nand U17817 (N_17817,N_11130,N_14788);
nor U17818 (N_17818,N_10022,N_11967);
or U17819 (N_17819,N_10176,N_12722);
or U17820 (N_17820,N_14692,N_12646);
nand U17821 (N_17821,N_12303,N_14498);
and U17822 (N_17822,N_11107,N_14374);
nor U17823 (N_17823,N_11514,N_10122);
and U17824 (N_17824,N_12508,N_13740);
nand U17825 (N_17825,N_14920,N_14453);
and U17826 (N_17826,N_14169,N_11672);
and U17827 (N_17827,N_12486,N_10872);
or U17828 (N_17828,N_12665,N_11012);
or U17829 (N_17829,N_14382,N_11402);
xnor U17830 (N_17830,N_14514,N_14592);
or U17831 (N_17831,N_11100,N_10911);
or U17832 (N_17832,N_11346,N_12420);
nand U17833 (N_17833,N_11988,N_12106);
or U17834 (N_17834,N_13747,N_11076);
nor U17835 (N_17835,N_10860,N_10388);
nor U17836 (N_17836,N_10172,N_14588);
and U17837 (N_17837,N_11598,N_14610);
nand U17838 (N_17838,N_10462,N_13639);
or U17839 (N_17839,N_12607,N_13670);
nand U17840 (N_17840,N_12095,N_12508);
or U17841 (N_17841,N_14838,N_11370);
and U17842 (N_17842,N_11328,N_12816);
and U17843 (N_17843,N_14905,N_14144);
nor U17844 (N_17844,N_14563,N_11376);
nor U17845 (N_17845,N_11656,N_14635);
and U17846 (N_17846,N_12653,N_12994);
or U17847 (N_17847,N_13094,N_13572);
or U17848 (N_17848,N_12371,N_13607);
nand U17849 (N_17849,N_13529,N_14236);
or U17850 (N_17850,N_12457,N_11950);
and U17851 (N_17851,N_11832,N_13263);
nand U17852 (N_17852,N_10550,N_13387);
nor U17853 (N_17853,N_14284,N_14550);
nor U17854 (N_17854,N_13313,N_12735);
nor U17855 (N_17855,N_13055,N_13174);
nand U17856 (N_17856,N_10182,N_13765);
nand U17857 (N_17857,N_14591,N_13201);
nor U17858 (N_17858,N_10455,N_14313);
and U17859 (N_17859,N_12658,N_13086);
nor U17860 (N_17860,N_12385,N_11051);
nand U17861 (N_17861,N_11997,N_11971);
nor U17862 (N_17862,N_12875,N_13897);
nor U17863 (N_17863,N_12067,N_10190);
or U17864 (N_17864,N_13438,N_12756);
nand U17865 (N_17865,N_10258,N_10437);
or U17866 (N_17866,N_10286,N_11479);
nor U17867 (N_17867,N_14427,N_11933);
nand U17868 (N_17868,N_11438,N_14428);
nor U17869 (N_17869,N_14611,N_14028);
nor U17870 (N_17870,N_13579,N_13123);
nand U17871 (N_17871,N_11814,N_12748);
xor U17872 (N_17872,N_13648,N_12837);
nor U17873 (N_17873,N_12591,N_11401);
nand U17874 (N_17874,N_11993,N_13858);
nor U17875 (N_17875,N_12836,N_12212);
nor U17876 (N_17876,N_13959,N_14880);
and U17877 (N_17877,N_10251,N_14054);
and U17878 (N_17878,N_12134,N_10783);
and U17879 (N_17879,N_11374,N_14284);
and U17880 (N_17880,N_13861,N_12102);
or U17881 (N_17881,N_10517,N_14266);
nor U17882 (N_17882,N_11666,N_14018);
and U17883 (N_17883,N_10043,N_14991);
or U17884 (N_17884,N_10811,N_11883);
nor U17885 (N_17885,N_11464,N_10724);
and U17886 (N_17886,N_11833,N_14383);
nor U17887 (N_17887,N_14168,N_13633);
nand U17888 (N_17888,N_13882,N_11269);
and U17889 (N_17889,N_11477,N_14826);
nor U17890 (N_17890,N_11311,N_11633);
and U17891 (N_17891,N_11343,N_14632);
and U17892 (N_17892,N_10404,N_11110);
nor U17893 (N_17893,N_12631,N_12589);
nand U17894 (N_17894,N_11821,N_12212);
nor U17895 (N_17895,N_12286,N_10828);
xnor U17896 (N_17896,N_14168,N_10367);
or U17897 (N_17897,N_11512,N_12190);
nor U17898 (N_17898,N_12009,N_12405);
or U17899 (N_17899,N_11877,N_13267);
or U17900 (N_17900,N_11412,N_10784);
or U17901 (N_17901,N_13798,N_12128);
and U17902 (N_17902,N_13690,N_13023);
or U17903 (N_17903,N_14103,N_10462);
nand U17904 (N_17904,N_11069,N_10754);
nor U17905 (N_17905,N_14355,N_12883);
and U17906 (N_17906,N_10787,N_12536);
nor U17907 (N_17907,N_14698,N_10002);
nor U17908 (N_17908,N_10764,N_11214);
nand U17909 (N_17909,N_10148,N_11805);
nand U17910 (N_17910,N_14601,N_11500);
nand U17911 (N_17911,N_10551,N_13370);
nand U17912 (N_17912,N_10545,N_10565);
and U17913 (N_17913,N_12414,N_14055);
or U17914 (N_17914,N_13255,N_13936);
nand U17915 (N_17915,N_11146,N_10999);
nor U17916 (N_17916,N_11702,N_12333);
or U17917 (N_17917,N_10253,N_14818);
nand U17918 (N_17918,N_11436,N_11413);
nand U17919 (N_17919,N_12013,N_10165);
nand U17920 (N_17920,N_13466,N_11194);
nor U17921 (N_17921,N_10128,N_11470);
or U17922 (N_17922,N_14512,N_14390);
or U17923 (N_17923,N_10404,N_13370);
or U17924 (N_17924,N_12909,N_10249);
nor U17925 (N_17925,N_13481,N_13111);
and U17926 (N_17926,N_13986,N_14351);
and U17927 (N_17927,N_14941,N_14957);
or U17928 (N_17928,N_10828,N_12193);
or U17929 (N_17929,N_11652,N_11935);
and U17930 (N_17930,N_13520,N_11056);
and U17931 (N_17931,N_12558,N_12689);
nand U17932 (N_17932,N_14780,N_12203);
nand U17933 (N_17933,N_12871,N_13961);
and U17934 (N_17934,N_12184,N_10877);
nor U17935 (N_17935,N_13770,N_10854);
or U17936 (N_17936,N_10762,N_14610);
and U17937 (N_17937,N_14845,N_13758);
nand U17938 (N_17938,N_14812,N_12090);
or U17939 (N_17939,N_11242,N_14832);
or U17940 (N_17940,N_11219,N_10734);
and U17941 (N_17941,N_10259,N_12988);
and U17942 (N_17942,N_11754,N_14868);
xnor U17943 (N_17943,N_14920,N_11177);
nand U17944 (N_17944,N_13706,N_10920);
and U17945 (N_17945,N_13497,N_11966);
or U17946 (N_17946,N_11097,N_11241);
or U17947 (N_17947,N_14411,N_10297);
nor U17948 (N_17948,N_10402,N_11135);
nor U17949 (N_17949,N_14122,N_13788);
and U17950 (N_17950,N_11763,N_12127);
nor U17951 (N_17951,N_14489,N_12430);
and U17952 (N_17952,N_10827,N_13608);
nor U17953 (N_17953,N_11754,N_10922);
nand U17954 (N_17954,N_11627,N_13238);
nor U17955 (N_17955,N_12020,N_12489);
and U17956 (N_17956,N_11109,N_12640);
nor U17957 (N_17957,N_13770,N_13517);
nand U17958 (N_17958,N_10121,N_10431);
and U17959 (N_17959,N_14640,N_13786);
or U17960 (N_17960,N_14379,N_14970);
and U17961 (N_17961,N_13101,N_14443);
nand U17962 (N_17962,N_14362,N_11827);
or U17963 (N_17963,N_12814,N_10473);
or U17964 (N_17964,N_14758,N_12897);
nor U17965 (N_17965,N_14624,N_10104);
or U17966 (N_17966,N_13047,N_14162);
and U17967 (N_17967,N_10875,N_11070);
or U17968 (N_17968,N_12801,N_12016);
or U17969 (N_17969,N_11548,N_13720);
and U17970 (N_17970,N_11146,N_14573);
and U17971 (N_17971,N_11561,N_10813);
and U17972 (N_17972,N_10172,N_10418);
and U17973 (N_17973,N_10295,N_14381);
nor U17974 (N_17974,N_14951,N_10666);
nor U17975 (N_17975,N_13863,N_11092);
or U17976 (N_17976,N_12699,N_11815);
and U17977 (N_17977,N_10891,N_13671);
nor U17978 (N_17978,N_14025,N_11080);
nor U17979 (N_17979,N_10697,N_11229);
or U17980 (N_17980,N_10771,N_14390);
or U17981 (N_17981,N_10613,N_13038);
and U17982 (N_17982,N_14062,N_11620);
nor U17983 (N_17983,N_14410,N_14415);
nand U17984 (N_17984,N_10817,N_12610);
or U17985 (N_17985,N_12533,N_12107);
and U17986 (N_17986,N_11983,N_12572);
and U17987 (N_17987,N_11674,N_14243);
and U17988 (N_17988,N_11660,N_12284);
nor U17989 (N_17989,N_12706,N_12584);
nor U17990 (N_17990,N_13390,N_12197);
or U17991 (N_17991,N_13522,N_13865);
nand U17992 (N_17992,N_14113,N_10182);
or U17993 (N_17993,N_10518,N_14889);
or U17994 (N_17994,N_12944,N_13782);
or U17995 (N_17995,N_11806,N_13867);
nand U17996 (N_17996,N_10532,N_14007);
nand U17997 (N_17997,N_10500,N_12491);
or U17998 (N_17998,N_14793,N_14836);
and U17999 (N_17999,N_12685,N_14239);
and U18000 (N_18000,N_13878,N_14241);
xnor U18001 (N_18001,N_12481,N_11325);
nor U18002 (N_18002,N_11325,N_14104);
and U18003 (N_18003,N_11945,N_14181);
or U18004 (N_18004,N_10965,N_11316);
and U18005 (N_18005,N_13615,N_11465);
or U18006 (N_18006,N_11708,N_12930);
and U18007 (N_18007,N_11804,N_12578);
or U18008 (N_18008,N_13111,N_10772);
or U18009 (N_18009,N_10502,N_14688);
or U18010 (N_18010,N_12337,N_13931);
xnor U18011 (N_18011,N_13157,N_14844);
nor U18012 (N_18012,N_14295,N_12292);
nor U18013 (N_18013,N_10227,N_11437);
and U18014 (N_18014,N_13150,N_11435);
nor U18015 (N_18015,N_11097,N_13366);
or U18016 (N_18016,N_12035,N_12344);
nor U18017 (N_18017,N_13140,N_12385);
nand U18018 (N_18018,N_12706,N_13513);
nor U18019 (N_18019,N_13448,N_14141);
nand U18020 (N_18020,N_14319,N_14020);
nand U18021 (N_18021,N_10912,N_12515);
nor U18022 (N_18022,N_14474,N_10238);
nand U18023 (N_18023,N_13000,N_14664);
and U18024 (N_18024,N_14628,N_10392);
or U18025 (N_18025,N_10810,N_14839);
nand U18026 (N_18026,N_12920,N_12886);
nor U18027 (N_18027,N_14702,N_14877);
nand U18028 (N_18028,N_10021,N_12316);
nor U18029 (N_18029,N_13720,N_13369);
and U18030 (N_18030,N_13012,N_10790);
or U18031 (N_18031,N_14142,N_12989);
and U18032 (N_18032,N_11441,N_14039);
and U18033 (N_18033,N_14550,N_11760);
and U18034 (N_18034,N_12532,N_13056);
nand U18035 (N_18035,N_11000,N_14743);
nor U18036 (N_18036,N_13604,N_13005);
and U18037 (N_18037,N_14135,N_13835);
nand U18038 (N_18038,N_13880,N_11919);
nor U18039 (N_18039,N_13747,N_14135);
or U18040 (N_18040,N_14688,N_13224);
nor U18041 (N_18041,N_14367,N_11131);
nor U18042 (N_18042,N_14036,N_12279);
and U18043 (N_18043,N_13609,N_12244);
or U18044 (N_18044,N_11306,N_13484);
and U18045 (N_18045,N_13158,N_14316);
nor U18046 (N_18046,N_13986,N_14432);
or U18047 (N_18047,N_10695,N_12409);
and U18048 (N_18048,N_13087,N_11963);
nand U18049 (N_18049,N_10936,N_10794);
nand U18050 (N_18050,N_13031,N_10372);
or U18051 (N_18051,N_12488,N_11588);
nor U18052 (N_18052,N_10873,N_12196);
and U18053 (N_18053,N_12687,N_14722);
and U18054 (N_18054,N_12412,N_13358);
and U18055 (N_18055,N_13748,N_14371);
nand U18056 (N_18056,N_13738,N_12738);
nor U18057 (N_18057,N_12534,N_11290);
nor U18058 (N_18058,N_14281,N_10373);
or U18059 (N_18059,N_11353,N_12738);
nor U18060 (N_18060,N_11091,N_11537);
nand U18061 (N_18061,N_13597,N_11760);
or U18062 (N_18062,N_12542,N_14096);
nor U18063 (N_18063,N_11222,N_13686);
nor U18064 (N_18064,N_10154,N_13680);
or U18065 (N_18065,N_10505,N_14403);
nor U18066 (N_18066,N_14214,N_10049);
or U18067 (N_18067,N_11721,N_11865);
or U18068 (N_18068,N_11591,N_11523);
nand U18069 (N_18069,N_14624,N_10447);
nand U18070 (N_18070,N_11153,N_10406);
or U18071 (N_18071,N_13053,N_12492);
or U18072 (N_18072,N_11532,N_13123);
nor U18073 (N_18073,N_14964,N_13254);
nor U18074 (N_18074,N_13923,N_13181);
or U18075 (N_18075,N_10763,N_12889);
nand U18076 (N_18076,N_11977,N_11875);
and U18077 (N_18077,N_12158,N_13830);
or U18078 (N_18078,N_10827,N_14613);
nor U18079 (N_18079,N_14712,N_14484);
and U18080 (N_18080,N_13224,N_11683);
nand U18081 (N_18081,N_13402,N_10715);
nor U18082 (N_18082,N_12977,N_10541);
nand U18083 (N_18083,N_10815,N_11652);
nand U18084 (N_18084,N_14949,N_14968);
or U18085 (N_18085,N_11016,N_10024);
nor U18086 (N_18086,N_11106,N_13096);
and U18087 (N_18087,N_10291,N_14323);
or U18088 (N_18088,N_12248,N_11245);
and U18089 (N_18089,N_13161,N_10499);
or U18090 (N_18090,N_10841,N_12621);
nand U18091 (N_18091,N_12381,N_14090);
and U18092 (N_18092,N_11798,N_14039);
and U18093 (N_18093,N_12812,N_13250);
nand U18094 (N_18094,N_11573,N_12180);
or U18095 (N_18095,N_10980,N_13793);
xor U18096 (N_18096,N_12138,N_14572);
or U18097 (N_18097,N_11266,N_12892);
nand U18098 (N_18098,N_14619,N_14574);
nand U18099 (N_18099,N_13732,N_10607);
nand U18100 (N_18100,N_11143,N_11606);
nand U18101 (N_18101,N_11971,N_13434);
or U18102 (N_18102,N_11301,N_14621);
nand U18103 (N_18103,N_13099,N_10842);
and U18104 (N_18104,N_10798,N_14136);
or U18105 (N_18105,N_13255,N_14587);
or U18106 (N_18106,N_12062,N_11618);
and U18107 (N_18107,N_14890,N_13210);
or U18108 (N_18108,N_12629,N_14174);
nand U18109 (N_18109,N_11527,N_11497);
nand U18110 (N_18110,N_13167,N_10497);
or U18111 (N_18111,N_14158,N_11478);
and U18112 (N_18112,N_12009,N_12474);
nor U18113 (N_18113,N_13060,N_10589);
nor U18114 (N_18114,N_13440,N_14006);
or U18115 (N_18115,N_12922,N_13736);
and U18116 (N_18116,N_11184,N_13613);
nand U18117 (N_18117,N_14464,N_12322);
nor U18118 (N_18118,N_11939,N_10593);
nand U18119 (N_18119,N_14370,N_12202);
nand U18120 (N_18120,N_10186,N_13458);
nand U18121 (N_18121,N_11903,N_12400);
nor U18122 (N_18122,N_13010,N_13898);
or U18123 (N_18123,N_11888,N_12798);
nand U18124 (N_18124,N_10440,N_13111);
nor U18125 (N_18125,N_14668,N_12668);
nor U18126 (N_18126,N_12246,N_12531);
nor U18127 (N_18127,N_11189,N_12300);
nand U18128 (N_18128,N_12945,N_13644);
or U18129 (N_18129,N_12302,N_13954);
nand U18130 (N_18130,N_14949,N_10141);
nor U18131 (N_18131,N_11917,N_14195);
nor U18132 (N_18132,N_10656,N_14720);
nand U18133 (N_18133,N_10761,N_14187);
and U18134 (N_18134,N_12045,N_12788);
nand U18135 (N_18135,N_14314,N_10969);
and U18136 (N_18136,N_13521,N_11600);
or U18137 (N_18137,N_11131,N_14175);
nor U18138 (N_18138,N_13948,N_11292);
nand U18139 (N_18139,N_14496,N_12935);
or U18140 (N_18140,N_10638,N_11328);
xnor U18141 (N_18141,N_10649,N_13315);
nand U18142 (N_18142,N_10307,N_13009);
nand U18143 (N_18143,N_12829,N_10165);
nand U18144 (N_18144,N_12379,N_13085);
and U18145 (N_18145,N_12630,N_13633);
nand U18146 (N_18146,N_14620,N_12794);
or U18147 (N_18147,N_11007,N_11888);
nor U18148 (N_18148,N_10921,N_10970);
nand U18149 (N_18149,N_14512,N_13558);
or U18150 (N_18150,N_10447,N_11100);
and U18151 (N_18151,N_13394,N_10676);
nor U18152 (N_18152,N_11768,N_14773);
and U18153 (N_18153,N_10513,N_13712);
and U18154 (N_18154,N_13435,N_10798);
and U18155 (N_18155,N_10799,N_14532);
or U18156 (N_18156,N_11278,N_14535);
nor U18157 (N_18157,N_14751,N_13471);
and U18158 (N_18158,N_14052,N_11095);
and U18159 (N_18159,N_14297,N_13134);
or U18160 (N_18160,N_13433,N_12043);
or U18161 (N_18161,N_14585,N_10665);
and U18162 (N_18162,N_13177,N_11063);
nand U18163 (N_18163,N_10593,N_11644);
nand U18164 (N_18164,N_10114,N_13939);
and U18165 (N_18165,N_14213,N_13326);
and U18166 (N_18166,N_14700,N_11040);
xor U18167 (N_18167,N_13813,N_13801);
nand U18168 (N_18168,N_10397,N_10186);
or U18169 (N_18169,N_13480,N_12329);
or U18170 (N_18170,N_11839,N_11485);
and U18171 (N_18171,N_14597,N_14527);
and U18172 (N_18172,N_13709,N_10549);
and U18173 (N_18173,N_11197,N_11395);
nand U18174 (N_18174,N_13691,N_13287);
nor U18175 (N_18175,N_13493,N_11398);
nor U18176 (N_18176,N_10415,N_10096);
and U18177 (N_18177,N_13749,N_11700);
or U18178 (N_18178,N_14716,N_11159);
nor U18179 (N_18179,N_11767,N_14438);
nand U18180 (N_18180,N_11154,N_10689);
nor U18181 (N_18181,N_12520,N_14289);
or U18182 (N_18182,N_14010,N_13897);
and U18183 (N_18183,N_11498,N_11684);
or U18184 (N_18184,N_14575,N_13241);
nor U18185 (N_18185,N_10479,N_12992);
and U18186 (N_18186,N_14040,N_11026);
and U18187 (N_18187,N_12154,N_12706);
nor U18188 (N_18188,N_13549,N_10354);
nor U18189 (N_18189,N_10590,N_12792);
and U18190 (N_18190,N_14487,N_14772);
or U18191 (N_18191,N_13963,N_10641);
or U18192 (N_18192,N_13646,N_14773);
or U18193 (N_18193,N_11472,N_12971);
nand U18194 (N_18194,N_12828,N_10486);
or U18195 (N_18195,N_12930,N_11612);
nand U18196 (N_18196,N_12413,N_11000);
nand U18197 (N_18197,N_11804,N_13555);
nor U18198 (N_18198,N_12543,N_11323);
nor U18199 (N_18199,N_14465,N_13630);
nand U18200 (N_18200,N_13380,N_14738);
and U18201 (N_18201,N_14071,N_12876);
nand U18202 (N_18202,N_12345,N_11080);
nand U18203 (N_18203,N_14443,N_11750);
or U18204 (N_18204,N_14675,N_11093);
or U18205 (N_18205,N_13785,N_13950);
nor U18206 (N_18206,N_14585,N_13612);
and U18207 (N_18207,N_10374,N_14003);
and U18208 (N_18208,N_12354,N_14244);
and U18209 (N_18209,N_13321,N_14949);
and U18210 (N_18210,N_10007,N_11777);
nand U18211 (N_18211,N_11451,N_11373);
and U18212 (N_18212,N_11737,N_11496);
nand U18213 (N_18213,N_11682,N_13433);
nor U18214 (N_18214,N_10338,N_10368);
and U18215 (N_18215,N_12061,N_13948);
nor U18216 (N_18216,N_12946,N_12415);
or U18217 (N_18217,N_12855,N_14313);
nor U18218 (N_18218,N_13295,N_14474);
and U18219 (N_18219,N_10608,N_10318);
nor U18220 (N_18220,N_11465,N_11612);
nor U18221 (N_18221,N_12073,N_14129);
nor U18222 (N_18222,N_14960,N_14810);
and U18223 (N_18223,N_10220,N_11369);
nand U18224 (N_18224,N_11602,N_13100);
nand U18225 (N_18225,N_10486,N_10783);
and U18226 (N_18226,N_11054,N_11676);
nor U18227 (N_18227,N_13161,N_12125);
and U18228 (N_18228,N_13112,N_13179);
and U18229 (N_18229,N_13687,N_14692);
nand U18230 (N_18230,N_14204,N_10172);
or U18231 (N_18231,N_11745,N_14424);
and U18232 (N_18232,N_14055,N_10195);
or U18233 (N_18233,N_11567,N_10538);
xnor U18234 (N_18234,N_10635,N_12604);
or U18235 (N_18235,N_13953,N_10413);
or U18236 (N_18236,N_13795,N_11450);
nor U18237 (N_18237,N_14615,N_11241);
or U18238 (N_18238,N_13979,N_14865);
and U18239 (N_18239,N_13692,N_14854);
nand U18240 (N_18240,N_11513,N_10270);
and U18241 (N_18241,N_12631,N_13824);
and U18242 (N_18242,N_11992,N_13510);
or U18243 (N_18243,N_12056,N_10565);
nand U18244 (N_18244,N_12563,N_11197);
nand U18245 (N_18245,N_10861,N_13868);
or U18246 (N_18246,N_10296,N_10532);
nor U18247 (N_18247,N_13110,N_10980);
or U18248 (N_18248,N_10335,N_10152);
or U18249 (N_18249,N_13051,N_13217);
or U18250 (N_18250,N_14079,N_14589);
and U18251 (N_18251,N_12014,N_14386);
and U18252 (N_18252,N_14687,N_13837);
nand U18253 (N_18253,N_11377,N_14609);
nand U18254 (N_18254,N_14126,N_11150);
nor U18255 (N_18255,N_11333,N_13849);
nor U18256 (N_18256,N_13236,N_13056);
nand U18257 (N_18257,N_12156,N_14105);
and U18258 (N_18258,N_11110,N_14598);
and U18259 (N_18259,N_13840,N_11629);
or U18260 (N_18260,N_14008,N_11766);
and U18261 (N_18261,N_14835,N_11655);
or U18262 (N_18262,N_10865,N_12837);
and U18263 (N_18263,N_13891,N_10649);
or U18264 (N_18264,N_13596,N_13102);
or U18265 (N_18265,N_13271,N_13341);
nor U18266 (N_18266,N_12635,N_14792);
nor U18267 (N_18267,N_11738,N_14421);
nor U18268 (N_18268,N_11437,N_13890);
or U18269 (N_18269,N_13185,N_10687);
and U18270 (N_18270,N_10115,N_14213);
nor U18271 (N_18271,N_12345,N_11261);
nand U18272 (N_18272,N_14878,N_10799);
and U18273 (N_18273,N_14595,N_13718);
nor U18274 (N_18274,N_13349,N_11798);
nand U18275 (N_18275,N_13190,N_10718);
nand U18276 (N_18276,N_14684,N_11949);
nand U18277 (N_18277,N_13060,N_11350);
nand U18278 (N_18278,N_10746,N_12919);
nor U18279 (N_18279,N_10801,N_11660);
nand U18280 (N_18280,N_13926,N_14738);
nand U18281 (N_18281,N_10038,N_12958);
nor U18282 (N_18282,N_11182,N_13886);
nand U18283 (N_18283,N_11976,N_14455);
and U18284 (N_18284,N_11572,N_11521);
or U18285 (N_18285,N_11539,N_13849);
nor U18286 (N_18286,N_14033,N_14766);
nor U18287 (N_18287,N_11622,N_14381);
nor U18288 (N_18288,N_11398,N_11513);
and U18289 (N_18289,N_10997,N_12420);
nor U18290 (N_18290,N_10109,N_11366);
and U18291 (N_18291,N_14999,N_10896);
nor U18292 (N_18292,N_10390,N_11134);
nor U18293 (N_18293,N_14934,N_11041);
or U18294 (N_18294,N_12051,N_14035);
and U18295 (N_18295,N_14657,N_10139);
nor U18296 (N_18296,N_12061,N_14735);
nand U18297 (N_18297,N_13466,N_11527);
xor U18298 (N_18298,N_10317,N_14263);
and U18299 (N_18299,N_11204,N_13854);
xnor U18300 (N_18300,N_13959,N_10584);
and U18301 (N_18301,N_11391,N_13008);
and U18302 (N_18302,N_10994,N_12905);
or U18303 (N_18303,N_11212,N_11529);
or U18304 (N_18304,N_10659,N_13697);
nor U18305 (N_18305,N_13468,N_10347);
and U18306 (N_18306,N_11425,N_12037);
or U18307 (N_18307,N_11357,N_11187);
and U18308 (N_18308,N_14196,N_11520);
nor U18309 (N_18309,N_14171,N_10505);
nor U18310 (N_18310,N_11756,N_12560);
nor U18311 (N_18311,N_10419,N_10058);
nand U18312 (N_18312,N_13847,N_12287);
and U18313 (N_18313,N_10918,N_12177);
nand U18314 (N_18314,N_10212,N_10483);
or U18315 (N_18315,N_13545,N_14045);
nor U18316 (N_18316,N_10400,N_10523);
nand U18317 (N_18317,N_14982,N_12506);
nand U18318 (N_18318,N_12498,N_14618);
nand U18319 (N_18319,N_10914,N_14474);
nor U18320 (N_18320,N_13175,N_14755);
and U18321 (N_18321,N_12657,N_13130);
nor U18322 (N_18322,N_10830,N_10472);
nor U18323 (N_18323,N_11250,N_14221);
nor U18324 (N_18324,N_10193,N_10317);
or U18325 (N_18325,N_12904,N_13831);
nor U18326 (N_18326,N_13289,N_14479);
or U18327 (N_18327,N_14776,N_12476);
and U18328 (N_18328,N_12154,N_13108);
and U18329 (N_18329,N_11609,N_10487);
nor U18330 (N_18330,N_11490,N_11009);
or U18331 (N_18331,N_14875,N_11436);
and U18332 (N_18332,N_10065,N_10490);
and U18333 (N_18333,N_11060,N_13608);
nor U18334 (N_18334,N_12563,N_12462);
nor U18335 (N_18335,N_10698,N_11346);
or U18336 (N_18336,N_12897,N_11042);
and U18337 (N_18337,N_13494,N_14791);
nor U18338 (N_18338,N_11852,N_14521);
or U18339 (N_18339,N_13264,N_10127);
and U18340 (N_18340,N_10278,N_12828);
nand U18341 (N_18341,N_12923,N_12649);
or U18342 (N_18342,N_12780,N_13893);
nand U18343 (N_18343,N_12837,N_14491);
and U18344 (N_18344,N_11050,N_12391);
and U18345 (N_18345,N_11193,N_13755);
and U18346 (N_18346,N_13771,N_10871);
or U18347 (N_18347,N_13778,N_10664);
nand U18348 (N_18348,N_13729,N_13199);
nor U18349 (N_18349,N_13511,N_12118);
and U18350 (N_18350,N_12936,N_10717);
nand U18351 (N_18351,N_12155,N_10036);
and U18352 (N_18352,N_14129,N_13259);
nor U18353 (N_18353,N_11794,N_13028);
nor U18354 (N_18354,N_10882,N_11588);
or U18355 (N_18355,N_13759,N_11799);
nor U18356 (N_18356,N_11078,N_11041);
or U18357 (N_18357,N_14443,N_13240);
or U18358 (N_18358,N_14458,N_10660);
and U18359 (N_18359,N_14204,N_13699);
nand U18360 (N_18360,N_14429,N_12278);
nand U18361 (N_18361,N_14933,N_10200);
nand U18362 (N_18362,N_10505,N_10559);
nor U18363 (N_18363,N_12646,N_10814);
nand U18364 (N_18364,N_11976,N_11739);
and U18365 (N_18365,N_14238,N_11863);
nand U18366 (N_18366,N_14674,N_13844);
and U18367 (N_18367,N_14013,N_14668);
and U18368 (N_18368,N_11598,N_10710);
and U18369 (N_18369,N_13118,N_12070);
nor U18370 (N_18370,N_12057,N_12819);
nand U18371 (N_18371,N_10778,N_12661);
and U18372 (N_18372,N_14027,N_12316);
or U18373 (N_18373,N_11965,N_10979);
or U18374 (N_18374,N_12309,N_13190);
nand U18375 (N_18375,N_14048,N_10544);
nor U18376 (N_18376,N_13016,N_14854);
nor U18377 (N_18377,N_12028,N_11435);
nor U18378 (N_18378,N_13700,N_13139);
nor U18379 (N_18379,N_11832,N_12887);
and U18380 (N_18380,N_11116,N_12218);
nor U18381 (N_18381,N_10617,N_12120);
nor U18382 (N_18382,N_11066,N_12791);
and U18383 (N_18383,N_10946,N_14687);
nor U18384 (N_18384,N_14811,N_10366);
nand U18385 (N_18385,N_12324,N_10476);
nand U18386 (N_18386,N_14724,N_10772);
nor U18387 (N_18387,N_12872,N_10569);
and U18388 (N_18388,N_12023,N_14626);
or U18389 (N_18389,N_11124,N_13984);
or U18390 (N_18390,N_10372,N_14769);
or U18391 (N_18391,N_14239,N_12792);
and U18392 (N_18392,N_13514,N_14778);
nor U18393 (N_18393,N_11998,N_13318);
and U18394 (N_18394,N_10552,N_13043);
and U18395 (N_18395,N_13538,N_11360);
nor U18396 (N_18396,N_13700,N_11902);
or U18397 (N_18397,N_10959,N_10870);
nor U18398 (N_18398,N_10002,N_12295);
nor U18399 (N_18399,N_11824,N_14778);
and U18400 (N_18400,N_12498,N_11402);
nor U18401 (N_18401,N_11448,N_12291);
and U18402 (N_18402,N_11484,N_11050);
nand U18403 (N_18403,N_11064,N_14983);
nand U18404 (N_18404,N_13015,N_14109);
nand U18405 (N_18405,N_11018,N_11021);
nor U18406 (N_18406,N_11199,N_11269);
nor U18407 (N_18407,N_10267,N_14815);
nand U18408 (N_18408,N_14692,N_12020);
or U18409 (N_18409,N_11725,N_10224);
and U18410 (N_18410,N_13036,N_11826);
or U18411 (N_18411,N_13506,N_10645);
nand U18412 (N_18412,N_11693,N_13890);
nor U18413 (N_18413,N_10725,N_14899);
nand U18414 (N_18414,N_13637,N_14200);
or U18415 (N_18415,N_12193,N_13463);
and U18416 (N_18416,N_13736,N_11438);
nand U18417 (N_18417,N_14723,N_11810);
and U18418 (N_18418,N_12738,N_14938);
and U18419 (N_18419,N_11424,N_14710);
and U18420 (N_18420,N_14848,N_11010);
nand U18421 (N_18421,N_12240,N_13471);
nand U18422 (N_18422,N_12558,N_10356);
or U18423 (N_18423,N_10857,N_12966);
nor U18424 (N_18424,N_12270,N_12533);
nand U18425 (N_18425,N_13213,N_13539);
or U18426 (N_18426,N_14512,N_14696);
and U18427 (N_18427,N_11399,N_12818);
nand U18428 (N_18428,N_14111,N_14836);
or U18429 (N_18429,N_12277,N_14055);
nor U18430 (N_18430,N_13726,N_14257);
and U18431 (N_18431,N_13806,N_13546);
or U18432 (N_18432,N_10060,N_14258);
xor U18433 (N_18433,N_14703,N_13326);
or U18434 (N_18434,N_10123,N_14074);
or U18435 (N_18435,N_13487,N_10965);
nand U18436 (N_18436,N_12216,N_11147);
and U18437 (N_18437,N_14896,N_13851);
or U18438 (N_18438,N_13601,N_14293);
nand U18439 (N_18439,N_13321,N_12592);
or U18440 (N_18440,N_13560,N_12523);
nor U18441 (N_18441,N_13434,N_14958);
and U18442 (N_18442,N_11533,N_14923);
nor U18443 (N_18443,N_10854,N_10204);
or U18444 (N_18444,N_11537,N_10050);
and U18445 (N_18445,N_12216,N_13393);
nand U18446 (N_18446,N_11471,N_13889);
nand U18447 (N_18447,N_12772,N_10566);
nor U18448 (N_18448,N_12094,N_12297);
and U18449 (N_18449,N_14653,N_12289);
nand U18450 (N_18450,N_11256,N_14957);
and U18451 (N_18451,N_12419,N_11822);
and U18452 (N_18452,N_11884,N_14094);
nand U18453 (N_18453,N_12351,N_12029);
and U18454 (N_18454,N_14983,N_11113);
or U18455 (N_18455,N_10568,N_13093);
or U18456 (N_18456,N_10943,N_12615);
and U18457 (N_18457,N_14369,N_12496);
nand U18458 (N_18458,N_13275,N_11031);
and U18459 (N_18459,N_10611,N_10977);
nor U18460 (N_18460,N_10496,N_14385);
nor U18461 (N_18461,N_11552,N_11463);
nand U18462 (N_18462,N_12795,N_14975);
nand U18463 (N_18463,N_13227,N_11669);
and U18464 (N_18464,N_12892,N_11827);
nand U18465 (N_18465,N_11355,N_11674);
or U18466 (N_18466,N_14498,N_13128);
and U18467 (N_18467,N_13981,N_11681);
nor U18468 (N_18468,N_12734,N_12575);
xnor U18469 (N_18469,N_10235,N_14590);
nand U18470 (N_18470,N_14548,N_10996);
or U18471 (N_18471,N_14172,N_14696);
nor U18472 (N_18472,N_10202,N_10634);
xnor U18473 (N_18473,N_13509,N_10816);
or U18474 (N_18474,N_13061,N_12792);
or U18475 (N_18475,N_13652,N_14702);
and U18476 (N_18476,N_14670,N_11615);
nor U18477 (N_18477,N_14944,N_14545);
and U18478 (N_18478,N_12360,N_13947);
or U18479 (N_18479,N_10387,N_10836);
nand U18480 (N_18480,N_12457,N_12195);
or U18481 (N_18481,N_13874,N_11462);
and U18482 (N_18482,N_14240,N_12537);
nor U18483 (N_18483,N_10797,N_14646);
nor U18484 (N_18484,N_14110,N_12970);
nor U18485 (N_18485,N_13475,N_14496);
nor U18486 (N_18486,N_12949,N_14447);
and U18487 (N_18487,N_14148,N_14546);
or U18488 (N_18488,N_11069,N_12658);
nand U18489 (N_18489,N_11450,N_13459);
and U18490 (N_18490,N_13942,N_11172);
or U18491 (N_18491,N_13288,N_14152);
nor U18492 (N_18492,N_10509,N_10761);
and U18493 (N_18493,N_11967,N_14029);
and U18494 (N_18494,N_14244,N_12971);
and U18495 (N_18495,N_13849,N_11186);
and U18496 (N_18496,N_14684,N_10232);
nand U18497 (N_18497,N_11800,N_11492);
nand U18498 (N_18498,N_13767,N_11558);
and U18499 (N_18499,N_12083,N_11600);
nand U18500 (N_18500,N_11220,N_14260);
or U18501 (N_18501,N_10629,N_10592);
nand U18502 (N_18502,N_11346,N_14022);
nand U18503 (N_18503,N_12878,N_14357);
and U18504 (N_18504,N_13475,N_13111);
nor U18505 (N_18505,N_12114,N_14299);
nor U18506 (N_18506,N_11161,N_13236);
and U18507 (N_18507,N_11913,N_12081);
or U18508 (N_18508,N_12168,N_13534);
nor U18509 (N_18509,N_14346,N_13363);
nand U18510 (N_18510,N_14842,N_12897);
and U18511 (N_18511,N_10029,N_13222);
and U18512 (N_18512,N_12286,N_13446);
and U18513 (N_18513,N_14845,N_10012);
nor U18514 (N_18514,N_11390,N_14106);
or U18515 (N_18515,N_11279,N_10378);
nand U18516 (N_18516,N_14454,N_12766);
nor U18517 (N_18517,N_10392,N_10277);
and U18518 (N_18518,N_14896,N_11796);
or U18519 (N_18519,N_11913,N_12805);
nor U18520 (N_18520,N_10966,N_14007);
nor U18521 (N_18521,N_11940,N_11055);
nor U18522 (N_18522,N_11151,N_10253);
or U18523 (N_18523,N_10907,N_14540);
or U18524 (N_18524,N_10682,N_11284);
or U18525 (N_18525,N_10276,N_11529);
or U18526 (N_18526,N_13603,N_10089);
nand U18527 (N_18527,N_11808,N_13750);
nand U18528 (N_18528,N_14375,N_12534);
or U18529 (N_18529,N_14722,N_13047);
nor U18530 (N_18530,N_10001,N_10562);
and U18531 (N_18531,N_13870,N_12248);
nor U18532 (N_18532,N_14128,N_12794);
or U18533 (N_18533,N_11919,N_13368);
nor U18534 (N_18534,N_12738,N_14476);
nand U18535 (N_18535,N_13711,N_12026);
and U18536 (N_18536,N_10636,N_13568);
or U18537 (N_18537,N_12875,N_10324);
xor U18538 (N_18538,N_12120,N_13514);
and U18539 (N_18539,N_12355,N_12455);
nand U18540 (N_18540,N_12307,N_12087);
nand U18541 (N_18541,N_12395,N_10840);
nor U18542 (N_18542,N_13987,N_14751);
or U18543 (N_18543,N_14622,N_14661);
nor U18544 (N_18544,N_13897,N_12209);
or U18545 (N_18545,N_14248,N_10042);
nand U18546 (N_18546,N_12717,N_12869);
or U18547 (N_18547,N_10843,N_12193);
nand U18548 (N_18548,N_14368,N_12119);
and U18549 (N_18549,N_13390,N_12059);
nor U18550 (N_18550,N_10642,N_11246);
or U18551 (N_18551,N_11541,N_14452);
and U18552 (N_18552,N_10967,N_11773);
nor U18553 (N_18553,N_13794,N_14974);
nor U18554 (N_18554,N_14887,N_13084);
and U18555 (N_18555,N_12585,N_14282);
nor U18556 (N_18556,N_12850,N_11455);
and U18557 (N_18557,N_13445,N_14498);
or U18558 (N_18558,N_14530,N_14127);
nand U18559 (N_18559,N_13020,N_10123);
nand U18560 (N_18560,N_13784,N_11837);
or U18561 (N_18561,N_14172,N_14936);
nor U18562 (N_18562,N_12623,N_13545);
and U18563 (N_18563,N_10106,N_11139);
and U18564 (N_18564,N_12563,N_12409);
nor U18565 (N_18565,N_11629,N_14267);
or U18566 (N_18566,N_14413,N_11731);
or U18567 (N_18567,N_13679,N_13058);
nand U18568 (N_18568,N_13731,N_14174);
nor U18569 (N_18569,N_12325,N_10519);
and U18570 (N_18570,N_14973,N_14717);
nand U18571 (N_18571,N_10770,N_13759);
nor U18572 (N_18572,N_10310,N_10851);
or U18573 (N_18573,N_14587,N_13243);
or U18574 (N_18574,N_10025,N_10574);
nand U18575 (N_18575,N_12554,N_12858);
nor U18576 (N_18576,N_11979,N_10912);
or U18577 (N_18577,N_10979,N_13566);
and U18578 (N_18578,N_12533,N_14087);
and U18579 (N_18579,N_13052,N_11029);
or U18580 (N_18580,N_10002,N_14115);
and U18581 (N_18581,N_10957,N_10701);
or U18582 (N_18582,N_12138,N_13645);
or U18583 (N_18583,N_13817,N_11441);
or U18584 (N_18584,N_10422,N_10165);
nand U18585 (N_18585,N_14933,N_12946);
xor U18586 (N_18586,N_10778,N_10976);
nand U18587 (N_18587,N_10042,N_11437);
nor U18588 (N_18588,N_10407,N_14518);
and U18589 (N_18589,N_10078,N_11236);
or U18590 (N_18590,N_13473,N_10930);
nor U18591 (N_18591,N_13431,N_12169);
nand U18592 (N_18592,N_13352,N_11815);
and U18593 (N_18593,N_13631,N_10444);
nand U18594 (N_18594,N_14251,N_10947);
or U18595 (N_18595,N_13908,N_13354);
nor U18596 (N_18596,N_12215,N_13336);
nor U18597 (N_18597,N_11593,N_14978);
or U18598 (N_18598,N_14176,N_11623);
or U18599 (N_18599,N_13200,N_11374);
nor U18600 (N_18600,N_13923,N_14315);
nand U18601 (N_18601,N_12327,N_14841);
or U18602 (N_18602,N_10466,N_12983);
and U18603 (N_18603,N_11254,N_13659);
and U18604 (N_18604,N_12682,N_12257);
nand U18605 (N_18605,N_11801,N_11521);
or U18606 (N_18606,N_14598,N_10597);
or U18607 (N_18607,N_13737,N_10797);
nand U18608 (N_18608,N_12147,N_13540);
nor U18609 (N_18609,N_12695,N_10640);
and U18610 (N_18610,N_12860,N_12461);
or U18611 (N_18611,N_11428,N_10809);
nand U18612 (N_18612,N_11904,N_11879);
or U18613 (N_18613,N_11650,N_13166);
or U18614 (N_18614,N_11121,N_13727);
or U18615 (N_18615,N_13135,N_12261);
nand U18616 (N_18616,N_11763,N_11088);
nor U18617 (N_18617,N_13995,N_10154);
or U18618 (N_18618,N_12852,N_13377);
nor U18619 (N_18619,N_10470,N_13068);
and U18620 (N_18620,N_14758,N_12661);
or U18621 (N_18621,N_12197,N_12388);
and U18622 (N_18622,N_10925,N_13754);
nand U18623 (N_18623,N_10637,N_11092);
or U18624 (N_18624,N_14351,N_10045);
nand U18625 (N_18625,N_12931,N_10483);
or U18626 (N_18626,N_10938,N_12132);
nand U18627 (N_18627,N_13119,N_13827);
or U18628 (N_18628,N_13789,N_10862);
and U18629 (N_18629,N_12182,N_12765);
and U18630 (N_18630,N_10049,N_13812);
and U18631 (N_18631,N_10946,N_14165);
nand U18632 (N_18632,N_11610,N_11491);
nand U18633 (N_18633,N_12722,N_11819);
nand U18634 (N_18634,N_10959,N_12618);
and U18635 (N_18635,N_10865,N_14283);
nand U18636 (N_18636,N_14207,N_13127);
or U18637 (N_18637,N_10117,N_12110);
nand U18638 (N_18638,N_10259,N_11552);
nor U18639 (N_18639,N_12757,N_13083);
or U18640 (N_18640,N_11540,N_11262);
and U18641 (N_18641,N_14303,N_11980);
nor U18642 (N_18642,N_10768,N_13508);
nand U18643 (N_18643,N_11378,N_11716);
or U18644 (N_18644,N_13382,N_11582);
nand U18645 (N_18645,N_11164,N_11589);
and U18646 (N_18646,N_11860,N_11106);
nor U18647 (N_18647,N_10385,N_11904);
or U18648 (N_18648,N_12057,N_14648);
nand U18649 (N_18649,N_11337,N_12650);
and U18650 (N_18650,N_11542,N_14690);
and U18651 (N_18651,N_10131,N_10326);
or U18652 (N_18652,N_14261,N_11336);
nand U18653 (N_18653,N_13622,N_14645);
nor U18654 (N_18654,N_13876,N_12359);
nor U18655 (N_18655,N_11255,N_11129);
nor U18656 (N_18656,N_12340,N_10287);
nor U18657 (N_18657,N_12186,N_13523);
or U18658 (N_18658,N_14019,N_13100);
and U18659 (N_18659,N_10397,N_10079);
nor U18660 (N_18660,N_13070,N_11432);
nor U18661 (N_18661,N_12651,N_11235);
and U18662 (N_18662,N_13448,N_13500);
and U18663 (N_18663,N_12674,N_10550);
or U18664 (N_18664,N_10044,N_14376);
or U18665 (N_18665,N_14597,N_11878);
nor U18666 (N_18666,N_14871,N_10086);
or U18667 (N_18667,N_13480,N_12565);
nor U18668 (N_18668,N_12583,N_14096);
and U18669 (N_18669,N_10931,N_13919);
nor U18670 (N_18670,N_13661,N_13302);
and U18671 (N_18671,N_11635,N_14982);
nor U18672 (N_18672,N_10247,N_13529);
and U18673 (N_18673,N_11284,N_12614);
nor U18674 (N_18674,N_12637,N_11071);
and U18675 (N_18675,N_10555,N_11023);
or U18676 (N_18676,N_10689,N_13471);
and U18677 (N_18677,N_10086,N_13902);
or U18678 (N_18678,N_11899,N_13910);
or U18679 (N_18679,N_12508,N_11031);
or U18680 (N_18680,N_12135,N_13794);
nor U18681 (N_18681,N_13035,N_13346);
and U18682 (N_18682,N_12146,N_14640);
and U18683 (N_18683,N_14250,N_12739);
nand U18684 (N_18684,N_11991,N_11360);
or U18685 (N_18685,N_13647,N_11491);
nor U18686 (N_18686,N_12810,N_10514);
and U18687 (N_18687,N_11299,N_11304);
nand U18688 (N_18688,N_12578,N_12330);
and U18689 (N_18689,N_14314,N_10136);
nand U18690 (N_18690,N_12124,N_12074);
nand U18691 (N_18691,N_11891,N_13710);
nor U18692 (N_18692,N_10978,N_10603);
nor U18693 (N_18693,N_11594,N_13946);
nand U18694 (N_18694,N_13086,N_11421);
nor U18695 (N_18695,N_12427,N_14115);
or U18696 (N_18696,N_14266,N_11975);
nor U18697 (N_18697,N_11733,N_11250);
nand U18698 (N_18698,N_12245,N_11126);
nor U18699 (N_18699,N_11433,N_11410);
nor U18700 (N_18700,N_13123,N_14256);
nand U18701 (N_18701,N_14793,N_13736);
and U18702 (N_18702,N_10356,N_10071);
nand U18703 (N_18703,N_12256,N_10565);
or U18704 (N_18704,N_13286,N_11247);
nor U18705 (N_18705,N_12623,N_11666);
nand U18706 (N_18706,N_14223,N_11133);
or U18707 (N_18707,N_13708,N_13025);
nand U18708 (N_18708,N_13177,N_12752);
or U18709 (N_18709,N_12596,N_14918);
and U18710 (N_18710,N_11794,N_12129);
and U18711 (N_18711,N_13850,N_10790);
nand U18712 (N_18712,N_14005,N_14748);
nor U18713 (N_18713,N_12829,N_12836);
xor U18714 (N_18714,N_12355,N_13156);
nand U18715 (N_18715,N_14756,N_11905);
or U18716 (N_18716,N_13631,N_10322);
nor U18717 (N_18717,N_14641,N_11284);
or U18718 (N_18718,N_13497,N_14552);
nor U18719 (N_18719,N_14507,N_10138);
nor U18720 (N_18720,N_14445,N_14118);
and U18721 (N_18721,N_10379,N_13562);
nor U18722 (N_18722,N_11142,N_10396);
nor U18723 (N_18723,N_12872,N_13348);
nor U18724 (N_18724,N_11308,N_12465);
or U18725 (N_18725,N_13677,N_12453);
nor U18726 (N_18726,N_11174,N_12332);
nand U18727 (N_18727,N_14848,N_11444);
and U18728 (N_18728,N_14388,N_13762);
and U18729 (N_18729,N_11176,N_13738);
nor U18730 (N_18730,N_12716,N_10311);
nand U18731 (N_18731,N_12459,N_12895);
and U18732 (N_18732,N_10518,N_13266);
or U18733 (N_18733,N_10036,N_11290);
and U18734 (N_18734,N_11184,N_14379);
nor U18735 (N_18735,N_10589,N_13971);
or U18736 (N_18736,N_10914,N_14530);
nand U18737 (N_18737,N_13254,N_13156);
nor U18738 (N_18738,N_12713,N_11659);
nor U18739 (N_18739,N_12109,N_12080);
nand U18740 (N_18740,N_12096,N_10651);
nor U18741 (N_18741,N_14176,N_11317);
and U18742 (N_18742,N_13650,N_11818);
nand U18743 (N_18743,N_13470,N_11804);
nand U18744 (N_18744,N_13531,N_12128);
and U18745 (N_18745,N_12824,N_10055);
and U18746 (N_18746,N_10886,N_13422);
or U18747 (N_18747,N_12916,N_13618);
nand U18748 (N_18748,N_11071,N_12015);
nor U18749 (N_18749,N_10679,N_11470);
and U18750 (N_18750,N_14397,N_14459);
or U18751 (N_18751,N_12120,N_12171);
and U18752 (N_18752,N_11154,N_12318);
xor U18753 (N_18753,N_10721,N_11184);
nor U18754 (N_18754,N_14416,N_12870);
nor U18755 (N_18755,N_11874,N_13271);
nor U18756 (N_18756,N_12027,N_14834);
or U18757 (N_18757,N_11802,N_11605);
nand U18758 (N_18758,N_10275,N_14615);
nand U18759 (N_18759,N_14318,N_14279);
and U18760 (N_18760,N_13274,N_10993);
nand U18761 (N_18761,N_14986,N_10640);
and U18762 (N_18762,N_12732,N_10509);
nand U18763 (N_18763,N_14312,N_13392);
nor U18764 (N_18764,N_10647,N_13385);
nand U18765 (N_18765,N_12190,N_12760);
and U18766 (N_18766,N_12210,N_12296);
or U18767 (N_18767,N_14862,N_12839);
nand U18768 (N_18768,N_12407,N_13005);
and U18769 (N_18769,N_12219,N_11696);
nor U18770 (N_18770,N_12359,N_12496);
nor U18771 (N_18771,N_11950,N_14389);
nor U18772 (N_18772,N_12779,N_11689);
and U18773 (N_18773,N_13085,N_10496);
or U18774 (N_18774,N_13849,N_13573);
and U18775 (N_18775,N_11996,N_10842);
or U18776 (N_18776,N_12405,N_12809);
nor U18777 (N_18777,N_11580,N_14819);
nand U18778 (N_18778,N_11263,N_10345);
nor U18779 (N_18779,N_10047,N_14636);
nor U18780 (N_18780,N_11124,N_12659);
nand U18781 (N_18781,N_13671,N_10855);
and U18782 (N_18782,N_11136,N_13608);
and U18783 (N_18783,N_14301,N_11217);
and U18784 (N_18784,N_13786,N_12623);
or U18785 (N_18785,N_12430,N_10250);
nand U18786 (N_18786,N_13334,N_11228);
or U18787 (N_18787,N_10155,N_12330);
nor U18788 (N_18788,N_12097,N_10262);
nor U18789 (N_18789,N_10357,N_13357);
nor U18790 (N_18790,N_12845,N_12208);
nor U18791 (N_18791,N_13629,N_10691);
and U18792 (N_18792,N_12233,N_11232);
nand U18793 (N_18793,N_13271,N_14807);
nor U18794 (N_18794,N_10364,N_13971);
or U18795 (N_18795,N_14336,N_10510);
and U18796 (N_18796,N_12118,N_14164);
or U18797 (N_18797,N_12215,N_12845);
and U18798 (N_18798,N_14858,N_14578);
nand U18799 (N_18799,N_12046,N_12832);
or U18800 (N_18800,N_10914,N_12455);
and U18801 (N_18801,N_14132,N_13248);
nand U18802 (N_18802,N_11301,N_10169);
or U18803 (N_18803,N_11033,N_11146);
and U18804 (N_18804,N_10610,N_14277);
nand U18805 (N_18805,N_10540,N_11661);
nand U18806 (N_18806,N_11344,N_10394);
or U18807 (N_18807,N_14647,N_12571);
nand U18808 (N_18808,N_11661,N_12173);
nand U18809 (N_18809,N_11693,N_12228);
and U18810 (N_18810,N_12537,N_12703);
and U18811 (N_18811,N_14643,N_10192);
or U18812 (N_18812,N_13683,N_12123);
and U18813 (N_18813,N_10312,N_14356);
nand U18814 (N_18814,N_13304,N_10976);
and U18815 (N_18815,N_12929,N_10099);
or U18816 (N_18816,N_10592,N_13583);
nor U18817 (N_18817,N_14000,N_14904);
and U18818 (N_18818,N_10795,N_11090);
nor U18819 (N_18819,N_14977,N_12450);
or U18820 (N_18820,N_13509,N_11660);
nand U18821 (N_18821,N_13691,N_12555);
nor U18822 (N_18822,N_13187,N_13293);
and U18823 (N_18823,N_12013,N_13124);
or U18824 (N_18824,N_13639,N_11291);
and U18825 (N_18825,N_12571,N_12680);
nor U18826 (N_18826,N_13203,N_10159);
or U18827 (N_18827,N_13442,N_11379);
and U18828 (N_18828,N_12287,N_13424);
and U18829 (N_18829,N_13213,N_13664);
nor U18830 (N_18830,N_14766,N_13553);
or U18831 (N_18831,N_12006,N_12995);
nor U18832 (N_18832,N_12623,N_13145);
or U18833 (N_18833,N_10313,N_11456);
nand U18834 (N_18834,N_10236,N_12122);
nor U18835 (N_18835,N_10942,N_10152);
nand U18836 (N_18836,N_12498,N_12683);
nor U18837 (N_18837,N_14198,N_13887);
nor U18838 (N_18838,N_12893,N_13294);
or U18839 (N_18839,N_14199,N_12697);
nand U18840 (N_18840,N_10124,N_14789);
nand U18841 (N_18841,N_11003,N_10289);
or U18842 (N_18842,N_11168,N_10032);
nor U18843 (N_18843,N_14092,N_14337);
and U18844 (N_18844,N_11595,N_13642);
and U18845 (N_18845,N_13739,N_11184);
and U18846 (N_18846,N_11333,N_13489);
or U18847 (N_18847,N_13431,N_14352);
nor U18848 (N_18848,N_12487,N_13243);
nand U18849 (N_18849,N_12610,N_12733);
nor U18850 (N_18850,N_14884,N_12704);
nor U18851 (N_18851,N_10466,N_14060);
nor U18852 (N_18852,N_14596,N_10317);
and U18853 (N_18853,N_13410,N_14227);
nor U18854 (N_18854,N_13147,N_14503);
or U18855 (N_18855,N_13049,N_13232);
nand U18856 (N_18856,N_14534,N_14076);
and U18857 (N_18857,N_10134,N_12435);
nor U18858 (N_18858,N_10226,N_14758);
and U18859 (N_18859,N_12322,N_13783);
nand U18860 (N_18860,N_14807,N_14957);
nand U18861 (N_18861,N_11207,N_11748);
and U18862 (N_18862,N_12979,N_12612);
or U18863 (N_18863,N_11453,N_10155);
nor U18864 (N_18864,N_13120,N_10033);
or U18865 (N_18865,N_12163,N_11723);
nand U18866 (N_18866,N_14633,N_14765);
nor U18867 (N_18867,N_11844,N_14917);
nor U18868 (N_18868,N_10450,N_12897);
nor U18869 (N_18869,N_14925,N_10281);
or U18870 (N_18870,N_12500,N_14673);
nand U18871 (N_18871,N_14283,N_10256);
or U18872 (N_18872,N_14838,N_13947);
or U18873 (N_18873,N_10085,N_11582);
nand U18874 (N_18874,N_13087,N_13758);
and U18875 (N_18875,N_10441,N_11619);
nand U18876 (N_18876,N_13873,N_14454);
and U18877 (N_18877,N_14588,N_12875);
nor U18878 (N_18878,N_12193,N_13895);
and U18879 (N_18879,N_14049,N_14347);
nor U18880 (N_18880,N_11105,N_13866);
nor U18881 (N_18881,N_11398,N_12952);
and U18882 (N_18882,N_14638,N_12784);
nor U18883 (N_18883,N_11910,N_10382);
nor U18884 (N_18884,N_12332,N_14798);
or U18885 (N_18885,N_14899,N_13279);
nor U18886 (N_18886,N_10261,N_13092);
or U18887 (N_18887,N_12139,N_10778);
nand U18888 (N_18888,N_11403,N_11682);
and U18889 (N_18889,N_14416,N_10424);
or U18890 (N_18890,N_11234,N_12179);
nand U18891 (N_18891,N_11773,N_12513);
nor U18892 (N_18892,N_14926,N_10887);
nand U18893 (N_18893,N_13481,N_10547);
and U18894 (N_18894,N_14475,N_11072);
nand U18895 (N_18895,N_14363,N_13193);
nor U18896 (N_18896,N_13801,N_12917);
xnor U18897 (N_18897,N_11700,N_14667);
and U18898 (N_18898,N_13737,N_14051);
nand U18899 (N_18899,N_10689,N_12753);
and U18900 (N_18900,N_12811,N_12104);
or U18901 (N_18901,N_14313,N_11190);
and U18902 (N_18902,N_12444,N_10044);
and U18903 (N_18903,N_13632,N_14963);
nor U18904 (N_18904,N_10042,N_12540);
nand U18905 (N_18905,N_13232,N_11385);
nor U18906 (N_18906,N_11015,N_13943);
nand U18907 (N_18907,N_13616,N_14388);
nor U18908 (N_18908,N_10910,N_14990);
nor U18909 (N_18909,N_14087,N_14487);
nor U18910 (N_18910,N_10116,N_14624);
or U18911 (N_18911,N_12104,N_13796);
and U18912 (N_18912,N_10893,N_13181);
or U18913 (N_18913,N_10726,N_10384);
or U18914 (N_18914,N_11993,N_10306);
nand U18915 (N_18915,N_12576,N_12802);
or U18916 (N_18916,N_12201,N_10493);
and U18917 (N_18917,N_12928,N_13109);
nor U18918 (N_18918,N_14025,N_12965);
nor U18919 (N_18919,N_10391,N_10507);
or U18920 (N_18920,N_13681,N_14640);
or U18921 (N_18921,N_13074,N_14927);
nor U18922 (N_18922,N_12687,N_14489);
or U18923 (N_18923,N_12524,N_12531);
or U18924 (N_18924,N_12588,N_10957);
and U18925 (N_18925,N_14460,N_12109);
nor U18926 (N_18926,N_12154,N_12095);
xnor U18927 (N_18927,N_11157,N_13350);
and U18928 (N_18928,N_10316,N_12408);
nor U18929 (N_18929,N_11147,N_14397);
nand U18930 (N_18930,N_13191,N_11025);
or U18931 (N_18931,N_14822,N_11581);
nor U18932 (N_18932,N_14545,N_12408);
nand U18933 (N_18933,N_12846,N_14343);
or U18934 (N_18934,N_11631,N_13461);
xnor U18935 (N_18935,N_11563,N_12104);
nor U18936 (N_18936,N_11782,N_11766);
nor U18937 (N_18937,N_13019,N_12276);
nand U18938 (N_18938,N_13475,N_13447);
or U18939 (N_18939,N_13132,N_11212);
nor U18940 (N_18940,N_14424,N_14958);
nand U18941 (N_18941,N_12944,N_10867);
or U18942 (N_18942,N_13094,N_13463);
and U18943 (N_18943,N_11840,N_12667);
nand U18944 (N_18944,N_13555,N_12887);
nor U18945 (N_18945,N_11983,N_12220);
nor U18946 (N_18946,N_10928,N_12090);
or U18947 (N_18947,N_14214,N_13012);
nand U18948 (N_18948,N_12288,N_10525);
nor U18949 (N_18949,N_12704,N_10387);
nor U18950 (N_18950,N_10532,N_10252);
or U18951 (N_18951,N_14785,N_10892);
or U18952 (N_18952,N_11228,N_14104);
nor U18953 (N_18953,N_11376,N_11133);
and U18954 (N_18954,N_12745,N_11127);
nand U18955 (N_18955,N_13817,N_10084);
nand U18956 (N_18956,N_10764,N_10399);
nor U18957 (N_18957,N_12978,N_14423);
nor U18958 (N_18958,N_13236,N_11337);
or U18959 (N_18959,N_13125,N_14190);
or U18960 (N_18960,N_12031,N_13720);
nand U18961 (N_18961,N_11350,N_13580);
and U18962 (N_18962,N_13007,N_10480);
nand U18963 (N_18963,N_13048,N_14066);
nand U18964 (N_18964,N_10238,N_10300);
and U18965 (N_18965,N_10015,N_10969);
and U18966 (N_18966,N_14905,N_14369);
nor U18967 (N_18967,N_10926,N_10818);
xor U18968 (N_18968,N_11704,N_12471);
nand U18969 (N_18969,N_11992,N_12628);
and U18970 (N_18970,N_10334,N_10015);
nand U18971 (N_18971,N_10262,N_14017);
and U18972 (N_18972,N_11759,N_13218);
and U18973 (N_18973,N_10400,N_14522);
nand U18974 (N_18974,N_14524,N_11166);
nand U18975 (N_18975,N_10886,N_10507);
nor U18976 (N_18976,N_10091,N_14736);
or U18977 (N_18977,N_10594,N_12130);
nand U18978 (N_18978,N_10443,N_12729);
nor U18979 (N_18979,N_11635,N_10305);
nor U18980 (N_18980,N_11428,N_13198);
nand U18981 (N_18981,N_14365,N_13884);
nand U18982 (N_18982,N_10284,N_13080);
xor U18983 (N_18983,N_10991,N_12072);
or U18984 (N_18984,N_11055,N_14021);
or U18985 (N_18985,N_13586,N_13182);
nand U18986 (N_18986,N_14074,N_12032);
or U18987 (N_18987,N_12652,N_14668);
or U18988 (N_18988,N_14106,N_12958);
or U18989 (N_18989,N_10559,N_13041);
nor U18990 (N_18990,N_10215,N_11935);
and U18991 (N_18991,N_13791,N_13394);
nand U18992 (N_18992,N_12393,N_10269);
and U18993 (N_18993,N_14317,N_11884);
or U18994 (N_18994,N_11410,N_14180);
or U18995 (N_18995,N_14281,N_13531);
nor U18996 (N_18996,N_13516,N_10918);
nand U18997 (N_18997,N_10152,N_12101);
nor U18998 (N_18998,N_12922,N_10934);
or U18999 (N_18999,N_14756,N_13347);
and U19000 (N_19000,N_14539,N_11502);
nand U19001 (N_19001,N_14857,N_13743);
and U19002 (N_19002,N_11172,N_14720);
or U19003 (N_19003,N_13028,N_12705);
nand U19004 (N_19004,N_11705,N_10609);
nand U19005 (N_19005,N_10851,N_11297);
and U19006 (N_19006,N_11003,N_14425);
and U19007 (N_19007,N_12564,N_12843);
nor U19008 (N_19008,N_12319,N_13205);
and U19009 (N_19009,N_11363,N_13554);
and U19010 (N_19010,N_11057,N_11428);
and U19011 (N_19011,N_13717,N_14509);
or U19012 (N_19012,N_10048,N_12361);
nand U19013 (N_19013,N_10227,N_11767);
and U19014 (N_19014,N_12003,N_11160);
and U19015 (N_19015,N_10600,N_12861);
nand U19016 (N_19016,N_13258,N_11057);
or U19017 (N_19017,N_13931,N_14700);
nand U19018 (N_19018,N_13169,N_10505);
xnor U19019 (N_19019,N_14883,N_14047);
nor U19020 (N_19020,N_14563,N_12667);
or U19021 (N_19021,N_10031,N_10966);
nor U19022 (N_19022,N_12896,N_12238);
or U19023 (N_19023,N_11323,N_13989);
or U19024 (N_19024,N_10592,N_10234);
and U19025 (N_19025,N_10382,N_10338);
or U19026 (N_19026,N_13819,N_10524);
and U19027 (N_19027,N_10690,N_14083);
nor U19028 (N_19028,N_11368,N_13724);
nor U19029 (N_19029,N_12565,N_14000);
nand U19030 (N_19030,N_13087,N_10300);
and U19031 (N_19031,N_13864,N_13933);
and U19032 (N_19032,N_14816,N_13983);
nand U19033 (N_19033,N_13101,N_14920);
or U19034 (N_19034,N_13201,N_12806);
nor U19035 (N_19035,N_14414,N_13865);
or U19036 (N_19036,N_14771,N_12133);
and U19037 (N_19037,N_12987,N_12480);
or U19038 (N_19038,N_12944,N_12492);
or U19039 (N_19039,N_12663,N_14837);
nor U19040 (N_19040,N_12241,N_12113);
or U19041 (N_19041,N_11915,N_13738);
or U19042 (N_19042,N_12696,N_13619);
and U19043 (N_19043,N_13654,N_13420);
or U19044 (N_19044,N_10898,N_13899);
and U19045 (N_19045,N_12587,N_11773);
and U19046 (N_19046,N_11977,N_13968);
and U19047 (N_19047,N_13650,N_14174);
and U19048 (N_19048,N_12000,N_11341);
or U19049 (N_19049,N_12164,N_13699);
nand U19050 (N_19050,N_10810,N_11581);
nor U19051 (N_19051,N_12254,N_10904);
nor U19052 (N_19052,N_10559,N_12551);
and U19053 (N_19053,N_13589,N_14081);
and U19054 (N_19054,N_12799,N_13293);
nand U19055 (N_19055,N_14661,N_10114);
and U19056 (N_19056,N_10035,N_10730);
nand U19057 (N_19057,N_10464,N_12026);
and U19058 (N_19058,N_14182,N_11260);
nand U19059 (N_19059,N_14441,N_14037);
or U19060 (N_19060,N_12106,N_14137);
nor U19061 (N_19061,N_14124,N_13372);
nor U19062 (N_19062,N_13956,N_12142);
nand U19063 (N_19063,N_11980,N_10088);
nor U19064 (N_19064,N_11185,N_13583);
or U19065 (N_19065,N_10686,N_10774);
and U19066 (N_19066,N_14487,N_12582);
or U19067 (N_19067,N_12740,N_14066);
and U19068 (N_19068,N_13025,N_11737);
and U19069 (N_19069,N_10257,N_14254);
and U19070 (N_19070,N_13348,N_12589);
xnor U19071 (N_19071,N_11728,N_14032);
nor U19072 (N_19072,N_10240,N_14206);
or U19073 (N_19073,N_13380,N_11986);
nor U19074 (N_19074,N_12558,N_12970);
nor U19075 (N_19075,N_13246,N_13973);
nor U19076 (N_19076,N_13192,N_11027);
or U19077 (N_19077,N_11650,N_11445);
nor U19078 (N_19078,N_14216,N_13891);
and U19079 (N_19079,N_11604,N_12258);
nand U19080 (N_19080,N_10748,N_12794);
nor U19081 (N_19081,N_14893,N_13594);
nand U19082 (N_19082,N_13966,N_11266);
or U19083 (N_19083,N_12747,N_10408);
and U19084 (N_19084,N_10423,N_14178);
or U19085 (N_19085,N_13685,N_11523);
nand U19086 (N_19086,N_10348,N_10751);
and U19087 (N_19087,N_10542,N_10058);
and U19088 (N_19088,N_12886,N_12793);
nor U19089 (N_19089,N_14643,N_14425);
and U19090 (N_19090,N_11721,N_13208);
and U19091 (N_19091,N_14779,N_13493);
xnor U19092 (N_19092,N_11284,N_14705);
and U19093 (N_19093,N_14845,N_13069);
or U19094 (N_19094,N_14931,N_10655);
and U19095 (N_19095,N_12924,N_11340);
and U19096 (N_19096,N_12595,N_11943);
nor U19097 (N_19097,N_12212,N_10771);
nor U19098 (N_19098,N_13334,N_10745);
nor U19099 (N_19099,N_10330,N_11481);
or U19100 (N_19100,N_11325,N_14581);
nor U19101 (N_19101,N_13077,N_10580);
nand U19102 (N_19102,N_12784,N_10851);
nand U19103 (N_19103,N_14221,N_14283);
or U19104 (N_19104,N_10106,N_10814);
nor U19105 (N_19105,N_11662,N_11209);
nand U19106 (N_19106,N_14059,N_12572);
nand U19107 (N_19107,N_10970,N_13454);
nand U19108 (N_19108,N_13828,N_10222);
or U19109 (N_19109,N_11503,N_10161);
nor U19110 (N_19110,N_14684,N_12708);
nand U19111 (N_19111,N_13557,N_13365);
nor U19112 (N_19112,N_12998,N_14540);
or U19113 (N_19113,N_11417,N_14677);
nor U19114 (N_19114,N_12688,N_10809);
xnor U19115 (N_19115,N_10255,N_10693);
nand U19116 (N_19116,N_14707,N_10645);
or U19117 (N_19117,N_11211,N_12736);
nor U19118 (N_19118,N_12512,N_10835);
and U19119 (N_19119,N_14617,N_13312);
nor U19120 (N_19120,N_14228,N_12180);
and U19121 (N_19121,N_14108,N_10169);
nand U19122 (N_19122,N_10613,N_14653);
nor U19123 (N_19123,N_10860,N_14656);
and U19124 (N_19124,N_11901,N_13567);
or U19125 (N_19125,N_12798,N_14480);
nand U19126 (N_19126,N_12811,N_12199);
or U19127 (N_19127,N_10610,N_10523);
nand U19128 (N_19128,N_10131,N_10142);
and U19129 (N_19129,N_12444,N_10344);
nor U19130 (N_19130,N_14309,N_13022);
nor U19131 (N_19131,N_11693,N_13488);
and U19132 (N_19132,N_14043,N_12685);
nor U19133 (N_19133,N_11997,N_11047);
or U19134 (N_19134,N_11301,N_11564);
or U19135 (N_19135,N_10995,N_14297);
and U19136 (N_19136,N_13421,N_10893);
and U19137 (N_19137,N_12189,N_12033);
nand U19138 (N_19138,N_13820,N_14194);
or U19139 (N_19139,N_14765,N_11193);
and U19140 (N_19140,N_14478,N_10024);
or U19141 (N_19141,N_14436,N_13101);
nand U19142 (N_19142,N_11116,N_13818);
or U19143 (N_19143,N_10214,N_14848);
nand U19144 (N_19144,N_11688,N_10886);
or U19145 (N_19145,N_14814,N_12511);
nand U19146 (N_19146,N_10481,N_14743);
and U19147 (N_19147,N_10742,N_10670);
nand U19148 (N_19148,N_14701,N_11778);
nor U19149 (N_19149,N_11609,N_12530);
nor U19150 (N_19150,N_13203,N_13670);
or U19151 (N_19151,N_13721,N_13224);
nand U19152 (N_19152,N_13311,N_12130);
nand U19153 (N_19153,N_13765,N_10238);
nand U19154 (N_19154,N_13910,N_13420);
nand U19155 (N_19155,N_12616,N_13809);
and U19156 (N_19156,N_12395,N_14122);
and U19157 (N_19157,N_13403,N_13224);
and U19158 (N_19158,N_10028,N_12012);
or U19159 (N_19159,N_11783,N_11120);
or U19160 (N_19160,N_10334,N_10704);
or U19161 (N_19161,N_11640,N_10040);
nor U19162 (N_19162,N_10518,N_14901);
or U19163 (N_19163,N_13400,N_10417);
and U19164 (N_19164,N_13553,N_10300);
and U19165 (N_19165,N_12498,N_11226);
or U19166 (N_19166,N_14623,N_10614);
nand U19167 (N_19167,N_13610,N_12877);
and U19168 (N_19168,N_10164,N_10913);
nand U19169 (N_19169,N_10887,N_11279);
and U19170 (N_19170,N_14304,N_14253);
nor U19171 (N_19171,N_11423,N_11831);
nor U19172 (N_19172,N_12904,N_11950);
nand U19173 (N_19173,N_13742,N_14732);
nor U19174 (N_19174,N_14617,N_10783);
and U19175 (N_19175,N_12599,N_10000);
nand U19176 (N_19176,N_13769,N_12030);
and U19177 (N_19177,N_13250,N_11945);
nand U19178 (N_19178,N_10427,N_10264);
nand U19179 (N_19179,N_10268,N_12144);
nand U19180 (N_19180,N_10116,N_11863);
nor U19181 (N_19181,N_10247,N_10119);
or U19182 (N_19182,N_10358,N_11456);
or U19183 (N_19183,N_13223,N_12161);
nor U19184 (N_19184,N_12266,N_13698);
and U19185 (N_19185,N_11821,N_14208);
nand U19186 (N_19186,N_13519,N_14251);
nand U19187 (N_19187,N_10392,N_11704);
or U19188 (N_19188,N_10554,N_10607);
nand U19189 (N_19189,N_10493,N_14192);
nand U19190 (N_19190,N_11930,N_12174);
or U19191 (N_19191,N_11174,N_12976);
nand U19192 (N_19192,N_12882,N_12980);
nand U19193 (N_19193,N_14510,N_14965);
and U19194 (N_19194,N_11587,N_10666);
and U19195 (N_19195,N_11802,N_12090);
nand U19196 (N_19196,N_11442,N_10276);
and U19197 (N_19197,N_12672,N_12844);
nand U19198 (N_19198,N_13152,N_14309);
nor U19199 (N_19199,N_10136,N_14854);
and U19200 (N_19200,N_11974,N_12907);
and U19201 (N_19201,N_12877,N_14561);
and U19202 (N_19202,N_11542,N_10638);
nor U19203 (N_19203,N_14815,N_12286);
nand U19204 (N_19204,N_12404,N_13062);
and U19205 (N_19205,N_13880,N_11867);
or U19206 (N_19206,N_11778,N_11532);
or U19207 (N_19207,N_11475,N_12170);
and U19208 (N_19208,N_14678,N_12337);
and U19209 (N_19209,N_10869,N_12690);
and U19210 (N_19210,N_10215,N_11643);
or U19211 (N_19211,N_13344,N_11488);
or U19212 (N_19212,N_12786,N_11398);
nand U19213 (N_19213,N_12132,N_11895);
nor U19214 (N_19214,N_11843,N_11851);
or U19215 (N_19215,N_14517,N_14698);
nor U19216 (N_19216,N_12293,N_11134);
nor U19217 (N_19217,N_12142,N_12178);
or U19218 (N_19218,N_13189,N_11133);
or U19219 (N_19219,N_11114,N_14843);
nor U19220 (N_19220,N_13122,N_13104);
and U19221 (N_19221,N_14419,N_13884);
nor U19222 (N_19222,N_14461,N_13861);
or U19223 (N_19223,N_10574,N_12679);
nor U19224 (N_19224,N_11974,N_10830);
and U19225 (N_19225,N_14877,N_10546);
and U19226 (N_19226,N_13354,N_11422);
or U19227 (N_19227,N_13000,N_12632);
or U19228 (N_19228,N_14447,N_10587);
xor U19229 (N_19229,N_13807,N_13718);
nand U19230 (N_19230,N_10083,N_11034);
nor U19231 (N_19231,N_12847,N_14804);
or U19232 (N_19232,N_11539,N_12458);
and U19233 (N_19233,N_11406,N_10073);
nand U19234 (N_19234,N_13949,N_11903);
nor U19235 (N_19235,N_14573,N_10468);
nor U19236 (N_19236,N_10650,N_11702);
nand U19237 (N_19237,N_14722,N_12634);
or U19238 (N_19238,N_10047,N_10246);
nand U19239 (N_19239,N_14496,N_12071);
nor U19240 (N_19240,N_11055,N_11763);
and U19241 (N_19241,N_12293,N_13756);
or U19242 (N_19242,N_10948,N_11602);
xnor U19243 (N_19243,N_12392,N_11795);
and U19244 (N_19244,N_12611,N_12805);
nor U19245 (N_19245,N_13103,N_10756);
and U19246 (N_19246,N_10476,N_10364);
or U19247 (N_19247,N_14617,N_13863);
or U19248 (N_19248,N_14410,N_14273);
nand U19249 (N_19249,N_11877,N_11986);
xor U19250 (N_19250,N_14870,N_14529);
nand U19251 (N_19251,N_10839,N_12111);
and U19252 (N_19252,N_13566,N_11700);
nand U19253 (N_19253,N_12848,N_13005);
and U19254 (N_19254,N_10946,N_14199);
and U19255 (N_19255,N_12871,N_13460);
and U19256 (N_19256,N_13741,N_14267);
nor U19257 (N_19257,N_11545,N_14528);
and U19258 (N_19258,N_12434,N_14036);
nand U19259 (N_19259,N_11664,N_11328);
nor U19260 (N_19260,N_12672,N_10580);
and U19261 (N_19261,N_12402,N_10082);
or U19262 (N_19262,N_12021,N_12504);
nand U19263 (N_19263,N_14299,N_14518);
nor U19264 (N_19264,N_10465,N_10753);
and U19265 (N_19265,N_10876,N_13793);
nand U19266 (N_19266,N_14893,N_14925);
nor U19267 (N_19267,N_13365,N_13784);
or U19268 (N_19268,N_12059,N_14833);
nor U19269 (N_19269,N_10462,N_14162);
nor U19270 (N_19270,N_13192,N_13314);
nor U19271 (N_19271,N_12656,N_12789);
or U19272 (N_19272,N_11684,N_10490);
or U19273 (N_19273,N_14571,N_13462);
nand U19274 (N_19274,N_11620,N_12883);
or U19275 (N_19275,N_10035,N_13879);
nand U19276 (N_19276,N_13308,N_11695);
and U19277 (N_19277,N_12080,N_14252);
nor U19278 (N_19278,N_11288,N_12654);
nand U19279 (N_19279,N_10166,N_12128);
nor U19280 (N_19280,N_14934,N_11264);
nor U19281 (N_19281,N_11969,N_11827);
nand U19282 (N_19282,N_14019,N_10759);
nand U19283 (N_19283,N_13334,N_14513);
or U19284 (N_19284,N_11250,N_10544);
nand U19285 (N_19285,N_13688,N_14984);
and U19286 (N_19286,N_11582,N_11960);
nor U19287 (N_19287,N_11294,N_14007);
nor U19288 (N_19288,N_10026,N_12197);
nor U19289 (N_19289,N_12715,N_11976);
and U19290 (N_19290,N_10601,N_14207);
and U19291 (N_19291,N_14009,N_12942);
and U19292 (N_19292,N_10850,N_14107);
nor U19293 (N_19293,N_10034,N_11569);
or U19294 (N_19294,N_14363,N_14450);
nor U19295 (N_19295,N_11386,N_14141);
nor U19296 (N_19296,N_12520,N_10898);
nor U19297 (N_19297,N_11880,N_13920);
and U19298 (N_19298,N_10057,N_13603);
and U19299 (N_19299,N_13452,N_14831);
nand U19300 (N_19300,N_11791,N_12681);
nor U19301 (N_19301,N_12468,N_11443);
and U19302 (N_19302,N_11032,N_13611);
or U19303 (N_19303,N_10107,N_11769);
nand U19304 (N_19304,N_10110,N_14843);
or U19305 (N_19305,N_10061,N_13096);
or U19306 (N_19306,N_14227,N_13658);
nor U19307 (N_19307,N_14921,N_12254);
or U19308 (N_19308,N_12464,N_12434);
nor U19309 (N_19309,N_12205,N_11833);
nor U19310 (N_19310,N_12692,N_13566);
or U19311 (N_19311,N_11288,N_11186);
or U19312 (N_19312,N_13084,N_13036);
nand U19313 (N_19313,N_10302,N_11013);
nor U19314 (N_19314,N_12771,N_12338);
and U19315 (N_19315,N_11356,N_13267);
and U19316 (N_19316,N_14925,N_13574);
and U19317 (N_19317,N_10158,N_10078);
nand U19318 (N_19318,N_11846,N_11442);
nor U19319 (N_19319,N_14851,N_14512);
and U19320 (N_19320,N_13038,N_12495);
or U19321 (N_19321,N_13634,N_11380);
and U19322 (N_19322,N_12137,N_13870);
and U19323 (N_19323,N_14352,N_10223);
and U19324 (N_19324,N_10482,N_11610);
or U19325 (N_19325,N_14382,N_14802);
and U19326 (N_19326,N_14634,N_13379);
or U19327 (N_19327,N_10013,N_10081);
or U19328 (N_19328,N_13363,N_12296);
or U19329 (N_19329,N_10874,N_13396);
nor U19330 (N_19330,N_12493,N_13214);
and U19331 (N_19331,N_13443,N_12492);
nor U19332 (N_19332,N_14171,N_14446);
nand U19333 (N_19333,N_12105,N_10252);
and U19334 (N_19334,N_14359,N_12959);
nand U19335 (N_19335,N_10975,N_14300);
or U19336 (N_19336,N_14794,N_11851);
and U19337 (N_19337,N_12095,N_11499);
and U19338 (N_19338,N_14144,N_13465);
nor U19339 (N_19339,N_11530,N_12274);
and U19340 (N_19340,N_12695,N_14496);
or U19341 (N_19341,N_11534,N_12860);
and U19342 (N_19342,N_11899,N_11579);
or U19343 (N_19343,N_10662,N_13069);
nand U19344 (N_19344,N_12739,N_10093);
or U19345 (N_19345,N_12271,N_13711);
or U19346 (N_19346,N_13601,N_14029);
or U19347 (N_19347,N_10273,N_14770);
nand U19348 (N_19348,N_13636,N_10791);
nand U19349 (N_19349,N_11894,N_11188);
or U19350 (N_19350,N_13578,N_11240);
nand U19351 (N_19351,N_11337,N_10989);
or U19352 (N_19352,N_10414,N_12103);
and U19353 (N_19353,N_13228,N_11697);
and U19354 (N_19354,N_10989,N_13357);
and U19355 (N_19355,N_13552,N_12794);
nand U19356 (N_19356,N_12702,N_13410);
nand U19357 (N_19357,N_11412,N_13695);
nor U19358 (N_19358,N_10430,N_14339);
nor U19359 (N_19359,N_14097,N_11929);
and U19360 (N_19360,N_13028,N_10204);
or U19361 (N_19361,N_10522,N_12799);
and U19362 (N_19362,N_11568,N_14151);
and U19363 (N_19363,N_13877,N_14648);
and U19364 (N_19364,N_14007,N_12493);
xor U19365 (N_19365,N_12096,N_13217);
nand U19366 (N_19366,N_13673,N_12217);
or U19367 (N_19367,N_13839,N_11691);
and U19368 (N_19368,N_12684,N_14455);
and U19369 (N_19369,N_10861,N_10562);
nand U19370 (N_19370,N_10426,N_12471);
and U19371 (N_19371,N_10287,N_10137);
nand U19372 (N_19372,N_10574,N_10341);
and U19373 (N_19373,N_11981,N_14771);
and U19374 (N_19374,N_10033,N_14889);
nand U19375 (N_19375,N_12395,N_11245);
nand U19376 (N_19376,N_14800,N_10187);
and U19377 (N_19377,N_11569,N_11386);
nor U19378 (N_19378,N_11768,N_10492);
nand U19379 (N_19379,N_13123,N_10805);
and U19380 (N_19380,N_13472,N_13979);
and U19381 (N_19381,N_13906,N_11600);
and U19382 (N_19382,N_13044,N_11742);
or U19383 (N_19383,N_12630,N_14802);
xnor U19384 (N_19384,N_14451,N_11638);
and U19385 (N_19385,N_11395,N_14888);
and U19386 (N_19386,N_10998,N_12048);
nand U19387 (N_19387,N_11650,N_11813);
or U19388 (N_19388,N_13482,N_10771);
nand U19389 (N_19389,N_10247,N_12389);
and U19390 (N_19390,N_10707,N_11879);
nand U19391 (N_19391,N_13185,N_10192);
or U19392 (N_19392,N_13998,N_14111);
nor U19393 (N_19393,N_12099,N_11543);
and U19394 (N_19394,N_14934,N_12870);
nand U19395 (N_19395,N_13762,N_12085);
nand U19396 (N_19396,N_13619,N_10935);
nor U19397 (N_19397,N_11480,N_13941);
and U19398 (N_19398,N_11342,N_10898);
and U19399 (N_19399,N_14059,N_14783);
nand U19400 (N_19400,N_10755,N_13136);
nand U19401 (N_19401,N_12658,N_10811);
nand U19402 (N_19402,N_10657,N_10487);
nand U19403 (N_19403,N_14308,N_11533);
nand U19404 (N_19404,N_14878,N_13007);
or U19405 (N_19405,N_14652,N_10894);
nand U19406 (N_19406,N_10945,N_12573);
and U19407 (N_19407,N_11817,N_12766);
and U19408 (N_19408,N_14076,N_12289);
or U19409 (N_19409,N_11060,N_13650);
and U19410 (N_19410,N_12729,N_11695);
or U19411 (N_19411,N_14138,N_14641);
nor U19412 (N_19412,N_13660,N_10616);
or U19413 (N_19413,N_14703,N_14858);
nand U19414 (N_19414,N_10401,N_10932);
nand U19415 (N_19415,N_12193,N_11319);
or U19416 (N_19416,N_12507,N_12426);
or U19417 (N_19417,N_11708,N_11267);
nor U19418 (N_19418,N_12328,N_11368);
nor U19419 (N_19419,N_13438,N_13457);
or U19420 (N_19420,N_12145,N_14924);
nor U19421 (N_19421,N_13084,N_10002);
nor U19422 (N_19422,N_12390,N_12668);
or U19423 (N_19423,N_14459,N_11224);
or U19424 (N_19424,N_13792,N_11676);
or U19425 (N_19425,N_10467,N_10667);
or U19426 (N_19426,N_11056,N_13777);
and U19427 (N_19427,N_13601,N_10974);
or U19428 (N_19428,N_13976,N_11252);
or U19429 (N_19429,N_12846,N_10215);
or U19430 (N_19430,N_10446,N_13485);
nand U19431 (N_19431,N_12902,N_10130);
and U19432 (N_19432,N_12706,N_10559);
nand U19433 (N_19433,N_11159,N_12671);
or U19434 (N_19434,N_12437,N_10634);
nand U19435 (N_19435,N_11120,N_11203);
and U19436 (N_19436,N_13645,N_13528);
nor U19437 (N_19437,N_14104,N_13799);
nor U19438 (N_19438,N_12970,N_13581);
and U19439 (N_19439,N_14744,N_11219);
or U19440 (N_19440,N_12038,N_10365);
nor U19441 (N_19441,N_11822,N_10664);
nor U19442 (N_19442,N_12904,N_12294);
or U19443 (N_19443,N_10609,N_13310);
nor U19444 (N_19444,N_10111,N_10682);
and U19445 (N_19445,N_12144,N_10168);
nand U19446 (N_19446,N_10152,N_10918);
or U19447 (N_19447,N_14889,N_14140);
and U19448 (N_19448,N_12998,N_14500);
or U19449 (N_19449,N_13549,N_14797);
nor U19450 (N_19450,N_12424,N_10934);
and U19451 (N_19451,N_13051,N_10356);
or U19452 (N_19452,N_10511,N_12698);
nand U19453 (N_19453,N_14768,N_12428);
and U19454 (N_19454,N_11691,N_14945);
nand U19455 (N_19455,N_12868,N_11905);
and U19456 (N_19456,N_12767,N_13190);
or U19457 (N_19457,N_11068,N_11376);
and U19458 (N_19458,N_10264,N_14653);
or U19459 (N_19459,N_14267,N_13821);
or U19460 (N_19460,N_11849,N_14933);
and U19461 (N_19461,N_10164,N_12058);
or U19462 (N_19462,N_14185,N_12941);
or U19463 (N_19463,N_13136,N_13223);
xor U19464 (N_19464,N_12434,N_14277);
nor U19465 (N_19465,N_10085,N_12175);
or U19466 (N_19466,N_12922,N_10638);
and U19467 (N_19467,N_11439,N_14174);
nand U19468 (N_19468,N_11400,N_14725);
nand U19469 (N_19469,N_10503,N_13205);
nor U19470 (N_19470,N_13394,N_14123);
and U19471 (N_19471,N_14592,N_13869);
nand U19472 (N_19472,N_14101,N_12245);
or U19473 (N_19473,N_11631,N_11422);
nand U19474 (N_19474,N_11248,N_11874);
or U19475 (N_19475,N_13794,N_11483);
and U19476 (N_19476,N_13781,N_13133);
or U19477 (N_19477,N_13793,N_12201);
nand U19478 (N_19478,N_10780,N_14100);
or U19479 (N_19479,N_11673,N_13636);
or U19480 (N_19480,N_11949,N_11212);
and U19481 (N_19481,N_11405,N_14676);
and U19482 (N_19482,N_13080,N_13047);
nor U19483 (N_19483,N_13426,N_11811);
and U19484 (N_19484,N_14340,N_10866);
and U19485 (N_19485,N_14607,N_12227);
or U19486 (N_19486,N_13984,N_13088);
and U19487 (N_19487,N_13584,N_14836);
nand U19488 (N_19488,N_14978,N_14708);
nor U19489 (N_19489,N_12379,N_13407);
nor U19490 (N_19490,N_11166,N_14392);
nand U19491 (N_19491,N_11628,N_10493);
and U19492 (N_19492,N_14538,N_13864);
and U19493 (N_19493,N_14774,N_12032);
and U19494 (N_19494,N_14564,N_10524);
or U19495 (N_19495,N_12522,N_10005);
nor U19496 (N_19496,N_10944,N_12685);
or U19497 (N_19497,N_14125,N_11551);
and U19498 (N_19498,N_13167,N_10363);
or U19499 (N_19499,N_13194,N_11113);
nor U19500 (N_19500,N_13916,N_11618);
nor U19501 (N_19501,N_12943,N_10961);
nand U19502 (N_19502,N_10042,N_14032);
nor U19503 (N_19503,N_13673,N_10899);
or U19504 (N_19504,N_12641,N_13732);
or U19505 (N_19505,N_11856,N_12394);
or U19506 (N_19506,N_10259,N_10523);
or U19507 (N_19507,N_13024,N_11749);
and U19508 (N_19508,N_11751,N_12128);
and U19509 (N_19509,N_14631,N_14234);
and U19510 (N_19510,N_11252,N_12277);
nand U19511 (N_19511,N_14752,N_14172);
nor U19512 (N_19512,N_14138,N_12381);
or U19513 (N_19513,N_13131,N_10303);
nand U19514 (N_19514,N_14070,N_14503);
nor U19515 (N_19515,N_14797,N_11858);
nor U19516 (N_19516,N_14478,N_12105);
or U19517 (N_19517,N_14688,N_14573);
or U19518 (N_19518,N_10533,N_14655);
and U19519 (N_19519,N_10967,N_10220);
nand U19520 (N_19520,N_10171,N_12092);
or U19521 (N_19521,N_14213,N_11344);
and U19522 (N_19522,N_14743,N_11577);
and U19523 (N_19523,N_13512,N_14834);
and U19524 (N_19524,N_12014,N_13625);
and U19525 (N_19525,N_13889,N_11916);
and U19526 (N_19526,N_13481,N_13265);
and U19527 (N_19527,N_10894,N_14912);
nand U19528 (N_19528,N_10063,N_12415);
nor U19529 (N_19529,N_11331,N_10046);
nand U19530 (N_19530,N_13402,N_10597);
nor U19531 (N_19531,N_13149,N_14183);
and U19532 (N_19532,N_14279,N_12373);
and U19533 (N_19533,N_12605,N_13940);
or U19534 (N_19534,N_10504,N_13793);
nand U19535 (N_19535,N_12164,N_13203);
or U19536 (N_19536,N_14097,N_12446);
nor U19537 (N_19537,N_11535,N_13740);
and U19538 (N_19538,N_10392,N_14842);
nand U19539 (N_19539,N_13972,N_10350);
or U19540 (N_19540,N_14734,N_10993);
or U19541 (N_19541,N_10766,N_11793);
nor U19542 (N_19542,N_11598,N_10100);
nor U19543 (N_19543,N_13255,N_11093);
nor U19544 (N_19544,N_13471,N_13731);
nand U19545 (N_19545,N_12641,N_12831);
nand U19546 (N_19546,N_13381,N_14638);
nor U19547 (N_19547,N_11111,N_14499);
nor U19548 (N_19548,N_10758,N_12956);
nand U19549 (N_19549,N_13862,N_11176);
or U19550 (N_19550,N_11720,N_10308);
nor U19551 (N_19551,N_10108,N_12790);
nand U19552 (N_19552,N_12157,N_11339);
and U19553 (N_19553,N_12301,N_12809);
nor U19554 (N_19554,N_13141,N_10763);
nor U19555 (N_19555,N_13964,N_13364);
xnor U19556 (N_19556,N_14806,N_11636);
nor U19557 (N_19557,N_10404,N_11101);
nand U19558 (N_19558,N_11721,N_10208);
or U19559 (N_19559,N_14420,N_13751);
nand U19560 (N_19560,N_13657,N_12112);
nor U19561 (N_19561,N_14682,N_10001);
nand U19562 (N_19562,N_12423,N_13397);
nor U19563 (N_19563,N_10100,N_13124);
and U19564 (N_19564,N_10037,N_13813);
nor U19565 (N_19565,N_12903,N_13408);
and U19566 (N_19566,N_11313,N_12298);
or U19567 (N_19567,N_14199,N_14860);
nor U19568 (N_19568,N_13806,N_10664);
or U19569 (N_19569,N_11542,N_14212);
and U19570 (N_19570,N_10232,N_14833);
or U19571 (N_19571,N_14382,N_13694);
and U19572 (N_19572,N_14525,N_12746);
and U19573 (N_19573,N_13228,N_12125);
and U19574 (N_19574,N_14885,N_14179);
and U19575 (N_19575,N_10032,N_14829);
nand U19576 (N_19576,N_12401,N_13725);
nand U19577 (N_19577,N_13290,N_12222);
nor U19578 (N_19578,N_11008,N_12950);
and U19579 (N_19579,N_10084,N_12571);
nor U19580 (N_19580,N_11378,N_11207);
nand U19581 (N_19581,N_10164,N_14035);
nand U19582 (N_19582,N_14468,N_14208);
nor U19583 (N_19583,N_13838,N_14326);
nor U19584 (N_19584,N_13925,N_13887);
or U19585 (N_19585,N_14574,N_10424);
nand U19586 (N_19586,N_11479,N_13584);
and U19587 (N_19587,N_11900,N_11589);
nor U19588 (N_19588,N_10112,N_10527);
nand U19589 (N_19589,N_12297,N_13265);
nand U19590 (N_19590,N_12121,N_12270);
and U19591 (N_19591,N_14716,N_14687);
nor U19592 (N_19592,N_12395,N_12288);
nand U19593 (N_19593,N_12789,N_10028);
nor U19594 (N_19594,N_11315,N_11670);
nor U19595 (N_19595,N_12950,N_13235);
nand U19596 (N_19596,N_11313,N_14378);
or U19597 (N_19597,N_14170,N_14555);
and U19598 (N_19598,N_13732,N_13428);
nor U19599 (N_19599,N_10779,N_14577);
nand U19600 (N_19600,N_14797,N_11105);
or U19601 (N_19601,N_12559,N_12658);
nand U19602 (N_19602,N_11943,N_14768);
or U19603 (N_19603,N_13137,N_13202);
or U19604 (N_19604,N_10893,N_12293);
nor U19605 (N_19605,N_13476,N_11983);
nand U19606 (N_19606,N_11004,N_13322);
and U19607 (N_19607,N_13959,N_14369);
nand U19608 (N_19608,N_12723,N_11027);
and U19609 (N_19609,N_10817,N_10471);
nor U19610 (N_19610,N_14159,N_12236);
or U19611 (N_19611,N_14913,N_13385);
and U19612 (N_19612,N_10928,N_13097);
and U19613 (N_19613,N_14150,N_10694);
nand U19614 (N_19614,N_14139,N_14931);
nor U19615 (N_19615,N_11247,N_12169);
nand U19616 (N_19616,N_12464,N_12719);
or U19617 (N_19617,N_14186,N_14694);
xnor U19618 (N_19618,N_11676,N_13415);
nor U19619 (N_19619,N_10455,N_10699);
and U19620 (N_19620,N_14017,N_10435);
or U19621 (N_19621,N_13177,N_14779);
nand U19622 (N_19622,N_11455,N_10443);
or U19623 (N_19623,N_13660,N_11598);
nor U19624 (N_19624,N_10821,N_12686);
or U19625 (N_19625,N_13432,N_14968);
nor U19626 (N_19626,N_11261,N_13142);
nand U19627 (N_19627,N_14989,N_10438);
nand U19628 (N_19628,N_12658,N_10738);
nand U19629 (N_19629,N_11953,N_14151);
nor U19630 (N_19630,N_14345,N_13470);
and U19631 (N_19631,N_11966,N_11579);
nand U19632 (N_19632,N_14548,N_11685);
or U19633 (N_19633,N_12480,N_11845);
nand U19634 (N_19634,N_11761,N_14309);
and U19635 (N_19635,N_13062,N_10431);
or U19636 (N_19636,N_10229,N_10684);
xnor U19637 (N_19637,N_14270,N_11293);
nor U19638 (N_19638,N_13525,N_12954);
nor U19639 (N_19639,N_10847,N_12444);
and U19640 (N_19640,N_14035,N_10206);
nand U19641 (N_19641,N_10475,N_10826);
nand U19642 (N_19642,N_12693,N_10179);
nor U19643 (N_19643,N_12278,N_11904);
or U19644 (N_19644,N_13420,N_11459);
nand U19645 (N_19645,N_14558,N_13756);
nor U19646 (N_19646,N_11625,N_12843);
or U19647 (N_19647,N_11332,N_11145);
or U19648 (N_19648,N_10879,N_12946);
nor U19649 (N_19649,N_10371,N_14148);
nor U19650 (N_19650,N_13128,N_10570);
nand U19651 (N_19651,N_14702,N_10954);
or U19652 (N_19652,N_11440,N_12264);
nor U19653 (N_19653,N_14002,N_10615);
and U19654 (N_19654,N_14186,N_12386);
and U19655 (N_19655,N_12237,N_13091);
nor U19656 (N_19656,N_13956,N_12170);
nand U19657 (N_19657,N_13036,N_10798);
nand U19658 (N_19658,N_13343,N_12885);
and U19659 (N_19659,N_10661,N_14976);
or U19660 (N_19660,N_12157,N_10238);
or U19661 (N_19661,N_10503,N_12428);
nand U19662 (N_19662,N_14351,N_10817);
nor U19663 (N_19663,N_14814,N_10917);
nand U19664 (N_19664,N_14226,N_14121);
nor U19665 (N_19665,N_11389,N_11937);
nor U19666 (N_19666,N_14831,N_12079);
nor U19667 (N_19667,N_11267,N_14484);
nor U19668 (N_19668,N_10417,N_11429);
nand U19669 (N_19669,N_13707,N_13905);
nor U19670 (N_19670,N_12743,N_11254);
nor U19671 (N_19671,N_12462,N_12925);
and U19672 (N_19672,N_14601,N_11931);
or U19673 (N_19673,N_10985,N_10370);
or U19674 (N_19674,N_12674,N_13299);
and U19675 (N_19675,N_14376,N_12825);
and U19676 (N_19676,N_14788,N_12272);
nor U19677 (N_19677,N_14767,N_12638);
and U19678 (N_19678,N_12380,N_10199);
or U19679 (N_19679,N_12668,N_11851);
nor U19680 (N_19680,N_12275,N_13240);
or U19681 (N_19681,N_11641,N_13641);
nand U19682 (N_19682,N_14433,N_13962);
and U19683 (N_19683,N_14152,N_12462);
nand U19684 (N_19684,N_13558,N_13971);
nor U19685 (N_19685,N_12898,N_13953);
nor U19686 (N_19686,N_14707,N_14122);
nand U19687 (N_19687,N_14560,N_11177);
and U19688 (N_19688,N_13222,N_12339);
and U19689 (N_19689,N_12903,N_13171);
and U19690 (N_19690,N_12992,N_14261);
or U19691 (N_19691,N_11435,N_11216);
or U19692 (N_19692,N_13924,N_11922);
and U19693 (N_19693,N_13380,N_12480);
or U19694 (N_19694,N_11389,N_12537);
or U19695 (N_19695,N_10671,N_13270);
or U19696 (N_19696,N_13431,N_12203);
and U19697 (N_19697,N_10334,N_10291);
and U19698 (N_19698,N_14719,N_14758);
nor U19699 (N_19699,N_13908,N_13327);
or U19700 (N_19700,N_11431,N_10865);
nand U19701 (N_19701,N_11620,N_14944);
and U19702 (N_19702,N_10003,N_10285);
or U19703 (N_19703,N_10925,N_10030);
or U19704 (N_19704,N_14467,N_10564);
nand U19705 (N_19705,N_14015,N_11946);
nand U19706 (N_19706,N_11255,N_13227);
nor U19707 (N_19707,N_10362,N_13959);
or U19708 (N_19708,N_14844,N_11318);
and U19709 (N_19709,N_12502,N_10916);
or U19710 (N_19710,N_13480,N_11156);
nand U19711 (N_19711,N_11812,N_12623);
or U19712 (N_19712,N_14751,N_12632);
or U19713 (N_19713,N_13432,N_10916);
and U19714 (N_19714,N_14217,N_12052);
nand U19715 (N_19715,N_11519,N_10850);
nor U19716 (N_19716,N_13394,N_13903);
nand U19717 (N_19717,N_10900,N_10030);
nor U19718 (N_19718,N_13427,N_12986);
nor U19719 (N_19719,N_10934,N_14017);
nand U19720 (N_19720,N_12989,N_10156);
nand U19721 (N_19721,N_12253,N_13885);
nor U19722 (N_19722,N_12469,N_11636);
nor U19723 (N_19723,N_13128,N_11750);
or U19724 (N_19724,N_11325,N_10650);
nand U19725 (N_19725,N_14570,N_11783);
and U19726 (N_19726,N_13911,N_10715);
or U19727 (N_19727,N_11110,N_14219);
nor U19728 (N_19728,N_14403,N_14095);
and U19729 (N_19729,N_12662,N_11630);
or U19730 (N_19730,N_10897,N_11648);
or U19731 (N_19731,N_11821,N_12684);
nand U19732 (N_19732,N_13918,N_10983);
nand U19733 (N_19733,N_14395,N_14110);
nor U19734 (N_19734,N_14459,N_13090);
or U19735 (N_19735,N_10888,N_10707);
or U19736 (N_19736,N_11531,N_10765);
or U19737 (N_19737,N_10091,N_13787);
or U19738 (N_19738,N_13008,N_11440);
nor U19739 (N_19739,N_12473,N_11436);
and U19740 (N_19740,N_13436,N_13031);
and U19741 (N_19741,N_12122,N_14650);
nand U19742 (N_19742,N_10402,N_14302);
nand U19743 (N_19743,N_12365,N_13471);
and U19744 (N_19744,N_10238,N_12386);
nand U19745 (N_19745,N_10234,N_11004);
nand U19746 (N_19746,N_11680,N_11660);
nand U19747 (N_19747,N_12296,N_12810);
nor U19748 (N_19748,N_13424,N_12963);
or U19749 (N_19749,N_10082,N_14102);
or U19750 (N_19750,N_14083,N_10890);
and U19751 (N_19751,N_11919,N_12082);
and U19752 (N_19752,N_14412,N_12014);
and U19753 (N_19753,N_10349,N_13344);
and U19754 (N_19754,N_13156,N_14479);
and U19755 (N_19755,N_14927,N_11505);
or U19756 (N_19756,N_13266,N_14743);
nor U19757 (N_19757,N_11682,N_12833);
nand U19758 (N_19758,N_14223,N_12874);
and U19759 (N_19759,N_13588,N_12386);
or U19760 (N_19760,N_10146,N_14543);
nand U19761 (N_19761,N_10676,N_12258);
and U19762 (N_19762,N_12878,N_13085);
nor U19763 (N_19763,N_14765,N_11905);
xnor U19764 (N_19764,N_14588,N_14302);
or U19765 (N_19765,N_12169,N_12648);
xnor U19766 (N_19766,N_11452,N_13097);
and U19767 (N_19767,N_11321,N_10455);
or U19768 (N_19768,N_12718,N_10189);
nor U19769 (N_19769,N_12894,N_13527);
nand U19770 (N_19770,N_14037,N_11554);
nand U19771 (N_19771,N_11778,N_14754);
nor U19772 (N_19772,N_14659,N_10017);
nor U19773 (N_19773,N_13536,N_11430);
or U19774 (N_19774,N_13032,N_10610);
and U19775 (N_19775,N_14888,N_14749);
nand U19776 (N_19776,N_11530,N_10110);
and U19777 (N_19777,N_12606,N_13850);
nand U19778 (N_19778,N_13178,N_14883);
or U19779 (N_19779,N_11603,N_11502);
or U19780 (N_19780,N_10705,N_12011);
or U19781 (N_19781,N_11525,N_11947);
nand U19782 (N_19782,N_11813,N_14266);
nand U19783 (N_19783,N_11157,N_14657);
nor U19784 (N_19784,N_14376,N_10815);
or U19785 (N_19785,N_14109,N_10203);
nor U19786 (N_19786,N_14530,N_14902);
nand U19787 (N_19787,N_10641,N_10469);
nand U19788 (N_19788,N_13259,N_11083);
or U19789 (N_19789,N_11674,N_11691);
nand U19790 (N_19790,N_10178,N_13007);
and U19791 (N_19791,N_13872,N_12147);
and U19792 (N_19792,N_14219,N_13547);
or U19793 (N_19793,N_14889,N_11332);
nor U19794 (N_19794,N_13855,N_13521);
nor U19795 (N_19795,N_13399,N_11884);
nand U19796 (N_19796,N_11783,N_12365);
and U19797 (N_19797,N_12094,N_13493);
nor U19798 (N_19798,N_13477,N_12961);
nand U19799 (N_19799,N_11951,N_14241);
or U19800 (N_19800,N_14092,N_11017);
nand U19801 (N_19801,N_12802,N_14092);
or U19802 (N_19802,N_11894,N_12283);
or U19803 (N_19803,N_12689,N_12483);
and U19804 (N_19804,N_10536,N_14210);
and U19805 (N_19805,N_14865,N_10526);
nor U19806 (N_19806,N_12182,N_10245);
xor U19807 (N_19807,N_11872,N_10787);
and U19808 (N_19808,N_14476,N_11879);
or U19809 (N_19809,N_14129,N_10843);
nand U19810 (N_19810,N_12470,N_14142);
nand U19811 (N_19811,N_11716,N_12134);
and U19812 (N_19812,N_12622,N_14302);
nand U19813 (N_19813,N_12996,N_14339);
nand U19814 (N_19814,N_10267,N_10810);
nor U19815 (N_19815,N_13433,N_12977);
nor U19816 (N_19816,N_14822,N_12412);
or U19817 (N_19817,N_13946,N_10869);
nor U19818 (N_19818,N_10435,N_12789);
or U19819 (N_19819,N_11149,N_10191);
or U19820 (N_19820,N_10486,N_11465);
nand U19821 (N_19821,N_11223,N_11143);
or U19822 (N_19822,N_14002,N_10417);
or U19823 (N_19823,N_14649,N_11661);
and U19824 (N_19824,N_10452,N_11733);
nor U19825 (N_19825,N_11910,N_13409);
and U19826 (N_19826,N_12390,N_12651);
nor U19827 (N_19827,N_14437,N_10077);
or U19828 (N_19828,N_13866,N_14906);
and U19829 (N_19829,N_10802,N_13288);
or U19830 (N_19830,N_13986,N_11043);
and U19831 (N_19831,N_13951,N_11754);
and U19832 (N_19832,N_14989,N_12596);
nor U19833 (N_19833,N_13112,N_13893);
nand U19834 (N_19834,N_12885,N_14441);
nor U19835 (N_19835,N_10526,N_11733);
nand U19836 (N_19836,N_13830,N_12955);
nand U19837 (N_19837,N_13711,N_14580);
nand U19838 (N_19838,N_11321,N_13735);
nor U19839 (N_19839,N_13976,N_10606);
nor U19840 (N_19840,N_10593,N_13319);
nand U19841 (N_19841,N_10334,N_12842);
nor U19842 (N_19842,N_12565,N_13636);
nand U19843 (N_19843,N_14284,N_10497);
nand U19844 (N_19844,N_11189,N_14197);
nand U19845 (N_19845,N_11609,N_12708);
nand U19846 (N_19846,N_11313,N_11218);
and U19847 (N_19847,N_10703,N_11557);
nor U19848 (N_19848,N_10549,N_11670);
and U19849 (N_19849,N_11378,N_13822);
and U19850 (N_19850,N_10809,N_11114);
and U19851 (N_19851,N_10551,N_12647);
nand U19852 (N_19852,N_10494,N_14626);
and U19853 (N_19853,N_11283,N_12661);
or U19854 (N_19854,N_12898,N_11604);
or U19855 (N_19855,N_12128,N_13359);
nand U19856 (N_19856,N_12541,N_10135);
or U19857 (N_19857,N_12022,N_14043);
nand U19858 (N_19858,N_11990,N_12747);
and U19859 (N_19859,N_11773,N_12003);
or U19860 (N_19860,N_14249,N_10852);
nand U19861 (N_19861,N_10905,N_12269);
and U19862 (N_19862,N_12788,N_13878);
or U19863 (N_19863,N_11289,N_11702);
and U19864 (N_19864,N_14512,N_13126);
nor U19865 (N_19865,N_14523,N_14979);
nand U19866 (N_19866,N_12150,N_12947);
or U19867 (N_19867,N_12576,N_14839);
nor U19868 (N_19868,N_10196,N_10087);
or U19869 (N_19869,N_13026,N_13742);
nor U19870 (N_19870,N_10060,N_14183);
or U19871 (N_19871,N_10474,N_12728);
and U19872 (N_19872,N_13295,N_10681);
and U19873 (N_19873,N_10321,N_10496);
and U19874 (N_19874,N_14784,N_13308);
nor U19875 (N_19875,N_10384,N_10539);
and U19876 (N_19876,N_11820,N_10691);
or U19877 (N_19877,N_12949,N_14328);
nand U19878 (N_19878,N_14744,N_13833);
nor U19879 (N_19879,N_13618,N_10179);
or U19880 (N_19880,N_13291,N_14681);
or U19881 (N_19881,N_13541,N_10169);
or U19882 (N_19882,N_12000,N_13925);
or U19883 (N_19883,N_10567,N_14383);
and U19884 (N_19884,N_14903,N_13577);
nor U19885 (N_19885,N_13467,N_14753);
nand U19886 (N_19886,N_11289,N_10427);
nand U19887 (N_19887,N_10024,N_12437);
or U19888 (N_19888,N_13946,N_10720);
or U19889 (N_19889,N_14129,N_10692);
or U19890 (N_19890,N_14165,N_10739);
nor U19891 (N_19891,N_11244,N_13091);
nor U19892 (N_19892,N_10532,N_10617);
or U19893 (N_19893,N_14623,N_10622);
and U19894 (N_19894,N_13378,N_10659);
and U19895 (N_19895,N_10792,N_11375);
or U19896 (N_19896,N_10249,N_11066);
or U19897 (N_19897,N_12510,N_11405);
nand U19898 (N_19898,N_11290,N_14045);
and U19899 (N_19899,N_11320,N_10731);
nand U19900 (N_19900,N_10237,N_14082);
nor U19901 (N_19901,N_13528,N_10890);
and U19902 (N_19902,N_13819,N_10630);
and U19903 (N_19903,N_12543,N_14913);
nor U19904 (N_19904,N_12670,N_11632);
and U19905 (N_19905,N_12283,N_11739);
or U19906 (N_19906,N_11201,N_12590);
nand U19907 (N_19907,N_11183,N_10083);
or U19908 (N_19908,N_11219,N_14356);
nor U19909 (N_19909,N_10265,N_13136);
or U19910 (N_19910,N_12267,N_14250);
nor U19911 (N_19911,N_11779,N_14608);
or U19912 (N_19912,N_14599,N_12106);
and U19913 (N_19913,N_11719,N_14098);
nor U19914 (N_19914,N_13307,N_14736);
nand U19915 (N_19915,N_11932,N_13417);
nand U19916 (N_19916,N_13670,N_13175);
or U19917 (N_19917,N_12249,N_11823);
or U19918 (N_19918,N_12371,N_13891);
and U19919 (N_19919,N_12070,N_10732);
or U19920 (N_19920,N_14762,N_12226);
nor U19921 (N_19921,N_12335,N_11619);
and U19922 (N_19922,N_12540,N_13083);
nor U19923 (N_19923,N_10865,N_13928);
and U19924 (N_19924,N_13529,N_12863);
or U19925 (N_19925,N_11476,N_14167);
or U19926 (N_19926,N_13361,N_12394);
and U19927 (N_19927,N_13279,N_14474);
nand U19928 (N_19928,N_10711,N_10551);
nor U19929 (N_19929,N_13529,N_14380);
nor U19930 (N_19930,N_14618,N_11304);
or U19931 (N_19931,N_10007,N_11187);
nand U19932 (N_19932,N_14118,N_11961);
and U19933 (N_19933,N_14523,N_10677);
nand U19934 (N_19934,N_12066,N_13945);
and U19935 (N_19935,N_12570,N_12324);
and U19936 (N_19936,N_12458,N_14468);
nor U19937 (N_19937,N_11136,N_13283);
nand U19938 (N_19938,N_12824,N_10812);
or U19939 (N_19939,N_13986,N_13183);
nand U19940 (N_19940,N_12365,N_11152);
and U19941 (N_19941,N_11998,N_10458);
or U19942 (N_19942,N_11129,N_14881);
or U19943 (N_19943,N_14298,N_12289);
and U19944 (N_19944,N_11487,N_10575);
or U19945 (N_19945,N_14264,N_11500);
or U19946 (N_19946,N_12002,N_12257);
nand U19947 (N_19947,N_12609,N_12784);
or U19948 (N_19948,N_10230,N_14107);
or U19949 (N_19949,N_11660,N_11006);
nor U19950 (N_19950,N_13610,N_12019);
and U19951 (N_19951,N_13757,N_14070);
nand U19952 (N_19952,N_11679,N_14872);
and U19953 (N_19953,N_11244,N_10910);
nand U19954 (N_19954,N_11242,N_12457);
or U19955 (N_19955,N_11147,N_13150);
and U19956 (N_19956,N_11886,N_14312);
nor U19957 (N_19957,N_11134,N_11051);
and U19958 (N_19958,N_12940,N_13627);
nand U19959 (N_19959,N_14066,N_11178);
nor U19960 (N_19960,N_11935,N_12489);
and U19961 (N_19961,N_12245,N_11709);
or U19962 (N_19962,N_13036,N_10214);
nor U19963 (N_19963,N_13477,N_13219);
nand U19964 (N_19964,N_14213,N_14824);
nand U19965 (N_19965,N_13939,N_14769);
nand U19966 (N_19966,N_12513,N_14884);
and U19967 (N_19967,N_10511,N_11059);
nor U19968 (N_19968,N_11034,N_10798);
or U19969 (N_19969,N_13050,N_14701);
nor U19970 (N_19970,N_13472,N_14292);
and U19971 (N_19971,N_13894,N_11787);
and U19972 (N_19972,N_12717,N_12574);
nand U19973 (N_19973,N_12920,N_14523);
and U19974 (N_19974,N_10795,N_12506);
xnor U19975 (N_19975,N_10717,N_13347);
nand U19976 (N_19976,N_10435,N_14067);
and U19977 (N_19977,N_14944,N_11925);
and U19978 (N_19978,N_14884,N_10628);
or U19979 (N_19979,N_11193,N_12321);
nor U19980 (N_19980,N_10157,N_13178);
and U19981 (N_19981,N_12519,N_14669);
nor U19982 (N_19982,N_14902,N_11243);
nor U19983 (N_19983,N_12334,N_13356);
and U19984 (N_19984,N_14743,N_13297);
and U19985 (N_19985,N_10543,N_12282);
and U19986 (N_19986,N_10685,N_10312);
nand U19987 (N_19987,N_13623,N_11092);
nor U19988 (N_19988,N_11851,N_14944);
nor U19989 (N_19989,N_14018,N_10985);
nand U19990 (N_19990,N_14837,N_14776);
nor U19991 (N_19991,N_14829,N_13682);
and U19992 (N_19992,N_12926,N_13836);
or U19993 (N_19993,N_11748,N_12231);
and U19994 (N_19994,N_14077,N_11002);
and U19995 (N_19995,N_10543,N_10648);
nand U19996 (N_19996,N_14170,N_13846);
nor U19997 (N_19997,N_11368,N_11202);
nand U19998 (N_19998,N_12878,N_11193);
nand U19999 (N_19999,N_11459,N_13752);
nand U20000 (N_20000,N_15851,N_17126);
nor U20001 (N_20001,N_17497,N_17862);
or U20002 (N_20002,N_18013,N_18202);
and U20003 (N_20003,N_19186,N_15106);
xnor U20004 (N_20004,N_18021,N_15618);
or U20005 (N_20005,N_17018,N_16332);
nand U20006 (N_20006,N_15627,N_15317);
or U20007 (N_20007,N_17581,N_17550);
or U20008 (N_20008,N_17778,N_18542);
nor U20009 (N_20009,N_16906,N_18274);
and U20010 (N_20010,N_19891,N_16593);
and U20011 (N_20011,N_16860,N_19430);
and U20012 (N_20012,N_17047,N_18303);
and U20013 (N_20013,N_19144,N_17881);
or U20014 (N_20014,N_16516,N_16165);
or U20015 (N_20015,N_15988,N_19505);
and U20016 (N_20016,N_19480,N_17678);
nor U20017 (N_20017,N_18623,N_19214);
nor U20018 (N_20018,N_16499,N_18036);
and U20019 (N_20019,N_17736,N_15378);
nor U20020 (N_20020,N_19721,N_18364);
xor U20021 (N_20021,N_19905,N_16340);
and U20022 (N_20022,N_15292,N_19051);
nor U20023 (N_20023,N_16067,N_18173);
and U20024 (N_20024,N_16954,N_19844);
and U20025 (N_20025,N_17857,N_15179);
nand U20026 (N_20026,N_17225,N_18317);
nand U20027 (N_20027,N_16508,N_17715);
nor U20028 (N_20028,N_19591,N_18095);
and U20029 (N_20029,N_18340,N_17615);
nand U20030 (N_20030,N_15725,N_18983);
nor U20031 (N_20031,N_19936,N_16733);
and U20032 (N_20032,N_16386,N_18804);
nand U20033 (N_20033,N_15981,N_17929);
nor U20034 (N_20034,N_16760,N_19823);
nor U20035 (N_20035,N_18357,N_18796);
nand U20036 (N_20036,N_16627,N_15726);
or U20037 (N_20037,N_18179,N_15533);
or U20038 (N_20038,N_16708,N_15503);
and U20039 (N_20039,N_19659,N_19162);
and U20040 (N_20040,N_18496,N_18833);
or U20041 (N_20041,N_17781,N_16767);
and U20042 (N_20042,N_19388,N_16958);
and U20043 (N_20043,N_17396,N_17183);
nand U20044 (N_20044,N_19319,N_19990);
nor U20045 (N_20045,N_16521,N_16607);
or U20046 (N_20046,N_18866,N_19366);
or U20047 (N_20047,N_16515,N_18053);
or U20048 (N_20048,N_15274,N_17888);
and U20049 (N_20049,N_19229,N_15285);
or U20050 (N_20050,N_18911,N_19190);
and U20051 (N_20051,N_16232,N_18138);
and U20052 (N_20052,N_18384,N_19998);
nand U20053 (N_20053,N_16898,N_18846);
nand U20054 (N_20054,N_17814,N_19027);
nor U20055 (N_20055,N_16376,N_16227);
nor U20056 (N_20056,N_18932,N_19638);
or U20057 (N_20057,N_18620,N_16625);
nor U20058 (N_20058,N_16098,N_19154);
nand U20059 (N_20059,N_19237,N_19083);
and U20060 (N_20060,N_19524,N_16604);
nor U20061 (N_20061,N_17574,N_15247);
nor U20062 (N_20062,N_15461,N_18997);
nand U20063 (N_20063,N_19254,N_16816);
or U20064 (N_20064,N_17690,N_15775);
nand U20065 (N_20065,N_17883,N_18280);
nor U20066 (N_20066,N_16002,N_19878);
and U20067 (N_20067,N_15468,N_17142);
or U20068 (N_20068,N_17505,N_16777);
or U20069 (N_20069,N_15566,N_18743);
nand U20070 (N_20070,N_16922,N_15642);
nor U20071 (N_20071,N_19618,N_16037);
nand U20072 (N_20072,N_16565,N_15058);
or U20073 (N_20073,N_19493,N_19651);
nor U20074 (N_20074,N_18577,N_15971);
nor U20075 (N_20075,N_18616,N_18321);
nand U20076 (N_20076,N_17792,N_19065);
and U20077 (N_20077,N_16281,N_19139);
or U20078 (N_20078,N_15753,N_18196);
nand U20079 (N_20079,N_15118,N_15928);
nor U20080 (N_20080,N_16448,N_17924);
nand U20081 (N_20081,N_15326,N_18417);
or U20082 (N_20082,N_19966,N_15758);
nand U20083 (N_20083,N_19403,N_16036);
and U20084 (N_20084,N_19017,N_18830);
or U20085 (N_20085,N_17956,N_15830);
or U20086 (N_20086,N_19794,N_16579);
and U20087 (N_20087,N_16520,N_15211);
nand U20088 (N_20088,N_17145,N_16907);
nor U20089 (N_20089,N_18176,N_18134);
nand U20090 (N_20090,N_19760,N_16852);
nand U20091 (N_20091,N_16892,N_16570);
nand U20092 (N_20092,N_16985,N_15575);
or U20093 (N_20093,N_17073,N_17930);
nand U20094 (N_20094,N_15246,N_15440);
nor U20095 (N_20095,N_19506,N_17703);
and U20096 (N_20096,N_19509,N_19642);
or U20097 (N_20097,N_16897,N_19255);
nand U20098 (N_20098,N_15587,N_17522);
nor U20099 (N_20099,N_15149,N_16877);
nor U20100 (N_20100,N_18604,N_18703);
nand U20101 (N_20101,N_17262,N_19071);
and U20102 (N_20102,N_15452,N_18211);
nand U20103 (N_20103,N_18860,N_17007);
and U20104 (N_20104,N_15644,N_17952);
or U20105 (N_20105,N_16189,N_16108);
and U20106 (N_20106,N_16632,N_15538);
xnor U20107 (N_20107,N_19290,N_16721);
or U20108 (N_20108,N_16353,N_19010);
nand U20109 (N_20109,N_19993,N_19151);
or U20110 (N_20110,N_15525,N_15572);
nor U20111 (N_20111,N_15252,N_19449);
nor U20112 (N_20112,N_15173,N_17812);
and U20113 (N_20113,N_15559,N_18404);
nor U20114 (N_20114,N_16710,N_19232);
nor U20115 (N_20115,N_17326,N_18193);
and U20116 (N_20116,N_15636,N_18988);
nor U20117 (N_20117,N_15332,N_17915);
and U20118 (N_20118,N_18166,N_18547);
or U20119 (N_20119,N_19196,N_16949);
or U20120 (N_20120,N_15773,N_17393);
xnor U20121 (N_20121,N_17169,N_17573);
nor U20122 (N_20122,N_15481,N_19287);
nor U20123 (N_20123,N_17314,N_18520);
nand U20124 (N_20124,N_17445,N_15685);
and U20125 (N_20125,N_15000,N_19678);
nand U20126 (N_20126,N_18019,N_15991);
and U20127 (N_20127,N_18493,N_15679);
and U20128 (N_20128,N_16619,N_18661);
nor U20129 (N_20129,N_16259,N_19826);
and U20130 (N_20130,N_19159,N_19341);
or U20131 (N_20131,N_17752,N_17996);
and U20132 (N_20132,N_17371,N_18259);
nor U20133 (N_20133,N_18687,N_16442);
nor U20134 (N_20134,N_16204,N_17217);
and U20135 (N_20135,N_18206,N_17348);
nor U20136 (N_20136,N_15713,N_19050);
nand U20137 (N_20137,N_18012,N_19349);
or U20138 (N_20138,N_16522,N_15848);
or U20139 (N_20139,N_16069,N_15518);
nand U20140 (N_20140,N_17936,N_17533);
nor U20141 (N_20141,N_19395,N_17489);
nor U20142 (N_20142,N_19728,N_15906);
nor U20143 (N_20143,N_15736,N_18028);
or U20144 (N_20144,N_16603,N_16480);
nor U20145 (N_20145,N_16928,N_19557);
nand U20146 (N_20146,N_17823,N_18635);
nand U20147 (N_20147,N_17295,N_16064);
or U20148 (N_20148,N_17825,N_19927);
and U20149 (N_20149,N_16459,N_15880);
and U20150 (N_20150,N_18597,N_17424);
nor U20151 (N_20151,N_17840,N_17232);
nor U20152 (N_20152,N_19979,N_18347);
nor U20153 (N_20153,N_15722,N_18697);
and U20154 (N_20154,N_15858,N_15426);
or U20155 (N_20155,N_19806,N_18397);
nor U20156 (N_20156,N_18982,N_17940);
or U20157 (N_20157,N_18595,N_19194);
nor U20158 (N_20158,N_16884,N_18401);
or U20159 (N_20159,N_19201,N_17218);
nand U20160 (N_20160,N_16719,N_16912);
nand U20161 (N_20161,N_16270,N_18224);
nand U20162 (N_20162,N_18184,N_17645);
or U20163 (N_20163,N_16830,N_19928);
nor U20164 (N_20164,N_19856,N_19894);
nor U20165 (N_20165,N_17874,N_16584);
nand U20166 (N_20166,N_18110,N_16226);
or U20167 (N_20167,N_16050,N_18862);
and U20168 (N_20168,N_16644,N_17836);
nand U20169 (N_20169,N_16378,N_17839);
nor U20170 (N_20170,N_16542,N_19846);
and U20171 (N_20171,N_15901,N_18261);
and U20172 (N_20172,N_16167,N_15793);
or U20173 (N_20173,N_17976,N_18773);
nand U20174 (N_20174,N_17762,N_18770);
nand U20175 (N_20175,N_19324,N_18768);
and U20176 (N_20176,N_16436,N_18423);
nand U20177 (N_20177,N_16605,N_17770);
and U20178 (N_20178,N_15478,N_16339);
nand U20179 (N_20179,N_16762,N_17155);
nor U20180 (N_20180,N_15315,N_15064);
nor U20181 (N_20181,N_15450,N_16717);
or U20182 (N_20182,N_18865,N_15719);
or U20183 (N_20183,N_16582,N_15879);
and U20184 (N_20184,N_19356,N_17561);
nor U20185 (N_20185,N_16789,N_18378);
nor U20186 (N_20186,N_15063,N_19696);
nand U20187 (N_20187,N_18854,N_18408);
or U20188 (N_20188,N_16836,N_16571);
nor U20189 (N_20189,N_18906,N_15714);
or U20190 (N_20190,N_17922,N_19776);
nand U20191 (N_20191,N_16311,N_16438);
and U20192 (N_20192,N_17401,N_18450);
and U20193 (N_20193,N_15894,N_16390);
nand U20194 (N_20194,N_15873,N_16279);
or U20195 (N_20195,N_16142,N_15921);
nor U20196 (N_20196,N_17198,N_16614);
nor U20197 (N_20197,N_16859,N_16406);
nand U20198 (N_20198,N_15394,N_16250);
or U20199 (N_20199,N_15025,N_17448);
and U20200 (N_20200,N_17794,N_19654);
nor U20201 (N_20201,N_18132,N_15129);
and U20202 (N_20202,N_15616,N_19748);
nor U20203 (N_20203,N_18396,N_15145);
nand U20204 (N_20204,N_17270,N_18667);
or U20205 (N_20205,N_18580,N_16796);
nor U20206 (N_20206,N_19016,N_16342);
or U20207 (N_20207,N_16564,N_15261);
nor U20208 (N_20208,N_15717,N_15663);
and U20209 (N_20209,N_15990,N_17032);
or U20210 (N_20210,N_18287,N_19398);
nor U20211 (N_20211,N_16829,N_18331);
or U20212 (N_20212,N_17651,N_17328);
or U20213 (N_20213,N_17769,N_17428);
or U20214 (N_20214,N_18322,N_15603);
nand U20215 (N_20215,N_18605,N_19167);
nand U20216 (N_20216,N_18674,N_19177);
nand U20217 (N_20217,N_16242,N_18112);
nand U20218 (N_20218,N_19835,N_18679);
or U20219 (N_20219,N_17946,N_16191);
nand U20220 (N_20220,N_15712,N_15865);
xnor U20221 (N_20221,N_15074,N_16078);
nor U20222 (N_20222,N_15267,N_19583);
and U20223 (N_20223,N_18850,N_15003);
nand U20224 (N_20224,N_15311,N_18839);
or U20225 (N_20225,N_16493,N_17159);
and U20226 (N_20226,N_17082,N_16421);
nor U20227 (N_20227,N_15859,N_16790);
nor U20228 (N_20228,N_19862,N_17433);
or U20229 (N_20229,N_16382,N_17526);
and U20230 (N_20230,N_15738,N_19981);
or U20231 (N_20231,N_16024,N_15776);
nand U20232 (N_20232,N_15205,N_16883);
nand U20233 (N_20233,N_17098,N_17056);
nand U20234 (N_20234,N_18663,N_16888);
nand U20235 (N_20235,N_16863,N_19864);
or U20236 (N_20236,N_16927,N_19005);
nor U20237 (N_20237,N_17015,N_19918);
nor U20238 (N_20238,N_15189,N_17067);
or U20239 (N_20239,N_15492,N_19714);
nor U20240 (N_20240,N_17285,N_16776);
nor U20241 (N_20241,N_16401,N_18717);
and U20242 (N_20242,N_15564,N_17455);
or U20243 (N_20243,N_19227,N_18135);
nor U20244 (N_20244,N_16249,N_15238);
nor U20245 (N_20245,N_16589,N_16947);
or U20246 (N_20246,N_19727,N_19160);
and U20247 (N_20247,N_15567,N_16514);
nor U20248 (N_20248,N_16546,N_19752);
nand U20249 (N_20249,N_16992,N_17064);
and U20250 (N_20250,N_18480,N_15602);
and U20251 (N_20251,N_15215,N_19963);
and U20252 (N_20252,N_19463,N_17879);
and U20253 (N_20253,N_15279,N_15711);
and U20254 (N_20254,N_18787,N_19560);
nand U20255 (N_20255,N_17058,N_17809);
nand U20256 (N_20256,N_17807,N_15384);
xor U20257 (N_20257,N_18394,N_15509);
nor U20258 (N_20258,N_18253,N_17207);
nand U20259 (N_20259,N_15624,N_15825);
nand U20260 (N_20260,N_16667,N_16697);
nor U20261 (N_20261,N_17452,N_15443);
and U20262 (N_20262,N_19683,N_15739);
and U20263 (N_20263,N_16322,N_17921);
nor U20264 (N_20264,N_15141,N_17030);
and U20265 (N_20265,N_17552,N_16865);
and U20266 (N_20266,N_16237,N_15073);
and U20267 (N_20267,N_16126,N_18505);
nand U20268 (N_20268,N_18751,N_19292);
nor U20269 (N_20269,N_16013,N_15237);
nand U20270 (N_20270,N_17346,N_19637);
and U20271 (N_20271,N_17160,N_19612);
xnor U20272 (N_20272,N_18897,N_18298);
and U20273 (N_20273,N_15229,N_16292);
or U20274 (N_20274,N_16951,N_17012);
nor U20275 (N_20275,N_19132,N_18526);
or U20276 (N_20276,N_17283,N_15275);
or U20277 (N_20277,N_15220,N_16545);
nand U20278 (N_20278,N_16723,N_19238);
nor U20279 (N_20279,N_18517,N_15159);
or U20280 (N_20280,N_15983,N_17780);
or U20281 (N_20281,N_15052,N_15797);
or U20282 (N_20282,N_15258,N_18150);
or U20283 (N_20283,N_16010,N_16425);
or U20284 (N_20284,N_17055,N_16294);
and U20285 (N_20285,N_18809,N_16964);
and U20286 (N_20286,N_15264,N_19023);
nor U20287 (N_20287,N_15397,N_17597);
nor U20288 (N_20288,N_15540,N_18676);
or U20289 (N_20289,N_15170,N_17543);
and U20290 (N_20290,N_19636,N_15150);
or U20291 (N_20291,N_17194,N_19185);
nand U20292 (N_20292,N_19249,N_17019);
nor U20293 (N_20293,N_16258,N_18617);
nor U20294 (N_20294,N_19623,N_15606);
or U20295 (N_20295,N_16680,N_17135);
and U20296 (N_20296,N_19175,N_18728);
and U20297 (N_20297,N_16929,N_15195);
or U20298 (N_20298,N_19073,N_18947);
nand U20299 (N_20299,N_15708,N_16117);
nor U20300 (N_20300,N_16186,N_19688);
nor U20301 (N_20301,N_19311,N_19985);
or U20302 (N_20302,N_19679,N_17759);
nand U20303 (N_20303,N_17258,N_18445);
nand U20304 (N_20304,N_19141,N_18569);
nand U20305 (N_20305,N_15032,N_18088);
or U20306 (N_20306,N_17634,N_16746);
nor U20307 (N_20307,N_15801,N_16356);
or U20308 (N_20308,N_16038,N_19992);
nor U20309 (N_20309,N_16278,N_19286);
nand U20310 (N_20310,N_15321,N_15556);
and U20311 (N_20311,N_18489,N_18941);
and U20312 (N_20312,N_16896,N_16007);
nor U20313 (N_20313,N_18197,N_15233);
and U20314 (N_20314,N_18822,N_16761);
nand U20315 (N_20315,N_19730,N_15455);
nand U20316 (N_20316,N_15764,N_15437);
and U20317 (N_20317,N_19074,N_15718);
or U20318 (N_20318,N_19487,N_18752);
nor U20319 (N_20319,N_17409,N_19359);
or U20320 (N_20320,N_16469,N_17379);
or U20321 (N_20321,N_19068,N_19416);
or U20322 (N_20322,N_18372,N_15916);
nor U20323 (N_20323,N_16235,N_17313);
nand U20324 (N_20324,N_15262,N_16567);
nor U20325 (N_20325,N_16337,N_17426);
nor U20326 (N_20326,N_15127,N_19042);
nor U20327 (N_20327,N_16984,N_15404);
or U20328 (N_20328,N_15263,N_17624);
and U20329 (N_20329,N_19582,N_15605);
and U20330 (N_20330,N_19814,N_18777);
nand U20331 (N_20331,N_17771,N_18811);
and U20332 (N_20332,N_17185,N_15245);
nand U20333 (N_20333,N_18502,N_19145);
or U20334 (N_20334,N_17721,N_15961);
and U20335 (N_20335,N_16478,N_15870);
nor U20336 (N_20336,N_16594,N_16638);
or U20337 (N_20337,N_16088,N_19500);
nor U20338 (N_20338,N_18943,N_18171);
nor U20339 (N_20339,N_15429,N_19469);
and U20340 (N_20340,N_17060,N_18734);
nor U20341 (N_20341,N_19378,N_15001);
or U20342 (N_20342,N_15885,N_19199);
and U20343 (N_20343,N_17876,N_18250);
and U20344 (N_20344,N_16335,N_15458);
nand U20345 (N_20345,N_18147,N_18286);
nor U20346 (N_20346,N_19233,N_17636);
nor U20347 (N_20347,N_15034,N_16405);
nor U20348 (N_20348,N_15439,N_16072);
and U20349 (N_20349,N_16135,N_19406);
and U20350 (N_20350,N_18884,N_19900);
nand U20351 (N_20351,N_18339,N_15909);
or U20352 (N_20352,N_15020,N_17711);
nor U20353 (N_20353,N_19126,N_16967);
nand U20354 (N_20354,N_18371,N_16657);
or U20355 (N_20355,N_15669,N_15590);
and U20356 (N_20356,N_16481,N_15899);
nand U20357 (N_20357,N_16653,N_17602);
and U20358 (N_20358,N_19765,N_16973);
nor U20359 (N_20359,N_15499,N_17478);
nand U20360 (N_20360,N_18653,N_19015);
and U20361 (N_20361,N_16736,N_17981);
nand U20362 (N_20362,N_18557,N_19741);
nor U20363 (N_20363,N_16160,N_15491);
nor U20364 (N_20364,N_16807,N_17008);
nor U20365 (N_20365,N_16841,N_17482);
and U20366 (N_20366,N_16170,N_17300);
nand U20367 (N_20367,N_19907,N_17399);
or U20368 (N_20368,N_17376,N_19011);
and U20369 (N_20369,N_15774,N_16641);
or U20370 (N_20370,N_19468,N_15382);
or U20371 (N_20371,N_19488,N_18488);
or U20372 (N_20372,N_17821,N_17892);
nand U20373 (N_20373,N_18103,N_19753);
or U20374 (N_20374,N_15345,N_18937);
and U20375 (N_20375,N_19067,N_17688);
xnor U20376 (N_20376,N_16316,N_18230);
xor U20377 (N_20377,N_19616,N_16096);
nor U20378 (N_20378,N_19497,N_16343);
nand U20379 (N_20379,N_15379,N_17087);
nor U20380 (N_20380,N_17534,N_17035);
nor U20381 (N_20381,N_15668,N_16960);
nand U20382 (N_20382,N_15386,N_19791);
or U20383 (N_20383,N_19135,N_16268);
or U20384 (N_20384,N_17389,N_16451);
or U20385 (N_20385,N_17919,N_15671);
and U20386 (N_20386,N_17254,N_19490);
nand U20387 (N_20387,N_19674,N_16113);
nor U20388 (N_20388,N_17620,N_15777);
and U20389 (N_20389,N_17692,N_17062);
nand U20390 (N_20390,N_19281,N_16755);
nand U20391 (N_20391,N_17971,N_18440);
or U20392 (N_20392,N_17789,N_16743);
and U20393 (N_20393,N_15219,N_16578);
nor U20394 (N_20394,N_15077,N_16592);
or U20395 (N_20395,N_15459,N_17527);
and U20396 (N_20396,N_15495,N_18903);
nor U20397 (N_20397,N_17354,N_17521);
nor U20398 (N_20398,N_18160,N_19841);
and U20399 (N_20399,N_17474,N_15530);
or U20400 (N_20400,N_18289,N_15059);
and U20401 (N_20401,N_16452,N_17223);
nand U20402 (N_20402,N_19917,N_18644);
or U20403 (N_20403,N_18336,N_19105);
nand U20404 (N_20404,N_18483,N_18931);
nand U20405 (N_20405,N_19353,N_15696);
and U20406 (N_20406,N_19842,N_19695);
or U20407 (N_20407,N_19411,N_18341);
nor U20408 (N_20408,N_17941,N_16940);
and U20409 (N_20409,N_19045,N_17180);
nor U20410 (N_20410,N_16781,N_19221);
nor U20411 (N_20411,N_19057,N_18098);
nand U20412 (N_20412,N_19946,N_19138);
nand U20413 (N_20413,N_19479,N_18583);
and U20414 (N_20414,N_15209,N_19451);
and U20415 (N_20415,N_17503,N_19409);
nand U20416 (N_20416,N_16369,N_17553);
nand U20417 (N_20417,N_18177,N_17483);
or U20418 (N_20418,N_19581,N_18040);
nor U20419 (N_20419,N_18352,N_19279);
and U20420 (N_20420,N_16751,N_19639);
nand U20421 (N_20421,N_18227,N_19439);
nand U20422 (N_20422,N_18541,N_16502);
or U20423 (N_20423,N_17037,N_15242);
or U20424 (N_20424,N_15053,N_19360);
and U20425 (N_20425,N_16419,N_16795);
and U20426 (N_20426,N_17631,N_15369);
and U20427 (N_20427,N_15920,N_18724);
or U20428 (N_20428,N_18835,N_16434);
nand U20429 (N_20429,N_17676,N_18958);
or U20430 (N_20430,N_18128,N_16428);
or U20431 (N_20431,N_16190,N_16246);
nor U20432 (N_20432,N_17495,N_16996);
nand U20433 (N_20433,N_15204,N_15732);
nand U20434 (N_20434,N_19383,N_18874);
or U20435 (N_20435,N_15178,N_16889);
or U20436 (N_20436,N_19455,N_16869);
nor U20437 (N_20437,N_19496,N_17211);
nand U20438 (N_20438,N_15863,N_15811);
nand U20439 (N_20439,N_16357,N_17935);
or U20440 (N_20440,N_15655,N_18965);
nor U20441 (N_20441,N_17950,N_18043);
nand U20442 (N_20442,N_18817,N_16934);
and U20443 (N_20443,N_16774,N_18882);
or U20444 (N_20444,N_15427,N_15787);
and U20445 (N_20445,N_18664,N_16747);
and U20446 (N_20446,N_16987,N_16082);
or U20447 (N_20447,N_19152,N_19458);
nand U20448 (N_20448,N_18618,N_19644);
or U20449 (N_20449,N_17493,N_18640);
or U20450 (N_20450,N_16989,N_16770);
and U20451 (N_20451,N_18689,N_16201);
nor U20452 (N_20452,N_19948,N_16349);
nand U20453 (N_20453,N_15888,N_19446);
or U20454 (N_20454,N_17820,N_19587);
nand U20455 (N_20455,N_17739,N_18570);
nor U20456 (N_20456,N_16044,N_19331);
nor U20457 (N_20457,N_17324,N_16718);
and U20458 (N_20458,N_19796,N_16547);
and U20459 (N_20459,N_19549,N_18561);
nor U20460 (N_20460,N_15822,N_16783);
nor U20461 (N_20461,N_15266,N_17933);
nand U20462 (N_20462,N_16909,N_15529);
nand U20463 (N_20463,N_18976,N_18099);
nor U20464 (N_20464,N_16660,N_17068);
or U20465 (N_20465,N_16352,N_15185);
or U20466 (N_20466,N_15339,N_17984);
nand U20467 (N_20467,N_18023,N_18969);
nand U20468 (N_20468,N_18825,N_17090);
and U20469 (N_20469,N_19402,N_17469);
nor U20470 (N_20470,N_17241,N_17910);
and U20471 (N_20471,N_17588,N_17375);
nand U20472 (N_20472,N_16129,N_18168);
and U20473 (N_20473,N_17303,N_16026);
and U20474 (N_20474,N_19112,N_17382);
nand U20475 (N_20475,N_15094,N_17992);
or U20476 (N_20476,N_19617,N_19556);
and U20477 (N_20477,N_18433,N_17041);
nor U20478 (N_20478,N_16599,N_15744);
nand U20479 (N_20479,N_18395,N_17078);
or U20480 (N_20480,N_19615,N_15436);
nand U20481 (N_20481,N_17989,N_15791);
and U20482 (N_20482,N_16656,N_15918);
nor U20483 (N_20483,N_19541,N_19210);
and U20484 (N_20484,N_16997,N_19022);
nor U20485 (N_20485,N_19664,N_17488);
nand U20486 (N_20486,N_18072,N_16346);
nand U20487 (N_20487,N_19951,N_19914);
nand U20488 (N_20488,N_19143,N_16474);
xor U20489 (N_20489,N_15114,N_19689);
and U20490 (N_20490,N_19829,N_16106);
or U20491 (N_20491,N_17234,N_16885);
and U20492 (N_20492,N_17325,N_18306);
nand U20493 (N_20493,N_16566,N_16409);
nor U20494 (N_20494,N_19825,N_17163);
nand U20495 (N_20495,N_17361,N_19875);
and U20496 (N_20496,N_16471,N_16152);
nand U20497 (N_20497,N_17684,N_19080);
or U20498 (N_20498,N_17181,N_15039);
nor U20499 (N_20499,N_19176,N_15402);
or U20500 (N_20500,N_19669,N_19342);
nand U20501 (N_20501,N_17102,N_17208);
nand U20502 (N_20502,N_17251,N_17465);
or U20503 (N_20503,N_16284,N_18466);
nand U20504 (N_20504,N_19770,N_19306);
and U20505 (N_20505,N_18469,N_19584);
or U20506 (N_20506,N_18592,N_19313);
nor U20507 (N_20507,N_18413,N_18393);
nor U20508 (N_20508,N_19253,N_17097);
and U20509 (N_20509,N_19116,N_17242);
nor U20510 (N_20510,N_18024,N_16341);
nor U20511 (N_20511,N_17914,N_15223);
or U20512 (N_20512,N_19048,N_17316);
or U20513 (N_20513,N_18984,N_17168);
nand U20514 (N_20514,N_17988,N_17682);
or U20515 (N_20515,N_16440,N_17993);
or U20516 (N_20516,N_16093,N_16629);
nor U20517 (N_20517,N_17898,N_17509);
nor U20518 (N_20518,N_17813,N_15103);
nand U20519 (N_20519,N_16663,N_18696);
xor U20520 (N_20520,N_16351,N_17105);
or U20521 (N_20521,N_15289,N_19943);
and U20522 (N_20522,N_16364,N_18879);
and U20523 (N_20523,N_18741,N_19813);
nor U20524 (N_20524,N_15995,N_15473);
and U20525 (N_20525,N_19327,N_18533);
and U20526 (N_20526,N_15098,N_17972);
and U20527 (N_20527,N_19231,N_19921);
or U20528 (N_20528,N_18022,N_15850);
nand U20529 (N_20529,N_15519,N_16703);
and U20530 (N_20530,N_15667,N_16931);
or U20531 (N_20531,N_15432,N_18824);
and U20532 (N_20532,N_19498,N_17043);
or U20533 (N_20533,N_17608,N_18386);
nor U20534 (N_20534,N_17166,N_16740);
or U20535 (N_20535,N_17530,N_18549);
nor U20536 (N_20536,N_16187,N_18332);
nor U20537 (N_20537,N_16127,N_19332);
and U20538 (N_20538,N_18175,N_17479);
nand U20539 (N_20539,N_15417,N_18630);
nor U20540 (N_20540,N_17754,N_18448);
and U20541 (N_20541,N_16487,N_16631);
nand U20542 (N_20542,N_17544,N_17909);
nor U20543 (N_20543,N_19106,N_17384);
nand U20544 (N_20544,N_15939,N_17931);
and U20545 (N_20545,N_17673,N_17617);
or U20546 (N_20546,N_16302,N_19586);
nand U20547 (N_20547,N_19973,N_18546);
nand U20548 (N_20548,N_19673,N_18161);
and U20549 (N_20549,N_17390,N_17427);
and U20550 (N_20550,N_17201,N_15087);
nand U20551 (N_20551,N_17350,N_18708);
nor U20552 (N_20552,N_17512,N_19899);
and U20553 (N_20553,N_15820,N_15212);
nand U20554 (N_20554,N_18144,N_18131);
and U20555 (N_20555,N_18079,N_18065);
or U20556 (N_20556,N_19876,N_16590);
nor U20557 (N_20557,N_19995,N_18819);
and U20558 (N_20558,N_15306,N_16433);
and U20559 (N_20559,N_16059,N_15552);
nand U20560 (N_20560,N_15839,N_19697);
and U20561 (N_20561,N_17942,N_18648);
nand U20562 (N_20562,N_15589,N_15115);
and U20563 (N_20563,N_18654,N_19565);
and U20564 (N_20564,N_19737,N_19168);
nand U20565 (N_20565,N_15090,N_19924);
nand U20566 (N_20566,N_19323,N_18148);
nand U20567 (N_20567,N_19745,N_18241);
and U20568 (N_20568,N_15962,N_17686);
and U20569 (N_20569,N_15778,N_19404);
nor U20570 (N_20570,N_18189,N_15779);
or U20571 (N_20571,N_15514,N_18463);
and U20572 (N_20572,N_16085,N_15194);
nor U20573 (N_20573,N_17985,N_19443);
nand U20574 (N_20574,N_15006,N_17829);
or U20575 (N_20575,N_17726,N_19653);
nor U20576 (N_20576,N_17405,N_18139);
nor U20577 (N_20577,N_15933,N_18344);
nor U20578 (N_20578,N_17546,N_19289);
and U20579 (N_20579,N_15631,N_17858);
and U20580 (N_20580,N_19179,N_18452);
nor U20581 (N_20581,N_15016,N_19103);
nand U20582 (N_20582,N_18153,N_17562);
nand U20583 (N_20583,N_17773,N_19710);
or U20584 (N_20584,N_19923,N_16900);
or U20585 (N_20585,N_15944,N_16465);
or U20586 (N_20586,N_16205,N_19125);
nand U20587 (N_20587,N_15381,N_19299);
nand U20588 (N_20588,N_19977,N_15903);
or U20589 (N_20589,N_15707,N_17963);
and U20590 (N_20590,N_15067,N_15451);
or U20591 (N_20591,N_19805,N_19808);
nor U20592 (N_20592,N_16001,N_18607);
and U20593 (N_20593,N_15336,N_17912);
nor U20594 (N_20594,N_16971,N_19206);
nor U20595 (N_20595,N_17681,N_19429);
or U20596 (N_20596,N_15011,N_19320);
or U20597 (N_20597,N_18149,N_16576);
and U20598 (N_20598,N_19599,N_15444);
or U20599 (N_20599,N_17171,N_18550);
or U20600 (N_20600,N_16503,N_15945);
nand U20601 (N_20601,N_15044,N_19364);
nor U20602 (N_20602,N_17498,N_15953);
nand U20603 (N_20603,N_16798,N_17657);
nor U20604 (N_20604,N_19460,N_17618);
and U20605 (N_20605,N_17591,N_15307);
or U20606 (N_20606,N_16846,N_16831);
nor U20607 (N_20607,N_17763,N_18789);
or U20608 (N_20608,N_15154,N_16286);
nor U20609 (N_20609,N_16468,N_18594);
nand U20610 (N_20610,N_18140,N_19118);
nand U20611 (N_20611,N_16837,N_16220);
or U20612 (N_20612,N_16785,N_18494);
nand U20613 (N_20613,N_18312,N_16388);
and U20614 (N_20614,N_18892,N_15425);
nand U20615 (N_20615,N_16475,N_15171);
and U20616 (N_20616,N_19114,N_19687);
nand U20617 (N_20617,N_17297,N_18170);
and U20618 (N_20618,N_15541,N_18904);
and U20619 (N_20619,N_18270,N_16042);
or U20620 (N_20620,N_17464,N_15320);
or U20621 (N_20621,N_17668,N_17407);
nor U20622 (N_20622,N_18702,N_19550);
nor U20623 (N_20623,N_19975,N_18226);
nor U20624 (N_20624,N_18338,N_15095);
or U20625 (N_20625,N_16528,N_16612);
or U20626 (N_20626,N_18478,N_19124);
nand U20627 (N_20627,N_19735,N_19881);
nand U20628 (N_20628,N_17709,N_16714);
and U20629 (N_20629,N_18962,N_19109);
nand U20630 (N_20630,N_17640,N_17628);
nand U20631 (N_20631,N_17607,N_18998);
nor U20632 (N_20632,N_17366,N_15890);
and U20633 (N_20633,N_16527,N_18519);
and U20634 (N_20634,N_16505,N_16454);
nor U20635 (N_20635,N_18802,N_19930);
or U20636 (N_20636,N_18553,N_16304);
xor U20637 (N_20637,N_17785,N_16060);
or U20638 (N_20638,N_15852,N_17106);
nand U20639 (N_20639,N_19534,N_18510);
or U20640 (N_20640,N_17450,N_15131);
nand U20641 (N_20641,N_18158,N_18536);
or U20642 (N_20642,N_16058,N_16266);
or U20643 (N_20643,N_17900,N_17968);
nand U20644 (N_20644,N_17793,N_19733);
nor U20645 (N_20645,N_17235,N_18125);
and U20646 (N_20646,N_17749,N_19997);
nor U20647 (N_20647,N_16397,N_15027);
or U20648 (N_20648,N_16192,N_19926);
nor U20649 (N_20649,N_19304,N_16924);
and U20650 (N_20650,N_18933,N_17432);
nand U20651 (N_20651,N_15490,N_17536);
nor U20652 (N_20652,N_19691,N_16417);
nand U20653 (N_20653,N_15536,N_19393);
or U20654 (N_20654,N_16470,N_15108);
nor U20655 (N_20655,N_15188,N_18497);
nor U20656 (N_20656,N_16043,N_15584);
nand U20657 (N_20657,N_18025,N_15116);
nor U20658 (N_20658,N_18133,N_19317);
nand U20659 (N_20659,N_19685,N_19062);
and U20660 (N_20660,N_17388,N_17265);
and U20661 (N_20661,N_15172,N_19037);
or U20662 (N_20662,N_16702,N_19431);
nand U20663 (N_20663,N_19508,N_16136);
or U20664 (N_20664,N_16618,N_18109);
nand U20665 (N_20665,N_16979,N_16856);
or U20666 (N_20666,N_19059,N_18720);
and U20667 (N_20667,N_17016,N_15482);
or U20668 (N_20668,N_19819,N_19056);
nor U20669 (N_20669,N_18426,N_19991);
nor U20670 (N_20670,N_15061,N_18380);
nand U20671 (N_20671,N_19285,N_16553);
or U20672 (N_20672,N_18849,N_16611);
or U20673 (N_20673,N_18070,N_19091);
or U20674 (N_20674,N_16509,N_19896);
nand U20675 (N_20675,N_15021,N_18283);
and U20676 (N_20676,N_17872,N_15558);
nand U20677 (N_20677,N_15002,N_15963);
or U20678 (N_20678,N_19643,N_19911);
nand U20679 (N_20679,N_18756,N_15226);
nand U20680 (N_20680,N_15388,N_18710);
nand U20681 (N_20681,N_16670,N_19161);
nor U20682 (N_20682,N_17095,N_17449);
or U20683 (N_20683,N_19193,N_18002);
or U20684 (N_20684,N_17116,N_19115);
nor U20685 (N_20685,N_17962,N_15010);
nand U20686 (N_20686,N_18467,N_17767);
and U20687 (N_20687,N_15065,N_15721);
and U20688 (N_20688,N_19605,N_16306);
nor U20689 (N_20689,N_18471,N_16876);
nand U20690 (N_20690,N_17480,N_16325);
and U20691 (N_20691,N_19839,N_17613);
nor U20692 (N_20692,N_15770,N_19055);
xnor U20693 (N_20693,N_16998,N_16529);
and U20694 (N_20694,N_17658,N_16832);
nor U20695 (N_20695,N_17685,N_15573);
and U20696 (N_20696,N_18246,N_18236);
nor U20697 (N_20697,N_19761,N_15686);
or U20698 (N_20698,N_19271,N_19379);
nor U20699 (N_20699,N_19163,N_18247);
nand U20700 (N_20700,N_17502,N_19511);
nand U20701 (N_20701,N_15372,N_16414);
nor U20702 (N_20702,N_15463,N_15562);
nor U20703 (N_20703,N_17511,N_17786);
nor U20704 (N_20704,N_17085,N_17093);
and U20705 (N_20705,N_18454,N_17118);
and U20706 (N_20706,N_18899,N_16683);
nor U20707 (N_20707,N_17013,N_17716);
or U20708 (N_20708,N_17378,N_15942);
nor U20709 (N_20709,N_17227,N_17923);
or U20710 (N_20710,N_17701,N_16238);
nor U20711 (N_20711,N_17387,N_16630);
nand U20712 (N_20712,N_15331,N_18470);
nand U20713 (N_20713,N_15768,N_17459);
and U20714 (N_20714,N_17299,N_16247);
or U20715 (N_20715,N_17939,N_19734);
or U20716 (N_20716,N_15142,N_17071);
nor U20717 (N_20717,N_17675,N_18037);
nor U20718 (N_20718,N_15222,N_17273);
or U20719 (N_20719,N_18412,N_16178);
and U20720 (N_20720,N_16957,N_18660);
nor U20721 (N_20721,N_19265,N_15485);
nand U20722 (N_20722,N_18085,N_17508);
and U20723 (N_20723,N_16328,N_15276);
and U20724 (N_20724,N_16915,N_19140);
nand U20725 (N_20725,N_19959,N_18758);
nor U20726 (N_20726,N_17137,N_18706);
nor U20727 (N_20727,N_17307,N_19656);
and U20728 (N_20728,N_17583,N_18766);
and U20729 (N_20729,N_15651,N_19272);
nand U20730 (N_20730,N_19006,N_18961);
nand U20731 (N_20731,N_15416,N_16150);
or U20732 (N_20732,N_16153,N_15965);
nand U20733 (N_20733,N_17304,N_18539);
nand U20734 (N_20734,N_16608,N_18754);
or U20735 (N_20735,N_19302,N_16051);
and U20736 (N_20736,N_17738,N_18381);
or U20737 (N_20737,N_17202,N_19408);
and U20738 (N_20738,N_15387,N_18692);
nand U20739 (N_20739,N_17730,N_16647);
and U20740 (N_20740,N_18633,N_15976);
or U20741 (N_20741,N_15399,N_19754);
or U20742 (N_20742,N_15472,N_19912);
or U20743 (N_20743,N_18968,N_17880);
and U20744 (N_20744,N_16444,N_15956);
nand U20745 (N_20745,N_17717,N_19343);
nor U20746 (N_20746,N_17854,N_17866);
or U20747 (N_20747,N_18365,N_19482);
and U20748 (N_20748,N_16119,N_19478);
nor U20749 (N_20749,N_15912,N_16519);
and U20750 (N_20750,N_16639,N_18512);
nor U20751 (N_20751,N_19686,N_18430);
or U20752 (N_20752,N_15043,N_17851);
nor U20753 (N_20753,N_15581,N_19635);
nand U20754 (N_20754,N_17293,N_18258);
nand U20755 (N_20755,N_17841,N_19779);
nand U20756 (N_20756,N_15288,N_19354);
or U20757 (N_20757,N_18377,N_19603);
or U20758 (N_20758,N_19020,N_17321);
nor U20759 (N_20759,N_18182,N_17664);
nand U20760 (N_20760,N_18513,N_16464);
and U20761 (N_20761,N_16559,N_17973);
and U20762 (N_20762,N_17486,N_18614);
nor U20763 (N_20763,N_16068,N_18925);
and U20764 (N_20764,N_15055,N_17236);
nor U20765 (N_20765,N_17302,N_15560);
and U20766 (N_20766,N_15075,N_17772);
nand U20767 (N_20767,N_18540,N_15695);
or U20768 (N_20768,N_16675,N_16336);
or U20769 (N_20769,N_19830,N_18468);
nor U20770 (N_20770,N_17949,N_17999);
or U20771 (N_20771,N_15782,N_19662);
and U20772 (N_20772,N_16431,N_16950);
or U20773 (N_20773,N_19525,N_17551);
or U20774 (N_20774,N_16219,N_18130);
nand U20775 (N_20775,N_16439,N_19377);
and U20776 (N_20776,N_16161,N_15740);
or U20777 (N_20777,N_19013,N_18083);
or U20778 (N_20778,N_15471,N_15601);
and U20779 (N_20779,N_18495,N_18711);
xor U20780 (N_20780,N_18039,N_15097);
or U20781 (N_20781,N_17395,N_19523);
nor U20782 (N_20782,N_16083,N_18069);
nand U20783 (N_20783,N_19775,N_19580);
or U20784 (N_20784,N_16695,N_16842);
nand U20785 (N_20785,N_18188,N_17959);
and U20786 (N_20786,N_18325,N_16651);
nand U20787 (N_20787,N_15517,N_19700);
nor U20788 (N_20788,N_16634,N_17059);
or U20789 (N_20789,N_18651,N_19241);
and U20790 (N_20790,N_18649,N_16504);
nand U20791 (N_20791,N_15521,N_18212);
or U20792 (N_20792,N_17490,N_15966);
nor U20793 (N_20793,N_17961,N_19502);
nand U20794 (N_20794,N_18054,N_18832);
or U20795 (N_20795,N_19305,N_15769);
or U20796 (N_20796,N_18889,N_16199);
nand U20797 (N_20797,N_19382,N_18808);
and U20798 (N_20798,N_16491,N_15843);
and U20799 (N_20799,N_16035,N_15138);
nor U20800 (N_20800,N_16792,N_18194);
and U20801 (N_20801,N_15346,N_17210);
or U20802 (N_20802,N_19270,N_18263);
or U20803 (N_20803,N_15897,N_19095);
nand U20804 (N_20804,N_15620,N_16895);
and U20805 (N_20805,N_16610,N_15329);
and U20806 (N_20806,N_19248,N_19625);
nor U20807 (N_20807,N_16348,N_17473);
nor U20808 (N_20808,N_17182,N_19465);
nand U20809 (N_20809,N_15368,N_18564);
nor U20810 (N_20810,N_16709,N_18068);
and U20811 (N_20811,N_18004,N_18639);
or U20812 (N_20812,N_18044,N_19983);
nor U20813 (N_20813,N_19442,N_17970);
nor U20814 (N_20814,N_17280,N_18299);
nor U20815 (N_20815,N_18006,N_18216);
and U20816 (N_20816,N_17817,N_16496);
or U20817 (N_20817,N_16075,N_19189);
or U20818 (N_20818,N_19804,N_19100);
or U20819 (N_20819,N_18684,N_17535);
nand U20820 (N_20820,N_16495,N_18558);
nor U20821 (N_20821,N_16794,N_19633);
nand U20822 (N_20822,N_19234,N_16029);
nand U20823 (N_20823,N_17885,N_15134);
or U20824 (N_20824,N_19444,N_16367);
xnor U20825 (N_20825,N_15751,N_16813);
nor U20826 (N_20826,N_15643,N_16012);
nand U20827 (N_20827,N_17156,N_17920);
and U20828 (N_20828,N_19613,N_19239);
nand U20829 (N_20829,N_17322,N_19107);
or U20830 (N_20830,N_17080,N_15723);
nand U20831 (N_20831,N_18629,N_17908);
or U20832 (N_20832,N_17878,N_15809);
or U20833 (N_20833,N_17955,N_19301);
nand U20834 (N_20834,N_17446,N_19812);
nand U20835 (N_20835,N_17609,N_16224);
or U20836 (N_20836,N_18042,N_17267);
nor U20837 (N_20837,N_18573,N_15089);
nand U20838 (N_20838,N_15255,N_18077);
and U20839 (N_20839,N_15265,N_15952);
nand U20840 (N_20840,N_16875,N_18940);
or U20841 (N_20841,N_18658,N_15414);
or U20842 (N_20842,N_17103,N_16974);
and U20843 (N_20843,N_19939,N_18441);
and U20844 (N_20844,N_17590,N_17121);
nor U20845 (N_20845,N_16968,N_18622);
nand U20846 (N_20846,N_19832,N_16206);
nor U20847 (N_20847,N_18875,N_17094);
nand U20848 (N_20848,N_15271,N_19242);
nand U20849 (N_20849,N_17006,N_18208);
nor U20850 (N_20850,N_18818,N_17604);
or U20851 (N_20851,N_17282,N_19381);
nand U20852 (N_20852,N_16398,N_15467);
nand U20853 (N_20853,N_15259,N_17117);
nor U20854 (N_20854,N_17727,N_19218);
nand U20855 (N_20855,N_16615,N_18733);
nor U20856 (N_20856,N_18278,N_17458);
or U20857 (N_20857,N_16548,N_19950);
nand U20858 (N_20858,N_19211,N_19528);
nor U20859 (N_20859,N_19494,N_18213);
or U20860 (N_20860,N_17330,N_18485);
nor U20861 (N_20861,N_15474,N_15254);
nor U20862 (N_20862,N_16103,N_17081);
or U20863 (N_20863,N_19085,N_15153);
nor U20864 (N_20864,N_18612,N_19003);
nand U20865 (N_20865,N_15698,N_18210);
nand U20866 (N_20866,N_16805,N_16664);
nor U20867 (N_20867,N_18857,N_18350);
nor U20868 (N_20868,N_16772,N_17170);
and U20869 (N_20869,N_18292,N_15224);
nand U20870 (N_20870,N_18816,N_15151);
nand U20871 (N_20871,N_16435,N_15690);
and U20872 (N_20872,N_16706,N_16966);
and U20873 (N_20873,N_19236,N_18214);
nand U20874 (N_20874,N_15130,N_15203);
nor U20875 (N_20875,N_18030,N_18453);
or U20876 (N_20876,N_16402,N_18672);
or U20877 (N_20877,N_16457,N_19053);
or U20878 (N_20878,N_17414,N_19676);
or U20879 (N_20879,N_18560,N_18265);
and U20880 (N_20880,N_17422,N_19561);
nand U20881 (N_20881,N_15922,N_17750);
or U20882 (N_20882,N_16624,N_15702);
and U20883 (N_20883,N_15729,N_15555);
nor U20884 (N_20884,N_17683,N_18319);
and U20885 (N_20885,N_16687,N_17927);
or U20886 (N_20886,N_18382,N_17296);
or U20887 (N_20887,N_18199,N_18238);
nand U20888 (N_20888,N_18121,N_16033);
xor U20889 (N_20889,N_19828,N_19858);
or U20890 (N_20890,N_16385,N_18279);
or U20891 (N_20891,N_19181,N_15585);
nand U20892 (N_20892,N_15756,N_17268);
and U20893 (N_20893,N_15406,N_17264);
or U20894 (N_20894,N_19553,N_17252);
nor U20895 (N_20895,N_16995,N_16383);
and U20896 (N_20896,N_18886,N_18503);
nand U20897 (N_20897,N_18231,N_16686);
or U20898 (N_20898,N_16045,N_19200);
nor U20899 (N_20899,N_17691,N_17053);
or U20900 (N_20900,N_18544,N_18106);
nand U20901 (N_20901,N_16130,N_15337);
nand U20902 (N_20902,N_19040,N_19136);
nor U20903 (N_20903,N_17089,N_17600);
nor U20904 (N_20904,N_18491,N_17842);
nand U20905 (N_20905,N_18535,N_16858);
and U20906 (N_20906,N_17625,N_18104);
nor U20907 (N_20907,N_18712,N_15613);
or U20908 (N_20908,N_17643,N_19682);
or U20909 (N_20909,N_15637,N_15528);
nand U20910 (N_20910,N_17958,N_18745);
and U20911 (N_20911,N_18017,N_16216);
nand U20912 (N_20912,N_19766,N_16313);
or U20913 (N_20913,N_19785,N_19759);
or U20914 (N_20914,N_17441,N_15042);
and U20915 (N_20915,N_17351,N_19207);
nand U20916 (N_20916,N_17203,N_16715);
nor U20917 (N_20917,N_15914,N_17826);
and U20918 (N_20918,N_15828,N_15084);
or U20919 (N_20919,N_17896,N_17832);
or U20920 (N_20920,N_19866,N_19361);
or U20921 (N_20921,N_19310,N_17246);
and U20922 (N_20922,N_19293,N_19447);
or U20923 (N_20923,N_17362,N_16039);
nor U20924 (N_20924,N_18093,N_19263);
and U20925 (N_20925,N_15826,N_15823);
or U20926 (N_20926,N_17569,N_16768);
and U20927 (N_20927,N_19256,N_15881);
xnor U20928 (N_20928,N_19032,N_15968);
nand U20929 (N_20929,N_17788,N_17494);
nor U20930 (N_20930,N_16466,N_15929);
nand U20931 (N_20931,N_18005,N_18971);
or U20932 (N_20932,N_18930,N_18081);
nand U20933 (N_20933,N_16563,N_19655);
nand U20934 (N_20934,N_15028,N_17266);
xor U20935 (N_20935,N_17753,N_16749);
or U20936 (N_20936,N_18888,N_17873);
or U20937 (N_20937,N_15278,N_17868);
or U20938 (N_20938,N_18082,N_15359);
nand U20939 (N_20939,N_17072,N_19061);
nor U20940 (N_20940,N_19960,N_15819);
and U20941 (N_20941,N_18716,N_18358);
nor U20942 (N_20942,N_18385,N_16473);
nor U20943 (N_20943,N_17065,N_17746);
nand U20944 (N_20944,N_16080,N_17579);
and U20945 (N_20945,N_16244,N_19345);
nor U20946 (N_20946,N_19099,N_17937);
nor U20947 (N_20947,N_18033,N_16769);
nor U20948 (N_20948,N_18007,N_18424);
nand U20949 (N_20949,N_18455,N_17063);
nand U20950 (N_20950,N_15814,N_17756);
nor U20951 (N_20951,N_16006,N_15632);
or U20952 (N_20952,N_18444,N_15941);
nand U20953 (N_20953,N_15849,N_19300);
or U20954 (N_20954,N_18859,N_16911);
or U20955 (N_20955,N_18388,N_17517);
nor U20956 (N_20956,N_18522,N_19504);
nand U20957 (N_20957,N_17837,N_17702);
and U20958 (N_20958,N_19827,N_16560);
nor U20959 (N_20959,N_19988,N_16289);
and U20960 (N_20960,N_17421,N_16175);
nand U20961 (N_20961,N_17694,N_18297);
nand U20962 (N_20962,N_16453,N_18329);
or U20963 (N_20963,N_19671,N_17442);
and U20964 (N_20964,N_15004,N_15269);
or U20965 (N_20965,N_15421,N_19554);
nand U20966 (N_20966,N_17475,N_17714);
and U20967 (N_20967,N_15048,N_19389);
or U20968 (N_20968,N_16598,N_15405);
nand U20969 (N_20969,N_19762,N_17356);
and U20970 (N_20970,N_17671,N_18235);
xnor U20971 (N_20971,N_17983,N_19243);
nand U20972 (N_20972,N_16555,N_18232);
or U20973 (N_20973,N_18829,N_15176);
nand U20974 (N_20974,N_18237,N_17110);
or U20975 (N_20975,N_15681,N_19984);
or U20976 (N_20976,N_17568,N_16355);
nor U20977 (N_20977,N_16811,N_18064);
and U20978 (N_20978,N_16182,N_18008);
nor U20979 (N_20979,N_15924,N_16828);
or U20980 (N_20980,N_17757,N_15547);
nand U20981 (N_20981,N_17644,N_17599);
nand U20982 (N_20982,N_19982,N_15597);
nor U20983 (N_20983,N_17518,N_15595);
nor U20984 (N_20984,N_19568,N_15855);
nor U20985 (N_20985,N_19276,N_18376);
or U20986 (N_20986,N_18366,N_19472);
and U20987 (N_20987,N_15476,N_17928);
and U20988 (N_20988,N_18234,N_19322);
or U20989 (N_20989,N_16260,N_16649);
and U20990 (N_20990,N_16447,N_19089);
xor U20991 (N_20991,N_19108,N_17444);
or U20992 (N_20992,N_17224,N_15750);
nand U20993 (N_20993,N_17134,N_19155);
or U20994 (N_20994,N_18508,N_17333);
nand U20995 (N_20995,N_19569,N_15993);
nor U20996 (N_20996,N_17687,N_18999);
or U20997 (N_20997,N_15070,N_16874);
nand U20998 (N_20998,N_16424,N_18567);
and U20999 (N_20999,N_17463,N_18119);
nor U21000 (N_21000,N_15700,N_17831);
and U21001 (N_21001,N_16163,N_15692);
or U21002 (N_21002,N_18146,N_19909);
nor U21003 (N_21003,N_16840,N_16738);
and U21004 (N_21004,N_17036,N_19543);
nor U21005 (N_21005,N_15082,N_17069);
nor U21006 (N_21006,N_18534,N_18791);
or U21007 (N_21007,N_18615,N_16120);
nor U21008 (N_21008,N_16637,N_17101);
and U21009 (N_21009,N_15904,N_16062);
and U21010 (N_21010,N_18219,N_18665);
and U21011 (N_21011,N_15391,N_18681);
or U21012 (N_21012,N_16234,N_15720);
or U21013 (N_21013,N_16020,N_15949);
nor U21014 (N_21014,N_15900,N_18885);
or U21015 (N_21015,N_19224,N_18559);
or U21016 (N_21016,N_18313,N_18113);
nand U21017 (N_21017,N_18272,N_18562);
nor U21018 (N_21018,N_15621,N_18511);
nand U21019 (N_21019,N_15504,N_15674);
and U21020 (N_21020,N_18746,N_16360);
and U21021 (N_21021,N_15121,N_17733);
or U21022 (N_21022,N_15759,N_18122);
nor U21023 (N_21023,N_18342,N_16507);
nand U21024 (N_21024,N_18102,N_16461);
nor U21025 (N_21025,N_17665,N_15907);
or U21026 (N_21026,N_17633,N_15433);
and U21027 (N_21027,N_15335,N_17337);
or U21028 (N_21028,N_19601,N_19001);
or U21029 (N_21029,N_15935,N_15979);
or U21030 (N_21030,N_19743,N_18990);
nand U21031 (N_21031,N_16955,N_18391);
xnor U21032 (N_21032,N_19158,N_19968);
nand U21033 (N_21033,N_15236,N_17806);
or U21034 (N_21034,N_17099,N_19720);
nand U21035 (N_21035,N_15169,N_18574);
or U21036 (N_21036,N_18736,N_15693);
and U21037 (N_21037,N_19432,N_17039);
nand U21038 (N_21038,N_19595,N_18281);
nor U21039 (N_21039,N_19367,N_19063);
nor U21040 (N_21040,N_15553,N_17277);
or U21041 (N_21041,N_18952,N_15520);
nand U21042 (N_21042,N_17986,N_19259);
and U21043 (N_21043,N_17798,N_16123);
nor U21044 (N_21044,N_18518,N_19640);
and U21045 (N_21045,N_17529,N_19087);
and U21046 (N_21046,N_15507,N_17706);
and U21047 (N_21047,N_16969,N_18403);
or U21048 (N_21048,N_19454,N_16802);
nand U21049 (N_21049,N_19481,N_17143);
and U21050 (N_21050,N_17696,N_17429);
nand U21051 (N_21051,N_16671,N_17434);
and U21052 (N_21052,N_16005,N_16374);
nor U21053 (N_21053,N_17849,N_16943);
nor U21054 (N_21054,N_18779,N_18507);
and U21055 (N_21055,N_17863,N_17086);
nand U21056 (N_21056,N_15792,N_18305);
nand U21057 (N_21057,N_18293,N_19967);
nand U21058 (N_21058,N_18326,N_18406);
and U21059 (N_21059,N_17172,N_19046);
and U21060 (N_21060,N_15876,N_15291);
and U21061 (N_21061,N_19729,N_19747);
nor U21062 (N_21062,N_19934,N_19575);
or U21063 (N_21063,N_19957,N_19713);
nor U21064 (N_21064,N_15634,N_19235);
nor U21065 (N_21065,N_19892,N_18691);
or U21066 (N_21066,N_16847,N_15854);
nor U21067 (N_21067,N_17623,N_18145);
and U21068 (N_21068,N_18016,N_18799);
nand U21069 (N_21069,N_17392,N_16867);
nand U21070 (N_21070,N_15570,N_15309);
and U21071 (N_21071,N_16228,N_18531);
and U21072 (N_21072,N_18307,N_19614);
and U21073 (N_21073,N_15926,N_15198);
xnor U21074 (N_21074,N_19098,N_19414);
xor U21075 (N_21075,N_16275,N_18020);
or U21076 (N_21076,N_19672,N_19373);
or U21077 (N_21077,N_18360,N_19886);
nor U21078 (N_21078,N_15295,N_15370);
nor U21079 (N_21079,N_18924,N_19312);
nor U21080 (N_21080,N_18101,N_17834);
and U21081 (N_21081,N_17221,N_19843);
nor U21082 (N_21082,N_17500,N_16698);
nand U21083 (N_21083,N_19536,N_18443);
nor U21084 (N_21084,N_17760,N_17260);
nor U21085 (N_21085,N_18100,N_17987);
nand U21086 (N_21086,N_19486,N_16483);
and U21087 (N_21087,N_15930,N_19538);
nor U21088 (N_21088,N_17461,N_15524);
nor U21089 (N_21089,N_17109,N_17233);
or U21090 (N_21090,N_19422,N_18229);
nor U21091 (N_21091,N_19316,N_16506);
and U21092 (N_21092,N_17758,N_16445);
and U21093 (N_21093,N_18917,N_16739);
nor U21094 (N_21094,N_18009,N_19592);
or U21095 (N_21095,N_19358,N_15676);
nand U21096 (N_21096,N_18723,N_15600);
nor U21097 (N_21097,N_19882,N_15649);
nor U21098 (N_21098,N_16845,N_18870);
and U21099 (N_21099,N_19703,N_17632);
nand U21100 (N_21100,N_18749,N_17196);
nor U21101 (N_21101,N_18163,N_19908);
and U21102 (N_21102,N_17050,N_18273);
or U21103 (N_21103,N_19712,N_15300);
nand U21104 (N_21104,N_16241,N_15762);
and U21105 (N_21105,N_15675,N_16371);
and U21106 (N_21106,N_15807,N_18221);
nand U21107 (N_21107,N_15652,N_15771);
nor U21108 (N_21108,N_18375,N_17943);
nor U21109 (N_21109,N_16700,N_18014);
nor U21110 (N_21110,N_18589,N_17642);
or U21111 (N_21111,N_17964,N_18137);
or U21112 (N_21112,N_17865,N_17272);
or U21113 (N_21113,N_18439,N_19453);
or U21114 (N_21114,N_19631,N_19518);
nor U21115 (N_21115,N_16623,N_19448);
or U21116 (N_21116,N_16427,N_19786);
nor U21117 (N_21117,N_18256,N_16054);
or U21118 (N_21118,N_19399,N_19902);
and U21119 (N_21119,N_18905,N_15287);
nand U21120 (N_21120,N_16728,N_17889);
and U21121 (N_21121,N_18349,N_16310);
nand U21122 (N_21122,N_19916,N_19947);
or U21123 (N_21123,N_15548,N_18049);
and U21124 (N_21124,N_16236,N_18090);
and U21125 (N_21125,N_15757,N_18744);
nor U21126 (N_21126,N_16430,N_16826);
nand U21127 (N_21127,N_16801,N_18609);
and U21128 (N_21128,N_16513,N_15522);
or U21129 (N_21129,N_19315,N_15895);
nand U21130 (N_21130,N_18159,N_19611);
or U21131 (N_21131,N_17707,N_17385);
or U21132 (N_21132,N_16626,N_17138);
and U21133 (N_21133,N_16025,N_16843);
and U21134 (N_21134,N_18330,N_19570);
nor U21135 (N_21135,N_19166,N_18271);
nor U21136 (N_21136,N_18715,N_17830);
nand U21137 (N_21137,N_15325,N_15161);
nor U21138 (N_21138,N_16918,N_18719);
nand U21139 (N_21139,N_18827,N_18089);
nand U21140 (N_21140,N_16838,N_18356);
or U21141 (N_21141,N_19146,N_19865);
or U21142 (N_21142,N_18774,N_16850);
xnor U21143 (N_21143,N_17125,N_16799);
or U21144 (N_21144,N_16621,N_19578);
and U21145 (N_21145,N_17435,N_19197);
and U21146 (N_21146,N_18432,N_18353);
and U21147 (N_21147,N_15569,N_16158);
or U21148 (N_21148,N_19417,N_15164);
nand U21149 (N_21149,N_17383,N_15308);
or U21150 (N_21150,N_16110,N_18920);
nand U21151 (N_21151,N_16285,N_16361);
nor U21152 (N_21152,N_16668,N_15500);
and U21153 (N_21153,N_17484,N_16945);
and U21154 (N_21154,N_17111,N_16484);
and U21155 (N_21155,N_19369,N_16791);
nor U21156 (N_21156,N_15327,N_18218);
and U21157 (N_21157,N_18967,N_15633);
or U21158 (N_21158,N_19275,N_17368);
nor U21159 (N_21159,N_15014,N_16834);
nand U21160 (N_21160,N_19607,N_15608);
and U21161 (N_21161,N_15422,N_17199);
nand U21162 (N_21162,N_17177,N_15697);
or U21163 (N_21163,N_16212,N_17660);
nor U21164 (N_21164,N_17466,N_15978);
nor U21165 (N_21165,N_19180,N_16937);
and U21166 (N_21166,N_17710,N_17250);
or U21167 (N_21167,N_17052,N_15544);
nor U21168 (N_21168,N_16551,N_16307);
nor U21169 (N_21169,N_16601,N_15506);
and U21170 (N_21170,N_19415,N_17720);
nand U21171 (N_21171,N_19773,N_15754);
nand U21172 (N_21172,N_19328,N_19532);
nand U21173 (N_21173,N_17291,N_18727);
nor U21174 (N_21174,N_19213,N_16899);
and U21175 (N_21175,N_15350,N_16173);
or U21176 (N_21176,N_18473,N_16084);
and U21177 (N_21177,N_18737,N_15746);
nor U21178 (N_21178,N_17237,N_15323);
nand U21179 (N_21179,N_16403,N_15927);
xor U21180 (N_21180,N_15371,N_17761);
xor U21181 (N_21181,N_19069,N_18625);
nand U21182 (N_21182,N_18370,N_18701);
or U21183 (N_21183,N_17635,N_17593);
or U21184 (N_21184,N_15395,N_19036);
nand U21185 (N_21185,N_18634,N_17144);
and U21186 (N_21186,N_16354,N_17589);
or U21187 (N_21187,N_19278,N_18498);
and U21188 (N_21188,N_15737,N_15206);
and U21189 (N_21189,N_17548,N_16839);
and U21190 (N_21190,N_15767,N_19357);
xor U21191 (N_21191,N_18041,N_19172);
nor U21192 (N_21192,N_15030,N_19044);
nor U21193 (N_21193,N_16269,N_19215);
nand U21194 (N_21194,N_17402,N_19262);
and U21195 (N_21195,N_19034,N_17001);
nor U21196 (N_21196,N_15488,N_19385);
nand U21197 (N_21197,N_19188,N_15166);
and U21198 (N_21198,N_18418,N_17311);
nor U21199 (N_21199,N_17524,N_17418);
or U21200 (N_21200,N_19028,N_18075);
or U21201 (N_21201,N_17537,N_18792);
nor U21202 (N_21202,N_16812,N_17519);
and U21203 (N_21203,N_15512,N_16366);
and U21204 (N_21204,N_16122,N_17074);
and U21205 (N_21205,N_18290,N_16982);
and U21206 (N_21206,N_16009,N_19183);
nor U21207 (N_21207,N_16942,N_16534);
nand U21208 (N_21208,N_16363,N_16140);
nand U21209 (N_21209,N_17777,N_17731);
and U21210 (N_21210,N_19260,N_15701);
nor U21211 (N_21211,N_16800,N_17980);
and U21212 (N_21212,N_15453,N_17229);
nand U21213 (N_21213,N_19970,N_17154);
and U21214 (N_21214,N_16196,N_15041);
nor U21215 (N_21215,N_15272,N_17309);
nand U21216 (N_21216,N_18031,N_16041);
and U21217 (N_21217,N_15344,N_18631);
or U21218 (N_21218,N_17092,N_19070);
nor U21219 (N_21219,N_15496,N_15457);
or U21220 (N_21220,N_15715,N_16713);
nand U21221 (N_21221,N_16111,N_15664);
and U21222 (N_21222,N_15977,N_18151);
nor U21223 (N_21223,N_16256,N_15046);
nand U21224 (N_21224,N_17584,N_17179);
or U21225 (N_21225,N_16049,N_17220);
or U21226 (N_21226,N_15580,N_16350);
and U21227 (N_21227,N_19309,N_18251);
nor U21228 (N_21228,N_19646,N_19503);
and U21229 (N_21229,N_15298,N_18078);
and U21230 (N_21230,N_19000,N_17038);
xnor U21231 (N_21231,N_15925,N_18914);
nand U21232 (N_21232,N_19527,N_16640);
nand U21233 (N_21233,N_17276,N_19076);
nor U21234 (N_21234,N_16494,N_17661);
nor U21235 (N_21235,N_16726,N_15314);
and U21236 (N_21236,N_19961,N_17852);
and U21237 (N_21237,N_15629,N_17165);
xnor U21238 (N_21238,N_18514,N_16074);
or U21239 (N_21239,N_16287,N_15889);
nand U21240 (N_21240,N_16384,N_15510);
and U21241 (N_21241,N_16392,N_15658);
and U21242 (N_21242,N_15360,N_18725);
nand U21243 (N_21243,N_17190,N_19329);
or U21244 (N_21244,N_16903,N_16823);
nand U21245 (N_21245,N_16021,N_18011);
or U21246 (N_21246,N_17400,N_17374);
and U21247 (N_21247,N_15341,N_16255);
or U21248 (N_21248,N_16855,N_18449);
or U21249 (N_21249,N_18071,N_16407);
or U21250 (N_21250,N_18656,N_16525);
nand U21251 (N_21251,N_19778,N_17114);
nand U21252 (N_21252,N_18447,N_17119);
nand U21253 (N_21253,N_17979,N_19420);
and U21254 (N_21254,N_16970,N_16991);
and U21255 (N_21255,N_19789,N_18249);
nand U21256 (N_21256,N_19799,N_19090);
or U21257 (N_21257,N_16891,N_16061);
nand U21258 (N_21258,N_19666,N_17735);
or U21259 (N_21259,N_18673,N_16331);
nand U21260 (N_21260,N_16011,N_16271);
nor U21261 (N_21261,N_15816,N_18456);
or U21262 (N_21262,N_19149,N_18051);
and U21263 (N_21263,N_19675,N_18765);
nand U21264 (N_21264,N_16132,N_16815);
or U21265 (N_21265,N_16930,N_18621);
or U21266 (N_21266,N_16377,N_17538);
nor U21267 (N_21267,N_16183,N_19749);
nand U21268 (N_21268,N_18026,N_18367);
nor U21269 (N_21269,N_17816,N_18645);
or U21270 (N_21270,N_19184,N_16264);
or U21271 (N_21271,N_15877,N_15688);
and U21272 (N_21272,N_18525,N_18437);
and U21273 (N_21273,N_17398,N_17528);
nand U21274 (N_21274,N_15598,N_15217);
nand U21275 (N_21275,N_15334,N_19269);
nand U21276 (N_21276,N_19499,N_19620);
nand U21277 (N_21277,N_15734,N_15012);
nand U21278 (N_21278,N_19370,N_17629);
nor U21279 (N_21279,N_15104,N_17948);
or U21280 (N_21280,N_15347,N_18436);
or U21281 (N_21281,N_18670,N_19120);
and U21282 (N_21282,N_18636,N_16833);
or U21283 (N_21283,N_15947,N_19840);
nand U21284 (N_21284,N_17795,N_17151);
and U21285 (N_21285,N_17286,N_15079);
nor U21286 (N_21286,N_17893,N_17158);
and U21287 (N_21287,N_17672,N_15837);
or U21288 (N_21288,N_16027,N_19958);
and U21289 (N_21289,N_18285,N_18185);
nand U21290 (N_21290,N_18610,N_15190);
and U21291 (N_21291,N_17228,N_15970);
or U21292 (N_21292,N_17501,N_17610);
nor U21293 (N_21293,N_17558,N_17123);
nor U21294 (N_21294,N_17443,N_16616);
nand U21295 (N_21295,N_16886,N_19980);
nor U21296 (N_21296,N_15328,N_15760);
and U21297 (N_21297,N_19392,N_15583);
and U21298 (N_21298,N_19093,N_16771);
nor U21299 (N_21299,N_19425,N_15408);
or U21300 (N_21300,N_18995,N_16116);
nand U21301 (N_21301,N_17247,N_19485);
and U21302 (N_21302,N_19555,N_17364);
nand U21303 (N_21303,N_17213,N_19634);
or U21304 (N_21304,N_19303,N_15745);
nand U21305 (N_21305,N_18555,N_18390);
nor U21306 (N_21306,N_15860,N_16999);
nand U21307 (N_21307,N_18050,N_16418);
nand U21308 (N_21308,N_16047,N_17187);
nor U21309 (N_21309,N_18162,N_16297);
nor U21310 (N_21310,N_18252,N_17355);
or U21311 (N_21311,N_19477,N_16946);
nand U21312 (N_21312,N_17596,N_19610);
nand U21313 (N_21313,N_15062,N_17011);
nand U21314 (N_21314,N_15973,N_18869);
nor U21315 (N_21315,N_18837,N_17148);
nor U21316 (N_21316,N_16780,N_19986);
and U21317 (N_21317,N_16081,N_15609);
nand U21318 (N_21318,N_17967,N_19718);
and U21319 (N_21319,N_19834,N_18001);
or U21320 (N_21320,N_15403,N_15919);
nor U21321 (N_21321,N_17797,N_19440);
and U21322 (N_21322,N_15709,N_15424);
and U21323 (N_21323,N_15200,N_17913);
and U21324 (N_21324,N_19931,N_18868);
or U21325 (N_21325,N_16214,N_17654);
nor U21326 (N_21326,N_15085,N_19913);
or U21327 (N_21327,N_19471,N_16577);
nand U21328 (N_21328,N_17046,N_17472);
nor U21329 (N_21329,N_18055,N_19857);
nand U21330 (N_21330,N_18883,N_15665);
and U21331 (N_21331,N_19413,N_18174);
nor U21332 (N_21332,N_16450,N_16416);
and U21333 (N_21333,N_16757,N_16203);
and U21334 (N_21334,N_18046,N_19470);
nand U21335 (N_21335,N_15821,N_19708);
nand U21336 (N_21336,N_16071,N_18552);
nor U21337 (N_21337,N_15940,N_15508);
nor U21338 (N_21338,N_19473,N_19376);
or U21339 (N_21339,N_18242,N_17077);
or U21340 (N_21340,N_15831,N_17365);
and U21341 (N_21341,N_17934,N_15460);
or U21342 (N_21342,N_16925,N_16939);
nor U21343 (N_21343,N_19520,N_18843);
and U21344 (N_21344,N_15165,N_16511);
and U21345 (N_21345,N_17157,N_16808);
nor U21346 (N_21346,N_16176,N_19953);
xor U21347 (N_21347,N_19552,N_19325);
and U21348 (N_21348,N_18142,N_18379);
or U21349 (N_21349,N_19877,N_16961);
and U21350 (N_21350,N_17310,N_18107);
nor U21351 (N_21351,N_15464,N_18815);
nand U21352 (N_21352,N_17215,N_15112);
and U21353 (N_21353,N_16517,N_16775);
nor U21354 (N_21354,N_16650,N_17347);
and U21355 (N_21355,N_17844,N_16097);
nor U21356 (N_21356,N_19895,N_17439);
or U21357 (N_21357,N_19711,N_18800);
or U21358 (N_21358,N_15982,N_17344);
or U21359 (N_21359,N_19940,N_17403);
nor U21360 (N_21360,N_18586,N_16308);
or U21361 (N_21361,N_18844,N_16362);
or U21362 (N_21362,N_16693,N_16375);
or U21363 (N_21363,N_16415,N_19545);
or U21364 (N_21364,N_16124,N_17630);
nor U21365 (N_21365,N_15462,N_18655);
nand U21366 (N_21366,N_15441,N_19333);
nor U21367 (N_21367,N_18204,N_16252);
xor U21368 (N_21368,N_16239,N_17663);
or U21369 (N_21369,N_15348,N_16787);
or U21370 (N_21370,N_15554,N_19787);
or U21371 (N_21371,N_19164,N_17884);
or U21372 (N_21372,N_19288,N_18076);
or U21373 (N_21373,N_18460,N_17005);
or U21374 (N_21374,N_17358,N_17381);
or U21375 (N_21375,N_17471,N_18624);
nand U21376 (N_21376,N_18217,N_17800);
nor U21377 (N_21377,N_15340,N_16128);
nand U21378 (N_21378,N_17891,N_15838);
nor U21379 (N_21379,N_16052,N_15516);
nor U21380 (N_21380,N_16864,N_19647);
nor U21381 (N_21381,N_17271,N_19626);
and U21382 (N_21382,N_18763,N_17025);
or U21383 (N_21383,N_19815,N_19261);
nor U21384 (N_21384,N_15931,N_15808);
or U21385 (N_21385,N_16569,N_19129);
nor U21386 (N_21386,N_15780,N_17743);
or U21387 (N_21387,N_17317,N_15670);
or U21388 (N_21388,N_16822,N_19049);
and U21389 (N_21389,N_19064,N_17741);
and U21390 (N_21390,N_15047,N_18501);
nand U21391 (N_21391,N_15096,N_15256);
nor U21392 (N_21392,N_15057,N_16880);
and U21393 (N_21393,N_16729,N_18354);
or U21394 (N_21394,N_15974,N_15727);
or U21395 (N_21395,N_19245,N_19648);
or U21396 (N_21396,N_18810,N_17886);
or U21397 (N_21397,N_19890,N_18891);
or U21398 (N_21398,N_19225,N_18545);
nor U21399 (N_21399,N_19294,N_15286);
or U21400 (N_21400,N_15282,N_18529);
nand U21401 (N_21401,N_19546,N_17178);
or U21402 (N_21402,N_17560,N_16463);
and U21403 (N_21403,N_16233,N_17742);
and U21404 (N_21404,N_18446,N_19014);
and U21405 (N_21405,N_19314,N_15594);
nand U21406 (N_21406,N_16536,N_17124);
and U21407 (N_21407,N_15051,N_17856);
nor U21408 (N_21408,N_16500,N_18267);
and U21409 (N_21409,N_15896,N_16678);
or U21410 (N_21410,N_15678,N_17150);
or U21411 (N_21411,N_16400,N_17577);
nand U21412 (N_21412,N_17516,N_19596);
and U21413 (N_21413,N_15550,N_18980);
and U21414 (N_21414,N_16759,N_15827);
or U21415 (N_21415,N_17897,N_17369);
or U21416 (N_21416,N_15635,N_19824);
nor U21417 (N_21417,N_18842,N_15486);
or U21418 (N_21418,N_17882,N_16048);
or U21419 (N_21419,N_18192,N_18683);
nor U21420 (N_21420,N_17724,N_17572);
nand U21421 (N_21421,N_19078,N_15842);
and U21422 (N_21422,N_19598,N_16109);
or U21423 (N_21423,N_19423,N_15273);
nor U21424 (N_21424,N_19933,N_18568);
or U21425 (N_21425,N_18813,N_16535);
or U21426 (N_21426,N_16090,N_19562);
and U21427 (N_21427,N_16184,N_19092);
nand U21428 (N_21428,N_19705,N_17335);
nand U21429 (N_21429,N_19716,N_16148);
and U21430 (N_21430,N_16854,N_17367);
nand U21431 (N_21431,N_18996,N_17197);
nor U21432 (N_21432,N_15883,N_15563);
and U21433 (N_21433,N_16391,N_19462);
nand U21434 (N_21434,N_18912,N_16526);
and U21435 (N_21435,N_16881,N_18411);
and U21436 (N_21436,N_17386,N_19915);
nand U21437 (N_21437,N_19863,N_18486);
nand U21438 (N_21438,N_17492,N_15019);
or U21439 (N_21439,N_17556,N_16334);
or U21440 (N_21440,N_16125,N_18318);
nand U21441 (N_21441,N_18492,N_19326);
nor U21442 (N_21442,N_18264,N_18954);
nand U21443 (N_21443,N_17859,N_15040);
or U21444 (N_21444,N_17627,N_15111);
and U21445 (N_21445,N_18855,N_19670);
or U21446 (N_21446,N_19165,N_19372);
or U21447 (N_21447,N_18215,N_18949);
nor U21448 (N_21448,N_17467,N_19203);
nor U21449 (N_21449,N_19445,N_19515);
or U21450 (N_21450,N_17481,N_17674);
nor U21451 (N_21451,N_17349,N_17510);
nand U21452 (N_21452,N_15833,N_19768);
or U21453 (N_21453,N_19740,N_16533);
and U21454 (N_21454,N_16358,N_15834);
and U21455 (N_21455,N_16793,N_15872);
and U21456 (N_21456,N_15662,N_18027);
nor U21457 (N_21457,N_17447,N_18591);
nor U21458 (N_21458,N_19297,N_17997);
nand U21459 (N_21459,N_18003,N_17894);
nor U21460 (N_21460,N_18985,N_15802);
or U21461 (N_21461,N_16014,N_17436);
nand U21462 (N_21462,N_17205,N_19809);
nand U21463 (N_21463,N_18035,N_18187);
nand U21464 (N_21464,N_15866,N_16413);
nand U21465 (N_21465,N_15730,N_16635);
and U21466 (N_21466,N_16394,N_19307);
nand U21467 (N_21467,N_15752,N_18092);
and U21468 (N_21468,N_16537,N_18977);
xnor U21469 (N_21469,N_19428,N_17002);
nor U21470 (N_21470,N_17057,N_17174);
nor U21471 (N_21471,N_16155,N_16673);
and U21472 (N_21472,N_16692,N_19410);
and U21473 (N_21473,N_16596,N_19820);
nor U21474 (N_21474,N_16684,N_16298);
or U21475 (N_21475,N_19767,N_16380);
and U21476 (N_21476,N_17782,N_15442);
nor U21477 (N_21477,N_16490,N_17747);
and U21478 (N_21478,N_15531,N_17128);
or U21479 (N_21479,N_15412,N_17222);
nor U21480 (N_21480,N_18785,N_15374);
nand U21481 (N_21481,N_18096,N_18838);
nor U21482 (N_21482,N_16449,N_15418);
nor U21483 (N_21483,N_16658,N_17212);
or U21484 (N_21484,N_19849,N_18907);
and U21485 (N_21485,N_19576,N_16784);
nor U21486 (N_21486,N_17622,N_19371);
and U21487 (N_21487,N_15761,N_19501);
or U21488 (N_21488,N_19362,N_16101);
nor U21489 (N_21489,N_15123,N_19938);
and U21490 (N_21490,N_18422,N_15270);
nor U21491 (N_21491,N_16742,N_15611);
nand U21492 (N_21492,N_15871,N_18585);
nand U21493 (N_21493,N_18619,N_18155);
or U21494 (N_21494,N_17470,N_17531);
and U21495 (N_21495,N_15551,N_17916);
and U21496 (N_21496,N_16157,N_19784);
nor U21497 (N_21497,N_16617,N_18167);
nand U21498 (N_21498,N_16185,N_19739);
and U21499 (N_21499,N_16754,N_16597);
nor U21500 (N_21500,N_19563,N_19384);
nor U21501 (N_21501,N_18686,N_18970);
or U21502 (N_21502,N_19663,N_17801);
nor U21503 (N_21503,N_15160,N_15013);
xnor U21504 (N_21504,N_19517,N_15625);
nand U21505 (N_21505,N_17342,N_16690);
nor U21506 (N_21506,N_16962,N_19956);
or U21507 (N_21507,N_18126,N_16073);
nand U21508 (N_21508,N_19171,N_19495);
and U21509 (N_21509,N_19771,N_18048);
and U21510 (N_21510,N_19929,N_15393);
or U21511 (N_21511,N_16586,N_19219);
and U21512 (N_21512,N_16017,N_18530);
nor U21513 (N_21513,N_17899,N_15392);
and U21514 (N_21514,N_15235,N_19441);
nor U21515 (N_21515,N_19476,N_18761);
or U21516 (N_21516,N_15703,N_16871);
nor U21517 (N_21517,N_17646,N_18626);
and U21518 (N_21518,N_17867,N_16121);
or U21519 (N_21519,N_18528,N_19608);
nand U21520 (N_21520,N_18275,N_17460);
nor U21521 (N_21521,N_15208,N_16210);
nor U21522 (N_21522,N_19084,N_16063);
nor U21523 (N_21523,N_19879,N_15840);
nor U21524 (N_21524,N_18183,N_17193);
and U21525 (N_21525,N_18601,N_15066);
and U21526 (N_21526,N_16395,N_16581);
and U21527 (N_21527,N_15356,N_19833);
nand U21528 (N_21528,N_16731,N_16904);
and U21529 (N_21529,N_16169,N_18566);
nor U21530 (N_21530,N_16530,N_18457);
or U21531 (N_21531,N_16538,N_19228);
nand U21532 (N_21532,N_16389,N_15354);
nand U21533 (N_21533,N_15197,N_19661);
and U21534 (N_21534,N_17539,N_16215);
or U21535 (N_21535,N_15296,N_16803);
and U21536 (N_21536,N_15362,N_19113);
and U21537 (N_21537,N_16568,N_15786);
or U21538 (N_21538,N_16315,N_16293);
and U21539 (N_21539,N_17656,N_18880);
and U21540 (N_21540,N_18255,N_15018);
or U21541 (N_21541,N_16099,N_19434);
or U21542 (N_21542,N_17244,N_18993);
or U21543 (N_21543,N_19296,N_18934);
or U21544 (N_21544,N_15281,N_15818);
or U21545 (N_21545,N_17957,N_16115);
or U21546 (N_21546,N_19746,N_15135);
and U21547 (N_21547,N_18465,N_17024);
nand U21548 (N_21548,N_15232,N_18671);
nor U21549 (N_21549,N_15023,N_17641);
nand U21550 (N_21550,N_16983,N_17245);
nor U21551 (N_21551,N_17828,N_19649);
and U21552 (N_21552,N_15647,N_19726);
nor U21553 (N_21553,N_18783,N_19937);
or U21554 (N_21554,N_19622,N_17281);
and U21555 (N_21555,N_18115,N_18127);
nand U21556 (N_21556,N_18282,N_15479);
nand U21557 (N_21557,N_17737,N_19855);
or U21558 (N_21558,N_15201,N_19025);
nand U21559 (N_21559,N_16411,N_19147);
nor U21560 (N_21560,N_15950,N_18828);
nor U21561 (N_21561,N_18459,N_16053);
nor U21562 (N_21562,N_17695,N_17843);
nor U21563 (N_21563,N_17667,N_16758);
xnor U21564 (N_21564,N_15413,N_18938);
nand U21565 (N_21565,N_17216,N_15365);
and U21566 (N_21566,N_18704,N_16628);
or U21567 (N_21567,N_19405,N_15133);
nand U21568 (N_21568,N_18588,N_19521);
nand U21569 (N_21569,N_17044,N_18419);
or U21570 (N_21570,N_19777,N_16540);
nor U21571 (N_21571,N_19602,N_16200);
nor U21572 (N_21572,N_15984,N_16825);
nand U21573 (N_21573,N_19365,N_16745);
nor U21574 (N_21574,N_17132,N_17612);
nor U21575 (N_21575,N_18355,N_19401);
nand U21576 (N_21576,N_19346,N_19464);
or U21577 (N_21577,N_15284,N_19334);
nor U21578 (N_21578,N_18926,N_19978);
nand U21579 (N_21579,N_17693,N_19060);
and U21580 (N_21580,N_15155,N_19588);
nor U21581 (N_21581,N_17079,N_19157);
and U21582 (N_21582,N_15101,N_15501);
nor U21583 (N_21583,N_18973,N_18490);
nor U21584 (N_21584,N_17017,N_16209);
and U21585 (N_21585,N_15136,N_17070);
nand U21586 (N_21586,N_19821,N_19321);
nand U21587 (N_21587,N_15125,N_16166);
nor U21588 (N_21588,N_18861,N_19531);
nand U21589 (N_21589,N_19910,N_18228);
or U21590 (N_21590,N_15290,N_19707);
and U21591 (N_21591,N_16732,N_15140);
and U21592 (N_21592,N_18853,N_15867);
or U21593 (N_21593,N_18801,N_17029);
and U21594 (N_21594,N_19650,N_17380);
nor U21595 (N_21595,N_15423,N_19573);
and U21596 (N_21596,N_15672,N_15005);
nand U21597 (N_21597,N_17278,N_19658);
nand U21598 (N_21598,N_17619,N_19002);
or U21599 (N_21599,N_18602,N_17827);
and U21600 (N_21600,N_17639,N_16549);
or U21601 (N_21601,N_17176,N_17666);
nor U21602 (N_21602,N_15297,N_17113);
nor U21603 (N_21603,N_16720,N_15253);
or U21604 (N_21604,N_18059,N_18695);
nand U21605 (N_21605,N_16112,N_18902);
nand U21606 (N_21606,N_18169,N_19660);
nand U21607 (N_21607,N_19267,N_17152);
and U21608 (N_21608,N_15857,N_19564);
nand U21609 (N_21609,N_16057,N_18034);
and U21610 (N_21610,N_18908,N_18878);
and U21611 (N_21611,N_16432,N_15967);
and U21612 (N_21612,N_19424,N_15446);
nor U21613 (N_21613,N_17890,N_16835);
nor U21614 (N_21614,N_16476,N_19629);
xor U21615 (N_21615,N_16202,N_16272);
nor U21616 (N_21616,N_16426,N_15578);
nor U21617 (N_21617,N_17188,N_17284);
nand U21618 (N_21618,N_16764,N_17975);
nand U21619 (N_21619,N_15694,N_16180);
and U21620 (N_21620,N_19461,N_16488);
or U21621 (N_21621,N_19681,N_16988);
nand U21622 (N_21622,N_17219,N_17066);
nand U21623 (N_21623,N_19435,N_16032);
nor U21624 (N_21624,N_18784,N_19363);
or U21625 (N_21625,N_15113,N_18499);
nand U21626 (N_21626,N_16257,N_18978);
and U21627 (N_21627,N_19955,N_16198);
or U21628 (N_21628,N_16978,N_17456);
and U21629 (N_21629,N_16066,N_18254);
nor U21630 (N_21630,N_19706,N_17605);
and U21631 (N_21631,N_18714,N_17732);
nand U21632 (N_21632,N_19021,N_15612);
and U21633 (N_21633,N_18659,N_15864);
and U21634 (N_21634,N_18548,N_16004);
or U21635 (N_21635,N_17520,N_15992);
nor U21636 (N_21636,N_18359,N_17575);
nor U21637 (N_21637,N_18807,N_18863);
or U21638 (N_21638,N_17226,N_16077);
or U21639 (N_21639,N_15431,N_15875);
nand U21640 (N_21640,N_18814,N_16437);
nand U21641 (N_21641,N_16820,N_15241);
or U21642 (N_21642,N_15862,N_17028);
nand U21643 (N_21643,N_15132,N_15545);
nor U21644 (N_21644,N_18538,N_16696);
nor U21645 (N_21645,N_18362,N_18554);
or U21646 (N_21646,N_19204,N_17545);
nor U21647 (N_21647,N_15557,N_16737);
or U21648 (N_21648,N_19699,N_17532);
nor U21649 (N_21649,N_19935,N_15333);
nor U21650 (N_21650,N_15093,N_18587);
or U21651 (N_21651,N_19559,N_17312);
nand U21652 (N_21652,N_16694,N_16089);
and U21653 (N_21653,N_16809,N_17822);
nand U21654 (N_21654,N_16095,N_19782);
or U21655 (N_21655,N_18296,N_17614);
and U21656 (N_21656,N_19964,N_15182);
xnor U21657 (N_21657,N_19268,N_17776);
nand U21658 (N_21658,N_18794,N_17255);
and U21659 (N_21659,N_15484,N_18244);
or U21660 (N_21660,N_19298,N_18721);
and U21661 (N_21661,N_16211,N_16913);
or U21662 (N_21662,N_17504,N_19208);
nor U21663 (N_21663,N_18154,N_15092);
nor U21664 (N_21664,N_19230,N_15910);
nand U21665 (N_21665,N_16179,N_15366);
and U21666 (N_21666,N_16149,N_17648);
nand U21667 (N_21667,N_18642,N_15251);
xor U21668 (N_21668,N_18543,N_15083);
and U21669 (N_21669,N_15659,N_17334);
or U21670 (N_21670,N_15152,N_16817);
nor U21671 (N_21671,N_17557,N_19510);
and U21672 (N_21672,N_15398,N_15948);
nor U21673 (N_21673,N_18343,N_15076);
nor U21674 (N_21674,N_15465,N_18475);
nor U21675 (N_21675,N_16722,N_19859);
nor U21676 (N_21676,N_18638,N_19457);
or U21677 (N_21677,N_16748,N_18111);
and U21678 (N_21678,N_17751,N_15614);
nand U21679 (N_21679,N_16251,N_16977);
nand U21680 (N_21680,N_16919,N_15080);
and U21681 (N_21681,N_16676,N_16303);
nand U21682 (N_21682,N_19282,N_15908);
or U21683 (N_21683,N_19551,N_18073);
and U21684 (N_21684,N_18901,N_19680);
xor U21685 (N_21685,N_16659,N_15168);
or U21686 (N_21686,N_16338,N_19870);
nor U21687 (N_21687,N_16741,N_15542);
nand U21688 (N_21688,N_17341,N_19033);
or U21689 (N_21689,N_18757,N_17506);
nor U21690 (N_21690,N_15078,N_15747);
or U21691 (N_21691,N_19535,N_18405);
nor U21692 (N_21692,N_15628,N_15299);
and U21693 (N_21693,N_17945,N_17184);
and U21694 (N_21694,N_17805,N_16359);
and U21695 (N_21695,N_19024,N_17670);
nor U21696 (N_21696,N_15072,N_19874);
nor U21697 (N_21697,N_18143,N_15313);
or U21698 (N_21698,N_15031,N_16217);
nand U21699 (N_21699,N_19810,N_17991);
nand U21700 (N_21700,N_16283,N_18876);
or U21701 (N_21701,N_15312,N_16092);
nand U21702 (N_21702,N_15537,N_16248);
nand U21703 (N_21703,N_19530,N_16655);
or U21704 (N_21704,N_19807,N_18923);
and U21705 (N_21705,N_15654,N_17256);
nand U21706 (N_21706,N_17042,N_19374);
and U21707 (N_21707,N_19698,N_18165);
xor U21708 (N_21708,N_15088,N_18288);
and U21709 (N_21709,N_18515,N_16824);
and U21710 (N_21710,N_16993,N_19548);
or U21711 (N_21711,N_19884,N_18120);
or U21712 (N_21712,N_18243,N_18798);
or U21713 (N_21713,N_18781,N_17243);
or U21714 (N_21714,N_15448,N_15174);
nand U21715 (N_21715,N_17343,N_18389);
and U21716 (N_21716,N_18939,N_18461);
or U21717 (N_21717,N_16441,N_19889);
nand U21718 (N_21718,N_17848,N_16019);
or U21719 (N_21719,N_16312,N_19954);
and U21720 (N_21720,N_15784,N_18759);
or U21721 (N_21721,N_17357,N_18316);
or U21722 (N_21722,N_19347,N_16065);
or U21723 (N_21723,N_18772,N_19308);
and U21724 (N_21724,N_18668,N_18598);
and U21725 (N_21725,N_17076,N_18080);
and U21726 (N_21726,N_16379,N_18233);
nor U21727 (N_21727,N_16345,N_17107);
nand U21728 (N_21728,N_15836,N_19352);
nor U21729 (N_21729,N_17112,N_18117);
nor U21730 (N_21730,N_19512,N_15785);
nor U21731 (N_21731,N_15546,N_18786);
nand U21732 (N_21732,N_15683,N_16498);
nand U21733 (N_21733,N_18482,N_16712);
nor U21734 (N_21734,N_17329,N_18209);
and U21735 (N_21735,N_17818,N_17186);
or U21736 (N_21736,N_15975,N_16572);
or U21737 (N_21737,N_15186,N_17127);
nor U21738 (N_21738,N_16245,N_15143);
xor U21739 (N_21739,N_17847,N_17336);
and U21740 (N_21740,N_15511,N_15230);
and U21741 (N_21741,N_15593,N_16107);
nand U21742 (N_21742,N_15026,N_15454);
nand U21743 (N_21743,N_18315,N_18707);
and U21744 (N_21744,N_15119,N_17491);
nor U21745 (N_21745,N_19004,N_15638);
nor U21746 (N_21746,N_15964,N_16944);
or U21747 (N_21747,N_16138,N_18957);
nand U21748 (N_21748,N_16622,N_17766);
or U21749 (N_21749,N_19018,N_16056);
and U21750 (N_21750,N_16222,N_17725);
nand U21751 (N_21751,N_19715,N_18058);
and U21752 (N_21752,N_19187,N_17431);
or U21753 (N_21753,N_17133,N_16486);
and U21754 (N_21754,N_16902,N_16410);
nand U21755 (N_21755,N_16920,N_18451);
nand U21756 (N_21756,N_18986,N_17339);
nor U21757 (N_21757,N_18652,N_16804);
nor U21758 (N_21758,N_19860,N_15527);
nor U21759 (N_21759,N_17306,N_19798);
or U21760 (N_21760,N_17570,N_16873);
and U21761 (N_21761,N_19170,N_19096);
and U21762 (N_21762,N_17729,N_18581);
nor U21763 (N_21763,N_16373,N_18532);
and U21764 (N_21764,N_16620,N_18415);
or U21765 (N_21765,N_17905,N_19594);
and U21766 (N_21766,N_16030,N_15845);
nor U21767 (N_21767,N_17440,N_17540);
or U21768 (N_21768,N_19169,N_17141);
and U21769 (N_21769,N_15630,N_17565);
nor U21770 (N_21770,N_18812,N_16558);
nand U21771 (N_21771,N_17499,N_18584);
and U21772 (N_21772,N_16642,N_17360);
or U21773 (N_21773,N_16975,N_16705);
or U21774 (N_21774,N_18363,N_15622);
xor U21775 (N_21775,N_18434,N_16782);
nor U21776 (N_21776,N_18500,N_15913);
or U21777 (N_21777,N_18414,N_19731);
or U21778 (N_21778,N_19123,N_16646);
nand U21779 (N_21779,N_16265,N_18556);
or U21780 (N_21780,N_17810,N_17130);
nor U21781 (N_21781,N_19174,N_15648);
nor U21782 (N_21782,N_17982,N_19348);
or U21783 (N_21783,N_16420,N_18563);
nand U21784 (N_21784,N_17363,N_17290);
nor U21785 (N_21785,N_19104,N_15943);
nand U21786 (N_21786,N_17734,N_19645);
nor U21787 (N_21787,N_16518,N_17845);
or U21788 (N_21788,N_17305,N_18086);
or U21789 (N_21789,N_15175,N_16550);
nor U21790 (N_21790,N_19566,N_17240);
and U21791 (N_21791,N_18729,N_19396);
nor U21792 (N_21792,N_15766,N_16477);
xnor U21793 (N_21793,N_19009,N_17161);
or U21794 (N_21794,N_15316,N_19008);
nand U21795 (N_21795,N_16662,N_15110);
nand U21796 (N_21796,N_15641,N_19148);
and U21797 (N_21797,N_15954,N_19941);
nand U21798 (N_21798,N_15579,N_16932);
nand U21799 (N_21799,N_18416,N_19209);
or U21800 (N_21800,N_18481,N_17288);
and U21801 (N_21801,N_15795,N_16677);
nor U21802 (N_21802,N_15137,N_18820);
or U21803 (N_21803,N_16102,N_19121);
xor U21804 (N_21804,N_19318,N_17698);
or U21805 (N_21805,N_19838,N_19632);
nor U21806 (N_21806,N_16326,N_17438);
and U21807 (N_21807,N_18311,N_19755);
nor U21808 (N_21808,N_15868,N_19277);
and U21809 (N_21809,N_15680,N_16666);
nor U21810 (N_21810,N_18700,N_15689);
nand U21811 (N_21811,N_19742,N_15202);
or U21812 (N_21812,N_18203,N_16309);
nor U21813 (N_21813,N_16763,N_17108);
nor U21814 (N_21814,N_17359,N_16844);
nand U21815 (N_21815,N_15483,N_15846);
nor U21816 (N_21816,N_19007,N_17662);
nand U21817 (N_21817,N_15666,N_15367);
or U21818 (N_21818,N_18788,N_16938);
and U21819 (N_21819,N_16156,N_15050);
nand U21820 (N_21820,N_18666,N_16554);
and U21821 (N_21821,N_19216,N_19965);
nor U21822 (N_21822,N_15475,N_16022);
nand U21823 (N_21823,N_15049,N_16512);
nand U21824 (N_21824,N_18579,N_18753);
and U21825 (N_21825,N_18944,N_16893);
and U21826 (N_21826,N_17140,N_15240);
nand U21827 (N_21827,N_17476,N_16299);
nand U21828 (N_21828,N_17824,N_15951);
and U21829 (N_21829,N_18928,N_16936);
and U21830 (N_21830,N_15887,N_16333);
nand U21831 (N_21831,N_15069,N_19919);
or U21832 (N_21832,N_17164,N_19537);
or U21833 (N_21833,N_15832,N_16347);
and U21834 (N_21834,N_18718,N_16171);
nand U21835 (N_21835,N_15163,N_15411);
and U21836 (N_21836,N_15248,N_16849);
nand U21837 (N_21837,N_15639,N_18851);
and U21838 (N_21838,N_16606,N_18871);
nor U21839 (N_21839,N_17040,N_19756);
nor U21840 (N_21840,N_17582,N_17911);
nor U21841 (N_21841,N_19240,N_17677);
and U21842 (N_21842,N_18310,N_18060);
and U21843 (N_21843,N_19226,N_18767);
nor U21844 (N_21844,N_17315,N_16008);
or U21845 (N_21845,N_16458,N_15710);
nand U21846 (N_21846,N_16645,N_17009);
nand U21847 (N_21847,N_18295,N_18172);
nor U21848 (N_21848,N_19212,N_19952);
nor U21849 (N_21849,N_18709,N_19994);
or U21850 (N_21850,N_17033,N_15755);
nor U21851 (N_21851,N_16291,N_19944);
or U21852 (N_21852,N_17679,N_16595);
nor U21853 (N_21853,N_18872,N_18410);
or U21854 (N_21854,N_15804,N_19797);
and U21855 (N_21855,N_16665,N_16055);
or U21856 (N_21856,N_17611,N_15893);
nand U21857 (N_21857,N_17853,N_18713);
nand U21858 (N_21858,N_15682,N_19526);
or U21859 (N_21859,N_18435,N_16105);
or U21860 (N_21860,N_17744,N_18896);
nand U21861 (N_21861,N_15812,N_19906);
nor U21862 (N_21862,N_17338,N_16585);
nand U21863 (N_21863,N_16948,N_18750);
and U21864 (N_21864,N_16561,N_15588);
nand U21865 (N_21865,N_15139,N_16669);
nand U21866 (N_21866,N_15054,N_17437);
nor U21867 (N_21867,N_15184,N_17319);
nor U21868 (N_21868,N_19029,N_18105);
or U21869 (N_21869,N_18314,N_17998);
and U21870 (N_21870,N_17051,N_16455);
nand U21871 (N_21871,N_15105,N_15310);
or U21872 (N_21872,N_15565,N_17713);
nor U21873 (N_21873,N_18895,N_18337);
nor U21874 (N_21874,N_16168,N_19848);
xor U21875 (N_21875,N_16573,N_15268);
nand U21876 (N_21876,N_19883,N_16862);
nand U21877 (N_21877,N_19335,N_19962);
nor U21878 (N_21878,N_15144,N_15960);
or U21879 (N_21879,N_18680,N_15905);
nor U21880 (N_21880,N_18732,N_18225);
and U21881 (N_21881,N_16797,N_16866);
or U21882 (N_21882,N_19407,N_19690);
nor U21883 (N_21883,N_15996,N_18823);
or U21884 (N_21884,N_16422,N_17327);
nor U21885 (N_21885,N_16253,N_16994);
nand U21886 (N_21886,N_15400,N_17860);
nor U21887 (N_21887,N_18537,N_15091);
nor U21888 (N_21888,N_16159,N_17292);
nor U21889 (N_21889,N_16381,N_15615);
nand U21890 (N_21890,N_18974,N_17764);
or U21891 (N_21891,N_15937,N_19131);
or U21892 (N_21892,N_16344,N_15790);
nor U21893 (N_21893,N_15874,N_19867);
or U21894 (N_21894,N_18094,N_18074);
nor U21895 (N_21895,N_19976,N_19544);
or U21896 (N_21896,N_19547,N_18881);
or U21897 (N_21897,N_19075,N_19266);
nand U21898 (N_21898,N_16654,N_16580);
or U21899 (N_21899,N_15294,N_16181);
nand U21900 (N_21900,N_19137,N_15428);
nand U21901 (N_21901,N_16818,N_19489);
or U21902 (N_21902,N_15607,N_15958);
nand U21903 (N_21903,N_17819,N_16076);
nor U21904 (N_21904,N_18726,N_19989);
nor U21905 (N_21905,N_17034,N_17397);
nand U21906 (N_21906,N_15591,N_15869);
and U21907 (N_21907,N_16482,N_16274);
and U21908 (N_21908,N_19793,N_15445);
and U21909 (N_21909,N_15994,N_19052);
or U21910 (N_21910,N_18521,N_15989);
and U21911 (N_21911,N_19514,N_17904);
nor U21912 (N_21912,N_17728,N_17320);
or U21913 (N_21913,N_16277,N_18979);
nor U21914 (N_21914,N_15936,N_15789);
and U21915 (N_21915,N_17238,N_18333);
and U21916 (N_21916,N_16935,N_19920);
or U21917 (N_21917,N_16146,N_17960);
or U21918 (N_21918,N_16321,N_17131);
and U21919 (N_21919,N_16319,N_19803);
and U21920 (N_21920,N_15687,N_15415);
nor U21921 (N_21921,N_16701,N_18464);
nand U21922 (N_21922,N_16288,N_19539);
or U21923 (N_21923,N_16221,N_16015);
or U21924 (N_21924,N_19094,N_16688);
nand U21925 (N_21925,N_18284,N_15319);
nor U21926 (N_21926,N_19871,N_18063);
nand U21927 (N_21927,N_15980,N_16541);
nand U21928 (N_21928,N_19492,N_19764);
nand U21929 (N_21929,N_15157,N_17779);
or U21930 (N_21930,N_19355,N_16894);
and U21931 (N_21931,N_15342,N_17647);
and U21932 (N_21932,N_18156,N_17425);
and U21933 (N_21933,N_17430,N_17091);
and U21934 (N_21934,N_15515,N_19330);
and U21935 (N_21935,N_18989,N_18922);
or U21936 (N_21936,N_15835,N_17454);
and U21937 (N_21937,N_18994,N_16679);
or U21938 (N_21938,N_19340,N_17953);
or U21939 (N_21939,N_15167,N_19250);
or U21940 (N_21940,N_16756,N_19942);
or U21941 (N_21941,N_15234,N_19012);
nand U21942 (N_21942,N_16699,N_19836);
nor U21943 (N_21943,N_19097,N_19127);
nor U21944 (N_21944,N_18826,N_17783);
nand U21945 (N_21945,N_15363,N_16557);
nor U21946 (N_21946,N_15571,N_17815);
and U21947 (N_21947,N_17652,N_19283);
and U21948 (N_21948,N_18066,N_19974);
nor U21949 (N_21949,N_16868,N_17592);
or U21950 (N_21950,N_15610,N_16091);
and U21951 (N_21951,N_18596,N_19437);
or U21952 (N_21952,N_18956,N_16523);
nand U21953 (N_21953,N_15704,N_18334);
nand U21954 (N_21954,N_19677,N_19725);
nand U21955 (N_21955,N_15177,N_17966);
and U21956 (N_21956,N_19571,N_18735);
nand U21957 (N_21957,N_15357,N_16556);
nand U21958 (N_21958,N_19054,N_17175);
xnor U21959 (N_21959,N_19873,N_16600);
and U21960 (N_21960,N_17048,N_16404);
or U21961 (N_21961,N_17554,N_15794);
or U21962 (N_21962,N_15466,N_15324);
nand U21963 (N_21963,N_18266,N_16857);
or U21964 (N_21964,N_19178,N_17722);
or U21965 (N_21965,N_17249,N_18946);
xnor U21966 (N_21966,N_16689,N_18038);
or U21967 (N_21967,N_17578,N_18611);
or U21968 (N_21968,N_19783,N_18056);
and U21969 (N_21969,N_15456,N_19630);
nor U21970 (N_21970,N_16118,N_19117);
nand U21971 (N_21971,N_18551,N_15071);
nand U21972 (N_21972,N_15351,N_19291);
and U21973 (N_21973,N_18887,N_17195);
and U21974 (N_21974,N_18178,N_16207);
nand U21975 (N_21975,N_15934,N_18936);
or U21976 (N_21976,N_16489,N_18361);
and U21977 (N_21977,N_19880,N_17918);
and U21978 (N_21978,N_17705,N_17765);
or U21979 (N_21979,N_15102,N_17791);
nor U21980 (N_21980,N_16100,N_16735);
and U21981 (N_21981,N_17938,N_18262);
nand U21982 (N_21982,N_18240,N_19621);
nor U21983 (N_21983,N_17925,N_16779);
nor U21984 (N_21984,N_17887,N_15037);
nand U21985 (N_21985,N_15841,N_19351);
and U21986 (N_21986,N_19452,N_18442);
and U21987 (N_21987,N_16539,N_18351);
or U21988 (N_21988,N_17514,N_16079);
and U21989 (N_21989,N_16143,N_19641);
nand U21990 (N_21990,N_15539,N_16497);
nand U21991 (N_21991,N_15502,N_19665);
nand U21992 (N_21992,N_15810,N_17294);
nor U21993 (N_21993,N_15645,N_16320);
nand U21994 (N_21994,N_17525,N_15068);
or U21995 (N_21995,N_19558,N_18852);
or U21996 (N_21996,N_18323,N_16368);
and U21997 (N_21997,N_19795,N_17370);
nand U21998 (N_21998,N_18987,N_17994);
and U21999 (N_21999,N_18198,N_18593);
or U22000 (N_22000,N_16965,N_17653);
nor U22001 (N_22001,N_18398,N_18399);
or U22002 (N_22002,N_17298,N_19652);
or U22003 (N_22003,N_16018,N_17808);
nor U22004 (N_22004,N_15029,N_19904);
or U22005 (N_22005,N_17790,N_17598);
nor U22006 (N_22006,N_15343,N_19072);
and U22007 (N_22007,N_16154,N_18775);
and U22008 (N_22008,N_17595,N_18220);
nor U22009 (N_22009,N_15959,N_18087);
and U22010 (N_22010,N_16028,N_15060);
nand U22011 (N_22011,N_17279,N_18308);
or U22012 (N_22012,N_16330,N_18067);
nand U22013 (N_22013,N_15932,N_18328);
nor U22014 (N_22014,N_17869,N_15100);
and U22015 (N_22015,N_17917,N_17340);
nand U22016 (N_22016,N_17638,N_15199);
nor U22017 (N_22017,N_15763,N_15653);
or U22018 (N_22018,N_17712,N_17191);
nor U22019 (N_22019,N_18945,N_15390);
and U22020 (N_22020,N_17616,N_15892);
nor U22021 (N_22021,N_18760,N_16575);
nand U22022 (N_22022,N_17926,N_18504);
nor U22023 (N_22023,N_15277,N_17239);
or U22024 (N_22024,N_15216,N_15293);
and U22025 (N_22025,N_18462,N_15419);
nor U22026 (N_22026,N_19047,N_15829);
or U22027 (N_22027,N_18276,N_19026);
and U22028 (N_22028,N_15489,N_17850);
nand U22029 (N_22029,N_17515,N_17901);
or U22030 (N_22030,N_19589,N_19150);
and U22031 (N_22031,N_16151,N_15302);
nor U22032 (N_22032,N_18320,N_15783);
and U22033 (N_22033,N_17689,N_17954);
nand U22034 (N_22034,N_19750,N_19781);
or U22035 (N_22035,N_19901,N_16262);
nand U22036 (N_22036,N_15045,N_18678);
nor U22037 (N_22037,N_18873,N_17944);
or U22038 (N_22038,N_18856,N_15748);
nand U22039 (N_22039,N_18136,N_17969);
and U22040 (N_22040,N_16423,N_18207);
and U22041 (N_22041,N_17585,N_16280);
and U22042 (N_22042,N_15438,N_15038);
or U22043 (N_22043,N_19368,N_18200);
nand U22044 (N_22044,N_19156,N_19375);
or U22045 (N_22045,N_16023,N_15009);
or U22046 (N_22046,N_16393,N_19426);
or U22047 (N_22047,N_17861,N_15086);
or U22048 (N_22048,N_18960,N_16562);
and U22049 (N_22049,N_17289,N_17787);
nand U22050 (N_22050,N_17907,N_18950);
and U22051 (N_22051,N_18608,N_17680);
or U22052 (N_22052,N_15986,N_16254);
nand U22053 (N_22053,N_16040,N_16643);
nand U22054 (N_22054,N_16914,N_17257);
nor U22055 (N_22055,N_19474,N_15358);
nor U22056 (N_22056,N_17571,N_17774);
or U22057 (N_22057,N_19038,N_18657);
and U22058 (N_22058,N_18575,N_19390);
or U22059 (N_22059,N_17353,N_15805);
nand U22060 (N_22060,N_16467,N_16188);
nor U22061 (N_22061,N_15800,N_17031);
or U22062 (N_22062,N_15923,N_16086);
or U22063 (N_22063,N_19110,N_16734);
nor U22064 (N_22064,N_18916,N_18010);
or U22065 (N_22065,N_19483,N_19142);
and U22066 (N_22066,N_18698,N_19822);
nor U22067 (N_22067,N_17004,N_17003);
or U22068 (N_22068,N_18738,N_16114);
nor U22069 (N_22069,N_16531,N_19019);
and U22070 (N_22070,N_18084,N_19872);
and U22071 (N_22071,N_16851,N_18909);
nor U22072 (N_22072,N_17206,N_15505);
nand U22073 (N_22073,N_19600,N_16910);
nor U22074 (N_22074,N_19893,N_15180);
nand U22075 (N_22075,N_19418,N_16821);
nor U22076 (N_22076,N_16208,N_18637);
and U22077 (N_22077,N_15228,N_17413);
nor U22078 (N_22078,N_19475,N_15305);
nand U22079 (N_22079,N_16901,N_19350);
and U22080 (N_22080,N_15765,N_15815);
and U22081 (N_22081,N_19252,N_18294);
and U22082 (N_22082,N_16323,N_18929);
nor U22083 (N_22083,N_15480,N_17189);
or U22084 (N_22084,N_19519,N_18045);
nand U22085 (N_22085,N_15191,N_18669);
nand U22086 (N_22086,N_16750,N_15117);
nor U22087 (N_22087,N_17740,N_18628);
and U22088 (N_22088,N_16691,N_15853);
nand U22089 (N_22089,N_17541,N_18476);
nor U22090 (N_22090,N_16365,N_15015);
nand U22091 (N_22091,N_18599,N_18291);
and U22092 (N_22092,N_19220,N_16609);
nand U22093 (N_22093,N_18867,N_15352);
nand U22094 (N_22094,N_19082,N_19339);
and U22095 (N_22095,N_17718,N_19043);
nor U22096 (N_22096,N_16492,N_15126);
or U22097 (N_22097,N_17871,N_19198);
or U22098 (N_22098,N_18722,N_18431);
nand U22099 (N_22099,N_19887,N_19898);
or U22100 (N_22100,N_15007,N_18764);
or U22101 (N_22101,N_16524,N_19450);
and U22102 (N_22102,N_15957,N_16652);
nand U22103 (N_22103,N_17951,N_17547);
or U22104 (N_22104,N_15878,N_18052);
nand U22105 (N_22105,N_16301,N_17621);
nor U22106 (N_22106,N_15498,N_19987);
and U22107 (N_22107,N_18778,N_19945);
and U22108 (N_22108,N_17054,N_15646);
and U22109 (N_22109,N_19903,N_17104);
nand U22110 (N_22110,N_18606,N_15799);
and U22111 (N_22111,N_15969,N_16318);
nor U22112 (N_22112,N_18730,N_18195);
or U22113 (N_22113,N_15187,N_16317);
or U22114 (N_22114,N_16890,N_18847);
nand U22115 (N_22115,N_18245,N_19722);
nand U22116 (N_22116,N_15494,N_17895);
or U22117 (N_22117,N_19717,N_15856);
nand U22118 (N_22118,N_18152,N_15221);
nand U22119 (N_22119,N_19609,N_15257);
and U22120 (N_22120,N_18425,N_16672);
or U22121 (N_22121,N_19467,N_16810);
nor U22122 (N_22122,N_18479,N_16704);
and U22123 (N_22123,N_18222,N_19572);
nor U22124 (N_22124,N_17373,N_16908);
and U22125 (N_22125,N_16716,N_17457);
and U22126 (N_22126,N_16990,N_18509);
or U22127 (N_22127,N_17462,N_16372);
nor U22128 (N_22128,N_19868,N_15513);
nor U22129 (N_22129,N_15844,N_18062);
or U22130 (N_22130,N_19195,N_18913);
nand U22131 (N_22131,N_15477,N_17864);
nor U22132 (N_22132,N_18747,N_17803);
or U22133 (N_22133,N_15376,N_15373);
and U22134 (N_22134,N_19295,N_17323);
nand U22135 (N_22135,N_18248,N_17855);
and U22136 (N_22136,N_16408,N_18918);
nand U22137 (N_22137,N_16070,N_18409);
and U22138 (N_22138,N_15218,N_15227);
and U22139 (N_22139,N_19540,N_17697);
nor U22140 (N_22140,N_19507,N_19086);
nor U22141 (N_22141,N_16429,N_18257);
xnor U22142 (N_22142,N_18894,N_19081);
nor U22143 (N_22143,N_17096,N_18646);
nand U22144 (N_22144,N_17153,N_16870);
and U22145 (N_22145,N_15781,N_19854);
nor U22146 (N_22146,N_16725,N_18309);
nor U22147 (N_22147,N_17146,N_17549);
nand U22148 (N_22148,N_15650,N_19251);
nor U22149 (N_22149,N_15617,N_19845);
or U22150 (N_22150,N_18685,N_19173);
nand U22151 (N_22151,N_17122,N_19529);
or U22152 (N_22152,N_19792,N_15260);
nor U22153 (N_22153,N_16963,N_17576);
and U22154 (N_22154,N_19567,N_15420);
nor U22155 (N_22155,N_15410,N_18201);
and U22156 (N_22156,N_19969,N_16956);
nor U22157 (N_22157,N_18731,N_16296);
and U22158 (N_22158,N_19780,N_16986);
nand U22159 (N_22159,N_18572,N_19419);
or U22160 (N_22160,N_18407,N_19579);
nor U22161 (N_22161,N_16134,N_18277);
or U22162 (N_22162,N_16786,N_19280);
and U22163 (N_22163,N_17412,N_15017);
nor U22164 (N_22164,N_16231,N_17978);
nand U22165 (N_22165,N_16711,N_15377);
and U22166 (N_22166,N_17100,N_16147);
and U22167 (N_22167,N_19101,N_15225);
nor U22168 (N_22168,N_19972,N_16456);
nor U22169 (N_22169,N_15207,N_15998);
nand U22170 (N_22170,N_17231,N_18427);
or U22171 (N_22171,N_19273,N_16753);
or U22172 (N_22172,N_17084,N_16602);
nor U22173 (N_22173,N_15813,N_17263);
nor U22174 (N_22174,N_18831,N_17875);
nor U22175 (N_22175,N_19624,N_15561);
or U22176 (N_22176,N_18565,N_19853);
nor U22177 (N_22177,N_15898,N_17587);
nor U22178 (N_22178,N_16933,N_18576);
nand U22179 (N_22179,N_17659,N_17332);
nor U22180 (N_22180,N_19119,N_15109);
and U22181 (N_22181,N_15146,N_18373);
and U22182 (N_22182,N_19744,N_18806);
or U22183 (N_22183,N_15987,N_19932);
nand U22184 (N_22184,N_19246,N_15733);
nand U22185 (N_22185,N_18239,N_15915);
nand U22186 (N_22186,N_15677,N_17477);
or U22187 (N_22187,N_18991,N_19925);
xnor U22188 (N_22188,N_18893,N_15599);
and U22189 (N_22189,N_16972,N_18643);
or U22190 (N_22190,N_15231,N_19466);
or U22191 (N_22191,N_17275,N_16648);
nor U22192 (N_22192,N_16921,N_19041);
nor U22193 (N_22193,N_18018,N_17745);
nor U22194 (N_22194,N_19391,N_19438);
nor U22195 (N_22195,N_18803,N_19153);
nand U22196 (N_22196,N_17906,N_16778);
nor U22197 (N_22197,N_17601,N_18029);
nand U22198 (N_22198,N_18345,N_15036);
or U22199 (N_22199,N_15806,N_17559);
nor U22200 (N_22200,N_16000,N_17352);
nor U22201 (N_22201,N_16633,N_15318);
or U22202 (N_22202,N_16225,N_16446);
or U22203 (N_22203,N_17542,N_15330);
or U22204 (N_22204,N_17650,N_17811);
or U22205 (N_22205,N_15882,N_16144);
nand U22206 (N_22206,N_19039,N_15303);
nand U22207 (N_22207,N_16574,N_16145);
nor U22208 (N_22208,N_19192,N_18335);
or U22209 (N_22209,N_15623,N_18910);
and U22210 (N_22210,N_19888,N_17021);
or U22211 (N_22211,N_15158,N_15449);
or U22212 (N_22212,N_15396,N_15353);
and U22213 (N_22213,N_18705,N_16674);
and U22214 (N_22214,N_16917,N_15884);
or U22215 (N_22215,N_15911,N_15543);
nor U22216 (N_22216,N_19344,N_16174);
nand U22217 (N_22217,N_16591,N_15470);
nor U22218 (N_22218,N_19258,N_16230);
or U22219 (N_22219,N_16976,N_17420);
nor U22220 (N_22220,N_16724,N_18662);
nand U22221 (N_22221,N_19694,N_16139);
nand U22222 (N_22222,N_18613,N_16141);
nand U22223 (N_22223,N_18157,N_16412);
nor U22224 (N_22224,N_18864,N_15081);
nor U22225 (N_22225,N_19456,N_18368);
nor U22226 (N_22226,N_17372,N_16229);
or U22227 (N_22227,N_19336,N_18782);
or U22228 (N_22228,N_18776,N_16387);
nor U22229 (N_22229,N_16479,N_19574);
and U22230 (N_22230,N_16707,N_16472);
nand U22231 (N_22231,N_15985,N_18164);
nor U22232 (N_22232,N_15534,N_17406);
and U22233 (N_22233,N_19122,N_18780);
nor U22234 (N_22234,N_19949,N_16137);
or U22235 (N_22235,N_15338,N_19922);
nor U22236 (N_22236,N_17075,N_15691);
or U22237 (N_22237,N_17230,N_18369);
nor U22238 (N_22238,N_18327,N_18061);
and U22239 (N_22239,N_18900,N_18972);
nor U22240 (N_22240,N_16848,N_16305);
and U22241 (N_22241,N_18769,N_16923);
nand U22242 (N_22242,N_19223,N_16853);
and U22243 (N_22243,N_15735,N_15586);
nor U22244 (N_22244,N_17563,N_16267);
or U22245 (N_22245,N_15434,N_17669);
and U22246 (N_22246,N_18845,N_17026);
nor U22247 (N_22247,N_19128,N_15604);
nand U22248 (N_22248,N_19831,N_15008);
and U22249 (N_22249,N_15582,N_15301);
and U22250 (N_22250,N_15684,N_19757);
or U22251 (N_22251,N_15035,N_17023);
nand U22252 (N_22252,N_18387,N_15938);
and U22253 (N_22253,N_18000,N_17377);
or U22254 (N_22254,N_16959,N_19619);
and U22255 (N_22255,N_15824,N_16370);
nand U22256 (N_22256,N_15592,N_18438);
nor U22257 (N_22257,N_15886,N_19133);
nand U22258 (N_22258,N_19800,N_17200);
and U22259 (N_22259,N_19182,N_16104);
nor U22260 (N_22260,N_15972,N_18223);
nand U22261 (N_22261,N_16766,N_17833);
or U22262 (N_22262,N_17022,N_16744);
and U22263 (N_22263,N_16583,N_19692);
or U22264 (N_22264,N_18740,N_17192);
nand U22265 (N_22265,N_17147,N_18992);
and U22266 (N_22266,N_19597,N_18472);
or U22267 (N_22267,N_18571,N_17248);
nor U22268 (N_22268,N_15706,N_18474);
nor U22269 (N_22269,N_17261,N_19077);
and U22270 (N_22270,N_16399,N_15997);
nor U22271 (N_22271,N_19542,N_18487);
xor U22272 (N_22272,N_18108,N_15657);
xnor U22273 (N_22273,N_18948,N_17977);
and U22274 (N_22274,N_17513,N_16243);
nor U22275 (N_22275,N_15124,N_18840);
nor U22276 (N_22276,N_15743,N_16905);
nand U22277 (N_22277,N_17149,N_17580);
or U22278 (N_22278,N_17416,N_19816);
nand U22279 (N_22279,N_15532,N_15239);
or U22280 (N_22280,N_18374,N_16263);
nor U22281 (N_22281,N_18975,N_16177);
nor U22282 (N_22282,N_18647,N_17626);
or U22283 (N_22283,N_18951,N_17301);
and U22284 (N_22284,N_18523,N_19801);
nor U22285 (N_22285,N_18790,N_17411);
nor U22286 (N_22286,N_18421,N_17719);
or U22287 (N_22287,N_18688,N_19257);
nor U22288 (N_22288,N_17699,N_19337);
or U22289 (N_22289,N_15056,N_17947);
nand U22290 (N_22290,N_17965,N_17404);
or U22291 (N_22291,N_18420,N_18458);
nand U22292 (N_22292,N_18524,N_16501);
nand U22293 (N_22293,N_15210,N_16730);
and U22294 (N_22294,N_19264,N_17010);
or U22295 (N_22295,N_15661,N_19869);
nor U22296 (N_22296,N_17162,N_18400);
nor U22297 (N_22297,N_15148,N_15128);
and U22298 (N_22298,N_15355,N_18346);
nor U22299 (N_22299,N_18795,N_19222);
nand U22300 (N_22300,N_15244,N_17204);
nor U22301 (N_22301,N_18260,N_19723);
nand U22302 (N_22302,N_17606,N_19338);
and U22303 (N_22303,N_15526,N_17408);
and U22304 (N_22304,N_17723,N_16329);
or U22305 (N_22305,N_19774,N_15389);
or U22306 (N_22306,N_16195,N_15122);
or U22307 (N_22307,N_15304,N_17507);
or U22308 (N_22308,N_15796,N_17000);
or U22309 (N_22309,N_19751,N_18981);
nor U22310 (N_22310,N_16131,N_19657);
and U22311 (N_22311,N_17995,N_17451);
and U22312 (N_22312,N_17594,N_19971);
or U22313 (N_22313,N_17468,N_18953);
and U22314 (N_22314,N_16172,N_19102);
nor U22315 (N_22315,N_17129,N_18963);
nor U22316 (N_22316,N_16887,N_18114);
nand U22317 (N_22317,N_17990,N_18693);
nor U22318 (N_22318,N_19058,N_18771);
or U22319 (N_22319,N_18805,N_15574);
or U22320 (N_22320,N_17555,N_17485);
nor U22321 (N_22321,N_17287,N_15162);
xor U22322 (N_22322,N_17139,N_15469);
nor U22323 (N_22323,N_18477,N_16276);
nand U22324 (N_22324,N_19030,N_15749);
or U22325 (N_22325,N_15497,N_15349);
and U22326 (N_22326,N_15435,N_16396);
and U22327 (N_22327,N_18677,N_17173);
and U22328 (N_22328,N_18186,N_18627);
or U22329 (N_22329,N_17061,N_15656);
or U22330 (N_22330,N_16727,N_19516);
or U22331 (N_22331,N_15024,N_19202);
or U22332 (N_22332,N_19513,N_16261);
or U22333 (N_22333,N_16327,N_16194);
and U22334 (N_22334,N_16827,N_19837);
or U22335 (N_22335,N_16240,N_15626);
nor U22336 (N_22336,N_16685,N_18269);
nor U22337 (N_22337,N_19585,N_19885);
nor U22338 (N_22338,N_19732,N_18582);
or U22339 (N_22339,N_15407,N_17564);
or U22340 (N_22340,N_16926,N_18675);
and U22341 (N_22341,N_17496,N_15619);
or U22342 (N_22342,N_19693,N_16031);
or U22343 (N_22343,N_16290,N_15731);
xnor U22344 (N_22344,N_18690,N_18748);
nor U22345 (N_22345,N_15099,N_18915);
nand U22346 (N_22346,N_15999,N_19627);
and U22347 (N_22347,N_18603,N_17775);
and U22348 (N_22348,N_16193,N_16460);
nand U22349 (N_22349,N_17410,N_18516);
nand U22350 (N_22350,N_19433,N_18797);
and U22351 (N_22351,N_18181,N_17419);
or U22352 (N_22352,N_15430,N_19847);
nor U22353 (N_22353,N_17417,N_18699);
and U22354 (N_22354,N_18682,N_18890);
nand U22355 (N_22355,N_18742,N_17974);
nor U22356 (N_22356,N_17603,N_18392);
and U22357 (N_22357,N_18877,N_18097);
nor U22358 (N_22358,N_18942,N_17269);
nor U22359 (N_22359,N_15147,N_15250);
and U22360 (N_22360,N_17796,N_16133);
nor U22361 (N_22361,N_18959,N_18527);
and U22362 (N_22362,N_17115,N_18015);
or U22363 (N_22363,N_17049,N_19394);
and U22364 (N_22364,N_19111,N_16752);
nor U22365 (N_22365,N_16510,N_15817);
nand U22366 (N_22366,N_15380,N_16861);
or U22367 (N_22367,N_18955,N_19205);
nand U22368 (N_22368,N_17259,N_17649);
or U22369 (N_22369,N_18793,N_18429);
nor U22370 (N_22370,N_18324,N_18821);
or U22371 (N_22371,N_18927,N_16016);
and U22372 (N_22372,N_18191,N_16613);
or U22373 (N_22373,N_16916,N_19802);
or U22374 (N_22374,N_17136,N_18428);
nand U22375 (N_22375,N_16765,N_19035);
nor U22376 (N_22376,N_15493,N_19386);
nand U22377 (N_22377,N_16087,N_18124);
nor U22378 (N_22378,N_17932,N_15283);
or U22379 (N_22379,N_18118,N_19491);
xnor U22380 (N_22380,N_17903,N_19817);
or U22381 (N_22381,N_19628,N_17088);
and U22382 (N_22382,N_19763,N_19522);
and U22383 (N_22383,N_16661,N_16814);
nand U22384 (N_22384,N_15568,N_18091);
nand U22385 (N_22385,N_16046,N_18694);
nand U22386 (N_22386,N_17802,N_19247);
nand U22387 (N_22387,N_17394,N_19996);
nand U22388 (N_22388,N_19704,N_19066);
nand U22389 (N_22389,N_16462,N_17784);
nor U22390 (N_22390,N_18935,N_17274);
nor U22391 (N_22391,N_16588,N_15487);
nor U22392 (N_22392,N_19079,N_15772);
nand U22393 (N_22393,N_19850,N_16213);
or U22394 (N_22394,N_19421,N_16980);
nand U22395 (N_22395,N_18402,N_19088);
or U22396 (N_22396,N_15660,N_19736);
nand U22397 (N_22397,N_17708,N_17214);
and U22398 (N_22398,N_18632,N_16295);
xnor U22399 (N_22399,N_18836,N_16636);
nor U22400 (N_22400,N_15181,N_19818);
nand U22401 (N_22401,N_17655,N_17487);
nand U22402 (N_22402,N_16300,N_19412);
nand U22403 (N_22403,N_16223,N_17768);
and U22404 (N_22404,N_18848,N_17877);
or U22405 (N_22405,N_19999,N_18032);
xor U22406 (N_22406,N_17423,N_16819);
nand U22407 (N_22407,N_15891,N_17027);
or U22408 (N_22408,N_16164,N_15214);
and U22409 (N_22409,N_15576,N_18304);
and U22410 (N_22410,N_16197,N_19387);
and U22411 (N_22411,N_15401,N_16218);
or U22412 (N_22412,N_17308,N_19702);
nor U22413 (N_22413,N_17748,N_19852);
nand U22414 (N_22414,N_18141,N_19769);
nand U22415 (N_22415,N_15673,N_15742);
nand U22416 (N_22416,N_15788,N_17846);
nand U22417 (N_22417,N_16872,N_17523);
or U22418 (N_22418,N_15120,N_17083);
nor U22419 (N_22419,N_15193,N_18205);
nor U22420 (N_22420,N_17804,N_16682);
nor U22421 (N_22421,N_15383,N_19459);
nand U22422 (N_22422,N_15249,N_15728);
nor U22423 (N_22423,N_15364,N_15902);
nand U22424 (N_22424,N_15375,N_17331);
and U22425 (N_22425,N_18641,N_18129);
or U22426 (N_22426,N_16953,N_18739);
nor U22427 (N_22427,N_18383,N_19709);
nor U22428 (N_22428,N_18484,N_17902);
or U22429 (N_22429,N_17567,N_15917);
nor U22430 (N_22430,N_15640,N_17345);
or U22431 (N_22431,N_19851,N_18190);
and U22432 (N_22432,N_18180,N_15243);
or U22433 (N_22433,N_15535,N_18116);
nand U22434 (N_22434,N_16882,N_17586);
nor U22435 (N_22435,N_19811,N_18898);
nand U22436 (N_22436,N_15033,N_19533);
or U22437 (N_22437,N_19244,N_19667);
nand U22438 (N_22438,N_19031,N_16273);
or U22439 (N_22439,N_15741,N_19590);
and U22440 (N_22440,N_19758,N_19217);
and U22441 (N_22441,N_15847,N_17253);
and U22442 (N_22442,N_16806,N_15361);
nor U22443 (N_22443,N_18858,N_16543);
nor U22444 (N_22444,N_17453,N_17014);
nor U22445 (N_22445,N_17120,N_18301);
or U22446 (N_22446,N_19790,N_17637);
and U22447 (N_22447,N_15385,N_19788);
or U22448 (N_22448,N_19577,N_15798);
nand U22449 (N_22449,N_16773,N_19738);
xnor U22450 (N_22450,N_16878,N_19604);
and U22451 (N_22451,N_15549,N_19772);
nor U22452 (N_22452,N_19684,N_19427);
nand U22453 (N_22453,N_15946,N_18762);
or U22454 (N_22454,N_19436,N_19400);
nor U22455 (N_22455,N_18966,N_15523);
and U22456 (N_22456,N_18300,N_16162);
or U22457 (N_22457,N_17704,N_16094);
nand U22458 (N_22458,N_15196,N_19897);
or U22459 (N_22459,N_18600,N_19191);
and U22460 (N_22460,N_19380,N_16485);
and U22461 (N_22461,N_15156,N_15803);
or U22462 (N_22462,N_17799,N_15213);
or U22463 (N_22463,N_15280,N_18964);
nand U22464 (N_22464,N_16324,N_15716);
nand U22465 (N_22465,N_16788,N_17318);
or U22466 (N_22466,N_15192,N_17045);
and U22467 (N_22467,N_19134,N_16314);
nor U22468 (N_22468,N_17167,N_17835);
or U22469 (N_22469,N_17020,N_18047);
nor U22470 (N_22470,N_17870,N_15447);
or U22471 (N_22471,N_18921,N_16952);
nor U22472 (N_22472,N_17755,N_18578);
xnor U22473 (N_22473,N_15409,N_15861);
nand U22474 (N_22474,N_16544,N_18841);
nand U22475 (N_22475,N_18302,N_19593);
nor U22476 (N_22476,N_18057,N_15705);
nor U22477 (N_22477,N_18506,N_15577);
and U22478 (N_22478,N_15183,N_19861);
nor U22479 (N_22479,N_17700,N_19397);
and U22480 (N_22480,N_17838,N_15955);
and U22481 (N_22481,N_19274,N_15699);
nand U22482 (N_22482,N_15322,N_19724);
nand U22483 (N_22483,N_15022,N_16587);
nor U22484 (N_22484,N_17209,N_17566);
or U22485 (N_22485,N_15107,N_19284);
nand U22486 (N_22486,N_19719,N_16941);
and U22487 (N_22487,N_19701,N_18268);
and U22488 (N_22488,N_15596,N_16681);
nand U22489 (N_22489,N_19130,N_16282);
and U22490 (N_22490,N_19484,N_18834);
xnor U22491 (N_22491,N_17391,N_18123);
and U22492 (N_22492,N_15724,N_19606);
nand U22493 (N_22493,N_16879,N_16034);
nor U22494 (N_22494,N_16532,N_16981);
or U22495 (N_22495,N_18755,N_18919);
nor U22496 (N_22496,N_16443,N_16552);
nor U22497 (N_22497,N_18650,N_18348);
nand U22498 (N_22498,N_19668,N_18590);
or U22499 (N_22499,N_16003,N_17415);
and U22500 (N_22500,N_16745,N_18391);
or U22501 (N_22501,N_17707,N_15501);
nor U22502 (N_22502,N_16778,N_17960);
nor U22503 (N_22503,N_16499,N_15436);
or U22504 (N_22504,N_15254,N_16803);
nor U22505 (N_22505,N_18372,N_15550);
or U22506 (N_22506,N_19490,N_15320);
or U22507 (N_22507,N_19196,N_15337);
and U22508 (N_22508,N_17533,N_18003);
nor U22509 (N_22509,N_17429,N_16134);
nor U22510 (N_22510,N_18141,N_15471);
and U22511 (N_22511,N_16246,N_19480);
nand U22512 (N_22512,N_19096,N_15682);
nor U22513 (N_22513,N_17661,N_19404);
nand U22514 (N_22514,N_19546,N_19110);
nand U22515 (N_22515,N_16408,N_17663);
nor U22516 (N_22516,N_16451,N_19920);
nand U22517 (N_22517,N_18042,N_15980);
and U22518 (N_22518,N_15515,N_15663);
nand U22519 (N_22519,N_15843,N_16049);
and U22520 (N_22520,N_17309,N_15186);
or U22521 (N_22521,N_16998,N_16545);
nand U22522 (N_22522,N_15427,N_18425);
nand U22523 (N_22523,N_16074,N_19160);
nor U22524 (N_22524,N_15595,N_15228);
nand U22525 (N_22525,N_18225,N_17140);
or U22526 (N_22526,N_18335,N_18314);
nor U22527 (N_22527,N_16239,N_16124);
or U22528 (N_22528,N_17869,N_16475);
nand U22529 (N_22529,N_18527,N_19373);
xnor U22530 (N_22530,N_17418,N_15199);
or U22531 (N_22531,N_18608,N_18991);
nand U22532 (N_22532,N_15190,N_17382);
or U22533 (N_22533,N_18873,N_15682);
or U22534 (N_22534,N_19072,N_19890);
or U22535 (N_22535,N_17687,N_19724);
nand U22536 (N_22536,N_19615,N_19632);
and U22537 (N_22537,N_19749,N_16707);
nor U22538 (N_22538,N_18436,N_19783);
nor U22539 (N_22539,N_18783,N_18076);
nor U22540 (N_22540,N_15375,N_18130);
nand U22541 (N_22541,N_15032,N_17199);
nor U22542 (N_22542,N_17482,N_17040);
nand U22543 (N_22543,N_18755,N_18720);
nor U22544 (N_22544,N_16665,N_17820);
or U22545 (N_22545,N_19047,N_18411);
nor U22546 (N_22546,N_18746,N_16065);
nand U22547 (N_22547,N_15949,N_19682);
and U22548 (N_22548,N_17429,N_18319);
or U22549 (N_22549,N_17884,N_15300);
nor U22550 (N_22550,N_15154,N_18788);
and U22551 (N_22551,N_18555,N_17384);
and U22552 (N_22552,N_18069,N_18875);
nor U22553 (N_22553,N_17482,N_17249);
or U22554 (N_22554,N_15278,N_18632);
and U22555 (N_22555,N_16860,N_15732);
and U22556 (N_22556,N_15595,N_19805);
and U22557 (N_22557,N_19348,N_15689);
and U22558 (N_22558,N_17903,N_17119);
nor U22559 (N_22559,N_17238,N_18475);
nand U22560 (N_22560,N_17570,N_16450);
nor U22561 (N_22561,N_18169,N_18225);
and U22562 (N_22562,N_16497,N_17320);
nor U22563 (N_22563,N_18998,N_19608);
and U22564 (N_22564,N_16358,N_19475);
and U22565 (N_22565,N_19697,N_18944);
or U22566 (N_22566,N_15151,N_15644);
nand U22567 (N_22567,N_18783,N_18459);
nor U22568 (N_22568,N_19889,N_17092);
and U22569 (N_22569,N_19921,N_18163);
and U22570 (N_22570,N_19235,N_17201);
and U22571 (N_22571,N_15888,N_19752);
and U22572 (N_22572,N_15515,N_19060);
or U22573 (N_22573,N_18024,N_17498);
nand U22574 (N_22574,N_17927,N_19990);
and U22575 (N_22575,N_16041,N_16133);
nand U22576 (N_22576,N_15798,N_17556);
nor U22577 (N_22577,N_15641,N_17321);
nor U22578 (N_22578,N_15994,N_19286);
or U22579 (N_22579,N_16249,N_16602);
or U22580 (N_22580,N_17410,N_15841);
and U22581 (N_22581,N_15805,N_18529);
and U22582 (N_22582,N_17613,N_15634);
nor U22583 (N_22583,N_15914,N_19933);
nor U22584 (N_22584,N_15984,N_18806);
and U22585 (N_22585,N_16629,N_18846);
nand U22586 (N_22586,N_19131,N_19900);
nand U22587 (N_22587,N_18047,N_19871);
or U22588 (N_22588,N_15058,N_15846);
nor U22589 (N_22589,N_15269,N_19130);
or U22590 (N_22590,N_18118,N_15718);
nand U22591 (N_22591,N_18104,N_18191);
and U22592 (N_22592,N_17457,N_18346);
nor U22593 (N_22593,N_17923,N_17900);
and U22594 (N_22594,N_18355,N_18356);
nor U22595 (N_22595,N_17673,N_19957);
or U22596 (N_22596,N_18131,N_18642);
or U22597 (N_22597,N_18955,N_18502);
nand U22598 (N_22598,N_17903,N_18567);
and U22599 (N_22599,N_15761,N_19352);
or U22600 (N_22600,N_15528,N_15126);
nand U22601 (N_22601,N_18685,N_16035);
nor U22602 (N_22602,N_15559,N_16383);
or U22603 (N_22603,N_15052,N_18468);
or U22604 (N_22604,N_18801,N_16411);
nand U22605 (N_22605,N_19724,N_17498);
nor U22606 (N_22606,N_18002,N_17595);
or U22607 (N_22607,N_19358,N_15958);
nor U22608 (N_22608,N_16002,N_16917);
nand U22609 (N_22609,N_19890,N_19157);
nor U22610 (N_22610,N_16170,N_17286);
nand U22611 (N_22611,N_16134,N_16125);
and U22612 (N_22612,N_18811,N_18033);
nand U22613 (N_22613,N_17204,N_16179);
nor U22614 (N_22614,N_18134,N_16511);
nor U22615 (N_22615,N_18122,N_15919);
nor U22616 (N_22616,N_18520,N_17227);
nor U22617 (N_22617,N_18003,N_17125);
and U22618 (N_22618,N_19111,N_16065);
nand U22619 (N_22619,N_19355,N_15530);
and U22620 (N_22620,N_18187,N_15109);
and U22621 (N_22621,N_17963,N_16181);
nor U22622 (N_22622,N_16145,N_15168);
nand U22623 (N_22623,N_18083,N_15705);
nor U22624 (N_22624,N_15922,N_17067);
or U22625 (N_22625,N_17425,N_15641);
nor U22626 (N_22626,N_15127,N_15506);
and U22627 (N_22627,N_17367,N_19477);
or U22628 (N_22628,N_19215,N_18257);
or U22629 (N_22629,N_16842,N_16898);
nand U22630 (N_22630,N_17476,N_19374);
nand U22631 (N_22631,N_16108,N_19342);
or U22632 (N_22632,N_18156,N_18887);
or U22633 (N_22633,N_16316,N_15771);
and U22634 (N_22634,N_19837,N_16900);
nand U22635 (N_22635,N_16139,N_16768);
nand U22636 (N_22636,N_18059,N_17071);
nor U22637 (N_22637,N_16670,N_16245);
nand U22638 (N_22638,N_16932,N_19031);
and U22639 (N_22639,N_19549,N_18913);
nand U22640 (N_22640,N_15711,N_17536);
or U22641 (N_22641,N_18190,N_15991);
or U22642 (N_22642,N_19504,N_16680);
and U22643 (N_22643,N_18040,N_15171);
nor U22644 (N_22644,N_17038,N_18561);
nor U22645 (N_22645,N_15444,N_18092);
or U22646 (N_22646,N_15954,N_19258);
nor U22647 (N_22647,N_15854,N_17042);
nor U22648 (N_22648,N_15451,N_18085);
nor U22649 (N_22649,N_19097,N_16733);
nand U22650 (N_22650,N_17156,N_15942);
nand U22651 (N_22651,N_19287,N_19028);
nor U22652 (N_22652,N_15849,N_18525);
nand U22653 (N_22653,N_18164,N_16230);
and U22654 (N_22654,N_17116,N_15021);
and U22655 (N_22655,N_16026,N_19759);
or U22656 (N_22656,N_17212,N_17846);
and U22657 (N_22657,N_17452,N_17038);
or U22658 (N_22658,N_17751,N_16177);
nor U22659 (N_22659,N_15648,N_17838);
or U22660 (N_22660,N_16486,N_18701);
or U22661 (N_22661,N_15763,N_17134);
and U22662 (N_22662,N_18922,N_15126);
nor U22663 (N_22663,N_15729,N_17197);
nand U22664 (N_22664,N_18458,N_15128);
nor U22665 (N_22665,N_19616,N_16262);
and U22666 (N_22666,N_16463,N_17904);
xnor U22667 (N_22667,N_17696,N_19583);
and U22668 (N_22668,N_16622,N_19597);
and U22669 (N_22669,N_17620,N_16647);
or U22670 (N_22670,N_17600,N_17518);
or U22671 (N_22671,N_19851,N_17455);
nor U22672 (N_22672,N_18111,N_18237);
nor U22673 (N_22673,N_19852,N_17114);
and U22674 (N_22674,N_19305,N_19015);
and U22675 (N_22675,N_16697,N_18267);
or U22676 (N_22676,N_16662,N_19061);
or U22677 (N_22677,N_17609,N_17317);
nand U22678 (N_22678,N_16456,N_19845);
nor U22679 (N_22679,N_16700,N_19188);
or U22680 (N_22680,N_17767,N_16231);
nand U22681 (N_22681,N_18177,N_19017);
and U22682 (N_22682,N_17897,N_18513);
nor U22683 (N_22683,N_19523,N_19409);
or U22684 (N_22684,N_18788,N_18251);
or U22685 (N_22685,N_15007,N_18755);
and U22686 (N_22686,N_17100,N_15523);
nand U22687 (N_22687,N_18546,N_18564);
nor U22688 (N_22688,N_15136,N_15996);
nor U22689 (N_22689,N_16014,N_16286);
or U22690 (N_22690,N_19914,N_18916);
or U22691 (N_22691,N_17270,N_19950);
nand U22692 (N_22692,N_18917,N_15387);
nand U22693 (N_22693,N_18661,N_16312);
or U22694 (N_22694,N_16287,N_17603);
or U22695 (N_22695,N_18181,N_17867);
and U22696 (N_22696,N_16949,N_18508);
or U22697 (N_22697,N_17370,N_18686);
or U22698 (N_22698,N_15693,N_18621);
and U22699 (N_22699,N_19795,N_18346);
or U22700 (N_22700,N_15219,N_18567);
and U22701 (N_22701,N_19110,N_16678);
or U22702 (N_22702,N_15099,N_15566);
nand U22703 (N_22703,N_16627,N_19982);
or U22704 (N_22704,N_18116,N_19162);
and U22705 (N_22705,N_17291,N_17160);
and U22706 (N_22706,N_18422,N_18492);
nand U22707 (N_22707,N_18806,N_18951);
nor U22708 (N_22708,N_16700,N_15732);
nor U22709 (N_22709,N_15281,N_19034);
or U22710 (N_22710,N_15031,N_15632);
or U22711 (N_22711,N_19701,N_19491);
nor U22712 (N_22712,N_16021,N_15376);
nor U22713 (N_22713,N_17309,N_18947);
or U22714 (N_22714,N_17035,N_17447);
nand U22715 (N_22715,N_15080,N_16976);
nand U22716 (N_22716,N_15297,N_16641);
nor U22717 (N_22717,N_19541,N_18237);
nor U22718 (N_22718,N_19961,N_17515);
and U22719 (N_22719,N_17087,N_15883);
nand U22720 (N_22720,N_18135,N_17305);
nor U22721 (N_22721,N_17346,N_16054);
nand U22722 (N_22722,N_15057,N_17829);
nor U22723 (N_22723,N_18928,N_16165);
nand U22724 (N_22724,N_15534,N_18137);
or U22725 (N_22725,N_15760,N_18369);
or U22726 (N_22726,N_16263,N_15558);
or U22727 (N_22727,N_19925,N_19309);
nor U22728 (N_22728,N_16262,N_16093);
and U22729 (N_22729,N_17289,N_17337);
or U22730 (N_22730,N_16072,N_18040);
nor U22731 (N_22731,N_19691,N_16588);
nor U22732 (N_22732,N_15408,N_15236);
nand U22733 (N_22733,N_19018,N_17819);
and U22734 (N_22734,N_19462,N_19734);
nand U22735 (N_22735,N_19956,N_19127);
nand U22736 (N_22736,N_19555,N_16734);
nor U22737 (N_22737,N_17983,N_16897);
or U22738 (N_22738,N_18626,N_19566);
and U22739 (N_22739,N_17504,N_19455);
and U22740 (N_22740,N_16816,N_17201);
and U22741 (N_22741,N_17717,N_16726);
or U22742 (N_22742,N_19909,N_18259);
or U22743 (N_22743,N_16127,N_18970);
and U22744 (N_22744,N_17126,N_18947);
nand U22745 (N_22745,N_19529,N_17686);
nand U22746 (N_22746,N_15358,N_18855);
or U22747 (N_22747,N_16741,N_18275);
or U22748 (N_22748,N_18350,N_19258);
and U22749 (N_22749,N_19343,N_16871);
nand U22750 (N_22750,N_18938,N_16646);
nand U22751 (N_22751,N_16698,N_16017);
nor U22752 (N_22752,N_15184,N_18006);
nor U22753 (N_22753,N_15601,N_17532);
nand U22754 (N_22754,N_18785,N_15530);
nor U22755 (N_22755,N_19879,N_18739);
and U22756 (N_22756,N_15546,N_15878);
or U22757 (N_22757,N_17329,N_16924);
xnor U22758 (N_22758,N_19798,N_16600);
nor U22759 (N_22759,N_18145,N_17738);
nor U22760 (N_22760,N_15638,N_15109);
nor U22761 (N_22761,N_15293,N_17077);
nand U22762 (N_22762,N_16129,N_15157);
nand U22763 (N_22763,N_15800,N_18081);
or U22764 (N_22764,N_19186,N_15761);
and U22765 (N_22765,N_16922,N_18260);
and U22766 (N_22766,N_17354,N_15248);
nand U22767 (N_22767,N_16255,N_19695);
nand U22768 (N_22768,N_17506,N_19887);
and U22769 (N_22769,N_19137,N_18654);
and U22770 (N_22770,N_17066,N_16198);
nand U22771 (N_22771,N_16399,N_19378);
or U22772 (N_22772,N_19733,N_17284);
or U22773 (N_22773,N_16516,N_17524);
or U22774 (N_22774,N_18769,N_15629);
nor U22775 (N_22775,N_19605,N_18463);
and U22776 (N_22776,N_16474,N_18464);
nand U22777 (N_22777,N_16992,N_18269);
or U22778 (N_22778,N_17627,N_17493);
and U22779 (N_22779,N_15228,N_15618);
and U22780 (N_22780,N_17829,N_18222);
or U22781 (N_22781,N_18660,N_15560);
or U22782 (N_22782,N_19802,N_19123);
and U22783 (N_22783,N_15418,N_19098);
xor U22784 (N_22784,N_19073,N_19628);
nand U22785 (N_22785,N_15611,N_16367);
or U22786 (N_22786,N_16845,N_18510);
or U22787 (N_22787,N_18331,N_18320);
nand U22788 (N_22788,N_15862,N_16940);
nor U22789 (N_22789,N_16878,N_17320);
nor U22790 (N_22790,N_17556,N_18417);
or U22791 (N_22791,N_15209,N_18347);
nor U22792 (N_22792,N_18089,N_17328);
nor U22793 (N_22793,N_15717,N_18470);
or U22794 (N_22794,N_17477,N_16957);
or U22795 (N_22795,N_19526,N_16420);
and U22796 (N_22796,N_16467,N_16473);
and U22797 (N_22797,N_19696,N_19838);
and U22798 (N_22798,N_16413,N_15276);
nor U22799 (N_22799,N_15538,N_15378);
nand U22800 (N_22800,N_17983,N_18319);
and U22801 (N_22801,N_15089,N_15317);
or U22802 (N_22802,N_15840,N_19153);
nor U22803 (N_22803,N_16377,N_18327);
and U22804 (N_22804,N_17314,N_16960);
or U22805 (N_22805,N_18034,N_19848);
and U22806 (N_22806,N_18149,N_18882);
nor U22807 (N_22807,N_15035,N_17788);
and U22808 (N_22808,N_18980,N_16362);
and U22809 (N_22809,N_16655,N_16526);
nand U22810 (N_22810,N_15874,N_19557);
nand U22811 (N_22811,N_18405,N_17089);
nor U22812 (N_22812,N_15464,N_15124);
nand U22813 (N_22813,N_16956,N_15792);
and U22814 (N_22814,N_19487,N_18657);
or U22815 (N_22815,N_19569,N_17919);
nor U22816 (N_22816,N_17640,N_16805);
nand U22817 (N_22817,N_17748,N_17059);
nor U22818 (N_22818,N_15446,N_16273);
xnor U22819 (N_22819,N_18626,N_19106);
or U22820 (N_22820,N_17061,N_17022);
and U22821 (N_22821,N_18992,N_18788);
nand U22822 (N_22822,N_16840,N_16050);
nand U22823 (N_22823,N_17301,N_19936);
and U22824 (N_22824,N_15483,N_15152);
and U22825 (N_22825,N_19683,N_17340);
and U22826 (N_22826,N_18757,N_18450);
or U22827 (N_22827,N_15256,N_19366);
nor U22828 (N_22828,N_17218,N_17828);
or U22829 (N_22829,N_16309,N_15194);
or U22830 (N_22830,N_18086,N_15905);
or U22831 (N_22831,N_15185,N_17193);
nor U22832 (N_22832,N_15836,N_19034);
or U22833 (N_22833,N_19232,N_19225);
nand U22834 (N_22834,N_17373,N_18577);
or U22835 (N_22835,N_18743,N_16276);
nand U22836 (N_22836,N_19365,N_15941);
nor U22837 (N_22837,N_19832,N_16394);
nor U22838 (N_22838,N_19342,N_17546);
nand U22839 (N_22839,N_19704,N_16363);
nor U22840 (N_22840,N_15049,N_17259);
nand U22841 (N_22841,N_19518,N_19333);
nor U22842 (N_22842,N_17728,N_15122);
and U22843 (N_22843,N_19838,N_15114);
and U22844 (N_22844,N_17837,N_15867);
and U22845 (N_22845,N_17510,N_15299);
or U22846 (N_22846,N_19752,N_19516);
nor U22847 (N_22847,N_17288,N_18969);
nor U22848 (N_22848,N_16937,N_17855);
and U22849 (N_22849,N_19073,N_16225);
and U22850 (N_22850,N_19728,N_17462);
nor U22851 (N_22851,N_16432,N_16129);
nor U22852 (N_22852,N_19025,N_16930);
nor U22853 (N_22853,N_16325,N_17032);
nand U22854 (N_22854,N_15699,N_16547);
nand U22855 (N_22855,N_17355,N_18303);
nor U22856 (N_22856,N_18769,N_18235);
or U22857 (N_22857,N_17982,N_19284);
nor U22858 (N_22858,N_15200,N_19193);
nor U22859 (N_22859,N_16912,N_16958);
nand U22860 (N_22860,N_18263,N_18548);
xnor U22861 (N_22861,N_15961,N_15302);
nor U22862 (N_22862,N_18797,N_18737);
and U22863 (N_22863,N_17182,N_19031);
or U22864 (N_22864,N_15418,N_16348);
nand U22865 (N_22865,N_16014,N_17218);
or U22866 (N_22866,N_18194,N_17413);
xnor U22867 (N_22867,N_19643,N_18931);
nor U22868 (N_22868,N_17040,N_15886);
or U22869 (N_22869,N_17485,N_15548);
or U22870 (N_22870,N_16447,N_17026);
nand U22871 (N_22871,N_18293,N_19547);
and U22872 (N_22872,N_18177,N_19474);
nand U22873 (N_22873,N_15212,N_17978);
or U22874 (N_22874,N_15562,N_15603);
and U22875 (N_22875,N_17909,N_18359);
and U22876 (N_22876,N_18930,N_17271);
nor U22877 (N_22877,N_15473,N_18108);
or U22878 (N_22878,N_16397,N_17784);
nand U22879 (N_22879,N_18178,N_18279);
or U22880 (N_22880,N_17309,N_18676);
or U22881 (N_22881,N_15375,N_15528);
nor U22882 (N_22882,N_18740,N_17827);
nand U22883 (N_22883,N_16445,N_17872);
and U22884 (N_22884,N_19528,N_16626);
and U22885 (N_22885,N_18335,N_18724);
nor U22886 (N_22886,N_18609,N_19245);
nor U22887 (N_22887,N_19132,N_19284);
and U22888 (N_22888,N_17772,N_18291);
nand U22889 (N_22889,N_15609,N_15348);
and U22890 (N_22890,N_17628,N_19841);
and U22891 (N_22891,N_18848,N_18668);
and U22892 (N_22892,N_18265,N_19760);
nor U22893 (N_22893,N_15505,N_19819);
nor U22894 (N_22894,N_19285,N_18363);
and U22895 (N_22895,N_15336,N_19944);
nor U22896 (N_22896,N_17243,N_19267);
or U22897 (N_22897,N_15653,N_19210);
nand U22898 (N_22898,N_18020,N_18935);
and U22899 (N_22899,N_18853,N_18642);
or U22900 (N_22900,N_19838,N_18435);
and U22901 (N_22901,N_16708,N_19899);
and U22902 (N_22902,N_18420,N_18855);
nand U22903 (N_22903,N_19664,N_19016);
nand U22904 (N_22904,N_18503,N_19782);
or U22905 (N_22905,N_19580,N_16985);
nand U22906 (N_22906,N_18097,N_19878);
nor U22907 (N_22907,N_15594,N_18527);
and U22908 (N_22908,N_16687,N_18531);
nand U22909 (N_22909,N_15883,N_15925);
nand U22910 (N_22910,N_15379,N_18075);
and U22911 (N_22911,N_15583,N_19524);
nor U22912 (N_22912,N_16529,N_17808);
or U22913 (N_22913,N_17451,N_19194);
nand U22914 (N_22914,N_15325,N_16467);
nor U22915 (N_22915,N_19491,N_15166);
nor U22916 (N_22916,N_18199,N_19417);
nor U22917 (N_22917,N_15768,N_19089);
nor U22918 (N_22918,N_19068,N_18240);
or U22919 (N_22919,N_16919,N_15553);
nand U22920 (N_22920,N_19478,N_18192);
nand U22921 (N_22921,N_17396,N_16474);
nor U22922 (N_22922,N_16686,N_15351);
and U22923 (N_22923,N_17470,N_15283);
nor U22924 (N_22924,N_18596,N_15346);
nand U22925 (N_22925,N_18499,N_16383);
nand U22926 (N_22926,N_15996,N_18496);
and U22927 (N_22927,N_18435,N_17661);
nor U22928 (N_22928,N_15350,N_17610);
nor U22929 (N_22929,N_16946,N_19244);
or U22930 (N_22930,N_18641,N_19327);
or U22931 (N_22931,N_15704,N_17721);
and U22932 (N_22932,N_15337,N_18778);
nor U22933 (N_22933,N_19895,N_19769);
nand U22934 (N_22934,N_19419,N_17819);
and U22935 (N_22935,N_15829,N_16298);
and U22936 (N_22936,N_16886,N_16149);
nand U22937 (N_22937,N_17832,N_18500);
or U22938 (N_22938,N_17353,N_15815);
nand U22939 (N_22939,N_16895,N_19006);
nor U22940 (N_22940,N_15761,N_16800);
and U22941 (N_22941,N_16596,N_15665);
nor U22942 (N_22942,N_15639,N_16652);
nor U22943 (N_22943,N_17494,N_16180);
nand U22944 (N_22944,N_16611,N_17303);
nand U22945 (N_22945,N_17747,N_17896);
or U22946 (N_22946,N_18722,N_18802);
nand U22947 (N_22947,N_18288,N_15773);
xnor U22948 (N_22948,N_16593,N_17020);
nand U22949 (N_22949,N_17806,N_19089);
and U22950 (N_22950,N_18913,N_16785);
and U22951 (N_22951,N_15695,N_17608);
xnor U22952 (N_22952,N_17966,N_16014);
and U22953 (N_22953,N_17172,N_19957);
nor U22954 (N_22954,N_19269,N_19300);
or U22955 (N_22955,N_17430,N_18154);
and U22956 (N_22956,N_17861,N_19210);
nor U22957 (N_22957,N_17964,N_15173);
and U22958 (N_22958,N_19915,N_16049);
or U22959 (N_22959,N_19234,N_17779);
or U22960 (N_22960,N_17376,N_15047);
and U22961 (N_22961,N_19330,N_18701);
nor U22962 (N_22962,N_15264,N_19024);
nor U22963 (N_22963,N_15228,N_16316);
or U22964 (N_22964,N_19035,N_17909);
and U22965 (N_22965,N_17322,N_17690);
or U22966 (N_22966,N_16317,N_16761);
and U22967 (N_22967,N_15144,N_18423);
nor U22968 (N_22968,N_17133,N_16066);
nor U22969 (N_22969,N_17266,N_16115);
or U22970 (N_22970,N_18222,N_15074);
and U22971 (N_22971,N_15803,N_17001);
and U22972 (N_22972,N_16048,N_17415);
nand U22973 (N_22973,N_19530,N_17744);
and U22974 (N_22974,N_19525,N_19082);
nor U22975 (N_22975,N_16125,N_15735);
or U22976 (N_22976,N_19231,N_15049);
or U22977 (N_22977,N_17078,N_17381);
and U22978 (N_22978,N_17726,N_16446);
or U22979 (N_22979,N_16240,N_17681);
nor U22980 (N_22980,N_18523,N_17846);
or U22981 (N_22981,N_19727,N_19879);
or U22982 (N_22982,N_17064,N_19362);
nand U22983 (N_22983,N_19762,N_19709);
or U22984 (N_22984,N_17952,N_18120);
nand U22985 (N_22985,N_18875,N_19225);
nand U22986 (N_22986,N_19740,N_18224);
nand U22987 (N_22987,N_19455,N_19632);
or U22988 (N_22988,N_19811,N_15775);
nor U22989 (N_22989,N_15905,N_18739);
and U22990 (N_22990,N_17773,N_16261);
nand U22991 (N_22991,N_18263,N_18845);
or U22992 (N_22992,N_15682,N_19578);
nand U22993 (N_22993,N_17541,N_18508);
and U22994 (N_22994,N_17886,N_16377);
nand U22995 (N_22995,N_16459,N_15685);
nor U22996 (N_22996,N_18446,N_17848);
and U22997 (N_22997,N_19213,N_19877);
or U22998 (N_22998,N_19509,N_16646);
and U22999 (N_22999,N_18003,N_19410);
nand U23000 (N_23000,N_19882,N_15962);
or U23001 (N_23001,N_16553,N_19309);
nor U23002 (N_23002,N_18564,N_19743);
nor U23003 (N_23003,N_16457,N_16862);
and U23004 (N_23004,N_18694,N_17810);
nor U23005 (N_23005,N_19823,N_18211);
or U23006 (N_23006,N_18864,N_19606);
or U23007 (N_23007,N_19401,N_16658);
and U23008 (N_23008,N_18613,N_18393);
nor U23009 (N_23009,N_15654,N_18760);
nor U23010 (N_23010,N_15533,N_19392);
nand U23011 (N_23011,N_19045,N_17798);
and U23012 (N_23012,N_19130,N_15231);
or U23013 (N_23013,N_17443,N_16648);
or U23014 (N_23014,N_18997,N_19892);
nor U23015 (N_23015,N_18770,N_18484);
and U23016 (N_23016,N_17086,N_15165);
or U23017 (N_23017,N_16810,N_19010);
nor U23018 (N_23018,N_19491,N_16550);
or U23019 (N_23019,N_16680,N_19146);
nand U23020 (N_23020,N_16272,N_19611);
nor U23021 (N_23021,N_15419,N_17932);
and U23022 (N_23022,N_17821,N_16565);
and U23023 (N_23023,N_17687,N_16290);
and U23024 (N_23024,N_18874,N_16660);
or U23025 (N_23025,N_19609,N_17486);
or U23026 (N_23026,N_15248,N_16010);
or U23027 (N_23027,N_17184,N_19865);
nor U23028 (N_23028,N_18793,N_18137);
nand U23029 (N_23029,N_19519,N_16775);
nor U23030 (N_23030,N_18525,N_15175);
and U23031 (N_23031,N_16076,N_15953);
nand U23032 (N_23032,N_19282,N_19924);
nor U23033 (N_23033,N_17417,N_15174);
or U23034 (N_23034,N_16300,N_18822);
nand U23035 (N_23035,N_19306,N_17119);
and U23036 (N_23036,N_18216,N_15091);
or U23037 (N_23037,N_18957,N_15795);
or U23038 (N_23038,N_18820,N_19076);
nand U23039 (N_23039,N_15743,N_17232);
or U23040 (N_23040,N_15026,N_15553);
nor U23041 (N_23041,N_18770,N_17828);
nand U23042 (N_23042,N_15152,N_18803);
and U23043 (N_23043,N_17447,N_19730);
nor U23044 (N_23044,N_15909,N_18035);
and U23045 (N_23045,N_15919,N_16777);
or U23046 (N_23046,N_15762,N_18024);
nand U23047 (N_23047,N_19947,N_17902);
and U23048 (N_23048,N_16386,N_16456);
nand U23049 (N_23049,N_17423,N_19758);
nand U23050 (N_23050,N_18941,N_19834);
nand U23051 (N_23051,N_16978,N_19668);
or U23052 (N_23052,N_16568,N_15780);
and U23053 (N_23053,N_19734,N_19372);
and U23054 (N_23054,N_17954,N_17910);
and U23055 (N_23055,N_15278,N_15689);
and U23056 (N_23056,N_17373,N_19482);
nor U23057 (N_23057,N_19357,N_15649);
and U23058 (N_23058,N_19091,N_17354);
xnor U23059 (N_23059,N_16570,N_18919);
and U23060 (N_23060,N_19682,N_17618);
nand U23061 (N_23061,N_18669,N_19208);
nor U23062 (N_23062,N_16492,N_16597);
xor U23063 (N_23063,N_16114,N_16599);
nand U23064 (N_23064,N_18428,N_16173);
nand U23065 (N_23065,N_15998,N_19510);
nor U23066 (N_23066,N_19031,N_17450);
or U23067 (N_23067,N_15337,N_19126);
nand U23068 (N_23068,N_17984,N_16808);
and U23069 (N_23069,N_19098,N_15967);
nand U23070 (N_23070,N_16179,N_19927);
or U23071 (N_23071,N_17193,N_19017);
nand U23072 (N_23072,N_15213,N_18159);
and U23073 (N_23073,N_18959,N_19042);
and U23074 (N_23074,N_15987,N_18158);
nor U23075 (N_23075,N_19414,N_18575);
or U23076 (N_23076,N_17190,N_19961);
or U23077 (N_23077,N_19053,N_18811);
nand U23078 (N_23078,N_15793,N_19773);
nor U23079 (N_23079,N_16784,N_17553);
nand U23080 (N_23080,N_17405,N_16428);
nand U23081 (N_23081,N_15615,N_15472);
and U23082 (N_23082,N_17651,N_16149);
nand U23083 (N_23083,N_16558,N_15942);
or U23084 (N_23084,N_16624,N_15499);
nor U23085 (N_23085,N_17683,N_16786);
and U23086 (N_23086,N_18860,N_16987);
nor U23087 (N_23087,N_19778,N_17333);
nor U23088 (N_23088,N_16836,N_17471);
or U23089 (N_23089,N_17026,N_18360);
or U23090 (N_23090,N_19381,N_16918);
or U23091 (N_23091,N_15616,N_18543);
xnor U23092 (N_23092,N_16323,N_19824);
nor U23093 (N_23093,N_15106,N_19595);
or U23094 (N_23094,N_15166,N_16519);
nand U23095 (N_23095,N_19898,N_19896);
nor U23096 (N_23096,N_17501,N_19224);
or U23097 (N_23097,N_15942,N_18532);
nand U23098 (N_23098,N_17216,N_16208);
nor U23099 (N_23099,N_16615,N_19207);
nand U23100 (N_23100,N_19616,N_19149);
and U23101 (N_23101,N_19840,N_18844);
nor U23102 (N_23102,N_18294,N_15849);
nand U23103 (N_23103,N_15906,N_15487);
or U23104 (N_23104,N_18257,N_15919);
or U23105 (N_23105,N_16364,N_18565);
nand U23106 (N_23106,N_17995,N_19258);
nor U23107 (N_23107,N_17020,N_15785);
and U23108 (N_23108,N_18961,N_16952);
or U23109 (N_23109,N_18662,N_19501);
and U23110 (N_23110,N_17252,N_17904);
nor U23111 (N_23111,N_16003,N_18622);
and U23112 (N_23112,N_17284,N_17703);
and U23113 (N_23113,N_17266,N_19346);
and U23114 (N_23114,N_16544,N_15370);
or U23115 (N_23115,N_16690,N_18329);
nand U23116 (N_23116,N_17362,N_16188);
or U23117 (N_23117,N_16170,N_15873);
nand U23118 (N_23118,N_17790,N_18263);
or U23119 (N_23119,N_18365,N_17607);
or U23120 (N_23120,N_17904,N_16276);
and U23121 (N_23121,N_16977,N_15841);
nor U23122 (N_23122,N_17614,N_17703);
nand U23123 (N_23123,N_18183,N_17967);
nor U23124 (N_23124,N_16492,N_17822);
and U23125 (N_23125,N_19819,N_17106);
nor U23126 (N_23126,N_18719,N_19236);
or U23127 (N_23127,N_17118,N_16726);
nor U23128 (N_23128,N_17233,N_18749);
or U23129 (N_23129,N_15448,N_17647);
or U23130 (N_23130,N_19361,N_16332);
and U23131 (N_23131,N_19143,N_18498);
nor U23132 (N_23132,N_15071,N_15866);
nor U23133 (N_23133,N_18292,N_16275);
and U23134 (N_23134,N_17730,N_17700);
or U23135 (N_23135,N_17526,N_17611);
and U23136 (N_23136,N_18705,N_18088);
and U23137 (N_23137,N_17844,N_16439);
and U23138 (N_23138,N_17338,N_17465);
nor U23139 (N_23139,N_16815,N_16553);
nand U23140 (N_23140,N_17502,N_15049);
nor U23141 (N_23141,N_17121,N_18431);
or U23142 (N_23142,N_16981,N_17029);
nor U23143 (N_23143,N_18368,N_15320);
or U23144 (N_23144,N_16720,N_16468);
nand U23145 (N_23145,N_16071,N_19816);
nor U23146 (N_23146,N_18204,N_19295);
and U23147 (N_23147,N_19673,N_19125);
or U23148 (N_23148,N_17197,N_15168);
nand U23149 (N_23149,N_15782,N_15269);
xnor U23150 (N_23150,N_18005,N_16474);
and U23151 (N_23151,N_16535,N_17602);
nand U23152 (N_23152,N_15814,N_18448);
or U23153 (N_23153,N_17566,N_18824);
or U23154 (N_23154,N_17044,N_19934);
and U23155 (N_23155,N_17824,N_19168);
or U23156 (N_23156,N_18525,N_19669);
nor U23157 (N_23157,N_18243,N_15052);
and U23158 (N_23158,N_15914,N_16388);
nand U23159 (N_23159,N_17177,N_18345);
or U23160 (N_23160,N_15228,N_19562);
nor U23161 (N_23161,N_16124,N_15115);
and U23162 (N_23162,N_18876,N_18954);
or U23163 (N_23163,N_19358,N_19991);
or U23164 (N_23164,N_17536,N_17081);
and U23165 (N_23165,N_19584,N_18977);
nor U23166 (N_23166,N_19770,N_19174);
nand U23167 (N_23167,N_17166,N_16619);
nand U23168 (N_23168,N_15123,N_18161);
and U23169 (N_23169,N_19810,N_17311);
nor U23170 (N_23170,N_17868,N_15148);
nand U23171 (N_23171,N_17953,N_19643);
nor U23172 (N_23172,N_15405,N_15798);
or U23173 (N_23173,N_15784,N_15579);
nor U23174 (N_23174,N_16528,N_19571);
nand U23175 (N_23175,N_17816,N_16398);
and U23176 (N_23176,N_17440,N_19283);
or U23177 (N_23177,N_18609,N_17549);
nor U23178 (N_23178,N_16785,N_18039);
nand U23179 (N_23179,N_16822,N_18243);
and U23180 (N_23180,N_19268,N_18330);
nand U23181 (N_23181,N_15248,N_19645);
nand U23182 (N_23182,N_18139,N_15356);
nand U23183 (N_23183,N_16087,N_15841);
nor U23184 (N_23184,N_15645,N_15932);
or U23185 (N_23185,N_16679,N_15466);
nor U23186 (N_23186,N_15969,N_17797);
nor U23187 (N_23187,N_16854,N_18420);
nor U23188 (N_23188,N_19497,N_15713);
nand U23189 (N_23189,N_16451,N_17849);
nand U23190 (N_23190,N_16262,N_19313);
and U23191 (N_23191,N_15734,N_17009);
or U23192 (N_23192,N_17661,N_18816);
nand U23193 (N_23193,N_17916,N_17435);
or U23194 (N_23194,N_15876,N_16975);
and U23195 (N_23195,N_18288,N_16417);
or U23196 (N_23196,N_15900,N_18779);
and U23197 (N_23197,N_15247,N_19918);
nor U23198 (N_23198,N_19478,N_16589);
and U23199 (N_23199,N_15971,N_16115);
nor U23200 (N_23200,N_15343,N_15000);
or U23201 (N_23201,N_15215,N_15073);
nor U23202 (N_23202,N_15761,N_19685);
nor U23203 (N_23203,N_17881,N_17922);
nand U23204 (N_23204,N_17927,N_17433);
nor U23205 (N_23205,N_17608,N_19164);
nand U23206 (N_23206,N_18752,N_17506);
or U23207 (N_23207,N_17397,N_16137);
nand U23208 (N_23208,N_18902,N_15028);
nor U23209 (N_23209,N_17113,N_17270);
nand U23210 (N_23210,N_15755,N_17601);
nor U23211 (N_23211,N_15923,N_19980);
nand U23212 (N_23212,N_16849,N_17282);
and U23213 (N_23213,N_17678,N_19051);
nand U23214 (N_23214,N_16118,N_17443);
nand U23215 (N_23215,N_18524,N_15290);
and U23216 (N_23216,N_19024,N_19175);
nor U23217 (N_23217,N_19172,N_18186);
nor U23218 (N_23218,N_15707,N_18094);
nand U23219 (N_23219,N_15577,N_17736);
or U23220 (N_23220,N_19322,N_19533);
and U23221 (N_23221,N_17840,N_19375);
or U23222 (N_23222,N_19351,N_18167);
nor U23223 (N_23223,N_16237,N_19014);
and U23224 (N_23224,N_17358,N_19668);
and U23225 (N_23225,N_15671,N_16645);
and U23226 (N_23226,N_15058,N_17715);
nand U23227 (N_23227,N_15206,N_19370);
nand U23228 (N_23228,N_19255,N_16383);
nand U23229 (N_23229,N_19707,N_18615);
and U23230 (N_23230,N_16953,N_17626);
and U23231 (N_23231,N_18309,N_19366);
or U23232 (N_23232,N_19177,N_17464);
nor U23233 (N_23233,N_17793,N_17020);
and U23234 (N_23234,N_15699,N_15179);
and U23235 (N_23235,N_19855,N_15199);
nor U23236 (N_23236,N_18347,N_18970);
nand U23237 (N_23237,N_16184,N_16138);
or U23238 (N_23238,N_16821,N_18665);
nor U23239 (N_23239,N_19504,N_17493);
or U23240 (N_23240,N_15227,N_15773);
or U23241 (N_23241,N_18654,N_17203);
and U23242 (N_23242,N_17811,N_18349);
or U23243 (N_23243,N_16710,N_19659);
and U23244 (N_23244,N_16189,N_16799);
and U23245 (N_23245,N_17996,N_16662);
and U23246 (N_23246,N_18828,N_15623);
nor U23247 (N_23247,N_16793,N_18133);
and U23248 (N_23248,N_17681,N_16521);
nand U23249 (N_23249,N_17505,N_18224);
and U23250 (N_23250,N_19837,N_19391);
nor U23251 (N_23251,N_15379,N_16809);
nand U23252 (N_23252,N_15371,N_17172);
or U23253 (N_23253,N_17549,N_15556);
and U23254 (N_23254,N_17208,N_17341);
nand U23255 (N_23255,N_15108,N_18038);
nor U23256 (N_23256,N_16836,N_15560);
or U23257 (N_23257,N_16023,N_16576);
or U23258 (N_23258,N_19319,N_16108);
and U23259 (N_23259,N_19159,N_17015);
nand U23260 (N_23260,N_19459,N_16642);
nand U23261 (N_23261,N_15550,N_16760);
nand U23262 (N_23262,N_18946,N_18407);
or U23263 (N_23263,N_18361,N_19961);
and U23264 (N_23264,N_18744,N_15949);
or U23265 (N_23265,N_16026,N_19643);
nor U23266 (N_23266,N_19509,N_18667);
and U23267 (N_23267,N_16164,N_16096);
nand U23268 (N_23268,N_17946,N_16330);
or U23269 (N_23269,N_18538,N_15455);
and U23270 (N_23270,N_15440,N_19041);
and U23271 (N_23271,N_18606,N_15576);
nand U23272 (N_23272,N_19651,N_15407);
nor U23273 (N_23273,N_17832,N_18523);
and U23274 (N_23274,N_18117,N_18605);
and U23275 (N_23275,N_16902,N_18145);
nor U23276 (N_23276,N_16127,N_19550);
nor U23277 (N_23277,N_18834,N_15121);
and U23278 (N_23278,N_19771,N_15713);
nand U23279 (N_23279,N_19881,N_16936);
and U23280 (N_23280,N_18642,N_15853);
nand U23281 (N_23281,N_18800,N_16204);
nor U23282 (N_23282,N_19242,N_19268);
nor U23283 (N_23283,N_19074,N_16590);
or U23284 (N_23284,N_15422,N_17246);
or U23285 (N_23285,N_16109,N_17185);
or U23286 (N_23286,N_19447,N_19200);
or U23287 (N_23287,N_19693,N_16905);
nor U23288 (N_23288,N_19217,N_16611);
nor U23289 (N_23289,N_18787,N_17984);
nand U23290 (N_23290,N_17315,N_16399);
or U23291 (N_23291,N_17049,N_16479);
and U23292 (N_23292,N_18445,N_17085);
and U23293 (N_23293,N_17604,N_16551);
or U23294 (N_23294,N_15119,N_19823);
nor U23295 (N_23295,N_19280,N_19609);
and U23296 (N_23296,N_15172,N_18709);
or U23297 (N_23297,N_17987,N_18560);
or U23298 (N_23298,N_17302,N_19087);
and U23299 (N_23299,N_17239,N_15311);
or U23300 (N_23300,N_19787,N_15779);
nor U23301 (N_23301,N_16400,N_16270);
nor U23302 (N_23302,N_17573,N_17982);
nor U23303 (N_23303,N_16002,N_19436);
nand U23304 (N_23304,N_15213,N_15751);
nor U23305 (N_23305,N_15746,N_15857);
nand U23306 (N_23306,N_15306,N_15964);
nor U23307 (N_23307,N_19442,N_18432);
nor U23308 (N_23308,N_18675,N_15612);
and U23309 (N_23309,N_16178,N_17408);
nand U23310 (N_23310,N_18385,N_15913);
or U23311 (N_23311,N_19857,N_16272);
and U23312 (N_23312,N_15384,N_19557);
nand U23313 (N_23313,N_15723,N_15553);
nor U23314 (N_23314,N_15498,N_17678);
and U23315 (N_23315,N_17441,N_19937);
and U23316 (N_23316,N_16409,N_15975);
or U23317 (N_23317,N_15031,N_15302);
nand U23318 (N_23318,N_16431,N_17224);
and U23319 (N_23319,N_17701,N_18668);
nand U23320 (N_23320,N_16966,N_18168);
nand U23321 (N_23321,N_17114,N_18263);
and U23322 (N_23322,N_19112,N_19810);
nand U23323 (N_23323,N_17759,N_16029);
and U23324 (N_23324,N_17444,N_18718);
and U23325 (N_23325,N_17327,N_19682);
nor U23326 (N_23326,N_18632,N_17178);
nor U23327 (N_23327,N_19863,N_15698);
nand U23328 (N_23328,N_19945,N_17813);
nor U23329 (N_23329,N_17257,N_16007);
and U23330 (N_23330,N_19999,N_19610);
nor U23331 (N_23331,N_17358,N_19483);
nand U23332 (N_23332,N_19618,N_16555);
nor U23333 (N_23333,N_15740,N_16273);
nand U23334 (N_23334,N_19671,N_16042);
nor U23335 (N_23335,N_19144,N_16221);
nand U23336 (N_23336,N_19638,N_15646);
nor U23337 (N_23337,N_15507,N_19142);
or U23338 (N_23338,N_16530,N_19543);
or U23339 (N_23339,N_15880,N_19066);
and U23340 (N_23340,N_17253,N_17316);
and U23341 (N_23341,N_17141,N_18908);
or U23342 (N_23342,N_15565,N_16579);
and U23343 (N_23343,N_19233,N_16088);
or U23344 (N_23344,N_15641,N_18207);
or U23345 (N_23345,N_15261,N_18870);
and U23346 (N_23346,N_15296,N_17939);
nor U23347 (N_23347,N_17087,N_19512);
nand U23348 (N_23348,N_18604,N_16803);
nor U23349 (N_23349,N_17485,N_17535);
nand U23350 (N_23350,N_15863,N_16805);
or U23351 (N_23351,N_18339,N_15047);
or U23352 (N_23352,N_19387,N_16049);
nor U23353 (N_23353,N_18303,N_19011);
nand U23354 (N_23354,N_15116,N_19332);
and U23355 (N_23355,N_16305,N_17892);
and U23356 (N_23356,N_17181,N_15544);
nor U23357 (N_23357,N_16452,N_17019);
or U23358 (N_23358,N_15466,N_17176);
and U23359 (N_23359,N_18938,N_17009);
and U23360 (N_23360,N_15559,N_19553);
nand U23361 (N_23361,N_16390,N_19908);
or U23362 (N_23362,N_15667,N_16411);
or U23363 (N_23363,N_17355,N_18061);
or U23364 (N_23364,N_15447,N_19891);
or U23365 (N_23365,N_16844,N_18668);
nor U23366 (N_23366,N_19909,N_16695);
and U23367 (N_23367,N_18973,N_19866);
nand U23368 (N_23368,N_16143,N_17915);
and U23369 (N_23369,N_16631,N_16233);
and U23370 (N_23370,N_19673,N_18658);
nand U23371 (N_23371,N_16090,N_19020);
nor U23372 (N_23372,N_18631,N_17164);
nor U23373 (N_23373,N_18814,N_16317);
and U23374 (N_23374,N_19752,N_17605);
or U23375 (N_23375,N_17062,N_18896);
and U23376 (N_23376,N_16310,N_17572);
nor U23377 (N_23377,N_16481,N_16277);
or U23378 (N_23378,N_15085,N_15442);
nor U23379 (N_23379,N_18922,N_17959);
and U23380 (N_23380,N_15826,N_17925);
or U23381 (N_23381,N_19554,N_15793);
and U23382 (N_23382,N_15252,N_18311);
nor U23383 (N_23383,N_16496,N_15147);
nor U23384 (N_23384,N_19500,N_17336);
and U23385 (N_23385,N_16627,N_18937);
nand U23386 (N_23386,N_19283,N_17889);
or U23387 (N_23387,N_16519,N_17354);
and U23388 (N_23388,N_18015,N_16554);
and U23389 (N_23389,N_18481,N_19028);
nor U23390 (N_23390,N_16376,N_15343);
nor U23391 (N_23391,N_16746,N_16014);
nor U23392 (N_23392,N_19046,N_18388);
nor U23393 (N_23393,N_17574,N_16830);
and U23394 (N_23394,N_16204,N_15210);
or U23395 (N_23395,N_17124,N_18880);
nor U23396 (N_23396,N_16484,N_16812);
and U23397 (N_23397,N_16122,N_15311);
nor U23398 (N_23398,N_18453,N_19298);
or U23399 (N_23399,N_17158,N_16041);
nand U23400 (N_23400,N_18931,N_15424);
or U23401 (N_23401,N_16929,N_15077);
and U23402 (N_23402,N_19435,N_19957);
xnor U23403 (N_23403,N_18497,N_17597);
nor U23404 (N_23404,N_17570,N_16759);
or U23405 (N_23405,N_16470,N_18215);
nor U23406 (N_23406,N_19166,N_17945);
nor U23407 (N_23407,N_16501,N_17818);
nor U23408 (N_23408,N_18573,N_16725);
or U23409 (N_23409,N_19075,N_19828);
and U23410 (N_23410,N_16566,N_19360);
or U23411 (N_23411,N_18006,N_18118);
or U23412 (N_23412,N_18472,N_17473);
and U23413 (N_23413,N_16062,N_15606);
nand U23414 (N_23414,N_18788,N_17844);
nand U23415 (N_23415,N_18204,N_17354);
nand U23416 (N_23416,N_19002,N_17089);
or U23417 (N_23417,N_15234,N_17099);
nand U23418 (N_23418,N_15416,N_16149);
and U23419 (N_23419,N_16570,N_17416);
nand U23420 (N_23420,N_18393,N_16638);
and U23421 (N_23421,N_19773,N_15508);
nor U23422 (N_23422,N_15424,N_19946);
nand U23423 (N_23423,N_16771,N_16654);
nand U23424 (N_23424,N_18544,N_19922);
or U23425 (N_23425,N_17382,N_16963);
nand U23426 (N_23426,N_18579,N_16511);
nor U23427 (N_23427,N_19491,N_15386);
nand U23428 (N_23428,N_19268,N_16777);
nor U23429 (N_23429,N_18622,N_19016);
nor U23430 (N_23430,N_16336,N_15549);
and U23431 (N_23431,N_16794,N_16256);
and U23432 (N_23432,N_19514,N_16643);
or U23433 (N_23433,N_17738,N_19652);
and U23434 (N_23434,N_15933,N_15941);
nor U23435 (N_23435,N_17202,N_16112);
nor U23436 (N_23436,N_15972,N_15381);
nor U23437 (N_23437,N_16350,N_19482);
and U23438 (N_23438,N_15256,N_16368);
nand U23439 (N_23439,N_17199,N_16569);
or U23440 (N_23440,N_16325,N_18472);
or U23441 (N_23441,N_16854,N_17229);
nand U23442 (N_23442,N_19455,N_15379);
xor U23443 (N_23443,N_18939,N_17258);
or U23444 (N_23444,N_19812,N_15911);
or U23445 (N_23445,N_16548,N_18419);
nor U23446 (N_23446,N_16288,N_17795);
nor U23447 (N_23447,N_15940,N_18170);
and U23448 (N_23448,N_18603,N_18191);
xnor U23449 (N_23449,N_19703,N_17177);
nand U23450 (N_23450,N_16929,N_18603);
and U23451 (N_23451,N_16711,N_17470);
or U23452 (N_23452,N_15348,N_16179);
nor U23453 (N_23453,N_16709,N_16739);
or U23454 (N_23454,N_15398,N_15991);
or U23455 (N_23455,N_19765,N_17803);
and U23456 (N_23456,N_15939,N_19682);
and U23457 (N_23457,N_15664,N_19802);
and U23458 (N_23458,N_16499,N_18631);
nand U23459 (N_23459,N_18624,N_16794);
nand U23460 (N_23460,N_17572,N_15406);
or U23461 (N_23461,N_19684,N_19379);
nor U23462 (N_23462,N_16311,N_16150);
nor U23463 (N_23463,N_16831,N_16230);
and U23464 (N_23464,N_19270,N_19116);
or U23465 (N_23465,N_17594,N_17610);
nand U23466 (N_23466,N_19840,N_16581);
or U23467 (N_23467,N_19229,N_17491);
and U23468 (N_23468,N_18817,N_16699);
nand U23469 (N_23469,N_15527,N_16000);
or U23470 (N_23470,N_15665,N_16258);
nor U23471 (N_23471,N_15651,N_16606);
and U23472 (N_23472,N_17693,N_18020);
nand U23473 (N_23473,N_15487,N_19859);
or U23474 (N_23474,N_19892,N_19698);
nand U23475 (N_23475,N_19795,N_19734);
nor U23476 (N_23476,N_16018,N_17669);
and U23477 (N_23477,N_16764,N_16666);
and U23478 (N_23478,N_18253,N_16920);
nand U23479 (N_23479,N_17074,N_17690);
and U23480 (N_23480,N_19808,N_16820);
or U23481 (N_23481,N_18557,N_17758);
or U23482 (N_23482,N_17135,N_19315);
and U23483 (N_23483,N_19834,N_15665);
nand U23484 (N_23484,N_18756,N_15354);
nor U23485 (N_23485,N_17248,N_18937);
or U23486 (N_23486,N_16748,N_17789);
nor U23487 (N_23487,N_16448,N_19271);
nor U23488 (N_23488,N_19677,N_17080);
nor U23489 (N_23489,N_19673,N_19496);
and U23490 (N_23490,N_16159,N_17312);
nand U23491 (N_23491,N_17471,N_15900);
or U23492 (N_23492,N_19934,N_16888);
or U23493 (N_23493,N_16666,N_16390);
and U23494 (N_23494,N_15342,N_15754);
nor U23495 (N_23495,N_15467,N_17199);
nand U23496 (N_23496,N_19097,N_17935);
or U23497 (N_23497,N_18079,N_18999);
or U23498 (N_23498,N_19766,N_16964);
nand U23499 (N_23499,N_16027,N_17107);
nor U23500 (N_23500,N_18862,N_15360);
and U23501 (N_23501,N_16141,N_16721);
nor U23502 (N_23502,N_17329,N_16983);
nor U23503 (N_23503,N_18531,N_16373);
and U23504 (N_23504,N_16541,N_19238);
and U23505 (N_23505,N_18499,N_17281);
or U23506 (N_23506,N_18473,N_19198);
and U23507 (N_23507,N_17054,N_18530);
or U23508 (N_23508,N_17082,N_18300);
nand U23509 (N_23509,N_19066,N_16602);
nand U23510 (N_23510,N_15228,N_17800);
nor U23511 (N_23511,N_16724,N_17030);
and U23512 (N_23512,N_19229,N_17507);
nand U23513 (N_23513,N_18291,N_19373);
and U23514 (N_23514,N_17408,N_19136);
nand U23515 (N_23515,N_17727,N_15033);
nand U23516 (N_23516,N_19518,N_15267);
or U23517 (N_23517,N_19854,N_15746);
and U23518 (N_23518,N_16386,N_16882);
and U23519 (N_23519,N_19878,N_17592);
or U23520 (N_23520,N_15984,N_16255);
nand U23521 (N_23521,N_15979,N_16432);
nand U23522 (N_23522,N_15115,N_16393);
and U23523 (N_23523,N_19261,N_15536);
or U23524 (N_23524,N_17085,N_17228);
nor U23525 (N_23525,N_19116,N_19280);
or U23526 (N_23526,N_16717,N_15232);
or U23527 (N_23527,N_15924,N_16008);
nand U23528 (N_23528,N_17804,N_16877);
nand U23529 (N_23529,N_18215,N_16268);
or U23530 (N_23530,N_15689,N_19014);
and U23531 (N_23531,N_16140,N_19986);
nor U23532 (N_23532,N_17946,N_19148);
or U23533 (N_23533,N_16479,N_16496);
and U23534 (N_23534,N_18049,N_19205);
or U23535 (N_23535,N_19193,N_16373);
nor U23536 (N_23536,N_16227,N_18305);
or U23537 (N_23537,N_16357,N_17843);
and U23538 (N_23538,N_16647,N_15859);
nor U23539 (N_23539,N_17138,N_16396);
nor U23540 (N_23540,N_18579,N_18474);
xor U23541 (N_23541,N_15867,N_19959);
nor U23542 (N_23542,N_18755,N_16128);
and U23543 (N_23543,N_18146,N_15632);
nand U23544 (N_23544,N_15975,N_15662);
nor U23545 (N_23545,N_19223,N_15615);
and U23546 (N_23546,N_16845,N_17186);
or U23547 (N_23547,N_16706,N_19295);
or U23548 (N_23548,N_16774,N_18501);
nand U23549 (N_23549,N_19573,N_19822);
nand U23550 (N_23550,N_16932,N_18815);
or U23551 (N_23551,N_17529,N_15669);
nor U23552 (N_23552,N_17358,N_18178);
nor U23553 (N_23553,N_19381,N_15351);
and U23554 (N_23554,N_16170,N_19205);
and U23555 (N_23555,N_17938,N_15688);
or U23556 (N_23556,N_15108,N_19288);
nor U23557 (N_23557,N_15093,N_18190);
or U23558 (N_23558,N_16012,N_17940);
and U23559 (N_23559,N_18032,N_17993);
or U23560 (N_23560,N_16963,N_17504);
or U23561 (N_23561,N_18102,N_17130);
or U23562 (N_23562,N_18113,N_18236);
or U23563 (N_23563,N_17391,N_15609);
nand U23564 (N_23564,N_18153,N_17657);
or U23565 (N_23565,N_18881,N_15674);
or U23566 (N_23566,N_17091,N_16429);
and U23567 (N_23567,N_17639,N_19566);
nor U23568 (N_23568,N_17308,N_16894);
nand U23569 (N_23569,N_16417,N_19136);
or U23570 (N_23570,N_18304,N_17447);
and U23571 (N_23571,N_18016,N_19416);
nor U23572 (N_23572,N_18455,N_18980);
nand U23573 (N_23573,N_19786,N_15073);
and U23574 (N_23574,N_16927,N_15208);
nor U23575 (N_23575,N_17659,N_19284);
nand U23576 (N_23576,N_16764,N_17408);
and U23577 (N_23577,N_19638,N_16057);
nand U23578 (N_23578,N_19019,N_18151);
nor U23579 (N_23579,N_15407,N_19207);
or U23580 (N_23580,N_18690,N_18136);
nand U23581 (N_23581,N_15189,N_16711);
and U23582 (N_23582,N_19840,N_15567);
and U23583 (N_23583,N_15908,N_17948);
nor U23584 (N_23584,N_16592,N_19147);
nor U23585 (N_23585,N_19365,N_18682);
or U23586 (N_23586,N_19943,N_18993);
or U23587 (N_23587,N_16822,N_18608);
nor U23588 (N_23588,N_17505,N_15776);
nor U23589 (N_23589,N_16975,N_19031);
or U23590 (N_23590,N_15086,N_17481);
and U23591 (N_23591,N_18044,N_16832);
nor U23592 (N_23592,N_16829,N_19708);
xor U23593 (N_23593,N_17857,N_19997);
nor U23594 (N_23594,N_17453,N_15959);
or U23595 (N_23595,N_16599,N_15702);
and U23596 (N_23596,N_19286,N_19062);
nor U23597 (N_23597,N_16508,N_19868);
nand U23598 (N_23598,N_16143,N_19418);
and U23599 (N_23599,N_19930,N_16497);
or U23600 (N_23600,N_16249,N_16262);
nor U23601 (N_23601,N_18207,N_15890);
or U23602 (N_23602,N_16381,N_16255);
nand U23603 (N_23603,N_17957,N_19665);
nand U23604 (N_23604,N_19850,N_17911);
and U23605 (N_23605,N_15544,N_17100);
nor U23606 (N_23606,N_18691,N_19953);
nor U23607 (N_23607,N_17853,N_17361);
nor U23608 (N_23608,N_17629,N_16884);
nand U23609 (N_23609,N_18869,N_17644);
or U23610 (N_23610,N_17159,N_17266);
or U23611 (N_23611,N_19882,N_19568);
nor U23612 (N_23612,N_17816,N_18467);
or U23613 (N_23613,N_18139,N_15846);
nor U23614 (N_23614,N_15003,N_18577);
and U23615 (N_23615,N_16612,N_19263);
or U23616 (N_23616,N_19466,N_17671);
or U23617 (N_23617,N_18712,N_16438);
and U23618 (N_23618,N_19446,N_16850);
nor U23619 (N_23619,N_16664,N_15830);
nand U23620 (N_23620,N_16607,N_18680);
or U23621 (N_23621,N_16156,N_19369);
xor U23622 (N_23622,N_17570,N_17020);
nand U23623 (N_23623,N_19582,N_15385);
nor U23624 (N_23624,N_19071,N_17168);
nor U23625 (N_23625,N_19313,N_17785);
and U23626 (N_23626,N_16758,N_15202);
and U23627 (N_23627,N_19814,N_19597);
nor U23628 (N_23628,N_17149,N_16940);
and U23629 (N_23629,N_17060,N_16043);
and U23630 (N_23630,N_17794,N_15560);
or U23631 (N_23631,N_15768,N_16367);
or U23632 (N_23632,N_16840,N_19869);
or U23633 (N_23633,N_19073,N_17692);
nor U23634 (N_23634,N_16443,N_15458);
or U23635 (N_23635,N_17299,N_17199);
nand U23636 (N_23636,N_18640,N_16604);
xnor U23637 (N_23637,N_16636,N_18334);
and U23638 (N_23638,N_17148,N_18941);
nor U23639 (N_23639,N_19159,N_16065);
nand U23640 (N_23640,N_16166,N_17228);
or U23641 (N_23641,N_16334,N_18529);
or U23642 (N_23642,N_18892,N_19910);
nor U23643 (N_23643,N_18733,N_18130);
nor U23644 (N_23644,N_18456,N_15917);
nor U23645 (N_23645,N_17715,N_18088);
nand U23646 (N_23646,N_15741,N_17694);
or U23647 (N_23647,N_15127,N_15077);
nand U23648 (N_23648,N_17882,N_18835);
and U23649 (N_23649,N_16885,N_15291);
nor U23650 (N_23650,N_17446,N_17257);
xor U23651 (N_23651,N_16356,N_18923);
nor U23652 (N_23652,N_15903,N_16173);
nor U23653 (N_23653,N_18010,N_16947);
nor U23654 (N_23654,N_17350,N_15542);
nor U23655 (N_23655,N_16079,N_19408);
nor U23656 (N_23656,N_18322,N_17209);
or U23657 (N_23657,N_15015,N_16165);
nand U23658 (N_23658,N_16968,N_16310);
or U23659 (N_23659,N_17122,N_17705);
nand U23660 (N_23660,N_16628,N_19786);
nand U23661 (N_23661,N_18700,N_17426);
and U23662 (N_23662,N_16869,N_18998);
nand U23663 (N_23663,N_18494,N_19001);
or U23664 (N_23664,N_16702,N_18331);
nand U23665 (N_23665,N_17973,N_18070);
nand U23666 (N_23666,N_16297,N_17297);
nor U23667 (N_23667,N_19070,N_18303);
or U23668 (N_23668,N_17038,N_17806);
or U23669 (N_23669,N_17771,N_19035);
or U23670 (N_23670,N_19791,N_18088);
nand U23671 (N_23671,N_17997,N_18592);
nand U23672 (N_23672,N_17635,N_17167);
and U23673 (N_23673,N_15356,N_19876);
nor U23674 (N_23674,N_15609,N_15290);
or U23675 (N_23675,N_15452,N_17779);
and U23676 (N_23676,N_15685,N_17765);
nand U23677 (N_23677,N_15239,N_16849);
and U23678 (N_23678,N_16276,N_18931);
nor U23679 (N_23679,N_18346,N_19091);
nand U23680 (N_23680,N_17085,N_18553);
or U23681 (N_23681,N_19580,N_17878);
and U23682 (N_23682,N_19608,N_18964);
nand U23683 (N_23683,N_19826,N_15360);
and U23684 (N_23684,N_17209,N_18634);
and U23685 (N_23685,N_16544,N_15968);
or U23686 (N_23686,N_18660,N_19822);
nor U23687 (N_23687,N_18916,N_18555);
nand U23688 (N_23688,N_16984,N_18656);
nor U23689 (N_23689,N_15211,N_15919);
or U23690 (N_23690,N_17111,N_19734);
nor U23691 (N_23691,N_18521,N_15735);
nand U23692 (N_23692,N_18366,N_19885);
or U23693 (N_23693,N_18277,N_15376);
nor U23694 (N_23694,N_16729,N_18379);
xor U23695 (N_23695,N_16900,N_19779);
nand U23696 (N_23696,N_19170,N_19421);
or U23697 (N_23697,N_19892,N_19244);
nor U23698 (N_23698,N_19436,N_15365);
nor U23699 (N_23699,N_16708,N_17692);
or U23700 (N_23700,N_17324,N_19031);
and U23701 (N_23701,N_16559,N_19235);
nor U23702 (N_23702,N_19620,N_16745);
and U23703 (N_23703,N_18410,N_16287);
nor U23704 (N_23704,N_19768,N_18800);
or U23705 (N_23705,N_18550,N_16626);
or U23706 (N_23706,N_19636,N_15216);
nand U23707 (N_23707,N_19250,N_17858);
nand U23708 (N_23708,N_15282,N_19385);
and U23709 (N_23709,N_15852,N_15408);
nand U23710 (N_23710,N_15941,N_19202);
xor U23711 (N_23711,N_19309,N_19179);
nand U23712 (N_23712,N_17112,N_18106);
nor U23713 (N_23713,N_19805,N_17744);
and U23714 (N_23714,N_16976,N_19222);
or U23715 (N_23715,N_16972,N_16785);
nand U23716 (N_23716,N_19988,N_19787);
nor U23717 (N_23717,N_18515,N_16500);
or U23718 (N_23718,N_18295,N_19867);
nand U23719 (N_23719,N_15870,N_19842);
nand U23720 (N_23720,N_15237,N_18660);
nand U23721 (N_23721,N_19786,N_17837);
or U23722 (N_23722,N_16693,N_18894);
nor U23723 (N_23723,N_16678,N_15096);
nand U23724 (N_23724,N_18276,N_17738);
or U23725 (N_23725,N_17478,N_19717);
or U23726 (N_23726,N_15641,N_17773);
nor U23727 (N_23727,N_15830,N_18390);
and U23728 (N_23728,N_17872,N_16768);
and U23729 (N_23729,N_18855,N_19232);
nor U23730 (N_23730,N_19569,N_16566);
or U23731 (N_23731,N_19597,N_16543);
nor U23732 (N_23732,N_15558,N_19454);
nor U23733 (N_23733,N_16105,N_17503);
nor U23734 (N_23734,N_17534,N_15212);
or U23735 (N_23735,N_15361,N_18007);
or U23736 (N_23736,N_15117,N_18893);
nand U23737 (N_23737,N_16833,N_19618);
and U23738 (N_23738,N_17056,N_18572);
or U23739 (N_23739,N_16973,N_16530);
nand U23740 (N_23740,N_19320,N_17933);
xnor U23741 (N_23741,N_16037,N_16376);
nor U23742 (N_23742,N_16487,N_19760);
nor U23743 (N_23743,N_19715,N_17087);
nor U23744 (N_23744,N_15022,N_18605);
nor U23745 (N_23745,N_15889,N_19228);
and U23746 (N_23746,N_15485,N_17628);
nor U23747 (N_23747,N_19167,N_16555);
and U23748 (N_23748,N_18941,N_17591);
or U23749 (N_23749,N_18906,N_18061);
nand U23750 (N_23750,N_15779,N_15865);
or U23751 (N_23751,N_15266,N_17464);
nand U23752 (N_23752,N_18995,N_16403);
nand U23753 (N_23753,N_18306,N_17735);
and U23754 (N_23754,N_18880,N_16694);
nand U23755 (N_23755,N_16904,N_18769);
and U23756 (N_23756,N_15686,N_19643);
and U23757 (N_23757,N_16815,N_17932);
nor U23758 (N_23758,N_16831,N_17915);
or U23759 (N_23759,N_17578,N_19205);
nand U23760 (N_23760,N_18040,N_15949);
nor U23761 (N_23761,N_16835,N_15350);
and U23762 (N_23762,N_19053,N_18772);
nor U23763 (N_23763,N_17562,N_16654);
or U23764 (N_23764,N_19899,N_17487);
or U23765 (N_23765,N_19700,N_18108);
and U23766 (N_23766,N_15378,N_18115);
and U23767 (N_23767,N_16488,N_18961);
nand U23768 (N_23768,N_15457,N_16375);
or U23769 (N_23769,N_17862,N_19024);
or U23770 (N_23770,N_19106,N_16936);
nor U23771 (N_23771,N_15031,N_18456);
nand U23772 (N_23772,N_17966,N_16846);
nor U23773 (N_23773,N_19451,N_16023);
or U23774 (N_23774,N_19423,N_16594);
and U23775 (N_23775,N_18887,N_15787);
and U23776 (N_23776,N_18385,N_18857);
or U23777 (N_23777,N_19812,N_15802);
or U23778 (N_23778,N_18131,N_19877);
nand U23779 (N_23779,N_17187,N_17933);
nor U23780 (N_23780,N_17354,N_19946);
nor U23781 (N_23781,N_19145,N_19141);
nor U23782 (N_23782,N_19403,N_18105);
nor U23783 (N_23783,N_16096,N_19014);
and U23784 (N_23784,N_15913,N_15727);
and U23785 (N_23785,N_17535,N_15410);
and U23786 (N_23786,N_19400,N_15128);
xor U23787 (N_23787,N_17023,N_15597);
nor U23788 (N_23788,N_15079,N_18597);
or U23789 (N_23789,N_15110,N_16432);
nor U23790 (N_23790,N_15986,N_19928);
nor U23791 (N_23791,N_15848,N_15855);
nor U23792 (N_23792,N_15133,N_15340);
nor U23793 (N_23793,N_16593,N_16079);
nand U23794 (N_23794,N_17167,N_17720);
or U23795 (N_23795,N_17411,N_16648);
nand U23796 (N_23796,N_15189,N_19349);
and U23797 (N_23797,N_18470,N_18479);
nand U23798 (N_23798,N_18734,N_19355);
nand U23799 (N_23799,N_16866,N_17861);
or U23800 (N_23800,N_17185,N_17772);
nand U23801 (N_23801,N_15327,N_17281);
nand U23802 (N_23802,N_19995,N_16654);
nand U23803 (N_23803,N_17291,N_18094);
nand U23804 (N_23804,N_18026,N_19555);
xnor U23805 (N_23805,N_18977,N_17736);
and U23806 (N_23806,N_19167,N_15143);
nand U23807 (N_23807,N_18095,N_16339);
nor U23808 (N_23808,N_17614,N_19904);
nor U23809 (N_23809,N_16893,N_17364);
nand U23810 (N_23810,N_19005,N_18895);
or U23811 (N_23811,N_19207,N_18248);
or U23812 (N_23812,N_15200,N_16415);
or U23813 (N_23813,N_19736,N_18330);
nor U23814 (N_23814,N_19753,N_17118);
nor U23815 (N_23815,N_16279,N_17749);
nand U23816 (N_23816,N_15455,N_17519);
or U23817 (N_23817,N_18230,N_16281);
nand U23818 (N_23818,N_17077,N_15077);
nor U23819 (N_23819,N_15935,N_19392);
nor U23820 (N_23820,N_19250,N_18160);
or U23821 (N_23821,N_15375,N_17394);
or U23822 (N_23822,N_16960,N_16286);
nand U23823 (N_23823,N_18953,N_17087);
nand U23824 (N_23824,N_17484,N_17595);
and U23825 (N_23825,N_18894,N_17373);
nor U23826 (N_23826,N_17949,N_17260);
and U23827 (N_23827,N_19213,N_19532);
or U23828 (N_23828,N_17307,N_16685);
nand U23829 (N_23829,N_17391,N_19710);
or U23830 (N_23830,N_15537,N_18587);
or U23831 (N_23831,N_17515,N_16764);
and U23832 (N_23832,N_17917,N_18800);
and U23833 (N_23833,N_17226,N_16487);
and U23834 (N_23834,N_16081,N_19470);
nand U23835 (N_23835,N_16361,N_16261);
or U23836 (N_23836,N_19795,N_19908);
or U23837 (N_23837,N_15246,N_19508);
and U23838 (N_23838,N_16308,N_17918);
and U23839 (N_23839,N_19120,N_17654);
nor U23840 (N_23840,N_17036,N_17467);
nand U23841 (N_23841,N_17782,N_16432);
or U23842 (N_23842,N_19502,N_15986);
nor U23843 (N_23843,N_17868,N_17755);
nand U23844 (N_23844,N_19394,N_18250);
nor U23845 (N_23845,N_19282,N_15732);
nand U23846 (N_23846,N_17076,N_19336);
xnor U23847 (N_23847,N_18491,N_17764);
or U23848 (N_23848,N_19122,N_19927);
or U23849 (N_23849,N_15635,N_17782);
nor U23850 (N_23850,N_18652,N_18488);
nand U23851 (N_23851,N_18333,N_18217);
and U23852 (N_23852,N_15150,N_19163);
nor U23853 (N_23853,N_18226,N_16474);
xor U23854 (N_23854,N_15322,N_18380);
nor U23855 (N_23855,N_15068,N_15803);
and U23856 (N_23856,N_19290,N_15420);
or U23857 (N_23857,N_19287,N_16665);
nor U23858 (N_23858,N_18398,N_15329);
or U23859 (N_23859,N_17307,N_15787);
nor U23860 (N_23860,N_19523,N_16611);
nor U23861 (N_23861,N_18775,N_19232);
or U23862 (N_23862,N_19738,N_18348);
nand U23863 (N_23863,N_17008,N_15643);
nand U23864 (N_23864,N_19308,N_16953);
nand U23865 (N_23865,N_17408,N_17038);
nor U23866 (N_23866,N_17252,N_19918);
nand U23867 (N_23867,N_17627,N_18399);
or U23868 (N_23868,N_16061,N_18423);
or U23869 (N_23869,N_17314,N_18274);
nor U23870 (N_23870,N_16426,N_16261);
and U23871 (N_23871,N_19406,N_15978);
nand U23872 (N_23872,N_19578,N_19850);
nor U23873 (N_23873,N_16123,N_17789);
nand U23874 (N_23874,N_16617,N_16428);
nand U23875 (N_23875,N_19902,N_18295);
and U23876 (N_23876,N_18723,N_15693);
or U23877 (N_23877,N_19900,N_19426);
or U23878 (N_23878,N_19129,N_16487);
and U23879 (N_23879,N_19297,N_18145);
or U23880 (N_23880,N_16436,N_17687);
and U23881 (N_23881,N_15303,N_15928);
and U23882 (N_23882,N_16790,N_15696);
nor U23883 (N_23883,N_16705,N_16486);
xor U23884 (N_23884,N_16323,N_17359);
and U23885 (N_23885,N_17243,N_17936);
and U23886 (N_23886,N_16838,N_19514);
or U23887 (N_23887,N_16001,N_18306);
or U23888 (N_23888,N_19283,N_18466);
nand U23889 (N_23889,N_15200,N_16956);
nand U23890 (N_23890,N_17544,N_19237);
nor U23891 (N_23891,N_17234,N_15745);
or U23892 (N_23892,N_19661,N_17557);
or U23893 (N_23893,N_17569,N_16845);
or U23894 (N_23894,N_18439,N_16084);
and U23895 (N_23895,N_15167,N_17979);
nand U23896 (N_23896,N_15185,N_18598);
nor U23897 (N_23897,N_18663,N_15075);
and U23898 (N_23898,N_15899,N_16260);
nand U23899 (N_23899,N_17938,N_18250);
and U23900 (N_23900,N_17224,N_15817);
nor U23901 (N_23901,N_19458,N_18420);
nand U23902 (N_23902,N_15996,N_17554);
and U23903 (N_23903,N_18908,N_16677);
nor U23904 (N_23904,N_18348,N_16292);
or U23905 (N_23905,N_18779,N_19287);
and U23906 (N_23906,N_15739,N_18270);
nor U23907 (N_23907,N_17000,N_17701);
and U23908 (N_23908,N_17403,N_18758);
and U23909 (N_23909,N_17105,N_16203);
nand U23910 (N_23910,N_19594,N_16622);
nor U23911 (N_23911,N_15868,N_15599);
nor U23912 (N_23912,N_15045,N_15077);
nor U23913 (N_23913,N_19248,N_15114);
nor U23914 (N_23914,N_17286,N_19208);
and U23915 (N_23915,N_18732,N_16757);
nand U23916 (N_23916,N_18418,N_16315);
nand U23917 (N_23917,N_19949,N_17038);
and U23918 (N_23918,N_19263,N_16472);
nor U23919 (N_23919,N_15292,N_18792);
or U23920 (N_23920,N_18802,N_17415);
or U23921 (N_23921,N_17592,N_15115);
nand U23922 (N_23922,N_17008,N_16513);
nand U23923 (N_23923,N_18142,N_18853);
nor U23924 (N_23924,N_17394,N_18611);
or U23925 (N_23925,N_16722,N_18718);
nor U23926 (N_23926,N_15983,N_15769);
or U23927 (N_23927,N_18674,N_16433);
nor U23928 (N_23928,N_19315,N_15755);
or U23929 (N_23929,N_18331,N_17832);
and U23930 (N_23930,N_19748,N_15115);
and U23931 (N_23931,N_19003,N_16425);
nand U23932 (N_23932,N_17192,N_15279);
nor U23933 (N_23933,N_17590,N_18702);
or U23934 (N_23934,N_18126,N_16871);
and U23935 (N_23935,N_17155,N_16610);
nor U23936 (N_23936,N_15190,N_16197);
nand U23937 (N_23937,N_16714,N_17153);
nand U23938 (N_23938,N_19171,N_18702);
or U23939 (N_23939,N_15302,N_15957);
nor U23940 (N_23940,N_15568,N_19082);
and U23941 (N_23941,N_17754,N_16237);
and U23942 (N_23942,N_17586,N_16731);
or U23943 (N_23943,N_17413,N_18521);
nand U23944 (N_23944,N_19034,N_19914);
nand U23945 (N_23945,N_15526,N_17145);
nor U23946 (N_23946,N_15796,N_15291);
nor U23947 (N_23947,N_19497,N_16539);
nor U23948 (N_23948,N_17734,N_15290);
and U23949 (N_23949,N_19350,N_15579);
or U23950 (N_23950,N_18771,N_17955);
nor U23951 (N_23951,N_17264,N_17780);
nand U23952 (N_23952,N_19281,N_18916);
and U23953 (N_23953,N_18340,N_16615);
nand U23954 (N_23954,N_18898,N_16081);
or U23955 (N_23955,N_16300,N_19156);
or U23956 (N_23956,N_17619,N_17226);
or U23957 (N_23957,N_16043,N_16897);
nand U23958 (N_23958,N_15184,N_17528);
and U23959 (N_23959,N_15779,N_17448);
nand U23960 (N_23960,N_16719,N_17923);
nand U23961 (N_23961,N_15593,N_18255);
and U23962 (N_23962,N_19775,N_15019);
nand U23963 (N_23963,N_16828,N_19015);
nand U23964 (N_23964,N_17477,N_15874);
or U23965 (N_23965,N_19927,N_18382);
or U23966 (N_23966,N_16631,N_17418);
nor U23967 (N_23967,N_17035,N_15411);
nor U23968 (N_23968,N_16898,N_16335);
xor U23969 (N_23969,N_17496,N_15531);
nor U23970 (N_23970,N_17606,N_18161);
and U23971 (N_23971,N_16401,N_19347);
nand U23972 (N_23972,N_17382,N_17287);
or U23973 (N_23973,N_19891,N_17548);
nand U23974 (N_23974,N_19217,N_17941);
nand U23975 (N_23975,N_16597,N_18641);
nor U23976 (N_23976,N_16763,N_17823);
nand U23977 (N_23977,N_17475,N_15066);
nor U23978 (N_23978,N_17728,N_17093);
or U23979 (N_23979,N_17001,N_15898);
nand U23980 (N_23980,N_15266,N_19795);
nand U23981 (N_23981,N_16614,N_15395);
nor U23982 (N_23982,N_16458,N_16944);
and U23983 (N_23983,N_16649,N_18978);
nand U23984 (N_23984,N_15039,N_17222);
or U23985 (N_23985,N_18649,N_18636);
nand U23986 (N_23986,N_15582,N_18219);
and U23987 (N_23987,N_16436,N_17568);
nand U23988 (N_23988,N_19957,N_18190);
nor U23989 (N_23989,N_19431,N_16882);
or U23990 (N_23990,N_19564,N_17288);
nor U23991 (N_23991,N_18895,N_19324);
or U23992 (N_23992,N_17933,N_15994);
nor U23993 (N_23993,N_17245,N_16167);
and U23994 (N_23994,N_15578,N_17825);
and U23995 (N_23995,N_16775,N_16089);
nand U23996 (N_23996,N_15956,N_15773);
nor U23997 (N_23997,N_17511,N_18000);
and U23998 (N_23998,N_19479,N_17245);
nor U23999 (N_23999,N_18863,N_19957);
nor U24000 (N_24000,N_18536,N_16812);
nor U24001 (N_24001,N_18505,N_16402);
nand U24002 (N_24002,N_18812,N_15742);
or U24003 (N_24003,N_18660,N_15416);
nor U24004 (N_24004,N_16630,N_17796);
and U24005 (N_24005,N_16358,N_19043);
nor U24006 (N_24006,N_15375,N_19804);
or U24007 (N_24007,N_18141,N_16368);
nor U24008 (N_24008,N_17728,N_17531);
nand U24009 (N_24009,N_19255,N_18739);
nand U24010 (N_24010,N_17384,N_16124);
and U24011 (N_24011,N_16789,N_17619);
nor U24012 (N_24012,N_19609,N_18770);
nand U24013 (N_24013,N_19542,N_15784);
nor U24014 (N_24014,N_18084,N_15450);
and U24015 (N_24015,N_19265,N_15111);
and U24016 (N_24016,N_19535,N_17686);
nand U24017 (N_24017,N_17770,N_16744);
nor U24018 (N_24018,N_19502,N_16851);
or U24019 (N_24019,N_17857,N_15299);
nand U24020 (N_24020,N_17902,N_19628);
and U24021 (N_24021,N_19894,N_15944);
and U24022 (N_24022,N_15357,N_17887);
nand U24023 (N_24023,N_16187,N_17613);
or U24024 (N_24024,N_16924,N_16490);
or U24025 (N_24025,N_18982,N_18032);
and U24026 (N_24026,N_15889,N_18104);
nor U24027 (N_24027,N_16047,N_17953);
nand U24028 (N_24028,N_17741,N_15364);
or U24029 (N_24029,N_17561,N_19439);
and U24030 (N_24030,N_15265,N_16680);
nor U24031 (N_24031,N_18279,N_15859);
and U24032 (N_24032,N_16820,N_18149);
nor U24033 (N_24033,N_15398,N_19965);
and U24034 (N_24034,N_15588,N_16838);
nor U24035 (N_24035,N_15059,N_18203);
nand U24036 (N_24036,N_16312,N_15363);
nand U24037 (N_24037,N_15997,N_16061);
nand U24038 (N_24038,N_15257,N_19178);
or U24039 (N_24039,N_17472,N_18404);
and U24040 (N_24040,N_17779,N_19658);
and U24041 (N_24041,N_15745,N_17836);
and U24042 (N_24042,N_16229,N_15292);
xor U24043 (N_24043,N_16297,N_16347);
nor U24044 (N_24044,N_19698,N_19491);
or U24045 (N_24045,N_17549,N_17529);
or U24046 (N_24046,N_15497,N_15552);
and U24047 (N_24047,N_15790,N_16187);
nor U24048 (N_24048,N_19410,N_15540);
nor U24049 (N_24049,N_18419,N_15268);
and U24050 (N_24050,N_18218,N_17695);
nor U24051 (N_24051,N_19225,N_16232);
nand U24052 (N_24052,N_17602,N_18815);
and U24053 (N_24053,N_16412,N_17593);
and U24054 (N_24054,N_19011,N_18700);
or U24055 (N_24055,N_16923,N_17049);
or U24056 (N_24056,N_18540,N_17219);
nand U24057 (N_24057,N_19310,N_18708);
and U24058 (N_24058,N_18804,N_18640);
and U24059 (N_24059,N_19519,N_18212);
or U24060 (N_24060,N_16729,N_18225);
nor U24061 (N_24061,N_17593,N_15574);
or U24062 (N_24062,N_19211,N_15677);
nand U24063 (N_24063,N_17689,N_19548);
nand U24064 (N_24064,N_19360,N_17358);
nand U24065 (N_24065,N_17745,N_17341);
nor U24066 (N_24066,N_16898,N_18895);
nor U24067 (N_24067,N_16760,N_17363);
and U24068 (N_24068,N_18526,N_15101);
or U24069 (N_24069,N_17071,N_19926);
nand U24070 (N_24070,N_15940,N_18400);
or U24071 (N_24071,N_19242,N_17419);
nand U24072 (N_24072,N_15674,N_15056);
nor U24073 (N_24073,N_17046,N_18321);
or U24074 (N_24074,N_16934,N_15497);
and U24075 (N_24075,N_17647,N_15001);
and U24076 (N_24076,N_18258,N_17626);
nor U24077 (N_24077,N_15622,N_18647);
and U24078 (N_24078,N_18367,N_15694);
and U24079 (N_24079,N_19068,N_19434);
and U24080 (N_24080,N_17269,N_17287);
nor U24081 (N_24081,N_18601,N_18456);
nor U24082 (N_24082,N_15921,N_19187);
nand U24083 (N_24083,N_15775,N_18285);
nand U24084 (N_24084,N_17411,N_18905);
nor U24085 (N_24085,N_18857,N_15663);
nor U24086 (N_24086,N_19998,N_19382);
nand U24087 (N_24087,N_19126,N_19581);
nand U24088 (N_24088,N_17663,N_19094);
or U24089 (N_24089,N_19945,N_16864);
nand U24090 (N_24090,N_15115,N_18686);
and U24091 (N_24091,N_17891,N_15769);
nor U24092 (N_24092,N_18923,N_18176);
and U24093 (N_24093,N_19087,N_15464);
and U24094 (N_24094,N_17741,N_16962);
nor U24095 (N_24095,N_19727,N_18560);
and U24096 (N_24096,N_19759,N_17533);
and U24097 (N_24097,N_16619,N_17762);
or U24098 (N_24098,N_16595,N_17451);
nor U24099 (N_24099,N_19140,N_18243);
or U24100 (N_24100,N_16890,N_15996);
and U24101 (N_24101,N_15684,N_17160);
nor U24102 (N_24102,N_19954,N_15822);
and U24103 (N_24103,N_15545,N_18194);
or U24104 (N_24104,N_16401,N_17312);
and U24105 (N_24105,N_19953,N_18561);
and U24106 (N_24106,N_15595,N_17709);
nor U24107 (N_24107,N_17971,N_15938);
nor U24108 (N_24108,N_15407,N_16563);
and U24109 (N_24109,N_15593,N_15223);
and U24110 (N_24110,N_18138,N_16152);
nor U24111 (N_24111,N_18338,N_19244);
and U24112 (N_24112,N_19333,N_19790);
nor U24113 (N_24113,N_18931,N_15425);
xor U24114 (N_24114,N_17387,N_15370);
and U24115 (N_24115,N_19640,N_19096);
or U24116 (N_24116,N_19696,N_19559);
nand U24117 (N_24117,N_15665,N_18441);
nand U24118 (N_24118,N_18411,N_19327);
nand U24119 (N_24119,N_17727,N_18611);
and U24120 (N_24120,N_18897,N_16628);
or U24121 (N_24121,N_17024,N_19265);
or U24122 (N_24122,N_19708,N_16681);
nor U24123 (N_24123,N_19305,N_17937);
or U24124 (N_24124,N_15010,N_15073);
nand U24125 (N_24125,N_17418,N_16374);
nor U24126 (N_24126,N_16027,N_19822);
or U24127 (N_24127,N_19510,N_16662);
nor U24128 (N_24128,N_18449,N_16551);
or U24129 (N_24129,N_16085,N_18715);
and U24130 (N_24130,N_18633,N_15166);
nand U24131 (N_24131,N_16998,N_16948);
nand U24132 (N_24132,N_19323,N_16382);
nor U24133 (N_24133,N_15175,N_15305);
nor U24134 (N_24134,N_15456,N_17131);
or U24135 (N_24135,N_17043,N_15939);
and U24136 (N_24136,N_19072,N_15601);
nand U24137 (N_24137,N_15534,N_17445);
nor U24138 (N_24138,N_18589,N_18431);
nor U24139 (N_24139,N_16172,N_19542);
nor U24140 (N_24140,N_19296,N_19964);
nor U24141 (N_24141,N_18700,N_18914);
nor U24142 (N_24142,N_18188,N_17096);
or U24143 (N_24143,N_18811,N_18394);
and U24144 (N_24144,N_17314,N_15506);
nor U24145 (N_24145,N_16977,N_19520);
and U24146 (N_24146,N_16305,N_16934);
nand U24147 (N_24147,N_19065,N_16627);
or U24148 (N_24148,N_16188,N_16593);
nor U24149 (N_24149,N_17097,N_18691);
and U24150 (N_24150,N_19435,N_16814);
nor U24151 (N_24151,N_19932,N_15216);
or U24152 (N_24152,N_18133,N_19800);
nand U24153 (N_24153,N_17221,N_16235);
or U24154 (N_24154,N_17165,N_19212);
nor U24155 (N_24155,N_18509,N_18135);
nor U24156 (N_24156,N_16595,N_18705);
and U24157 (N_24157,N_16604,N_17930);
nor U24158 (N_24158,N_16017,N_17981);
and U24159 (N_24159,N_16392,N_18670);
and U24160 (N_24160,N_19770,N_15753);
or U24161 (N_24161,N_19656,N_17321);
nand U24162 (N_24162,N_18199,N_16190);
nand U24163 (N_24163,N_16614,N_15279);
and U24164 (N_24164,N_18645,N_15444);
and U24165 (N_24165,N_18372,N_16000);
nand U24166 (N_24166,N_16877,N_15309);
and U24167 (N_24167,N_15421,N_19508);
nand U24168 (N_24168,N_18617,N_18783);
or U24169 (N_24169,N_19461,N_16383);
nand U24170 (N_24170,N_15633,N_18979);
nand U24171 (N_24171,N_17040,N_15690);
and U24172 (N_24172,N_18319,N_16247);
or U24173 (N_24173,N_17533,N_19585);
and U24174 (N_24174,N_19656,N_17781);
nand U24175 (N_24175,N_15413,N_19478);
nand U24176 (N_24176,N_18299,N_19843);
or U24177 (N_24177,N_17302,N_19937);
nor U24178 (N_24178,N_17787,N_18405);
nand U24179 (N_24179,N_19978,N_17331);
and U24180 (N_24180,N_16553,N_18457);
nand U24181 (N_24181,N_16361,N_19606);
or U24182 (N_24182,N_18224,N_15599);
nor U24183 (N_24183,N_15790,N_17056);
nor U24184 (N_24184,N_19499,N_19261);
nor U24185 (N_24185,N_17671,N_16505);
or U24186 (N_24186,N_18630,N_16992);
nand U24187 (N_24187,N_16203,N_15839);
and U24188 (N_24188,N_17628,N_16461);
nor U24189 (N_24189,N_16434,N_18458);
nand U24190 (N_24190,N_16949,N_17302);
nand U24191 (N_24191,N_16644,N_17033);
nand U24192 (N_24192,N_19283,N_15283);
and U24193 (N_24193,N_19002,N_17215);
and U24194 (N_24194,N_15621,N_15410);
and U24195 (N_24195,N_17422,N_19735);
nor U24196 (N_24196,N_19851,N_18334);
or U24197 (N_24197,N_19781,N_16663);
xor U24198 (N_24198,N_17913,N_19972);
nor U24199 (N_24199,N_16365,N_16473);
and U24200 (N_24200,N_17482,N_17964);
and U24201 (N_24201,N_17127,N_19223);
nand U24202 (N_24202,N_17161,N_17390);
nor U24203 (N_24203,N_17161,N_19518);
and U24204 (N_24204,N_19667,N_16498);
nand U24205 (N_24205,N_16506,N_18703);
nor U24206 (N_24206,N_19404,N_17421);
xor U24207 (N_24207,N_15841,N_19972);
and U24208 (N_24208,N_16424,N_15796);
nand U24209 (N_24209,N_17472,N_16628);
nand U24210 (N_24210,N_16230,N_19243);
or U24211 (N_24211,N_18248,N_19226);
or U24212 (N_24212,N_16767,N_17554);
nand U24213 (N_24213,N_19150,N_17513);
nor U24214 (N_24214,N_16277,N_19972);
nand U24215 (N_24215,N_16442,N_15254);
nand U24216 (N_24216,N_18836,N_19727);
nor U24217 (N_24217,N_18171,N_15247);
nor U24218 (N_24218,N_16273,N_16443);
nor U24219 (N_24219,N_16307,N_16642);
and U24220 (N_24220,N_18415,N_18508);
nor U24221 (N_24221,N_17398,N_15971);
nor U24222 (N_24222,N_19127,N_17499);
nand U24223 (N_24223,N_15128,N_19083);
or U24224 (N_24224,N_19001,N_19757);
nand U24225 (N_24225,N_15647,N_18897);
nor U24226 (N_24226,N_17657,N_19377);
nand U24227 (N_24227,N_17334,N_15476);
nor U24228 (N_24228,N_19445,N_18834);
or U24229 (N_24229,N_15264,N_15665);
nand U24230 (N_24230,N_17744,N_17786);
or U24231 (N_24231,N_16438,N_15446);
nor U24232 (N_24232,N_16563,N_19915);
and U24233 (N_24233,N_18047,N_17543);
nand U24234 (N_24234,N_19505,N_19360);
nand U24235 (N_24235,N_15131,N_18557);
nor U24236 (N_24236,N_18100,N_15958);
or U24237 (N_24237,N_16332,N_17641);
and U24238 (N_24238,N_18044,N_17093);
nor U24239 (N_24239,N_17783,N_15948);
nor U24240 (N_24240,N_16025,N_15010);
nand U24241 (N_24241,N_16715,N_15730);
nand U24242 (N_24242,N_19434,N_17056);
nor U24243 (N_24243,N_16240,N_18904);
or U24244 (N_24244,N_18502,N_19660);
or U24245 (N_24245,N_16528,N_16865);
xnor U24246 (N_24246,N_15609,N_16818);
nand U24247 (N_24247,N_17235,N_16204);
nor U24248 (N_24248,N_17478,N_17819);
and U24249 (N_24249,N_19487,N_18812);
and U24250 (N_24250,N_19173,N_17812);
and U24251 (N_24251,N_19088,N_15112);
nand U24252 (N_24252,N_15157,N_15117);
or U24253 (N_24253,N_15313,N_19771);
nor U24254 (N_24254,N_19879,N_17848);
or U24255 (N_24255,N_19418,N_19641);
nand U24256 (N_24256,N_19471,N_18409);
nor U24257 (N_24257,N_15463,N_17407);
or U24258 (N_24258,N_19704,N_17480);
and U24259 (N_24259,N_18847,N_18559);
nor U24260 (N_24260,N_15007,N_17353);
and U24261 (N_24261,N_18008,N_17121);
nand U24262 (N_24262,N_15393,N_16050);
or U24263 (N_24263,N_18887,N_19484);
nand U24264 (N_24264,N_15299,N_17212);
or U24265 (N_24265,N_16495,N_16496);
nor U24266 (N_24266,N_16375,N_18960);
nor U24267 (N_24267,N_18805,N_16304);
and U24268 (N_24268,N_17248,N_17748);
and U24269 (N_24269,N_16416,N_18853);
nand U24270 (N_24270,N_19183,N_15515);
nand U24271 (N_24271,N_16986,N_16799);
nor U24272 (N_24272,N_15520,N_18329);
nor U24273 (N_24273,N_16124,N_17545);
nor U24274 (N_24274,N_16366,N_17434);
nor U24275 (N_24275,N_17191,N_18896);
nand U24276 (N_24276,N_17169,N_19309);
nand U24277 (N_24277,N_15784,N_16433);
and U24278 (N_24278,N_15839,N_17773);
nand U24279 (N_24279,N_15190,N_18464);
nor U24280 (N_24280,N_18205,N_15306);
nor U24281 (N_24281,N_16071,N_17426);
or U24282 (N_24282,N_19017,N_17925);
nand U24283 (N_24283,N_19098,N_15407);
and U24284 (N_24284,N_18398,N_15046);
xor U24285 (N_24285,N_16443,N_19714);
nor U24286 (N_24286,N_16365,N_15687);
and U24287 (N_24287,N_17563,N_17250);
or U24288 (N_24288,N_15603,N_18715);
nor U24289 (N_24289,N_18654,N_15968);
or U24290 (N_24290,N_18732,N_17148);
or U24291 (N_24291,N_16532,N_19954);
nand U24292 (N_24292,N_17371,N_19403);
and U24293 (N_24293,N_15518,N_17148);
nand U24294 (N_24294,N_18660,N_18224);
and U24295 (N_24295,N_16441,N_16719);
nor U24296 (N_24296,N_16390,N_15261);
and U24297 (N_24297,N_19729,N_15822);
nand U24298 (N_24298,N_16740,N_16925);
nor U24299 (N_24299,N_18700,N_17513);
nand U24300 (N_24300,N_15387,N_18478);
nor U24301 (N_24301,N_17037,N_19298);
or U24302 (N_24302,N_16412,N_17745);
and U24303 (N_24303,N_18044,N_15377);
or U24304 (N_24304,N_17739,N_16038);
and U24305 (N_24305,N_16241,N_15896);
nand U24306 (N_24306,N_19720,N_19794);
nand U24307 (N_24307,N_18989,N_17202);
or U24308 (N_24308,N_19308,N_19530);
nand U24309 (N_24309,N_17673,N_16090);
nor U24310 (N_24310,N_16163,N_18058);
nand U24311 (N_24311,N_15396,N_18938);
nand U24312 (N_24312,N_19565,N_16541);
and U24313 (N_24313,N_18791,N_19374);
nand U24314 (N_24314,N_16287,N_19793);
nand U24315 (N_24315,N_17881,N_15584);
nand U24316 (N_24316,N_18886,N_19144);
and U24317 (N_24317,N_15500,N_17205);
nor U24318 (N_24318,N_18903,N_16790);
and U24319 (N_24319,N_19133,N_18279);
nand U24320 (N_24320,N_17930,N_18400);
and U24321 (N_24321,N_18674,N_18419);
or U24322 (N_24322,N_18700,N_17486);
nor U24323 (N_24323,N_18594,N_19567);
nor U24324 (N_24324,N_17020,N_15569);
and U24325 (N_24325,N_16179,N_18572);
nor U24326 (N_24326,N_16524,N_16339);
nand U24327 (N_24327,N_15406,N_17291);
nand U24328 (N_24328,N_18150,N_18292);
and U24329 (N_24329,N_18017,N_15997);
and U24330 (N_24330,N_19237,N_18285);
and U24331 (N_24331,N_17358,N_18281);
nor U24332 (N_24332,N_18356,N_18329);
nor U24333 (N_24333,N_17738,N_17558);
and U24334 (N_24334,N_16864,N_19377);
nor U24335 (N_24335,N_16271,N_19626);
nand U24336 (N_24336,N_15657,N_19310);
and U24337 (N_24337,N_18005,N_18292);
nand U24338 (N_24338,N_15465,N_18473);
nand U24339 (N_24339,N_18937,N_17665);
and U24340 (N_24340,N_19201,N_17499);
nor U24341 (N_24341,N_15944,N_16753);
and U24342 (N_24342,N_18116,N_15084);
nor U24343 (N_24343,N_17874,N_15958);
nand U24344 (N_24344,N_16597,N_17318);
and U24345 (N_24345,N_16227,N_15753);
and U24346 (N_24346,N_18766,N_18643);
and U24347 (N_24347,N_16452,N_17535);
nand U24348 (N_24348,N_17270,N_18824);
nand U24349 (N_24349,N_16543,N_16557);
nand U24350 (N_24350,N_15439,N_15393);
or U24351 (N_24351,N_17042,N_15043);
nor U24352 (N_24352,N_19644,N_18211);
or U24353 (N_24353,N_19665,N_19330);
nor U24354 (N_24354,N_15831,N_16605);
nand U24355 (N_24355,N_19216,N_16577);
and U24356 (N_24356,N_15752,N_18788);
and U24357 (N_24357,N_15553,N_15644);
and U24358 (N_24358,N_19294,N_17278);
nor U24359 (N_24359,N_16772,N_19755);
and U24360 (N_24360,N_17673,N_19385);
or U24361 (N_24361,N_17339,N_15543);
nor U24362 (N_24362,N_17461,N_16173);
nand U24363 (N_24363,N_19037,N_16852);
nor U24364 (N_24364,N_17024,N_19620);
or U24365 (N_24365,N_15302,N_19218);
or U24366 (N_24366,N_18668,N_16452);
nor U24367 (N_24367,N_19055,N_16126);
or U24368 (N_24368,N_18073,N_18039);
nor U24369 (N_24369,N_16024,N_16861);
and U24370 (N_24370,N_18150,N_16181);
and U24371 (N_24371,N_17492,N_18766);
nand U24372 (N_24372,N_16054,N_18837);
and U24373 (N_24373,N_18416,N_16171);
nor U24374 (N_24374,N_18444,N_19088);
nor U24375 (N_24375,N_16551,N_18878);
or U24376 (N_24376,N_17668,N_19403);
xnor U24377 (N_24377,N_17446,N_18981);
nor U24378 (N_24378,N_17827,N_16550);
and U24379 (N_24379,N_19546,N_16363);
nand U24380 (N_24380,N_16411,N_15000);
and U24381 (N_24381,N_15827,N_16714);
or U24382 (N_24382,N_16143,N_18505);
nand U24383 (N_24383,N_19992,N_16826);
or U24384 (N_24384,N_17439,N_15103);
nand U24385 (N_24385,N_18610,N_16830);
or U24386 (N_24386,N_19352,N_19624);
nor U24387 (N_24387,N_17216,N_16692);
and U24388 (N_24388,N_17808,N_17262);
or U24389 (N_24389,N_15075,N_15621);
nor U24390 (N_24390,N_19631,N_16109);
or U24391 (N_24391,N_15383,N_18473);
nand U24392 (N_24392,N_16624,N_18017);
nand U24393 (N_24393,N_15124,N_17516);
and U24394 (N_24394,N_19366,N_15083);
and U24395 (N_24395,N_18832,N_16938);
nor U24396 (N_24396,N_17809,N_17098);
or U24397 (N_24397,N_18900,N_17903);
nor U24398 (N_24398,N_17644,N_16436);
nor U24399 (N_24399,N_19287,N_19308);
or U24400 (N_24400,N_16908,N_18650);
nand U24401 (N_24401,N_19218,N_19314);
nand U24402 (N_24402,N_17035,N_15322);
nor U24403 (N_24403,N_19622,N_15064);
nand U24404 (N_24404,N_17411,N_17949);
and U24405 (N_24405,N_17482,N_17795);
nand U24406 (N_24406,N_19999,N_19774);
nand U24407 (N_24407,N_18469,N_18713);
nor U24408 (N_24408,N_16430,N_19426);
or U24409 (N_24409,N_15719,N_17141);
or U24410 (N_24410,N_18380,N_15221);
and U24411 (N_24411,N_17064,N_16099);
nand U24412 (N_24412,N_16668,N_19924);
or U24413 (N_24413,N_18110,N_17162);
nor U24414 (N_24414,N_18610,N_16966);
or U24415 (N_24415,N_18241,N_19603);
and U24416 (N_24416,N_19968,N_15335);
and U24417 (N_24417,N_15865,N_16356);
nor U24418 (N_24418,N_16348,N_16178);
and U24419 (N_24419,N_19958,N_17566);
and U24420 (N_24420,N_18050,N_15218);
or U24421 (N_24421,N_15572,N_16064);
nand U24422 (N_24422,N_18998,N_17252);
nand U24423 (N_24423,N_16003,N_17034);
nand U24424 (N_24424,N_18146,N_15217);
xnor U24425 (N_24425,N_18714,N_18871);
xor U24426 (N_24426,N_19134,N_15873);
or U24427 (N_24427,N_16609,N_15476);
nand U24428 (N_24428,N_17043,N_16192);
nor U24429 (N_24429,N_17360,N_17565);
nand U24430 (N_24430,N_16913,N_17707);
nor U24431 (N_24431,N_15486,N_16099);
or U24432 (N_24432,N_17279,N_19821);
nor U24433 (N_24433,N_15241,N_18224);
nand U24434 (N_24434,N_16269,N_17574);
nand U24435 (N_24435,N_17387,N_19995);
nor U24436 (N_24436,N_17049,N_15787);
and U24437 (N_24437,N_18605,N_15762);
or U24438 (N_24438,N_16943,N_17323);
nor U24439 (N_24439,N_17537,N_17771);
or U24440 (N_24440,N_19886,N_15379);
and U24441 (N_24441,N_19506,N_16391);
or U24442 (N_24442,N_18596,N_15027);
or U24443 (N_24443,N_19647,N_15246);
and U24444 (N_24444,N_16931,N_17585);
nor U24445 (N_24445,N_17031,N_16227);
nand U24446 (N_24446,N_18529,N_19723);
and U24447 (N_24447,N_17636,N_19426);
nand U24448 (N_24448,N_16379,N_17998);
or U24449 (N_24449,N_16759,N_17690);
nor U24450 (N_24450,N_18047,N_19501);
nor U24451 (N_24451,N_19450,N_19290);
nor U24452 (N_24452,N_19354,N_15833);
nand U24453 (N_24453,N_17360,N_15891);
and U24454 (N_24454,N_19356,N_15483);
or U24455 (N_24455,N_19225,N_19131);
nor U24456 (N_24456,N_18331,N_17679);
and U24457 (N_24457,N_18011,N_19357);
and U24458 (N_24458,N_17193,N_19923);
and U24459 (N_24459,N_19934,N_15041);
nand U24460 (N_24460,N_17039,N_16703);
nor U24461 (N_24461,N_15896,N_16682);
and U24462 (N_24462,N_15743,N_18978);
or U24463 (N_24463,N_17431,N_15677);
and U24464 (N_24464,N_16610,N_15429);
nand U24465 (N_24465,N_18565,N_18414);
nor U24466 (N_24466,N_15600,N_15510);
nor U24467 (N_24467,N_15185,N_18022);
or U24468 (N_24468,N_16851,N_17818);
nand U24469 (N_24469,N_15407,N_16451);
nor U24470 (N_24470,N_17336,N_18506);
nor U24471 (N_24471,N_15856,N_15048);
nor U24472 (N_24472,N_18566,N_19326);
nor U24473 (N_24473,N_18309,N_19302);
nand U24474 (N_24474,N_17189,N_16772);
and U24475 (N_24475,N_18872,N_15037);
and U24476 (N_24476,N_18262,N_17225);
or U24477 (N_24477,N_15314,N_15152);
nand U24478 (N_24478,N_18401,N_15802);
or U24479 (N_24479,N_19495,N_15471);
and U24480 (N_24480,N_17766,N_17247);
or U24481 (N_24481,N_19689,N_15576);
nand U24482 (N_24482,N_18909,N_16489);
and U24483 (N_24483,N_17767,N_18149);
or U24484 (N_24484,N_17676,N_17657);
and U24485 (N_24485,N_19117,N_15330);
nand U24486 (N_24486,N_19481,N_16111);
nor U24487 (N_24487,N_15064,N_17940);
nand U24488 (N_24488,N_19380,N_18285);
nand U24489 (N_24489,N_15675,N_19218);
nor U24490 (N_24490,N_15245,N_15610);
nor U24491 (N_24491,N_15104,N_15376);
nor U24492 (N_24492,N_17717,N_18286);
nor U24493 (N_24493,N_18781,N_18300);
nand U24494 (N_24494,N_15452,N_19502);
nand U24495 (N_24495,N_19255,N_15957);
and U24496 (N_24496,N_15685,N_15340);
and U24497 (N_24497,N_18350,N_16025);
or U24498 (N_24498,N_18613,N_19691);
nand U24499 (N_24499,N_16657,N_16675);
and U24500 (N_24500,N_19905,N_17459);
and U24501 (N_24501,N_19236,N_15893);
nor U24502 (N_24502,N_18472,N_17701);
or U24503 (N_24503,N_18878,N_15617);
nand U24504 (N_24504,N_19881,N_19506);
nand U24505 (N_24505,N_15175,N_15519);
nand U24506 (N_24506,N_17251,N_15283);
nor U24507 (N_24507,N_19775,N_19351);
and U24508 (N_24508,N_18662,N_16021);
nor U24509 (N_24509,N_18583,N_18233);
nand U24510 (N_24510,N_18671,N_19617);
nor U24511 (N_24511,N_18242,N_16734);
and U24512 (N_24512,N_17250,N_16456);
and U24513 (N_24513,N_17295,N_15294);
nand U24514 (N_24514,N_18937,N_16847);
and U24515 (N_24515,N_18525,N_19753);
or U24516 (N_24516,N_17148,N_17236);
nor U24517 (N_24517,N_16022,N_18138);
and U24518 (N_24518,N_18512,N_19720);
or U24519 (N_24519,N_17957,N_16501);
or U24520 (N_24520,N_17430,N_17702);
nand U24521 (N_24521,N_16488,N_19022);
and U24522 (N_24522,N_16895,N_19372);
nor U24523 (N_24523,N_17958,N_16262);
nand U24524 (N_24524,N_18531,N_17015);
nand U24525 (N_24525,N_19333,N_15821);
or U24526 (N_24526,N_16485,N_16582);
nand U24527 (N_24527,N_15750,N_17394);
nand U24528 (N_24528,N_19872,N_15578);
or U24529 (N_24529,N_15841,N_19336);
nor U24530 (N_24530,N_15888,N_17775);
nor U24531 (N_24531,N_15615,N_18941);
and U24532 (N_24532,N_19396,N_16699);
or U24533 (N_24533,N_15135,N_18264);
or U24534 (N_24534,N_19286,N_19383);
nand U24535 (N_24535,N_18989,N_15994);
nor U24536 (N_24536,N_16273,N_19774);
and U24537 (N_24537,N_16073,N_16695);
or U24538 (N_24538,N_19846,N_18125);
nand U24539 (N_24539,N_18477,N_16705);
nor U24540 (N_24540,N_16728,N_17935);
and U24541 (N_24541,N_15508,N_15055);
or U24542 (N_24542,N_15721,N_18215);
nor U24543 (N_24543,N_16690,N_17884);
and U24544 (N_24544,N_16874,N_16865);
nor U24545 (N_24545,N_19009,N_16057);
nor U24546 (N_24546,N_17267,N_19143);
and U24547 (N_24547,N_19660,N_17227);
and U24548 (N_24548,N_19233,N_18156);
nor U24549 (N_24549,N_16341,N_16782);
nand U24550 (N_24550,N_15949,N_16161);
or U24551 (N_24551,N_17320,N_19202);
or U24552 (N_24552,N_15348,N_15887);
and U24553 (N_24553,N_15521,N_16830);
nand U24554 (N_24554,N_16945,N_16267);
or U24555 (N_24555,N_15084,N_16331);
or U24556 (N_24556,N_17873,N_18034);
or U24557 (N_24557,N_19404,N_16100);
or U24558 (N_24558,N_19246,N_17057);
and U24559 (N_24559,N_15224,N_17856);
nor U24560 (N_24560,N_16301,N_16694);
nor U24561 (N_24561,N_19962,N_18290);
and U24562 (N_24562,N_19039,N_15633);
and U24563 (N_24563,N_15998,N_15080);
nand U24564 (N_24564,N_15663,N_17027);
nor U24565 (N_24565,N_16892,N_15272);
nand U24566 (N_24566,N_15794,N_16878);
nand U24567 (N_24567,N_15350,N_19591);
or U24568 (N_24568,N_17059,N_15977);
or U24569 (N_24569,N_17151,N_16823);
and U24570 (N_24570,N_15342,N_17261);
and U24571 (N_24571,N_17194,N_18668);
or U24572 (N_24572,N_19251,N_16271);
nor U24573 (N_24573,N_19742,N_19861);
or U24574 (N_24574,N_17694,N_16598);
or U24575 (N_24575,N_19410,N_17314);
and U24576 (N_24576,N_19775,N_19372);
or U24577 (N_24577,N_18734,N_18261);
or U24578 (N_24578,N_18583,N_18117);
or U24579 (N_24579,N_19057,N_15141);
and U24580 (N_24580,N_15034,N_16856);
nand U24581 (N_24581,N_18356,N_16676);
and U24582 (N_24582,N_15147,N_15211);
nor U24583 (N_24583,N_17215,N_16736);
and U24584 (N_24584,N_18699,N_19616);
and U24585 (N_24585,N_15860,N_18701);
and U24586 (N_24586,N_19731,N_16492);
or U24587 (N_24587,N_18027,N_15897);
nand U24588 (N_24588,N_19104,N_19715);
or U24589 (N_24589,N_17799,N_19775);
or U24590 (N_24590,N_16865,N_19902);
nand U24591 (N_24591,N_19790,N_16120);
and U24592 (N_24592,N_16668,N_19267);
or U24593 (N_24593,N_19091,N_16874);
nor U24594 (N_24594,N_16486,N_15004);
or U24595 (N_24595,N_15021,N_17437);
and U24596 (N_24596,N_19693,N_16800);
and U24597 (N_24597,N_15668,N_19428);
and U24598 (N_24598,N_18997,N_16929);
nand U24599 (N_24599,N_16787,N_18851);
or U24600 (N_24600,N_19948,N_19197);
nor U24601 (N_24601,N_19335,N_19513);
or U24602 (N_24602,N_16819,N_18751);
xor U24603 (N_24603,N_16265,N_19607);
nand U24604 (N_24604,N_16321,N_17921);
nor U24605 (N_24605,N_17343,N_19485);
and U24606 (N_24606,N_16270,N_18594);
or U24607 (N_24607,N_17076,N_19061);
nand U24608 (N_24608,N_17944,N_18314);
nor U24609 (N_24609,N_17358,N_17308);
nand U24610 (N_24610,N_15237,N_16084);
nor U24611 (N_24611,N_16321,N_17206);
nand U24612 (N_24612,N_15529,N_19569);
and U24613 (N_24613,N_16999,N_17289);
nand U24614 (N_24614,N_18047,N_18446);
or U24615 (N_24615,N_16127,N_17487);
and U24616 (N_24616,N_18195,N_16362);
or U24617 (N_24617,N_16049,N_17574);
or U24618 (N_24618,N_16305,N_19514);
and U24619 (N_24619,N_19593,N_18450);
or U24620 (N_24620,N_19608,N_15883);
and U24621 (N_24621,N_18855,N_16910);
nor U24622 (N_24622,N_19570,N_18284);
or U24623 (N_24623,N_19729,N_15288);
and U24624 (N_24624,N_18919,N_18574);
and U24625 (N_24625,N_19530,N_15133);
or U24626 (N_24626,N_17429,N_15144);
nand U24627 (N_24627,N_16949,N_16701);
nand U24628 (N_24628,N_18703,N_16840);
or U24629 (N_24629,N_19560,N_15772);
nor U24630 (N_24630,N_17086,N_19026);
or U24631 (N_24631,N_17624,N_17601);
and U24632 (N_24632,N_19001,N_18835);
nand U24633 (N_24633,N_16005,N_17213);
or U24634 (N_24634,N_19996,N_17844);
nand U24635 (N_24635,N_15358,N_15737);
or U24636 (N_24636,N_18511,N_18376);
and U24637 (N_24637,N_15709,N_17433);
and U24638 (N_24638,N_17440,N_15586);
and U24639 (N_24639,N_15089,N_19784);
nor U24640 (N_24640,N_18400,N_16045);
or U24641 (N_24641,N_15245,N_15892);
and U24642 (N_24642,N_18919,N_15345);
nand U24643 (N_24643,N_15452,N_15273);
nor U24644 (N_24644,N_18118,N_15417);
nand U24645 (N_24645,N_16848,N_16704);
and U24646 (N_24646,N_15135,N_19561);
or U24647 (N_24647,N_16297,N_15402);
nand U24648 (N_24648,N_17131,N_19224);
xor U24649 (N_24649,N_18549,N_16851);
xnor U24650 (N_24650,N_16112,N_15380);
or U24651 (N_24651,N_17201,N_15103);
or U24652 (N_24652,N_19716,N_16946);
nand U24653 (N_24653,N_15660,N_17792);
or U24654 (N_24654,N_15851,N_16012);
nand U24655 (N_24655,N_18915,N_17526);
nand U24656 (N_24656,N_18461,N_19306);
and U24657 (N_24657,N_15860,N_15952);
or U24658 (N_24658,N_19977,N_15773);
nor U24659 (N_24659,N_16200,N_15570);
nand U24660 (N_24660,N_15526,N_16803);
and U24661 (N_24661,N_15688,N_16788);
and U24662 (N_24662,N_19196,N_18552);
and U24663 (N_24663,N_15342,N_17854);
nand U24664 (N_24664,N_15119,N_17215);
nor U24665 (N_24665,N_17793,N_18107);
nand U24666 (N_24666,N_16210,N_16407);
or U24667 (N_24667,N_19913,N_17268);
nor U24668 (N_24668,N_18256,N_17465);
nor U24669 (N_24669,N_19136,N_19531);
and U24670 (N_24670,N_15498,N_16059);
nor U24671 (N_24671,N_18664,N_16576);
and U24672 (N_24672,N_18948,N_15263);
nand U24673 (N_24673,N_16650,N_15892);
or U24674 (N_24674,N_18475,N_18762);
and U24675 (N_24675,N_15920,N_18811);
nor U24676 (N_24676,N_19221,N_19620);
nand U24677 (N_24677,N_17560,N_17024);
or U24678 (N_24678,N_17060,N_18472);
nor U24679 (N_24679,N_19795,N_17289);
nor U24680 (N_24680,N_19403,N_16499);
nand U24681 (N_24681,N_18333,N_18167);
nor U24682 (N_24682,N_15075,N_17654);
nand U24683 (N_24683,N_15026,N_16198);
nor U24684 (N_24684,N_16098,N_19428);
nor U24685 (N_24685,N_16405,N_19394);
and U24686 (N_24686,N_19806,N_16251);
nand U24687 (N_24687,N_19523,N_18715);
nor U24688 (N_24688,N_16670,N_15738);
and U24689 (N_24689,N_16694,N_17216);
and U24690 (N_24690,N_15672,N_18912);
and U24691 (N_24691,N_15741,N_17378);
xnor U24692 (N_24692,N_15895,N_19663);
nor U24693 (N_24693,N_15697,N_15444);
nand U24694 (N_24694,N_18057,N_16868);
nand U24695 (N_24695,N_16495,N_16000);
nor U24696 (N_24696,N_19117,N_18304);
and U24697 (N_24697,N_16223,N_18938);
nor U24698 (N_24698,N_15240,N_15988);
and U24699 (N_24699,N_15131,N_17905);
or U24700 (N_24700,N_17827,N_18788);
nand U24701 (N_24701,N_15088,N_15434);
and U24702 (N_24702,N_16602,N_17663);
or U24703 (N_24703,N_17907,N_18071);
or U24704 (N_24704,N_15660,N_19156);
and U24705 (N_24705,N_17040,N_15848);
nor U24706 (N_24706,N_18131,N_16817);
or U24707 (N_24707,N_17158,N_15369);
nor U24708 (N_24708,N_15924,N_19287);
nand U24709 (N_24709,N_16171,N_16225);
or U24710 (N_24710,N_16607,N_15920);
nand U24711 (N_24711,N_19836,N_18939);
nand U24712 (N_24712,N_16061,N_19508);
nand U24713 (N_24713,N_19553,N_19110);
nor U24714 (N_24714,N_17042,N_15779);
or U24715 (N_24715,N_16928,N_18574);
and U24716 (N_24716,N_16571,N_16529);
and U24717 (N_24717,N_19427,N_15658);
nand U24718 (N_24718,N_15594,N_15347);
and U24719 (N_24719,N_15571,N_17276);
or U24720 (N_24720,N_17155,N_17996);
or U24721 (N_24721,N_17604,N_16858);
and U24722 (N_24722,N_15888,N_16799);
and U24723 (N_24723,N_19099,N_19213);
nor U24724 (N_24724,N_16765,N_16476);
nand U24725 (N_24725,N_19257,N_18721);
nor U24726 (N_24726,N_17392,N_15001);
or U24727 (N_24727,N_15606,N_16255);
or U24728 (N_24728,N_17691,N_18660);
nor U24729 (N_24729,N_16333,N_17632);
nor U24730 (N_24730,N_18673,N_17329);
or U24731 (N_24731,N_18161,N_18942);
and U24732 (N_24732,N_18346,N_19920);
nand U24733 (N_24733,N_19154,N_18457);
or U24734 (N_24734,N_18681,N_16728);
or U24735 (N_24735,N_19716,N_18483);
nor U24736 (N_24736,N_19786,N_16578);
or U24737 (N_24737,N_19841,N_17761);
and U24738 (N_24738,N_19137,N_17361);
or U24739 (N_24739,N_19467,N_16304);
and U24740 (N_24740,N_17821,N_17048);
nand U24741 (N_24741,N_16796,N_19489);
nand U24742 (N_24742,N_17096,N_15325);
nor U24743 (N_24743,N_15600,N_15591);
nor U24744 (N_24744,N_16880,N_16215);
nor U24745 (N_24745,N_18083,N_19334);
or U24746 (N_24746,N_15456,N_16580);
nand U24747 (N_24747,N_19079,N_19393);
or U24748 (N_24748,N_17303,N_18640);
and U24749 (N_24749,N_17519,N_15623);
nand U24750 (N_24750,N_19041,N_17647);
xor U24751 (N_24751,N_18122,N_17581);
nor U24752 (N_24752,N_17307,N_18356);
or U24753 (N_24753,N_18719,N_17699);
nor U24754 (N_24754,N_16418,N_15345);
and U24755 (N_24755,N_17254,N_17205);
nand U24756 (N_24756,N_15233,N_18650);
nor U24757 (N_24757,N_15493,N_15660);
or U24758 (N_24758,N_15189,N_16014);
nand U24759 (N_24759,N_17401,N_18152);
nand U24760 (N_24760,N_17641,N_15267);
or U24761 (N_24761,N_16811,N_16557);
nor U24762 (N_24762,N_18479,N_17283);
nor U24763 (N_24763,N_16629,N_18378);
nand U24764 (N_24764,N_18542,N_16791);
and U24765 (N_24765,N_18520,N_19649);
nand U24766 (N_24766,N_15673,N_19783);
xnor U24767 (N_24767,N_19119,N_15343);
and U24768 (N_24768,N_18582,N_18431);
and U24769 (N_24769,N_19965,N_17608);
nand U24770 (N_24770,N_18058,N_16518);
nand U24771 (N_24771,N_17057,N_15941);
nor U24772 (N_24772,N_19767,N_19203);
and U24773 (N_24773,N_19213,N_16423);
and U24774 (N_24774,N_15204,N_19472);
or U24775 (N_24775,N_16647,N_19506);
nor U24776 (N_24776,N_15133,N_18736);
nor U24777 (N_24777,N_19772,N_18057);
and U24778 (N_24778,N_15843,N_16264);
and U24779 (N_24779,N_18116,N_16590);
nand U24780 (N_24780,N_16062,N_17015);
or U24781 (N_24781,N_19738,N_17837);
and U24782 (N_24782,N_15442,N_19827);
or U24783 (N_24783,N_17693,N_19793);
and U24784 (N_24784,N_16352,N_15007);
nand U24785 (N_24785,N_15638,N_19739);
nand U24786 (N_24786,N_18361,N_16323);
nand U24787 (N_24787,N_18181,N_16964);
or U24788 (N_24788,N_17623,N_17954);
and U24789 (N_24789,N_16087,N_15899);
or U24790 (N_24790,N_15071,N_15599);
nand U24791 (N_24791,N_19360,N_15316);
nor U24792 (N_24792,N_18251,N_18435);
nand U24793 (N_24793,N_15456,N_18126);
and U24794 (N_24794,N_17129,N_16737);
or U24795 (N_24795,N_17376,N_19668);
nand U24796 (N_24796,N_17153,N_17764);
or U24797 (N_24797,N_18049,N_18669);
and U24798 (N_24798,N_16196,N_16078);
and U24799 (N_24799,N_19456,N_19335);
nor U24800 (N_24800,N_19065,N_15005);
nor U24801 (N_24801,N_18364,N_17007);
or U24802 (N_24802,N_18198,N_16195);
or U24803 (N_24803,N_16863,N_18184);
nor U24804 (N_24804,N_19195,N_18601);
nand U24805 (N_24805,N_17646,N_18528);
nor U24806 (N_24806,N_16570,N_16611);
nor U24807 (N_24807,N_15386,N_16194);
or U24808 (N_24808,N_18520,N_19889);
nor U24809 (N_24809,N_19195,N_16218);
nand U24810 (N_24810,N_18188,N_15644);
nor U24811 (N_24811,N_17863,N_15469);
or U24812 (N_24812,N_18749,N_16217);
and U24813 (N_24813,N_17134,N_18270);
and U24814 (N_24814,N_16731,N_18901);
or U24815 (N_24815,N_18433,N_18903);
nor U24816 (N_24816,N_19371,N_18833);
nand U24817 (N_24817,N_15971,N_19764);
nor U24818 (N_24818,N_15044,N_19418);
or U24819 (N_24819,N_16806,N_17677);
or U24820 (N_24820,N_17756,N_17443);
nor U24821 (N_24821,N_16199,N_16123);
nand U24822 (N_24822,N_15858,N_19757);
nand U24823 (N_24823,N_19638,N_17476);
and U24824 (N_24824,N_17121,N_19397);
or U24825 (N_24825,N_15979,N_19355);
nor U24826 (N_24826,N_16833,N_16902);
nor U24827 (N_24827,N_15548,N_19708);
nor U24828 (N_24828,N_16579,N_18164);
or U24829 (N_24829,N_19231,N_19357);
nand U24830 (N_24830,N_18250,N_16930);
or U24831 (N_24831,N_16487,N_17569);
nor U24832 (N_24832,N_15062,N_18101);
nand U24833 (N_24833,N_16478,N_15130);
and U24834 (N_24834,N_19127,N_19370);
and U24835 (N_24835,N_19970,N_17270);
nor U24836 (N_24836,N_15534,N_15096);
and U24837 (N_24837,N_15802,N_19198);
and U24838 (N_24838,N_19778,N_15781);
nor U24839 (N_24839,N_18324,N_18169);
and U24840 (N_24840,N_16182,N_15205);
or U24841 (N_24841,N_16621,N_15485);
nor U24842 (N_24842,N_19256,N_18300);
nor U24843 (N_24843,N_18639,N_18967);
nand U24844 (N_24844,N_18203,N_17382);
and U24845 (N_24845,N_15550,N_19761);
or U24846 (N_24846,N_19815,N_17998);
or U24847 (N_24847,N_19112,N_16942);
nor U24848 (N_24848,N_17429,N_15425);
or U24849 (N_24849,N_17655,N_16594);
nand U24850 (N_24850,N_15989,N_19824);
xor U24851 (N_24851,N_16521,N_18435);
nor U24852 (N_24852,N_19329,N_15649);
or U24853 (N_24853,N_15078,N_19780);
or U24854 (N_24854,N_15329,N_15863);
nor U24855 (N_24855,N_19944,N_17179);
or U24856 (N_24856,N_19371,N_17506);
or U24857 (N_24857,N_17135,N_18593);
or U24858 (N_24858,N_18172,N_16765);
nand U24859 (N_24859,N_15184,N_19400);
nor U24860 (N_24860,N_18236,N_19214);
or U24861 (N_24861,N_17880,N_17311);
and U24862 (N_24862,N_16145,N_17213);
nor U24863 (N_24863,N_15069,N_17427);
and U24864 (N_24864,N_19269,N_16617);
or U24865 (N_24865,N_16276,N_19695);
nor U24866 (N_24866,N_16781,N_18846);
nand U24867 (N_24867,N_17401,N_19625);
and U24868 (N_24868,N_19148,N_15712);
nor U24869 (N_24869,N_19550,N_16007);
nor U24870 (N_24870,N_16704,N_16070);
nand U24871 (N_24871,N_17531,N_15275);
and U24872 (N_24872,N_15584,N_15847);
or U24873 (N_24873,N_18127,N_15914);
and U24874 (N_24874,N_15261,N_16478);
nand U24875 (N_24875,N_18419,N_17911);
nor U24876 (N_24876,N_18255,N_16112);
nor U24877 (N_24877,N_17369,N_19957);
nor U24878 (N_24878,N_19851,N_18633);
or U24879 (N_24879,N_18713,N_19643);
nor U24880 (N_24880,N_19112,N_15823);
or U24881 (N_24881,N_18020,N_16405);
nand U24882 (N_24882,N_17439,N_19030);
or U24883 (N_24883,N_19565,N_15008);
nand U24884 (N_24884,N_18397,N_19336);
and U24885 (N_24885,N_15313,N_15855);
or U24886 (N_24886,N_16959,N_17097);
nand U24887 (N_24887,N_19427,N_17905);
and U24888 (N_24888,N_17604,N_18099);
and U24889 (N_24889,N_17292,N_18565);
nand U24890 (N_24890,N_15178,N_17471);
nand U24891 (N_24891,N_19513,N_16709);
and U24892 (N_24892,N_18873,N_16767);
and U24893 (N_24893,N_19679,N_16135);
xor U24894 (N_24894,N_15570,N_18803);
nand U24895 (N_24895,N_18140,N_17631);
and U24896 (N_24896,N_15924,N_17440);
nor U24897 (N_24897,N_18534,N_16531);
nor U24898 (N_24898,N_19790,N_19484);
nand U24899 (N_24899,N_17656,N_18757);
or U24900 (N_24900,N_18580,N_18636);
or U24901 (N_24901,N_18488,N_16226);
nor U24902 (N_24902,N_18916,N_16037);
and U24903 (N_24903,N_17274,N_19352);
or U24904 (N_24904,N_16339,N_15463);
and U24905 (N_24905,N_16548,N_15495);
nor U24906 (N_24906,N_16169,N_17242);
and U24907 (N_24907,N_18325,N_16197);
nor U24908 (N_24908,N_17433,N_15529);
nor U24909 (N_24909,N_18233,N_16357);
and U24910 (N_24910,N_17780,N_17219);
and U24911 (N_24911,N_17248,N_19625);
and U24912 (N_24912,N_19000,N_15027);
and U24913 (N_24913,N_16102,N_16661);
nor U24914 (N_24914,N_19584,N_17113);
nand U24915 (N_24915,N_16889,N_19527);
or U24916 (N_24916,N_17813,N_16882);
and U24917 (N_24917,N_19155,N_19805);
nor U24918 (N_24918,N_15467,N_17868);
and U24919 (N_24919,N_18055,N_17967);
and U24920 (N_24920,N_19332,N_18834);
nor U24921 (N_24921,N_19130,N_18315);
or U24922 (N_24922,N_17230,N_16311);
or U24923 (N_24923,N_17049,N_15724);
nand U24924 (N_24924,N_15231,N_16776);
nand U24925 (N_24925,N_19039,N_18615);
nand U24926 (N_24926,N_16033,N_18915);
nor U24927 (N_24927,N_17225,N_19869);
or U24928 (N_24928,N_19264,N_19467);
or U24929 (N_24929,N_15527,N_15995);
or U24930 (N_24930,N_18544,N_17416);
nand U24931 (N_24931,N_16543,N_16036);
nand U24932 (N_24932,N_17500,N_17052);
nor U24933 (N_24933,N_17543,N_15571);
and U24934 (N_24934,N_19142,N_19032);
and U24935 (N_24935,N_18113,N_17200);
or U24936 (N_24936,N_16009,N_16653);
or U24937 (N_24937,N_18682,N_17632);
nand U24938 (N_24938,N_15600,N_15341);
and U24939 (N_24939,N_18694,N_18017);
nand U24940 (N_24940,N_18475,N_16506);
and U24941 (N_24941,N_17566,N_17268);
nor U24942 (N_24942,N_19734,N_15001);
nand U24943 (N_24943,N_19897,N_19864);
nor U24944 (N_24944,N_19309,N_19799);
nand U24945 (N_24945,N_16520,N_17508);
nor U24946 (N_24946,N_17924,N_19488);
nand U24947 (N_24947,N_18491,N_18140);
nand U24948 (N_24948,N_18489,N_18186);
nor U24949 (N_24949,N_15162,N_15485);
or U24950 (N_24950,N_16665,N_15403);
and U24951 (N_24951,N_15428,N_16849);
and U24952 (N_24952,N_16597,N_17212);
nor U24953 (N_24953,N_15668,N_19047);
and U24954 (N_24954,N_19587,N_15912);
nand U24955 (N_24955,N_15464,N_15661);
and U24956 (N_24956,N_18312,N_17464);
nand U24957 (N_24957,N_15052,N_18302);
and U24958 (N_24958,N_18139,N_17794);
xor U24959 (N_24959,N_16709,N_16101);
nand U24960 (N_24960,N_17521,N_17658);
and U24961 (N_24961,N_19310,N_19361);
and U24962 (N_24962,N_19710,N_16899);
and U24963 (N_24963,N_17966,N_15926);
nand U24964 (N_24964,N_15705,N_17060);
and U24965 (N_24965,N_19551,N_19105);
and U24966 (N_24966,N_18607,N_15558);
and U24967 (N_24967,N_17651,N_16027);
or U24968 (N_24968,N_19029,N_18147);
nand U24969 (N_24969,N_19537,N_16528);
or U24970 (N_24970,N_17339,N_17919);
or U24971 (N_24971,N_17205,N_17709);
nand U24972 (N_24972,N_18868,N_18619);
nand U24973 (N_24973,N_19566,N_16126);
or U24974 (N_24974,N_18050,N_19757);
nor U24975 (N_24975,N_17606,N_15351);
nor U24976 (N_24976,N_18324,N_18682);
nand U24977 (N_24977,N_15156,N_18010);
and U24978 (N_24978,N_16667,N_16804);
or U24979 (N_24979,N_18062,N_15200);
or U24980 (N_24980,N_17234,N_19359);
or U24981 (N_24981,N_16799,N_16933);
nor U24982 (N_24982,N_15066,N_19724);
nand U24983 (N_24983,N_19703,N_19766);
and U24984 (N_24984,N_16782,N_17789);
xnor U24985 (N_24985,N_15276,N_16180);
or U24986 (N_24986,N_19006,N_19274);
nor U24987 (N_24987,N_18384,N_18342);
nor U24988 (N_24988,N_18486,N_18567);
or U24989 (N_24989,N_19163,N_18720);
or U24990 (N_24990,N_16177,N_15157);
nor U24991 (N_24991,N_18267,N_19603);
or U24992 (N_24992,N_15092,N_16411);
nand U24993 (N_24993,N_16491,N_19310);
and U24994 (N_24994,N_16455,N_16558);
or U24995 (N_24995,N_18213,N_18448);
or U24996 (N_24996,N_18923,N_19103);
nand U24997 (N_24997,N_15169,N_19323);
or U24998 (N_24998,N_15905,N_16295);
nor U24999 (N_24999,N_17489,N_19597);
nor U25000 (N_25000,N_21259,N_21874);
or U25001 (N_25001,N_24463,N_20707);
and U25002 (N_25002,N_21854,N_22514);
nand U25003 (N_25003,N_21521,N_24930);
or U25004 (N_25004,N_24975,N_20934);
nor U25005 (N_25005,N_23101,N_21714);
nand U25006 (N_25006,N_24137,N_23932);
and U25007 (N_25007,N_23148,N_21876);
or U25008 (N_25008,N_22876,N_24038);
and U25009 (N_25009,N_24406,N_21536);
nand U25010 (N_25010,N_23455,N_22340);
or U25011 (N_25011,N_23430,N_24007);
or U25012 (N_25012,N_23575,N_21716);
nor U25013 (N_25013,N_24123,N_24452);
or U25014 (N_25014,N_20981,N_22626);
or U25015 (N_25015,N_23404,N_24099);
nand U25016 (N_25016,N_24497,N_20401);
nand U25017 (N_25017,N_24556,N_20792);
and U25018 (N_25018,N_22446,N_22616);
nor U25019 (N_25019,N_21687,N_23301);
and U25020 (N_25020,N_20008,N_20869);
nor U25021 (N_25021,N_24086,N_24034);
and U25022 (N_25022,N_23297,N_20931);
nand U25023 (N_25023,N_22144,N_22305);
nand U25024 (N_25024,N_20431,N_20246);
and U25025 (N_25025,N_21050,N_22973);
and U25026 (N_25026,N_20814,N_24672);
nor U25027 (N_25027,N_24052,N_20985);
or U25028 (N_25028,N_21590,N_24788);
and U25029 (N_25029,N_22176,N_24013);
nand U25030 (N_25030,N_23832,N_22563);
nand U25031 (N_25031,N_22078,N_24195);
nand U25032 (N_25032,N_23522,N_22063);
nor U25033 (N_25033,N_22875,N_22966);
and U25034 (N_25034,N_24302,N_21072);
and U25035 (N_25035,N_22957,N_21111);
and U25036 (N_25036,N_23966,N_22062);
nand U25037 (N_25037,N_21449,N_24541);
and U25038 (N_25038,N_20871,N_23850);
or U25039 (N_25039,N_20258,N_24805);
and U25040 (N_25040,N_23459,N_20171);
or U25041 (N_25041,N_24927,N_22800);
or U25042 (N_25042,N_21244,N_23720);
or U25043 (N_25043,N_24409,N_20457);
nand U25044 (N_25044,N_24383,N_23130);
and U25045 (N_25045,N_22233,N_20413);
nor U25046 (N_25046,N_21282,N_23080);
and U25047 (N_25047,N_23047,N_23512);
and U25048 (N_25048,N_24702,N_24339);
or U25049 (N_25049,N_24667,N_24689);
nand U25050 (N_25050,N_20343,N_23225);
nor U25051 (N_25051,N_21517,N_20631);
xnor U25052 (N_25052,N_22110,N_23372);
and U25053 (N_25053,N_22343,N_23154);
and U25054 (N_25054,N_24859,N_20020);
or U25055 (N_25055,N_24062,N_23040);
and U25056 (N_25056,N_24109,N_21226);
or U25057 (N_25057,N_20203,N_24374);
or U25058 (N_25058,N_24950,N_24048);
nor U25059 (N_25059,N_20714,N_21289);
nand U25060 (N_25060,N_23883,N_24447);
and U25061 (N_25061,N_22022,N_24111);
or U25062 (N_25062,N_23707,N_21948);
and U25063 (N_25063,N_24278,N_22678);
nand U25064 (N_25064,N_22808,N_20658);
xnor U25065 (N_25065,N_21233,N_21713);
or U25066 (N_25066,N_20201,N_20996);
nand U25067 (N_25067,N_24623,N_21011);
nand U25068 (N_25068,N_21090,N_24558);
nand U25069 (N_25069,N_20582,N_21962);
nand U25070 (N_25070,N_23897,N_24790);
nand U25071 (N_25071,N_20085,N_24305);
and U25072 (N_25072,N_20075,N_23807);
nand U25073 (N_25073,N_24885,N_21618);
nand U25074 (N_25074,N_23476,N_20746);
or U25075 (N_25075,N_21048,N_23066);
or U25076 (N_25076,N_22243,N_23083);
nand U25077 (N_25077,N_24008,N_21775);
or U25078 (N_25078,N_20054,N_20173);
and U25079 (N_25079,N_20143,N_24088);
nand U25080 (N_25080,N_24502,N_22758);
or U25081 (N_25081,N_22101,N_22042);
nor U25082 (N_25082,N_20100,N_23598);
nand U25083 (N_25083,N_23835,N_23642);
and U25084 (N_25084,N_23032,N_22996);
and U25085 (N_25085,N_24389,N_23189);
or U25086 (N_25086,N_22267,N_21062);
and U25087 (N_25087,N_20466,N_20838);
and U25088 (N_25088,N_21969,N_20427);
nand U25089 (N_25089,N_22582,N_22304);
nor U25090 (N_25090,N_21341,N_23857);
nand U25091 (N_25091,N_21475,N_23118);
or U25092 (N_25092,N_20149,N_23442);
or U25093 (N_25093,N_20526,N_24629);
nand U25094 (N_25094,N_21607,N_23361);
or U25095 (N_25095,N_22794,N_20412);
or U25096 (N_25096,N_20467,N_20132);
or U25097 (N_25097,N_21350,N_24036);
nand U25098 (N_25098,N_23576,N_20529);
and U25099 (N_25099,N_21515,N_21381);
nand U25100 (N_25100,N_22231,N_20933);
nor U25101 (N_25101,N_21802,N_24711);
nor U25102 (N_25102,N_22845,N_24323);
and U25103 (N_25103,N_24461,N_20523);
nand U25104 (N_25104,N_21942,N_23466);
nand U25105 (N_25105,N_24953,N_20177);
nand U25106 (N_25106,N_23098,N_20053);
and U25107 (N_25107,N_23216,N_24526);
and U25108 (N_25108,N_21330,N_23096);
or U25109 (N_25109,N_23458,N_21260);
nor U25110 (N_25110,N_22874,N_22494);
xnor U25111 (N_25111,N_23457,N_20879);
and U25112 (N_25112,N_23518,N_22672);
and U25113 (N_25113,N_24103,N_24039);
nor U25114 (N_25114,N_21809,N_24946);
or U25115 (N_25115,N_20596,N_23676);
and U25116 (N_25116,N_21280,N_22722);
nand U25117 (N_25117,N_22697,N_20813);
nand U25118 (N_25118,N_22389,N_23015);
nor U25119 (N_25119,N_23157,N_24366);
or U25120 (N_25120,N_23334,N_22791);
or U25121 (N_25121,N_24763,N_22702);
nand U25122 (N_25122,N_24792,N_20041);
nor U25123 (N_25123,N_23163,N_24731);
nor U25124 (N_25124,N_23043,N_21377);
nor U25125 (N_25125,N_22669,N_23123);
or U25126 (N_25126,N_22869,N_23462);
and U25127 (N_25127,N_22493,N_22162);
and U25128 (N_25128,N_23552,N_22727);
and U25129 (N_25129,N_21547,N_21840);
and U25130 (N_25130,N_23740,N_22490);
and U25131 (N_25131,N_20946,N_22547);
nor U25132 (N_25132,N_23531,N_22204);
or U25133 (N_25133,N_23501,N_21999);
nor U25134 (N_25134,N_20122,N_21872);
or U25135 (N_25135,N_20183,N_21975);
and U25136 (N_25136,N_20265,N_23197);
nor U25137 (N_25137,N_22263,N_22437);
or U25138 (N_25138,N_22578,N_20205);
nand U25139 (N_25139,N_22533,N_22030);
and U25140 (N_25140,N_24414,N_20924);
nand U25141 (N_25141,N_23823,N_20007);
nand U25142 (N_25142,N_22034,N_21830);
and U25143 (N_25143,N_20713,N_22409);
and U25144 (N_25144,N_24830,N_20352);
nor U25145 (N_25145,N_24379,N_22019);
or U25146 (N_25146,N_21225,N_21601);
or U25147 (N_25147,N_20182,N_21451);
nor U25148 (N_25148,N_20620,N_22033);
and U25149 (N_25149,N_22926,N_23687);
or U25150 (N_25150,N_24733,N_23326);
nand U25151 (N_25151,N_22510,N_20668);
and U25152 (N_25152,N_24259,N_23323);
nor U25153 (N_25153,N_24184,N_21262);
nor U25154 (N_25154,N_23618,N_24762);
nor U25155 (N_25155,N_24954,N_22045);
xor U25156 (N_25156,N_23960,N_23675);
and U25157 (N_25157,N_21976,N_22659);
or U25158 (N_25158,N_20046,N_21150);
nor U25159 (N_25159,N_20174,N_21166);
or U25160 (N_25160,N_24043,N_23600);
or U25161 (N_25161,N_24605,N_24349);
and U25162 (N_25162,N_22413,N_22764);
and U25163 (N_25163,N_20514,N_20312);
nor U25164 (N_25164,N_23848,N_21651);
nor U25165 (N_25165,N_24411,N_22217);
and U25166 (N_25166,N_21699,N_21881);
or U25167 (N_25167,N_24201,N_24371);
or U25168 (N_25168,N_24094,N_20134);
and U25169 (N_25169,N_20801,N_21044);
and U25170 (N_25170,N_20135,N_21479);
or U25171 (N_25171,N_24944,N_22350);
nand U25172 (N_25172,N_21167,N_22431);
or U25173 (N_25173,N_24855,N_21819);
nand U25174 (N_25174,N_22603,N_22576);
and U25175 (N_25175,N_20224,N_23917);
nor U25176 (N_25176,N_21100,N_22302);
and U25177 (N_25177,N_22282,N_24124);
nor U25178 (N_25178,N_24955,N_21114);
and U25179 (N_25179,N_22763,N_24532);
and U25180 (N_25180,N_20260,N_20383);
nand U25181 (N_25181,N_24085,N_21949);
nor U25182 (N_25182,N_22214,N_23093);
and U25183 (N_25183,N_21973,N_23677);
or U25184 (N_25184,N_23353,N_22587);
nor U25185 (N_25185,N_21678,N_22462);
nand U25186 (N_25186,N_23790,N_21439);
nand U25187 (N_25187,N_22887,N_23131);
nand U25188 (N_25188,N_22558,N_21194);
and U25189 (N_25189,N_21836,N_22293);
nand U25190 (N_25190,N_21243,N_20589);
and U25191 (N_25191,N_20039,N_22332);
xor U25192 (N_25192,N_23035,N_23105);
or U25193 (N_25193,N_22347,N_20706);
and U25194 (N_25194,N_21732,N_21423);
nor U25195 (N_25195,N_21772,N_22106);
and U25196 (N_25196,N_21288,N_20870);
or U25197 (N_25197,N_23227,N_21777);
nor U25198 (N_25198,N_20697,N_22252);
or U25199 (N_25199,N_24920,N_24990);
and U25200 (N_25200,N_22219,N_22757);
nor U25201 (N_25201,N_24503,N_20510);
or U25202 (N_25202,N_20210,N_21595);
or U25203 (N_25203,N_22661,N_24555);
and U25204 (N_25204,N_22318,N_22049);
nor U25205 (N_25205,N_23210,N_24444);
nand U25206 (N_25206,N_20393,N_20095);
nor U25207 (N_25207,N_22885,N_20344);
nor U25208 (N_25208,N_22944,N_22084);
nand U25209 (N_25209,N_23138,N_20536);
nand U25210 (N_25210,N_22701,N_24829);
or U25211 (N_25211,N_24773,N_20220);
nor U25212 (N_25212,N_20287,N_21932);
and U25213 (N_25213,N_21118,N_23426);
and U25214 (N_25214,N_23274,N_22386);
nand U25215 (N_25215,N_21035,N_24397);
nand U25216 (N_25216,N_22184,N_20378);
nor U25217 (N_25217,N_23039,N_22141);
nand U25218 (N_25218,N_22333,N_23965);
nand U25219 (N_25219,N_20004,N_23681);
or U25220 (N_25220,N_21101,N_23099);
nor U25221 (N_25221,N_21444,N_20580);
and U25222 (N_25222,N_22325,N_21319);
and U25223 (N_25223,N_24675,N_20573);
xor U25224 (N_25224,N_23029,N_23867);
and U25225 (N_25225,N_24678,N_23170);
or U25226 (N_25226,N_23621,N_21303);
or U25227 (N_25227,N_22767,N_21163);
or U25228 (N_25228,N_20402,N_22164);
nor U25229 (N_25229,N_20010,N_22053);
nand U25230 (N_25230,N_23958,N_20684);
and U25231 (N_25231,N_23436,N_22893);
xnor U25232 (N_25232,N_22391,N_20902);
nor U25233 (N_25233,N_21641,N_22234);
or U25234 (N_25234,N_21508,N_21220);
nor U25235 (N_25235,N_24440,N_22657);
or U25236 (N_25236,N_22301,N_20708);
and U25237 (N_25237,N_20883,N_21941);
nor U25238 (N_25238,N_22650,N_24127);
nor U25239 (N_25239,N_24272,N_22313);
and U25240 (N_25240,N_24893,N_22590);
or U25241 (N_25241,N_23308,N_22262);
and U25242 (N_25242,N_24016,N_21206);
or U25243 (N_25243,N_23685,N_21522);
or U25244 (N_25244,N_22731,N_20281);
nor U25245 (N_25245,N_22930,N_23581);
and U25246 (N_25246,N_24213,N_22645);
or U25247 (N_25247,N_20877,N_20284);
and U25248 (N_25248,N_24514,N_21008);
nor U25249 (N_25249,N_23049,N_24998);
and U25250 (N_25250,N_22883,N_21749);
and U25251 (N_25251,N_21174,N_22717);
nor U25252 (N_25252,N_23403,N_23657);
or U25253 (N_25253,N_21299,N_24698);
or U25254 (N_25254,N_20669,N_24049);
nand U25255 (N_25255,N_21593,N_21895);
and U25256 (N_25256,N_22120,N_22221);
nor U25257 (N_25257,N_21838,N_22787);
xor U25258 (N_25258,N_21145,N_23635);
nor U25259 (N_25259,N_24084,N_23505);
nor U25260 (N_25260,N_24076,N_23938);
or U25261 (N_25261,N_23587,N_23388);
nor U25262 (N_25262,N_22422,N_24751);
nor U25263 (N_25263,N_23773,N_20787);
nand U25264 (N_25264,N_20055,N_20463);
nor U25265 (N_25265,N_22864,N_22173);
and U25266 (N_25266,N_22884,N_20125);
and U25267 (N_25267,N_22891,N_23650);
and U25268 (N_25268,N_22246,N_20590);
or U25269 (N_25269,N_20730,N_24317);
and U25270 (N_25270,N_22297,N_23922);
and U25271 (N_25271,N_22820,N_21318);
nand U25272 (N_25272,N_22421,N_21870);
and U25273 (N_25273,N_24017,N_23482);
and U25274 (N_25274,N_22192,N_22753);
and U25275 (N_25275,N_23427,N_23864);
nor U25276 (N_25276,N_22855,N_23293);
nor U25277 (N_25277,N_23964,N_22236);
and U25278 (N_25278,N_21605,N_23437);
nor U25279 (N_25279,N_21889,N_23846);
nor U25280 (N_25280,N_21834,N_20900);
nand U25281 (N_25281,N_24246,N_22248);
nand U25282 (N_25282,N_24091,N_22417);
and U25283 (N_25283,N_22224,N_24493);
nor U25284 (N_25284,N_20938,N_20334);
and U25285 (N_25285,N_21027,N_24492);
nor U25286 (N_25286,N_20285,N_20718);
nand U25287 (N_25287,N_24468,N_24442);
or U25288 (N_25288,N_20111,N_21129);
nand U25289 (N_25289,N_20929,N_20023);
or U25290 (N_25290,N_22760,N_20342);
and U25291 (N_25291,N_22037,N_24135);
and U25292 (N_25292,N_24288,N_20650);
nor U25293 (N_25293,N_22719,N_24077);
nand U25294 (N_25294,N_24642,N_21457);
and U25295 (N_25295,N_21395,N_21121);
xnor U25296 (N_25296,N_21216,N_24163);
or U25297 (N_25297,N_23934,N_20110);
and U25298 (N_25298,N_23181,N_24289);
nor U25299 (N_25299,N_23557,N_24165);
nand U25300 (N_25300,N_24544,N_20230);
or U25301 (N_25301,N_23012,N_24981);
nand U25302 (N_25302,N_20876,N_20719);
and U25303 (N_25303,N_22088,N_24173);
and U25304 (N_25304,N_21015,N_24237);
or U25305 (N_25305,N_20569,N_21806);
nand U25306 (N_25306,N_21599,N_20915);
or U25307 (N_25307,N_23754,N_20836);
nor U25308 (N_25308,N_20222,N_21738);
nor U25309 (N_25309,N_21655,N_22668);
nand U25310 (N_25310,N_24931,N_20350);
or U25311 (N_25311,N_22539,N_22593);
nor U25312 (N_25312,N_20227,N_22715);
or U25313 (N_25313,N_21446,N_22782);
nand U25314 (N_25314,N_20070,N_24400);
nor U25315 (N_25315,N_22423,N_23777);
or U25316 (N_25316,N_20537,N_20791);
nor U25317 (N_25317,N_23359,N_23381);
and U25318 (N_25318,N_23000,N_24121);
and U25319 (N_25319,N_21630,N_23240);
xnor U25320 (N_25320,N_21789,N_20614);
nor U25321 (N_25321,N_22210,N_23986);
nor U25322 (N_25322,N_20190,N_20442);
or U25323 (N_25323,N_24636,N_21316);
and U25324 (N_25324,N_23726,N_20270);
xnor U25325 (N_25325,N_21549,N_21940);
nor U25326 (N_25326,N_22512,N_20256);
or U25327 (N_25327,N_20586,N_22823);
or U25328 (N_25328,N_21074,N_24102);
and U25329 (N_25329,N_21808,N_20408);
nor U25330 (N_25330,N_20865,N_23653);
and U25331 (N_25331,N_23818,N_20616);
nand U25332 (N_25332,N_21211,N_21017);
and U25333 (N_25333,N_20675,N_22553);
or U25334 (N_25334,N_24772,N_23881);
or U25335 (N_25335,N_22759,N_24546);
nand U25336 (N_25336,N_22693,N_21826);
and U25337 (N_25337,N_22003,N_20604);
and U25338 (N_25338,N_21463,N_21705);
and U25339 (N_25339,N_23627,N_23943);
and U25340 (N_25340,N_22390,N_23034);
nor U25341 (N_25341,N_22433,N_20180);
nand U25342 (N_25342,N_23752,N_21286);
nor U25343 (N_25343,N_22906,N_20678);
nor U25344 (N_25344,N_22972,N_21231);
nand U25345 (N_25345,N_23324,N_23314);
nor U25346 (N_25346,N_23787,N_23448);
nor U25347 (N_25347,N_23561,N_23959);
and U25348 (N_25348,N_20819,N_20138);
xor U25349 (N_25349,N_22359,N_20123);
nand U25350 (N_25350,N_24040,N_23056);
and U25351 (N_25351,N_22048,N_23254);
nor U25352 (N_25352,N_21223,N_20083);
and U25353 (N_25353,N_23780,N_23363);
nor U25354 (N_25354,N_20490,N_21077);
or U25355 (N_25355,N_22070,N_23665);
and U25356 (N_25356,N_21563,N_22707);
nor U25357 (N_25357,N_24391,N_22994);
and U25358 (N_25358,N_20047,N_23534);
nor U25359 (N_25359,N_20269,N_22969);
or U25360 (N_25360,N_20237,N_23304);
and U25361 (N_25361,N_20852,N_21425);
nor U25362 (N_25362,N_23615,N_24941);
nand U25363 (N_25363,N_21113,N_22585);
or U25364 (N_25364,N_20120,N_23198);
or U25365 (N_25365,N_23266,N_23348);
and U25366 (N_25366,N_20729,N_21695);
or U25367 (N_25367,N_20919,N_20331);
nor U25368 (N_25368,N_22206,N_24224);
and U25369 (N_25369,N_21155,N_22240);
or U25370 (N_25370,N_23262,N_23494);
and U25371 (N_25371,N_24670,N_20608);
or U25372 (N_25372,N_21362,N_20997);
nand U25373 (N_25373,N_20844,N_24153);
and U25374 (N_25374,N_24175,N_20420);
nand U25375 (N_25375,N_23102,N_22145);
nor U25376 (N_25376,N_20648,N_24136);
nor U25377 (N_25377,N_23340,N_20019);
nand U25378 (N_25378,N_24170,N_23866);
or U25379 (N_25379,N_20323,N_21963);
and U25380 (N_25380,N_20519,N_22244);
nand U25381 (N_25381,N_21723,N_24186);
and U25382 (N_25382,N_21068,N_21614);
or U25383 (N_25383,N_23994,N_22600);
nor U25384 (N_25384,N_20228,N_24700);
nor U25385 (N_25385,N_23120,N_23202);
and U25386 (N_25386,N_20073,N_23828);
nor U25387 (N_25387,N_22150,N_20610);
and U25388 (N_25388,N_22382,N_21409);
nor U25389 (N_25389,N_21421,N_21082);
or U25390 (N_25390,N_24467,N_24756);
nor U25391 (N_25391,N_23239,N_20563);
or U25392 (N_25392,N_21739,N_20759);
or U25393 (N_25393,N_20899,N_20179);
and U25394 (N_25394,N_24348,N_21671);
nand U25395 (N_25395,N_24735,N_23298);
or U25396 (N_25396,N_23774,N_21525);
nor U25397 (N_25397,N_22454,N_21904);
nand U25398 (N_25398,N_22928,N_24612);
and U25399 (N_25399,N_22812,N_21915);
or U25400 (N_25400,N_20845,N_21060);
or U25401 (N_25401,N_24239,N_24316);
nand U25402 (N_25402,N_21368,N_20487);
nand U25403 (N_25403,N_24872,N_21825);
and U25404 (N_25404,N_24852,N_24067);
nor U25405 (N_25405,N_24697,N_21300);
nand U25406 (N_25406,N_21755,N_22843);
nand U25407 (N_25407,N_21589,N_24041);
and U25408 (N_25408,N_21136,N_20984);
nand U25409 (N_25409,N_20327,N_22771);
nor U25410 (N_25410,N_24641,N_22324);
and U25411 (N_25411,N_21091,N_20722);
or U25412 (N_25412,N_22021,N_21038);
or U25413 (N_25413,N_23954,N_23387);
nor U25414 (N_25414,N_23259,N_20990);
nand U25415 (N_25415,N_24842,N_20705);
or U25416 (N_25416,N_24659,N_23710);
nor U25417 (N_25417,N_21222,N_21663);
nand U25418 (N_25418,N_22830,N_24505);
nor U25419 (N_25419,N_21466,N_20375);
nand U25420 (N_25420,N_20198,N_23977);
nand U25421 (N_25421,N_22504,N_22071);
and U25422 (N_25422,N_20065,N_21752);
and U25423 (N_25423,N_21415,N_24285);
or U25424 (N_25424,N_23516,N_20774);
nand U25425 (N_25425,N_21042,N_22201);
nand U25426 (N_25426,N_20704,N_23059);
nand U25427 (N_25427,N_22414,N_23868);
or U25428 (N_25428,N_21748,N_23729);
and U25429 (N_25429,N_23432,N_23255);
and U25430 (N_25430,N_22054,N_23944);
and U25431 (N_25431,N_22117,N_24644);
and U25432 (N_25432,N_22841,N_20379);
and U25433 (N_25433,N_23822,N_24064);
nand U25434 (N_25434,N_21472,N_24924);
and U25435 (N_25435,N_22997,N_21998);
nor U25436 (N_25436,N_20479,N_21712);
nand U25437 (N_25437,N_24340,N_24079);
nand U25438 (N_25438,N_21363,N_20766);
nand U25439 (N_25439,N_21458,N_20346);
nand U25440 (N_25440,N_24897,N_21721);
and U25441 (N_25441,N_21551,N_24147);
nand U25442 (N_25442,N_21600,N_23444);
nor U25443 (N_25443,N_22136,N_24128);
nor U25444 (N_25444,N_21147,N_21644);
nor U25445 (N_25445,N_23305,N_20967);
nand U25446 (N_25446,N_20842,N_21546);
nand U25447 (N_25447,N_24158,N_23660);
nand U25448 (N_25448,N_21627,N_20016);
and U25449 (N_25449,N_20347,N_24218);
or U25450 (N_25450,N_22113,N_23160);
nor U25451 (N_25451,N_23052,N_24949);
or U25452 (N_25452,N_21428,N_23833);
or U25453 (N_25453,N_23510,N_23941);
nand U25454 (N_25454,N_20630,N_24032);
nor U25455 (N_25455,N_20821,N_24011);
nand U25456 (N_25456,N_23747,N_22082);
nand U25457 (N_25457,N_22599,N_22962);
and U25458 (N_25458,N_23915,N_21844);
or U25459 (N_25459,N_23018,N_23357);
or U25460 (N_25460,N_20611,N_24940);
and U25461 (N_25461,N_20504,N_20175);
or U25462 (N_25462,N_24705,N_22889);
nor U25463 (N_25463,N_23139,N_21394);
nand U25464 (N_25464,N_21726,N_24899);
and U25465 (N_25465,N_21464,N_20460);
nand U25466 (N_25466,N_22641,N_22909);
nand U25467 (N_25467,N_23711,N_21424);
nand U25468 (N_25468,N_24009,N_20196);
nor U25469 (N_25469,N_23208,N_21661);
or U25470 (N_25470,N_22220,N_21445);
nor U25471 (N_25471,N_24518,N_20989);
nor U25472 (N_25472,N_23005,N_24042);
nand U25473 (N_25473,N_20006,N_23634);
or U25474 (N_25474,N_21568,N_21304);
nor U25475 (N_25475,N_23321,N_22270);
xor U25476 (N_25476,N_21725,N_23639);
nor U25477 (N_25477,N_23555,N_24531);
nor U25478 (N_25478,N_22087,N_21039);
and U25479 (N_25479,N_21153,N_23733);
and U25480 (N_25480,N_21855,N_23011);
nand U25481 (N_25481,N_20937,N_20142);
or U25482 (N_25482,N_22654,N_24807);
nand U25483 (N_25483,N_21139,N_24879);
nor U25484 (N_25484,N_20002,N_20394);
or U25485 (N_25485,N_20272,N_23767);
or U25486 (N_25486,N_24203,N_20374);
or U25487 (N_25487,N_22061,N_23036);
or U25488 (N_25488,N_22663,N_20325);
and U25489 (N_25489,N_23182,N_21189);
and U25490 (N_25490,N_22676,N_23207);
nor U25491 (N_25491,N_23471,N_23201);
nand U25492 (N_25492,N_23511,N_24806);
nand U25493 (N_25493,N_24620,N_23153);
and U25494 (N_25494,N_22026,N_20191);
nor U25495 (N_25495,N_23873,N_22074);
nor U25496 (N_25496,N_22273,N_20972);
or U25497 (N_25497,N_23434,N_24567);
nand U25498 (N_25498,N_21970,N_20619);
nor U25499 (N_25499,N_23062,N_22059);
nor U25500 (N_25500,N_22964,N_23535);
or U25501 (N_25501,N_20570,N_24537);
or U25502 (N_25502,N_21078,N_22961);
nor U25503 (N_25503,N_22230,N_20715);
nand U25504 (N_25504,N_23452,N_24972);
nor U25505 (N_25505,N_24129,N_20951);
nor U25506 (N_25506,N_23423,N_22981);
nand U25507 (N_25507,N_22942,N_21996);
and U25508 (N_25508,N_22465,N_20056);
nor U25509 (N_25509,N_20238,N_23662);
nand U25510 (N_25510,N_22695,N_24797);
or U25511 (N_25511,N_22453,N_20261);
and U25512 (N_25512,N_20979,N_21388);
and U25513 (N_25513,N_20508,N_23741);
nor U25514 (N_25514,N_24631,N_24568);
nand U25515 (N_25515,N_21640,N_23050);
nand U25516 (N_25516,N_22369,N_21955);
and U25517 (N_25517,N_20927,N_23414);
and U25518 (N_25518,N_24704,N_22259);
nor U25519 (N_25519,N_23933,N_24789);
and U25520 (N_25520,N_22000,N_23316);
and U25521 (N_25521,N_22796,N_21240);
nand U25522 (N_25522,N_20126,N_21376);
nand U25523 (N_25523,N_20782,N_20396);
nor U25524 (N_25524,N_20683,N_20109);
and U25525 (N_25525,N_20738,N_22484);
nor U25526 (N_25526,N_24952,N_23593);
or U25527 (N_25527,N_23547,N_22967);
or U25528 (N_25528,N_23900,N_21771);
and U25529 (N_25529,N_24291,N_23121);
or U25530 (N_25530,N_23158,N_22403);
nand U25531 (N_25531,N_24725,N_24833);
and U25532 (N_25532,N_23524,N_24404);
nand U25533 (N_25533,N_22529,N_22451);
and U25534 (N_25534,N_23185,N_20674);
xor U25535 (N_25535,N_20806,N_22648);
or U25536 (N_25536,N_20425,N_24431);
nand U25537 (N_25537,N_21993,N_23808);
and U25538 (N_25538,N_22188,N_24583);
nand U25539 (N_25539,N_22570,N_20890);
nor U25540 (N_25540,N_21140,N_23537);
nor U25541 (N_25541,N_21403,N_22773);
nand U25542 (N_25542,N_22573,N_21953);
nor U25543 (N_25543,N_20688,N_21681);
nand U25544 (N_25544,N_20308,N_22847);
nor U25545 (N_25545,N_22017,N_24607);
nor U25546 (N_25546,N_23124,N_24309);
or U25547 (N_25547,N_20816,N_21770);
nor U25548 (N_25548,N_22480,N_22018);
or U25549 (N_25549,N_24880,N_21071);
and U25550 (N_25550,N_20213,N_20454);
nor U25551 (N_25551,N_24988,N_20363);
nand U25552 (N_25552,N_20236,N_23195);
nand U25553 (N_25553,N_23186,N_20861);
nor U25554 (N_25554,N_24914,N_22671);
or U25555 (N_25555,N_21615,N_24318);
nand U25556 (N_25556,N_21542,N_20282);
nor U25557 (N_25557,N_23284,N_20702);
nand U25558 (N_25558,N_20037,N_20194);
and U25559 (N_25559,N_21971,N_22726);
nand U25560 (N_25560,N_20133,N_23987);
or U25561 (N_25561,N_21559,N_21359);
nor U25562 (N_25562,N_23193,N_22025);
nor U25563 (N_25563,N_20313,N_22163);
and U25564 (N_25564,N_22742,N_20263);
or U25565 (N_25565,N_24822,N_22829);
or U25566 (N_25566,N_24257,N_21528);
nor U25567 (N_25567,N_23990,N_24143);
nor U25568 (N_25568,N_20072,N_24621);
and U25569 (N_25569,N_24229,N_21910);
nor U25570 (N_25570,N_21053,N_22099);
or U25571 (N_25571,N_22860,N_20680);
nor U25572 (N_25572,N_21676,N_24437);
or U25573 (N_25573,N_22354,N_23451);
or U25574 (N_25574,N_20975,N_23885);
and U25575 (N_25575,N_22900,N_22276);
nand U25576 (N_25576,N_21985,N_20485);
nand U25577 (N_25577,N_22550,N_20643);
nor U25578 (N_25578,N_23863,N_24301);
and U25579 (N_25579,N_21566,N_23980);
xnor U25580 (N_25580,N_24275,N_21076);
nand U25581 (N_25581,N_20336,N_21503);
and U25582 (N_25582,N_24392,N_24581);
nor U25583 (N_25583,N_22769,N_23378);
and U25584 (N_25584,N_20847,N_22039);
nand U25585 (N_25585,N_21779,N_24355);
nor U25586 (N_25586,N_24610,N_24458);
and U25587 (N_25587,N_24650,N_24554);
nor U25588 (N_25588,N_24274,N_24664);
and U25589 (N_25589,N_20435,N_20048);
or U25590 (N_25590,N_24489,N_24139);
and U25591 (N_25591,N_21407,N_20184);
and U25592 (N_25592,N_24867,N_23289);
nor U25593 (N_25593,N_20851,N_24810);
or U25594 (N_25594,N_22666,N_24796);
or U25595 (N_25595,N_22687,N_20728);
or U25596 (N_25596,N_23930,N_23415);
nand U25597 (N_25597,N_24417,N_22924);
nand U25598 (N_25598,N_20763,N_23375);
nand U25599 (N_25599,N_24480,N_21786);
nor U25600 (N_25600,N_23486,N_20044);
or U25601 (N_25601,N_22473,N_24324);
nand U25602 (N_25602,N_20148,N_20274);
or U25603 (N_25603,N_20178,N_23242);
and U25604 (N_25604,N_23901,N_22457);
nor U25605 (N_25605,N_21518,N_24277);
nor U25606 (N_25606,N_22915,N_20321);
and U25607 (N_25607,N_20038,N_23580);
nor U25608 (N_25608,N_22850,N_24179);
nor U25609 (N_25609,N_21670,N_22128);
and U25610 (N_25610,N_22890,N_21979);
and U25611 (N_25611,N_22977,N_21656);
nor U25612 (N_25612,N_22978,N_23241);
or U25613 (N_25613,N_23602,N_22310);
nand U25614 (N_25614,N_24821,N_21711);
nor U25615 (N_25615,N_23596,N_23995);
and U25616 (N_25616,N_22186,N_22351);
nor U25617 (N_25617,N_21398,N_23608);
or U25618 (N_25618,N_22694,N_22381);
nor U25619 (N_25619,N_24826,N_22225);
and U25620 (N_25620,N_23936,N_24803);
or U25621 (N_25621,N_24742,N_23125);
and U25622 (N_25622,N_23290,N_24611);
and U25623 (N_25623,N_22873,N_24584);
or U25624 (N_25624,N_20219,N_20468);
nor U25625 (N_25625,N_24044,N_23057);
xor U25626 (N_25626,N_22211,N_20369);
or U25627 (N_25627,N_24881,N_24385);
nor U25628 (N_25628,N_21096,N_22877);
nor U25629 (N_25629,N_23558,N_21066);
and U25630 (N_25630,N_23709,N_22713);
or U25631 (N_25631,N_20243,N_23858);
nor U25632 (N_25632,N_24222,N_24134);
or U25633 (N_25633,N_21850,N_23560);
nor U25634 (N_25634,N_21019,N_21702);
and U25635 (N_25635,N_23470,N_23276);
and U25636 (N_25636,N_23073,N_22430);
and U25637 (N_25637,N_24622,N_21724);
nand U25638 (N_25638,N_23519,N_21258);
and U25639 (N_25639,N_24529,N_21868);
or U25640 (N_25640,N_22126,N_24980);
nand U25641 (N_25641,N_20864,N_21583);
nand U25642 (N_25642,N_24767,N_20241);
nor U25643 (N_25643,N_20885,N_21734);
or U25644 (N_25644,N_21162,N_21137);
or U25645 (N_25645,N_20493,N_24652);
nor U25646 (N_25646,N_21089,N_21190);
nor U25647 (N_25647,N_24818,N_24341);
nor U25648 (N_25648,N_21875,N_22828);
nor U25649 (N_25649,N_21731,N_21498);
and U25650 (N_25650,N_21433,N_23887);
nor U25651 (N_25651,N_23937,N_23700);
and U25652 (N_25652,N_21146,N_20654);
or U25653 (N_25653,N_24591,N_23795);
nand U25654 (N_25654,N_20306,N_24096);
nor U25655 (N_25655,N_24978,N_24560);
nor U25656 (N_25656,N_24466,N_23076);
nand U25657 (N_25657,N_21894,N_20686);
or U25658 (N_25658,N_21954,N_20949);
nor U25659 (N_25659,N_22254,N_24926);
or U25660 (N_25660,N_24979,N_21584);
nand U25661 (N_25661,N_22119,N_20857);
or U25662 (N_25662,N_21818,N_22315);
or U25663 (N_25663,N_22849,N_24194);
or U25664 (N_25664,N_22478,N_20469);
or U25665 (N_25665,N_20348,N_24423);
or U25666 (N_25666,N_24888,N_23142);
nor U25667 (N_25667,N_23703,N_24148);
and U25668 (N_25668,N_23604,N_23801);
nand U25669 (N_25669,N_20925,N_21758);
nor U25670 (N_25670,N_22709,N_22999);
and U25671 (N_25671,N_21925,N_20271);
and U25672 (N_25672,N_23295,N_24401);
nand U25673 (N_25673,N_20944,N_23312);
and U25674 (N_25674,N_21672,N_23691);
nor U25675 (N_25675,N_24308,N_23758);
or U25676 (N_25676,N_23380,N_24112);
nand U25677 (N_25677,N_20330,N_20316);
or U25678 (N_25678,N_20474,N_21392);
and U25679 (N_25679,N_24247,N_24310);
xor U25680 (N_25680,N_22123,N_24633);
and U25681 (N_25681,N_22639,N_23008);
or U25682 (N_25682,N_22443,N_23238);
xnor U25683 (N_25683,N_23410,N_22840);
or U25684 (N_25684,N_20226,N_23332);
nand U25685 (N_25685,N_23134,N_20058);
xnor U25686 (N_25686,N_23661,N_24072);
and U25687 (N_25687,N_22073,N_24066);
or U25688 (N_25688,N_22072,N_22602);
nand U25689 (N_25689,N_20696,N_24696);
nand U25690 (N_25690,N_23496,N_21345);
nand U25691 (N_25691,N_23659,N_20693);
nor U25692 (N_25692,N_21582,N_24413);
and U25693 (N_25693,N_22816,N_22203);
or U25694 (N_25694,N_20388,N_20455);
nor U25695 (N_25695,N_23506,N_24080);
nor U25696 (N_25696,N_22245,N_22392);
nand U25697 (N_25697,N_21497,N_21324);
nand U25698 (N_25698,N_24189,N_20558);
nor U25699 (N_25699,N_22502,N_24669);
or U25700 (N_25700,N_23893,N_20986);
and U25701 (N_25701,N_20912,N_20419);
nor U25702 (N_25702,N_21866,N_24595);
nand U25703 (N_25703,N_21252,N_23465);
nor U25704 (N_25704,N_22817,N_23956);
and U25705 (N_25705,N_20862,N_20494);
and U25706 (N_25706,N_21863,N_20541);
or U25707 (N_25707,N_22095,N_21108);
or U25708 (N_25708,N_23009,N_22776);
and U25709 (N_25709,N_24019,N_24215);
nand U25710 (N_25710,N_20968,N_21097);
or U25711 (N_25711,N_23344,N_24145);
or U25712 (N_25712,N_23004,N_21307);
nand U25713 (N_25713,N_23870,N_20128);
or U25714 (N_25714,N_23667,N_21922);
or U25715 (N_25715,N_21624,N_24601);
nor U25716 (N_25716,N_22407,N_23408);
nor U25717 (N_25717,N_21513,N_22482);
nand U25718 (N_25718,N_21440,N_22945);
nand U25719 (N_25719,N_23983,N_23513);
nand U25720 (N_25720,N_22975,N_20682);
or U25721 (N_25721,N_21063,N_24837);
and U25722 (N_25722,N_24098,N_20145);
and U25723 (N_25723,N_24439,N_21170);
nor U25724 (N_25724,N_23477,N_22290);
and U25725 (N_25725,N_23281,N_23840);
or U25726 (N_25726,N_22257,N_23841);
or U25727 (N_25727,N_24875,N_21411);
or U25728 (N_25728,N_20600,N_22345);
or U25729 (N_25729,N_24684,N_21093);
nand U25730 (N_25730,N_24845,N_21893);
and U25731 (N_25731,N_22135,N_22207);
or U25732 (N_25732,N_21117,N_20429);
nand U25733 (N_25733,N_23027,N_22452);
nor U25734 (N_25734,N_21061,N_21543);
and U25735 (N_25735,N_24478,N_21857);
or U25736 (N_25736,N_22867,N_21294);
nor U25737 (N_25737,N_22744,N_24198);
nand U25738 (N_25738,N_20562,N_21249);
nand U25739 (N_25739,N_24053,N_24045);
or U25740 (N_25740,N_22598,N_23540);
or U25741 (N_25741,N_21340,N_23542);
nand U25742 (N_25742,N_23765,N_24917);
and U25743 (N_25743,N_24510,N_24766);
nor U25744 (N_25744,N_24590,N_21805);
nor U25745 (N_25745,N_20119,N_24866);
and U25746 (N_25746,N_22634,N_23178);
and U25747 (N_25747,N_21933,N_20141);
nor U25748 (N_25748,N_24242,N_23699);
nand U25749 (N_25749,N_22294,N_23500);
xor U25750 (N_25750,N_20507,N_22109);
or U25751 (N_25751,N_23782,N_21968);
and U25752 (N_25752,N_20601,N_22652);
nand U25753 (N_25753,N_21196,N_23069);
nor U25754 (N_25754,N_23683,N_20303);
nand U25755 (N_25755,N_23212,N_22295);
and U25756 (N_25756,N_22683,N_21256);
nor U25757 (N_25757,N_21852,N_23368);
or U25758 (N_25758,N_20011,N_23632);
or U25759 (N_25759,N_23784,N_20955);
or U25760 (N_25760,N_20703,N_23815);
and U25761 (N_25761,N_22266,N_23313);
nand U25762 (N_25762,N_20999,N_22689);
nor U25763 (N_25763,N_23251,N_21247);
or U25764 (N_25764,N_20913,N_22498);
nand U25765 (N_25765,N_24566,N_21759);
or U25766 (N_25766,N_20181,N_20595);
or U25767 (N_25767,N_23628,N_24942);
nand U25768 (N_25768,N_21210,N_21760);
and U25769 (N_25769,N_23859,N_22752);
and U25770 (N_25770,N_22948,N_20607);
and U25771 (N_25771,N_21810,N_22277);
nand U25772 (N_25772,N_24141,N_24002);
and U25773 (N_25773,N_22447,N_23961);
xnor U25774 (N_25774,N_20948,N_21138);
nor U25775 (N_25775,N_23695,N_24270);
and U25776 (N_25776,N_22339,N_23847);
and U25777 (N_25777,N_24811,N_20077);
nand U25778 (N_25778,N_21682,N_21966);
or U25779 (N_25779,N_24192,N_22564);
nand U25780 (N_25780,N_21718,N_24450);
nand U25781 (N_25781,N_23345,N_21023);
nand U25782 (N_25782,N_20176,N_20547);
and U25783 (N_25783,N_21329,N_21353);
and U25784 (N_25784,N_24857,N_21529);
or U25785 (N_25785,N_20403,N_21990);
and U25786 (N_25786,N_20150,N_21199);
nor U25787 (N_25787,N_20473,N_24630);
nand U25788 (N_25788,N_22559,N_22953);
or U25789 (N_25789,N_20297,N_21418);
or U25790 (N_25790,N_23971,N_21310);
nand U25791 (N_25791,N_20893,N_24187);
and U25792 (N_25792,N_24527,N_24370);
nand U25793 (N_25793,N_24848,N_24312);
and U25794 (N_25794,N_23217,N_23493);
nor U25795 (N_25795,N_20815,N_23809);
nand U25796 (N_25796,N_23713,N_23963);
nor U25797 (N_25797,N_21505,N_24538);
or U25798 (N_25798,N_24759,N_21822);
and U25799 (N_25799,N_20755,N_22515);
or U25800 (N_25800,N_20882,N_24435);
nand U25801 (N_25801,N_24543,N_22699);
nand U25802 (N_25802,N_24364,N_21526);
or U25803 (N_25803,N_23294,N_23164);
and U25804 (N_25804,N_21030,N_24655);
and U25805 (N_25805,N_22517,N_24516);
or U25806 (N_25806,N_21198,N_24369);
nand U25807 (N_25807,N_22762,N_22610);
nor U25808 (N_25808,N_22894,N_21031);
nand U25809 (N_25809,N_21331,N_21467);
nand U25810 (N_25810,N_23722,N_22024);
nand U25811 (N_25811,N_20209,N_24280);
and U25812 (N_25812,N_23146,N_24345);
or U25813 (N_25813,N_22066,N_24779);
and U25814 (N_25814,N_23439,N_22436);
nand U25815 (N_25815,N_22432,N_22910);
nor U25816 (N_25816,N_22971,N_22079);
xnor U25817 (N_25817,N_22187,N_20254);
nand U25818 (N_25818,N_23655,N_22834);
and U25819 (N_25819,N_20302,N_20012);
or U25820 (N_25820,N_21301,N_21311);
nor U25821 (N_25821,N_22611,N_23222);
nand U25822 (N_25822,N_23053,N_24376);
and U25823 (N_25823,N_20521,N_23258);
or U25824 (N_25824,N_21654,N_21719);
or U25825 (N_25825,N_21264,N_23233);
nand U25826 (N_25826,N_24943,N_20822);
nand U25827 (N_25827,N_23834,N_22623);
or U25828 (N_25828,N_22756,N_24271);
and U25829 (N_25829,N_21184,N_24107);
and U25830 (N_25830,N_21846,N_23243);
nor U25831 (N_25831,N_21486,N_24281);
and U25832 (N_25832,N_20780,N_22835);
nand U25833 (N_25833,N_24081,N_20300);
nor U25834 (N_25834,N_22068,N_21176);
nand U25835 (N_25835,N_21860,N_20994);
nand U25836 (N_25836,N_24434,N_21187);
nand U25837 (N_25837,N_20160,N_24232);
nand U25838 (N_25838,N_22229,N_22179);
or U25839 (N_25839,N_22007,N_24801);
or U25840 (N_25840,N_23640,N_20377);
nand U25841 (N_25841,N_24416,N_24718);
nor U25842 (N_25842,N_23256,N_20731);
and U25843 (N_25843,N_24230,N_20456);
nand U25844 (N_25844,N_22822,N_20118);
or U25845 (N_25845,N_20362,N_22441);
nor U25846 (N_25846,N_20291,N_21130);
nor U25847 (N_25847,N_22704,N_20089);
nor U25848 (N_25848,N_22985,N_23637);
or U25849 (N_25849,N_23589,N_22196);
or U25850 (N_25850,N_21983,N_22781);
or U25851 (N_25851,N_22253,N_22525);
nor U25852 (N_25852,N_21765,N_21177);
and U25853 (N_25853,N_21004,N_21132);
or U25854 (N_25854,N_22786,N_21046);
nor U25855 (N_25855,N_24637,N_23910);
or U25856 (N_25856,N_24286,N_20840);
nor U25857 (N_25857,N_24344,N_24551);
or U25858 (N_25858,N_23422,N_21858);
nor U25859 (N_25859,N_21685,N_22537);
and U25860 (N_25860,N_24562,N_21692);
nand U25861 (N_25861,N_21427,N_20627);
nor U25862 (N_25862,N_21065,N_21814);
nand U25863 (N_25863,N_24732,N_22631);
or U25864 (N_25864,N_24891,N_20671);
nand U25865 (N_25865,N_23539,N_23371);
nor U25866 (N_25866,N_20169,N_24329);
nand U25867 (N_25867,N_21828,N_21164);
nand U25868 (N_25868,N_22425,N_20954);
nor U25869 (N_25869,N_22083,N_22991);
nor U25870 (N_25870,N_21709,N_24282);
and U25871 (N_25871,N_20699,N_21235);
nor U25872 (N_25872,N_23369,N_20672);
or U25873 (N_25873,N_23664,N_20908);
and U25874 (N_25874,N_22530,N_22401);
and U25875 (N_25875,N_22788,N_23877);
or U25876 (N_25876,N_23112,N_23612);
nor U25877 (N_25877,N_20170,N_20633);
nor U25878 (N_25878,N_22092,N_21124);
or U25879 (N_25879,N_20794,N_23952);
nand U25880 (N_25880,N_24075,N_24074);
nand U25881 (N_25881,N_20475,N_24656);
and U25882 (N_25882,N_24907,N_23122);
and U25883 (N_25883,N_24105,N_21401);
and U25884 (N_25884,N_23578,N_21609);
and U25885 (N_25885,N_23646,N_21965);
and U25886 (N_25886,N_24304,N_21763);
and U25887 (N_25887,N_22222,N_20584);
and U25888 (N_25888,N_21684,N_21084);
or U25889 (N_25889,N_24812,N_22522);
or U25890 (N_25890,N_21354,N_20232);
nand U25891 (N_25891,N_24559,N_24660);
nor U25892 (N_25892,N_20761,N_24033);
nand U25893 (N_25893,N_24156,N_20542);
or U25894 (N_25894,N_22040,N_20154);
or U25895 (N_25895,N_24248,N_20317);
nand U25896 (N_25896,N_23443,N_23853);
and U25897 (N_25897,N_22698,N_21613);
or U25898 (N_25898,N_24328,N_20886);
and U25899 (N_25899,N_20881,N_23268);
nor U25900 (N_25900,N_23606,N_23614);
nand U25901 (N_25901,N_22851,N_23727);
nand U25902 (N_25902,N_22151,N_21835);
and U25903 (N_25903,N_21183,N_20267);
nand U25904 (N_25904,N_21298,N_21790);
nor U25905 (N_25905,N_21144,N_22632);
nand U25906 (N_25906,N_20197,N_22004);
or U25907 (N_25907,N_21921,N_22922);
nor U25908 (N_25908,N_23065,N_21861);
nand U25909 (N_25909,N_21813,N_24266);
or U25910 (N_25910,N_24739,N_22583);
nor U25911 (N_25911,N_24178,N_20543);
and U25912 (N_25912,N_24500,N_24018);
nor U25913 (N_25913,N_23082,N_20292);
and U25914 (N_25914,N_23409,N_23947);
and U25915 (N_25915,N_22387,N_20528);
nand U25916 (N_25916,N_21195,N_22655);
nand U25917 (N_25917,N_24983,N_23309);
nor U25918 (N_25918,N_20634,N_23137);
nor U25919 (N_25919,N_23147,N_20288);
and U25920 (N_25920,N_24149,N_23026);
and U25921 (N_25921,N_20914,N_22677);
nand U25922 (N_25922,N_22614,N_24984);
nand U25923 (N_25923,N_23191,N_21273);
or U25924 (N_25924,N_21891,N_21978);
or U25925 (N_25925,N_21477,N_22597);
nand U25926 (N_25926,N_24494,N_21639);
and U25927 (N_25927,N_21625,N_22296);
and U25928 (N_25928,N_24545,N_22509);
and U25929 (N_25929,N_23802,N_23090);
or U25930 (N_25930,N_22912,N_24429);
nand U25931 (N_25931,N_20422,N_22714);
or U25932 (N_25932,N_22384,N_23880);
and U25933 (N_25933,N_20767,N_21629);
nor U25934 (N_25934,N_22388,N_22907);
nand U25935 (N_25935,N_22197,N_24864);
and U25936 (N_25936,N_24381,N_20640);
or U25937 (N_25937,N_24342,N_21634);
nand U25938 (N_25938,N_24746,N_22419);
nor U25939 (N_25939,N_24150,N_22335);
nand U25940 (N_25940,N_21504,N_20112);
nor U25941 (N_25941,N_23678,N_23166);
and U25942 (N_25942,N_20834,N_20962);
nand U25943 (N_25943,N_23920,N_23748);
nor U25944 (N_25944,N_23224,N_24957);
and U25945 (N_25945,N_24575,N_22194);
nand U25946 (N_25946,N_24691,N_22705);
nor U25947 (N_25947,N_24923,N_23079);
and U25948 (N_25948,N_21553,N_22751);
or U25949 (N_25949,N_24771,N_24540);
or U25950 (N_25950,N_20527,N_22002);
or U25951 (N_25951,N_20653,N_20549);
nand U25952 (N_25952,N_23303,N_23742);
or U25953 (N_25953,N_20404,N_23872);
and U25954 (N_25954,N_23844,N_22142);
nand U25955 (N_25955,N_22501,N_22056);
or U25956 (N_25956,N_21218,N_20152);
and U25957 (N_25957,N_22132,N_24116);
nor U25958 (N_25958,N_23060,N_21156);
nor U25959 (N_25959,N_21902,N_23636);
nor U25960 (N_25960,N_21913,N_22306);
nand U25961 (N_25961,N_22466,N_22256);
or U25962 (N_25962,N_22356,N_21767);
and U25963 (N_25963,N_24915,N_22483);
nand U25964 (N_25964,N_23236,N_24330);
or U25965 (N_25965,N_21356,N_23374);
nand U25966 (N_25966,N_24542,N_22638);
or U25967 (N_25967,N_23405,N_23939);
nand U25968 (N_25968,N_21783,N_24006);
or U25969 (N_25969,N_24491,N_21265);
or U25970 (N_25970,N_21766,N_20874);
nand U25971 (N_25971,N_20613,N_20200);
nor U25972 (N_25972,N_21831,N_21730);
nor U25973 (N_25973,N_20561,N_23450);
and U25974 (N_25974,N_21419,N_24479);
and U25975 (N_25975,N_22226,N_21069);
nand U25976 (N_25976,N_20033,N_23925);
or U25977 (N_25977,N_20775,N_21886);
nand U25978 (N_25978,N_21664,N_22935);
and U25979 (N_25979,N_22814,N_22491);
and U25980 (N_25980,N_24101,N_20739);
nor U25981 (N_25981,N_24420,N_21010);
nand U25982 (N_25982,N_21537,N_24892);
or U25983 (N_25983,N_22983,N_23187);
nand U25984 (N_25984,N_22797,N_21452);
and U25985 (N_25985,N_24368,N_21351);
or U25986 (N_25986,N_22821,N_21865);
and U25987 (N_25987,N_23485,N_22080);
xnor U25988 (N_25988,N_24850,N_21271);
and U25989 (N_25989,N_21987,N_24947);
nand U25990 (N_25990,N_24573,N_21510);
nor U25991 (N_25991,N_23688,N_20745);
or U25992 (N_25992,N_23908,N_22215);
and U25993 (N_25993,N_20305,N_23649);
nand U25994 (N_25994,N_24707,N_21579);
nor U25995 (N_25995,N_21268,N_24182);
nand U25996 (N_25996,N_22023,N_24676);
nand U25997 (N_25997,N_23739,N_20478);
nand U25998 (N_25998,N_24951,N_23622);
nor U25999 (N_25999,N_21095,N_22519);
or U26000 (N_26000,N_23230,N_23473);
nand U26001 (N_26001,N_24152,N_24776);
nor U26002 (N_26002,N_23416,N_22223);
and U26003 (N_26003,N_22011,N_23972);
or U26004 (N_26004,N_21575,N_21864);
nor U26005 (N_26005,N_24015,N_21753);
or U26006 (N_26006,N_23209,N_21276);
and U26007 (N_26007,N_20823,N_23095);
nand U26008 (N_26008,N_21047,N_21088);
nor U26009 (N_26009,N_20779,N_22868);
nand U26010 (N_26010,N_24958,N_21366);
nor U26011 (N_26011,N_21572,N_20677);
nand U26012 (N_26012,N_22383,N_20036);
nand U26013 (N_26013,N_22970,N_23989);
nand U26014 (N_26014,N_20096,N_21745);
and U26015 (N_26015,N_21000,N_24055);
nor U26016 (N_26016,N_22327,N_21320);
or U26017 (N_26017,N_20355,N_23136);
nand U26018 (N_26018,N_24606,N_24130);
nor U26019 (N_26019,N_22567,N_21246);
nor U26020 (N_26020,N_20628,N_24319);
nand U26021 (N_26021,N_21157,N_24456);
nand U26022 (N_26022,N_22331,N_22097);
nand U26023 (N_26023,N_23968,N_21033);
nand U26024 (N_26024,N_20952,N_23753);
nor U26025 (N_26025,N_24588,N_23889);
and U26026 (N_26026,N_20635,N_20311);
nor U26027 (N_26027,N_20373,N_20151);
nor U26028 (N_26028,N_20009,N_20511);
nand U26029 (N_26029,N_21434,N_22342);
or U26030 (N_26030,N_22947,N_23734);
nand U26031 (N_26031,N_22959,N_23328);
and U26032 (N_26032,N_22129,N_22122);
and U26033 (N_26033,N_21169,N_21029);
nand U26034 (N_26034,N_22976,N_24635);
nor U26035 (N_26035,N_22172,N_20642);
and U26036 (N_26036,N_24122,N_21454);
and U26037 (N_26037,N_22601,N_22743);
nand U26038 (N_26038,N_23367,N_24068);
or U26039 (N_26039,N_20364,N_23024);
and U26040 (N_26040,N_21533,N_24936);
or U26041 (N_26041,N_23672,N_20698);
nor U26042 (N_26042,N_23998,N_22495);
nor U26043 (N_26043,N_21637,N_22989);
and U26044 (N_26044,N_20907,N_24521);
or U26045 (N_26045,N_24726,N_24024);
nand U26046 (N_26046,N_20651,N_23517);
or U26047 (N_26047,N_23982,N_23022);
nor U26048 (N_26048,N_24168,N_22212);
nor U26049 (N_26049,N_21611,N_22939);
or U26050 (N_26050,N_21608,N_20295);
and U26051 (N_26051,N_21784,N_23194);
nor U26052 (N_26052,N_23694,N_20500);
nand U26053 (N_26053,N_20920,N_24063);
and U26054 (N_26054,N_21591,N_21621);
nor U26055 (N_26055,N_24267,N_23504);
nor U26056 (N_26056,N_23548,N_21493);
or U26057 (N_26057,N_21290,N_23526);
nor U26058 (N_26058,N_23469,N_20587);
nand U26059 (N_26059,N_23633,N_23292);
xor U26060 (N_26060,N_21799,N_21250);
nand U26061 (N_26061,N_22549,N_20935);
and U26062 (N_26062,N_21580,N_24240);
nand U26063 (N_26063,N_22543,N_22399);
nand U26064 (N_26064,N_22156,N_23180);
nand U26065 (N_26065,N_21414,N_23584);
or U26066 (N_26066,N_23383,N_23007);
or U26067 (N_26067,N_23669,N_24155);
nor U26068 (N_26068,N_22833,N_21741);
and U26069 (N_26069,N_22311,N_22029);
or U26070 (N_26070,N_24475,N_24351);
nor U26071 (N_26071,N_21385,N_23413);
or U26072 (N_26072,N_21647,N_21135);
nor U26073 (N_26073,N_24501,N_21565);
nand U26074 (N_26074,N_21312,N_23257);
nand U26075 (N_26075,N_21610,N_23338);
or U26076 (N_26076,N_23502,N_21279);
nand U26077 (N_26077,N_21022,N_20855);
and U26078 (N_26078,N_24490,N_22198);
and U26079 (N_26079,N_22801,N_20884);
or U26080 (N_26080,N_20656,N_23988);
and U26081 (N_26081,N_24905,N_22918);
and U26082 (N_26082,N_22028,N_24146);
nand U26083 (N_26083,N_22487,N_20695);
or U26084 (N_26084,N_23690,N_20810);
nor U26085 (N_26085,N_23824,N_20385);
and U26086 (N_26086,N_24264,N_20636);
and U26087 (N_26087,N_23962,N_22552);
or U26088 (N_26088,N_20923,N_21314);
and U26089 (N_26089,N_20410,N_20805);
nor U26090 (N_26090,N_21412,N_24469);
and U26091 (N_26091,N_22418,N_24530);
and U26092 (N_26092,N_24314,N_24679);
or U26093 (N_26093,N_20606,N_21213);
nand U26094 (N_26094,N_21906,N_23566);
and U26095 (N_26095,N_22588,N_22052);
and U26096 (N_26096,N_21612,N_21085);
or U26097 (N_26097,N_24306,N_23322);
nand U26098 (N_26098,N_22577,N_23111);
and U26099 (N_26099,N_22400,N_20488);
or U26100 (N_26100,N_22363,N_22832);
nor U26101 (N_26101,N_23395,N_21358);
nand U26102 (N_26102,N_20480,N_21847);
or U26103 (N_26103,N_22861,N_20769);
nor U26104 (N_26104,N_24372,N_23161);
or U26105 (N_26105,N_20848,N_22810);
or U26106 (N_26106,N_21406,N_21960);
and U26107 (N_26107,N_20661,N_23503);
nand U26108 (N_26108,N_24863,N_22516);
nor U26109 (N_26109,N_20911,N_24909);
nor U26110 (N_26110,N_20974,N_20242);
or U26111 (N_26111,N_22933,N_21148);
and U26112 (N_26112,N_22545,N_22497);
or U26113 (N_26113,N_24421,N_24765);
and U26114 (N_26114,N_23385,N_22937);
nor U26115 (N_26115,N_23674,N_20392);
nor U26116 (N_26116,N_23006,N_22958);
and U26117 (N_26117,N_24512,N_22809);
nor U26118 (N_26118,N_24586,N_24465);
or U26119 (N_26119,N_23250,N_21733);
and U26120 (N_26120,N_24577,N_24966);
nor U26121 (N_26121,N_22474,N_20206);
nand U26122 (N_26122,N_23811,N_21762);
and U26123 (N_26123,N_23400,N_24065);
nand U26124 (N_26124,N_23031,N_20034);
or U26125 (N_26125,N_22020,N_24322);
or U26126 (N_26126,N_23619,N_24585);
nor U26127 (N_26127,N_23103,N_22837);
xnor U26128 (N_26128,N_23406,N_22353);
nor U26129 (N_26129,N_24774,N_22395);
or U26130 (N_26130,N_20799,N_23789);
and U26131 (N_26131,N_22708,N_22299);
and U26132 (N_26132,N_24142,N_21512);
nand U26133 (N_26133,N_22775,N_20942);
nor U26134 (N_26134,N_22660,N_22825);
or U26135 (N_26135,N_20117,N_24384);
nand U26136 (N_26136,N_20843,N_23311);
nor U26137 (N_26137,N_24430,N_23058);
nor U26138 (N_26138,N_21207,N_20788);
and U26139 (N_26139,N_22729,N_21125);
and U26140 (N_26140,N_20262,N_21727);
nor U26141 (N_26141,N_21142,N_24030);
and U26142 (N_26142,N_22155,N_23192);
nand U26143 (N_26143,N_21594,N_21507);
nand U26144 (N_26144,N_21168,N_21643);
and U26145 (N_26145,N_20691,N_20853);
and U26146 (N_26146,N_21483,N_24519);
nor U26147 (N_26147,N_23425,N_22147);
nor U26148 (N_26148,N_21717,N_20540);
or U26149 (N_26149,N_24407,N_24073);
and U26150 (N_26150,N_24900,N_24448);
and U26151 (N_26151,N_23527,N_20064);
nand U26152 (N_26152,N_22047,N_24580);
and U26153 (N_26153,N_21511,N_22902);
nor U26154 (N_26154,N_20849,N_21494);
nand U26155 (N_26155,N_23762,N_20789);
nand U26156 (N_26156,N_22795,N_23226);
nor U26157 (N_26157,N_21179,N_22337);
nor U26158 (N_26158,N_23806,N_20027);
or U26159 (N_26159,N_24028,N_22093);
or U26160 (N_26160,N_21746,N_24861);
and U26161 (N_26161,N_23140,N_21253);
or U26162 (N_26162,N_22067,N_21680);
and U26163 (N_26163,N_21899,N_24238);
nor U26164 (N_26164,N_21110,N_23264);
or U26165 (N_26165,N_24313,N_24484);
nor U26166 (N_26166,N_20103,N_20666);
nor U26167 (N_26167,N_23843,N_21662);
and U26168 (N_26168,N_24365,N_21578);
and U26169 (N_26169,N_23921,N_21555);
nor U26170 (N_26170,N_23515,N_21172);
and U26171 (N_26171,N_22427,N_23876);
or U26172 (N_26172,N_24798,N_22901);
nand U26173 (N_26173,N_23750,N_20797);
and U26174 (N_26174,N_23658,N_20391);
nor U26175 (N_26175,N_23100,N_23755);
nor U26176 (N_26176,N_20644,N_23821);
nor U26177 (N_26177,N_21040,N_22541);
or U26178 (N_26178,N_24300,N_20520);
or U26179 (N_26179,N_23279,N_22807);
and U26180 (N_26180,N_21842,N_24970);
nor U26181 (N_26181,N_20659,N_23306);
or U26182 (N_26182,N_23010,N_24738);
and U26183 (N_26183,N_21495,N_21496);
nor U26184 (N_26184,N_23686,N_23856);
and U26185 (N_26185,N_20215,N_24446);
or U26186 (N_26186,N_24665,N_23151);
and U26187 (N_26187,N_21205,N_22496);
or U26188 (N_26188,N_21238,N_24311);
or U26189 (N_26189,N_24874,N_22209);
nand U26190 (N_26190,N_23668,N_24154);
and U26191 (N_26191,N_21191,N_24550);
and U26192 (N_26192,N_21947,N_22846);
nor U26193 (N_26193,N_24939,N_23086);
nor U26194 (N_26194,N_22555,N_20501);
nand U26195 (N_26195,N_21897,N_22450);
or U26196 (N_26196,N_22247,N_23756);
and U26197 (N_26197,N_21880,N_24353);
nor U26198 (N_26198,N_23698,N_24254);
nand U26199 (N_26199,N_22500,N_23913);
nand U26200 (N_26200,N_22035,N_20868);
nor U26201 (N_26201,N_22105,N_21935);
nand U26202 (N_26202,N_22724,N_21173);
and U26203 (N_26203,N_21550,N_20168);
or U26204 (N_26204,N_22152,N_20240);
nor U26205 (N_26205,N_20958,N_21843);
or U26206 (N_26206,N_20817,N_23556);
and U26207 (N_26207,N_23769,N_21219);
nand U26208 (N_26208,N_22789,N_24360);
or U26209 (N_26209,N_20436,N_21245);
nor U26210 (N_26210,N_22362,N_22249);
and U26211 (N_26211,N_20199,N_24828);
nor U26212 (N_26212,N_21720,N_23247);
or U26213 (N_26213,N_20097,N_20107);
and U26214 (N_26214,N_20098,N_22565);
nor U26215 (N_26215,N_24321,N_24445);
or U26216 (N_26216,N_23364,N_20552);
or U26217 (N_26217,N_23116,N_24906);
nor U26218 (N_26218,N_23623,N_22728);
or U26219 (N_26219,N_21548,N_23579);
or U26220 (N_26220,N_21491,N_24347);
or U26221 (N_26221,N_23089,N_22946);
or U26222 (N_26222,N_23261,N_21602);
nor U26223 (N_26223,N_24557,N_23955);
and U26224 (N_26224,N_22168,N_24326);
nand U26225 (N_26225,N_21051,N_23214);
and U26226 (N_26226,N_21490,N_22269);
and U26227 (N_26227,N_22927,N_23331);
nor U26228 (N_26228,N_23641,N_20244);
and U26229 (N_26229,N_24834,N_24110);
or U26230 (N_26230,N_23759,N_21119);
nor U26231 (N_26231,N_24873,N_22520);
or U26232 (N_26232,N_24159,N_23333);
and U26233 (N_26233,N_20496,N_23042);
or U26234 (N_26234,N_24724,N_22014);
nor U26235 (N_26235,N_23176,N_21502);
nor U26236 (N_26236,N_24177,N_23075);
nor U26237 (N_26237,N_23016,N_24451);
nand U26238 (N_26238,N_20398,N_20898);
nor U26239 (N_26239,N_20449,N_23014);
nand U26240 (N_26240,N_23162,N_24320);
nor U26241 (N_26241,N_20785,N_22905);
nand U26242 (N_26242,N_23757,N_23975);
and U26243 (N_26243,N_22954,N_20825);
nor U26244 (N_26244,N_24093,N_21686);
nand U26245 (N_26245,N_24350,N_20188);
and U26246 (N_26246,N_23145,N_24843);
and U26247 (N_26247,N_22200,N_24377);
nand U26248 (N_26248,N_21372,N_24730);
and U26249 (N_26249,N_20776,N_23595);
and U26250 (N_26250,N_23356,N_23967);
nand U26251 (N_26251,N_20370,N_20525);
nand U26252 (N_26252,N_22380,N_21957);
nor U26253 (N_26253,N_20195,N_21438);
or U26254 (N_26254,N_21012,N_20904);
and U26255 (N_26255,N_21901,N_21021);
and U26256 (N_26256,N_22191,N_20146);
and U26257 (N_26257,N_24059,N_22951);
or U26258 (N_26258,N_20087,N_20926);
or U26259 (N_26259,N_23970,N_21393);
nand U26260 (N_26260,N_21079,N_21032);
or U26261 (N_26261,N_20014,N_20296);
or U26262 (N_26262,N_21120,N_20366);
nand U26263 (N_26263,N_23277,N_24564);
nor U26264 (N_26264,N_23914,N_22393);
nand U26265 (N_26265,N_21016,N_24375);
nor U26266 (N_26266,N_23745,N_23945);
nor U26267 (N_26267,N_24534,N_21086);
and U26268 (N_26268,N_23567,N_20597);
nand U26269 (N_26269,N_24574,N_22154);
nor U26270 (N_26270,N_20918,N_21787);
nor U26271 (N_26271,N_23030,N_22960);
and U26272 (N_26272,N_21269,N_24962);
and U26273 (N_26273,N_22334,N_24989);
and U26274 (N_26274,N_21928,N_23999);
nand U26275 (N_26275,N_23928,N_21339);
nor U26276 (N_26276,N_23390,N_24785);
or U26277 (N_26277,N_21558,N_22675);
nor U26278 (N_26278,N_24378,N_24921);
or U26279 (N_26279,N_24904,N_20042);
nor U26280 (N_26280,N_21796,N_24749);
and U26281 (N_26281,N_24615,N_21441);
nor U26282 (N_26282,N_20859,N_20320);
or U26283 (N_26283,N_22085,N_22131);
and U26284 (N_26284,N_21693,N_20916);
nor U26285 (N_26285,N_23479,N_21005);
nand U26286 (N_26286,N_21691,N_20057);
or U26287 (N_26287,N_21750,N_24925);
nand U26288 (N_26288,N_21820,N_24515);
nand U26289 (N_26289,N_24119,N_21284);
nand U26290 (N_26290,N_23283,N_20421);
nor U26291 (N_26291,N_22813,N_21984);
nand U26292 (N_26292,N_24624,N_24223);
nand U26293 (N_26293,N_24202,N_22280);
nor U26294 (N_26294,N_20786,N_24598);
nand U26295 (N_26295,N_22308,N_24035);
or U26296 (N_26296,N_24231,N_21267);
and U26297 (N_26297,N_21665,N_20516);
nand U26298 (N_26298,N_21569,N_22826);
or U26299 (N_26299,N_24387,N_21480);
nor U26300 (N_26300,N_23401,N_23565);
and U26301 (N_26301,N_20754,N_20533);
nand U26302 (N_26302,N_20770,N_22319);
nand U26303 (N_26303,N_22346,N_22524);
nor U26304 (N_26304,N_21270,N_20283);
or U26305 (N_26305,N_20185,N_22321);
nor U26306 (N_26306,N_21337,N_20624);
nor U26307 (N_26307,N_20778,N_23020);
and U26308 (N_26308,N_22548,N_22896);
nand U26309 (N_26309,N_24938,N_21952);
or U26310 (N_26310,N_22718,N_21336);
nand U26311 (N_26311,N_24386,N_20647);
nand U26312 (N_26312,N_22103,N_24960);
or U26313 (N_26313,N_24511,N_20161);
nor U26314 (N_26314,N_23940,N_22546);
or U26315 (N_26315,N_23159,N_21795);
and U26316 (N_26316,N_21674,N_22137);
or U26317 (N_26317,N_23523,N_20084);
and U26318 (N_26318,N_24056,N_21241);
nor U26319 (N_26319,N_23884,N_21014);
nand U26320 (N_26320,N_21527,N_20172);
or U26321 (N_26321,N_22853,N_24169);
or U26322 (N_26322,N_22086,N_20318);
nand U26323 (N_26323,N_22998,N_20957);
and U26324 (N_26324,N_24226,N_21499);
nor U26325 (N_26325,N_20551,N_22171);
nor U26326 (N_26326,N_24959,N_23771);
nor U26327 (N_26327,N_22284,N_24131);
and U26328 (N_26328,N_22489,N_22010);
and U26329 (N_26329,N_24536,N_22199);
or U26330 (N_26330,N_20328,N_21981);
and U26331 (N_26331,N_20502,N_21747);
nor U26332 (N_26332,N_21573,N_20359);
nand U26333 (N_26333,N_20846,N_23398);
nor U26334 (N_26334,N_24332,N_23092);
and U26335 (N_26335,N_22526,N_24325);
and U26336 (N_26336,N_21669,N_20062);
and U26337 (N_26337,N_21485,N_20692);
or U26338 (N_26338,N_20987,N_23172);
nor U26339 (N_26339,N_20005,N_24114);
and U26340 (N_26340,N_21500,N_24997);
and U26341 (N_26341,N_24804,N_23845);
or U26342 (N_26342,N_21227,N_22507);
nand U26343 (N_26343,N_20026,N_20030);
and U26344 (N_26344,N_21489,N_21800);
and U26345 (N_26345,N_21476,N_20255);
nand U26346 (N_26346,N_20670,N_22372);
nor U26347 (N_26347,N_20681,N_21251);
and U26348 (N_26348,N_20880,N_23577);
nand U26349 (N_26349,N_20453,N_20687);
nand U26350 (N_26350,N_23775,N_23330);
nand U26351 (N_26351,N_23165,N_24654);
or U26352 (N_26352,N_23594,N_21375);
and U26353 (N_26353,N_20603,N_21154);
and U26354 (N_26354,N_20451,N_24528);
nand U26355 (N_26355,N_20998,N_20091);
and U26356 (N_26356,N_24268,N_23144);
nor U26357 (N_26357,N_23573,N_22298);
nand U26358 (N_26358,N_21416,N_23453);
and U26359 (N_26359,N_21516,N_23842);
nor U26360 (N_26360,N_23791,N_20711);
nand U26361 (N_26361,N_23611,N_24100);
nand U26362 (N_26362,N_21400,N_21126);
nor U26363 (N_26363,N_20622,N_21064);
and U26364 (N_26364,N_23196,N_24258);
or U26365 (N_26365,N_22920,N_20461);
and U26366 (N_26366,N_20564,N_20632);
nor U26367 (N_26367,N_24918,N_23671);
nor U26368 (N_26368,N_21898,N_22069);
or U26369 (N_26369,N_23013,N_20079);
or U26370 (N_26370,N_24481,N_21234);
nor U26371 (N_26371,N_22904,N_23267);
nor U26372 (N_26372,N_23564,N_21343);
and U26373 (N_26373,N_24294,N_24750);
and U26374 (N_26374,N_23084,N_23310);
and U26375 (N_26375,N_24117,N_23435);
nor U26376 (N_26376,N_23445,N_21352);
nand U26377 (N_26377,N_21931,N_20554);
or U26378 (N_26378,N_21632,N_24934);
and U26379 (N_26379,N_24343,N_21160);
and U26380 (N_26380,N_20351,N_22158);
and U26381 (N_26381,N_20784,N_21141);
or U26382 (N_26382,N_24273,N_20214);
and U26383 (N_26383,N_20094,N_23454);
and U26384 (N_26384,N_21275,N_21567);
or U26385 (N_26385,N_23643,N_23129);
and U26386 (N_26386,N_24964,N_23064);
xnor U26387 (N_26387,N_22605,N_21841);
and U26388 (N_26388,N_23113,N_22684);
nor U26389 (N_26389,N_24509,N_22077);
and U26390 (N_26390,N_21967,N_21212);
or U26391 (N_26391,N_21530,N_23973);
nor U26392 (N_26392,N_24057,N_24617);
nor U26393 (N_26393,N_24996,N_21884);
or U26394 (N_26394,N_24686,N_20139);
and U26395 (N_26395,N_21853,N_24786);
or U26396 (N_26396,N_24403,N_23273);
or U26397 (N_26397,N_24825,N_21523);
or U26398 (N_26398,N_20790,N_21909);
nand U26399 (N_26399,N_21055,N_20484);
nor U26400 (N_26400,N_20086,N_24994);
nand U26401 (N_26401,N_21539,N_22242);
and U26402 (N_26402,N_24552,N_22316);
nand U26403 (N_26403,N_22323,N_23411);
and U26404 (N_26404,N_21815,N_22768);
nand U26405 (N_26405,N_22159,N_21323);
and U26406 (N_26406,N_21636,N_21003);
and U26407 (N_26407,N_24572,N_22736);
nand U26408 (N_26408,N_21389,N_22213);
nand U26409 (N_26409,N_21959,N_22492);
nand U26410 (N_26410,N_21099,N_20018);
and U26411 (N_26411,N_24171,N_21018);
nor U26412 (N_26412,N_23772,N_21938);
and U26413 (N_26413,N_21379,N_24813);
or U26414 (N_26414,N_22089,N_24090);
and U26415 (N_26415,N_23896,N_22749);
and U26416 (N_26416,N_22531,N_22568);
nor U26417 (N_26417,N_20389,N_20565);
nor U26418 (N_26418,N_23715,N_21562);
or U26419 (N_26419,N_23948,N_23156);
or U26420 (N_26420,N_22625,N_24221);
nand U26421 (N_26421,N_20572,N_20649);
nor U26422 (N_26422,N_20906,N_22338);
or U26423 (N_26423,N_20444,N_24303);
or U26424 (N_26424,N_22175,N_22856);
nor U26425 (N_26425,N_21255,N_20399);
nor U26426 (N_26426,N_22218,N_21239);
or U26427 (N_26427,N_20625,N_23586);
or U26428 (N_26428,N_21471,N_23085);
or U26429 (N_26429,N_23441,N_24884);
nand U26430 (N_26430,N_23705,N_22644);
or U26431 (N_26431,N_23630,N_21652);
nor U26432 (N_26432,N_22748,N_21020);
nand U26433 (N_26433,N_20273,N_22838);
or U26434 (N_26434,N_24592,N_20820);
and U26435 (N_26435,N_20189,N_21916);
nand U26436 (N_26436,N_23554,N_24214);
nor U26437 (N_26437,N_20963,N_24380);
nand U26438 (N_26438,N_21488,N_20381);
nand U26439 (N_26439,N_24477,N_24699);
nand U26440 (N_26440,N_24535,N_20594);
or U26441 (N_26441,N_20734,N_22470);
and U26442 (N_26442,N_20646,N_20136);
and U26443 (N_26443,N_22091,N_21204);
nand U26444 (N_26444,N_21202,N_22250);
or U26445 (N_26445,N_23440,N_22031);
or U26446 (N_26446,N_21892,N_24604);
and U26447 (N_26447,N_21367,N_20462);
nand U26448 (N_26448,N_24547,N_24851);
nor U26449 (N_26449,N_20575,N_24089);
and U26450 (N_26450,N_22015,N_20867);
or U26451 (N_26451,N_20137,N_23926);
xnor U26452 (N_26452,N_21365,N_22551);
or U26453 (N_26453,N_22361,N_22656);
nor U26454 (N_26454,N_20660,N_20465);
and U26455 (N_26455,N_20101,N_24003);
nor U26456 (N_26456,N_21764,N_24844);
or U26457 (N_26457,N_20583,N_22952);
xor U26458 (N_26458,N_21722,N_21571);
nor U26459 (N_26459,N_24719,N_20207);
and U26460 (N_26460,N_23354,N_21193);
nor U26461 (N_26461,N_20940,N_21792);
nor U26462 (N_26462,N_20777,N_24060);
and U26463 (N_26463,N_23981,N_21254);
nand U26464 (N_26464,N_23543,N_20259);
nand U26465 (N_26465,N_22897,N_24399);
xnor U26466 (N_26466,N_23478,N_24438);
or U26467 (N_26467,N_22357,N_24118);
or U26468 (N_26468,N_20216,N_20294);
nand U26469 (N_26469,N_24903,N_22574);
or U26470 (N_26470,N_23133,N_20723);
and U26471 (N_26471,N_22686,N_24973);
and U26472 (N_26472,N_21509,N_23909);
and U26473 (N_26473,N_20387,N_20483);
nand U26474 (N_26474,N_24183,N_23472);
nor U26475 (N_26475,N_24176,N_21776);
and U26476 (N_26476,N_20618,N_24298);
nand U26477 (N_26477,N_23091,N_22892);
nor U26478 (N_26478,N_22178,N_22076);
nor U26479 (N_26479,N_23021,N_24012);
nor U26480 (N_26480,N_22355,N_21710);
nor U26481 (N_26481,N_22737,N_22286);
xor U26482 (N_26482,N_21879,N_24051);
or U26483 (N_26483,N_20229,N_22278);
nand U26484 (N_26484,N_22870,N_23585);
nand U26485 (N_26485,N_22376,N_22375);
or U26486 (N_26486,N_21185,N_21704);
or U26487 (N_26487,N_20903,N_20556);
and U26488 (N_26488,N_24722,N_21729);
nand U26489 (N_26489,N_20252,N_24929);
and U26490 (N_26490,N_24428,N_20752);
and U26491 (N_26491,N_20247,N_24634);
nand U26492 (N_26492,N_22673,N_21896);
nand U26493 (N_26493,N_20268,N_23248);
nor U26494 (N_26494,N_24396,N_23061);
nand U26495 (N_26495,N_22857,N_24354);
nand U26496 (N_26496,N_21606,N_22618);
nand U26497 (N_26497,N_22001,N_23521);
and U26498 (N_26498,N_23574,N_23071);
nand U26499 (N_26499,N_24087,N_22114);
nand U26500 (N_26500,N_21313,N_20943);
nand U26501 (N_26501,N_24910,N_24729);
nor U26502 (N_26502,N_21360,N_23078);
nor U26503 (N_26503,N_24894,N_22637);
and U26504 (N_26504,N_23396,N_20973);
nor U26505 (N_26505,N_23054,N_21951);
xnor U26506 (N_26506,N_20124,N_22992);
nand U26507 (N_26507,N_20165,N_22289);
nand U26508 (N_26508,N_20505,N_23067);
nand U26509 (N_26509,N_23362,N_20811);
or U26510 (N_26510,N_22566,N_24922);
nand U26511 (N_26511,N_20166,N_24985);
and U26512 (N_26512,N_22662,N_22292);
nor U26513 (N_26513,N_22405,N_22365);
nand U26514 (N_26514,N_24235,N_24014);
nor U26515 (N_26515,N_23692,N_23391);
and U26516 (N_26516,N_22096,N_21435);
or U26517 (N_26517,N_24299,N_23916);
nand U26518 (N_26518,N_23342,N_22505);
or U26519 (N_26519,N_23597,N_22777);
nand U26520 (N_26520,N_23514,N_23839);
and U26521 (N_26521,N_23953,N_20524);
nor U26522 (N_26522,N_20341,N_24474);
nand U26523 (N_26523,N_20315,N_21429);
or U26524 (N_26524,N_24928,N_24078);
nand U26525 (N_26525,N_22862,N_21442);
and U26526 (N_26526,N_23902,N_21751);
nand U26527 (N_26527,N_24251,N_21073);
or U26528 (N_26528,N_24295,N_20314);
nor U26529 (N_26529,N_21737,N_23786);
nand U26530 (N_26530,N_20832,N_22750);
or U26531 (N_26531,N_20187,N_21092);
or U26532 (N_26532,N_23349,N_24579);
or U26533 (N_26533,N_21371,N_20052);
nor U26534 (N_26534,N_20440,N_24196);
or U26535 (N_26535,N_20411,N_21657);
and U26536 (N_26536,N_23017,N_21581);
nor U26537 (N_26537,N_22943,N_21420);
or U26538 (N_26538,N_23702,N_22903);
xor U26539 (N_26539,N_23693,N_24279);
nand U26540 (N_26540,N_20059,N_23246);
nor U26541 (N_26541,N_23898,N_20591);
or U26542 (N_26542,N_24787,N_24640);
nor U26543 (N_26543,N_24255,N_24382);
nand U26544 (N_26544,N_21437,N_23249);
or U26545 (N_26545,N_22963,N_24668);
nand U26546 (N_26546,N_21570,N_20031);
or U26547 (N_26547,N_20930,N_20497);
nor U26548 (N_26548,N_21788,N_21348);
and U26549 (N_26549,N_24359,N_20685);
or U26550 (N_26550,N_20980,N_20433);
nor U26551 (N_26551,N_22766,N_22921);
nand U26552 (N_26552,N_20337,N_22561);
nand U26553 (N_26553,N_21742,N_20550);
nor U26554 (N_26554,N_24290,N_23798);
nor U26555 (N_26555,N_23218,N_21378);
nand U26556 (N_26556,N_21057,N_22016);
nand U26557 (N_26557,N_20266,N_24106);
nor U26558 (N_26558,N_23829,N_22326);
and U26559 (N_26559,N_22649,N_22404);
nor U26560 (N_26560,N_24882,N_20623);
nor U26561 (N_26561,N_20655,N_23638);
and U26562 (N_26562,N_21939,N_20744);
nor U26563 (N_26563,N_22202,N_20000);
nor U26564 (N_26564,N_21645,N_24619);
or U26565 (N_26565,N_23697,N_22745);
nand U26566 (N_26566,N_21780,N_21399);
or U26567 (N_26567,N_21431,N_24005);
or U26568 (N_26568,N_24902,N_21851);
nand U26569 (N_26569,N_21349,N_24361);
nand U26570 (N_26570,N_20515,N_21134);
nand U26571 (N_26571,N_20414,N_24197);
nand U26572 (N_26572,N_24871,N_21041);
and U26573 (N_26573,N_23231,N_21448);
nor U26574 (N_26574,N_21237,N_22785);
and U26575 (N_26575,N_24459,N_20129);
nor U26576 (N_26576,N_24188,N_23271);
or U26577 (N_26577,N_23317,N_23270);
nand U26578 (N_26578,N_22169,N_23785);
nor U26579 (N_26579,N_24261,N_24138);
nand U26580 (N_26580,N_21585,N_20131);
or U26581 (N_26581,N_23179,N_22798);
or U26582 (N_26582,N_24754,N_22532);
or U26583 (N_26583,N_24933,N_24436);
nand U26584 (N_26584,N_22396,N_23770);
nand U26585 (N_26585,N_22646,N_24715);
and U26586 (N_26586,N_22081,N_21087);
or U26587 (N_26587,N_24853,N_23384);
or U26588 (N_26588,N_23991,N_22036);
nor U26589 (N_26589,N_22974,N_21383);
and U26590 (N_26590,N_23431,N_22586);
or U26591 (N_26591,N_22449,N_23204);
and U26592 (N_26592,N_24433,N_21650);
and U26593 (N_26593,N_22232,N_21903);
and U26594 (N_26594,N_20333,N_21520);
nand U26595 (N_26595,N_21703,N_22848);
or U26596 (N_26596,N_21105,N_21677);
or U26597 (N_26597,N_23553,N_22271);
nor U26598 (N_26598,N_22990,N_22348);
or U26599 (N_26599,N_24674,N_23942);
nor U26600 (N_26600,N_24688,N_24362);
and U26601 (N_26601,N_24854,N_23291);
or U26602 (N_26602,N_20158,N_24662);
and U26603 (N_26603,N_22476,N_22886);
nand U26604 (N_26604,N_21519,N_21122);
nand U26605 (N_26605,N_22622,N_24071);
nor U26606 (N_26606,N_20969,N_24808);
nor U26607 (N_26607,N_20275,N_21364);
and U26608 (N_26608,N_23546,N_23978);
or U26609 (N_26609,N_20557,N_20961);
nor U26610 (N_26610,N_21098,N_24761);
or U26611 (N_26611,N_21744,N_24838);
and U26612 (N_26612,N_22434,N_21832);
nor U26613 (N_26613,N_21778,N_24741);
nor U26614 (N_26614,N_22941,N_23969);
nand U26615 (N_26615,N_20796,N_22367);
and U26616 (N_26616,N_20225,N_21192);
nor U26617 (N_26617,N_21673,N_23421);
or U26618 (N_26618,N_20917,N_22183);
or U26619 (N_26619,N_20159,N_20756);
nand U26620 (N_26620,N_23325,N_23286);
nand U26621 (N_26621,N_24334,N_23446);
or U26622 (N_26622,N_21460,N_23984);
and U26623 (N_26623,N_20804,N_23820);
or U26624 (N_26624,N_21623,N_22806);
nand U26625 (N_26625,N_20021,N_24709);
nand U26626 (N_26626,N_22934,N_21128);
or U26627 (N_26627,N_23696,N_23763);
or U26628 (N_26628,N_23234,N_23074);
and U26629 (N_26629,N_20099,N_24778);
nor U26630 (N_26630,N_21283,N_21107);
and U26631 (N_26631,N_21200,N_23714);
and U26632 (N_26632,N_20024,N_23895);
and U26633 (N_26633,N_22579,N_24393);
and U26634 (N_26634,N_24755,N_22503);
or U26635 (N_26635,N_21588,N_22397);
and U26636 (N_26636,N_23680,N_20971);
or U26637 (N_26637,N_24216,N_20092);
nor U26638 (N_26638,N_21811,N_24422);
or U26639 (N_26639,N_23272,N_20888);
nand U26640 (N_26640,N_23352,N_20539);
and U26641 (N_26641,N_21342,N_22630);
nand U26642 (N_26642,N_21706,N_24549);
and U26643 (N_26643,N_20800,N_20694);
nand U26644 (N_26644,N_24356,N_21455);
and U26645 (N_26645,N_23666,N_23190);
or U26646 (N_26646,N_22613,N_20673);
nand U26647 (N_26647,N_24472,N_22712);
nor U26648 (N_26648,N_23002,N_23508);
nand U26649 (N_26649,N_21785,N_24570);
nor U26650 (N_26650,N_20409,N_23203);
or U26651 (N_26651,N_24022,N_23223);
nand U26652 (N_26652,N_23860,N_20544);
nand U26653 (N_26653,N_24648,N_22783);
nor U26654 (N_26654,N_21943,N_23051);
and U26655 (N_26655,N_20726,N_22255);
or U26656 (N_26656,N_21700,N_21402);
and U26657 (N_26657,N_20495,N_21478);
nor U26658 (N_26658,N_24253,N_21215);
or U26659 (N_26659,N_22472,N_21689);
nand U26660 (N_26660,N_23648,N_23287);
nor U26661 (N_26661,N_20443,N_23716);
nand U26662 (N_26662,N_23899,N_22774);
nand U26663 (N_26663,N_23591,N_22792);
nand U26664 (N_26664,N_20576,N_20891);
or U26665 (N_26665,N_24185,N_22157);
or U26666 (N_26666,N_23447,N_21604);
nor U26667 (N_26667,N_23652,N_23200);
nor U26668 (N_26668,N_21413,N_21469);
and U26669 (N_26669,N_24626,N_22620);
nand U26670 (N_26670,N_21995,N_22571);
or U26671 (N_26671,N_20700,N_21824);
nor U26672 (N_26672,N_23149,N_21067);
and U26673 (N_26673,N_21598,N_20757);
and U26674 (N_26674,N_24457,N_21054);
and U26675 (N_26675,N_20153,N_20966);
and U26676 (N_26676,N_22402,N_24663);
nand U26677 (N_26677,N_24513,N_22125);
nor U26678 (N_26678,N_21631,N_21292);
nand U26679 (N_26679,N_24569,N_20750);
nand U26680 (N_26680,N_22540,N_22349);
nand U26681 (N_26681,N_21103,N_22898);
or U26682 (N_26682,N_21013,N_23379);
or U26683 (N_26683,N_22455,N_20446);
nor U26684 (N_26684,N_24991,N_20217);
nor U26685 (N_26685,N_21859,N_24346);
xor U26686 (N_26686,N_23019,N_24132);
nor U26687 (N_26687,N_24363,N_23799);
nand U26688 (N_26688,N_24708,N_20415);
and U26689 (N_26689,N_20995,N_20249);
or U26690 (N_26690,N_22272,N_20878);
or U26691 (N_26691,N_20947,N_23732);
nand U26692 (N_26692,N_23358,N_23533);
nand U26693 (N_26693,N_24204,N_21878);
and U26694 (N_26694,N_22189,N_21620);
or U26695 (N_26695,N_24208,N_20901);
nor U26696 (N_26696,N_20802,N_23307);
or U26697 (N_26697,N_24207,N_21635);
nor U26698 (N_26698,N_23875,N_22881);
or U26699 (N_26699,N_20081,N_24398);
or U26700 (N_26700,N_23282,N_20167);
and U26701 (N_26701,N_20424,N_20895);
nand U26702 (N_26702,N_22647,N_23794);
or U26703 (N_26703,N_23803,N_20448);
or U26704 (N_26704,N_22008,N_21116);
nand U26705 (N_26705,N_23890,N_22366);
and U26706 (N_26706,N_24054,N_24886);
or U26707 (N_26707,N_21257,N_20830);
and U26708 (N_26708,N_24681,N_24760);
nand U26709 (N_26709,N_23810,N_24868);
nor U26710 (N_26710,N_20489,N_23736);
or U26711 (N_26711,N_20090,N_22195);
nor U26712 (N_26712,N_21592,N_24336);
or U26713 (N_26713,N_22445,N_24263);
nor U26714 (N_26714,N_20748,N_23174);
nand U26715 (N_26715,N_20432,N_22006);
and U26716 (N_26716,N_21538,N_21807);
nand U26717 (N_26717,N_24744,N_24104);
nand U26718 (N_26718,N_21912,N_21334);
nor U26719 (N_26719,N_22261,N_24233);
nand U26720 (N_26720,N_24293,N_21326);
or U26721 (N_26721,N_22448,N_22486);
nand U26722 (N_26722,N_22439,N_21178);
nand U26723 (N_26723,N_23475,N_20066);
nand U26724 (N_26724,N_21006,N_21817);
and U26725 (N_26725,N_21821,N_21660);
and U26726 (N_26726,N_22761,N_20553);
nand U26727 (N_26727,N_24092,N_20737);
or U26728 (N_26728,N_23682,N_20076);
nor U26729 (N_26729,N_24483,N_23428);
and U26730 (N_26730,N_21285,N_22238);
nor U26731 (N_26731,N_20063,N_23525);
and U26732 (N_26732,N_22980,N_23997);
nand U26733 (N_26733,N_21081,N_23171);
and U26734 (N_26734,N_22415,N_22790);
nand U26735 (N_26735,N_24671,N_24728);
nor U26736 (N_26736,N_23520,N_22710);
and U26737 (N_26737,N_21002,N_22916);
or U26738 (N_26738,N_20959,N_24782);
and U26739 (N_26739,N_20645,N_22274);
or U26740 (N_26740,N_20186,N_20509);
or U26741 (N_26741,N_23386,N_23721);
and U26742 (N_26742,N_24666,N_24419);
nor U26743 (N_26743,N_21295,N_20253);
or U26744 (N_26744,N_24249,N_24000);
nand U26745 (N_26745,N_23001,N_24865);
or U26746 (N_26746,N_24687,N_21911);
and U26747 (N_26747,N_21232,N_24794);
nor U26748 (N_26748,N_24029,N_23571);
and U26749 (N_26749,N_20491,N_20872);
nand U26750 (N_26750,N_20234,N_22177);
or U26751 (N_26751,N_21950,N_24315);
and U26752 (N_26752,N_21524,N_20950);
nor U26753 (N_26753,N_21325,N_24913);
nand U26754 (N_26754,N_24661,N_23532);
and U26755 (N_26755,N_24602,N_22596);
and U26756 (N_26756,N_20279,N_20162);
nand U26757 (N_26757,N_24878,N_22050);
xnor U26758 (N_26758,N_20922,N_23854);
or U26759 (N_26759,N_21989,N_24770);
nor U26760 (N_26760,N_22251,N_23812);
or U26761 (N_26761,N_23737,N_20025);
and U26762 (N_26762,N_21462,N_24408);
nor U26763 (N_26763,N_20276,N_20909);
or U26764 (N_26764,N_22895,N_24734);
or U26765 (N_26765,N_23779,N_24614);
nand U26766 (N_26766,N_20818,N_24963);
nand U26767 (N_26767,N_22398,N_21208);
nand U26768 (N_26768,N_20577,N_20835);
and U26769 (N_26769,N_20758,N_22711);
nor U26770 (N_26770,N_24780,N_24394);
xnor U26771 (N_26771,N_22241,N_24824);
nand U26772 (N_26772,N_24217,N_23874);
and U26773 (N_26773,N_22911,N_23894);
nor U26774 (N_26774,N_24524,N_20003);
nor U26775 (N_26775,N_20307,N_23783);
and U26776 (N_26776,N_24680,N_24956);
nand U26777 (N_26777,N_22041,N_20405);
nand U26778 (N_26778,N_23184,N_23985);
nor U26779 (N_26779,N_22205,N_23215);
nand U26780 (N_26780,N_23350,N_21958);
or U26781 (N_26781,N_22406,N_20992);
nand U26782 (N_26782,N_22300,N_22442);
and U26783 (N_26783,N_20144,N_22658);
nand U26784 (N_26784,N_22852,N_24172);
nand U26785 (N_26785,N_24522,N_24495);
and U26786 (N_26786,N_24593,N_22377);
and U26787 (N_26787,N_22595,N_20905);
or U26788 (N_26788,N_21278,N_21649);
nand U26789 (N_26789,N_20028,N_22370);
xor U26790 (N_26790,N_23464,N_22584);
or U26791 (N_26791,N_23237,N_23041);
and U26792 (N_26792,N_22461,N_22842);
and U26793 (N_26793,N_23861,N_20599);
and U26794 (N_26794,N_22444,N_23568);
nor U26795 (N_26795,N_24307,N_21026);
or U26796 (N_26796,N_21887,N_21740);
nand U26797 (N_26797,N_23206,N_24870);
or U26798 (N_26798,N_23228,N_20082);
nand U26799 (N_26799,N_21856,N_24737);
nor U26800 (N_26800,N_23582,N_23045);
and U26801 (N_26801,N_24908,N_23629);
or U26802 (N_26802,N_23768,N_21236);
nand U26803 (N_26803,N_22408,N_21373);
and U26804 (N_26804,N_20045,N_21335);
or U26805 (N_26805,N_24464,N_21228);
or U26806 (N_26806,N_23420,N_24199);
nand U26807 (N_26807,N_24140,N_24802);
nor U26808 (N_26808,N_20860,N_23152);
nand U26809 (N_26809,N_21396,N_24021);
and U26810 (N_26810,N_20212,N_24553);
nand U26811 (N_26811,N_24367,N_20140);
nor U26812 (N_26812,N_23529,N_23625);
nand U26813 (N_26813,N_20795,N_22358);
or U26814 (N_26814,N_23869,N_20017);
and U26815 (N_26815,N_23624,N_21230);
or U26816 (N_26816,N_24645,N_23563);
nor U26817 (N_26817,N_21422,N_21397);
nor U26818 (N_26818,N_23626,N_23603);
or U26819 (N_26819,N_24205,N_21827);
nand U26820 (N_26820,N_24082,N_24133);
or U26821 (N_26821,N_23911,N_24847);
nor U26822 (N_26822,N_20858,N_21123);
and U26823 (N_26823,N_21180,N_20049);
and U26824 (N_26824,N_24795,N_21556);
or U26825 (N_26825,N_24262,N_20727);
or U26826 (N_26826,N_22181,N_20472);
and U26827 (N_26827,N_22138,N_20639);
nand U26828 (N_26828,N_20765,N_21514);
and U26829 (N_26829,N_20067,N_22464);
or U26830 (N_26830,N_20567,N_24058);
and U26831 (N_26831,N_24161,N_23538);
and U26832 (N_26832,N_22908,N_21197);
nand U26833 (N_26833,N_23831,N_20102);
nor U26834 (N_26834,N_23253,N_23132);
and U26835 (N_26835,N_23484,N_21024);
nor U26836 (N_26836,N_21628,N_21261);
nand U26837 (N_26837,N_20932,N_24831);
nor U26838 (N_26838,N_22336,N_24333);
nor U26839 (N_26839,N_22170,N_21736);
or U26840 (N_26840,N_24948,N_22239);
and U26841 (N_26841,N_21274,N_23570);
or U26842 (N_26842,N_21165,N_22544);
or U26843 (N_26843,N_23607,N_22373);
or U26844 (N_26844,N_20841,N_23679);
nand U26845 (N_26845,N_21837,N_24757);
or U26846 (N_26846,N_20760,N_22780);
and U26847 (N_26847,N_20407,N_22854);
and U26848 (N_26848,N_20278,N_23480);
nor U26849 (N_26849,N_21317,N_22688);
or U26850 (N_26850,N_22872,N_22703);
and U26851 (N_26851,N_23793,N_22467);
and U26852 (N_26852,N_21094,N_20335);
and U26853 (N_26853,N_20740,N_23651);
nor U26854 (N_26854,N_22995,N_22917);
and U26855 (N_26855,N_23946,N_23706);
nand U26856 (N_26856,N_23394,N_24352);
or U26857 (N_26857,N_20050,N_23731);
nor U26858 (N_26858,N_22435,N_23852);
nor U26859 (N_26859,N_22320,N_21058);
nand U26860 (N_26860,N_22322,N_20248);
nand U26861 (N_26861,N_24234,N_20069);
nand U26862 (N_26862,N_24673,N_21405);
and U26863 (N_26863,N_24701,N_22317);
nand U26864 (N_26864,N_21266,N_21390);
and U26865 (N_26865,N_24209,N_22118);
nand U26866 (N_26866,N_23028,N_23562);
nor U26867 (N_26867,N_24775,N_21754);
nand U26868 (N_26868,N_23302,N_23044);
or U26869 (N_26869,N_23429,N_22193);
and U26870 (N_26870,N_20733,N_23487);
and U26871 (N_26871,N_24628,N_22228);
nor U26872 (N_26872,N_22778,N_20264);
or U26873 (N_26873,N_24769,N_22420);
nor U26874 (N_26874,N_21470,N_22746);
nand U26875 (N_26875,N_24632,N_20657);
nor U26876 (N_26876,N_22643,N_20447);
nand U26877 (N_26877,N_21781,N_22108);
nor U26878 (N_26878,N_24603,N_22621);
and U26879 (N_26879,N_22804,N_23778);
or U26880 (N_26880,N_22281,N_20637);
nor U26881 (N_26881,N_20793,N_21080);
nor U26882 (N_26882,N_22374,N_23025);
or U26883 (N_26883,N_23337,N_24582);
xnor U26884 (N_26884,N_22051,N_22460);
nor U26885 (N_26885,N_21839,N_20114);
or U26886 (N_26886,N_20807,N_24020);
or U26887 (N_26887,N_20476,N_20470);
and U26888 (N_26888,N_22344,N_24695);
nor U26889 (N_26889,N_20751,N_22784);
nand U26890 (N_26890,N_24945,N_23609);
nor U26891 (N_26891,N_21302,N_23141);
or U26892 (N_26892,N_22866,N_22779);
nand U26893 (N_26893,N_21297,N_21001);
nand U26894 (N_26894,N_24174,N_23488);
nor U26895 (N_26895,N_22615,N_22032);
or U26896 (N_26896,N_23830,N_24473);
or U26897 (N_26897,N_20725,N_20384);
and U26898 (N_26898,N_24982,N_23188);
nor U26899 (N_26899,N_22312,N_22844);
nand U26900 (N_26900,N_20221,N_22765);
and U26901 (N_26901,N_20571,N_22481);
and U26902 (N_26902,N_23544,N_24476);
nand U26903 (N_26903,N_21201,N_22477);
nand U26904 (N_26904,N_23235,N_22986);
and U26905 (N_26905,N_22260,N_24256);
or U26906 (N_26906,N_22730,N_23826);
nand U26907 (N_26907,N_23389,N_23906);
or U26908 (N_26908,N_20231,N_22556);
or U26909 (N_26909,N_20665,N_23838);
nand U26910 (N_26910,N_24410,N_23927);
nand U26911 (N_26911,N_22949,N_21934);
and U26912 (N_26912,N_22919,N_21338);
nand U26913 (N_26913,N_22681,N_20043);
nand U26914 (N_26914,N_20116,N_24533);
or U26915 (N_26915,N_23351,N_23068);
nor U26916 (N_26916,N_21083,N_22116);
and U26917 (N_26917,N_22064,N_20301);
nor U26918 (N_26918,N_21248,N_21683);
nor U26919 (N_26919,N_22878,N_21321);
nor U26920 (N_26920,N_21862,N_21992);
or U26921 (N_26921,N_21112,N_24995);
or U26922 (N_26922,N_21075,N_24969);
and U26923 (N_26923,N_23205,N_24703);
nand U26924 (N_26924,N_23583,N_23491);
or U26925 (N_26925,N_20299,N_21369);
or U26926 (N_26926,N_21919,N_20245);
nand U26927 (N_26927,N_24539,N_23879);
or U26928 (N_26928,N_21964,N_22058);
nand U26929 (N_26929,N_21143,N_20809);
or U26930 (N_26930,N_24357,N_23613);
nor U26931 (N_26931,N_20482,N_23468);
xnor U26932 (N_26932,N_23265,N_22836);
or U26933 (N_26933,N_24783,N_24682);
nand U26934 (N_26934,N_21596,N_20368);
or U26935 (N_26935,N_20896,N_21355);
nand U26936 (N_26936,N_23087,N_24883);
nor U26937 (N_26937,N_21465,N_23918);
nand U26938 (N_26938,N_24823,N_23498);
nor U26939 (N_26939,N_22185,N_21944);
nand U26940 (N_26940,N_22925,N_23979);
xnor U26941 (N_26941,N_24212,N_22819);
and U26942 (N_26942,N_22914,N_20218);
and U26943 (N_26943,N_24485,N_21049);
nor U26944 (N_26944,N_21133,N_24243);
nor U26945 (N_26945,N_20239,N_22107);
nand U26946 (N_26946,N_24935,N_23097);
or U26947 (N_26947,N_22479,N_22094);
nor U26948 (N_26948,N_22581,N_21417);
or U26949 (N_26949,N_23460,N_21501);
nor U26950 (N_26950,N_23849,N_20223);
nand U26951 (N_26951,N_21506,N_23951);
nand U26952 (N_26952,N_24869,N_21690);
nand U26953 (N_26953,N_24283,N_23418);
xnor U26954 (N_26954,N_20701,N_21456);
nand U26955 (N_26955,N_21638,N_23169);
nor U26956 (N_26956,N_20720,N_20939);
nor U26957 (N_26957,N_24968,N_24896);
or U26958 (N_26958,N_21104,N_20319);
nor U26959 (N_26959,N_20829,N_20982);
nor U26960 (N_26960,N_22100,N_21564);
or U26961 (N_26961,N_24499,N_20357);
or U26962 (N_26962,N_24548,N_24265);
nand U26963 (N_26963,N_20664,N_21158);
or U26964 (N_26964,N_24563,N_20371);
or U26965 (N_26965,N_22640,N_24200);
nand U26966 (N_26966,N_22165,N_21642);
or U26967 (N_26967,N_24596,N_22664);
nor U26968 (N_26968,N_22005,N_22429);
nand U26969 (N_26969,N_22352,N_21597);
nor U26970 (N_26970,N_21937,N_22394);
nor U26971 (N_26971,N_23851,N_21812);
nand U26972 (N_26972,N_20837,N_24269);
nor U26973 (N_26973,N_23760,N_24520);
and U26974 (N_26974,N_20771,N_20345);
or U26975 (N_26975,N_24287,N_23800);
nor U26976 (N_26976,N_22831,N_21291);
nand U26977 (N_26977,N_22385,N_21037);
nor U26978 (N_26978,N_21793,N_22121);
nand U26979 (N_26979,N_24252,N_24608);
nor U26980 (N_26980,N_24496,N_24889);
nand U26981 (N_26981,N_21961,N_22674);
nand U26982 (N_26982,N_20626,N_22929);
nand U26983 (N_26983,N_21203,N_23329);
and U26984 (N_26984,N_21209,N_21773);
or U26985 (N_26985,N_20894,N_21774);
nor U26986 (N_26986,N_20233,N_22265);
and U26987 (N_26987,N_20293,N_20250);
nand U26988 (N_26988,N_24206,N_22591);
nand U26989 (N_26989,N_21890,N_20360);
and U26990 (N_26990,N_23360,N_20964);
nor U26991 (N_26991,N_21391,N_20753);
nand U26992 (N_26992,N_23684,N_24576);
and U26993 (N_26993,N_23128,N_22965);
nor U26994 (N_26994,N_24565,N_22747);
and U26995 (N_26995,N_24424,N_22950);
or U26996 (N_26996,N_21461,N_23788);
nor U26997 (N_26997,N_20538,N_21616);
xor U26998 (N_26998,N_24219,N_21927);
and U26999 (N_26999,N_22379,N_22521);
nand U27000 (N_27000,N_20689,N_20298);
and U27001 (N_27001,N_23229,N_23081);
nor U27002 (N_27002,N_23976,N_22235);
and U27003 (N_27003,N_20621,N_21036);
xor U27004 (N_27004,N_24061,N_21106);
nand U27005 (N_27005,N_20013,N_22148);
nor U27006 (N_27006,N_24095,N_21991);
nor U27007 (N_27007,N_22863,N_24578);
nor U27008 (N_27008,N_20326,N_21804);
xnor U27009 (N_27009,N_23463,N_23088);
or U27010 (N_27010,N_24025,N_23796);
nand U27011 (N_27011,N_24685,N_24971);
or U27012 (N_27012,N_21761,N_22955);
nor U27013 (N_27013,N_21918,N_20193);
nand U27014 (N_27014,N_20061,N_23689);
nor U27015 (N_27015,N_22592,N_23220);
or U27016 (N_27016,N_22130,N_24720);
nand U27017 (N_27017,N_23336,N_22670);
nor U27018 (N_27018,N_24712,N_22858);
and U27019 (N_27019,N_22440,N_21272);
nor U27020 (N_27020,N_22987,N_22629);
and U27021 (N_27021,N_23219,N_24745);
and U27022 (N_27022,N_20093,N_23499);
or U27023 (N_27023,N_22594,N_21281);
and U27024 (N_27024,N_21994,N_21535);
nand U27025 (N_27025,N_24441,N_23929);
nand U27026 (N_27026,N_23923,N_23605);
nand U27027 (N_27027,N_22279,N_24827);
nor U27028 (N_27028,N_20015,N_20304);
nor U27029 (N_27029,N_20581,N_22865);
nand U27030 (N_27030,N_21408,N_21436);
xnor U27031 (N_27031,N_23199,N_22416);
nor U27032 (N_27032,N_21357,N_22938);
or U27033 (N_27033,N_21484,N_21344);
nand U27034 (N_27034,N_21648,N_20492);
nor U27035 (N_27035,N_20078,N_21277);
and U27036 (N_27036,N_23805,N_21982);
nor U27037 (N_27037,N_21956,N_23263);
and U27038 (N_27038,N_21873,N_22988);
and U27039 (N_27039,N_20452,N_24658);
nand U27040 (N_27040,N_21468,N_22124);
nor U27041 (N_27041,N_20535,N_22499);
or U27042 (N_27042,N_22667,N_24507);
or U27043 (N_27043,N_21586,N_23735);
or U27044 (N_27044,N_21361,N_24992);
or U27045 (N_27045,N_21988,N_23836);
nor U27046 (N_27046,N_24228,N_21974);
nand U27047 (N_27047,N_20423,N_24781);
or U27048 (N_27048,N_20662,N_22307);
nor U27049 (N_27049,N_20309,N_22636);
nor U27050 (N_27050,N_22696,N_20742);
or U27051 (N_27051,N_22770,N_21540);
nor U27052 (N_27052,N_23817,N_23104);
nand U27053 (N_27053,N_21387,N_23751);
and U27054 (N_27054,N_20029,N_23601);
nand U27055 (N_27055,N_24427,N_21541);
or U27056 (N_27056,N_24225,N_20071);
and U27057 (N_27057,N_23509,N_24327);
and U27058 (N_27058,N_21848,N_24412);
nand U27059 (N_27059,N_21287,N_22716);
and U27060 (N_27060,N_20873,N_20155);
nand U27061 (N_27061,N_22793,N_20390);
nand U27062 (N_27062,N_24638,N_24587);
and U27063 (N_27063,N_21327,N_23886);
or U27064 (N_27064,N_24026,N_22115);
and U27065 (N_27065,N_22411,N_21869);
nand U27066 (N_27066,N_22133,N_20977);
nor U27067 (N_27067,N_22090,N_21305);
and U27068 (N_27068,N_24653,N_23109);
nor U27069 (N_27069,N_23905,N_21045);
or U27070 (N_27070,N_22665,N_22364);
nor U27071 (N_27071,N_22127,N_20690);
nand U27072 (N_27072,N_24418,N_20332);
nand U27073 (N_27073,N_23766,N_24753);
nand U27074 (N_27074,N_22149,N_23647);
nor U27075 (N_27075,N_23327,N_21845);
and U27076 (N_27076,N_21430,N_24764);
nor U27077 (N_27077,N_23530,N_21306);
nor U27078 (N_27078,N_24561,N_22839);
nor U27079 (N_27079,N_24919,N_23117);
and U27080 (N_27080,N_24193,N_22143);
nand U27081 (N_27081,N_22161,N_21798);
nor U27082 (N_27082,N_23481,N_21025);
nor U27083 (N_27083,N_24331,N_24010);
nor U27084 (N_27084,N_21459,N_20612);
nand U27085 (N_27085,N_24250,N_24877);
nor U27086 (N_27086,N_22237,N_20400);
nor U27087 (N_27087,N_20741,N_20856);
nor U27088 (N_27088,N_23339,N_24613);
and U27089 (N_27089,N_24657,N_22923);
xnor U27090 (N_27090,N_22368,N_24395);
nor U27091 (N_27091,N_22805,N_21102);
or U27092 (N_27092,N_22799,N_23717);
or U27093 (N_27093,N_23814,N_24862);
nor U27094 (N_27094,N_22216,N_22827);
or U27095 (N_27095,N_22166,N_21646);
nor U27096 (N_27096,N_22635,N_20824);
nand U27097 (N_27097,N_21930,N_21214);
nand U27098 (N_27098,N_22468,N_24839);
nand U27099 (N_27099,N_22075,N_21577);
and U27100 (N_27100,N_24717,N_22642);
and U27101 (N_27101,N_20068,N_21473);
or U27102 (N_27102,N_24517,N_23907);
and U27103 (N_27103,N_20743,N_20667);
or U27104 (N_27104,N_20941,N_24358);
nand U27105 (N_27105,N_23046,N_22060);
nand U27106 (N_27106,N_20709,N_23610);
and U27107 (N_27107,N_23280,N_20910);
nand U27108 (N_27108,N_23559,N_23670);
nand U27109 (N_27109,N_22735,N_22140);
nor U27110 (N_27110,N_20717,N_23992);
nor U27111 (N_27111,N_20710,N_20450);
nor U27112 (N_27112,N_23320,N_24693);
or U27113 (N_27113,N_21877,N_22739);
and U27114 (N_27114,N_21945,N_22275);
nor U27115 (N_27115,N_21309,N_21384);
nand U27116 (N_27116,N_20376,N_21474);
nor U27117 (N_27117,N_23931,N_23865);
and U27118 (N_27118,N_24126,N_21617);
or U27119 (N_27119,N_20286,N_20164);
and U27120 (N_27120,N_24817,N_22732);
nor U27121 (N_27121,N_20839,N_24937);
or U27122 (N_27122,N_23211,N_24470);
and U27123 (N_27123,N_21986,N_22055);
and U27124 (N_27124,N_20531,N_21905);
or U27125 (N_27125,N_23393,N_21374);
or U27126 (N_27126,N_21920,N_20638);
nor U27127 (N_27127,N_20106,N_20104);
or U27128 (N_27128,N_20202,N_20498);
nor U27129 (N_27129,N_24710,N_22682);
and U27130 (N_27130,N_24647,N_22824);
or U27131 (N_27131,N_24144,N_24292);
and U27132 (N_27132,N_23299,N_21242);
nand U27133 (N_27133,N_24692,N_21554);
nand U27134 (N_27134,N_24651,N_20956);
or U27135 (N_27135,N_20532,N_23541);
and U27136 (N_27136,N_20828,N_23723);
and U27137 (N_27137,N_21224,N_21263);
nand U27138 (N_27138,N_20593,N_23724);
nand U27139 (N_27139,N_23616,N_23495);
nand U27140 (N_27140,N_24832,N_24809);
nand U27141 (N_27141,N_23346,N_23347);
and U27142 (N_27142,N_20988,N_24236);
nor U27143 (N_27143,N_21109,N_20147);
nand U27144 (N_27144,N_22984,N_22174);
and U27145 (N_27145,N_22913,N_21115);
or U27146 (N_27146,N_21587,N_24597);
and U27147 (N_27147,N_24070,N_22485);
or U27148 (N_27148,N_20372,N_21679);
or U27149 (N_27149,N_23155,N_24426);
or U27150 (N_27150,N_23366,N_20545);
or U27151 (N_27151,N_21152,N_21221);
or U27152 (N_27152,N_24245,N_20808);
or U27153 (N_27153,N_24151,N_22542);
nand U27154 (N_27154,N_23467,N_20798);
nand U27155 (N_27155,N_20080,N_20354);
nor U27156 (N_27156,N_24455,N_20762);
and U27157 (N_27157,N_21532,N_20663);
nand U27158 (N_27158,N_23957,N_24716);
nand U27159 (N_27159,N_23424,N_23545);
and U27160 (N_27160,N_24643,N_21404);
nand U27161 (N_27161,N_24841,N_20609);
or U27162 (N_27162,N_20641,N_21545);
or U27163 (N_27163,N_22378,N_24846);
nor U27164 (N_27164,N_24504,N_23761);
or U27165 (N_27165,N_24820,N_23536);
nand U27166 (N_27166,N_23038,N_23776);
or U27167 (N_27167,N_24784,N_22772);
and U27168 (N_27168,N_20113,N_20568);
nand U27169 (N_27169,N_22309,N_20060);
nand U27170 (N_27170,N_23269,N_22167);
nand U27171 (N_27171,N_24986,N_21666);
nor U27172 (N_27172,N_24220,N_23106);
nand U27173 (N_27173,N_22438,N_23888);
or U27174 (N_27174,N_24974,N_21557);
and U27175 (N_27175,N_20781,N_24373);
and U27176 (N_27176,N_21328,N_24706);
nand U27177 (N_27177,N_22412,N_22627);
nand U27178 (N_27178,N_24125,N_20978);
and U27179 (N_27179,N_20991,N_24713);
nand U27180 (N_27180,N_24911,N_23813);
and U27181 (N_27181,N_20976,N_22633);
and U27182 (N_27182,N_24599,N_21603);
and U27183 (N_27183,N_20434,N_21308);
or U27184 (N_27184,N_23701,N_22685);
and U27185 (N_27185,N_22227,N_22569);
nor U27186 (N_27186,N_24836,N_20887);
or U27187 (N_27187,N_20022,N_20428);
or U27188 (N_27188,N_23135,N_22303);
or U27189 (N_27189,N_22624,N_24191);
nand U27190 (N_27190,N_20156,N_23300);
nand U27191 (N_27191,N_24777,N_23260);
nor U27192 (N_27192,N_21883,N_23115);
and U27193 (N_27193,N_20459,N_24895);
or U27194 (N_27194,N_20897,N_20324);
nor U27195 (N_27195,N_20406,N_21735);
nor U27196 (N_27196,N_24190,N_21728);
or U27197 (N_27197,N_23392,N_22979);
nand U27198 (N_27198,N_23792,N_23315);
nor U27199 (N_27199,N_21923,N_20983);
nand U27200 (N_27200,N_23797,N_22936);
nor U27201 (N_27201,N_23048,N_22859);
or U27202 (N_27202,N_23744,N_24618);
or U27203 (N_27203,N_23474,N_24840);
and U27204 (N_27204,N_24181,N_23070);
or U27205 (N_27205,N_20854,N_24816);
and U27206 (N_27206,N_20579,N_22208);
or U27207 (N_27207,N_24525,N_24589);
nand U27208 (N_27208,N_21782,N_20277);
xnor U27209 (N_27209,N_24967,N_22888);
and U27210 (N_27210,N_24097,N_20464);
nor U27211 (N_27211,N_22410,N_22459);
and U27212 (N_27212,N_22557,N_23382);
nand U27213 (N_27213,N_24083,N_22043);
nor U27214 (N_27214,N_20074,N_24752);
xnor U27215 (N_27215,N_24164,N_20105);
or U27216 (N_27216,N_24901,N_23213);
and U27217 (N_27217,N_20035,N_21410);
nand U27218 (N_27218,N_21980,N_24594);
and U27219 (N_27219,N_21380,N_21694);
or U27220 (N_27220,N_21009,N_23592);
or U27221 (N_27221,N_20289,N_24649);
or U27222 (N_27222,N_24488,N_24211);
and U27223 (N_27223,N_20773,N_20522);
and U27224 (N_27224,N_21181,N_24887);
or U27225 (N_27225,N_22471,N_20395);
or U27226 (N_27226,N_21127,N_23177);
and U27227 (N_27227,N_20439,N_22811);
nand U27228 (N_27228,N_24487,N_24727);
or U27229 (N_27229,N_21332,N_23376);
nor U27230 (N_27230,N_24120,N_23993);
and U27231 (N_27231,N_23878,N_22523);
nand U27232 (N_27232,N_21229,N_23296);
nor U27233 (N_27233,N_20290,N_24390);
and U27234 (N_27234,N_23950,N_21668);
and U27235 (N_27235,N_23037,N_23528);
nor U27236 (N_27236,N_20945,N_24747);
nand U27237 (N_27237,N_23407,N_23419);
and U27238 (N_27238,N_23127,N_21653);
or U27239 (N_27239,N_24987,N_20257);
or U27240 (N_27240,N_21833,N_23507);
nand U27241 (N_27241,N_20617,N_20716);
and U27242 (N_27242,N_23110,N_20481);
and U27243 (N_27243,N_24860,N_24748);
and U27244 (N_27244,N_24453,N_21346);
nor U27245 (N_27245,N_22057,N_21059);
or U27246 (N_27246,N_22733,N_23150);
nand U27247 (N_27247,N_22721,N_20712);
nand U27248 (N_27248,N_20430,N_24157);
nand U27249 (N_27249,N_24166,N_20251);
and U27250 (N_27250,N_21829,N_24284);
nand U27251 (N_27251,N_23764,N_21382);
and U27252 (N_27252,N_22098,N_21182);
and U27253 (N_27253,N_21622,N_22738);
or U27254 (N_27254,N_21443,N_23819);
or U27255 (N_27255,N_23126,N_24162);
or U27256 (N_27256,N_23245,N_22146);
and U27257 (N_27257,N_21175,N_20340);
nor U27258 (N_27258,N_22968,N_22536);
nor U27259 (N_27259,N_23003,N_24815);
nand U27260 (N_27260,N_22285,N_24916);
nor U27261 (N_27261,N_22488,N_20380);
nand U27262 (N_27262,N_23244,N_21151);
nand U27263 (N_27263,N_23402,N_22899);
nor U27264 (N_27264,N_22691,N_20812);
nand U27265 (N_27265,N_20735,N_22264);
nand U27266 (N_27266,N_24023,N_20965);
and U27267 (N_27267,N_24571,N_22511);
nand U27268 (N_27268,N_22982,N_23114);
or U27269 (N_27269,N_20749,N_23143);
nor U27270 (N_27270,N_22802,N_20953);
or U27271 (N_27271,N_22463,N_24849);
nor U27272 (N_27272,N_20426,N_21492);
nor U27273 (N_27273,N_23855,N_22617);
and U27274 (N_27274,N_20108,N_20418);
and U27275 (N_27275,N_22815,N_24405);
nor U27276 (N_27276,N_21707,N_22871);
nor U27277 (N_27277,N_23572,N_21715);
nand U27278 (N_27278,N_24037,N_21867);
nand U27279 (N_27279,N_23072,N_20513);
and U27280 (N_27280,N_24723,N_21487);
nor U27281 (N_27281,N_21052,N_24819);
and U27282 (N_27282,N_23617,N_24443);
nor U27283 (N_27283,N_20555,N_20445);
nor U27284 (N_27284,N_23871,N_22679);
or U27285 (N_27285,N_22190,N_21453);
nor U27286 (N_27286,N_20339,N_24462);
and U27287 (N_27287,N_22734,N_21658);
nor U27288 (N_27288,N_21296,N_24004);
or U27289 (N_27289,N_22044,N_20127);
or U27290 (N_27290,N_24677,N_21797);
nor U27291 (N_27291,N_23949,N_24160);
and U27292 (N_27292,N_22535,N_22528);
nand U27293 (N_27293,N_23549,N_22580);
or U27294 (N_27294,N_24609,N_20192);
nor U27295 (N_27295,N_22012,N_20417);
xnor U27296 (N_27296,N_20578,N_24482);
or U27297 (N_27297,N_22330,N_23278);
nor U27298 (N_27298,N_24714,N_20993);
and U27299 (N_27299,N_23399,N_23119);
nand U27300 (N_27300,N_23023,N_23497);
nor U27301 (N_27301,N_22562,N_20960);
nand U27302 (N_27302,N_22604,N_22723);
nor U27303 (N_27303,N_21698,N_23620);
nand U27304 (N_27304,N_24388,N_20503);
and U27305 (N_27305,N_20679,N_22013);
and U27306 (N_27306,N_20921,N_21450);
nand U27307 (N_27307,N_20936,N_23974);
nor U27308 (N_27308,N_21293,N_22956);
nor U27309 (N_27309,N_21900,N_20546);
nand U27310 (N_27310,N_24498,N_21171);
nand U27311 (N_27311,N_23924,N_21816);
and U27312 (N_27312,N_21561,N_20863);
nand U27313 (N_27313,N_20477,N_20349);
or U27314 (N_27314,N_22258,N_24486);
nor U27315 (N_27315,N_23718,N_22102);
xor U27316 (N_27316,N_21159,N_21043);
or U27317 (N_27317,N_21481,N_23168);
and U27318 (N_27318,N_23077,N_21188);
nand U27319 (N_27319,N_22606,N_22424);
nand U27320 (N_27320,N_21007,N_22371);
nand U27321 (N_27321,N_21186,N_20280);
and U27322 (N_27322,N_24449,N_21675);
or U27323 (N_27323,N_20598,N_23749);
or U27324 (N_27324,N_23550,N_23730);
nor U27325 (N_27325,N_20386,N_22554);
and U27326 (N_27326,N_20365,N_21696);
nor U27327 (N_27327,N_22518,N_22287);
or U27328 (N_27328,N_23663,N_21801);
and U27329 (N_27329,N_20530,N_23412);
or U27330 (N_27330,N_20512,N_20416);
nand U27331 (N_27331,N_24296,N_22993);
nor U27332 (N_27332,N_24047,N_23417);
and U27333 (N_27333,N_21552,N_20115);
nor U27334 (N_27334,N_23644,N_24999);
nor U27335 (N_27335,N_23654,N_22268);
nand U27336 (N_27336,N_23631,N_20970);
and U27337 (N_27337,N_22754,N_20721);
nand U27338 (N_27338,N_24965,N_24800);
or U27339 (N_27339,N_22180,N_24402);
and U27340 (N_27340,N_22720,N_23728);
and U27341 (N_27341,N_21849,N_24180);
nor U27342 (N_27342,N_24961,N_20040);
nand U27343 (N_27343,N_23891,N_23397);
nor U27344 (N_27344,N_22426,N_21482);
or U27345 (N_27345,N_24415,N_24297);
nor U27346 (N_27346,N_21914,N_20850);
or U27347 (N_27347,N_23252,N_24425);
or U27348 (N_27348,N_24890,N_24876);
or U27349 (N_27349,N_21070,N_22879);
and U27350 (N_27350,N_23433,N_23492);
nor U27351 (N_27351,N_21823,N_23275);
nor U27352 (N_27352,N_20130,N_20592);
or U27353 (N_27353,N_23094,N_24736);
and U27354 (N_27354,N_22508,N_20382);
and U27355 (N_27355,N_21701,N_24646);
or U27356 (N_27356,N_20574,N_23599);
nand U27357 (N_27357,N_24768,N_23449);
nand U27358 (N_27358,N_23781,N_24227);
nand U27359 (N_27359,N_23746,N_20560);
or U27360 (N_27360,N_22314,N_21791);
nor U27361 (N_27361,N_24740,N_24793);
or U27362 (N_27362,N_20157,N_21769);
and U27363 (N_27363,N_24031,N_23719);
and U27364 (N_27364,N_24616,N_24627);
and U27365 (N_27365,N_23656,N_21997);
or U27366 (N_27366,N_22527,N_24050);
nor U27367 (N_27367,N_22283,N_20397);
or U27368 (N_27368,N_20471,N_20163);
nor U27369 (N_27369,N_23033,N_20517);
or U27370 (N_27370,N_22182,N_22680);
and U27371 (N_27371,N_23461,N_24506);
and U27372 (N_27372,N_20585,N_21370);
or U27373 (N_27373,N_22940,N_21688);
nor U27374 (N_27374,N_24260,N_22112);
and U27375 (N_27375,N_20001,N_22572);
nand U27376 (N_27376,N_22651,N_24976);
nand U27377 (N_27377,N_24523,N_24508);
nand U27378 (N_27378,N_21034,N_20724);
or U27379 (N_27379,N_22931,N_24241);
nor U27380 (N_27380,N_21626,N_20559);
nor U27381 (N_27381,N_24027,N_23183);
and U27382 (N_27382,N_22741,N_24835);
and U27383 (N_27383,N_22328,N_20458);
nor U27384 (N_27384,N_21924,N_24113);
nor U27385 (N_27385,N_24721,N_21768);
and U27386 (N_27386,N_20518,N_21659);
nand U27387 (N_27387,N_21888,N_23903);
nand U27388 (N_27388,N_21534,N_24471);
or U27389 (N_27389,N_20438,N_22469);
or U27390 (N_27390,N_20499,N_24694);
nor U27391 (N_27391,N_23355,N_22134);
nand U27392 (N_27392,N_20928,N_20437);
or U27393 (N_27393,N_22153,N_24758);
nor U27394 (N_27394,N_23588,N_21574);
nor U27395 (N_27395,N_23456,N_21131);
nand U27396 (N_27396,N_20889,N_21882);
nand U27397 (N_27397,N_24799,N_20310);
or U27398 (N_27398,N_24932,N_20783);
nor U27399 (N_27399,N_21926,N_24858);
nand U27400 (N_27400,N_21917,N_22111);
or U27401 (N_27401,N_22560,N_23996);
nor U27402 (N_27402,N_20235,N_24639);
nand U27403 (N_27403,N_20506,N_23483);
nand U27404 (N_27404,N_23335,N_21333);
nor U27405 (N_27405,N_21149,N_21426);
nor U27406 (N_27406,N_24898,N_24454);
or U27407 (N_27407,N_22329,N_20772);
and U27408 (N_27408,N_22475,N_24600);
or U27409 (N_27409,N_24276,N_21576);
nor U27410 (N_27410,N_20736,N_21619);
nand U27411 (N_27411,N_22803,N_24743);
xnor U27412 (N_27412,N_22065,N_20875);
and U27413 (N_27413,N_22740,N_22139);
nand U27414 (N_27414,N_21743,N_22288);
nand U27415 (N_27415,N_22755,N_23370);
or U27416 (N_27416,N_22534,N_20356);
or U27417 (N_27417,N_24337,N_23569);
or U27418 (N_27418,N_23438,N_20588);
nand U27419 (N_27419,N_21977,N_21161);
and U27420 (N_27420,N_20329,N_24977);
nand U27421 (N_27421,N_23551,N_22160);
nor U27422 (N_27422,N_21871,N_21560);
nand U27423 (N_27423,N_23738,N_24856);
nor U27424 (N_27424,N_20548,N_24244);
and U27425 (N_27425,N_22608,N_22458);
nor U27426 (N_27426,N_21972,N_22607);
and U27427 (N_27427,N_22818,N_21432);
xor U27428 (N_27428,N_20121,N_22880);
and U27429 (N_27429,N_23673,N_24108);
or U27430 (N_27430,N_20764,N_23825);
or U27431 (N_27431,N_22428,N_22046);
and U27432 (N_27432,N_22538,N_23173);
nor U27433 (N_27433,N_20358,N_20629);
nand U27434 (N_27434,N_20322,N_23882);
nor U27435 (N_27435,N_24814,N_22692);
nand U27436 (N_27436,N_20831,N_24167);
nand U27437 (N_27437,N_20768,N_23935);
or U27438 (N_27438,N_20833,N_22653);
or U27439 (N_27439,N_22027,N_23167);
nor U27440 (N_27440,N_24335,N_24912);
or U27441 (N_27441,N_22513,N_23373);
or U27442 (N_27442,N_21697,N_24460);
or U27443 (N_27443,N_22291,N_23919);
xnor U27444 (N_27444,N_22009,N_20615);
and U27445 (N_27445,N_20803,N_22589);
and U27446 (N_27446,N_23063,N_22456);
nand U27447 (N_27447,N_23862,N_21315);
or U27448 (N_27448,N_23912,N_23285);
and U27449 (N_27449,N_22619,N_24432);
nor U27450 (N_27450,N_22628,N_20892);
or U27451 (N_27451,N_21347,N_20566);
nor U27452 (N_27452,N_23704,N_20826);
and U27453 (N_27453,N_20652,N_24001);
or U27454 (N_27454,N_23232,N_20676);
nand U27455 (N_27455,N_23377,N_23904);
nor U27456 (N_27456,N_21708,N_23837);
or U27457 (N_27457,N_20827,N_24338);
or U27458 (N_27458,N_24210,N_23107);
and U27459 (N_27459,N_21794,N_21757);
nand U27460 (N_27460,N_22706,N_23892);
nand U27461 (N_27461,N_23490,N_24993);
nor U27462 (N_27462,N_20602,N_20338);
and U27463 (N_27463,N_23175,N_24625);
or U27464 (N_27464,N_22360,N_24046);
and U27465 (N_27465,N_21667,N_22104);
nand U27466 (N_27466,N_22038,N_22506);
nand U27467 (N_27467,N_20866,N_23108);
nor U27468 (N_27468,N_24690,N_21929);
and U27469 (N_27469,N_21028,N_20051);
and U27470 (N_27470,N_21907,N_24791);
nand U27471 (N_27471,N_24069,N_23827);
or U27472 (N_27472,N_20367,N_20605);
nand U27473 (N_27473,N_21908,N_21544);
nor U27474 (N_27474,N_20208,N_23708);
nor U27475 (N_27475,N_20088,N_22932);
nor U27476 (N_27476,N_21322,N_20732);
xor U27477 (N_27477,N_23343,N_23318);
or U27478 (N_27478,N_23816,N_21885);
or U27479 (N_27479,N_23590,N_21531);
nor U27480 (N_27480,N_22700,N_21936);
or U27481 (N_27481,N_20032,N_21056);
nor U27482 (N_27482,N_23645,N_23725);
nand U27483 (N_27483,N_21447,N_20211);
nand U27484 (N_27484,N_22575,N_21633);
and U27485 (N_27485,N_20747,N_20361);
or U27486 (N_27486,N_20353,N_20486);
nor U27487 (N_27487,N_22612,N_23319);
and U27488 (N_27488,N_23221,N_24683);
or U27489 (N_27489,N_21386,N_21756);
nor U27490 (N_27490,N_24115,N_23489);
nand U27491 (N_27491,N_23288,N_20441);
or U27492 (N_27492,N_20534,N_23804);
and U27493 (N_27493,N_21803,N_22609);
nor U27494 (N_27494,N_23055,N_21217);
and U27495 (N_27495,N_22690,N_20204);
nor U27496 (N_27496,N_21946,N_22725);
nand U27497 (N_27497,N_22882,N_22341);
nor U27498 (N_27498,N_23341,N_23712);
or U27499 (N_27499,N_23743,N_23365);
nor U27500 (N_27500,N_22670,N_22229);
nand U27501 (N_27501,N_22608,N_23021);
or U27502 (N_27502,N_20018,N_22399);
or U27503 (N_27503,N_22896,N_22532);
or U27504 (N_27504,N_20593,N_22081);
and U27505 (N_27505,N_21468,N_23384);
and U27506 (N_27506,N_23378,N_23571);
nand U27507 (N_27507,N_20585,N_20550);
or U27508 (N_27508,N_24229,N_24862);
nor U27509 (N_27509,N_20343,N_23514);
nor U27510 (N_27510,N_20572,N_23100);
or U27511 (N_27511,N_21529,N_20718);
or U27512 (N_27512,N_23699,N_21451);
or U27513 (N_27513,N_23084,N_22327);
or U27514 (N_27514,N_21661,N_24460);
or U27515 (N_27515,N_20413,N_24130);
or U27516 (N_27516,N_21753,N_22213);
or U27517 (N_27517,N_22025,N_20523);
and U27518 (N_27518,N_21404,N_23329);
and U27519 (N_27519,N_20696,N_21686);
or U27520 (N_27520,N_23702,N_22848);
nand U27521 (N_27521,N_20328,N_22642);
and U27522 (N_27522,N_20388,N_22543);
or U27523 (N_27523,N_22783,N_24047);
and U27524 (N_27524,N_21084,N_22502);
or U27525 (N_27525,N_21644,N_22987);
nor U27526 (N_27526,N_20782,N_23405);
nand U27527 (N_27527,N_21234,N_21866);
or U27528 (N_27528,N_22914,N_24574);
or U27529 (N_27529,N_21058,N_24136);
nand U27530 (N_27530,N_24391,N_24298);
and U27531 (N_27531,N_22381,N_24436);
nand U27532 (N_27532,N_24329,N_23970);
nand U27533 (N_27533,N_21825,N_20368);
or U27534 (N_27534,N_21430,N_22942);
and U27535 (N_27535,N_20954,N_22243);
and U27536 (N_27536,N_23317,N_23017);
and U27537 (N_27537,N_20786,N_22918);
nor U27538 (N_27538,N_24812,N_23543);
or U27539 (N_27539,N_21605,N_20519);
nor U27540 (N_27540,N_22907,N_20912);
or U27541 (N_27541,N_21205,N_22159);
nand U27542 (N_27542,N_21820,N_23185);
nand U27543 (N_27543,N_21894,N_24736);
or U27544 (N_27544,N_23556,N_22188);
and U27545 (N_27545,N_20738,N_20723);
nor U27546 (N_27546,N_22478,N_21590);
or U27547 (N_27547,N_20372,N_24222);
or U27548 (N_27548,N_20350,N_20392);
and U27549 (N_27549,N_24380,N_21244);
nand U27550 (N_27550,N_23078,N_22024);
xnor U27551 (N_27551,N_24889,N_21531);
nand U27552 (N_27552,N_24393,N_22031);
or U27553 (N_27553,N_24429,N_22537);
or U27554 (N_27554,N_20737,N_23403);
nor U27555 (N_27555,N_22921,N_21935);
and U27556 (N_27556,N_22431,N_21986);
nand U27557 (N_27557,N_24917,N_23200);
nor U27558 (N_27558,N_21945,N_22918);
nand U27559 (N_27559,N_21981,N_23982);
or U27560 (N_27560,N_24490,N_20247);
nand U27561 (N_27561,N_24354,N_20019);
or U27562 (N_27562,N_21419,N_23988);
nand U27563 (N_27563,N_22288,N_24360);
or U27564 (N_27564,N_21804,N_23834);
nor U27565 (N_27565,N_22978,N_21976);
nand U27566 (N_27566,N_20243,N_21608);
nor U27567 (N_27567,N_23247,N_20139);
and U27568 (N_27568,N_20229,N_20889);
and U27569 (N_27569,N_21575,N_22618);
nor U27570 (N_27570,N_24121,N_22021);
nand U27571 (N_27571,N_23860,N_24309);
nor U27572 (N_27572,N_23788,N_23647);
or U27573 (N_27573,N_24183,N_21866);
and U27574 (N_27574,N_22129,N_20203);
and U27575 (N_27575,N_22996,N_20307);
and U27576 (N_27576,N_23915,N_22087);
or U27577 (N_27577,N_20988,N_21978);
and U27578 (N_27578,N_21242,N_20439);
nand U27579 (N_27579,N_24377,N_20171);
or U27580 (N_27580,N_20650,N_24208);
nor U27581 (N_27581,N_22563,N_23417);
and U27582 (N_27582,N_20954,N_22099);
nor U27583 (N_27583,N_23583,N_21668);
nand U27584 (N_27584,N_23485,N_20249);
xnor U27585 (N_27585,N_24153,N_22658);
and U27586 (N_27586,N_22767,N_22100);
or U27587 (N_27587,N_23365,N_23145);
and U27588 (N_27588,N_23763,N_23137);
or U27589 (N_27589,N_22540,N_20600);
xor U27590 (N_27590,N_21581,N_23496);
nand U27591 (N_27591,N_22700,N_23046);
nor U27592 (N_27592,N_23578,N_23217);
or U27593 (N_27593,N_24161,N_20322);
nor U27594 (N_27594,N_23816,N_20171);
nand U27595 (N_27595,N_21794,N_23593);
or U27596 (N_27596,N_20886,N_23372);
nand U27597 (N_27597,N_23981,N_22183);
nand U27598 (N_27598,N_21133,N_20442);
and U27599 (N_27599,N_24571,N_20127);
nor U27600 (N_27600,N_21527,N_23587);
nand U27601 (N_27601,N_20374,N_22519);
or U27602 (N_27602,N_23357,N_21070);
nand U27603 (N_27603,N_22000,N_22650);
nand U27604 (N_27604,N_22239,N_20151);
nor U27605 (N_27605,N_24388,N_22526);
and U27606 (N_27606,N_22872,N_22818);
or U27607 (N_27607,N_21020,N_23797);
nand U27608 (N_27608,N_21181,N_20986);
and U27609 (N_27609,N_22602,N_23130);
and U27610 (N_27610,N_22943,N_24750);
nand U27611 (N_27611,N_22194,N_22732);
nor U27612 (N_27612,N_23958,N_22792);
and U27613 (N_27613,N_23353,N_23066);
or U27614 (N_27614,N_20586,N_22183);
nand U27615 (N_27615,N_22748,N_24740);
nand U27616 (N_27616,N_22796,N_23084);
nand U27617 (N_27617,N_22469,N_23866);
nand U27618 (N_27618,N_23807,N_21315);
nor U27619 (N_27619,N_24366,N_23069);
or U27620 (N_27620,N_23666,N_24930);
nand U27621 (N_27621,N_21597,N_22472);
nor U27622 (N_27622,N_24657,N_22223);
or U27623 (N_27623,N_22646,N_22350);
and U27624 (N_27624,N_22710,N_23706);
nand U27625 (N_27625,N_20934,N_24404);
nand U27626 (N_27626,N_23386,N_20845);
and U27627 (N_27627,N_21625,N_20443);
or U27628 (N_27628,N_22989,N_21864);
and U27629 (N_27629,N_24745,N_22907);
and U27630 (N_27630,N_22562,N_20839);
and U27631 (N_27631,N_23990,N_23430);
nand U27632 (N_27632,N_22096,N_24243);
nor U27633 (N_27633,N_21672,N_22878);
and U27634 (N_27634,N_23606,N_24735);
nor U27635 (N_27635,N_21900,N_23080);
nor U27636 (N_27636,N_22132,N_23650);
nor U27637 (N_27637,N_21485,N_22412);
and U27638 (N_27638,N_24995,N_21745);
or U27639 (N_27639,N_23983,N_20763);
and U27640 (N_27640,N_21905,N_24394);
nor U27641 (N_27641,N_23022,N_22115);
nand U27642 (N_27642,N_22793,N_20129);
nor U27643 (N_27643,N_22515,N_23398);
or U27644 (N_27644,N_20108,N_20885);
nand U27645 (N_27645,N_24129,N_21215);
and U27646 (N_27646,N_24382,N_23129);
nor U27647 (N_27647,N_22989,N_22897);
nor U27648 (N_27648,N_22558,N_22412);
and U27649 (N_27649,N_24889,N_24397);
or U27650 (N_27650,N_24519,N_22590);
or U27651 (N_27651,N_23889,N_21363);
nor U27652 (N_27652,N_21456,N_22803);
nor U27653 (N_27653,N_22300,N_21091);
or U27654 (N_27654,N_23130,N_24003);
nand U27655 (N_27655,N_21571,N_20277);
nor U27656 (N_27656,N_20303,N_23205);
or U27657 (N_27657,N_24202,N_21514);
and U27658 (N_27658,N_23275,N_21426);
and U27659 (N_27659,N_23371,N_20417);
or U27660 (N_27660,N_21242,N_24946);
nor U27661 (N_27661,N_20132,N_23115);
nor U27662 (N_27662,N_21449,N_20750);
and U27663 (N_27663,N_23272,N_24478);
nand U27664 (N_27664,N_24650,N_23778);
nor U27665 (N_27665,N_24160,N_23615);
nor U27666 (N_27666,N_20652,N_21722);
or U27667 (N_27667,N_22660,N_23774);
or U27668 (N_27668,N_24918,N_22849);
and U27669 (N_27669,N_23613,N_21631);
nand U27670 (N_27670,N_22556,N_24681);
nand U27671 (N_27671,N_22472,N_23739);
nand U27672 (N_27672,N_20012,N_22820);
and U27673 (N_27673,N_23187,N_21850);
or U27674 (N_27674,N_20950,N_20297);
nor U27675 (N_27675,N_24687,N_20948);
nand U27676 (N_27676,N_22494,N_23964);
and U27677 (N_27677,N_24474,N_20250);
nor U27678 (N_27678,N_22178,N_21562);
and U27679 (N_27679,N_23106,N_20658);
and U27680 (N_27680,N_21440,N_23783);
nor U27681 (N_27681,N_24910,N_20392);
xor U27682 (N_27682,N_20515,N_22568);
nand U27683 (N_27683,N_20125,N_21329);
and U27684 (N_27684,N_21912,N_24116);
nor U27685 (N_27685,N_20927,N_23916);
and U27686 (N_27686,N_21785,N_23858);
and U27687 (N_27687,N_22683,N_22300);
nand U27688 (N_27688,N_20036,N_23614);
nand U27689 (N_27689,N_24294,N_23935);
and U27690 (N_27690,N_21499,N_22775);
or U27691 (N_27691,N_23672,N_22295);
nor U27692 (N_27692,N_21705,N_22190);
or U27693 (N_27693,N_24514,N_23926);
nor U27694 (N_27694,N_24716,N_23403);
nor U27695 (N_27695,N_21250,N_23899);
or U27696 (N_27696,N_20786,N_20234);
nand U27697 (N_27697,N_21426,N_22590);
nor U27698 (N_27698,N_22698,N_21669);
and U27699 (N_27699,N_20868,N_20861);
and U27700 (N_27700,N_20685,N_24125);
nand U27701 (N_27701,N_24773,N_23401);
or U27702 (N_27702,N_22968,N_21544);
nor U27703 (N_27703,N_22215,N_22055);
xor U27704 (N_27704,N_23799,N_23750);
and U27705 (N_27705,N_24314,N_24926);
nand U27706 (N_27706,N_24709,N_20559);
or U27707 (N_27707,N_24566,N_22263);
and U27708 (N_27708,N_21375,N_23177);
or U27709 (N_27709,N_23187,N_23140);
nand U27710 (N_27710,N_20565,N_21392);
nor U27711 (N_27711,N_22242,N_21152);
nor U27712 (N_27712,N_23054,N_21499);
nand U27713 (N_27713,N_20676,N_23974);
nand U27714 (N_27714,N_23710,N_24790);
nor U27715 (N_27715,N_21940,N_23448);
nor U27716 (N_27716,N_20205,N_20580);
and U27717 (N_27717,N_21534,N_23109);
or U27718 (N_27718,N_24735,N_23775);
and U27719 (N_27719,N_20524,N_22783);
and U27720 (N_27720,N_21017,N_20293);
nor U27721 (N_27721,N_20143,N_22397);
nor U27722 (N_27722,N_22442,N_23328);
nor U27723 (N_27723,N_21125,N_24317);
nand U27724 (N_27724,N_23739,N_24461);
nand U27725 (N_27725,N_20948,N_20111);
nand U27726 (N_27726,N_22248,N_24036);
and U27727 (N_27727,N_20449,N_24318);
nor U27728 (N_27728,N_24673,N_23045);
or U27729 (N_27729,N_23128,N_20059);
nand U27730 (N_27730,N_23922,N_21164);
and U27731 (N_27731,N_21587,N_23276);
nand U27732 (N_27732,N_22730,N_20194);
nand U27733 (N_27733,N_20081,N_21835);
or U27734 (N_27734,N_21132,N_21792);
nor U27735 (N_27735,N_20944,N_24971);
nand U27736 (N_27736,N_24330,N_24759);
and U27737 (N_27737,N_24985,N_21336);
nand U27738 (N_27738,N_23320,N_20484);
and U27739 (N_27739,N_23149,N_22547);
or U27740 (N_27740,N_21312,N_22086);
and U27741 (N_27741,N_20566,N_20614);
nand U27742 (N_27742,N_21760,N_22903);
nor U27743 (N_27743,N_23923,N_20628);
nand U27744 (N_27744,N_24586,N_23092);
nand U27745 (N_27745,N_23525,N_20110);
nand U27746 (N_27746,N_24865,N_21814);
and U27747 (N_27747,N_21399,N_23933);
or U27748 (N_27748,N_24327,N_23505);
and U27749 (N_27749,N_22979,N_21862);
and U27750 (N_27750,N_21348,N_21625);
nor U27751 (N_27751,N_21218,N_20914);
nor U27752 (N_27752,N_22635,N_24686);
or U27753 (N_27753,N_21663,N_23595);
nor U27754 (N_27754,N_23244,N_23491);
nand U27755 (N_27755,N_20269,N_22717);
nand U27756 (N_27756,N_20462,N_22292);
nand U27757 (N_27757,N_23365,N_20505);
or U27758 (N_27758,N_24075,N_22613);
nor U27759 (N_27759,N_21178,N_24681);
nor U27760 (N_27760,N_24640,N_22797);
nand U27761 (N_27761,N_22460,N_21136);
nor U27762 (N_27762,N_23501,N_22727);
nand U27763 (N_27763,N_23608,N_23144);
nand U27764 (N_27764,N_24585,N_24178);
and U27765 (N_27765,N_22940,N_23237);
or U27766 (N_27766,N_22139,N_23772);
or U27767 (N_27767,N_22609,N_21706);
or U27768 (N_27768,N_20775,N_20475);
or U27769 (N_27769,N_24457,N_20626);
nor U27770 (N_27770,N_24663,N_20901);
nor U27771 (N_27771,N_23775,N_20851);
nand U27772 (N_27772,N_22455,N_21877);
or U27773 (N_27773,N_21561,N_21140);
nand U27774 (N_27774,N_24229,N_20567);
or U27775 (N_27775,N_23063,N_24186);
nor U27776 (N_27776,N_24566,N_20183);
or U27777 (N_27777,N_20515,N_24323);
and U27778 (N_27778,N_22915,N_23503);
and U27779 (N_27779,N_22006,N_24306);
or U27780 (N_27780,N_20188,N_22129);
nand U27781 (N_27781,N_21410,N_23341);
nor U27782 (N_27782,N_23095,N_24462);
nor U27783 (N_27783,N_24013,N_22519);
and U27784 (N_27784,N_22502,N_23077);
nor U27785 (N_27785,N_22971,N_22249);
and U27786 (N_27786,N_22564,N_23904);
or U27787 (N_27787,N_21318,N_22888);
and U27788 (N_27788,N_20016,N_21842);
nand U27789 (N_27789,N_22925,N_22034);
nand U27790 (N_27790,N_21629,N_22215);
nand U27791 (N_27791,N_20782,N_23774);
xnor U27792 (N_27792,N_20111,N_21469);
nand U27793 (N_27793,N_21417,N_23367);
or U27794 (N_27794,N_20472,N_23301);
nor U27795 (N_27795,N_20665,N_23789);
nand U27796 (N_27796,N_22354,N_23314);
nand U27797 (N_27797,N_21628,N_24687);
nand U27798 (N_27798,N_22362,N_24051);
nand U27799 (N_27799,N_20762,N_20126);
nand U27800 (N_27800,N_24211,N_22598);
nand U27801 (N_27801,N_24253,N_20457);
and U27802 (N_27802,N_23794,N_21243);
nor U27803 (N_27803,N_21298,N_20131);
nor U27804 (N_27804,N_21929,N_21723);
or U27805 (N_27805,N_22782,N_22224);
nand U27806 (N_27806,N_22292,N_20499);
nand U27807 (N_27807,N_20662,N_20855);
and U27808 (N_27808,N_24333,N_20942);
nand U27809 (N_27809,N_20278,N_21499);
nor U27810 (N_27810,N_24993,N_22580);
nor U27811 (N_27811,N_20632,N_24120);
nand U27812 (N_27812,N_21812,N_24382);
nand U27813 (N_27813,N_23811,N_24056);
or U27814 (N_27814,N_23027,N_22929);
or U27815 (N_27815,N_24713,N_23300);
nor U27816 (N_27816,N_22617,N_22858);
and U27817 (N_27817,N_24361,N_23674);
nand U27818 (N_27818,N_20261,N_24195);
or U27819 (N_27819,N_22162,N_23921);
or U27820 (N_27820,N_20279,N_21689);
nand U27821 (N_27821,N_20943,N_21623);
and U27822 (N_27822,N_23035,N_20881);
or U27823 (N_27823,N_21916,N_20637);
and U27824 (N_27824,N_23489,N_24743);
nand U27825 (N_27825,N_23730,N_20187);
or U27826 (N_27826,N_20528,N_24877);
nor U27827 (N_27827,N_22547,N_23897);
or U27828 (N_27828,N_23065,N_21401);
and U27829 (N_27829,N_20050,N_21870);
and U27830 (N_27830,N_21121,N_21278);
nor U27831 (N_27831,N_23772,N_24657);
or U27832 (N_27832,N_24775,N_21098);
xor U27833 (N_27833,N_22757,N_23278);
and U27834 (N_27834,N_23802,N_21350);
and U27835 (N_27835,N_23070,N_24992);
or U27836 (N_27836,N_24268,N_22256);
nand U27837 (N_27837,N_22540,N_20220);
and U27838 (N_27838,N_23404,N_24964);
nand U27839 (N_27839,N_21310,N_24325);
or U27840 (N_27840,N_21385,N_24739);
nand U27841 (N_27841,N_21487,N_20563);
and U27842 (N_27842,N_22846,N_20257);
nand U27843 (N_27843,N_24191,N_23995);
or U27844 (N_27844,N_24074,N_22286);
and U27845 (N_27845,N_21401,N_24416);
nand U27846 (N_27846,N_20192,N_23464);
or U27847 (N_27847,N_22358,N_21130);
nand U27848 (N_27848,N_22225,N_21363);
nor U27849 (N_27849,N_23202,N_24011);
nand U27850 (N_27850,N_24981,N_22814);
nand U27851 (N_27851,N_20125,N_24291);
nand U27852 (N_27852,N_22154,N_20404);
or U27853 (N_27853,N_21694,N_20540);
and U27854 (N_27854,N_21185,N_23648);
nand U27855 (N_27855,N_23337,N_23225);
and U27856 (N_27856,N_21266,N_24011);
nand U27857 (N_27857,N_23232,N_21206);
or U27858 (N_27858,N_20078,N_22111);
or U27859 (N_27859,N_22278,N_24112);
and U27860 (N_27860,N_23042,N_22816);
and U27861 (N_27861,N_22143,N_24884);
or U27862 (N_27862,N_24207,N_23236);
nand U27863 (N_27863,N_21040,N_24956);
or U27864 (N_27864,N_23995,N_20570);
nand U27865 (N_27865,N_20295,N_21606);
nand U27866 (N_27866,N_22819,N_22748);
nand U27867 (N_27867,N_20345,N_23306);
or U27868 (N_27868,N_24959,N_21606);
nor U27869 (N_27869,N_23210,N_22088);
nand U27870 (N_27870,N_22512,N_24064);
nand U27871 (N_27871,N_23473,N_23815);
nor U27872 (N_27872,N_23052,N_22256);
or U27873 (N_27873,N_23594,N_23995);
or U27874 (N_27874,N_21577,N_20681);
nor U27875 (N_27875,N_20596,N_21694);
or U27876 (N_27876,N_22246,N_24146);
nor U27877 (N_27877,N_23779,N_23155);
nand U27878 (N_27878,N_20213,N_24304);
nor U27879 (N_27879,N_21011,N_22686);
nor U27880 (N_27880,N_23018,N_20022);
and U27881 (N_27881,N_23136,N_22516);
or U27882 (N_27882,N_23924,N_21468);
or U27883 (N_27883,N_20985,N_23531);
and U27884 (N_27884,N_24527,N_20304);
or U27885 (N_27885,N_20621,N_23035);
nand U27886 (N_27886,N_20530,N_22066);
nand U27887 (N_27887,N_22595,N_21704);
nand U27888 (N_27888,N_21098,N_22786);
or U27889 (N_27889,N_22032,N_21289);
or U27890 (N_27890,N_23369,N_20737);
nand U27891 (N_27891,N_22158,N_22939);
or U27892 (N_27892,N_24528,N_23360);
nor U27893 (N_27893,N_22454,N_20455);
and U27894 (N_27894,N_21583,N_24004);
and U27895 (N_27895,N_23324,N_23670);
nand U27896 (N_27896,N_23034,N_20882);
nor U27897 (N_27897,N_24477,N_24182);
or U27898 (N_27898,N_23112,N_21222);
or U27899 (N_27899,N_24658,N_22942);
and U27900 (N_27900,N_23034,N_22392);
or U27901 (N_27901,N_22089,N_21334);
or U27902 (N_27902,N_24101,N_24802);
and U27903 (N_27903,N_20613,N_20430);
nand U27904 (N_27904,N_22165,N_21170);
nand U27905 (N_27905,N_23559,N_23576);
or U27906 (N_27906,N_23958,N_21530);
nand U27907 (N_27907,N_22195,N_20450);
nand U27908 (N_27908,N_22932,N_23052);
nand U27909 (N_27909,N_24575,N_21749);
nor U27910 (N_27910,N_22652,N_24844);
nand U27911 (N_27911,N_23085,N_21166);
nand U27912 (N_27912,N_24616,N_22064);
or U27913 (N_27913,N_24260,N_21629);
nand U27914 (N_27914,N_20362,N_22834);
nor U27915 (N_27915,N_20892,N_24598);
and U27916 (N_27916,N_24826,N_23050);
or U27917 (N_27917,N_21947,N_22893);
nand U27918 (N_27918,N_23891,N_23284);
and U27919 (N_27919,N_23538,N_23702);
nor U27920 (N_27920,N_20481,N_24300);
and U27921 (N_27921,N_24561,N_23619);
nor U27922 (N_27922,N_23804,N_24101);
and U27923 (N_27923,N_23529,N_23172);
and U27924 (N_27924,N_22072,N_21336);
and U27925 (N_27925,N_20424,N_20296);
nor U27926 (N_27926,N_20291,N_24439);
and U27927 (N_27927,N_20580,N_24335);
or U27928 (N_27928,N_24887,N_23300);
nand U27929 (N_27929,N_21788,N_22833);
or U27930 (N_27930,N_22732,N_21160);
or U27931 (N_27931,N_23143,N_23609);
and U27932 (N_27932,N_22162,N_22329);
or U27933 (N_27933,N_23705,N_23791);
nand U27934 (N_27934,N_23146,N_23519);
and U27935 (N_27935,N_21706,N_24587);
or U27936 (N_27936,N_22801,N_22649);
or U27937 (N_27937,N_21046,N_20567);
and U27938 (N_27938,N_22010,N_22767);
nand U27939 (N_27939,N_22696,N_24269);
nor U27940 (N_27940,N_22595,N_24947);
nand U27941 (N_27941,N_24298,N_21198);
or U27942 (N_27942,N_21913,N_23751);
or U27943 (N_27943,N_24441,N_24170);
and U27944 (N_27944,N_21218,N_22489);
and U27945 (N_27945,N_22854,N_24537);
nor U27946 (N_27946,N_24573,N_21086);
and U27947 (N_27947,N_23952,N_23523);
nand U27948 (N_27948,N_21147,N_24938);
or U27949 (N_27949,N_23611,N_23432);
nand U27950 (N_27950,N_21399,N_23955);
nor U27951 (N_27951,N_23373,N_22157);
and U27952 (N_27952,N_21487,N_22063);
and U27953 (N_27953,N_22311,N_20197);
or U27954 (N_27954,N_22920,N_24996);
nand U27955 (N_27955,N_20930,N_22309);
or U27956 (N_27956,N_24962,N_22158);
nor U27957 (N_27957,N_23650,N_22903);
nand U27958 (N_27958,N_20956,N_21321);
or U27959 (N_27959,N_21086,N_24734);
nor U27960 (N_27960,N_21969,N_24110);
nand U27961 (N_27961,N_24029,N_24225);
and U27962 (N_27962,N_23326,N_22533);
or U27963 (N_27963,N_20341,N_21412);
nand U27964 (N_27964,N_20749,N_22937);
and U27965 (N_27965,N_20439,N_24609);
nand U27966 (N_27966,N_23034,N_21816);
nand U27967 (N_27967,N_22453,N_21186);
nor U27968 (N_27968,N_24382,N_20909);
or U27969 (N_27969,N_24475,N_21033);
and U27970 (N_27970,N_21285,N_24768);
and U27971 (N_27971,N_23994,N_24984);
nor U27972 (N_27972,N_24491,N_24736);
nor U27973 (N_27973,N_23431,N_21436);
and U27974 (N_27974,N_20236,N_21996);
nand U27975 (N_27975,N_21490,N_23566);
nand U27976 (N_27976,N_22890,N_21250);
or U27977 (N_27977,N_24763,N_23635);
and U27978 (N_27978,N_23499,N_20061);
xor U27979 (N_27979,N_24192,N_23323);
nand U27980 (N_27980,N_24453,N_24272);
or U27981 (N_27981,N_20227,N_22948);
or U27982 (N_27982,N_21665,N_20959);
nand U27983 (N_27983,N_24543,N_23302);
or U27984 (N_27984,N_22109,N_24834);
or U27985 (N_27985,N_24718,N_21916);
nand U27986 (N_27986,N_21120,N_24664);
nor U27987 (N_27987,N_23425,N_22151);
nor U27988 (N_27988,N_21934,N_22431);
nand U27989 (N_27989,N_23627,N_21609);
and U27990 (N_27990,N_23313,N_22684);
or U27991 (N_27991,N_20027,N_23079);
and U27992 (N_27992,N_20526,N_21658);
nand U27993 (N_27993,N_24051,N_21721);
and U27994 (N_27994,N_24414,N_20818);
and U27995 (N_27995,N_21759,N_24153);
nor U27996 (N_27996,N_23648,N_21803);
or U27997 (N_27997,N_20237,N_22891);
nand U27998 (N_27998,N_20934,N_23181);
and U27999 (N_27999,N_21998,N_21621);
nand U28000 (N_28000,N_24184,N_21369);
nand U28001 (N_28001,N_20594,N_21973);
nand U28002 (N_28002,N_20872,N_22609);
nor U28003 (N_28003,N_24290,N_23931);
nor U28004 (N_28004,N_22736,N_23832);
or U28005 (N_28005,N_20567,N_21394);
or U28006 (N_28006,N_20798,N_20065);
and U28007 (N_28007,N_21384,N_23839);
nand U28008 (N_28008,N_22284,N_24512);
nor U28009 (N_28009,N_21829,N_24098);
or U28010 (N_28010,N_21183,N_23531);
nor U28011 (N_28011,N_21334,N_23311);
and U28012 (N_28012,N_23464,N_24649);
or U28013 (N_28013,N_24316,N_23530);
nor U28014 (N_28014,N_23119,N_20687);
and U28015 (N_28015,N_20817,N_24151);
nand U28016 (N_28016,N_24372,N_22521);
or U28017 (N_28017,N_24016,N_20748);
and U28018 (N_28018,N_24179,N_22115);
or U28019 (N_28019,N_20253,N_23899);
nor U28020 (N_28020,N_21179,N_20493);
nor U28021 (N_28021,N_21713,N_23068);
nand U28022 (N_28022,N_23994,N_21684);
or U28023 (N_28023,N_21930,N_24700);
nand U28024 (N_28024,N_22855,N_24188);
nor U28025 (N_28025,N_22605,N_24577);
and U28026 (N_28026,N_24321,N_21033);
nor U28027 (N_28027,N_23127,N_21666);
and U28028 (N_28028,N_22329,N_23910);
or U28029 (N_28029,N_20530,N_22699);
or U28030 (N_28030,N_22812,N_24880);
and U28031 (N_28031,N_21346,N_22437);
or U28032 (N_28032,N_20600,N_24519);
nor U28033 (N_28033,N_22194,N_22239);
nor U28034 (N_28034,N_21932,N_20487);
nor U28035 (N_28035,N_24146,N_21790);
nor U28036 (N_28036,N_20870,N_23737);
and U28037 (N_28037,N_21884,N_24450);
nor U28038 (N_28038,N_21539,N_20205);
xor U28039 (N_28039,N_23201,N_21983);
and U28040 (N_28040,N_24271,N_24110);
nor U28041 (N_28041,N_21518,N_24655);
nand U28042 (N_28042,N_20697,N_20899);
nor U28043 (N_28043,N_22166,N_21020);
and U28044 (N_28044,N_22863,N_23071);
nor U28045 (N_28045,N_20415,N_24570);
and U28046 (N_28046,N_21382,N_23240);
and U28047 (N_28047,N_20393,N_24389);
nor U28048 (N_28048,N_21859,N_24912);
and U28049 (N_28049,N_20316,N_20496);
nand U28050 (N_28050,N_22837,N_20960);
or U28051 (N_28051,N_23795,N_23359);
nor U28052 (N_28052,N_23566,N_22855);
or U28053 (N_28053,N_24340,N_21139);
or U28054 (N_28054,N_24310,N_24349);
nor U28055 (N_28055,N_23567,N_24992);
nand U28056 (N_28056,N_22740,N_23846);
or U28057 (N_28057,N_22585,N_21181);
or U28058 (N_28058,N_22106,N_20681);
and U28059 (N_28059,N_20009,N_23568);
and U28060 (N_28060,N_23445,N_22049);
or U28061 (N_28061,N_23545,N_24837);
or U28062 (N_28062,N_23315,N_24932);
nor U28063 (N_28063,N_22901,N_23860);
nand U28064 (N_28064,N_21972,N_21316);
or U28065 (N_28065,N_23207,N_23767);
nor U28066 (N_28066,N_21992,N_21300);
or U28067 (N_28067,N_21752,N_22386);
and U28068 (N_28068,N_22745,N_23164);
nand U28069 (N_28069,N_24892,N_24451);
nor U28070 (N_28070,N_24041,N_21003);
nor U28071 (N_28071,N_20191,N_24837);
and U28072 (N_28072,N_20063,N_20655);
or U28073 (N_28073,N_23747,N_21951);
nor U28074 (N_28074,N_20423,N_24011);
or U28075 (N_28075,N_23662,N_20542);
nor U28076 (N_28076,N_24312,N_20196);
or U28077 (N_28077,N_22617,N_21628);
or U28078 (N_28078,N_24364,N_22596);
and U28079 (N_28079,N_21327,N_21570);
nor U28080 (N_28080,N_20740,N_21429);
nand U28081 (N_28081,N_20989,N_23956);
or U28082 (N_28082,N_23882,N_21045);
and U28083 (N_28083,N_20743,N_20916);
or U28084 (N_28084,N_21339,N_21625);
or U28085 (N_28085,N_20806,N_20645);
and U28086 (N_28086,N_21520,N_22372);
and U28087 (N_28087,N_20588,N_22307);
nand U28088 (N_28088,N_20568,N_20327);
or U28089 (N_28089,N_24417,N_20185);
and U28090 (N_28090,N_21858,N_23660);
nor U28091 (N_28091,N_22058,N_20573);
nor U28092 (N_28092,N_23115,N_22091);
and U28093 (N_28093,N_22032,N_20088);
nor U28094 (N_28094,N_21386,N_24836);
and U28095 (N_28095,N_24885,N_22118);
nand U28096 (N_28096,N_22177,N_20832);
and U28097 (N_28097,N_21529,N_20498);
and U28098 (N_28098,N_21958,N_22122);
nand U28099 (N_28099,N_24264,N_23589);
nand U28100 (N_28100,N_22120,N_24740);
nand U28101 (N_28101,N_23974,N_24416);
or U28102 (N_28102,N_23276,N_22887);
or U28103 (N_28103,N_24097,N_21364);
nor U28104 (N_28104,N_20246,N_24458);
and U28105 (N_28105,N_21183,N_20161);
and U28106 (N_28106,N_23855,N_21557);
and U28107 (N_28107,N_23453,N_22531);
or U28108 (N_28108,N_20699,N_24802);
and U28109 (N_28109,N_22840,N_23368);
nand U28110 (N_28110,N_20826,N_23252);
nand U28111 (N_28111,N_24135,N_22716);
nand U28112 (N_28112,N_21518,N_22581);
nor U28113 (N_28113,N_20479,N_21724);
nor U28114 (N_28114,N_20936,N_24675);
nor U28115 (N_28115,N_21239,N_22970);
nor U28116 (N_28116,N_23320,N_24969);
and U28117 (N_28117,N_23742,N_24611);
nor U28118 (N_28118,N_24013,N_22012);
nor U28119 (N_28119,N_23276,N_20921);
or U28120 (N_28120,N_20037,N_21500);
or U28121 (N_28121,N_21461,N_20565);
nor U28122 (N_28122,N_24766,N_21343);
nor U28123 (N_28123,N_24670,N_22539);
nand U28124 (N_28124,N_20902,N_24241);
nand U28125 (N_28125,N_21640,N_21468);
nor U28126 (N_28126,N_20288,N_22784);
nor U28127 (N_28127,N_20666,N_23215);
or U28128 (N_28128,N_24157,N_23978);
or U28129 (N_28129,N_21488,N_22067);
or U28130 (N_28130,N_20970,N_24097);
or U28131 (N_28131,N_22449,N_23521);
or U28132 (N_28132,N_23849,N_22102);
and U28133 (N_28133,N_22949,N_20560);
and U28134 (N_28134,N_20403,N_21285);
and U28135 (N_28135,N_22633,N_22186);
and U28136 (N_28136,N_23067,N_21747);
nor U28137 (N_28137,N_20475,N_23170);
or U28138 (N_28138,N_21459,N_20915);
and U28139 (N_28139,N_21306,N_23728);
nor U28140 (N_28140,N_22205,N_23876);
and U28141 (N_28141,N_21312,N_20314);
nand U28142 (N_28142,N_23843,N_24750);
nand U28143 (N_28143,N_24713,N_23091);
or U28144 (N_28144,N_20432,N_20379);
nand U28145 (N_28145,N_22272,N_22574);
or U28146 (N_28146,N_23299,N_22424);
nand U28147 (N_28147,N_20933,N_20441);
nor U28148 (N_28148,N_23394,N_20665);
and U28149 (N_28149,N_22036,N_23706);
and U28150 (N_28150,N_23890,N_22890);
and U28151 (N_28151,N_23035,N_20244);
nor U28152 (N_28152,N_21270,N_24249);
nor U28153 (N_28153,N_22573,N_23356);
and U28154 (N_28154,N_21868,N_23078);
and U28155 (N_28155,N_21750,N_20434);
and U28156 (N_28156,N_21404,N_24795);
nand U28157 (N_28157,N_22023,N_21677);
and U28158 (N_28158,N_22684,N_21374);
or U28159 (N_28159,N_20630,N_24789);
or U28160 (N_28160,N_23871,N_21948);
and U28161 (N_28161,N_22071,N_23458);
or U28162 (N_28162,N_24916,N_20479);
nand U28163 (N_28163,N_23180,N_21099);
and U28164 (N_28164,N_21877,N_23379);
and U28165 (N_28165,N_21932,N_24520);
or U28166 (N_28166,N_22990,N_22867);
nand U28167 (N_28167,N_24176,N_24995);
nand U28168 (N_28168,N_23292,N_20333);
nand U28169 (N_28169,N_22122,N_22834);
or U28170 (N_28170,N_23565,N_20618);
and U28171 (N_28171,N_23169,N_23907);
and U28172 (N_28172,N_22804,N_24802);
and U28173 (N_28173,N_21252,N_23882);
nand U28174 (N_28174,N_23188,N_20593);
nor U28175 (N_28175,N_21543,N_21156);
nor U28176 (N_28176,N_20948,N_24659);
or U28177 (N_28177,N_23050,N_21025);
nor U28178 (N_28178,N_22765,N_24851);
and U28179 (N_28179,N_23897,N_21910);
and U28180 (N_28180,N_20382,N_21019);
nor U28181 (N_28181,N_24353,N_23653);
nand U28182 (N_28182,N_20846,N_23480);
nand U28183 (N_28183,N_24248,N_21550);
or U28184 (N_28184,N_22440,N_23060);
nand U28185 (N_28185,N_24863,N_24441);
or U28186 (N_28186,N_23011,N_22641);
and U28187 (N_28187,N_23344,N_23984);
nand U28188 (N_28188,N_23684,N_24455);
and U28189 (N_28189,N_22028,N_21133);
nand U28190 (N_28190,N_21708,N_24871);
or U28191 (N_28191,N_22530,N_22947);
nand U28192 (N_28192,N_20734,N_21456);
or U28193 (N_28193,N_23750,N_21370);
or U28194 (N_28194,N_23245,N_23754);
and U28195 (N_28195,N_24424,N_20208);
or U28196 (N_28196,N_23077,N_22456);
or U28197 (N_28197,N_22042,N_21443);
and U28198 (N_28198,N_22145,N_22340);
nor U28199 (N_28199,N_21027,N_23441);
nand U28200 (N_28200,N_22598,N_21203);
or U28201 (N_28201,N_20018,N_20371);
nor U28202 (N_28202,N_23443,N_23434);
nor U28203 (N_28203,N_23687,N_23450);
nand U28204 (N_28204,N_21818,N_24737);
and U28205 (N_28205,N_24598,N_22270);
nor U28206 (N_28206,N_24891,N_24511);
or U28207 (N_28207,N_22346,N_21753);
nor U28208 (N_28208,N_24051,N_24018);
and U28209 (N_28209,N_20423,N_23135);
and U28210 (N_28210,N_24319,N_22391);
and U28211 (N_28211,N_23355,N_20406);
nor U28212 (N_28212,N_24697,N_21623);
or U28213 (N_28213,N_22433,N_22544);
nand U28214 (N_28214,N_24686,N_21655);
and U28215 (N_28215,N_20897,N_24658);
or U28216 (N_28216,N_23830,N_23694);
or U28217 (N_28217,N_24247,N_23019);
and U28218 (N_28218,N_21001,N_20391);
and U28219 (N_28219,N_23199,N_22251);
or U28220 (N_28220,N_24124,N_23178);
and U28221 (N_28221,N_20642,N_23211);
nor U28222 (N_28222,N_23993,N_23101);
nand U28223 (N_28223,N_24491,N_23725);
or U28224 (N_28224,N_22868,N_24616);
and U28225 (N_28225,N_21451,N_21912);
or U28226 (N_28226,N_23567,N_20090);
nand U28227 (N_28227,N_23774,N_24443);
nand U28228 (N_28228,N_20568,N_23733);
xor U28229 (N_28229,N_20859,N_22984);
or U28230 (N_28230,N_21878,N_21187);
and U28231 (N_28231,N_20794,N_20140);
nand U28232 (N_28232,N_23701,N_23366);
nor U28233 (N_28233,N_20448,N_22906);
nand U28234 (N_28234,N_20325,N_20548);
and U28235 (N_28235,N_20143,N_23751);
nor U28236 (N_28236,N_23104,N_21170);
nor U28237 (N_28237,N_23415,N_21874);
or U28238 (N_28238,N_22605,N_23313);
nand U28239 (N_28239,N_20560,N_23345);
nand U28240 (N_28240,N_22023,N_20344);
nand U28241 (N_28241,N_22811,N_22710);
and U28242 (N_28242,N_22173,N_21286);
nand U28243 (N_28243,N_20985,N_22554);
or U28244 (N_28244,N_24865,N_24898);
nor U28245 (N_28245,N_20507,N_21527);
nor U28246 (N_28246,N_20779,N_22024);
or U28247 (N_28247,N_21604,N_20354);
and U28248 (N_28248,N_24514,N_20320);
and U28249 (N_28249,N_22713,N_23641);
nor U28250 (N_28250,N_22733,N_23778);
or U28251 (N_28251,N_21955,N_23874);
and U28252 (N_28252,N_23141,N_24864);
and U28253 (N_28253,N_24862,N_22223);
nand U28254 (N_28254,N_20709,N_23395);
and U28255 (N_28255,N_22454,N_23562);
nand U28256 (N_28256,N_24227,N_24593);
and U28257 (N_28257,N_22165,N_24122);
nor U28258 (N_28258,N_21240,N_24774);
nor U28259 (N_28259,N_20439,N_21539);
nor U28260 (N_28260,N_21109,N_24933);
or U28261 (N_28261,N_23023,N_21518);
and U28262 (N_28262,N_22218,N_22961);
nor U28263 (N_28263,N_21077,N_24285);
nand U28264 (N_28264,N_20705,N_22563);
nor U28265 (N_28265,N_24897,N_23092);
nor U28266 (N_28266,N_21576,N_23997);
and U28267 (N_28267,N_21636,N_22193);
or U28268 (N_28268,N_24658,N_21867);
nand U28269 (N_28269,N_23968,N_24176);
or U28270 (N_28270,N_24724,N_24002);
nor U28271 (N_28271,N_21515,N_23883);
nand U28272 (N_28272,N_20166,N_23557);
nor U28273 (N_28273,N_21051,N_23515);
nor U28274 (N_28274,N_24354,N_22688);
nand U28275 (N_28275,N_23844,N_21827);
and U28276 (N_28276,N_24719,N_20411);
nor U28277 (N_28277,N_23372,N_22564);
or U28278 (N_28278,N_23306,N_22268);
and U28279 (N_28279,N_22027,N_22666);
and U28280 (N_28280,N_24616,N_23516);
nand U28281 (N_28281,N_22155,N_22019);
nor U28282 (N_28282,N_23119,N_20288);
and U28283 (N_28283,N_20797,N_23175);
nor U28284 (N_28284,N_21154,N_20328);
or U28285 (N_28285,N_20017,N_24628);
nand U28286 (N_28286,N_24656,N_22503);
nand U28287 (N_28287,N_22653,N_24387);
nand U28288 (N_28288,N_23940,N_22293);
nor U28289 (N_28289,N_21341,N_20951);
nor U28290 (N_28290,N_20170,N_20078);
or U28291 (N_28291,N_23999,N_20388);
nand U28292 (N_28292,N_21846,N_24775);
and U28293 (N_28293,N_20559,N_23858);
nor U28294 (N_28294,N_20659,N_20160);
or U28295 (N_28295,N_21618,N_22147);
nor U28296 (N_28296,N_21964,N_22413);
or U28297 (N_28297,N_21510,N_20356);
nor U28298 (N_28298,N_21746,N_22880);
nor U28299 (N_28299,N_23930,N_21655);
and U28300 (N_28300,N_23492,N_22761);
nand U28301 (N_28301,N_20559,N_23177);
nor U28302 (N_28302,N_24907,N_24178);
and U28303 (N_28303,N_22134,N_22412);
nand U28304 (N_28304,N_23530,N_24487);
and U28305 (N_28305,N_23845,N_24185);
and U28306 (N_28306,N_23832,N_22345);
nand U28307 (N_28307,N_24964,N_22584);
or U28308 (N_28308,N_24693,N_21907);
or U28309 (N_28309,N_20103,N_23219);
or U28310 (N_28310,N_20736,N_24246);
nor U28311 (N_28311,N_23923,N_21265);
or U28312 (N_28312,N_22321,N_20460);
or U28313 (N_28313,N_20570,N_21233);
nor U28314 (N_28314,N_21860,N_23633);
nand U28315 (N_28315,N_22573,N_24320);
or U28316 (N_28316,N_22672,N_21322);
and U28317 (N_28317,N_23496,N_21443);
or U28318 (N_28318,N_20628,N_23851);
or U28319 (N_28319,N_21727,N_22840);
and U28320 (N_28320,N_22758,N_20341);
or U28321 (N_28321,N_21723,N_22342);
or U28322 (N_28322,N_24859,N_22546);
nand U28323 (N_28323,N_20382,N_22324);
or U28324 (N_28324,N_20456,N_23630);
or U28325 (N_28325,N_22924,N_23322);
and U28326 (N_28326,N_21721,N_22010);
or U28327 (N_28327,N_22360,N_24714);
nor U28328 (N_28328,N_23321,N_22774);
nor U28329 (N_28329,N_21628,N_22205);
nor U28330 (N_28330,N_24089,N_24667);
or U28331 (N_28331,N_22416,N_22230);
or U28332 (N_28332,N_21716,N_21916);
and U28333 (N_28333,N_20109,N_22772);
and U28334 (N_28334,N_24261,N_23223);
and U28335 (N_28335,N_23800,N_20560);
and U28336 (N_28336,N_23081,N_23725);
nand U28337 (N_28337,N_23169,N_24569);
and U28338 (N_28338,N_21763,N_23606);
nor U28339 (N_28339,N_20170,N_20382);
and U28340 (N_28340,N_21400,N_21561);
and U28341 (N_28341,N_24079,N_24283);
and U28342 (N_28342,N_24439,N_20350);
or U28343 (N_28343,N_22222,N_21800);
or U28344 (N_28344,N_23702,N_20132);
or U28345 (N_28345,N_22413,N_22398);
nor U28346 (N_28346,N_23341,N_23138);
and U28347 (N_28347,N_20703,N_20232);
or U28348 (N_28348,N_22575,N_21989);
nor U28349 (N_28349,N_20301,N_21832);
or U28350 (N_28350,N_23222,N_20203);
nand U28351 (N_28351,N_23553,N_21225);
nor U28352 (N_28352,N_21455,N_23176);
nor U28353 (N_28353,N_22731,N_22977);
and U28354 (N_28354,N_21342,N_20392);
or U28355 (N_28355,N_23271,N_20023);
nor U28356 (N_28356,N_24091,N_22122);
and U28357 (N_28357,N_24430,N_24432);
nor U28358 (N_28358,N_23895,N_20282);
nand U28359 (N_28359,N_23416,N_22536);
nor U28360 (N_28360,N_24944,N_23830);
nand U28361 (N_28361,N_22253,N_22561);
nor U28362 (N_28362,N_24317,N_20357);
and U28363 (N_28363,N_20227,N_24558);
nand U28364 (N_28364,N_21874,N_20639);
and U28365 (N_28365,N_23771,N_22444);
or U28366 (N_28366,N_23119,N_24437);
or U28367 (N_28367,N_23823,N_24390);
nand U28368 (N_28368,N_21821,N_20094);
and U28369 (N_28369,N_22989,N_21560);
or U28370 (N_28370,N_24340,N_24330);
or U28371 (N_28371,N_21174,N_24308);
nand U28372 (N_28372,N_22283,N_24971);
or U28373 (N_28373,N_21120,N_22346);
and U28374 (N_28374,N_20959,N_21356);
and U28375 (N_28375,N_20877,N_20771);
xnor U28376 (N_28376,N_23147,N_22729);
or U28377 (N_28377,N_21175,N_23945);
nor U28378 (N_28378,N_24727,N_24179);
or U28379 (N_28379,N_22967,N_24793);
and U28380 (N_28380,N_23554,N_20378);
nor U28381 (N_28381,N_22705,N_24189);
nand U28382 (N_28382,N_24814,N_21043);
nor U28383 (N_28383,N_20337,N_24687);
or U28384 (N_28384,N_24034,N_24316);
nor U28385 (N_28385,N_23104,N_20286);
or U28386 (N_28386,N_23292,N_24099);
and U28387 (N_28387,N_24667,N_22890);
nand U28388 (N_28388,N_24258,N_22308);
or U28389 (N_28389,N_23340,N_23649);
or U28390 (N_28390,N_24427,N_20553);
and U28391 (N_28391,N_22136,N_21812);
nor U28392 (N_28392,N_24411,N_20890);
nor U28393 (N_28393,N_20126,N_21786);
nand U28394 (N_28394,N_23275,N_22220);
nand U28395 (N_28395,N_21611,N_23939);
nor U28396 (N_28396,N_24844,N_24246);
or U28397 (N_28397,N_24604,N_24822);
and U28398 (N_28398,N_21001,N_22507);
or U28399 (N_28399,N_20533,N_24833);
or U28400 (N_28400,N_23934,N_20106);
nor U28401 (N_28401,N_22337,N_22792);
and U28402 (N_28402,N_24979,N_22702);
or U28403 (N_28403,N_24534,N_20794);
and U28404 (N_28404,N_23525,N_21114);
or U28405 (N_28405,N_21868,N_24900);
nand U28406 (N_28406,N_20083,N_22709);
nand U28407 (N_28407,N_20627,N_23621);
or U28408 (N_28408,N_21243,N_20876);
nor U28409 (N_28409,N_23050,N_22435);
and U28410 (N_28410,N_20464,N_20541);
nand U28411 (N_28411,N_21071,N_21252);
nor U28412 (N_28412,N_22457,N_23428);
and U28413 (N_28413,N_21890,N_22541);
nor U28414 (N_28414,N_24723,N_22241);
nor U28415 (N_28415,N_24340,N_24873);
and U28416 (N_28416,N_20215,N_22140);
and U28417 (N_28417,N_23281,N_24987);
and U28418 (N_28418,N_20728,N_23841);
nand U28419 (N_28419,N_22028,N_23937);
and U28420 (N_28420,N_20321,N_22699);
and U28421 (N_28421,N_21220,N_21024);
nand U28422 (N_28422,N_21487,N_20881);
nor U28423 (N_28423,N_21678,N_23705);
xor U28424 (N_28424,N_24266,N_22872);
nor U28425 (N_28425,N_21146,N_20560);
nor U28426 (N_28426,N_23031,N_24459);
or U28427 (N_28427,N_23564,N_23464);
and U28428 (N_28428,N_22159,N_23525);
or U28429 (N_28429,N_22550,N_22040);
or U28430 (N_28430,N_20277,N_21664);
and U28431 (N_28431,N_23419,N_23878);
and U28432 (N_28432,N_24182,N_22901);
nor U28433 (N_28433,N_23725,N_21202);
nor U28434 (N_28434,N_20525,N_21403);
and U28435 (N_28435,N_22272,N_21761);
nand U28436 (N_28436,N_21871,N_20026);
nand U28437 (N_28437,N_24594,N_23495);
nor U28438 (N_28438,N_22521,N_20246);
nand U28439 (N_28439,N_23725,N_21646);
nand U28440 (N_28440,N_22521,N_24129);
nand U28441 (N_28441,N_22230,N_23512);
and U28442 (N_28442,N_21075,N_21499);
nand U28443 (N_28443,N_22141,N_20285);
and U28444 (N_28444,N_24985,N_23565);
nand U28445 (N_28445,N_22156,N_21560);
or U28446 (N_28446,N_23377,N_22382);
nand U28447 (N_28447,N_22991,N_20257);
nand U28448 (N_28448,N_23997,N_24604);
or U28449 (N_28449,N_22749,N_24215);
nand U28450 (N_28450,N_20238,N_22667);
nand U28451 (N_28451,N_21735,N_21028);
and U28452 (N_28452,N_20750,N_20814);
and U28453 (N_28453,N_24433,N_22498);
nor U28454 (N_28454,N_21306,N_23316);
and U28455 (N_28455,N_21232,N_22072);
and U28456 (N_28456,N_22824,N_23219);
nor U28457 (N_28457,N_24753,N_22284);
nor U28458 (N_28458,N_23047,N_22863);
xnor U28459 (N_28459,N_23246,N_22673);
and U28460 (N_28460,N_23128,N_24467);
or U28461 (N_28461,N_21816,N_24762);
nand U28462 (N_28462,N_23717,N_24364);
nand U28463 (N_28463,N_22283,N_23478);
or U28464 (N_28464,N_21302,N_20644);
nand U28465 (N_28465,N_22824,N_21799);
nand U28466 (N_28466,N_20890,N_23981);
and U28467 (N_28467,N_24072,N_24038);
and U28468 (N_28468,N_21449,N_21731);
nor U28469 (N_28469,N_22470,N_20193);
or U28470 (N_28470,N_20535,N_20009);
nor U28471 (N_28471,N_24657,N_23827);
nand U28472 (N_28472,N_20355,N_20029);
nor U28473 (N_28473,N_22669,N_23018);
nand U28474 (N_28474,N_24974,N_24542);
or U28475 (N_28475,N_22153,N_22075);
nand U28476 (N_28476,N_22447,N_20506);
or U28477 (N_28477,N_21186,N_23831);
nor U28478 (N_28478,N_22166,N_22332);
nor U28479 (N_28479,N_22469,N_22110);
and U28480 (N_28480,N_21386,N_22163);
nor U28481 (N_28481,N_24770,N_21419);
nor U28482 (N_28482,N_21661,N_21870);
and U28483 (N_28483,N_21558,N_24092);
nand U28484 (N_28484,N_21667,N_22004);
and U28485 (N_28485,N_23187,N_20334);
or U28486 (N_28486,N_23099,N_23758);
nand U28487 (N_28487,N_21042,N_20034);
nand U28488 (N_28488,N_23108,N_22004);
nor U28489 (N_28489,N_20304,N_24775);
or U28490 (N_28490,N_22494,N_21712);
nand U28491 (N_28491,N_21237,N_24895);
and U28492 (N_28492,N_21660,N_20786);
or U28493 (N_28493,N_21940,N_24903);
nor U28494 (N_28494,N_21694,N_21356);
nor U28495 (N_28495,N_20353,N_20389);
nor U28496 (N_28496,N_22241,N_24731);
and U28497 (N_28497,N_22046,N_24745);
nand U28498 (N_28498,N_22289,N_23738);
nor U28499 (N_28499,N_21894,N_21310);
nor U28500 (N_28500,N_21667,N_22752);
nor U28501 (N_28501,N_23422,N_20731);
nor U28502 (N_28502,N_21320,N_22406);
and U28503 (N_28503,N_22035,N_22750);
nor U28504 (N_28504,N_22212,N_23551);
nor U28505 (N_28505,N_24252,N_23169);
or U28506 (N_28506,N_20902,N_22424);
or U28507 (N_28507,N_24266,N_20728);
nand U28508 (N_28508,N_21709,N_21833);
nand U28509 (N_28509,N_23806,N_22451);
nand U28510 (N_28510,N_24694,N_23941);
or U28511 (N_28511,N_24353,N_23062);
nor U28512 (N_28512,N_22075,N_24418);
nor U28513 (N_28513,N_20946,N_24912);
nor U28514 (N_28514,N_24067,N_24966);
nor U28515 (N_28515,N_21785,N_23760);
or U28516 (N_28516,N_22401,N_23794);
or U28517 (N_28517,N_22005,N_23857);
xor U28518 (N_28518,N_23875,N_22851);
nand U28519 (N_28519,N_20297,N_22844);
and U28520 (N_28520,N_21282,N_20483);
and U28521 (N_28521,N_23836,N_22874);
or U28522 (N_28522,N_23124,N_24653);
nand U28523 (N_28523,N_23831,N_22668);
and U28524 (N_28524,N_24908,N_20237);
or U28525 (N_28525,N_21511,N_22931);
or U28526 (N_28526,N_24727,N_24659);
nor U28527 (N_28527,N_23838,N_21201);
nor U28528 (N_28528,N_21610,N_23198);
nor U28529 (N_28529,N_24140,N_21343);
nor U28530 (N_28530,N_24802,N_20910);
nor U28531 (N_28531,N_23693,N_21071);
nor U28532 (N_28532,N_23370,N_22579);
and U28533 (N_28533,N_23732,N_20860);
xor U28534 (N_28534,N_23127,N_20608);
nand U28535 (N_28535,N_21892,N_23333);
nor U28536 (N_28536,N_24268,N_22196);
and U28537 (N_28537,N_23691,N_21717);
or U28538 (N_28538,N_21504,N_23777);
and U28539 (N_28539,N_21074,N_23772);
nor U28540 (N_28540,N_23598,N_22488);
nor U28541 (N_28541,N_20619,N_22571);
or U28542 (N_28542,N_21973,N_21438);
or U28543 (N_28543,N_20297,N_20507);
nand U28544 (N_28544,N_24446,N_24766);
nand U28545 (N_28545,N_22951,N_22744);
nand U28546 (N_28546,N_23559,N_23641);
or U28547 (N_28547,N_24447,N_24377);
nand U28548 (N_28548,N_22437,N_24616);
nand U28549 (N_28549,N_23741,N_20447);
and U28550 (N_28550,N_24786,N_22825);
and U28551 (N_28551,N_22769,N_22759);
nand U28552 (N_28552,N_21725,N_23779);
nor U28553 (N_28553,N_24547,N_24695);
nor U28554 (N_28554,N_21881,N_22173);
and U28555 (N_28555,N_21532,N_21486);
or U28556 (N_28556,N_20952,N_22012);
nor U28557 (N_28557,N_21049,N_21096);
or U28558 (N_28558,N_20346,N_20585);
nand U28559 (N_28559,N_23867,N_21848);
and U28560 (N_28560,N_21841,N_20962);
or U28561 (N_28561,N_22221,N_24872);
and U28562 (N_28562,N_20167,N_24792);
and U28563 (N_28563,N_24427,N_24963);
nand U28564 (N_28564,N_21199,N_21205);
xor U28565 (N_28565,N_20441,N_22460);
nor U28566 (N_28566,N_20397,N_20183);
and U28567 (N_28567,N_22139,N_20474);
or U28568 (N_28568,N_20619,N_24122);
and U28569 (N_28569,N_24620,N_21368);
or U28570 (N_28570,N_22469,N_24167);
and U28571 (N_28571,N_20922,N_24835);
or U28572 (N_28572,N_21219,N_23370);
and U28573 (N_28573,N_21015,N_22686);
nor U28574 (N_28574,N_20469,N_22883);
or U28575 (N_28575,N_20211,N_20300);
xor U28576 (N_28576,N_21550,N_22752);
or U28577 (N_28577,N_22935,N_20273);
nand U28578 (N_28578,N_23769,N_20365);
and U28579 (N_28579,N_23450,N_22540);
nand U28580 (N_28580,N_21160,N_20903);
nor U28581 (N_28581,N_24188,N_23893);
nor U28582 (N_28582,N_22257,N_24009);
or U28583 (N_28583,N_24609,N_24508);
or U28584 (N_28584,N_21113,N_23667);
nor U28585 (N_28585,N_22458,N_22478);
or U28586 (N_28586,N_24560,N_22028);
and U28587 (N_28587,N_20964,N_21759);
nand U28588 (N_28588,N_21385,N_20161);
and U28589 (N_28589,N_23778,N_23150);
and U28590 (N_28590,N_20228,N_23646);
and U28591 (N_28591,N_22649,N_21373);
nor U28592 (N_28592,N_22336,N_22676);
or U28593 (N_28593,N_22340,N_23487);
nor U28594 (N_28594,N_23394,N_20413);
nor U28595 (N_28595,N_23318,N_23921);
or U28596 (N_28596,N_20714,N_20273);
nor U28597 (N_28597,N_22617,N_20487);
nor U28598 (N_28598,N_23147,N_24715);
and U28599 (N_28599,N_23876,N_20444);
or U28600 (N_28600,N_22183,N_20380);
nor U28601 (N_28601,N_24951,N_22851);
and U28602 (N_28602,N_20892,N_21760);
or U28603 (N_28603,N_24515,N_21434);
nor U28604 (N_28604,N_20282,N_24854);
nor U28605 (N_28605,N_20650,N_21225);
nor U28606 (N_28606,N_24771,N_21117);
xor U28607 (N_28607,N_23959,N_20833);
nor U28608 (N_28608,N_24371,N_24071);
nand U28609 (N_28609,N_22046,N_21347);
or U28610 (N_28610,N_23021,N_23053);
nor U28611 (N_28611,N_23153,N_22349);
or U28612 (N_28612,N_23749,N_21013);
nor U28613 (N_28613,N_21083,N_20586);
nand U28614 (N_28614,N_20384,N_22098);
and U28615 (N_28615,N_20522,N_23347);
nand U28616 (N_28616,N_23152,N_20349);
and U28617 (N_28617,N_22673,N_20168);
or U28618 (N_28618,N_22218,N_22081);
nand U28619 (N_28619,N_22490,N_24841);
and U28620 (N_28620,N_21474,N_21037);
nand U28621 (N_28621,N_23292,N_22365);
or U28622 (N_28622,N_21782,N_23451);
xnor U28623 (N_28623,N_22425,N_22592);
nor U28624 (N_28624,N_22459,N_22133);
nand U28625 (N_28625,N_21232,N_21585);
nor U28626 (N_28626,N_22218,N_23553);
nor U28627 (N_28627,N_23120,N_21175);
nand U28628 (N_28628,N_24477,N_23542);
nor U28629 (N_28629,N_22359,N_22429);
nor U28630 (N_28630,N_20563,N_20417);
and U28631 (N_28631,N_22566,N_21187);
nor U28632 (N_28632,N_23199,N_24659);
nand U28633 (N_28633,N_20853,N_21569);
nor U28634 (N_28634,N_24294,N_24877);
nor U28635 (N_28635,N_22148,N_24834);
nand U28636 (N_28636,N_21728,N_22298);
and U28637 (N_28637,N_21104,N_20201);
or U28638 (N_28638,N_22367,N_20282);
nor U28639 (N_28639,N_22016,N_23855);
nand U28640 (N_28640,N_24312,N_23879);
nand U28641 (N_28641,N_22570,N_23928);
nand U28642 (N_28642,N_22821,N_21237);
xor U28643 (N_28643,N_23963,N_21585);
and U28644 (N_28644,N_22687,N_24511);
or U28645 (N_28645,N_22076,N_20114);
and U28646 (N_28646,N_24081,N_22641);
and U28647 (N_28647,N_23842,N_22325);
and U28648 (N_28648,N_23744,N_22411);
nor U28649 (N_28649,N_22130,N_21659);
nand U28650 (N_28650,N_24041,N_20513);
nand U28651 (N_28651,N_23110,N_22974);
or U28652 (N_28652,N_20902,N_21123);
nand U28653 (N_28653,N_21488,N_24603);
or U28654 (N_28654,N_23299,N_21809);
and U28655 (N_28655,N_22920,N_22188);
and U28656 (N_28656,N_23019,N_20966);
and U28657 (N_28657,N_21201,N_22264);
or U28658 (N_28658,N_20522,N_21482);
or U28659 (N_28659,N_20681,N_22851);
or U28660 (N_28660,N_24074,N_20044);
and U28661 (N_28661,N_22233,N_22779);
or U28662 (N_28662,N_22732,N_22079);
nor U28663 (N_28663,N_23832,N_20054);
and U28664 (N_28664,N_20454,N_22035);
xor U28665 (N_28665,N_21911,N_20390);
nand U28666 (N_28666,N_24369,N_20534);
nor U28667 (N_28667,N_21002,N_22002);
xnor U28668 (N_28668,N_24526,N_22598);
and U28669 (N_28669,N_23903,N_23726);
nor U28670 (N_28670,N_23646,N_22384);
nor U28671 (N_28671,N_21164,N_24397);
or U28672 (N_28672,N_24599,N_21932);
and U28673 (N_28673,N_20806,N_21507);
xnor U28674 (N_28674,N_23868,N_24012);
nor U28675 (N_28675,N_20941,N_24173);
and U28676 (N_28676,N_23818,N_24718);
or U28677 (N_28677,N_22680,N_24833);
or U28678 (N_28678,N_22414,N_21616);
or U28679 (N_28679,N_20289,N_23800);
or U28680 (N_28680,N_24410,N_22121);
nor U28681 (N_28681,N_23883,N_22449);
nor U28682 (N_28682,N_22574,N_21741);
nor U28683 (N_28683,N_21662,N_21568);
nor U28684 (N_28684,N_23559,N_23337);
nand U28685 (N_28685,N_23268,N_23053);
and U28686 (N_28686,N_23673,N_23666);
xor U28687 (N_28687,N_20102,N_23075);
nand U28688 (N_28688,N_22049,N_24149);
nand U28689 (N_28689,N_23364,N_21797);
nand U28690 (N_28690,N_24516,N_24667);
or U28691 (N_28691,N_24047,N_24214);
and U28692 (N_28692,N_24499,N_23941);
and U28693 (N_28693,N_23941,N_22896);
and U28694 (N_28694,N_22248,N_21238);
nand U28695 (N_28695,N_24135,N_22999);
nor U28696 (N_28696,N_24920,N_24202);
or U28697 (N_28697,N_23299,N_20338);
and U28698 (N_28698,N_22822,N_23754);
xnor U28699 (N_28699,N_23700,N_20286);
and U28700 (N_28700,N_23989,N_23145);
or U28701 (N_28701,N_21912,N_21124);
nand U28702 (N_28702,N_20049,N_24997);
nor U28703 (N_28703,N_20221,N_23438);
and U28704 (N_28704,N_21544,N_22567);
nand U28705 (N_28705,N_21778,N_24850);
nor U28706 (N_28706,N_22180,N_21335);
or U28707 (N_28707,N_24867,N_23662);
nand U28708 (N_28708,N_22398,N_22462);
or U28709 (N_28709,N_24718,N_21119);
or U28710 (N_28710,N_21839,N_20708);
nand U28711 (N_28711,N_20694,N_24386);
nor U28712 (N_28712,N_22648,N_21130);
nor U28713 (N_28713,N_22153,N_23333);
and U28714 (N_28714,N_21840,N_20602);
nor U28715 (N_28715,N_24357,N_21838);
nor U28716 (N_28716,N_20855,N_20470);
and U28717 (N_28717,N_21712,N_23180);
or U28718 (N_28718,N_22331,N_22128);
or U28719 (N_28719,N_23182,N_21965);
or U28720 (N_28720,N_22969,N_22600);
nand U28721 (N_28721,N_24400,N_21240);
or U28722 (N_28722,N_23408,N_23329);
nor U28723 (N_28723,N_24001,N_22156);
xor U28724 (N_28724,N_24829,N_22780);
or U28725 (N_28725,N_23174,N_23780);
nand U28726 (N_28726,N_23133,N_22348);
and U28727 (N_28727,N_22937,N_23979);
nor U28728 (N_28728,N_23969,N_21414);
or U28729 (N_28729,N_23042,N_21396);
nor U28730 (N_28730,N_21872,N_23121);
or U28731 (N_28731,N_20031,N_24230);
and U28732 (N_28732,N_20499,N_24333);
nor U28733 (N_28733,N_24450,N_22539);
nand U28734 (N_28734,N_24344,N_22157);
or U28735 (N_28735,N_24301,N_22841);
nor U28736 (N_28736,N_24014,N_22924);
nand U28737 (N_28737,N_24449,N_22845);
or U28738 (N_28738,N_23818,N_24721);
and U28739 (N_28739,N_20112,N_24176);
nor U28740 (N_28740,N_23297,N_22270);
or U28741 (N_28741,N_21312,N_20713);
nand U28742 (N_28742,N_22409,N_21417);
or U28743 (N_28743,N_21360,N_21754);
nor U28744 (N_28744,N_22368,N_22305);
and U28745 (N_28745,N_23106,N_23424);
nand U28746 (N_28746,N_24939,N_23002);
or U28747 (N_28747,N_20018,N_21770);
and U28748 (N_28748,N_24140,N_22607);
nand U28749 (N_28749,N_24814,N_20574);
nor U28750 (N_28750,N_23998,N_24769);
nand U28751 (N_28751,N_23493,N_24779);
and U28752 (N_28752,N_24493,N_24783);
nor U28753 (N_28753,N_24296,N_21661);
and U28754 (N_28754,N_22605,N_22414);
or U28755 (N_28755,N_22034,N_23732);
and U28756 (N_28756,N_24700,N_21225);
or U28757 (N_28757,N_24624,N_24032);
or U28758 (N_28758,N_22192,N_22529);
or U28759 (N_28759,N_23467,N_21041);
and U28760 (N_28760,N_22389,N_20934);
or U28761 (N_28761,N_23803,N_22809);
nand U28762 (N_28762,N_24534,N_21143);
or U28763 (N_28763,N_23090,N_22262);
or U28764 (N_28764,N_21914,N_24982);
or U28765 (N_28765,N_24254,N_23701);
nand U28766 (N_28766,N_20627,N_21788);
xor U28767 (N_28767,N_24299,N_22358);
nor U28768 (N_28768,N_23240,N_24276);
and U28769 (N_28769,N_21309,N_22076);
and U28770 (N_28770,N_23059,N_21904);
nand U28771 (N_28771,N_23550,N_22635);
nor U28772 (N_28772,N_21828,N_24929);
or U28773 (N_28773,N_20698,N_24906);
and U28774 (N_28774,N_24863,N_20034);
nor U28775 (N_28775,N_24293,N_20574);
nor U28776 (N_28776,N_22977,N_22992);
or U28777 (N_28777,N_22651,N_23949);
and U28778 (N_28778,N_23010,N_22836);
nand U28779 (N_28779,N_21414,N_23187);
nand U28780 (N_28780,N_23826,N_21841);
or U28781 (N_28781,N_20787,N_23379);
and U28782 (N_28782,N_22622,N_20909);
nand U28783 (N_28783,N_24954,N_22091);
xnor U28784 (N_28784,N_22818,N_22510);
and U28785 (N_28785,N_24219,N_23360);
nand U28786 (N_28786,N_21617,N_22447);
or U28787 (N_28787,N_22414,N_24371);
nor U28788 (N_28788,N_20181,N_20374);
and U28789 (N_28789,N_23902,N_20340);
nor U28790 (N_28790,N_21407,N_23813);
nor U28791 (N_28791,N_22219,N_24192);
nand U28792 (N_28792,N_23473,N_24882);
nor U28793 (N_28793,N_21364,N_23009);
nand U28794 (N_28794,N_20850,N_20680);
nand U28795 (N_28795,N_21431,N_24983);
or U28796 (N_28796,N_21013,N_23251);
nand U28797 (N_28797,N_22108,N_23979);
nor U28798 (N_28798,N_23831,N_21230);
nand U28799 (N_28799,N_24855,N_22905);
and U28800 (N_28800,N_23286,N_22068);
nor U28801 (N_28801,N_20254,N_20070);
nor U28802 (N_28802,N_22934,N_24002);
nand U28803 (N_28803,N_22210,N_24659);
nor U28804 (N_28804,N_21269,N_24793);
nand U28805 (N_28805,N_20072,N_23985);
nand U28806 (N_28806,N_23721,N_22414);
nor U28807 (N_28807,N_22843,N_21802);
or U28808 (N_28808,N_24180,N_20263);
nand U28809 (N_28809,N_24850,N_21086);
and U28810 (N_28810,N_20392,N_21402);
nor U28811 (N_28811,N_21553,N_21325);
nand U28812 (N_28812,N_22726,N_23876);
and U28813 (N_28813,N_24451,N_20127);
and U28814 (N_28814,N_24297,N_23439);
and U28815 (N_28815,N_21647,N_22528);
and U28816 (N_28816,N_23987,N_22011);
and U28817 (N_28817,N_20798,N_20232);
or U28818 (N_28818,N_23039,N_22721);
nand U28819 (N_28819,N_22872,N_22398);
or U28820 (N_28820,N_21515,N_21120);
and U28821 (N_28821,N_23302,N_23494);
or U28822 (N_28822,N_22380,N_23035);
and U28823 (N_28823,N_21667,N_22828);
nand U28824 (N_28824,N_24272,N_24986);
and U28825 (N_28825,N_20945,N_20488);
nor U28826 (N_28826,N_23054,N_21260);
nor U28827 (N_28827,N_24037,N_21792);
nor U28828 (N_28828,N_22441,N_20709);
and U28829 (N_28829,N_23989,N_23225);
xnor U28830 (N_28830,N_24354,N_23868);
nor U28831 (N_28831,N_24599,N_21193);
or U28832 (N_28832,N_24134,N_20571);
and U28833 (N_28833,N_23901,N_21792);
or U28834 (N_28834,N_23692,N_20288);
nand U28835 (N_28835,N_23193,N_20413);
nor U28836 (N_28836,N_23187,N_20674);
or U28837 (N_28837,N_22951,N_23708);
nor U28838 (N_28838,N_23226,N_22254);
or U28839 (N_28839,N_24311,N_24631);
and U28840 (N_28840,N_24931,N_23353);
nand U28841 (N_28841,N_24909,N_24224);
and U28842 (N_28842,N_20132,N_22138);
nand U28843 (N_28843,N_20066,N_23050);
or U28844 (N_28844,N_23628,N_21139);
or U28845 (N_28845,N_22237,N_23767);
and U28846 (N_28846,N_23701,N_20859);
or U28847 (N_28847,N_20136,N_23022);
nor U28848 (N_28848,N_24677,N_24983);
nor U28849 (N_28849,N_22218,N_20062);
or U28850 (N_28850,N_20770,N_22039);
or U28851 (N_28851,N_21702,N_20060);
and U28852 (N_28852,N_21350,N_22556);
nand U28853 (N_28853,N_21945,N_20680);
or U28854 (N_28854,N_22030,N_22538);
nand U28855 (N_28855,N_24567,N_24472);
or U28856 (N_28856,N_21058,N_23632);
and U28857 (N_28857,N_20741,N_22439);
nand U28858 (N_28858,N_22836,N_22091);
and U28859 (N_28859,N_23936,N_22697);
nor U28860 (N_28860,N_22407,N_24501);
nor U28861 (N_28861,N_21140,N_24657);
nor U28862 (N_28862,N_20818,N_24235);
nor U28863 (N_28863,N_20353,N_24443);
nor U28864 (N_28864,N_24973,N_21854);
and U28865 (N_28865,N_20986,N_23087);
nand U28866 (N_28866,N_24554,N_22642);
and U28867 (N_28867,N_23856,N_20375);
nor U28868 (N_28868,N_21094,N_23112);
nand U28869 (N_28869,N_24823,N_20233);
or U28870 (N_28870,N_20037,N_21760);
nor U28871 (N_28871,N_22709,N_23062);
or U28872 (N_28872,N_23465,N_20001);
and U28873 (N_28873,N_22686,N_20250);
nor U28874 (N_28874,N_23487,N_21236);
nor U28875 (N_28875,N_24843,N_20684);
and U28876 (N_28876,N_24322,N_20912);
nand U28877 (N_28877,N_21525,N_24783);
or U28878 (N_28878,N_20772,N_20765);
or U28879 (N_28879,N_24337,N_24906);
or U28880 (N_28880,N_23791,N_21961);
nand U28881 (N_28881,N_23080,N_22090);
and U28882 (N_28882,N_22812,N_24586);
nor U28883 (N_28883,N_24579,N_20395);
and U28884 (N_28884,N_23202,N_24740);
nand U28885 (N_28885,N_22898,N_24759);
nor U28886 (N_28886,N_23636,N_21342);
and U28887 (N_28887,N_20812,N_23999);
and U28888 (N_28888,N_20676,N_20289);
nand U28889 (N_28889,N_21618,N_21806);
or U28890 (N_28890,N_21532,N_20075);
and U28891 (N_28891,N_21711,N_24231);
nor U28892 (N_28892,N_20284,N_20527);
or U28893 (N_28893,N_24575,N_24854);
nor U28894 (N_28894,N_22776,N_24379);
nand U28895 (N_28895,N_21680,N_24086);
nor U28896 (N_28896,N_24291,N_23498);
and U28897 (N_28897,N_24730,N_22361);
nor U28898 (N_28898,N_20985,N_24572);
and U28899 (N_28899,N_24064,N_20874);
and U28900 (N_28900,N_24525,N_22808);
nor U28901 (N_28901,N_24905,N_23103);
nand U28902 (N_28902,N_21020,N_22091);
nor U28903 (N_28903,N_21407,N_20099);
and U28904 (N_28904,N_22237,N_23175);
nand U28905 (N_28905,N_20074,N_22899);
and U28906 (N_28906,N_20870,N_24729);
and U28907 (N_28907,N_20412,N_24062);
and U28908 (N_28908,N_20094,N_23055);
nand U28909 (N_28909,N_21812,N_22252);
and U28910 (N_28910,N_20274,N_22231);
or U28911 (N_28911,N_23219,N_24926);
and U28912 (N_28912,N_20844,N_22629);
and U28913 (N_28913,N_20753,N_24118);
and U28914 (N_28914,N_22082,N_20662);
nor U28915 (N_28915,N_20306,N_23797);
or U28916 (N_28916,N_22531,N_22681);
or U28917 (N_28917,N_23149,N_23051);
nand U28918 (N_28918,N_24167,N_20227);
nor U28919 (N_28919,N_21183,N_22655);
nand U28920 (N_28920,N_24064,N_24090);
or U28921 (N_28921,N_22732,N_21050);
and U28922 (N_28922,N_21815,N_23748);
and U28923 (N_28923,N_24781,N_24902);
nor U28924 (N_28924,N_20935,N_23012);
and U28925 (N_28925,N_21707,N_20959);
or U28926 (N_28926,N_20003,N_22790);
or U28927 (N_28927,N_23817,N_21653);
nor U28928 (N_28928,N_24527,N_21784);
nor U28929 (N_28929,N_21710,N_21720);
and U28930 (N_28930,N_21226,N_22830);
nand U28931 (N_28931,N_20346,N_24126);
and U28932 (N_28932,N_22616,N_21857);
nand U28933 (N_28933,N_22179,N_22315);
and U28934 (N_28934,N_22420,N_20569);
nor U28935 (N_28935,N_24402,N_22841);
nor U28936 (N_28936,N_21415,N_20568);
nand U28937 (N_28937,N_20500,N_23922);
nand U28938 (N_28938,N_24847,N_21518);
nor U28939 (N_28939,N_24748,N_23713);
nor U28940 (N_28940,N_24033,N_23824);
nor U28941 (N_28941,N_22204,N_24516);
xor U28942 (N_28942,N_20665,N_20652);
or U28943 (N_28943,N_22505,N_22562);
and U28944 (N_28944,N_20060,N_24953);
nor U28945 (N_28945,N_21427,N_22155);
nand U28946 (N_28946,N_22522,N_23522);
nor U28947 (N_28947,N_21542,N_21800);
nand U28948 (N_28948,N_20807,N_20030);
nor U28949 (N_28949,N_21866,N_24011);
and U28950 (N_28950,N_22183,N_21722);
or U28951 (N_28951,N_23091,N_23020);
or U28952 (N_28952,N_22975,N_23069);
xor U28953 (N_28953,N_24767,N_21716);
and U28954 (N_28954,N_20239,N_22948);
and U28955 (N_28955,N_24191,N_21540);
nand U28956 (N_28956,N_21861,N_22626);
nand U28957 (N_28957,N_23905,N_20988);
and U28958 (N_28958,N_22812,N_24888);
or U28959 (N_28959,N_21725,N_24822);
nand U28960 (N_28960,N_23211,N_23879);
or U28961 (N_28961,N_20979,N_23428);
nand U28962 (N_28962,N_20318,N_24646);
nor U28963 (N_28963,N_20222,N_20986);
or U28964 (N_28964,N_23942,N_20025);
nor U28965 (N_28965,N_22894,N_22185);
nand U28966 (N_28966,N_23758,N_24612);
nor U28967 (N_28967,N_22447,N_20249);
nand U28968 (N_28968,N_23048,N_22393);
nor U28969 (N_28969,N_20482,N_24080);
nand U28970 (N_28970,N_21334,N_21011);
or U28971 (N_28971,N_23851,N_24379);
nand U28972 (N_28972,N_24542,N_20304);
xor U28973 (N_28973,N_20325,N_22747);
or U28974 (N_28974,N_24405,N_24875);
nor U28975 (N_28975,N_20856,N_22873);
nor U28976 (N_28976,N_22984,N_21154);
and U28977 (N_28977,N_20739,N_20186);
nand U28978 (N_28978,N_24758,N_23883);
nor U28979 (N_28979,N_24346,N_22839);
nor U28980 (N_28980,N_21091,N_22050);
and U28981 (N_28981,N_21561,N_24485);
nor U28982 (N_28982,N_21581,N_24635);
nand U28983 (N_28983,N_22565,N_22442);
and U28984 (N_28984,N_20081,N_21148);
nand U28985 (N_28985,N_23647,N_23721);
or U28986 (N_28986,N_20591,N_21841);
nor U28987 (N_28987,N_21589,N_24713);
nor U28988 (N_28988,N_20005,N_22435);
nand U28989 (N_28989,N_23696,N_24516);
nor U28990 (N_28990,N_24855,N_24863);
nand U28991 (N_28991,N_21677,N_20028);
or U28992 (N_28992,N_22662,N_22478);
and U28993 (N_28993,N_22575,N_20536);
and U28994 (N_28994,N_23865,N_20157);
xor U28995 (N_28995,N_23399,N_24863);
nor U28996 (N_28996,N_22582,N_23955);
or U28997 (N_28997,N_21249,N_23755);
and U28998 (N_28998,N_22692,N_23312);
nor U28999 (N_28999,N_21572,N_21188);
or U29000 (N_29000,N_21463,N_23751);
or U29001 (N_29001,N_23512,N_23681);
nor U29002 (N_29002,N_24551,N_20298);
nand U29003 (N_29003,N_24892,N_20941);
and U29004 (N_29004,N_20683,N_22932);
nand U29005 (N_29005,N_23074,N_21998);
nand U29006 (N_29006,N_20364,N_21624);
nor U29007 (N_29007,N_21330,N_23600);
nor U29008 (N_29008,N_21678,N_23633);
nand U29009 (N_29009,N_20673,N_23324);
or U29010 (N_29010,N_20346,N_22170);
nand U29011 (N_29011,N_24008,N_24750);
nand U29012 (N_29012,N_22658,N_24923);
xnor U29013 (N_29013,N_21532,N_20137);
nand U29014 (N_29014,N_23326,N_23776);
nand U29015 (N_29015,N_20383,N_23967);
and U29016 (N_29016,N_24168,N_20608);
nor U29017 (N_29017,N_20083,N_23778);
and U29018 (N_29018,N_20997,N_22157);
nor U29019 (N_29019,N_23126,N_20700);
nor U29020 (N_29020,N_21386,N_23582);
nand U29021 (N_29021,N_21393,N_22688);
nor U29022 (N_29022,N_23481,N_23110);
nand U29023 (N_29023,N_22721,N_20159);
nand U29024 (N_29024,N_21214,N_20362);
nor U29025 (N_29025,N_21638,N_22623);
or U29026 (N_29026,N_24391,N_24051);
or U29027 (N_29027,N_24867,N_23053);
and U29028 (N_29028,N_20032,N_22429);
and U29029 (N_29029,N_22928,N_20595);
and U29030 (N_29030,N_21650,N_24783);
nor U29031 (N_29031,N_23512,N_22691);
and U29032 (N_29032,N_23746,N_23229);
and U29033 (N_29033,N_23641,N_22086);
and U29034 (N_29034,N_22570,N_22247);
nand U29035 (N_29035,N_20085,N_21930);
nand U29036 (N_29036,N_22321,N_23981);
nand U29037 (N_29037,N_23890,N_22741);
nand U29038 (N_29038,N_22183,N_23321);
and U29039 (N_29039,N_20403,N_21995);
and U29040 (N_29040,N_24351,N_20113);
and U29041 (N_29041,N_24022,N_22935);
nand U29042 (N_29042,N_22768,N_23146);
nor U29043 (N_29043,N_20325,N_23691);
nand U29044 (N_29044,N_21188,N_21148);
nor U29045 (N_29045,N_22115,N_21751);
nand U29046 (N_29046,N_24796,N_23314);
or U29047 (N_29047,N_23127,N_20419);
nand U29048 (N_29048,N_20600,N_24673);
nand U29049 (N_29049,N_24219,N_22029);
or U29050 (N_29050,N_20210,N_23533);
or U29051 (N_29051,N_22404,N_21458);
and U29052 (N_29052,N_23470,N_22246);
nor U29053 (N_29053,N_22410,N_24791);
and U29054 (N_29054,N_20293,N_22096);
nand U29055 (N_29055,N_24214,N_21178);
nand U29056 (N_29056,N_21010,N_21839);
or U29057 (N_29057,N_23395,N_23447);
nand U29058 (N_29058,N_22542,N_24245);
nand U29059 (N_29059,N_24392,N_22188);
and U29060 (N_29060,N_21313,N_24935);
nor U29061 (N_29061,N_20223,N_22767);
and U29062 (N_29062,N_22500,N_22432);
and U29063 (N_29063,N_24483,N_22161);
nand U29064 (N_29064,N_24713,N_24691);
or U29065 (N_29065,N_20613,N_23176);
and U29066 (N_29066,N_23874,N_22428);
nor U29067 (N_29067,N_21322,N_23860);
nand U29068 (N_29068,N_22809,N_21562);
and U29069 (N_29069,N_23170,N_20452);
nor U29070 (N_29070,N_23955,N_24711);
nand U29071 (N_29071,N_23329,N_23835);
nor U29072 (N_29072,N_24373,N_21178);
nor U29073 (N_29073,N_22840,N_23619);
and U29074 (N_29074,N_20794,N_24289);
nor U29075 (N_29075,N_20248,N_20770);
and U29076 (N_29076,N_20952,N_23698);
nand U29077 (N_29077,N_23039,N_21612);
nor U29078 (N_29078,N_23000,N_22448);
nor U29079 (N_29079,N_24710,N_21715);
and U29080 (N_29080,N_23918,N_20910);
and U29081 (N_29081,N_20822,N_24684);
and U29082 (N_29082,N_22700,N_20038);
or U29083 (N_29083,N_21952,N_22002);
or U29084 (N_29084,N_20055,N_21506);
nand U29085 (N_29085,N_24707,N_22456);
nand U29086 (N_29086,N_23402,N_21245);
or U29087 (N_29087,N_22601,N_21384);
nor U29088 (N_29088,N_21911,N_21673);
and U29089 (N_29089,N_20554,N_21996);
and U29090 (N_29090,N_20475,N_24963);
nor U29091 (N_29091,N_24313,N_22618);
and U29092 (N_29092,N_21189,N_24344);
or U29093 (N_29093,N_24748,N_23836);
or U29094 (N_29094,N_21343,N_21748);
nor U29095 (N_29095,N_20033,N_22626);
nand U29096 (N_29096,N_21030,N_23721);
or U29097 (N_29097,N_24143,N_24947);
and U29098 (N_29098,N_20696,N_22349);
nor U29099 (N_29099,N_23499,N_23735);
nand U29100 (N_29100,N_24725,N_24507);
or U29101 (N_29101,N_24213,N_24722);
or U29102 (N_29102,N_24476,N_21577);
or U29103 (N_29103,N_20787,N_24769);
and U29104 (N_29104,N_24221,N_21801);
and U29105 (N_29105,N_20372,N_21738);
nor U29106 (N_29106,N_24808,N_20882);
xnor U29107 (N_29107,N_21317,N_21981);
nand U29108 (N_29108,N_21252,N_23213);
or U29109 (N_29109,N_22624,N_24835);
and U29110 (N_29110,N_22176,N_23878);
and U29111 (N_29111,N_23641,N_24868);
nor U29112 (N_29112,N_20823,N_23631);
nand U29113 (N_29113,N_21747,N_20009);
and U29114 (N_29114,N_22860,N_24088);
and U29115 (N_29115,N_21105,N_23810);
or U29116 (N_29116,N_21911,N_23947);
and U29117 (N_29117,N_21705,N_23026);
and U29118 (N_29118,N_24668,N_22810);
nand U29119 (N_29119,N_21088,N_23013);
nor U29120 (N_29120,N_23229,N_23683);
or U29121 (N_29121,N_20113,N_23835);
nand U29122 (N_29122,N_23948,N_20491);
nand U29123 (N_29123,N_21175,N_23807);
or U29124 (N_29124,N_24977,N_24217);
nor U29125 (N_29125,N_21411,N_22063);
and U29126 (N_29126,N_23957,N_24860);
nand U29127 (N_29127,N_20826,N_20870);
xor U29128 (N_29128,N_24529,N_23258);
or U29129 (N_29129,N_23062,N_20106);
nand U29130 (N_29130,N_22708,N_23078);
or U29131 (N_29131,N_24982,N_24769);
or U29132 (N_29132,N_20040,N_20716);
nor U29133 (N_29133,N_21168,N_20342);
nor U29134 (N_29134,N_22987,N_23592);
nand U29135 (N_29135,N_21683,N_22285);
and U29136 (N_29136,N_22969,N_21731);
and U29137 (N_29137,N_21817,N_20787);
nand U29138 (N_29138,N_21427,N_23541);
or U29139 (N_29139,N_21742,N_24238);
nand U29140 (N_29140,N_21645,N_24131);
and U29141 (N_29141,N_22385,N_23252);
nand U29142 (N_29142,N_23857,N_24084);
nor U29143 (N_29143,N_24491,N_24940);
or U29144 (N_29144,N_24138,N_22575);
nand U29145 (N_29145,N_22892,N_23830);
nand U29146 (N_29146,N_24036,N_21128);
nor U29147 (N_29147,N_24526,N_24970);
nor U29148 (N_29148,N_24688,N_22287);
and U29149 (N_29149,N_21437,N_23297);
nand U29150 (N_29150,N_21460,N_23927);
or U29151 (N_29151,N_22387,N_21441);
and U29152 (N_29152,N_20624,N_22562);
nor U29153 (N_29153,N_20305,N_21174);
and U29154 (N_29154,N_21730,N_24870);
nor U29155 (N_29155,N_24484,N_23486);
or U29156 (N_29156,N_23630,N_22572);
nor U29157 (N_29157,N_22427,N_21846);
and U29158 (N_29158,N_21234,N_24911);
and U29159 (N_29159,N_22415,N_22559);
or U29160 (N_29160,N_21718,N_22772);
nand U29161 (N_29161,N_24460,N_21528);
and U29162 (N_29162,N_22409,N_23836);
nand U29163 (N_29163,N_21404,N_24949);
or U29164 (N_29164,N_21745,N_22498);
nor U29165 (N_29165,N_24136,N_20095);
nand U29166 (N_29166,N_22217,N_24695);
and U29167 (N_29167,N_20581,N_24882);
nand U29168 (N_29168,N_23868,N_24472);
and U29169 (N_29169,N_24363,N_23626);
nor U29170 (N_29170,N_22508,N_23101);
and U29171 (N_29171,N_23080,N_23735);
xor U29172 (N_29172,N_21148,N_20208);
or U29173 (N_29173,N_23992,N_20073);
and U29174 (N_29174,N_23933,N_24285);
nor U29175 (N_29175,N_24919,N_20271);
nor U29176 (N_29176,N_22284,N_23316);
nor U29177 (N_29177,N_24501,N_24395);
or U29178 (N_29178,N_21996,N_23699);
nor U29179 (N_29179,N_22675,N_22199);
and U29180 (N_29180,N_21146,N_20440);
nor U29181 (N_29181,N_21968,N_21350);
or U29182 (N_29182,N_20795,N_24871);
or U29183 (N_29183,N_21532,N_24834);
nand U29184 (N_29184,N_20875,N_22806);
or U29185 (N_29185,N_24644,N_20542);
or U29186 (N_29186,N_22225,N_22582);
nand U29187 (N_29187,N_21473,N_21555);
nand U29188 (N_29188,N_20326,N_24645);
nor U29189 (N_29189,N_23337,N_20191);
or U29190 (N_29190,N_23039,N_20816);
and U29191 (N_29191,N_24063,N_24097);
nand U29192 (N_29192,N_24692,N_23649);
nor U29193 (N_29193,N_22780,N_22474);
and U29194 (N_29194,N_22442,N_22504);
nand U29195 (N_29195,N_22074,N_21713);
nor U29196 (N_29196,N_20170,N_21300);
nand U29197 (N_29197,N_23431,N_24795);
nor U29198 (N_29198,N_23256,N_22798);
and U29199 (N_29199,N_23911,N_22459);
nor U29200 (N_29200,N_21791,N_24405);
nand U29201 (N_29201,N_23083,N_23768);
or U29202 (N_29202,N_24498,N_21792);
nand U29203 (N_29203,N_20528,N_22539);
nor U29204 (N_29204,N_22561,N_21489);
nand U29205 (N_29205,N_20650,N_21689);
nor U29206 (N_29206,N_23788,N_21962);
nor U29207 (N_29207,N_23671,N_22844);
nand U29208 (N_29208,N_22411,N_20678);
nor U29209 (N_29209,N_22485,N_22431);
and U29210 (N_29210,N_20600,N_23434);
and U29211 (N_29211,N_22661,N_22685);
and U29212 (N_29212,N_22023,N_24489);
nand U29213 (N_29213,N_20188,N_21464);
nor U29214 (N_29214,N_23006,N_20946);
nor U29215 (N_29215,N_21921,N_23932);
nor U29216 (N_29216,N_24125,N_20584);
or U29217 (N_29217,N_23103,N_23758);
nand U29218 (N_29218,N_23384,N_20913);
nor U29219 (N_29219,N_20056,N_23107);
nand U29220 (N_29220,N_20908,N_20712);
or U29221 (N_29221,N_23322,N_21599);
or U29222 (N_29222,N_24026,N_21932);
or U29223 (N_29223,N_24044,N_23606);
nor U29224 (N_29224,N_20799,N_20033);
or U29225 (N_29225,N_22916,N_24985);
and U29226 (N_29226,N_24445,N_22453);
and U29227 (N_29227,N_21689,N_24806);
and U29228 (N_29228,N_22780,N_20943);
and U29229 (N_29229,N_22796,N_23368);
nand U29230 (N_29230,N_24388,N_23322);
or U29231 (N_29231,N_22873,N_24363);
nand U29232 (N_29232,N_20193,N_20530);
nand U29233 (N_29233,N_20028,N_23294);
or U29234 (N_29234,N_24500,N_22692);
nand U29235 (N_29235,N_22337,N_22338);
or U29236 (N_29236,N_20379,N_24664);
or U29237 (N_29237,N_21111,N_24339);
or U29238 (N_29238,N_24124,N_20445);
and U29239 (N_29239,N_20572,N_21059);
nor U29240 (N_29240,N_22386,N_20507);
or U29241 (N_29241,N_23005,N_23441);
nand U29242 (N_29242,N_20677,N_23367);
nand U29243 (N_29243,N_20915,N_22501);
nand U29244 (N_29244,N_24807,N_21749);
nor U29245 (N_29245,N_22148,N_22188);
nor U29246 (N_29246,N_21176,N_23068);
nand U29247 (N_29247,N_21129,N_20593);
nand U29248 (N_29248,N_21564,N_21279);
and U29249 (N_29249,N_24575,N_24369);
nor U29250 (N_29250,N_22359,N_24321);
nor U29251 (N_29251,N_24487,N_20085);
nor U29252 (N_29252,N_22090,N_20891);
nand U29253 (N_29253,N_20375,N_21102);
or U29254 (N_29254,N_22036,N_20559);
or U29255 (N_29255,N_21624,N_21180);
nand U29256 (N_29256,N_24787,N_23473);
and U29257 (N_29257,N_20153,N_24601);
nor U29258 (N_29258,N_22512,N_24408);
or U29259 (N_29259,N_20606,N_24334);
and U29260 (N_29260,N_22531,N_22202);
nand U29261 (N_29261,N_22256,N_21202);
nand U29262 (N_29262,N_21068,N_20032);
or U29263 (N_29263,N_21678,N_20923);
and U29264 (N_29264,N_20727,N_20144);
nand U29265 (N_29265,N_20687,N_23041);
nor U29266 (N_29266,N_23801,N_24032);
nor U29267 (N_29267,N_20905,N_22635);
and U29268 (N_29268,N_21584,N_23590);
xor U29269 (N_29269,N_22129,N_24901);
and U29270 (N_29270,N_22886,N_21951);
nand U29271 (N_29271,N_22382,N_22969);
nand U29272 (N_29272,N_23006,N_21777);
nor U29273 (N_29273,N_23021,N_23766);
or U29274 (N_29274,N_23674,N_21336);
and U29275 (N_29275,N_24738,N_23287);
nand U29276 (N_29276,N_22134,N_22714);
nor U29277 (N_29277,N_20705,N_24487);
nand U29278 (N_29278,N_21944,N_21015);
and U29279 (N_29279,N_21077,N_23354);
and U29280 (N_29280,N_24558,N_24169);
nand U29281 (N_29281,N_24771,N_24355);
nor U29282 (N_29282,N_21023,N_23379);
nor U29283 (N_29283,N_22608,N_23973);
nand U29284 (N_29284,N_24375,N_22215);
nor U29285 (N_29285,N_23464,N_24987);
and U29286 (N_29286,N_20003,N_24412);
and U29287 (N_29287,N_20975,N_22647);
nor U29288 (N_29288,N_21892,N_23762);
nor U29289 (N_29289,N_22901,N_23501);
nor U29290 (N_29290,N_20569,N_21145);
or U29291 (N_29291,N_21702,N_24999);
nor U29292 (N_29292,N_22207,N_23434);
or U29293 (N_29293,N_24188,N_24072);
nor U29294 (N_29294,N_23190,N_22251);
nand U29295 (N_29295,N_24132,N_23767);
and U29296 (N_29296,N_22485,N_20588);
and U29297 (N_29297,N_22860,N_24380);
and U29298 (N_29298,N_24355,N_24738);
and U29299 (N_29299,N_24755,N_20903);
and U29300 (N_29300,N_21338,N_24146);
and U29301 (N_29301,N_23850,N_24392);
nand U29302 (N_29302,N_24496,N_24396);
or U29303 (N_29303,N_21327,N_21263);
nand U29304 (N_29304,N_24899,N_24906);
and U29305 (N_29305,N_21506,N_23276);
and U29306 (N_29306,N_23094,N_22180);
and U29307 (N_29307,N_22187,N_21957);
nor U29308 (N_29308,N_23258,N_22705);
or U29309 (N_29309,N_23133,N_20470);
nand U29310 (N_29310,N_22110,N_20549);
and U29311 (N_29311,N_24966,N_24382);
and U29312 (N_29312,N_21659,N_22224);
xnor U29313 (N_29313,N_23912,N_21457);
and U29314 (N_29314,N_21155,N_20533);
and U29315 (N_29315,N_22024,N_22085);
nor U29316 (N_29316,N_21531,N_22919);
nand U29317 (N_29317,N_23158,N_24470);
or U29318 (N_29318,N_21379,N_20423);
or U29319 (N_29319,N_20032,N_24045);
nor U29320 (N_29320,N_24688,N_22727);
and U29321 (N_29321,N_21101,N_22796);
and U29322 (N_29322,N_24322,N_22802);
nor U29323 (N_29323,N_23344,N_21050);
and U29324 (N_29324,N_21889,N_21395);
nand U29325 (N_29325,N_24445,N_22288);
nand U29326 (N_29326,N_24855,N_21121);
nand U29327 (N_29327,N_20799,N_21165);
and U29328 (N_29328,N_22586,N_20177);
nor U29329 (N_29329,N_23582,N_21205);
and U29330 (N_29330,N_21014,N_20470);
or U29331 (N_29331,N_23258,N_22720);
or U29332 (N_29332,N_20837,N_24881);
and U29333 (N_29333,N_23226,N_24245);
or U29334 (N_29334,N_21736,N_22825);
nor U29335 (N_29335,N_20247,N_22276);
nor U29336 (N_29336,N_23887,N_23254);
and U29337 (N_29337,N_20424,N_22664);
nor U29338 (N_29338,N_24245,N_23154);
nor U29339 (N_29339,N_23995,N_24262);
nor U29340 (N_29340,N_24632,N_21814);
or U29341 (N_29341,N_21085,N_20907);
and U29342 (N_29342,N_20671,N_21446);
and U29343 (N_29343,N_22236,N_20009);
nor U29344 (N_29344,N_22683,N_22366);
nand U29345 (N_29345,N_22150,N_22078);
nor U29346 (N_29346,N_21404,N_21691);
or U29347 (N_29347,N_23341,N_23077);
nand U29348 (N_29348,N_22389,N_23294);
nor U29349 (N_29349,N_21461,N_21235);
nor U29350 (N_29350,N_22031,N_20462);
nand U29351 (N_29351,N_20382,N_24945);
nand U29352 (N_29352,N_20854,N_23173);
nand U29353 (N_29353,N_20034,N_24936);
and U29354 (N_29354,N_23957,N_23388);
nand U29355 (N_29355,N_23833,N_24503);
nand U29356 (N_29356,N_23686,N_21782);
nand U29357 (N_29357,N_24157,N_22865);
nand U29358 (N_29358,N_22888,N_24918);
nor U29359 (N_29359,N_22760,N_21549);
nor U29360 (N_29360,N_20792,N_22784);
or U29361 (N_29361,N_23158,N_23741);
nand U29362 (N_29362,N_20372,N_21076);
nor U29363 (N_29363,N_24251,N_24989);
nand U29364 (N_29364,N_22330,N_20927);
and U29365 (N_29365,N_22203,N_24169);
or U29366 (N_29366,N_22404,N_22109);
nand U29367 (N_29367,N_21044,N_20371);
nor U29368 (N_29368,N_22173,N_24206);
nor U29369 (N_29369,N_20198,N_21983);
nand U29370 (N_29370,N_23551,N_21960);
nand U29371 (N_29371,N_23497,N_20102);
nand U29372 (N_29372,N_22622,N_20920);
nor U29373 (N_29373,N_21508,N_24445);
nand U29374 (N_29374,N_21548,N_22311);
nand U29375 (N_29375,N_23021,N_23343);
and U29376 (N_29376,N_22196,N_20412);
nand U29377 (N_29377,N_21890,N_20009);
and U29378 (N_29378,N_23303,N_24952);
or U29379 (N_29379,N_22973,N_23141);
nand U29380 (N_29380,N_20312,N_21651);
or U29381 (N_29381,N_23853,N_24842);
and U29382 (N_29382,N_23656,N_23734);
nor U29383 (N_29383,N_24209,N_24667);
or U29384 (N_29384,N_21680,N_20911);
or U29385 (N_29385,N_20791,N_20251);
and U29386 (N_29386,N_22654,N_22966);
nor U29387 (N_29387,N_22632,N_21039);
or U29388 (N_29388,N_21486,N_23197);
and U29389 (N_29389,N_22878,N_23248);
or U29390 (N_29390,N_21298,N_20748);
and U29391 (N_29391,N_21385,N_24094);
nor U29392 (N_29392,N_22520,N_24465);
nor U29393 (N_29393,N_20539,N_22508);
and U29394 (N_29394,N_24231,N_24912);
nor U29395 (N_29395,N_20226,N_21892);
and U29396 (N_29396,N_22053,N_21555);
or U29397 (N_29397,N_20715,N_20373);
or U29398 (N_29398,N_23756,N_24227);
and U29399 (N_29399,N_21840,N_23702);
nor U29400 (N_29400,N_24042,N_24804);
nand U29401 (N_29401,N_21020,N_24038);
or U29402 (N_29402,N_23219,N_23718);
and U29403 (N_29403,N_20130,N_24128);
or U29404 (N_29404,N_23066,N_23030);
or U29405 (N_29405,N_23967,N_22275);
nor U29406 (N_29406,N_20052,N_20059);
nand U29407 (N_29407,N_21570,N_22243);
nand U29408 (N_29408,N_21597,N_20780);
or U29409 (N_29409,N_24536,N_23802);
nor U29410 (N_29410,N_22103,N_22116);
or U29411 (N_29411,N_24285,N_24394);
nand U29412 (N_29412,N_22987,N_22706);
and U29413 (N_29413,N_24759,N_24078);
and U29414 (N_29414,N_22785,N_20976);
or U29415 (N_29415,N_20928,N_20789);
nor U29416 (N_29416,N_21576,N_24395);
nor U29417 (N_29417,N_24669,N_20015);
or U29418 (N_29418,N_24634,N_22154);
and U29419 (N_29419,N_23422,N_22366);
and U29420 (N_29420,N_22542,N_21882);
or U29421 (N_29421,N_24906,N_21215);
or U29422 (N_29422,N_20518,N_22089);
nor U29423 (N_29423,N_24565,N_24514);
nand U29424 (N_29424,N_20002,N_21644);
and U29425 (N_29425,N_21301,N_20559);
nor U29426 (N_29426,N_23868,N_21407);
and U29427 (N_29427,N_24450,N_20149);
and U29428 (N_29428,N_24964,N_21232);
and U29429 (N_29429,N_23446,N_20743);
nand U29430 (N_29430,N_23418,N_23615);
or U29431 (N_29431,N_23203,N_23488);
nand U29432 (N_29432,N_21001,N_24773);
nor U29433 (N_29433,N_24585,N_20144);
nand U29434 (N_29434,N_20781,N_24736);
or U29435 (N_29435,N_21301,N_20457);
nor U29436 (N_29436,N_24057,N_20976);
nand U29437 (N_29437,N_22771,N_20150);
xor U29438 (N_29438,N_20238,N_20733);
and U29439 (N_29439,N_22488,N_22934);
nor U29440 (N_29440,N_20807,N_20160);
nand U29441 (N_29441,N_23580,N_22742);
nand U29442 (N_29442,N_21737,N_24132);
nor U29443 (N_29443,N_21959,N_22491);
nor U29444 (N_29444,N_23448,N_23311);
or U29445 (N_29445,N_20512,N_23902);
or U29446 (N_29446,N_20289,N_22927);
nor U29447 (N_29447,N_20557,N_23436);
nand U29448 (N_29448,N_21272,N_22136);
nand U29449 (N_29449,N_21870,N_21505);
nor U29450 (N_29450,N_21388,N_22646);
nand U29451 (N_29451,N_21747,N_24902);
nand U29452 (N_29452,N_24582,N_20626);
nor U29453 (N_29453,N_20726,N_22828);
nor U29454 (N_29454,N_24791,N_23990);
and U29455 (N_29455,N_20077,N_23121);
and U29456 (N_29456,N_21134,N_22869);
nand U29457 (N_29457,N_22449,N_23597);
nor U29458 (N_29458,N_21351,N_20579);
or U29459 (N_29459,N_23321,N_23561);
nor U29460 (N_29460,N_21673,N_20659);
nand U29461 (N_29461,N_24880,N_23171);
and U29462 (N_29462,N_21621,N_22696);
and U29463 (N_29463,N_23474,N_22553);
and U29464 (N_29464,N_20193,N_21169);
nor U29465 (N_29465,N_21400,N_23318);
or U29466 (N_29466,N_20395,N_22506);
xor U29467 (N_29467,N_20097,N_21953);
nor U29468 (N_29468,N_24962,N_21113);
and U29469 (N_29469,N_24615,N_21185);
or U29470 (N_29470,N_23785,N_23758);
and U29471 (N_29471,N_24527,N_23678);
nor U29472 (N_29472,N_23217,N_21451);
nor U29473 (N_29473,N_20583,N_20092);
and U29474 (N_29474,N_23666,N_24428);
or U29475 (N_29475,N_22241,N_24140);
nor U29476 (N_29476,N_21978,N_23436);
nand U29477 (N_29477,N_23979,N_23777);
and U29478 (N_29478,N_20075,N_24434);
or U29479 (N_29479,N_20490,N_20619);
nor U29480 (N_29480,N_20897,N_24344);
and U29481 (N_29481,N_23490,N_24718);
nand U29482 (N_29482,N_24616,N_22330);
nor U29483 (N_29483,N_20798,N_21817);
nand U29484 (N_29484,N_22145,N_20460);
nand U29485 (N_29485,N_23692,N_22550);
nor U29486 (N_29486,N_20809,N_23047);
and U29487 (N_29487,N_20271,N_21779);
and U29488 (N_29488,N_24044,N_23642);
and U29489 (N_29489,N_24922,N_20666);
or U29490 (N_29490,N_23943,N_21540);
nor U29491 (N_29491,N_23211,N_24209);
or U29492 (N_29492,N_24829,N_22159);
and U29493 (N_29493,N_20082,N_20254);
and U29494 (N_29494,N_24220,N_21503);
xor U29495 (N_29495,N_21819,N_23388);
or U29496 (N_29496,N_22721,N_24106);
or U29497 (N_29497,N_21461,N_23741);
or U29498 (N_29498,N_23393,N_22472);
and U29499 (N_29499,N_20661,N_20877);
nand U29500 (N_29500,N_21682,N_23446);
xnor U29501 (N_29501,N_21470,N_22477);
nand U29502 (N_29502,N_21907,N_20711);
and U29503 (N_29503,N_21557,N_21970);
or U29504 (N_29504,N_20061,N_24315);
and U29505 (N_29505,N_20586,N_23928);
and U29506 (N_29506,N_20099,N_22411);
or U29507 (N_29507,N_23401,N_21243);
or U29508 (N_29508,N_21391,N_24498);
or U29509 (N_29509,N_22310,N_23511);
nand U29510 (N_29510,N_21915,N_20028);
nand U29511 (N_29511,N_21252,N_24508);
nor U29512 (N_29512,N_24538,N_20519);
nand U29513 (N_29513,N_20301,N_24699);
or U29514 (N_29514,N_22999,N_23445);
nand U29515 (N_29515,N_24753,N_20407);
or U29516 (N_29516,N_21989,N_21103);
nand U29517 (N_29517,N_21227,N_21920);
or U29518 (N_29518,N_23750,N_24224);
nor U29519 (N_29519,N_23520,N_21967);
nand U29520 (N_29520,N_22846,N_24415);
nor U29521 (N_29521,N_20800,N_23604);
nand U29522 (N_29522,N_23021,N_20075);
or U29523 (N_29523,N_23324,N_23716);
and U29524 (N_29524,N_23418,N_23831);
and U29525 (N_29525,N_20865,N_20863);
and U29526 (N_29526,N_20808,N_24496);
nand U29527 (N_29527,N_21414,N_22672);
or U29528 (N_29528,N_21138,N_24365);
or U29529 (N_29529,N_20547,N_24190);
nand U29530 (N_29530,N_20579,N_22431);
nand U29531 (N_29531,N_20559,N_22862);
nand U29532 (N_29532,N_23190,N_20058);
nand U29533 (N_29533,N_20209,N_20233);
nand U29534 (N_29534,N_20731,N_22421);
and U29535 (N_29535,N_23354,N_21474);
and U29536 (N_29536,N_24035,N_22639);
nand U29537 (N_29537,N_21683,N_20155);
nand U29538 (N_29538,N_24930,N_21027);
nand U29539 (N_29539,N_22477,N_24082);
and U29540 (N_29540,N_22721,N_20588);
nor U29541 (N_29541,N_24088,N_24972);
nand U29542 (N_29542,N_21777,N_23456);
or U29543 (N_29543,N_23619,N_23509);
or U29544 (N_29544,N_24099,N_22251);
nor U29545 (N_29545,N_23392,N_23633);
nand U29546 (N_29546,N_24664,N_21574);
nand U29547 (N_29547,N_23396,N_21679);
and U29548 (N_29548,N_20283,N_24041);
nand U29549 (N_29549,N_22500,N_22084);
nand U29550 (N_29550,N_24483,N_22471);
or U29551 (N_29551,N_21630,N_21229);
nand U29552 (N_29552,N_23164,N_22641);
nand U29553 (N_29553,N_22505,N_23706);
nand U29554 (N_29554,N_24629,N_24565);
or U29555 (N_29555,N_22633,N_24290);
nand U29556 (N_29556,N_21839,N_23963);
and U29557 (N_29557,N_21986,N_22243);
and U29558 (N_29558,N_22608,N_24569);
nand U29559 (N_29559,N_20720,N_20669);
and U29560 (N_29560,N_20238,N_21515);
nor U29561 (N_29561,N_23662,N_23212);
nand U29562 (N_29562,N_20926,N_22226);
or U29563 (N_29563,N_24755,N_21224);
and U29564 (N_29564,N_24278,N_22739);
and U29565 (N_29565,N_22293,N_22554);
or U29566 (N_29566,N_24173,N_23417);
nor U29567 (N_29567,N_22244,N_20567);
nand U29568 (N_29568,N_20079,N_22034);
nor U29569 (N_29569,N_24713,N_20585);
nor U29570 (N_29570,N_24248,N_23492);
and U29571 (N_29571,N_21431,N_22900);
or U29572 (N_29572,N_20816,N_21290);
nand U29573 (N_29573,N_21134,N_21201);
and U29574 (N_29574,N_24118,N_24319);
or U29575 (N_29575,N_21056,N_22255);
nor U29576 (N_29576,N_24147,N_20257);
and U29577 (N_29577,N_20974,N_22117);
nand U29578 (N_29578,N_22562,N_22339);
nand U29579 (N_29579,N_20080,N_23283);
or U29580 (N_29580,N_24645,N_23279);
nand U29581 (N_29581,N_24415,N_20393);
nor U29582 (N_29582,N_20755,N_22702);
nor U29583 (N_29583,N_21237,N_21902);
or U29584 (N_29584,N_24848,N_22752);
and U29585 (N_29585,N_22152,N_20945);
nand U29586 (N_29586,N_20579,N_22963);
and U29587 (N_29587,N_22300,N_20749);
nor U29588 (N_29588,N_23808,N_24709);
or U29589 (N_29589,N_22213,N_22825);
nand U29590 (N_29590,N_24353,N_21718);
and U29591 (N_29591,N_22744,N_20990);
nor U29592 (N_29592,N_24638,N_20314);
and U29593 (N_29593,N_24881,N_23748);
and U29594 (N_29594,N_24748,N_24299);
and U29595 (N_29595,N_22264,N_20347);
or U29596 (N_29596,N_20250,N_24250);
nor U29597 (N_29597,N_20680,N_24967);
nor U29598 (N_29598,N_24150,N_22867);
nor U29599 (N_29599,N_21408,N_24467);
nor U29600 (N_29600,N_22240,N_23979);
or U29601 (N_29601,N_20200,N_20915);
or U29602 (N_29602,N_20812,N_20387);
and U29603 (N_29603,N_20711,N_23265);
or U29604 (N_29604,N_20659,N_23704);
nand U29605 (N_29605,N_22639,N_20363);
nand U29606 (N_29606,N_23614,N_21044);
or U29607 (N_29607,N_20749,N_20096);
or U29608 (N_29608,N_20150,N_22159);
and U29609 (N_29609,N_20550,N_24504);
and U29610 (N_29610,N_22278,N_23537);
nand U29611 (N_29611,N_23162,N_23419);
nor U29612 (N_29612,N_24227,N_20956);
and U29613 (N_29613,N_23636,N_24818);
and U29614 (N_29614,N_24766,N_24421);
or U29615 (N_29615,N_22554,N_20756);
nand U29616 (N_29616,N_24162,N_23052);
nor U29617 (N_29617,N_20753,N_21060);
nor U29618 (N_29618,N_24924,N_22886);
nor U29619 (N_29619,N_20212,N_23349);
nand U29620 (N_29620,N_24455,N_22239);
xor U29621 (N_29621,N_24345,N_23617);
or U29622 (N_29622,N_24256,N_23875);
nand U29623 (N_29623,N_22557,N_21163);
nand U29624 (N_29624,N_20778,N_23458);
or U29625 (N_29625,N_23732,N_24963);
and U29626 (N_29626,N_20568,N_22169);
nand U29627 (N_29627,N_20272,N_21966);
and U29628 (N_29628,N_22261,N_22410);
nand U29629 (N_29629,N_20381,N_21340);
or U29630 (N_29630,N_22066,N_22249);
or U29631 (N_29631,N_22209,N_20173);
nand U29632 (N_29632,N_22011,N_23370);
or U29633 (N_29633,N_20210,N_23694);
and U29634 (N_29634,N_20719,N_23777);
and U29635 (N_29635,N_20223,N_20644);
nand U29636 (N_29636,N_24654,N_22833);
nor U29637 (N_29637,N_24211,N_20735);
nor U29638 (N_29638,N_23801,N_24003);
or U29639 (N_29639,N_22495,N_21792);
or U29640 (N_29640,N_23608,N_22705);
and U29641 (N_29641,N_21093,N_23843);
and U29642 (N_29642,N_20126,N_21798);
nor U29643 (N_29643,N_23383,N_22315);
or U29644 (N_29644,N_22749,N_22096);
nor U29645 (N_29645,N_21810,N_20705);
or U29646 (N_29646,N_20584,N_21963);
nand U29647 (N_29647,N_22065,N_21440);
nand U29648 (N_29648,N_20862,N_23426);
and U29649 (N_29649,N_23698,N_22352);
nand U29650 (N_29650,N_21080,N_23387);
nor U29651 (N_29651,N_23530,N_20508);
or U29652 (N_29652,N_24930,N_22664);
and U29653 (N_29653,N_24035,N_24656);
nand U29654 (N_29654,N_21108,N_20841);
xnor U29655 (N_29655,N_21171,N_23524);
nand U29656 (N_29656,N_21994,N_20965);
or U29657 (N_29657,N_24330,N_21377);
nor U29658 (N_29658,N_24601,N_23695);
nand U29659 (N_29659,N_21998,N_24231);
and U29660 (N_29660,N_23233,N_21344);
nand U29661 (N_29661,N_22608,N_21948);
nand U29662 (N_29662,N_21741,N_22195);
nor U29663 (N_29663,N_22724,N_22267);
nand U29664 (N_29664,N_21910,N_23393);
and U29665 (N_29665,N_21270,N_20137);
or U29666 (N_29666,N_20598,N_22339);
nand U29667 (N_29667,N_22160,N_21277);
and U29668 (N_29668,N_21852,N_23736);
nand U29669 (N_29669,N_20588,N_23129);
or U29670 (N_29670,N_22623,N_24221);
and U29671 (N_29671,N_20855,N_22838);
and U29672 (N_29672,N_23663,N_21651);
and U29673 (N_29673,N_21303,N_20214);
nor U29674 (N_29674,N_20321,N_23652);
or U29675 (N_29675,N_21655,N_21840);
nand U29676 (N_29676,N_23321,N_20355);
and U29677 (N_29677,N_22578,N_23330);
nand U29678 (N_29678,N_20946,N_22481);
nand U29679 (N_29679,N_24486,N_24632);
or U29680 (N_29680,N_22973,N_22657);
nand U29681 (N_29681,N_24129,N_21213);
nand U29682 (N_29682,N_24829,N_21195);
nor U29683 (N_29683,N_23090,N_21325);
or U29684 (N_29684,N_22295,N_21406);
or U29685 (N_29685,N_24763,N_20068);
nor U29686 (N_29686,N_20286,N_21420);
nor U29687 (N_29687,N_24839,N_20833);
nor U29688 (N_29688,N_24226,N_20422);
and U29689 (N_29689,N_21019,N_21392);
nor U29690 (N_29690,N_22474,N_23748);
and U29691 (N_29691,N_22862,N_21876);
nor U29692 (N_29692,N_22547,N_24152);
nand U29693 (N_29693,N_24258,N_24809);
or U29694 (N_29694,N_21829,N_23692);
and U29695 (N_29695,N_22681,N_21033);
or U29696 (N_29696,N_21706,N_23574);
nand U29697 (N_29697,N_20937,N_23455);
and U29698 (N_29698,N_24675,N_20795);
nand U29699 (N_29699,N_24565,N_20357);
nand U29700 (N_29700,N_24063,N_20160);
xor U29701 (N_29701,N_21175,N_20913);
or U29702 (N_29702,N_24550,N_21349);
and U29703 (N_29703,N_21792,N_23086);
and U29704 (N_29704,N_21569,N_22063);
or U29705 (N_29705,N_20952,N_23987);
nand U29706 (N_29706,N_24180,N_24283);
nand U29707 (N_29707,N_21720,N_21337);
nor U29708 (N_29708,N_20159,N_23545);
nand U29709 (N_29709,N_22600,N_22730);
or U29710 (N_29710,N_22890,N_22963);
nor U29711 (N_29711,N_22060,N_21639);
and U29712 (N_29712,N_24308,N_24229);
or U29713 (N_29713,N_24358,N_24864);
nand U29714 (N_29714,N_23847,N_24185);
or U29715 (N_29715,N_23737,N_24526);
nor U29716 (N_29716,N_24117,N_24922);
nand U29717 (N_29717,N_20872,N_23049);
and U29718 (N_29718,N_20751,N_21765);
nand U29719 (N_29719,N_24667,N_22285);
nand U29720 (N_29720,N_22672,N_20910);
and U29721 (N_29721,N_21334,N_21275);
nand U29722 (N_29722,N_23029,N_20262);
nor U29723 (N_29723,N_23264,N_20856);
nor U29724 (N_29724,N_20623,N_22006);
xor U29725 (N_29725,N_22859,N_21854);
or U29726 (N_29726,N_24857,N_21737);
nor U29727 (N_29727,N_23422,N_23901);
nor U29728 (N_29728,N_22812,N_22706);
nor U29729 (N_29729,N_24823,N_22757);
nor U29730 (N_29730,N_20962,N_21704);
and U29731 (N_29731,N_22092,N_21785);
xor U29732 (N_29732,N_24871,N_22843);
or U29733 (N_29733,N_22361,N_21154);
and U29734 (N_29734,N_21361,N_23083);
nand U29735 (N_29735,N_22893,N_20525);
nor U29736 (N_29736,N_21786,N_22819);
or U29737 (N_29737,N_21099,N_20086);
or U29738 (N_29738,N_23130,N_24417);
and U29739 (N_29739,N_21278,N_22073);
and U29740 (N_29740,N_22656,N_24621);
and U29741 (N_29741,N_21642,N_22629);
nor U29742 (N_29742,N_24901,N_23122);
or U29743 (N_29743,N_23169,N_23366);
nand U29744 (N_29744,N_23460,N_23122);
or U29745 (N_29745,N_23449,N_20582);
or U29746 (N_29746,N_21722,N_20983);
nand U29747 (N_29747,N_23357,N_21165);
xnor U29748 (N_29748,N_21411,N_22353);
or U29749 (N_29749,N_21969,N_21516);
nand U29750 (N_29750,N_24569,N_21130);
and U29751 (N_29751,N_22385,N_20953);
nor U29752 (N_29752,N_22093,N_24768);
and U29753 (N_29753,N_24740,N_20894);
nand U29754 (N_29754,N_20146,N_21069);
and U29755 (N_29755,N_22641,N_22012);
nor U29756 (N_29756,N_22311,N_20650);
or U29757 (N_29757,N_22958,N_23378);
nand U29758 (N_29758,N_20669,N_22995);
or U29759 (N_29759,N_21970,N_23371);
or U29760 (N_29760,N_23195,N_20087);
nor U29761 (N_29761,N_22613,N_24215);
or U29762 (N_29762,N_22957,N_20253);
or U29763 (N_29763,N_21451,N_21543);
and U29764 (N_29764,N_23808,N_22783);
or U29765 (N_29765,N_21851,N_20286);
and U29766 (N_29766,N_23270,N_22511);
nand U29767 (N_29767,N_22931,N_22028);
nand U29768 (N_29768,N_23519,N_23345);
or U29769 (N_29769,N_20332,N_22818);
or U29770 (N_29770,N_24212,N_20468);
and U29771 (N_29771,N_23564,N_21229);
xor U29772 (N_29772,N_20056,N_23203);
nor U29773 (N_29773,N_21352,N_24766);
nand U29774 (N_29774,N_24622,N_24418);
nand U29775 (N_29775,N_22905,N_21317);
nor U29776 (N_29776,N_22417,N_20508);
nor U29777 (N_29777,N_23995,N_20270);
or U29778 (N_29778,N_24913,N_22406);
and U29779 (N_29779,N_24563,N_20478);
nor U29780 (N_29780,N_23136,N_22764);
nor U29781 (N_29781,N_24426,N_22867);
or U29782 (N_29782,N_21447,N_23252);
and U29783 (N_29783,N_21062,N_22236);
or U29784 (N_29784,N_24565,N_20829);
nand U29785 (N_29785,N_23601,N_24238);
nor U29786 (N_29786,N_23240,N_24484);
and U29787 (N_29787,N_21993,N_22709);
or U29788 (N_29788,N_23555,N_20630);
nor U29789 (N_29789,N_22322,N_21611);
nand U29790 (N_29790,N_20649,N_20041);
nor U29791 (N_29791,N_23979,N_20832);
or U29792 (N_29792,N_23963,N_23166);
or U29793 (N_29793,N_23054,N_23708);
and U29794 (N_29794,N_22279,N_22019);
or U29795 (N_29795,N_23567,N_24484);
or U29796 (N_29796,N_22765,N_23404);
or U29797 (N_29797,N_24670,N_22656);
nand U29798 (N_29798,N_21971,N_21705);
nor U29799 (N_29799,N_20291,N_21239);
and U29800 (N_29800,N_22850,N_24103);
nor U29801 (N_29801,N_22709,N_24852);
or U29802 (N_29802,N_23112,N_20334);
nor U29803 (N_29803,N_24694,N_21536);
nor U29804 (N_29804,N_24012,N_20400);
nand U29805 (N_29805,N_21578,N_24630);
nand U29806 (N_29806,N_24258,N_22163);
and U29807 (N_29807,N_24257,N_24081);
nor U29808 (N_29808,N_22521,N_20569);
or U29809 (N_29809,N_22067,N_21375);
or U29810 (N_29810,N_20677,N_24060);
nand U29811 (N_29811,N_21051,N_23134);
or U29812 (N_29812,N_21366,N_22341);
nand U29813 (N_29813,N_23845,N_21221);
and U29814 (N_29814,N_22122,N_20177);
or U29815 (N_29815,N_23814,N_24082);
or U29816 (N_29816,N_23616,N_22783);
or U29817 (N_29817,N_21257,N_24984);
or U29818 (N_29818,N_22667,N_20199);
or U29819 (N_29819,N_21045,N_24104);
nor U29820 (N_29820,N_22255,N_24588);
or U29821 (N_29821,N_21872,N_21471);
nor U29822 (N_29822,N_20931,N_23402);
nor U29823 (N_29823,N_22587,N_20968);
nor U29824 (N_29824,N_22624,N_23128);
nand U29825 (N_29825,N_24811,N_23102);
or U29826 (N_29826,N_23693,N_22837);
nand U29827 (N_29827,N_20219,N_21851);
or U29828 (N_29828,N_24477,N_23200);
and U29829 (N_29829,N_23913,N_21635);
or U29830 (N_29830,N_21327,N_24810);
or U29831 (N_29831,N_23681,N_23704);
and U29832 (N_29832,N_21269,N_22597);
nor U29833 (N_29833,N_23810,N_21358);
and U29834 (N_29834,N_22224,N_23598);
nand U29835 (N_29835,N_23173,N_24826);
and U29836 (N_29836,N_20047,N_23872);
nor U29837 (N_29837,N_21944,N_22256);
nand U29838 (N_29838,N_24841,N_24412);
or U29839 (N_29839,N_20088,N_21981);
nor U29840 (N_29840,N_21527,N_20578);
or U29841 (N_29841,N_20672,N_24609);
nor U29842 (N_29842,N_22317,N_24309);
nor U29843 (N_29843,N_23581,N_24210);
or U29844 (N_29844,N_23476,N_20915);
nand U29845 (N_29845,N_21044,N_20669);
or U29846 (N_29846,N_20996,N_23031);
or U29847 (N_29847,N_23283,N_20517);
or U29848 (N_29848,N_22094,N_22183);
and U29849 (N_29849,N_24250,N_23921);
nor U29850 (N_29850,N_24399,N_24489);
or U29851 (N_29851,N_21912,N_22495);
nor U29852 (N_29852,N_24695,N_23766);
and U29853 (N_29853,N_23506,N_24210);
or U29854 (N_29854,N_22987,N_24653);
or U29855 (N_29855,N_21606,N_21864);
nor U29856 (N_29856,N_24608,N_20925);
and U29857 (N_29857,N_21876,N_22704);
nor U29858 (N_29858,N_20984,N_21633);
nand U29859 (N_29859,N_22004,N_23574);
or U29860 (N_29860,N_23389,N_20055);
nand U29861 (N_29861,N_20248,N_22544);
nand U29862 (N_29862,N_22028,N_22446);
or U29863 (N_29863,N_21535,N_24868);
nand U29864 (N_29864,N_21906,N_22879);
or U29865 (N_29865,N_20829,N_22853);
nor U29866 (N_29866,N_22018,N_21896);
nor U29867 (N_29867,N_22359,N_21345);
and U29868 (N_29868,N_24766,N_22329);
or U29869 (N_29869,N_24393,N_24693);
nor U29870 (N_29870,N_24215,N_20825);
or U29871 (N_29871,N_23190,N_21783);
nand U29872 (N_29872,N_24414,N_20200);
or U29873 (N_29873,N_20880,N_21070);
nand U29874 (N_29874,N_23801,N_21510);
nor U29875 (N_29875,N_24532,N_22137);
or U29876 (N_29876,N_20017,N_23533);
nand U29877 (N_29877,N_23800,N_20348);
and U29878 (N_29878,N_20877,N_23959);
nor U29879 (N_29879,N_21364,N_23845);
and U29880 (N_29880,N_23334,N_23629);
or U29881 (N_29881,N_24879,N_24679);
nand U29882 (N_29882,N_23908,N_21995);
nand U29883 (N_29883,N_22552,N_22564);
nor U29884 (N_29884,N_21365,N_23584);
nand U29885 (N_29885,N_20256,N_21516);
xor U29886 (N_29886,N_24582,N_20254);
nor U29887 (N_29887,N_22332,N_21563);
nor U29888 (N_29888,N_22628,N_20043);
or U29889 (N_29889,N_23557,N_23548);
nand U29890 (N_29890,N_23206,N_22450);
nor U29891 (N_29891,N_22298,N_21446);
or U29892 (N_29892,N_20435,N_21919);
nand U29893 (N_29893,N_21818,N_22758);
or U29894 (N_29894,N_23547,N_23416);
nand U29895 (N_29895,N_24334,N_22231);
and U29896 (N_29896,N_24044,N_23000);
nor U29897 (N_29897,N_23657,N_24137);
and U29898 (N_29898,N_20386,N_23744);
and U29899 (N_29899,N_24521,N_24010);
nand U29900 (N_29900,N_23338,N_24681);
and U29901 (N_29901,N_22037,N_21769);
or U29902 (N_29902,N_21600,N_23952);
nor U29903 (N_29903,N_21399,N_21009);
xnor U29904 (N_29904,N_22202,N_24468);
or U29905 (N_29905,N_21695,N_23494);
nand U29906 (N_29906,N_21529,N_22379);
and U29907 (N_29907,N_20148,N_23822);
or U29908 (N_29908,N_22460,N_23212);
or U29909 (N_29909,N_23395,N_24576);
nor U29910 (N_29910,N_20562,N_20070);
nand U29911 (N_29911,N_21070,N_22489);
and U29912 (N_29912,N_22976,N_23747);
or U29913 (N_29913,N_24134,N_21525);
nor U29914 (N_29914,N_22235,N_22144);
or U29915 (N_29915,N_24808,N_20486);
nor U29916 (N_29916,N_21601,N_20926);
or U29917 (N_29917,N_20011,N_24316);
nand U29918 (N_29918,N_23780,N_22518);
nor U29919 (N_29919,N_20014,N_20276);
and U29920 (N_29920,N_23295,N_22256);
nor U29921 (N_29921,N_21727,N_24392);
and U29922 (N_29922,N_24836,N_23121);
nor U29923 (N_29923,N_21604,N_22529);
nand U29924 (N_29924,N_24406,N_24204);
and U29925 (N_29925,N_22797,N_21604);
nor U29926 (N_29926,N_21885,N_21577);
nand U29927 (N_29927,N_20000,N_20732);
and U29928 (N_29928,N_24605,N_23745);
nand U29929 (N_29929,N_20148,N_24032);
nor U29930 (N_29930,N_23923,N_20914);
nor U29931 (N_29931,N_21234,N_20181);
nor U29932 (N_29932,N_23207,N_23915);
and U29933 (N_29933,N_21731,N_21073);
nor U29934 (N_29934,N_24238,N_24054);
nand U29935 (N_29935,N_24438,N_22526);
nor U29936 (N_29936,N_22216,N_22007);
and U29937 (N_29937,N_20462,N_23074);
xnor U29938 (N_29938,N_24245,N_23916);
and U29939 (N_29939,N_22550,N_21736);
nand U29940 (N_29940,N_24840,N_20190);
and U29941 (N_29941,N_20242,N_22666);
nor U29942 (N_29942,N_23199,N_24221);
and U29943 (N_29943,N_23881,N_24168);
nor U29944 (N_29944,N_20633,N_22293);
and U29945 (N_29945,N_22507,N_23205);
or U29946 (N_29946,N_24052,N_20422);
nor U29947 (N_29947,N_21836,N_20886);
nand U29948 (N_29948,N_23049,N_23192);
or U29949 (N_29949,N_20628,N_24483);
nor U29950 (N_29950,N_22188,N_21569);
and U29951 (N_29951,N_24735,N_22099);
or U29952 (N_29952,N_23913,N_23800);
nand U29953 (N_29953,N_23594,N_24805);
or U29954 (N_29954,N_21955,N_23221);
or U29955 (N_29955,N_24379,N_24507);
nand U29956 (N_29956,N_20654,N_24260);
or U29957 (N_29957,N_23572,N_24997);
and U29958 (N_29958,N_23966,N_24783);
nand U29959 (N_29959,N_22690,N_20550);
and U29960 (N_29960,N_20102,N_23581);
and U29961 (N_29961,N_21304,N_21209);
nand U29962 (N_29962,N_23908,N_21384);
and U29963 (N_29963,N_21541,N_21261);
nor U29964 (N_29964,N_23585,N_24586);
nor U29965 (N_29965,N_20207,N_24837);
or U29966 (N_29966,N_23220,N_24733);
nor U29967 (N_29967,N_22704,N_22291);
nor U29968 (N_29968,N_20704,N_22072);
or U29969 (N_29969,N_24369,N_23646);
or U29970 (N_29970,N_22011,N_24264);
and U29971 (N_29971,N_20512,N_22841);
and U29972 (N_29972,N_23799,N_22598);
and U29973 (N_29973,N_24735,N_23214);
or U29974 (N_29974,N_24227,N_24453);
or U29975 (N_29975,N_23466,N_24860);
nand U29976 (N_29976,N_20536,N_22859);
and U29977 (N_29977,N_23149,N_23456);
or U29978 (N_29978,N_23151,N_23524);
and U29979 (N_29979,N_24511,N_24221);
nor U29980 (N_29980,N_20073,N_22776);
nor U29981 (N_29981,N_24272,N_20400);
and U29982 (N_29982,N_20873,N_24950);
nand U29983 (N_29983,N_22454,N_23327);
nor U29984 (N_29984,N_23969,N_20344);
nand U29985 (N_29985,N_24886,N_20297);
nor U29986 (N_29986,N_20926,N_20550);
or U29987 (N_29987,N_22588,N_23585);
nand U29988 (N_29988,N_24399,N_22990);
or U29989 (N_29989,N_21653,N_22978);
or U29990 (N_29990,N_22955,N_21626);
and U29991 (N_29991,N_21434,N_24905);
and U29992 (N_29992,N_22591,N_20151);
or U29993 (N_29993,N_21683,N_24300);
nor U29994 (N_29994,N_22828,N_22736);
and U29995 (N_29995,N_23040,N_23465);
and U29996 (N_29996,N_24000,N_20702);
nand U29997 (N_29997,N_24529,N_20099);
and U29998 (N_29998,N_21276,N_23285);
nor U29999 (N_29999,N_22145,N_22271);
or UO_0 (O_0,N_29917,N_27711);
nor UO_1 (O_1,N_28590,N_27087);
and UO_2 (O_2,N_25038,N_29393);
or UO_3 (O_3,N_25750,N_25494);
nor UO_4 (O_4,N_28958,N_26226);
nand UO_5 (O_5,N_25702,N_25086);
nor UO_6 (O_6,N_26788,N_26518);
nor UO_7 (O_7,N_29907,N_28623);
and UO_8 (O_8,N_26279,N_25272);
xnor UO_9 (O_9,N_29378,N_29718);
or UO_10 (O_10,N_29660,N_28896);
nor UO_11 (O_11,N_27192,N_28625);
and UO_12 (O_12,N_28082,N_28575);
nor UO_13 (O_13,N_26417,N_28968);
and UO_14 (O_14,N_26013,N_26478);
and UO_15 (O_15,N_28318,N_29515);
or UO_16 (O_16,N_27196,N_27907);
or UO_17 (O_17,N_25168,N_28086);
and UO_18 (O_18,N_25119,N_28023);
or UO_19 (O_19,N_29412,N_29291);
and UO_20 (O_20,N_25626,N_25635);
nor UO_21 (O_21,N_27623,N_28038);
and UO_22 (O_22,N_26908,N_27575);
nor UO_23 (O_23,N_25928,N_26935);
nor UO_24 (O_24,N_28397,N_27181);
nor UO_25 (O_25,N_29890,N_25584);
nand UO_26 (O_26,N_27870,N_26324);
nand UO_27 (O_27,N_25137,N_27313);
or UO_28 (O_28,N_29128,N_27372);
nor UO_29 (O_29,N_26234,N_25638);
nand UO_30 (O_30,N_28889,N_28765);
or UO_31 (O_31,N_29292,N_25955);
and UO_32 (O_32,N_28155,N_26099);
or UO_33 (O_33,N_29299,N_26424);
nor UO_34 (O_34,N_27285,N_29851);
nand UO_35 (O_35,N_28634,N_26427);
or UO_36 (O_36,N_27074,N_27107);
and UO_37 (O_37,N_26799,N_27947);
nor UO_38 (O_38,N_29894,N_28714);
or UO_39 (O_39,N_29102,N_26214);
nor UO_40 (O_40,N_27662,N_28261);
and UO_41 (O_41,N_27164,N_29290);
or UO_42 (O_42,N_28532,N_26028);
nor UO_43 (O_43,N_29664,N_29263);
and UO_44 (O_44,N_28972,N_27396);
nor UO_45 (O_45,N_26253,N_29830);
nand UO_46 (O_46,N_27780,N_27893);
nand UO_47 (O_47,N_25158,N_28276);
or UO_48 (O_48,N_27763,N_29641);
and UO_49 (O_49,N_27162,N_25256);
and UO_50 (O_50,N_28867,N_25355);
nor UO_51 (O_51,N_27266,N_26561);
and UO_52 (O_52,N_26108,N_28761);
nor UO_53 (O_53,N_25399,N_25043);
nand UO_54 (O_54,N_26785,N_28418);
nor UO_55 (O_55,N_28738,N_27900);
nand UO_56 (O_56,N_27543,N_29705);
and UO_57 (O_57,N_28736,N_27448);
or UO_58 (O_58,N_26490,N_29261);
or UO_59 (O_59,N_27921,N_28823);
nor UO_60 (O_60,N_27265,N_29346);
or UO_61 (O_61,N_29151,N_25593);
or UO_62 (O_62,N_25010,N_28419);
nor UO_63 (O_63,N_28204,N_29413);
and UO_64 (O_64,N_28747,N_25837);
nand UO_65 (O_65,N_25933,N_28335);
nand UO_66 (O_66,N_28391,N_27059);
or UO_67 (O_67,N_29030,N_29268);
nor UO_68 (O_68,N_29795,N_26900);
nand UO_69 (O_69,N_27830,N_28321);
nor UO_70 (O_70,N_29174,N_27225);
nor UO_71 (O_71,N_25711,N_29309);
or UO_72 (O_72,N_28196,N_29879);
nand UO_73 (O_73,N_28721,N_29588);
nor UO_74 (O_74,N_29672,N_29853);
or UO_75 (O_75,N_27823,N_29583);
and UO_76 (O_76,N_28599,N_26633);
nand UO_77 (O_77,N_27776,N_28710);
or UO_78 (O_78,N_29329,N_25329);
nand UO_79 (O_79,N_28413,N_28331);
nor UO_80 (O_80,N_26601,N_27946);
nand UO_81 (O_81,N_28030,N_28212);
nand UO_82 (O_82,N_29791,N_29304);
or UO_83 (O_83,N_26005,N_26513);
or UO_84 (O_84,N_29365,N_27938);
nor UO_85 (O_85,N_29167,N_26575);
nand UO_86 (O_86,N_28778,N_25846);
or UO_87 (O_87,N_27844,N_27046);
nand UO_88 (O_88,N_25896,N_27995);
and UO_89 (O_89,N_28956,N_27510);
xnor UO_90 (O_90,N_26700,N_25143);
nor UO_91 (O_91,N_27483,N_25686);
nand UO_92 (O_92,N_25989,N_26847);
nor UO_93 (O_93,N_25182,N_28632);
nor UO_94 (O_94,N_27463,N_26964);
nor UO_95 (O_95,N_28617,N_27210);
nor UO_96 (O_96,N_25948,N_26155);
and UO_97 (O_97,N_29944,N_29199);
nand UO_98 (O_98,N_26292,N_29311);
and UO_99 (O_99,N_25585,N_27125);
and UO_100 (O_100,N_29046,N_25284);
and UO_101 (O_101,N_28344,N_26041);
xor UO_102 (O_102,N_26418,N_27215);
nor UO_103 (O_103,N_29020,N_28270);
nor UO_104 (O_104,N_26072,N_26469);
or UO_105 (O_105,N_28376,N_25135);
and UO_106 (O_106,N_25788,N_25558);
or UO_107 (O_107,N_27614,N_25311);
or UO_108 (O_108,N_27977,N_26716);
and UO_109 (O_109,N_27580,N_25792);
nand UO_110 (O_110,N_29258,N_28474);
nor UO_111 (O_111,N_26649,N_28804);
nand UO_112 (O_112,N_27885,N_29658);
nand UO_113 (O_113,N_29691,N_29081);
and UO_114 (O_114,N_27010,N_29508);
or UO_115 (O_115,N_27650,N_26530);
nand UO_116 (O_116,N_28537,N_26846);
nor UO_117 (O_117,N_28272,N_28871);
nand UO_118 (O_118,N_28337,N_27479);
and UO_119 (O_119,N_27677,N_26824);
nand UO_120 (O_120,N_28002,N_25688);
or UO_121 (O_121,N_25631,N_28696);
and UO_122 (O_122,N_29009,N_27993);
nand UO_123 (O_123,N_28910,N_25213);
nor UO_124 (O_124,N_25348,N_25965);
nor UO_125 (O_125,N_25561,N_28458);
nand UO_126 (O_126,N_29903,N_29127);
nor UO_127 (O_127,N_25861,N_28529);
nor UO_128 (O_128,N_27268,N_25198);
nor UO_129 (O_129,N_25496,N_27682);
nor UO_130 (O_130,N_26671,N_28745);
nor UO_131 (O_131,N_27332,N_29112);
or UO_132 (O_132,N_27040,N_28841);
nor UO_133 (O_133,N_27950,N_27916);
xor UO_134 (O_134,N_26163,N_28184);
nand UO_135 (O_135,N_28589,N_29667);
nand UO_136 (O_136,N_28917,N_28789);
nor UO_137 (O_137,N_25733,N_25465);
nand UO_138 (O_138,N_28366,N_29482);
or UO_139 (O_139,N_28856,N_26133);
or UO_140 (O_140,N_29527,N_27604);
and UO_141 (O_141,N_25338,N_27974);
or UO_142 (O_142,N_25673,N_26722);
and UO_143 (O_143,N_25128,N_25124);
and UO_144 (O_144,N_28894,N_27175);
and UO_145 (O_145,N_28223,N_26567);
nand UO_146 (O_146,N_29395,N_28785);
or UO_147 (O_147,N_26614,N_29981);
or UO_148 (O_148,N_27718,N_29007);
nand UO_149 (O_149,N_26387,N_27457);
nor UO_150 (O_150,N_26886,N_26271);
or UO_151 (O_151,N_28729,N_28467);
nand UO_152 (O_152,N_25061,N_26910);
nor UO_153 (O_153,N_28959,N_26458);
nand UO_154 (O_154,N_29977,N_27169);
or UO_155 (O_155,N_26315,N_28020);
or UO_156 (O_156,N_27636,N_27300);
and UO_157 (O_157,N_27739,N_28058);
nor UO_158 (O_158,N_26980,N_27027);
and UO_159 (O_159,N_29699,N_28792);
or UO_160 (O_160,N_27085,N_28843);
and UO_161 (O_161,N_28567,N_26025);
nor UO_162 (O_162,N_27451,N_27983);
or UO_163 (O_163,N_26540,N_29845);
nor UO_164 (O_164,N_28647,N_29695);
nor UO_165 (O_165,N_28147,N_25344);
nor UO_166 (O_166,N_27366,N_26479);
or UO_167 (O_167,N_26002,N_29088);
nand UO_168 (O_168,N_26423,N_29473);
and UO_169 (O_169,N_27425,N_28516);
or UO_170 (O_170,N_27480,N_28370);
or UO_171 (O_171,N_28062,N_27088);
nor UO_172 (O_172,N_27081,N_27506);
nor UO_173 (O_173,N_29563,N_29130);
nand UO_174 (O_174,N_26851,N_29760);
nor UO_175 (O_175,N_25277,N_28495);
nand UO_176 (O_176,N_25574,N_29840);
and UO_177 (O_177,N_26573,N_25629);
nand UO_178 (O_178,N_28712,N_25562);
or UO_179 (O_179,N_25567,N_29385);
nand UO_180 (O_180,N_28648,N_25588);
and UO_181 (O_181,N_29421,N_25375);
and UO_182 (O_182,N_25620,N_25110);
and UO_183 (O_183,N_26791,N_26285);
and UO_184 (O_184,N_29864,N_25359);
or UO_185 (O_185,N_29051,N_25007);
nor UO_186 (O_186,N_29049,N_25270);
or UO_187 (O_187,N_26061,N_25217);
and UO_188 (O_188,N_29679,N_26263);
and UO_189 (O_189,N_26245,N_27436);
or UO_190 (O_190,N_26773,N_27752);
nor UO_191 (O_191,N_29888,N_28796);
or UO_192 (O_192,N_28387,N_28128);
or UO_193 (O_193,N_27291,N_28024);
nand UO_194 (O_194,N_27554,N_25508);
nor UO_195 (O_195,N_28597,N_29033);
nor UO_196 (O_196,N_27020,N_25615);
or UO_197 (O_197,N_29838,N_26820);
xor UO_198 (O_198,N_28072,N_26294);
or UO_199 (O_199,N_28156,N_28362);
or UO_200 (O_200,N_29477,N_26859);
nor UO_201 (O_201,N_26645,N_26465);
and UO_202 (O_202,N_27850,N_27271);
or UO_203 (O_203,N_28669,N_29294);
nand UO_204 (O_204,N_26166,N_28799);
nand UO_205 (O_205,N_28787,N_26686);
nor UO_206 (O_206,N_29459,N_28868);
xor UO_207 (O_207,N_28578,N_25319);
xnor UO_208 (O_208,N_27854,N_25790);
or UO_209 (O_209,N_26201,N_26351);
and UO_210 (O_210,N_26734,N_25192);
or UO_211 (O_211,N_26943,N_25550);
nand UO_212 (O_212,N_25824,N_29735);
nor UO_213 (O_213,N_26728,N_27043);
and UO_214 (O_214,N_25781,N_25899);
and UO_215 (O_215,N_27367,N_27527);
nor UO_216 (O_216,N_29204,N_28472);
nand UO_217 (O_217,N_27464,N_28970);
and UO_218 (O_218,N_27061,N_26938);
and UO_219 (O_219,N_26709,N_26221);
nand UO_220 (O_220,N_27174,N_25041);
nor UO_221 (O_221,N_27454,N_27129);
and UO_222 (O_222,N_26774,N_26874);
and UO_223 (O_223,N_26555,N_26589);
or UO_224 (O_224,N_29195,N_25647);
and UO_225 (O_225,N_26492,N_29752);
nand UO_226 (O_226,N_29178,N_29974);
and UO_227 (O_227,N_28498,N_29017);
nand UO_228 (O_228,N_29420,N_28766);
nor UO_229 (O_229,N_26995,N_29465);
nand UO_230 (O_230,N_26924,N_27672);
and UO_231 (O_231,N_26339,N_29690);
nand UO_232 (O_232,N_26616,N_28011);
or UO_233 (O_233,N_25268,N_27071);
and UO_234 (O_234,N_28887,N_25705);
or UO_235 (O_235,N_27775,N_29483);
and UO_236 (O_236,N_28506,N_27132);
nor UO_237 (O_237,N_26477,N_29629);
nand UO_238 (O_238,N_27991,N_29436);
nor UO_239 (O_239,N_29933,N_27701);
or UO_240 (O_240,N_28838,N_29739);
nand UO_241 (O_241,N_28189,N_27449);
nand UO_242 (O_242,N_25822,N_26993);
or UO_243 (O_243,N_27504,N_25808);
or UO_244 (O_244,N_25358,N_25935);
nand UO_245 (O_245,N_27298,N_27104);
and UO_246 (O_246,N_28649,N_27564);
and UO_247 (O_247,N_26176,N_26172);
nand UO_248 (O_248,N_27136,N_25627);
nor UO_249 (O_249,N_27676,N_26033);
and UO_250 (O_250,N_25022,N_29676);
and UO_251 (O_251,N_26243,N_28754);
nor UO_252 (O_252,N_25271,N_27640);
nand UO_253 (O_253,N_26648,N_29960);
nand UO_254 (O_254,N_28012,N_28350);
nand UO_255 (O_255,N_29861,N_26766);
nor UO_256 (O_256,N_29991,N_27121);
nor UO_257 (O_257,N_27688,N_27748);
or UO_258 (O_258,N_26174,N_27001);
nor UO_259 (O_259,N_26703,N_25551);
and UO_260 (O_260,N_25547,N_27227);
or UO_261 (O_261,N_26609,N_29332);
and UO_262 (O_262,N_26067,N_26157);
and UO_263 (O_263,N_25873,N_28517);
or UO_264 (O_264,N_25067,N_29580);
or UO_265 (O_265,N_28888,N_25829);
and UO_266 (O_266,N_27857,N_29463);
and UO_267 (O_267,N_29634,N_27557);
nor UO_268 (O_268,N_29249,N_27545);
nand UO_269 (O_269,N_29386,N_29206);
and UO_270 (O_270,N_28361,N_29132);
and UO_271 (O_271,N_26866,N_26485);
and UO_272 (O_272,N_28586,N_27526);
nand UO_273 (O_273,N_27028,N_29498);
nor UO_274 (O_274,N_27865,N_29996);
and UO_275 (O_275,N_29955,N_28760);
nor UO_276 (O_276,N_25764,N_26738);
and UO_277 (O_277,N_27073,N_27660);
or UO_278 (O_278,N_26447,N_26336);
and UO_279 (O_279,N_28298,N_27864);
nand UO_280 (O_280,N_29554,N_27962);
and UO_281 (O_281,N_29601,N_29157);
nand UO_282 (O_282,N_27612,N_27301);
or UO_283 (O_283,N_28149,N_26739);
or UO_284 (O_284,N_26302,N_26317);
and UO_285 (O_285,N_27394,N_26737);
nand UO_286 (O_286,N_25078,N_26319);
and UO_287 (O_287,N_26096,N_27333);
or UO_288 (O_288,N_25062,N_29942);
nand UO_289 (O_289,N_26660,N_27245);
or UO_290 (O_290,N_29243,N_25720);
nor UO_291 (O_291,N_28866,N_29417);
or UO_292 (O_292,N_25579,N_26316);
xor UO_293 (O_293,N_25658,N_26974);
or UO_294 (O_294,N_28192,N_29700);
and UO_295 (O_295,N_29817,N_29442);
and UO_296 (O_296,N_27972,N_29107);
nor UO_297 (O_297,N_29466,N_27751);
and UO_298 (O_298,N_25232,N_27744);
xor UO_299 (O_299,N_26014,N_28892);
nor UO_300 (O_300,N_26957,N_28167);
nor UO_301 (O_301,N_29771,N_28718);
nand UO_302 (O_302,N_28975,N_27171);
and UO_303 (O_303,N_28333,N_29059);
nand UO_304 (O_304,N_27696,N_29574);
nand UO_305 (O_305,N_25677,N_27511);
or UO_306 (O_306,N_27737,N_25501);
nor UO_307 (O_307,N_28724,N_25102);
nand UO_308 (O_308,N_25976,N_28522);
and UO_309 (O_309,N_28832,N_29550);
nand UO_310 (O_310,N_29828,N_29627);
nand UO_311 (O_311,N_29837,N_28946);
or UO_312 (O_312,N_26335,N_28314);
or UO_313 (O_313,N_29284,N_26576);
nand UO_314 (O_314,N_29624,N_27212);
or UO_315 (O_315,N_29392,N_26835);
or UO_316 (O_316,N_25390,N_25998);
nand UO_317 (O_317,N_29802,N_27323);
or UO_318 (O_318,N_29834,N_29098);
nand UO_319 (O_319,N_27615,N_25587);
or UO_320 (O_320,N_28997,N_26466);
or UO_321 (O_321,N_27383,N_28682);
nand UO_322 (O_322,N_28905,N_25307);
nand UO_323 (O_323,N_29135,N_29164);
or UO_324 (O_324,N_28595,N_27118);
nor UO_325 (O_325,N_28142,N_29532);
and UO_326 (O_326,N_26329,N_26801);
or UO_327 (O_327,N_26556,N_26147);
nor UO_328 (O_328,N_25662,N_25690);
nand UO_329 (O_329,N_26797,N_29433);
nand UO_330 (O_330,N_28043,N_26699);
and UO_331 (O_331,N_28004,N_27869);
nand UO_332 (O_332,N_28406,N_27729);
nor UO_333 (O_333,N_25954,N_27205);
and UO_334 (O_334,N_28334,N_29697);
nand UO_335 (O_335,N_25258,N_25616);
and UO_336 (O_336,N_27016,N_25893);
or UO_337 (O_337,N_28213,N_26448);
or UO_338 (O_338,N_25057,N_25224);
nand UO_339 (O_339,N_26714,N_25586);
or UO_340 (O_340,N_28576,N_25595);
and UO_341 (O_341,N_29564,N_27595);
nand UO_342 (O_342,N_25167,N_26973);
and UO_343 (O_343,N_27208,N_26507);
or UO_344 (O_344,N_27646,N_25836);
nand UO_345 (O_345,N_29447,N_26044);
or UO_346 (O_346,N_25623,N_27815);
nor UO_347 (O_347,N_28502,N_28010);
nand UO_348 (O_348,N_28372,N_27159);
nor UO_349 (O_349,N_26624,N_28955);
nand UO_350 (O_350,N_25147,N_27387);
nor UO_351 (O_351,N_25719,N_26111);
nor UO_352 (O_352,N_28249,N_26313);
nor UO_353 (O_353,N_25517,N_28715);
nand UO_354 (O_354,N_28216,N_25709);
or UO_355 (O_355,N_25816,N_26262);
nand UO_356 (O_356,N_29087,N_25883);
nand UO_357 (O_357,N_28728,N_27134);
nor UO_358 (O_358,N_27097,N_25862);
nor UO_359 (O_359,N_26275,N_25019);
and UO_360 (O_360,N_27937,N_29998);
nand UO_361 (O_361,N_26443,N_28433);
and UO_362 (O_362,N_29862,N_25591);
nand UO_363 (O_363,N_26167,N_25944);
nor UO_364 (O_364,N_28425,N_26211);
or UO_365 (O_365,N_29053,N_28533);
and UO_366 (O_366,N_25911,N_27546);
nand UO_367 (O_367,N_27541,N_25756);
or UO_368 (O_368,N_26073,N_29772);
nor UO_369 (O_369,N_27742,N_27655);
nor UO_370 (O_370,N_26008,N_27335);
and UO_371 (O_371,N_28230,N_28929);
nand UO_372 (O_372,N_26265,N_27474);
nor UO_373 (O_373,N_25710,N_27851);
and UO_374 (O_374,N_28412,N_28371);
nor UO_375 (O_375,N_27379,N_26121);
nand UO_376 (O_376,N_28443,N_25646);
nor UO_377 (O_377,N_27812,N_26459);
or UO_378 (O_378,N_28114,N_28503);
or UO_379 (O_379,N_27643,N_27503);
nand UO_380 (O_380,N_28515,N_28731);
nand UO_381 (O_381,N_25885,N_27190);
or UO_382 (O_382,N_27127,N_29505);
or UO_383 (O_383,N_27072,N_29632);
or UO_384 (O_384,N_25323,N_25146);
nand UO_385 (O_385,N_27499,N_29720);
or UO_386 (O_386,N_27060,N_28379);
or UO_387 (O_387,N_27876,N_28007);
and UO_388 (O_388,N_28709,N_26701);
nand UO_389 (O_389,N_27350,N_29794);
or UO_390 (O_390,N_25197,N_27579);
nor UO_391 (O_391,N_26752,N_25308);
nor UO_392 (O_392,N_28422,N_26128);
and UO_393 (O_393,N_26710,N_29060);
and UO_394 (O_394,N_26487,N_25990);
and UO_395 (O_395,N_25956,N_27610);
or UO_396 (O_396,N_27684,N_26227);
and UO_397 (O_397,N_26607,N_26720);
and UO_398 (O_398,N_27337,N_27468);
nand UO_399 (O_399,N_27030,N_25231);
nor UO_400 (O_400,N_26353,N_27585);
nand UO_401 (O_401,N_25863,N_26305);
and UO_402 (O_402,N_29653,N_26963);
and UO_403 (O_403,N_25510,N_27182);
and UO_404 (O_404,N_28779,N_26257);
and UO_405 (O_405,N_26978,N_28873);
nor UO_406 (O_406,N_26168,N_25054);
nor UO_407 (O_407,N_25384,N_25092);
and UO_408 (O_408,N_28199,N_26162);
and UO_409 (O_409,N_27009,N_29230);
and UO_410 (O_410,N_29723,N_26250);
xnor UO_411 (O_411,N_26220,N_27845);
nand UO_412 (O_412,N_28982,N_27941);
nand UO_413 (O_413,N_26876,N_27374);
nor UO_414 (O_414,N_26732,N_28036);
or UO_415 (O_415,N_25503,N_28901);
and UO_416 (O_416,N_27793,N_27658);
nor UO_417 (O_417,N_27805,N_25749);
nor UO_418 (O_418,N_28540,N_28803);
or UO_419 (O_419,N_27879,N_25907);
nor UO_420 (O_420,N_29429,N_28568);
and UO_421 (O_421,N_26454,N_29809);
nor UO_422 (O_422,N_27819,N_28313);
nand UO_423 (O_423,N_28879,N_28463);
nor UO_424 (O_424,N_29786,N_25388);
or UO_425 (O_425,N_28159,N_26094);
nor UO_426 (O_426,N_28525,N_26665);
nor UO_427 (O_427,N_28756,N_29491);
nor UO_428 (O_428,N_29201,N_29185);
nand UO_429 (O_429,N_25763,N_25821);
or UO_430 (O_430,N_29927,N_25652);
or UO_431 (O_431,N_26307,N_26798);
nor UO_432 (O_432,N_25009,N_28478);
and UO_433 (O_433,N_28040,N_26890);
nand UO_434 (O_434,N_28198,N_29486);
and UO_435 (O_435,N_25064,N_27259);
nand UO_436 (O_436,N_29878,N_27814);
nor UO_437 (O_437,N_25035,N_25691);
and UO_438 (O_438,N_27173,N_27553);
and UO_439 (O_439,N_29757,N_29096);
nor UO_440 (O_440,N_27172,N_25859);
nand UO_441 (O_441,N_29576,N_28208);
nor UO_442 (O_442,N_26105,N_27438);
nor UO_443 (O_443,N_25172,N_29022);
and UO_444 (O_444,N_27424,N_27958);
or UO_445 (O_445,N_27154,N_27209);
and UO_446 (O_446,N_26658,N_26228);
nor UO_447 (O_447,N_29360,N_29971);
and UO_448 (O_448,N_28014,N_28903);
nor UO_449 (O_449,N_28624,N_29635);
and UO_450 (O_450,N_29470,N_29343);
and UO_451 (O_451,N_29921,N_26537);
nor UO_452 (O_452,N_26190,N_26429);
or UO_453 (O_453,N_29617,N_27068);
nand UO_454 (O_454,N_26051,N_29396);
nand UO_455 (O_455,N_26457,N_27976);
or UO_456 (O_456,N_27908,N_28153);
or UO_457 (O_457,N_26297,N_26596);
nand UO_458 (O_458,N_29811,N_27703);
or UO_459 (O_459,N_28950,N_28426);
or UO_460 (O_460,N_25296,N_25336);
nand UO_461 (O_461,N_29685,N_27822);
nand UO_462 (O_462,N_25222,N_27138);
nand UO_463 (O_463,N_26237,N_26539);
or UO_464 (O_464,N_27693,N_28197);
and UO_465 (O_465,N_28446,N_27421);
nor UO_466 (O_466,N_26613,N_27710);
or UO_467 (O_467,N_26894,N_29605);
nor UO_468 (O_468,N_26634,N_29613);
nand UO_469 (O_469,N_26743,N_26154);
nand UO_470 (O_470,N_29101,N_29001);
or UO_471 (O_471,N_26212,N_28242);
and UO_472 (O_472,N_26364,N_25671);
and UO_473 (O_473,N_25314,N_28559);
nor UO_474 (O_474,N_27102,N_27914);
nor UO_475 (O_475,N_25648,N_28630);
nor UO_476 (O_476,N_27967,N_28442);
or UO_477 (O_477,N_28694,N_27600);
or UO_478 (O_478,N_28863,N_26723);
nor UO_479 (O_479,N_25347,N_25618);
nor UO_480 (O_480,N_26225,N_27122);
nor UO_481 (O_481,N_25984,N_26661);
or UO_482 (O_482,N_28570,N_27019);
xnor UO_483 (O_483,N_27390,N_25127);
nor UO_484 (O_484,N_26006,N_26652);
or UO_485 (O_485,N_26503,N_26127);
or UO_486 (O_486,N_25016,N_26148);
nor UO_487 (O_487,N_29246,N_29621);
or UO_488 (O_488,N_29298,N_29902);
nand UO_489 (O_489,N_28671,N_25825);
nand UO_490 (O_490,N_29598,N_25403);
nand UO_491 (O_491,N_29286,N_25809);
and UO_492 (O_492,N_28175,N_29031);
or UO_493 (O_493,N_29171,N_25968);
nand UO_494 (O_494,N_27011,N_25576);
nand UO_495 (O_495,N_27269,N_29631);
and UO_496 (O_496,N_28755,N_28947);
and UO_497 (O_497,N_27005,N_29595);
or UO_498 (O_498,N_27891,N_26713);
nor UO_499 (O_499,N_27423,N_29644);
nor UO_500 (O_500,N_29591,N_26425);
or UO_501 (O_501,N_28684,N_27351);
and UO_502 (O_502,N_26996,N_29095);
nor UO_503 (O_503,N_28822,N_27530);
xor UO_504 (O_504,N_26373,N_25495);
nand UO_505 (O_505,N_25869,N_25523);
and UO_506 (O_506,N_29218,N_29846);
and UO_507 (O_507,N_28703,N_25947);
and UO_508 (O_508,N_29227,N_27177);
and UO_509 (O_509,N_25729,N_26551);
and UO_510 (O_510,N_25276,N_28436);
or UO_511 (O_511,N_29481,N_28757);
and UO_512 (O_512,N_25530,N_27875);
nand UO_513 (O_513,N_28759,N_27082);
nor UO_514 (O_514,N_26455,N_25298);
nor UO_515 (O_515,N_25538,N_28716);
nor UO_516 (O_516,N_26625,N_27147);
nand UO_517 (O_517,N_28250,N_26793);
and UO_518 (O_518,N_27596,N_26406);
and UO_519 (O_519,N_27149,N_25129);
nor UO_520 (O_520,N_29962,N_29992);
nand UO_521 (O_521,N_25675,N_27145);
nand UO_522 (O_522,N_27569,N_25751);
or UO_523 (O_523,N_28557,N_28166);
or UO_524 (O_524,N_27708,N_27768);
nand UO_525 (O_525,N_26204,N_29321);
and UO_526 (O_526,N_27874,N_29989);
or UO_527 (O_527,N_29086,N_25292);
nor UO_528 (O_528,N_28553,N_26236);
and UO_529 (O_529,N_26927,N_28116);
nor UO_530 (O_530,N_27685,N_28163);
and UO_531 (O_531,N_27095,N_29147);
nor UO_532 (O_532,N_27289,N_29972);
nor UO_533 (O_533,N_28654,N_28807);
nor UO_534 (O_534,N_29920,N_26309);
or UO_535 (O_535,N_28848,N_29288);
nand UO_536 (O_536,N_29525,N_28942);
and UO_537 (O_537,N_25044,N_25519);
nor UO_538 (O_538,N_25216,N_29694);
and UO_539 (O_539,N_27312,N_27741);
or UO_540 (O_540,N_29889,N_29381);
nor UO_541 (O_541,N_28727,N_29016);
and UO_542 (O_542,N_29616,N_25818);
nor UO_543 (O_543,N_25261,N_27199);
or UO_544 (O_544,N_27369,N_26925);
nand UO_545 (O_545,N_26343,N_27645);
nor UO_546 (O_546,N_28750,N_29746);
and UO_547 (O_547,N_28211,N_29200);
nand UO_548 (O_548,N_27112,N_25234);
and UO_549 (O_549,N_28369,N_29484);
and UO_550 (O_550,N_25505,N_25194);
and UO_551 (O_551,N_25225,N_29380);
nand UO_552 (O_552,N_28162,N_26134);
and UO_553 (O_553,N_27894,N_25978);
or UO_554 (O_554,N_27518,N_29500);
nor UO_555 (O_555,N_26171,N_25798);
nor UO_556 (O_556,N_26502,N_27012);
or UO_557 (O_557,N_25186,N_25326);
and UO_558 (O_558,N_25082,N_28429);
or UO_559 (O_559,N_28386,N_27613);
nor UO_560 (O_560,N_29727,N_26695);
nand UO_561 (O_561,N_25188,N_29659);
or UO_562 (O_562,N_29626,N_28994);
and UO_563 (O_563,N_26850,N_29540);
or UO_564 (O_564,N_29255,N_29344);
and UO_565 (O_565,N_25867,N_29820);
nor UO_566 (O_566,N_29010,N_29538);
and UO_567 (O_567,N_28118,N_25649);
and UO_568 (O_568,N_29984,N_28833);
nand UO_569 (O_569,N_25785,N_25299);
and UO_570 (O_570,N_29041,N_25760);
or UO_571 (O_571,N_29331,N_28229);
nor UO_572 (O_572,N_28884,N_25476);
nor UO_573 (O_573,N_27512,N_27563);
nor UO_574 (O_574,N_26623,N_25783);
xor UO_575 (O_575,N_25117,N_29796);
nor UO_576 (O_576,N_28107,N_29136);
nor UO_577 (O_577,N_28178,N_27856);
and UO_578 (O_578,N_28157,N_26708);
nor UO_579 (O_579,N_25927,N_25274);
and UO_580 (O_580,N_29006,N_25775);
nor UO_581 (O_581,N_28238,N_27970);
nor UO_582 (O_582,N_28845,N_27244);
or UO_583 (O_583,N_27843,N_28733);
and UO_584 (O_584,N_25696,N_27290);
and UO_585 (O_585,N_25952,N_29352);
nand UO_586 (O_586,N_28679,N_29349);
nor UO_587 (O_587,N_27036,N_26078);
nor UO_588 (O_588,N_28626,N_28122);
and UO_589 (O_589,N_29979,N_26246);
nor UO_590 (O_590,N_26875,N_25118);
nand UO_591 (O_591,N_29698,N_27920);
nand UO_592 (O_592,N_26340,N_27607);
and UO_593 (O_593,N_27537,N_29747);
nand UO_594 (O_594,N_29389,N_29761);
and UO_595 (O_595,N_26783,N_25628);
nor UO_596 (O_596,N_25714,N_25778);
and UO_597 (O_597,N_26143,N_27898);
nor UO_598 (O_598,N_27411,N_29109);
nand UO_599 (O_599,N_28875,N_29182);
nand UO_600 (O_600,N_28561,N_26568);
and UO_601 (O_601,N_29448,N_27481);
nand UO_602 (O_602,N_26563,N_27884);
nor UO_603 (O_603,N_26140,N_29662);
xor UO_604 (O_604,N_27928,N_28047);
or UO_605 (O_605,N_26419,N_26928);
nor UO_606 (O_606,N_27339,N_26291);
or UO_607 (O_607,N_27140,N_29600);
or UO_608 (O_608,N_28610,N_28963);
and UO_609 (O_609,N_25050,N_28151);
or UO_610 (O_610,N_25287,N_28349);
and UO_611 (O_611,N_25126,N_26735);
and UO_612 (O_612,N_25932,N_25712);
nor UO_613 (O_613,N_29541,N_27853);
and UO_614 (O_614,N_28605,N_25722);
nor UO_615 (O_615,N_28902,N_28535);
or UO_616 (O_616,N_27458,N_28551);
or UO_617 (O_617,N_25553,N_29637);
nand UO_618 (O_618,N_25380,N_29640);
nand UO_619 (O_619,N_29511,N_27628);
nand UO_620 (O_620,N_27505,N_25625);
nor UO_621 (O_621,N_26296,N_25811);
nand UO_622 (O_622,N_26552,N_26192);
nor UO_623 (O_623,N_25684,N_28234);
and UO_624 (O_624,N_28965,N_26177);
and UO_625 (O_625,N_27889,N_25419);
or UO_626 (O_626,N_29356,N_27077);
and UO_627 (O_627,N_29252,N_29247);
and UO_628 (O_628,N_27373,N_25685);
nand UO_629 (O_629,N_25247,N_27398);
and UO_630 (O_630,N_27392,N_27432);
nor UO_631 (O_631,N_26277,N_28734);
nor UO_632 (O_632,N_29993,N_29765);
nand UO_633 (O_633,N_27930,N_28554);
and UO_634 (O_634,N_27559,N_26322);
and UO_635 (O_635,N_29899,N_29742);
nand UO_636 (O_636,N_29083,N_26161);
nor UO_637 (O_637,N_27525,N_29975);
or UO_638 (O_638,N_29722,N_29797);
or UO_639 (O_639,N_26853,N_27280);
nand UO_640 (O_640,N_28740,N_27611);
or UO_641 (O_641,N_29868,N_28585);
nor UO_642 (O_642,N_28794,N_28039);
and UO_643 (O_643,N_25526,N_29622);
nand UO_644 (O_644,N_26170,N_29887);
and UO_645 (O_645,N_27841,N_27796);
and UO_646 (O_646,N_28080,N_25423);
and UO_647 (O_647,N_26580,N_27862);
or UO_648 (O_648,N_25999,N_25048);
nand UO_649 (O_649,N_25847,N_28279);
and UO_650 (O_650,N_25085,N_27355);
and UO_651 (O_651,N_28672,N_29731);
nor UO_652 (O_652,N_26433,N_26348);
nor UO_653 (O_653,N_27802,N_26053);
nand UO_654 (O_654,N_28592,N_29058);
or UO_655 (O_655,N_25972,N_28129);
nor UO_656 (O_656,N_25100,N_29823);
nor UO_657 (O_657,N_27778,N_29625);
nand UO_658 (O_658,N_28051,N_28636);
or UO_659 (O_659,N_26112,N_26389);
nor UO_660 (O_660,N_28777,N_25400);
nor UO_661 (O_661,N_29229,N_29044);
nand UO_662 (O_662,N_25269,N_26464);
nand UO_663 (O_663,N_27382,N_29213);
nand UO_664 (O_664,N_27069,N_26102);
nor UO_665 (O_665,N_27288,N_28056);
or UO_666 (O_666,N_28384,N_28662);
or UO_667 (O_667,N_28292,N_27193);
nor UO_668 (O_668,N_26666,N_25704);
or UO_669 (O_669,N_27041,N_26440);
nor UO_670 (O_670,N_28133,N_29814);
nand UO_671 (O_671,N_27434,N_25349);
or UO_672 (O_672,N_29825,N_29148);
or UO_673 (O_673,N_29176,N_25754);
xor UO_674 (O_674,N_28539,N_26870);
and UO_675 (O_675,N_25393,N_25427);
nor UO_676 (O_676,N_28365,N_25563);
nand UO_677 (O_677,N_25404,N_28323);
or UO_678 (O_678,N_27376,N_27996);
nand UO_679 (O_679,N_29589,N_25945);
nor UO_680 (O_680,N_28915,N_25919);
nor UO_681 (O_681,N_27038,N_26426);
nor UO_682 (O_682,N_27086,N_29592);
nor UO_683 (O_683,N_28035,N_25464);
nand UO_684 (O_684,N_25189,N_27080);
and UO_685 (O_685,N_25732,N_28784);
or UO_686 (O_686,N_25521,N_25145);
and UO_687 (O_687,N_29582,N_26131);
nor UO_688 (O_688,N_25334,N_26361);
or UO_689 (O_689,N_28643,N_27932);
nand UO_690 (O_690,N_28158,N_26873);
nand UO_691 (O_691,N_26060,N_29638);
nor UO_692 (O_692,N_27630,N_27709);
nor UO_693 (O_693,N_25068,N_27877);
nor UO_694 (O_694,N_29910,N_25376);
or UO_695 (O_695,N_29335,N_27949);
or UO_696 (O_696,N_29019,N_28248);
and UO_697 (O_697,N_29674,N_25665);
nor UO_698 (O_698,N_27599,N_27723);
nor UO_699 (O_699,N_28251,N_28849);
nor UO_700 (O_700,N_26653,N_28825);
or UO_701 (O_701,N_25929,N_28960);
or UO_702 (O_702,N_29451,N_28019);
or UO_703 (O_703,N_28457,N_29264);
nand UO_704 (O_704,N_25148,N_29168);
and UO_705 (O_705,N_26919,N_25875);
nor UO_706 (O_706,N_29560,N_28231);
or UO_707 (O_707,N_26488,N_26579);
or UO_708 (O_708,N_26349,N_27324);
and UO_709 (O_709,N_26266,N_26508);
or UO_710 (O_710,N_25957,N_25333);
or UO_711 (O_711,N_28492,N_26981);
nor UO_712 (O_712,N_25417,N_27321);
nor UO_713 (O_713,N_29021,N_25654);
and UO_714 (O_714,N_27766,N_29454);
or UO_715 (O_715,N_27251,N_27531);
nor UO_716 (O_716,N_27584,N_29280);
nand UO_717 (O_717,N_27389,N_29287);
nor UO_718 (O_718,N_25904,N_28859);
nor UO_719 (O_719,N_26932,N_26615);
nor UO_720 (O_720,N_26827,N_27574);
nand UO_721 (O_721,N_27101,N_29568);
nor UO_722 (O_722,N_28299,N_28346);
and UO_723 (O_723,N_29877,N_29602);
nand UO_724 (O_724,N_28444,N_29943);
or UO_725 (O_725,N_29918,N_26618);
nand UO_726 (O_726,N_28943,N_27444);
or UO_727 (O_727,N_27632,N_25747);
nor UO_728 (O_728,N_26282,N_26662);
and UO_729 (O_729,N_26318,N_27325);
and UO_730 (O_730,N_29440,N_28753);
nand UO_731 (O_731,N_28432,N_26116);
nand UO_732 (O_732,N_26958,N_27327);
and UO_733 (O_733,N_25446,N_27756);
and UO_734 (O_734,N_27590,N_28670);
or UO_735 (O_735,N_27261,N_27178);
or UO_736 (O_736,N_25557,N_29004);
and UO_737 (O_737,N_25395,N_27230);
or UO_738 (O_738,N_29951,N_28053);
or UO_739 (O_739,N_29313,N_25692);
nand UO_740 (O_740,N_28698,N_26145);
or UO_741 (O_741,N_27275,N_26578);
nor UO_742 (O_742,N_27202,N_25275);
nand UO_743 (O_743,N_25037,N_25004);
nand UO_744 (O_744,N_26394,N_28860);
or UO_745 (O_745,N_25367,N_25969);
and UO_746 (O_746,N_29383,N_27477);
nand UO_747 (O_747,N_28066,N_27568);
and UO_748 (O_748,N_29278,N_28507);
and UO_749 (O_749,N_28600,N_29111);
and UO_750 (O_750,N_27320,N_25727);
nand UO_751 (O_751,N_27186,N_25116);
nor UO_752 (O_752,N_28409,N_25500);
and UO_753 (O_753,N_27963,N_25250);
or UO_754 (O_754,N_29710,N_28593);
and UO_755 (O_755,N_29520,N_25529);
nand UO_756 (O_756,N_29117,N_26989);
and UO_757 (O_757,N_27591,N_28497);
nor UO_758 (O_758,N_25995,N_25280);
nor UO_759 (O_759,N_28885,N_28338);
and UO_760 (O_760,N_29854,N_28601);
nand UO_761 (O_761,N_27179,N_26706);
xnor UO_762 (O_762,N_25909,N_29150);
or UO_763 (O_763,N_27226,N_28459);
nand UO_764 (O_764,N_26586,N_27135);
xor UO_765 (O_765,N_27765,N_26311);
or UO_766 (O_766,N_28665,N_28691);
and UO_767 (O_767,N_26481,N_26822);
or UO_768 (O_768,N_26790,N_25089);
and UO_769 (O_769,N_27385,N_25015);
nor UO_770 (O_770,N_27375,N_27808);
nor UO_771 (O_771,N_25622,N_25152);
nor UO_772 (O_772,N_28961,N_26554);
nor UO_773 (O_773,N_26251,N_27529);
nor UO_774 (O_774,N_27381,N_26705);
or UO_775 (O_775,N_26681,N_27256);
nor UO_776 (O_776,N_26617,N_26016);
and UO_777 (O_777,N_26949,N_27453);
and UO_778 (O_778,N_26628,N_28854);
nand UO_779 (O_779,N_28966,N_25734);
or UO_780 (O_780,N_26179,N_25439);
or UO_781 (O_781,N_27260,N_28044);
or UO_782 (O_782,N_27840,N_29374);
nor UO_783 (O_783,N_26858,N_26125);
and UO_784 (O_784,N_27990,N_25220);
or UO_785 (O_785,N_28180,N_25407);
nand UO_786 (O_786,N_29359,N_28233);
nor UO_787 (O_787,N_28031,N_29897);
or UO_788 (O_788,N_29729,N_27727);
or UO_789 (O_789,N_25977,N_26438);
and UO_790 (O_790,N_27706,N_25724);
nor UO_791 (O_791,N_25819,N_26259);
or UO_792 (O_792,N_25573,N_26972);
or UO_793 (O_793,N_29183,N_29898);
nand UO_794 (O_794,N_28106,N_29682);
and UO_795 (O_795,N_26453,N_25872);
nor UO_796 (O_796,N_29408,N_29935);
nand UO_797 (O_797,N_28685,N_26986);
or UO_798 (O_798,N_25537,N_29522);
or UO_799 (O_799,N_28844,N_28435);
or UO_800 (O_800,N_29196,N_26521);
or UO_801 (O_801,N_28828,N_25497);
or UO_802 (O_802,N_27922,N_29648);
nand UO_803 (O_803,N_26441,N_26206);
or UO_804 (O_804,N_29000,N_25599);
nor UO_805 (O_805,N_26505,N_27400);
or UO_806 (O_806,N_28664,N_25916);
or UO_807 (O_807,N_27331,N_26274);
or UO_808 (O_808,N_26805,N_28059);
or UO_809 (O_809,N_25803,N_29347);
nor UO_810 (O_810,N_27006,N_28953);
nand UO_811 (O_811,N_28098,N_29061);
and UO_812 (O_812,N_25003,N_25243);
nor UO_813 (O_813,N_25239,N_27698);
nor UO_814 (O_814,N_27833,N_25981);
nand UO_815 (O_815,N_28326,N_28775);
and UO_816 (O_816,N_26040,N_26534);
xor UO_817 (O_817,N_28919,N_26435);
and UO_818 (O_818,N_29961,N_29963);
nor UO_819 (O_819,N_28661,N_28909);
nand UO_820 (O_820,N_27806,N_28687);
and UO_821 (O_821,N_26347,N_29162);
or UO_822 (O_822,N_27746,N_28900);
nor UO_823 (O_823,N_27999,N_29431);
nor UO_824 (O_824,N_29769,N_25207);
and UO_825 (O_825,N_27418,N_28154);
or UO_826 (O_826,N_29620,N_27948);
and UO_827 (O_827,N_29566,N_27605);
nand UO_828 (O_828,N_28341,N_26982);
nand UO_829 (O_829,N_27745,N_26470);
nand UO_830 (O_830,N_28914,N_25743);
nand UO_831 (O_831,N_28453,N_28227);
and UO_832 (O_832,N_29467,N_28316);
nor UO_833 (O_833,N_29211,N_27832);
and UO_834 (O_834,N_28751,N_26840);
nand UO_835 (O_835,N_29896,N_27728);
nor UO_836 (O_836,N_28124,N_26402);
nor UO_837 (O_837,N_27446,N_26178);
nor UO_838 (O_838,N_27460,N_28990);
nor UO_839 (O_839,N_28646,N_29253);
or UO_840 (O_840,N_25876,N_26019);
nand UO_841 (O_841,N_25156,N_28222);
nor UO_842 (O_842,N_26393,N_25154);
nand UO_843 (O_843,N_29725,N_25249);
nor UO_844 (O_844,N_28455,N_28374);
or UO_845 (O_845,N_25300,N_27826);
nand UO_846 (O_846,N_27795,N_25485);
nand UO_847 (O_847,N_25676,N_25934);
nor UO_848 (O_848,N_27044,N_28544);
or UO_849 (O_849,N_29874,N_25366);
nor UO_850 (O_850,N_29726,N_29488);
or UO_851 (O_851,N_28113,N_28441);
and UO_852 (O_852,N_29988,N_29575);
or UO_853 (O_853,N_27824,N_28588);
nor UO_854 (O_854,N_29552,N_29609);
nor UO_855 (O_855,N_27522,N_27116);
and UO_856 (O_856,N_25210,N_25378);
or UO_857 (O_857,N_27555,N_26895);
and UO_858 (O_858,N_26592,N_27049);
xor UO_859 (O_859,N_25894,N_28389);
nand UO_860 (O_860,N_29784,N_27702);
or UO_861 (O_861,N_25242,N_28752);
or UO_862 (O_862,N_25679,N_29003);
nor UO_863 (O_863,N_25583,N_25470);
nand UO_864 (O_864,N_27544,N_29557);
and UO_865 (O_865,N_29390,N_28851);
nor UO_866 (O_866,N_27194,N_25093);
nand UO_867 (O_867,N_27328,N_29173);
or UO_868 (O_868,N_26930,N_25340);
or UO_869 (O_869,N_29934,N_29733);
and UO_870 (O_870,N_29741,N_26562);
nand UO_871 (O_871,N_26475,N_29929);
nand UO_872 (O_872,N_28602,N_25569);
nor UO_873 (O_873,N_27573,N_28944);
and UO_874 (O_874,N_26385,N_27831);
and UO_875 (O_875,N_29906,N_25660);
and UO_876 (O_876,N_26542,N_29015);
nand UO_877 (O_877,N_26794,N_26907);
and UO_878 (O_878,N_28280,N_26988);
or UO_879 (O_879,N_27263,N_29461);
nand UO_880 (O_880,N_25752,N_29224);
or UO_881 (O_881,N_28484,N_25346);
nor UO_882 (O_882,N_25964,N_27887);
or UO_883 (O_883,N_26522,N_26800);
or UO_884 (O_884,N_27281,N_28028);
nand UO_885 (O_885,N_27769,N_25203);
nor UO_886 (O_886,N_28847,N_26704);
nand UO_887 (O_887,N_25240,N_25603);
or UO_888 (O_888,N_26594,N_29005);
nand UO_889 (O_889,N_29869,N_29317);
or UO_890 (O_890,N_26249,N_26730);
or UO_891 (O_891,N_27359,N_26533);
and UO_892 (O_892,N_25866,N_25960);
or UO_893 (O_893,N_29054,N_25914);
nor UO_894 (O_894,N_26381,N_26081);
nand UO_895 (O_895,N_28291,N_29145);
or UO_896 (O_896,N_26770,N_26825);
nor UO_897 (O_897,N_29368,N_27786);
or UO_898 (O_898,N_26321,N_25480);
nand UO_899 (O_899,N_29543,N_28808);
nand UO_900 (O_900,N_29832,N_25549);
or UO_901 (O_901,N_28583,N_28219);
nand UO_902 (O_902,N_29954,N_28266);
nand UO_903 (O_903,N_28976,N_27692);
and UO_904 (O_904,N_28795,N_25028);
and UO_905 (O_905,N_25060,N_27878);
and UO_906 (O_906,N_27975,N_25328);
nor UO_907 (O_907,N_29842,N_26331);
or UO_908 (O_908,N_29803,N_27652);
and UO_909 (O_909,N_25244,N_28818);
or UO_910 (O_910,N_27743,N_29753);
nor UO_911 (O_911,N_29158,N_29257);
and UO_912 (O_912,N_25918,N_29822);
or UO_913 (O_913,N_28528,N_26223);
nand UO_914 (O_914,N_26693,N_26446);
nor UO_915 (O_915,N_27435,N_28934);
or UO_916 (O_916,N_26077,N_25416);
or UO_917 (O_917,N_29704,N_28256);
nand UO_918 (O_918,N_25744,N_28852);
and UO_919 (O_919,N_25475,N_29093);
or UO_920 (O_920,N_26380,N_28489);
nor UO_921 (O_921,N_29275,N_29155);
and UO_922 (O_922,N_26276,N_25176);
or UO_923 (O_923,N_28301,N_25657);
nor UO_924 (O_924,N_25221,N_29203);
nand UO_925 (O_925,N_28075,N_26199);
nor UO_926 (O_926,N_27397,N_27307);
nor UO_927 (O_927,N_27731,N_29342);
nand UO_928 (O_928,N_28657,N_25024);
nand UO_929 (O_929,N_27098,N_29892);
nor UO_930 (O_930,N_27143,N_28878);
and UO_931 (O_931,N_26630,N_26672);
nor UO_932 (O_932,N_27232,N_29394);
and UO_933 (O_933,N_25312,N_28464);
and UO_934 (O_934,N_27620,N_28102);
or UO_935 (O_935,N_25609,N_29692);
nand UO_936 (O_936,N_27103,N_27258);
or UO_937 (O_937,N_25008,N_25920);
nor UO_938 (O_938,N_26320,N_25365);
nand UO_939 (O_939,N_26138,N_28991);
or UO_940 (O_940,N_27609,N_26621);
or UO_941 (O_941,N_28355,N_28725);
nand UO_942 (O_942,N_26629,N_27195);
nor UO_943 (O_943,N_28835,N_29762);
nor UO_944 (O_944,N_29133,N_27661);
and UO_945 (O_945,N_25073,N_27665);
or UO_946 (O_946,N_28566,N_28300);
or UO_947 (O_947,N_28771,N_27836);
nor UO_948 (O_948,N_26655,N_26208);
or UO_949 (O_949,N_26191,N_28836);
and UO_950 (O_950,N_28631,N_25000);
nand UO_951 (O_951,N_25578,N_25436);
nand UO_952 (O_952,N_25432,N_27773);
nor UO_953 (O_953,N_25159,N_26113);
nand UO_954 (O_954,N_27964,N_25528);
nor UO_955 (O_955,N_28311,N_27777);
and UO_956 (O_956,N_27189,N_29324);
nor UO_957 (O_957,N_27602,N_28534);
or UO_958 (O_958,N_26998,N_29103);
or UO_959 (O_959,N_26480,N_29404);
nand UO_960 (O_960,N_25580,N_28842);
nand UO_961 (O_961,N_28550,N_25917);
and UO_962 (O_962,N_29501,N_25149);
and UO_963 (O_963,N_25058,N_26602);
nand UO_964 (O_964,N_28837,N_25049);
nand UO_965 (O_965,N_29315,N_29661);
nor UO_966 (O_966,N_28772,N_29065);
nor UO_967 (O_967,N_29367,N_25780);
and UO_968 (O_968,N_29684,N_27549);
xnor UO_969 (O_969,N_29032,N_26195);
nand UO_970 (O_970,N_29956,N_29238);
or UO_971 (O_971,N_27021,N_28547);
nor UO_972 (O_972,N_26961,N_29867);
or UO_973 (O_973,N_28603,N_28026);
nor UO_974 (O_974,N_25504,N_26779);
or UO_975 (O_975,N_27167,N_27386);
nor UO_976 (O_976,N_28660,N_29131);
nand UO_977 (O_977,N_29947,N_27165);
or UO_978 (O_978,N_26577,N_25971);
nand UO_979 (O_979,N_27648,N_27306);
or UO_980 (O_980,N_27551,N_27264);
or UO_981 (O_981,N_27821,N_27310);
and UO_982 (O_982,N_27694,N_28278);
nand UO_983 (O_983,N_28295,N_27699);
or UO_984 (O_984,N_25437,N_28317);
nor UO_985 (O_985,N_28992,N_29376);
nor UO_986 (O_986,N_29715,N_28115);
nand UO_987 (O_987,N_26549,N_29489);
or UO_988 (O_988,N_27861,N_28812);
nand UO_989 (O_989,N_26205,N_25033);
and UO_990 (O_990,N_27142,N_29248);
and UO_991 (O_991,N_26129,N_28834);
or UO_992 (O_992,N_29847,N_27911);
and UO_993 (O_993,N_28741,N_27755);
and UO_994 (O_994,N_28452,N_26287);
and UO_995 (O_995,N_27931,N_29293);
nand UO_996 (O_996,N_28579,N_27528);
nor UO_997 (O_997,N_26872,N_27634);
or UO_998 (O_998,N_26467,N_28615);
nand UO_999 (O_999,N_25939,N_28050);
or UO_1000 (O_1000,N_25858,N_28325);
or UO_1001 (O_1001,N_26795,N_26144);
nor UO_1002 (O_1002,N_28070,N_26009);
or UO_1003 (O_1003,N_26350,N_27126);
or UO_1004 (O_1004,N_29785,N_26564);
nor UO_1005 (O_1005,N_27978,N_25106);
nor UO_1006 (O_1006,N_28281,N_25717);
and UO_1007 (O_1007,N_27203,N_29756);
nand UO_1008 (O_1008,N_29529,N_28273);
nor UO_1009 (O_1009,N_25350,N_29076);
nand UO_1010 (O_1010,N_26119,N_28531);
and UO_1011 (O_1011,N_25518,N_29070);
and UO_1012 (O_1012,N_29423,N_25291);
nor UO_1013 (O_1013,N_26565,N_25229);
nand UO_1014 (O_1014,N_29804,N_26823);
nor UO_1015 (O_1015,N_25499,N_27393);
or UO_1016 (O_1016,N_25838,N_27788);
and UO_1017 (O_1017,N_25762,N_28587);
and UO_1018 (O_1018,N_26526,N_28538);
nor UO_1019 (O_1019,N_27183,N_26359);
nor UO_1020 (O_1020,N_26891,N_25305);
nor UO_1021 (O_1021,N_25398,N_25111);
and UO_1022 (O_1022,N_27638,N_29455);
and UO_1023 (O_1023,N_28078,N_26657);
nand UO_1024 (O_1024,N_28009,N_26889);
nand UO_1025 (O_1025,N_26405,N_28037);
and UO_1026 (O_1026,N_28486,N_26392);
nand UO_1027 (O_1027,N_29793,N_29140);
or UO_1028 (O_1028,N_29748,N_29351);
nand UO_1029 (O_1029,N_29370,N_26036);
nand UO_1030 (O_1030,N_25993,N_25443);
or UO_1031 (O_1031,N_26740,N_26056);
nand UO_1032 (O_1032,N_29881,N_29789);
or UO_1033 (O_1033,N_25982,N_29444);
or UO_1034 (O_1034,N_29296,N_28673);
and UO_1035 (O_1035,N_27031,N_29503);
nor UO_1036 (O_1036,N_29928,N_29456);
or UO_1037 (O_1037,N_27762,N_26772);
nand UO_1038 (O_1038,N_26240,N_26627);
nor UO_1039 (O_1039,N_29276,N_27115);
and UO_1040 (O_1040,N_29403,N_28117);
nand UO_1041 (O_1041,N_25897,N_27988);
nor UO_1042 (O_1042,N_26697,N_29615);
nor UO_1043 (O_1043,N_26581,N_29815);
nand UO_1044 (O_1044,N_25489,N_29328);
or UO_1045 (O_1045,N_26202,N_27033);
nor UO_1046 (O_1046,N_27747,N_28096);
xor UO_1047 (O_1047,N_28666,N_27083);
nor UO_1048 (O_1048,N_28148,N_27188);
nor UO_1049 (O_1049,N_25817,N_28177);
and UO_1050 (O_1050,N_28708,N_25449);
or UO_1051 (O_1051,N_28285,N_25236);
xnor UO_1052 (O_1052,N_29371,N_25949);
nand UO_1053 (O_1053,N_28695,N_27730);
nor UO_1054 (O_1054,N_25900,N_26999);
or UO_1055 (O_1055,N_28171,N_29909);
nor UO_1056 (O_1056,N_25612,N_25986);
and UO_1057 (O_1057,N_29023,N_25162);
nand UO_1058 (O_1058,N_26386,N_25565);
or UO_1059 (O_1059,N_26304,N_26216);
nand UO_1060 (O_1060,N_27410,N_27586);
nor UO_1061 (O_1061,N_27299,N_28013);
nand UO_1062 (O_1062,N_29310,N_25130);
and UO_1063 (O_1063,N_27007,N_27368);
nand UO_1064 (O_1064,N_27344,N_26656);
nor UO_1065 (O_1065,N_29713,N_25386);
xnor UO_1066 (O_1066,N_28514,N_26075);
nor UO_1067 (O_1067,N_26369,N_28933);
nand UO_1068 (O_1068,N_26523,N_26885);
xnor UO_1069 (O_1069,N_27475,N_25815);
and UO_1070 (O_1070,N_28591,N_29189);
nor UO_1071 (O_1071,N_29039,N_27034);
and UO_1072 (O_1072,N_25703,N_29024);
nand UO_1073 (O_1073,N_28581,N_27152);
nand UO_1074 (O_1074,N_26905,N_27303);
nand UO_1075 (O_1075,N_26409,N_27278);
nor UO_1076 (O_1076,N_29400,N_29068);
nand UO_1077 (O_1077,N_27587,N_27919);
nor UO_1078 (O_1078,N_26494,N_25746);
or UO_1079 (O_1079,N_26018,N_27686);
nand UO_1080 (O_1080,N_29027,N_27532);
nor UO_1081 (O_1081,N_25757,N_28241);
nor UO_1082 (O_1082,N_25921,N_25520);
nor UO_1083 (O_1083,N_26235,N_27637);
and UO_1084 (O_1084,N_26954,N_25555);
or UO_1085 (O_1085,N_27114,N_29740);
nand UO_1086 (O_1086,N_29236,N_27733);
nand UO_1087 (O_1087,N_27997,N_28003);
and UO_1088 (O_1088,N_29764,N_26482);
or UO_1089 (O_1089,N_26132,N_27065);
nand UO_1090 (O_1090,N_27940,N_29870);
nor UO_1091 (O_1091,N_29721,N_28141);
and UO_1092 (O_1092,N_28895,N_29479);
or UO_1093 (O_1093,N_26074,N_25516);
nor UO_1094 (O_1094,N_29561,N_26936);
or UO_1095 (O_1095,N_28368,N_25823);
nor UO_1096 (O_1096,N_25796,N_28074);
nor UO_1097 (O_1097,N_29063,N_25257);
nand UO_1098 (O_1098,N_27029,N_26501);
nand UO_1099 (O_1099,N_27500,N_28552);
and UO_1100 (O_1100,N_29940,N_25339);
or UO_1101 (O_1101,N_28642,N_26404);
nor UO_1102 (O_1102,N_28555,N_28726);
nor UO_1103 (O_1103,N_25619,N_25201);
nand UO_1104 (O_1104,N_27054,N_29297);
xor UO_1105 (O_1105,N_28343,N_26940);
nor UO_1106 (O_1106,N_28088,N_28411);
or UO_1107 (O_1107,N_29521,N_26869);
and UO_1108 (O_1108,N_25071,N_29755);
and UO_1109 (O_1109,N_27669,N_25721);
or UO_1110 (O_1110,N_28618,N_27255);
nand UO_1111 (O_1111,N_28530,N_29596);
nor UO_1112 (O_1112,N_25218,N_29355);
nor UO_1113 (O_1113,N_26215,N_29379);
nand UO_1114 (O_1114,N_25105,N_28342);
and UO_1115 (O_1115,N_27986,N_27516);
and UO_1116 (O_1116,N_27413,N_27357);
nand UO_1117 (O_1117,N_27234,N_28306);
nand UO_1118 (O_1118,N_25248,N_26504);
nand UO_1119 (O_1119,N_29821,N_29469);
nand UO_1120 (O_1120,N_27811,N_26611);
nor UO_1121 (O_1121,N_27957,N_29337);
and UO_1122 (O_1122,N_27903,N_29208);
or UO_1123 (O_1123,N_29673,N_25381);
and UO_1124 (O_1124,N_27117,N_25786);
nand UO_1125 (O_1125,N_27465,N_27880);
or UO_1126 (O_1126,N_25341,N_25535);
xor UO_1127 (O_1127,N_28179,N_25109);
nor UO_1128 (O_1128,N_27576,N_29530);
and UO_1129 (O_1129,N_25539,N_28428);
and UO_1130 (O_1130,N_27025,N_27295);
xnor UO_1131 (O_1131,N_28193,N_26007);
nor UO_1132 (O_1132,N_26947,N_28005);
nor UO_1133 (O_1133,N_27047,N_29593);
nand UO_1134 (O_1134,N_25051,N_26151);
nor UO_1135 (O_1135,N_29364,N_28941);
and UO_1136 (O_1136,N_29205,N_27317);
nor UO_1137 (O_1137,N_25463,N_27156);
nor UO_1138 (O_1138,N_25951,N_28758);
nand UO_1139 (O_1139,N_26509,N_25546);
and UO_1140 (O_1140,N_27863,N_27774);
and UO_1141 (O_1141,N_29146,N_28651);
nor UO_1142 (O_1142,N_26841,N_26310);
or UO_1143 (O_1143,N_27895,N_28265);
and UO_1144 (O_1144,N_28144,N_25473);
nor UO_1145 (O_1145,N_26754,N_27944);
nand UO_1146 (O_1146,N_29657,N_27960);
nand UO_1147 (O_1147,N_29363,N_28111);
nor UO_1148 (O_1148,N_25942,N_29327);
or UO_1149 (O_1149,N_28109,N_28025);
or UO_1150 (O_1150,N_26638,N_28033);
nand UO_1151 (O_1151,N_25868,N_28319);
nand UO_1152 (O_1152,N_26432,N_27236);
and UO_1153 (O_1153,N_29079,N_25133);
nand UO_1154 (O_1154,N_28399,N_28469);
nand UO_1155 (O_1155,N_26864,N_25506);
nand UO_1156 (O_1156,N_29274,N_26558);
nand UO_1157 (O_1157,N_26345,N_26300);
or UO_1158 (O_1158,N_29018,N_25488);
or UO_1159 (O_1159,N_29165,N_29573);
nand UO_1160 (O_1160,N_26828,N_26400);
nand UO_1161 (O_1161,N_28239,N_28987);
and UO_1162 (O_1162,N_27354,N_27137);
and UO_1163 (O_1163,N_26917,N_26519);
nand UO_1164 (O_1164,N_29428,N_29405);
or UO_1165 (O_1165,N_26767,N_25878);
nand UO_1166 (O_1166,N_25075,N_25533);
and UO_1167 (O_1167,N_27829,N_28329);
xor UO_1168 (O_1168,N_28264,N_26198);
and UO_1169 (O_1169,N_29671,N_26230);
nand UO_1170 (O_1170,N_26232,N_26367);
nor UO_1171 (O_1171,N_29750,N_29209);
and UO_1172 (O_1172,N_25332,N_28348);
and UO_1173 (O_1173,N_29075,N_27915);
nand UO_1174 (O_1174,N_26585,N_28932);
or UO_1175 (O_1175,N_28485,N_28081);
nor UO_1176 (O_1176,N_29553,N_26280);
and UO_1177 (O_1177,N_25633,N_27514);
and UO_1178 (O_1178,N_28403,N_28161);
nor UO_1179 (O_1179,N_27714,N_27197);
nand UO_1180 (O_1180,N_28678,N_25369);
nor UO_1181 (O_1181,N_26979,N_28999);
or UO_1182 (O_1182,N_29528,N_28322);
and UO_1183 (O_1183,N_25362,N_27933);
or UO_1184 (O_1184,N_27109,N_26354);
nor UO_1185 (O_1185,N_29724,N_25226);
and UO_1186 (O_1186,N_28957,N_29234);
or UO_1187 (O_1187,N_29606,N_27716);
nor UO_1188 (O_1188,N_28993,N_28995);
nor UO_1189 (O_1189,N_29578,N_26118);
nor UO_1190 (O_1190,N_29410,N_26817);
nand UO_1191 (O_1191,N_25157,N_29244);
nor UO_1192 (O_1192,N_26356,N_26374);
xnor UO_1193 (O_1193,N_28491,N_25379);
and UO_1194 (O_1194,N_29985,N_26346);
nand UO_1195 (O_1195,N_25422,N_28164);
nor UO_1196 (O_1196,N_27037,N_27023);
or UO_1197 (O_1197,N_26021,N_26852);
nand UO_1198 (O_1198,N_25214,N_26584);
and UO_1199 (O_1199,N_25014,N_28099);
and UO_1200 (O_1200,N_28542,N_25233);
or UO_1201 (O_1201,N_27560,N_25509);
and UO_1202 (O_1202,N_26059,N_27128);
and UO_1203 (O_1203,N_26802,N_28681);
nor UO_1204 (O_1204,N_25175,N_26860);
nand UO_1205 (O_1205,N_29841,N_27370);
nand UO_1206 (O_1206,N_26626,N_26698);
or UO_1207 (O_1207,N_28255,N_25782);
or UO_1208 (O_1208,N_25923,N_29348);
nand UO_1209 (O_1209,N_29539,N_25834);
and UO_1210 (O_1210,N_29980,N_27308);
and UO_1211 (O_1211,N_28782,N_28562);
and UO_1212 (O_1212,N_25870,N_25178);
or UO_1213 (O_1213,N_29119,N_29011);
nand UO_1214 (O_1214,N_27316,N_27835);
nor UO_1215 (O_1215,N_25596,N_29240);
nor UO_1216 (O_1216,N_29267,N_26511);
nand UO_1217 (O_1217,N_26641,N_27550);
and UO_1218 (O_1218,N_26254,N_27356);
or UO_1219 (O_1219,N_26436,N_27253);
nor UO_1220 (O_1220,N_27489,N_27971);
and UO_1221 (O_1221,N_28936,N_26736);
nand UO_1222 (O_1222,N_26023,N_29964);
and UO_1223 (O_1223,N_29824,N_27048);
or UO_1224 (O_1224,N_25467,N_28176);
or UO_1225 (O_1225,N_29050,N_27057);
nand UO_1226 (O_1226,N_26525,N_25205);
nor UO_1227 (O_1227,N_26955,N_29468);
nand UO_1228 (O_1228,N_27262,N_29537);
nor UO_1229 (O_1229,N_25513,N_27621);
and UO_1230 (O_1230,N_29774,N_28083);
and UO_1231 (O_1231,N_27433,N_27346);
or UO_1232 (O_1232,N_27759,N_28174);
nand UO_1233 (O_1233,N_26532,N_29122);
nand UO_1234 (O_1234,N_25810,N_26854);
nor UO_1235 (O_1235,N_29670,N_28481);
nor UO_1236 (O_1236,N_25795,N_29677);
or UO_1237 (O_1237,N_25794,N_28454);
or UO_1238 (O_1238,N_25938,N_29818);
nor UO_1239 (O_1239,N_28819,N_28471);
nand UO_1240 (O_1240,N_28482,N_27473);
nand UO_1241 (O_1241,N_29078,N_25084);
nor UO_1242 (O_1242,N_28560,N_27405);
nand UO_1243 (O_1243,N_29860,N_29608);
nor UO_1244 (O_1244,N_25030,N_25812);
or UO_1245 (O_1245,N_29029,N_27070);
nor UO_1246 (O_1246,N_26923,N_25912);
nand UO_1247 (O_1247,N_28477,N_26213);
or UO_1248 (O_1248,N_25854,N_29357);
nand UO_1249 (O_1249,N_25020,N_25726);
nand UO_1250 (O_1250,N_25027,N_25211);
nand UO_1251 (O_1251,N_27635,N_26985);
nor UO_1252 (O_1252,N_27849,N_25886);
nor UO_1253 (O_1253,N_25766,N_26375);
and UO_1254 (O_1254,N_25301,N_27540);
and UO_1255 (O_1255,N_26210,N_25493);
nor UO_1256 (O_1256,N_27890,N_27455);
nor UO_1257 (O_1257,N_28018,N_29398);
nor UO_1258 (O_1258,N_29219,N_26902);
and UO_1259 (O_1259,N_25013,N_27148);
and UO_1260 (O_1260,N_28706,N_26775);
or UO_1261 (O_1261,N_26691,N_26548);
and UO_1262 (O_1262,N_25161,N_26175);
nand UO_1263 (O_1263,N_25699,N_26027);
nor UO_1264 (O_1264,N_28644,N_28185);
nor UO_1265 (O_1265,N_28434,N_25430);
or UO_1266 (O_1266,N_29743,N_29693);
nor UO_1267 (O_1267,N_28652,N_26493);
nand UO_1268 (O_1268,N_26644,N_26939);
and UO_1269 (O_1269,N_26295,N_28451);
and UO_1270 (O_1270,N_25125,N_25941);
nand UO_1271 (O_1271,N_29490,N_25052);
and UO_1272 (O_1272,N_26952,N_25356);
nand UO_1273 (O_1273,N_25471,N_28855);
or UO_1274 (O_1274,N_27616,N_26004);
nand UO_1275 (O_1275,N_29754,N_28347);
nand UO_1276 (O_1276,N_29265,N_27905);
or UO_1277 (O_1277,N_25435,N_27272);
nand UO_1278 (O_1278,N_29773,N_29056);
and UO_1279 (O_1279,N_27521,N_29435);
and UO_1280 (O_1280,N_25065,N_29787);
nand UO_1281 (O_1281,N_26971,N_25571);
or UO_1282 (O_1282,N_29549,N_25429);
or UO_1283 (O_1283,N_25974,N_29665);
or UO_1284 (O_1284,N_28830,N_25313);
nor UO_1285 (O_1285,N_27799,N_28675);
or UO_1286 (O_1286,N_29948,N_27319);
and UO_1287 (O_1287,N_26063,N_28077);
nand UO_1288 (O_1288,N_25245,N_28565);
and UO_1289 (O_1289,N_26524,N_28816);
or UO_1290 (O_1290,N_29544,N_25352);
nand UO_1291 (O_1291,N_26781,N_25302);
and UO_1292 (O_1292,N_27956,N_28924);
nand UO_1293 (O_1293,N_29905,N_26451);
and UO_1294 (O_1294,N_27484,N_27784);
nor UO_1295 (O_1295,N_25434,N_25104);
nor UO_1296 (O_1296,N_27798,N_28577);
or UO_1297 (O_1297,N_28120,N_29100);
nor UO_1298 (O_1298,N_27334,N_28723);
or UO_1299 (O_1299,N_25689,N_25840);
nor UO_1300 (O_1300,N_26283,N_28686);
and UO_1301 (O_1301,N_29636,N_27523);
nand UO_1302 (O_1302,N_29425,N_27583);
and UO_1303 (O_1303,N_27690,N_25115);
and UO_1304 (O_1304,N_29322,N_27214);
or UO_1305 (O_1305,N_27282,N_26871);
and UO_1306 (O_1306,N_27639,N_25641);
nand UO_1307 (O_1307,N_26692,N_26683);
nand UO_1308 (O_1308,N_29472,N_27211);
nand UO_1309 (O_1309,N_25253,N_25830);
nand UO_1310 (O_1310,N_28421,N_27237);
nand UO_1311 (O_1311,N_26401,N_25267);
or UO_1312 (O_1312,N_26583,N_26599);
and UO_1313 (O_1313,N_28876,N_29190);
or UO_1314 (O_1314,N_27984,N_28259);
and UO_1315 (O_1315,N_28465,N_28396);
nand UO_1316 (O_1316,N_27399,N_27666);
nand UO_1317 (O_1317,N_29301,N_27430);
or UO_1318 (O_1318,N_26867,N_27341);
or UO_1319 (O_1319,N_25611,N_28302);
nand UO_1320 (O_1320,N_25606,N_25731);
or UO_1321 (O_1321,N_26269,N_25871);
and UO_1322 (O_1322,N_27772,N_25967);
or UO_1323 (O_1323,N_28996,N_29099);
and UO_1324 (O_1324,N_28351,N_28069);
and UO_1325 (O_1325,N_28979,N_28582);
and UO_1326 (O_1326,N_29849,N_28312);
or UO_1327 (O_1327,N_29210,N_25005);
nor UO_1328 (O_1328,N_27653,N_29025);
nor UO_1329 (O_1329,N_28339,N_26619);
or UO_1330 (O_1330,N_28095,N_26137);
and UO_1331 (O_1331,N_28382,N_25572);
nor UO_1332 (O_1332,N_29958,N_27131);
or UO_1333 (O_1333,N_26677,N_29114);
or UO_1334 (O_1334,N_27695,N_27644);
and UO_1335 (O_1335,N_28214,N_27445);
or UO_1336 (O_1336,N_25723,N_28309);
nor UO_1337 (O_1337,N_28543,N_25887);
nand UO_1338 (O_1338,N_29458,N_27032);
nor UO_1339 (O_1339,N_26038,N_25693);
nor UO_1340 (O_1340,N_27342,N_26396);
or UO_1341 (O_1341,N_27257,N_28813);
nand UO_1342 (O_1342,N_26877,N_27439);
nand UO_1343 (O_1343,N_25479,N_28110);
or UO_1344 (O_1344,N_29709,N_28890);
nand UO_1345 (O_1345,N_29217,N_26541);
or UO_1346 (O_1346,N_25482,N_29161);
and UO_1347 (O_1347,N_25460,N_26286);
nand UO_1348 (O_1348,N_27093,N_27384);
nor UO_1349 (O_1349,N_28296,N_29453);
and UO_1350 (O_1350,N_28354,N_29936);
or UO_1351 (O_1351,N_26516,N_27314);
nand UO_1352 (O_1352,N_25556,N_29040);
nand UO_1353 (O_1353,N_27429,N_25402);
nand UO_1354 (O_1354,N_28202,N_26444);
and UO_1355 (O_1355,N_29207,N_29776);
nand UO_1356 (O_1356,N_29353,N_26141);
nor UO_1357 (O_1357,N_29221,N_28460);
and UO_1358 (O_1358,N_29326,N_27318);
and UO_1359 (O_1359,N_25445,N_25001);
nand UO_1360 (O_1360,N_28898,N_26514);
nor UO_1361 (O_1361,N_28417,N_29042);
or UO_1362 (O_1362,N_27213,N_29308);
nor UO_1363 (O_1363,N_25548,N_27807);
nor UO_1364 (O_1364,N_27363,N_29303);
or UO_1365 (O_1365,N_29952,N_28810);
nand UO_1366 (O_1366,N_28500,N_26065);
and UO_1367 (O_1367,N_29926,N_26643);
nand UO_1368 (O_1368,N_29026,N_26120);
or UO_1369 (O_1369,N_25122,N_25943);
nor UO_1370 (O_1370,N_29325,N_28473);
or UO_1371 (O_1371,N_28345,N_29427);
or UO_1372 (O_1372,N_25730,N_26090);
nand UO_1373 (O_1373,N_28262,N_25282);
nand UO_1374 (O_1374,N_27791,N_27163);
and UO_1375 (O_1375,N_29137,N_25209);
or UO_1376 (O_1376,N_26670,N_26363);
or UO_1377 (O_1377,N_29045,N_28742);
nor UO_1378 (O_1378,N_26142,N_28639);
nor UO_1379 (O_1379,N_26612,N_29758);
or UO_1380 (O_1380,N_26410,N_28536);
nor UO_1381 (O_1381,N_28101,N_25630);
nand UO_1382 (O_1382,N_28000,N_29216);
nand UO_1383 (O_1383,N_28456,N_25190);
or UO_1384 (O_1384,N_28861,N_29939);
nand UO_1385 (O_1385,N_26252,N_25246);
and UO_1386 (O_1386,N_28650,N_25056);
or UO_1387 (O_1387,N_29212,N_29973);
and UO_1388 (O_1388,N_28420,N_29402);
nand UO_1389 (O_1389,N_28392,N_28548);
or UO_1390 (O_1390,N_28377,N_26083);
and UO_1391 (O_1391,N_29969,N_27024);
and UO_1392 (O_1392,N_28136,N_29816);
and UO_1393 (O_1393,N_29449,N_25672);
nor UO_1394 (O_1394,N_27834,N_29884);
nand UO_1395 (O_1395,N_27113,N_26391);
and UO_1396 (O_1396,N_26070,N_29316);
or UO_1397 (O_1397,N_29829,N_27783);
nand UO_1398 (O_1398,N_27302,N_25483);
or UO_1399 (O_1399,N_26085,N_29307);
and UO_1400 (O_1400,N_28702,N_26593);
and UO_1401 (O_1401,N_27534,N_25036);
nor UO_1402 (O_1402,N_27067,N_25079);
nor UO_1403 (O_1403,N_27601,N_28257);
nor UO_1404 (O_1404,N_25151,N_27817);
nand UO_1405 (O_1405,N_29037,N_25653);
nor UO_1406 (O_1406,N_29106,N_26921);
or UO_1407 (O_1407,N_28209,N_27909);
nor UO_1408 (O_1408,N_29492,N_25095);
and UO_1409 (O_1409,N_25908,N_29139);
nand UO_1410 (O_1410,N_29999,N_27917);
nand UO_1411 (O_1411,N_25173,N_29945);
and UO_1412 (O_1412,N_27204,N_25659);
nor UO_1413 (O_1413,N_27248,N_28130);
and UO_1414 (O_1414,N_27642,N_27478);
nand UO_1415 (O_1415,N_28640,N_26024);
or UO_1416 (O_1416,N_25184,N_25108);
or UO_1417 (O_1417,N_25985,N_26682);
and UO_1418 (O_1418,N_27051,N_27969);
or UO_1419 (O_1419,N_28187,N_28041);
and UO_1420 (O_1420,N_29806,N_29603);
or UO_1421 (O_1421,N_28732,N_25624);
nand UO_1422 (O_1422,N_29272,N_25559);
nor UO_1423 (O_1423,N_28806,N_25979);
nand UO_1424 (O_1424,N_28108,N_26990);
nor UO_1425 (O_1425,N_28394,N_25180);
nand UO_1426 (O_1426,N_25601,N_27228);
and UO_1427 (O_1427,N_27670,N_25966);
and UO_1428 (O_1428,N_27790,N_29536);
nor UO_1429 (O_1429,N_29882,N_27954);
and UO_1430 (O_1430,N_29865,N_25975);
or UO_1431 (O_1431,N_26742,N_28667);
xnor UO_1432 (O_1432,N_26603,N_25678);
or UO_1433 (O_1433,N_25797,N_27519);
nor UO_1434 (O_1434,N_25791,N_25279);
nor UO_1435 (O_1435,N_28092,N_26442);
nand UO_1436 (O_1436,N_26718,N_26545);
or UO_1437 (O_1437,N_28388,N_25017);
and UO_1438 (O_1438,N_25925,N_28549);
nor UO_1439 (O_1439,N_25592,N_26413);
or UO_1440 (O_1440,N_25373,N_28563);
and UO_1441 (O_1441,N_28607,N_28152);
or UO_1442 (O_1442,N_29839,N_28305);
and UO_1443 (O_1443,N_25040,N_25011);
or UO_1444 (O_1444,N_26093,N_25820);
nor UO_1445 (O_1445,N_25802,N_25514);
or UO_1446 (O_1446,N_25228,N_28235);
nor UO_1447 (O_1447,N_28527,N_26833);
and UO_1448 (O_1448,N_29250,N_28513);
xor UO_1449 (O_1449,N_26054,N_26273);
nor UO_1450 (O_1450,N_27858,N_25937);
xor UO_1451 (O_1451,N_29689,N_29607);
or UO_1452 (O_1452,N_25640,N_27571);
or UO_1453 (O_1453,N_28405,N_25826);
nor UO_1454 (O_1454,N_28218,N_29857);
or UO_1455 (O_1455,N_26069,N_29445);
or UO_1456 (O_1456,N_25991,N_27207);
nor UO_1457 (O_1457,N_27249,N_26983);
nand UO_1458 (O_1458,N_29160,N_28016);
nor UO_1459 (O_1459,N_28308,N_28768);
and UO_1460 (O_1460,N_25983,N_25166);
nor UO_1461 (O_1461,N_28923,N_29623);
and UO_1462 (O_1462,N_27520,N_29064);
nand UO_1463 (O_1463,N_26358,N_26527);
xnor UO_1464 (O_1464,N_27304,N_25297);
nand UO_1465 (O_1465,N_29339,N_28303);
or UO_1466 (O_1466,N_27594,N_26844);
nand UO_1467 (O_1467,N_27442,N_27925);
nor UO_1468 (O_1468,N_29916,N_29900);
or UO_1469 (O_1469,N_26904,N_26842);
or UO_1470 (O_1470,N_27825,N_25842);
nor UO_1471 (O_1471,N_26922,N_25444);
or UO_1472 (O_1472,N_29120,N_28183);
or UO_1473 (O_1473,N_26039,N_26572);
nand UO_1474 (O_1474,N_25063,N_25610);
nor UO_1475 (O_1475,N_28505,N_27221);
xnor UO_1476 (O_1476,N_29066,N_26651);
and UO_1477 (O_1477,N_28921,N_27035);
nand UO_1478 (O_1478,N_25382,N_29597);
or UO_1479 (O_1479,N_27813,N_26664);
or UO_1480 (O_1480,N_26557,N_27629);
xnor UO_1481 (O_1481,N_27459,N_28693);
or UO_1482 (O_1482,N_25543,N_27254);
nand UO_1483 (O_1483,N_25706,N_28762);
nand UO_1484 (O_1484,N_25150,N_29464);
or UO_1485 (O_1485,N_25087,N_29594);
nand UO_1486 (O_1486,N_28320,N_27124);
and UO_1487 (O_1487,N_29893,N_26546);
and UO_1488 (O_1488,N_26372,N_26476);
xor UO_1489 (O_1489,N_25950,N_27004);
or UO_1490 (O_1490,N_26780,N_25905);
or UO_1491 (O_1491,N_26637,N_29232);
nor UO_1492 (O_1492,N_27980,N_25860);
or UO_1493 (O_1493,N_29911,N_25487);
and UO_1494 (O_1494,N_28770,N_27414);
nand UO_1495 (O_1495,N_28638,N_25097);
nor UO_1496 (O_1496,N_26760,N_28021);
or UO_1497 (O_1497,N_28774,N_25674);
or UO_1498 (O_1498,N_29450,N_29844);
nor UO_1499 (O_1499,N_27570,N_29908);
nor UO_1500 (O_1500,N_28430,N_25895);
nand UO_1501 (O_1501,N_26344,N_25740);
nand UO_1502 (O_1502,N_28791,N_25621);
and UO_1503 (O_1503,N_25397,N_29281);
nand UO_1504 (O_1504,N_28268,N_26719);
or UO_1505 (O_1505,N_26646,N_27886);
nor UO_1506 (O_1506,N_26849,N_28614);
and UO_1507 (O_1507,N_25183,N_26164);
or UO_1508 (O_1508,N_28191,N_26379);
or UO_1509 (O_1509,N_26945,N_26969);
nand UO_1510 (O_1510,N_26528,N_27713);
nand UO_1511 (O_1511,N_26746,N_26725);
nand UO_1512 (O_1512,N_26333,N_29186);
or UO_1513 (O_1513,N_27691,N_25492);
and UO_1514 (O_1514,N_27697,N_29237);
or UO_1515 (O_1515,N_29924,N_29245);
and UO_1516 (O_1516,N_25639,N_25177);
nor UO_1517 (O_1517,N_28501,N_26768);
nor UO_1518 (O_1518,N_26160,N_28206);
nand UO_1519 (O_1519,N_27440,N_26231);
and UO_1520 (O_1520,N_25806,N_28140);
or UO_1521 (O_1521,N_25607,N_25132);
or UO_1522 (O_1522,N_29514,N_26590);
or UO_1523 (O_1523,N_26412,N_26043);
or UO_1524 (O_1524,N_25163,N_27968);
and UO_1525 (O_1525,N_29885,N_26196);
and UO_1526 (O_1526,N_29399,N_26431);
or UO_1527 (O_1527,N_27839,N_25294);
nor UO_1528 (O_1528,N_25374,N_26032);
nand UO_1529 (O_1529,N_29696,N_28217);
nand UO_1530 (O_1530,N_25099,N_28690);
and UO_1531 (O_1531,N_29289,N_28606);
nor UO_1532 (O_1532,N_28483,N_29418);
nor UO_1533 (O_1533,N_25090,N_29493);
or UO_1534 (O_1534,N_28100,N_27287);
nor UO_1535 (O_1535,N_27656,N_25902);
or UO_1536 (O_1536,N_26109,N_26654);
nand UO_1537 (O_1537,N_29319,N_28052);
or UO_1538 (O_1538,N_27598,N_29014);
nor UO_1539 (O_1539,N_25669,N_29462);
and UO_1540 (O_1540,N_26071,N_25428);
and UO_1541 (O_1541,N_26893,N_25290);
or UO_1542 (O_1542,N_27654,N_29231);
and UO_1543 (O_1543,N_27494,N_29270);
nor UO_1544 (O_1544,N_27872,N_25389);
or UO_1545 (O_1545,N_25667,N_27593);
and UO_1546 (O_1546,N_25915,N_27781);
nand UO_1547 (O_1547,N_25459,N_28635);
nand UO_1548 (O_1548,N_25739,N_26830);
nor UO_1549 (O_1549,N_28237,N_26382);
nor UO_1550 (O_1550,N_28079,N_29937);
nor UO_1551 (O_1551,N_25088,N_28945);
and UO_1552 (O_1552,N_25888,N_25227);
nor UO_1553 (O_1553,N_27501,N_28713);
or UO_1554 (O_1554,N_27482,N_25771);
nand UO_1555 (O_1555,N_25021,N_26636);
or UO_1556 (O_1556,N_29512,N_28150);
and UO_1557 (O_1557,N_25442,N_29669);
nor UO_1558 (O_1558,N_29649,N_28939);
and UO_1559 (O_1559,N_26491,N_28574);
or UO_1560 (O_1560,N_28359,N_27326);
nor UO_1561 (O_1561,N_29968,N_26684);
or UO_1562 (O_1562,N_26903,N_27592);
and UO_1563 (O_1563,N_28493,N_28907);
or UO_1564 (O_1564,N_29737,N_29931);
and UO_1565 (O_1565,N_27315,N_28699);
and UO_1566 (O_1566,N_28683,N_28707);
or UO_1567 (O_1567,N_29121,N_29226);
and UO_1568 (O_1568,N_27848,N_27402);
and UO_1569 (O_1569,N_27075,N_29519);
nor UO_1570 (O_1570,N_26510,N_29599);
and UO_1571 (O_1571,N_27929,N_27243);
nor UO_1572 (O_1572,N_28032,N_28290);
nand UO_1573 (O_1573,N_26550,N_27943);
and UO_1574 (O_1574,N_26920,N_28719);
nor UO_1575 (O_1575,N_28104,N_29434);
or UO_1576 (O_1576,N_28402,N_27353);
nand UO_1577 (O_1577,N_25411,N_26298);
nand UO_1578 (O_1578,N_25169,N_27426);
nor UO_1579 (O_1579,N_26135,N_26011);
and UO_1580 (O_1580,N_25185,N_27608);
nor UO_1581 (O_1581,N_29749,N_27141);
or UO_1582 (O_1582,N_26771,N_25114);
nor UO_1583 (O_1583,N_29866,N_29770);
nand UO_1584 (O_1584,N_25262,N_28244);
nor UO_1585 (O_1585,N_28746,N_25716);
or UO_1586 (O_1586,N_25681,N_28061);
nor UO_1587 (O_1587,N_25032,N_29089);
nand UO_1588 (O_1588,N_27417,N_26640);
and UO_1589 (O_1589,N_29668,N_28701);
and UO_1590 (O_1590,N_25324,N_29619);
and UO_1591 (O_1591,N_28912,N_26189);
and UO_1592 (O_1592,N_29886,N_27064);
nor UO_1593 (O_1593,N_25160,N_27000);
nand UO_1594 (O_1594,N_29338,N_26092);
or UO_1595 (O_1595,N_28207,N_28829);
or UO_1596 (O_1596,N_28616,N_26942);
or UO_1597 (O_1597,N_29138,N_27539);
and UO_1598 (O_1598,N_25632,N_26535);
nand UO_1599 (O_1599,N_25181,N_28438);
nand UO_1600 (O_1600,N_27558,N_29744);
nand UO_1601 (O_1601,N_26721,N_26258);
or UO_1602 (O_1602,N_28508,N_26489);
and UO_1603 (O_1603,N_26150,N_29502);
nor UO_1604 (O_1604,N_27090,N_29559);
or UO_1605 (O_1605,N_27735,N_27329);
nor UO_1606 (O_1606,N_27631,N_26712);
and UO_1607 (O_1607,N_27486,N_26560);
xnor UO_1608 (O_1608,N_25101,N_25682);
nand UO_1609 (O_1609,N_26222,N_25098);
nor UO_1610 (O_1610,N_25570,N_26553);
or UO_1611 (O_1611,N_25385,N_29071);
nor UO_1612 (O_1612,N_27882,N_26868);
nand UO_1613 (O_1613,N_28826,N_25718);
and UO_1614 (O_1614,N_25608,N_29932);
nor UO_1615 (O_1615,N_27562,N_25767);
nand UO_1616 (O_1616,N_26763,N_26897);
or UO_1617 (O_1617,N_29730,N_27588);
nand UO_1618 (O_1618,N_27657,N_26764);
nand UO_1619 (O_1619,N_25447,N_28415);
and UO_1620 (O_1620,N_26635,N_26610);
and UO_1621 (O_1621,N_28857,N_27091);
and UO_1622 (O_1622,N_25396,N_25708);
or UO_1623 (O_1623,N_29330,N_27797);
nand UO_1624 (O_1624,N_27241,N_29334);
and UO_1625 (O_1625,N_25544,N_29369);
nand UO_1626 (O_1626,N_26430,N_27801);
or UO_1627 (O_1627,N_26804,N_29652);
or UO_1628 (O_1628,N_29441,N_26659);
and UO_1629 (O_1629,N_26806,N_25963);
or UO_1630 (O_1630,N_26089,N_28870);
or UO_1631 (O_1631,N_29533,N_29306);
or UO_1632 (O_1632,N_26156,N_26029);
and UO_1633 (O_1633,N_29612,N_29072);
or UO_1634 (O_1634,N_27092,N_29504);
or UO_1635 (O_1635,N_26574,N_27026);
and UO_1636 (O_1636,N_28173,N_29957);
nand UO_1637 (O_1637,N_25401,N_28980);
and UO_1638 (O_1638,N_25787,N_25613);
nand UO_1639 (O_1639,N_29125,N_29047);
nand UO_1640 (O_1640,N_25992,N_26384);
or UO_1641 (O_1641,N_26499,N_27626);
nor UO_1642 (O_1642,N_25758,N_25910);
or UO_1643 (O_1643,N_26328,N_27022);
and UO_1644 (O_1644,N_25074,N_28793);
or UO_1645 (O_1645,N_29628,N_28363);
or UO_1646 (O_1646,N_28034,N_27056);
nor UO_1647 (O_1647,N_29728,N_25409);
or UO_1648 (O_1648,N_28243,N_25552);
nor UO_1649 (O_1649,N_28143,N_26676);
and UO_1650 (O_1650,N_27063,N_29411);
or UO_1651 (O_1651,N_27897,N_29738);
nand UO_1652 (O_1652,N_29191,N_28881);
or UO_1653 (O_1653,N_25053,N_26474);
or UO_1654 (O_1654,N_26122,N_25091);
and UO_1655 (O_1655,N_25605,N_28287);
and UO_1656 (O_1656,N_29873,N_26293);
or UO_1657 (O_1657,N_29013,N_28949);
or UO_1658 (O_1658,N_29166,N_28367);
and UO_1659 (O_1659,N_25451,N_26256);
nor UO_1660 (O_1660,N_27816,N_27771);
nand UO_1661 (O_1661,N_29997,N_28802);
and UO_1662 (O_1662,N_28226,N_29366);
nor UO_1663 (O_1663,N_29946,N_27039);
or UO_1664 (O_1664,N_28596,N_25850);
or UO_1665 (O_1665,N_25031,N_26582);
or UO_1666 (O_1666,N_27896,N_27238);
xor UO_1667 (O_1667,N_27416,N_25354);
or UO_1668 (O_1668,N_27567,N_25852);
or UO_1669 (O_1669,N_27360,N_27358);
or UO_1670 (O_1670,N_26414,N_28358);
or UO_1671 (O_1671,N_26813,N_28008);
or UO_1672 (O_1672,N_27247,N_29716);
nor UO_1673 (O_1673,N_26468,N_27428);
and UO_1674 (O_1674,N_28275,N_26290);
and UO_1675 (O_1675,N_28228,N_29994);
and UO_1676 (O_1676,N_27447,N_29767);
or UO_1677 (O_1677,N_25002,N_25283);
and UO_1678 (O_1678,N_28908,N_26727);
or UO_1679 (O_1679,N_28315,N_26679);
or UO_1680 (O_1680,N_26608,N_28267);
nand UO_1681 (O_1681,N_26184,N_25759);
nand UO_1682 (O_1682,N_27720,N_27927);
or UO_1683 (O_1683,N_27873,N_28628);
nand UO_1684 (O_1684,N_26244,N_28668);
nand UO_1685 (O_1685,N_25996,N_26862);
and UO_1686 (O_1686,N_28336,N_26437);
or UO_1687 (O_1687,N_26086,N_26741);
nand UO_1688 (O_1688,N_26789,N_26052);
or UO_1689 (O_1689,N_28604,N_25564);
and UO_1690 (O_1690,N_25317,N_25164);
nand UO_1691 (O_1691,N_26383,N_26010);
nand UO_1692 (O_1692,N_25889,N_28824);
nand UO_1693 (O_1693,N_26334,N_27239);
nor UO_1694 (O_1694,N_29546,N_28811);
nand UO_1695 (O_1695,N_28978,N_29260);
or UO_1696 (O_1696,N_28969,N_26807);
nor UO_1697 (O_1697,N_27231,N_25394);
nand UO_1698 (O_1698,N_28764,N_27153);
or UO_1699 (O_1699,N_27942,N_27191);
and UO_1700 (O_1700,N_29855,N_26631);
and UO_1701 (O_1701,N_25458,N_25377);
and UO_1702 (O_1702,N_26366,N_25779);
nand UO_1703 (O_1703,N_27536,N_28084);
nand UO_1704 (O_1704,N_26055,N_26749);
nor UO_1705 (O_1705,N_26777,N_28286);
or UO_1706 (O_1706,N_26994,N_26729);
nand UO_1707 (O_1707,N_25426,N_29976);
nor UO_1708 (O_1708,N_25498,N_25325);
nand UO_1709 (O_1709,N_29302,N_29542);
and UO_1710 (O_1710,N_27939,N_27496);
and UO_1711 (O_1711,N_29792,N_28656);
and UO_1712 (O_1712,N_26784,N_28042);
nor UO_1713 (O_1713,N_25424,N_27517);
nand UO_1714 (O_1714,N_28139,N_26194);
nand UO_1715 (O_1715,N_27078,N_26110);
and UO_1716 (O_1716,N_29113,N_25713);
nand UO_1717 (O_1717,N_26733,N_25363);
and UO_1718 (O_1718,N_28781,N_28526);
nor UO_1719 (O_1719,N_25066,N_27412);
or UO_1720 (O_1720,N_26976,N_28479);
or UO_1721 (O_1721,N_26515,N_26416);
nor UO_1722 (O_1722,N_28930,N_26678);
and UO_1723 (O_1723,N_25940,N_29215);
nand UO_1724 (O_1724,N_29967,N_29711);
nor UO_1725 (O_1725,N_27641,N_26731);
nor UO_1726 (O_1726,N_25241,N_25805);
or UO_1727 (O_1727,N_26224,N_29852);
nor UO_1728 (O_1728,N_25252,N_29719);
and UO_1729 (O_1729,N_29225,N_26026);
nor UO_1730 (O_1730,N_27467,N_27981);
nor UO_1731 (O_1731,N_26126,N_27362);
or UO_1732 (O_1732,N_26332,N_26570);
and UO_1733 (O_1733,N_27216,N_25337);
and UO_1734 (O_1734,N_29055,N_25532);
and UO_1735 (O_1735,N_27419,N_28653);
xnor UO_1736 (O_1736,N_28254,N_25701);
nand UO_1737 (O_1737,N_25372,N_25364);
nor UO_1738 (O_1738,N_25512,N_27055);
nand UO_1739 (O_1739,N_29094,N_26124);
nor UO_1740 (O_1740,N_26153,N_26878);
nand UO_1741 (O_1741,N_28165,N_27336);
nor UO_1742 (O_1742,N_27422,N_25490);
nand UO_1743 (O_1743,N_29300,N_28692);
nand UO_1744 (O_1744,N_28556,N_25081);
or UO_1745 (O_1745,N_25472,N_27305);
nand UO_1746 (O_1746,N_28404,N_25542);
nor UO_1747 (O_1747,N_27270,N_25594);
nor UO_1748 (O_1748,N_27294,N_25457);
nand UO_1749 (O_1749,N_27338,N_28236);
or UO_1750 (O_1750,N_26717,N_25351);
or UO_1751 (O_1751,N_26434,N_25531);
or UO_1752 (O_1752,N_25315,N_29775);
nor UO_1753 (O_1753,N_27488,N_28283);
xnor UO_1754 (O_1754,N_28450,N_27687);
nand UO_1755 (O_1755,N_25687,N_28967);
nor UO_1756 (O_1756,N_29904,N_27918);
nor UO_1757 (O_1757,N_25962,N_29036);
or UO_1758 (O_1758,N_25174,N_27431);
or UO_1759 (O_1759,N_26209,N_26861);
and UO_1760 (O_1760,N_26068,N_29159);
nand UO_1761 (O_1761,N_29800,N_28988);
and UO_1762 (O_1762,N_28737,N_26473);
nand UO_1763 (O_1763,N_25961,N_25345);
nor UO_1764 (O_1764,N_27754,N_28629);
or UO_1765 (O_1765,N_27561,N_26918);
or UO_1766 (O_1766,N_29269,N_28641);
or UO_1767 (O_1767,N_29833,N_26984);
or UO_1768 (O_1768,N_25425,N_28584);
nand UO_1769 (O_1769,N_29361,N_27330);
nand UO_1770 (O_1770,N_26588,N_29534);
nor UO_1771 (O_1771,N_25025,N_25874);
nand UO_1772 (O_1772,N_27297,N_26260);
nand UO_1773 (O_1773,N_28475,N_29759);
or UO_1774 (O_1774,N_28971,N_27487);
xnor UO_1775 (O_1775,N_26776,N_25855);
or UO_1776 (O_1776,N_25431,N_26544);
or UO_1777 (O_1777,N_26064,N_25454);
and UO_1778 (O_1778,N_25784,N_27973);
and UO_1779 (O_1779,N_28401,N_26130);
and UO_1780 (O_1780,N_28307,N_26188);
nand UO_1781 (O_1781,N_25171,N_26031);
or UO_1782 (O_1782,N_25469,N_29251);
and UO_1783 (O_1783,N_25230,N_29476);
or UO_1784 (O_1784,N_29656,N_25391);
and UO_1785 (O_1785,N_26308,N_28938);
or UO_1786 (O_1786,N_28676,N_27180);
nor UO_1787 (O_1787,N_26811,N_29314);
nor UO_1788 (O_1788,N_29555,N_28918);
or UO_1789 (O_1789,N_27403,N_27108);
nand UO_1790 (O_1790,N_27985,N_27347);
nand UO_1791 (O_1791,N_27705,N_25450);
nor UO_1792 (O_1792,N_28815,N_28973);
nand UO_1793 (O_1793,N_29305,N_26242);
nor UO_1794 (O_1794,N_29650,N_28049);
nor UO_1795 (O_1795,N_25970,N_27150);
nor UO_1796 (O_1796,N_28769,N_25994);
and UO_1797 (O_1797,N_27160,N_25799);
nand UO_1798 (O_1798,N_27782,N_25330);
and UO_1799 (O_1799,N_25540,N_27472);
or UO_1800 (O_1800,N_25215,N_28380);
and UO_1801 (O_1801,N_26674,N_27994);
and UO_1802 (O_1802,N_26916,N_28488);
or UO_1803 (O_1803,N_29571,N_28720);
nand UO_1804 (O_1804,N_27734,N_25959);
and UO_1805 (O_1805,N_26261,N_26330);
and UO_1806 (O_1806,N_28893,N_29077);
nor UO_1807 (O_1807,N_27284,N_28293);
nor UO_1808 (O_1808,N_26977,N_29115);
nor UO_1809 (O_1809,N_26987,N_27681);
or UO_1810 (O_1810,N_27155,N_26193);
and UO_1811 (O_1811,N_26845,N_28225);
nor UO_1812 (O_1812,N_25103,N_29152);
xor UO_1813 (O_1813,N_25600,N_28085);
nor UO_1814 (O_1814,N_28447,N_25769);
and UO_1815 (O_1815,N_28437,N_25288);
nand UO_1816 (O_1816,N_25865,N_29949);
and UO_1817 (O_1817,N_26883,N_25881);
nand UO_1818 (O_1818,N_27094,N_26229);
nor UO_1819 (O_1819,N_26865,N_26696);
nand UO_1820 (O_1820,N_29586,N_29651);
nor UO_1821 (O_1821,N_25440,N_29930);
nand UO_1822 (O_1822,N_28252,N_27617);
and UO_1823 (O_1823,N_25112,N_28470);
and UO_1824 (O_1824,N_29262,N_28297);
nor UO_1825 (O_1825,N_25804,N_25293);
or UO_1826 (O_1826,N_27998,N_26272);
and UO_1827 (O_1827,N_26325,N_28922);
and UO_1828 (O_1828,N_26035,N_27151);
nand UO_1829 (O_1829,N_26832,N_25879);
nor UO_1830 (O_1830,N_28680,N_27838);
nor UO_1831 (O_1831,N_29686,N_29883);
or UO_1832 (O_1832,N_28797,N_26559);
nand UO_1833 (O_1833,N_27721,N_28891);
and UO_1834 (O_1834,N_25832,N_26888);
nand UO_1835 (O_1835,N_28496,N_29585);
nor UO_1836 (O_1836,N_29777,N_25387);
and UO_1837 (O_1837,N_25012,N_26837);
nor UO_1838 (O_1838,N_26388,N_29333);
and UO_1839 (O_1839,N_25361,N_29734);
or UO_1840 (O_1840,N_29478,N_26669);
and UO_1841 (O_1841,N_29358,N_29801);
nand UO_1842 (O_1842,N_29082,N_26887);
or UO_1843 (O_1843,N_27935,N_28093);
and UO_1844 (O_1844,N_25987,N_27185);
or UO_1845 (O_1845,N_29614,N_25536);
nand UO_1846 (O_1846,N_29277,N_29126);
nand UO_1847 (O_1847,N_26115,N_27764);
nand UO_1848 (O_1848,N_29558,N_28620);
nand UO_1849 (O_1849,N_27792,N_27058);
nor UO_1850 (O_1850,N_25670,N_29681);
nor UO_1851 (O_1851,N_25202,N_27725);
nor UO_1852 (O_1852,N_28869,N_26856);
nand UO_1853 (O_1853,N_25698,N_28289);
or UO_1854 (O_1854,N_26066,N_26057);
nor UO_1855 (O_1855,N_25884,N_25083);
and UO_1856 (O_1856,N_29663,N_26107);
nand UO_1857 (O_1857,N_26049,N_29584);
nand UO_1858 (O_1858,N_26829,N_28190);
or UO_1859 (O_1859,N_25694,N_28511);
or UO_1860 (O_1860,N_25206,N_28060);
nor UO_1861 (O_1861,N_25080,N_27246);
nor UO_1862 (O_1862,N_26471,N_26663);
nand UO_1863 (O_1863,N_27274,N_25833);
nor UO_1864 (O_1864,N_27015,N_28134);
nor UO_1865 (O_1865,N_26848,N_27673);
or UO_1866 (O_1866,N_29798,N_25170);
nand UO_1867 (O_1867,N_27779,N_28573);
nand UO_1868 (O_1868,N_25254,N_26101);
and UO_1869 (O_1869,N_27906,N_28215);
and UO_1870 (O_1870,N_25235,N_25903);
and UO_1871 (O_1871,N_28160,N_27606);
nor UO_1872 (O_1872,N_29485,N_25462);
nor UO_1873 (O_1873,N_29108,N_26792);
or UO_1874 (O_1874,N_27566,N_28221);
or UO_1875 (O_1875,N_27452,N_28029);
nand UO_1876 (O_1876,N_27292,N_27461);
nor UO_1877 (O_1877,N_26341,N_25848);
nor UO_1878 (O_1878,N_27535,N_25793);
or UO_1879 (O_1879,N_25891,N_26882);
nor UO_1880 (O_1880,N_27502,N_25193);
and UO_1881 (O_1881,N_29110,N_25856);
or UO_1882 (O_1882,N_29443,N_26838);
or UO_1883 (O_1883,N_28364,N_26506);
or UO_1884 (O_1884,N_28258,N_26604);
or UO_1885 (O_1885,N_27952,N_28046);
and UO_1886 (O_1886,N_29407,N_26407);
nor UO_1887 (O_1887,N_26080,N_26834);
or UO_1888 (O_1888,N_29487,N_29577);
or UO_1889 (O_1889,N_26218,N_26517);
and UO_1890 (O_1890,N_26707,N_29282);
nor UO_1891 (O_1891,N_29535,N_27166);
or UO_1892 (O_1892,N_28448,N_27881);
and UO_1893 (O_1893,N_29439,N_28814);
and UO_1894 (O_1894,N_26000,N_28874);
nor UO_1895 (O_1895,N_26787,N_26726);
nor UO_1896 (O_1896,N_26450,N_27089);
nor UO_1897 (O_1897,N_28697,N_27493);
nor UO_1898 (O_1898,N_27556,N_29923);
nor UO_1899 (O_1899,N_28985,N_28094);
and UO_1900 (O_1900,N_25997,N_29545);
or UO_1901 (O_1901,N_29419,N_25789);
or UO_1902 (O_1902,N_26360,N_27668);
or UO_1903 (O_1903,N_28423,N_25776);
nand UO_1904 (O_1904,N_26512,N_27406);
and UO_1905 (O_1905,N_29384,N_26342);
nand UO_1906 (O_1906,N_25645,N_26050);
nand UO_1907 (O_1907,N_25138,N_27538);
and UO_1908 (O_1908,N_25930,N_26370);
or UO_1909 (O_1909,N_26566,N_26687);
nand UO_1910 (O_1910,N_28373,N_26758);
and UO_1911 (O_1911,N_26042,N_28240);
nor UO_1912 (O_1912,N_27123,N_28461);
or UO_1913 (O_1913,N_25481,N_28087);
nand UO_1914 (O_1914,N_28194,N_25368);
or UO_1915 (O_1915,N_26529,N_25029);
and UO_1916 (O_1916,N_26747,N_28304);
or UO_1917 (O_1917,N_29788,N_27794);
nor UO_1918 (O_1918,N_29069,N_28022);
nor UO_1919 (O_1919,N_28131,N_28181);
nor UO_1920 (O_1920,N_28288,N_28986);
or UO_1921 (O_1921,N_27409,N_25144);
nand UO_1922 (O_1922,N_26724,N_25901);
and UO_1923 (O_1923,N_25931,N_28105);
nand UO_1924 (O_1924,N_26062,N_25281);
nand UO_1925 (O_1925,N_29052,N_26088);
or UO_1926 (O_1926,N_28523,N_26183);
or UO_1927 (O_1927,N_26934,N_27388);
or UO_1928 (O_1928,N_26808,N_26826);
nand UO_1929 (O_1929,N_26180,N_27176);
and UO_1930 (O_1930,N_26909,N_29002);
or UO_1931 (O_1931,N_29717,N_28916);
and UO_1932 (O_1932,N_29452,N_25958);
nor UO_1933 (O_1933,N_25697,N_26185);
and UO_1934 (O_1934,N_27513,N_28853);
and UO_1935 (O_1935,N_26668,N_27924);
or UO_1936 (O_1936,N_28705,N_28414);
nand UO_1937 (O_1937,N_25773,N_28801);
xor UO_1938 (O_1938,N_29982,N_26046);
or UO_1939 (O_1939,N_28904,N_27407);
nor UO_1940 (O_1940,N_25845,N_25331);
nor UO_1941 (O_1941,N_26301,N_27867);
or UO_1942 (O_1942,N_26759,N_25844);
xor UO_1943 (O_1943,N_28659,N_28984);
nor UO_1944 (O_1944,N_27902,N_28356);
nand UO_1945 (O_1945,N_28232,N_26606);
or UO_1946 (O_1946,N_27624,N_26933);
or UO_1947 (O_1947,N_29779,N_28512);
xor UO_1948 (O_1948,N_25059,N_25511);
nor UO_1949 (O_1949,N_27597,N_29506);
nor UO_1950 (O_1950,N_27348,N_28383);
and UO_1951 (O_1951,N_29090,N_27017);
nand UO_1952 (O_1952,N_29850,N_27470);
nor UO_1953 (O_1953,N_29712,N_26403);
or UO_1954 (O_1954,N_29156,N_27749);
or UO_1955 (O_1955,N_26968,N_29460);
nor UO_1956 (O_1956,N_26571,N_25491);
or UO_1957 (O_1957,N_25303,N_25289);
nand UO_1958 (O_1958,N_29978,N_29766);
nand UO_1959 (O_1959,N_25707,N_26100);
and UO_1960 (O_1960,N_25266,N_28126);
or UO_1961 (O_1961,N_27490,N_25768);
nor UO_1962 (O_1962,N_26169,N_25882);
nor UO_1963 (O_1963,N_26884,N_29523);
nor UO_1964 (O_1964,N_27066,N_29675);
nor UO_1965 (O_1965,N_28119,N_26632);
or UO_1966 (O_1966,N_25525,N_27820);
and UO_1967 (O_1967,N_29507,N_28324);
nand UO_1968 (O_1968,N_26762,N_26863);
nand UO_1969 (O_1969,N_29875,N_26087);
or UO_1970 (O_1970,N_29254,N_28598);
nand UO_1971 (O_1971,N_28862,N_28271);
or UO_1972 (O_1972,N_26255,N_27408);
and UO_1973 (O_1973,N_28146,N_28569);
nand UO_1974 (O_1974,N_26690,N_28998);
nor UO_1975 (O_1975,N_25661,N_26323);
and UO_1976 (O_1976,N_26428,N_28440);
nand UO_1977 (O_1977,N_29516,N_26268);
nand UO_1978 (O_1978,N_29105,N_29214);
or UO_1979 (O_1979,N_27250,N_29350);
nand UO_1980 (O_1980,N_25843,N_28519);
or UO_1981 (O_1981,N_27828,N_28462);
or UO_1982 (O_1982,N_28594,N_27633);
or UO_1983 (O_1983,N_29556,N_26751);
or UO_1984 (O_1984,N_26030,N_28809);
nand UO_1985 (O_1985,N_25828,N_26965);
and UO_1986 (O_1986,N_26911,N_25936);
and UO_1987 (O_1987,N_29666,N_29643);
nand UO_1988 (O_1988,N_25433,N_25456);
or UO_1989 (O_1989,N_25849,N_25039);
and UO_1990 (O_1990,N_28188,N_25597);
or UO_1991 (O_1991,N_27712,N_27084);
and UO_1992 (O_1992,N_28263,N_25643);
xor UO_1993 (O_1993,N_25278,N_25839);
nand UO_1994 (O_1994,N_29925,N_27619);
nand UO_1995 (O_1995,N_29859,N_29318);
and UO_1996 (O_1996,N_26956,N_26203);
nand UO_1997 (O_1997,N_25683,N_28743);
or UO_1998 (O_1998,N_28253,N_25327);
or UO_1999 (O_1999,N_28048,N_29745);
nand UO_2000 (O_2000,N_25522,N_27809);
and UO_2001 (O_2001,N_26536,N_28865);
or UO_2002 (O_2002,N_25853,N_29922);
and UO_2003 (O_2003,N_26992,N_26538);
nand UO_2004 (O_2004,N_29782,N_29480);
nor UO_2005 (O_2005,N_26267,N_25953);
nand UO_2006 (O_2006,N_26200,N_29805);
and UO_2007 (O_2007,N_27508,N_26461);
nor UO_2008 (O_2008,N_25055,N_28132);
or UO_2009 (O_2009,N_29285,N_26881);
nor UO_2010 (O_2010,N_27961,N_27524);
nor UO_2011 (O_2011,N_26796,N_28951);
and UO_2012 (O_2012,N_26197,N_26667);
or UO_2013 (O_2013,N_29708,N_27161);
or UO_2014 (O_2014,N_25320,N_28282);
and UO_2015 (O_2015,N_27045,N_28172);
nor UO_2016 (O_2016,N_27492,N_28739);
nor UO_2017 (O_2017,N_26247,N_26338);
or UO_2018 (O_2018,N_26915,N_26547);
nor UO_2019 (O_2019,N_26642,N_29172);
nand UO_2020 (O_2020,N_28071,N_26650);
nor UO_2021 (O_2021,N_29184,N_25913);
nor UO_2022 (O_2022,N_27548,N_27267);
nor UO_2023 (O_2023,N_29581,N_28468);
and UO_2024 (O_2024,N_29382,N_29323);
and UO_2025 (O_2025,N_26456,N_25835);
nor UO_2026 (O_2026,N_26821,N_25072);
nand UO_2027 (O_2027,N_25589,N_29143);
or UO_2028 (O_2028,N_25371,N_29987);
or UO_2029 (O_2029,N_29526,N_29880);
nand UO_2030 (O_2030,N_27509,N_29474);
xnor UO_2031 (O_2031,N_25264,N_26914);
or UO_2032 (O_2032,N_27842,N_29714);
nor UO_2033 (O_2033,N_29179,N_28400);
and UO_2034 (O_2034,N_25413,N_26531);
nor UO_2035 (O_2035,N_28798,N_28294);
or UO_2036 (O_2036,N_26020,N_25196);
and UO_2037 (O_2037,N_25741,N_27218);
nand UO_2038 (O_2038,N_27761,N_25343);
and UO_2039 (O_2039,N_29633,N_29397);
nor UO_2040 (O_2040,N_25255,N_26326);
or UO_2041 (O_2041,N_29073,N_28637);
nand UO_2042 (O_2042,N_27675,N_27233);
nand UO_2043 (O_2043,N_28928,N_29256);
nand UO_2044 (O_2044,N_26314,N_28408);
nor UO_2045 (O_2045,N_27456,N_29446);
nand UO_2046 (O_2046,N_28911,N_28135);
nand UO_2047 (O_2047,N_25273,N_27717);
or UO_2048 (O_2048,N_29187,N_28103);
nand UO_2049 (O_2049,N_25263,N_25841);
nor UO_2050 (O_2050,N_26012,N_27757);
nor UO_2051 (O_2051,N_29499,N_29116);
nor UO_2052 (O_2052,N_26104,N_29154);
and UO_2053 (O_2053,N_29414,N_25617);
or UO_2054 (O_2054,N_26449,N_29170);
and UO_2055 (O_2055,N_25321,N_26913);
or UO_2056 (O_2056,N_27846,N_25123);
nand UO_2057 (O_2057,N_27110,N_28260);
nor UO_2058 (O_2058,N_29426,N_28564);
nand UO_2059 (O_2059,N_26689,N_26929);
or UO_2060 (O_2060,N_25208,N_25650);
nor UO_2061 (O_2061,N_29415,N_27982);
nand UO_2062 (O_2062,N_27133,N_27235);
nand UO_2063 (O_2063,N_29129,N_27667);
and UO_2064 (O_2064,N_29970,N_29639);
or UO_2065 (O_2065,N_28689,N_27377);
or UO_2066 (O_2066,N_25880,N_29876);
and UO_2067 (O_2067,N_26017,N_28717);
nor UO_2068 (O_2068,N_27837,N_29062);
or UO_2069 (O_2069,N_29222,N_27674);
nor UO_2070 (O_2070,N_25199,N_25353);
or UO_2071 (O_2071,N_29241,N_29074);
xnor UO_2072 (O_2072,N_26500,N_27860);
nand UO_2073 (O_2073,N_27901,N_26803);
and UO_2074 (O_2074,N_28820,N_28518);
and UO_2075 (O_2075,N_25644,N_28800);
and UO_2076 (O_2076,N_27719,N_29475);
nor UO_2077 (O_2077,N_29048,N_26587);
nand UO_2078 (O_2078,N_26357,N_29028);
nor UO_2079 (O_2079,N_25357,N_25034);
nand UO_2080 (O_2080,N_26281,N_26673);
or UO_2081 (O_2081,N_25219,N_25575);
or UO_2082 (O_2082,N_27715,N_26855);
nor UO_2083 (O_2083,N_25486,N_28284);
nor UO_2084 (O_2084,N_28839,N_29938);
and UO_2085 (O_2085,N_27945,N_28006);
nand UO_2086 (O_2086,N_27401,N_29831);
nor UO_2087 (O_2087,N_28121,N_25306);
and UO_2088 (O_2088,N_28395,N_27293);
and UO_2089 (O_2089,N_27404,N_26149);
nand UO_2090 (O_2090,N_29198,N_29531);
nor UO_2091 (O_2091,N_29430,N_26912);
or UO_2092 (O_2092,N_26103,N_26496);
or UO_2093 (O_2093,N_25545,N_27219);
or UO_2094 (O_2094,N_27678,N_28327);
nand UO_2095 (O_2095,N_27096,N_27170);
and UO_2096 (O_2096,N_25412,N_28073);
xor UO_2097 (O_2097,N_26289,N_27100);
and UO_2098 (O_2098,N_26352,N_29259);
nand UO_2099 (O_2099,N_27450,N_25113);
nand UO_2100 (O_2100,N_28790,N_26836);
nor UO_2101 (O_2101,N_26815,N_25094);
nor UO_2102 (O_2102,N_29618,N_27014);
nand UO_2103 (O_2103,N_26398,N_26819);
and UO_2104 (O_2104,N_27365,N_27158);
or UO_2105 (O_2105,N_29959,N_25077);
nor UO_2106 (O_2106,N_25566,N_28926);
or UO_2107 (O_2107,N_28091,N_29688);
nor UO_2108 (O_2108,N_25614,N_28977);
and UO_2109 (O_2109,N_26880,N_26483);
nand UO_2110 (O_2110,N_29895,N_25295);
nand UO_2111 (O_2111,N_28494,N_27471);
nor UO_2112 (O_2112,N_27507,N_25468);
or UO_2113 (O_2113,N_28883,N_27785);
nor UO_2114 (O_2114,N_26001,N_29604);
or UO_2115 (O_2115,N_25179,N_28385);
and UO_2116 (O_2116,N_29914,N_28954);
and UO_2117 (O_2117,N_28168,N_25636);
or UO_2118 (O_2118,N_27934,N_26892);
and UO_2119 (O_2119,N_26809,N_29843);
and UO_2120 (O_2120,N_29320,N_26187);
nor UO_2121 (O_2121,N_26415,N_26495);
nand UO_2122 (O_2122,N_28277,N_26970);
or UO_2123 (O_2123,N_26962,N_26139);
nand UO_2124 (O_2124,N_27062,N_25285);
nor UO_2125 (O_2125,N_28749,N_28246);
and UO_2126 (O_2126,N_25634,N_29197);
nand UO_2127 (O_2127,N_25259,N_29872);
nor UO_2128 (O_2128,N_29362,N_29863);
or UO_2129 (O_2129,N_27871,N_27892);
xor UO_2130 (O_2130,N_25590,N_25924);
or UO_2131 (O_2131,N_29995,N_27659);
and UO_2132 (O_2132,N_29565,N_29642);
and UO_2133 (O_2133,N_26946,N_28989);
and UO_2134 (O_2134,N_27552,N_27750);
nand UO_2135 (O_2135,N_28730,N_28619);
or UO_2136 (O_2136,N_27724,N_29233);
or UO_2137 (O_2137,N_27352,N_28541);
nor UO_2138 (O_2138,N_29655,N_28877);
and UO_2139 (O_2139,N_26091,N_29983);
or UO_2140 (O_2140,N_27965,N_27462);
nor UO_2141 (O_2141,N_25745,N_26486);
or UO_2142 (O_2142,N_27732,N_27187);
or UO_2143 (O_2143,N_27625,N_28427);
nand UO_2144 (O_2144,N_29810,N_28089);
nor UO_2145 (O_2145,N_28964,N_27497);
nand UO_2146 (O_2146,N_26233,N_26926);
nand UO_2147 (O_2147,N_25461,N_27252);
nand UO_2148 (O_2148,N_26378,N_25335);
or UO_2149 (O_2149,N_27224,N_26814);
nand UO_2150 (O_2150,N_28476,N_29494);
and UO_2151 (O_2151,N_25448,N_29340);
and UO_2152 (O_2152,N_29965,N_28353);
nor UO_2153 (O_2153,N_25541,N_27018);
or UO_2154 (O_2154,N_27758,N_29057);
nor UO_2155 (O_2155,N_28906,N_28449);
nor UO_2156 (O_2156,N_25737,N_25023);
and UO_2157 (O_2157,N_25831,N_28613);
or UO_2158 (O_2158,N_25554,N_26165);
nor UO_2159 (O_2159,N_27003,N_25577);
nand UO_2160 (O_2160,N_26598,N_27738);
nand UO_2161 (O_2161,N_25046,N_26181);
nor UO_2162 (O_2162,N_28330,N_29192);
nand UO_2163 (O_2163,N_25304,N_26097);
or UO_2164 (O_2164,N_29827,N_29856);
nand UO_2165 (O_2165,N_29548,N_26238);
nor UO_2166 (O_2166,N_27050,N_29647);
nand UO_2167 (O_2167,N_25742,N_27201);
and UO_2168 (O_2168,N_27953,N_25582);
nand UO_2169 (O_2169,N_27076,N_28520);
and UO_2170 (O_2170,N_29790,N_27627);
or UO_2171 (O_2171,N_28981,N_26146);
nand UO_2172 (O_2172,N_27053,N_28328);
nand UO_2173 (O_2173,N_25801,N_26399);
and UO_2174 (O_2174,N_26186,N_26744);
or UO_2175 (O_2175,N_26960,N_29495);
and UO_2176 (O_2176,N_27979,N_28398);
nor UO_2177 (O_2177,N_28269,N_28123);
nor UO_2178 (O_2178,N_28920,N_28310);
nand UO_2179 (O_2179,N_27144,N_25069);
or UO_2180 (O_2180,N_26217,N_27904);
and UO_2181 (O_2181,N_28663,N_25265);
and UO_2182 (O_2182,N_26748,N_28201);
nand UO_2183 (O_2183,N_25725,N_29808);
nor UO_2184 (O_2184,N_25466,N_29572);
nor UO_2185 (O_2185,N_25076,N_26136);
or UO_2186 (O_2186,N_26622,N_28169);
nand UO_2187 (O_2187,N_25238,N_26284);
or UO_2188 (O_2188,N_27577,N_26022);
or UO_2189 (O_2189,N_26076,N_29799);
nor UO_2190 (O_2190,N_26337,N_27787);
nor UO_2191 (O_2191,N_25453,N_29142);
and UO_2192 (O_2192,N_28763,N_29124);
nand UO_2193 (O_2193,N_27343,N_28203);
nand UO_2194 (O_2194,N_27565,N_26395);
nand UO_2195 (O_2195,N_29097,N_26597);
nor UO_2196 (O_2196,N_28431,N_25455);
and UO_2197 (O_2197,N_25414,N_28360);
nor UO_2198 (O_2198,N_27810,N_29701);
and UO_2199 (O_2199,N_29953,N_29228);
nand UO_2200 (O_2200,N_29587,N_26411);
nor UO_2201 (O_2201,N_28067,N_26753);
nor UO_2202 (O_2202,N_26408,N_29118);
or UO_2203 (O_2203,N_28063,N_27966);
and UO_2204 (O_2204,N_26058,N_29813);
or UO_2205 (O_2205,N_26048,N_27923);
or UO_2206 (O_2206,N_27223,N_26967);
and UO_2207 (O_2207,N_28786,N_26765);
and UO_2208 (O_2208,N_27198,N_25946);
nand UO_2209 (O_2209,N_27498,N_25604);
nand UO_2210 (O_2210,N_29590,N_26839);
and UO_2211 (O_2211,N_26675,N_29891);
nor UO_2212 (O_2212,N_26569,N_29312);
and UO_2213 (O_2213,N_28580,N_26991);
nand UO_2214 (O_2214,N_29067,N_26472);
nand UO_2215 (O_2215,N_28840,N_28805);
and UO_2216 (O_2216,N_27283,N_27847);
nor UO_2217 (O_2217,N_26778,N_27485);
and UO_2218 (O_2218,N_26812,N_29912);
or UO_2219 (O_2219,N_28510,N_26931);
nor UO_2220 (O_2220,N_25738,N_28864);
nor UO_2221 (O_2221,N_28622,N_28466);
nor UO_2222 (O_2222,N_26376,N_26079);
nor UO_2223 (O_2223,N_25121,N_27296);
nor UO_2224 (O_2224,N_26605,N_29812);
and UO_2225 (O_2225,N_27683,N_25026);
and UO_2226 (O_2226,N_27105,N_28521);
or UO_2227 (O_2227,N_28899,N_25524);
nor UO_2228 (O_2228,N_28195,N_27649);
and UO_2229 (O_2229,N_27420,N_29941);
nor UO_2230 (O_2230,N_29202,N_29966);
or UO_2231 (O_2231,N_27542,N_29645);
nand UO_2232 (O_2232,N_25864,N_29336);
nor UO_2233 (O_2233,N_29736,N_26937);
or UO_2234 (O_2234,N_26106,N_27726);
nand UO_2235 (O_2235,N_29807,N_29416);
and UO_2236 (O_2236,N_29432,N_29524);
nor UO_2237 (O_2237,N_29283,N_29092);
nor UO_2238 (O_2238,N_28937,N_28674);
nor UO_2239 (O_2239,N_28880,N_28045);
nor UO_2240 (O_2240,N_28780,N_29683);
nand UO_2241 (O_2241,N_28210,N_29509);
nand UO_2242 (O_2242,N_26843,N_27818);
and UO_2243 (O_2243,N_28783,N_28407);
and UO_2244 (O_2244,N_28925,N_25318);
and UO_2245 (O_2245,N_27495,N_28611);
or UO_2246 (O_2246,N_29763,N_27533);
and UO_2247 (O_2247,N_28017,N_27581);
and UO_2248 (O_2248,N_28487,N_25441);
xor UO_2249 (O_2249,N_26463,N_25642);
nor UO_2250 (O_2250,N_29134,N_29373);
nor UO_2251 (O_2251,N_28125,N_28490);
or UO_2252 (O_2252,N_25655,N_29517);
and UO_2253 (O_2253,N_27146,N_27859);
nand UO_2254 (O_2254,N_26702,N_27910);
or UO_2255 (O_2255,N_25070,N_29035);
and UO_2256 (O_2256,N_26278,N_27168);
and UO_2257 (O_2257,N_27111,N_26786);
nand UO_2258 (O_2258,N_25857,N_27371);
nand UO_2259 (O_2259,N_26422,N_29646);
xnor UO_2260 (O_2260,N_27222,N_26715);
or UO_2261 (O_2261,N_26299,N_26595);
and UO_2262 (O_2262,N_29510,N_26906);
or UO_2263 (O_2263,N_26003,N_28846);
nand UO_2264 (O_2264,N_25187,N_25973);
nor UO_2265 (O_2265,N_27770,N_26520);
nor UO_2266 (O_2266,N_27008,N_26015);
and UO_2267 (O_2267,N_25560,N_28247);
or UO_2268 (O_2268,N_27803,N_27883);
or UO_2269 (O_2269,N_27789,N_28952);
or UO_2270 (O_2270,N_27760,N_25695);
or UO_2271 (O_2271,N_28186,N_28711);
and UO_2272 (O_2272,N_28393,N_26421);
nor UO_2273 (O_2273,N_29341,N_25140);
or UO_2274 (O_2274,N_29279,N_25484);
or UO_2275 (O_2275,N_29012,N_25602);
nand UO_2276 (O_2276,N_27349,N_28065);
and UO_2277 (O_2277,N_29438,N_26098);
nand UO_2278 (O_2278,N_25477,N_29901);
and UO_2279 (O_2279,N_27767,N_27912);
nand UO_2280 (O_2280,N_27184,N_29678);
and UO_2281 (O_2281,N_28524,N_27340);
nor UO_2282 (O_2282,N_25045,N_25664);
nand UO_2283 (O_2283,N_26397,N_28633);
and UO_2284 (O_2284,N_29354,N_27052);
nor UO_2285 (O_2285,N_29104,N_27951);
nor UO_2286 (O_2286,N_25418,N_25772);
nor UO_2287 (O_2287,N_28609,N_27099);
nor UO_2288 (O_2288,N_28509,N_25807);
or UO_2289 (O_2289,N_27888,N_29144);
nand UO_2290 (O_2290,N_27242,N_28424);
nor UO_2291 (O_2291,N_27651,N_28572);
nor UO_2292 (O_2292,N_26685,N_29819);
nand UO_2293 (O_2293,N_28145,N_29266);
nand UO_2294 (O_2294,N_27002,N_28137);
or UO_2295 (O_2295,N_26950,N_25581);
and UO_2296 (O_2296,N_25096,N_26966);
and UO_2297 (O_2297,N_28224,N_27578);
nor UO_2298 (O_2298,N_26241,N_29570);
nor UO_2299 (O_2299,N_29497,N_25408);
nand UO_2300 (O_2300,N_29008,N_25700);
nand UO_2301 (O_2301,N_29579,N_29377);
or UO_2302 (O_2302,N_29220,N_29123);
or UO_2303 (O_2303,N_26498,N_29239);
or UO_2304 (O_2304,N_26462,N_26782);
nor UO_2305 (O_2305,N_27926,N_26312);
nor UO_2306 (O_2306,N_26270,N_29630);
and UO_2307 (O_2307,N_26152,N_25980);
or UO_2308 (O_2308,N_28068,N_25141);
and UO_2309 (O_2309,N_26755,N_29080);
nor UO_2310 (O_2310,N_29295,N_29551);
nand UO_2311 (O_2311,N_29732,N_27130);
and UO_2312 (O_2312,N_27680,N_28645);
nand UO_2313 (O_2313,N_25383,N_25507);
nand UO_2314 (O_2314,N_28205,N_25370);
nor UO_2315 (O_2315,N_29707,N_26941);
nand UO_2316 (O_2316,N_29188,N_29687);
or UO_2317 (O_2317,N_26158,N_25988);
or UO_2318 (O_2318,N_27395,N_29871);
and UO_2319 (O_2319,N_26355,N_28182);
nand UO_2320 (O_2320,N_27689,N_29567);
or UO_2321 (O_2321,N_29223,N_29781);
nor UO_2322 (O_2322,N_25598,N_28927);
or UO_2323 (O_2323,N_28935,N_25134);
or UO_2324 (O_2324,N_28962,N_28913);
and UO_2325 (O_2325,N_29513,N_29193);
nand UO_2326 (O_2326,N_25006,N_25527);
nor UO_2327 (O_2327,N_25316,N_26082);
or UO_2328 (O_2328,N_28112,N_26750);
xnor UO_2329 (O_2329,N_25410,N_26239);
and UO_2330 (O_2330,N_26975,N_28886);
nor UO_2331 (O_2331,N_26620,N_27345);
nor UO_2332 (O_2332,N_27679,N_29242);
nand UO_2333 (O_2333,N_29273,N_25748);
or UO_2334 (O_2334,N_25191,N_28817);
nor UO_2335 (O_2335,N_26898,N_28170);
nand UO_2336 (O_2336,N_27391,N_26953);
nand UO_2337 (O_2337,N_25251,N_29703);
and UO_2338 (O_2338,N_29038,N_25309);
xnor UO_2339 (O_2339,N_26114,N_26047);
nand UO_2340 (O_2340,N_29950,N_25342);
nand UO_2341 (O_2341,N_27868,N_28546);
nor UO_2342 (O_2342,N_25502,N_27279);
and UO_2343 (O_2343,N_28700,N_26600);
or UO_2344 (O_2344,N_27106,N_25814);
nor UO_2345 (O_2345,N_27441,N_28352);
nand UO_2346 (O_2346,N_25765,N_28612);
and UO_2347 (O_2347,N_26420,N_26816);
and UO_2348 (O_2348,N_28658,N_27120);
and UO_2349 (O_2349,N_27378,N_28621);
nand UO_2350 (O_2350,N_26484,N_25680);
and UO_2351 (O_2351,N_25813,N_27437);
or UO_2352 (O_2352,N_28340,N_26219);
or UO_2353 (O_2353,N_26497,N_26857);
or UO_2354 (O_2354,N_29424,N_26959);
nor UO_2355 (O_2355,N_27855,N_25515);
or UO_2356 (O_2356,N_29177,N_27200);
and UO_2357 (O_2357,N_29375,N_25651);
nor UO_2358 (O_2358,N_27469,N_27959);
and UO_2359 (O_2359,N_26680,N_27217);
nand UO_2360 (O_2360,N_28821,N_28677);
and UO_2361 (O_2361,N_27547,N_26365);
nor UO_2362 (O_2362,N_25755,N_25534);
or UO_2363 (O_2363,N_28357,N_25656);
nand UO_2364 (O_2364,N_27582,N_25906);
and UO_2365 (O_2365,N_29387,N_27220);
and UO_2366 (O_2366,N_28974,N_27671);
and UO_2367 (O_2367,N_27936,N_26390);
and UO_2368 (O_2368,N_28274,N_25286);
nor UO_2369 (O_2369,N_29084,N_25042);
nor UO_2370 (O_2370,N_25736,N_28245);
and UO_2371 (O_2371,N_25107,N_25735);
or UO_2372 (O_2372,N_28571,N_29175);
nand UO_2373 (O_2373,N_29085,N_29547);
and UO_2374 (O_2374,N_27987,N_27206);
or UO_2375 (O_2375,N_27427,N_29778);
or UO_2376 (O_2376,N_29826,N_25777);
nor UO_2377 (O_2377,N_29194,N_25478);
nand UO_2378 (O_2378,N_28558,N_29372);
or UO_2379 (O_2379,N_25392,N_28416);
and UO_2380 (O_2380,N_29611,N_27276);
and UO_2381 (O_2381,N_29783,N_27415);
nand UO_2382 (O_2382,N_25260,N_25668);
nor UO_2383 (O_2383,N_26951,N_29986);
nor UO_2384 (O_2384,N_28850,N_28748);
and UO_2385 (O_2385,N_25898,N_25405);
and UO_2386 (O_2386,N_26694,N_27647);
nand UO_2387 (O_2387,N_28090,N_29562);
nand UO_2388 (O_2388,N_28545,N_26034);
nand UO_2389 (O_2389,N_27079,N_26362);
nor UO_2390 (O_2390,N_28220,N_25761);
nand UO_2391 (O_2391,N_27603,N_28827);
nand UO_2392 (O_2392,N_25474,N_26182);
nand UO_2393 (O_2393,N_28608,N_25415);
nor UO_2394 (O_2394,N_29835,N_29913);
and UO_2395 (O_2395,N_26306,N_25452);
nand UO_2396 (O_2396,N_26123,N_27955);
nor UO_2397 (O_2397,N_29836,N_28655);
nand UO_2398 (O_2398,N_25877,N_29149);
nor UO_2399 (O_2399,N_26445,N_26460);
nor UO_2400 (O_2400,N_27618,N_29043);
and UO_2401 (O_2401,N_26117,N_25753);
and UO_2402 (O_2402,N_28200,N_27476);
nand UO_2403 (O_2403,N_25200,N_26769);
xnor UO_2404 (O_2404,N_29169,N_28127);
nor UO_2405 (O_2405,N_25851,N_28897);
and UO_2406 (O_2406,N_25047,N_26439);
and UO_2407 (O_2407,N_25165,N_29271);
and UO_2408 (O_2408,N_27899,N_26037);
nor UO_2409 (O_2409,N_26818,N_28831);
xnor UO_2410 (O_2410,N_25212,N_28940);
nand UO_2411 (O_2411,N_28948,N_28931);
nand UO_2412 (O_2412,N_25142,N_26761);
and UO_2413 (O_2413,N_26639,N_28983);
nand UO_2414 (O_2414,N_28445,N_26084);
and UO_2415 (O_2415,N_25153,N_25926);
nand UO_2416 (O_2416,N_29654,N_29768);
or UO_2417 (O_2417,N_26371,N_26997);
and UO_2418 (O_2418,N_27804,N_25420);
nand UO_2419 (O_2419,N_27273,N_28504);
nor UO_2420 (O_2420,N_25890,N_29034);
nor UO_2421 (O_2421,N_27866,N_27992);
nor UO_2422 (O_2422,N_26757,N_26288);
nor UO_2423 (O_2423,N_28776,N_28381);
or UO_2424 (O_2424,N_27515,N_29919);
nand UO_2425 (O_2425,N_27722,N_26368);
or UO_2426 (O_2426,N_28704,N_29780);
or UO_2427 (O_2427,N_25827,N_27989);
or UO_2428 (O_2428,N_25136,N_27042);
or UO_2429 (O_2429,N_29180,N_29422);
and UO_2430 (O_2430,N_29496,N_29706);
and UO_2431 (O_2431,N_25155,N_27753);
or UO_2432 (O_2432,N_29388,N_27913);
nand UO_2433 (O_2433,N_25421,N_26810);
nor UO_2434 (O_2434,N_29457,N_28057);
or UO_2435 (O_2435,N_29610,N_27277);
nand UO_2436 (O_2436,N_28788,N_27740);
or UO_2437 (O_2437,N_25663,N_26831);
nand UO_2438 (O_2438,N_29401,N_26901);
nor UO_2439 (O_2439,N_28378,N_27013);
nand UO_2440 (O_2440,N_27664,N_26948);
nand UO_2441 (O_2441,N_28001,N_25568);
or UO_2442 (O_2442,N_25728,N_29181);
or UO_2443 (O_2443,N_26327,N_25139);
or UO_2444 (O_2444,N_27800,N_26896);
xnor UO_2445 (O_2445,N_26879,N_25131);
nor UO_2446 (O_2446,N_29751,N_29153);
nand UO_2447 (O_2447,N_26591,N_27707);
nor UO_2448 (O_2448,N_29235,N_27622);
nand UO_2449 (O_2449,N_26377,N_27361);
nor UO_2450 (O_2450,N_27443,N_26711);
or UO_2451 (O_2451,N_27311,N_28439);
or UO_2452 (O_2452,N_27704,N_25637);
and UO_2453 (O_2453,N_28499,N_26264);
and UO_2454 (O_2454,N_28767,N_26899);
nand UO_2455 (O_2455,N_27663,N_26452);
and UO_2456 (O_2456,N_25770,N_25310);
or UO_2457 (O_2457,N_28097,N_28688);
nand UO_2458 (O_2458,N_29915,N_29406);
nand UO_2459 (O_2459,N_25406,N_29091);
and UO_2460 (O_2460,N_27240,N_29437);
nand UO_2461 (O_2461,N_27572,N_26207);
or UO_2462 (O_2462,N_25223,N_25666);
or UO_2463 (O_2463,N_28872,N_28390);
xnor UO_2464 (O_2464,N_28076,N_25800);
and UO_2465 (O_2465,N_29680,N_25892);
nor UO_2466 (O_2466,N_25237,N_29345);
nand UO_2467 (O_2467,N_25922,N_26173);
nor UO_2468 (O_2468,N_27589,N_25018);
and UO_2469 (O_2469,N_26688,N_29163);
or UO_2470 (O_2470,N_25438,N_27736);
or UO_2471 (O_2471,N_28882,N_28480);
and UO_2472 (O_2472,N_28773,N_28055);
nand UO_2473 (O_2473,N_27380,N_28735);
nand UO_2474 (O_2474,N_27286,N_26756);
and UO_2475 (O_2475,N_27491,N_29702);
nor UO_2476 (O_2476,N_29569,N_29848);
nor UO_2477 (O_2477,N_28332,N_26944);
or UO_2478 (O_2478,N_27827,N_27157);
nor UO_2479 (O_2479,N_27322,N_29141);
nand UO_2480 (O_2480,N_29391,N_27119);
nor UO_2481 (O_2481,N_27700,N_28410);
nand UO_2482 (O_2482,N_27229,N_28054);
or UO_2483 (O_2483,N_27364,N_28138);
nand UO_2484 (O_2484,N_25360,N_29990);
nand UO_2485 (O_2485,N_29409,N_27466);
nor UO_2486 (O_2486,N_28722,N_28858);
nand UO_2487 (O_2487,N_25774,N_25120);
or UO_2488 (O_2488,N_26248,N_28015);
or UO_2489 (O_2489,N_28027,N_28064);
and UO_2490 (O_2490,N_28744,N_27852);
or UO_2491 (O_2491,N_27309,N_27139);
nand UO_2492 (O_2492,N_28375,N_26045);
or UO_2493 (O_2493,N_29471,N_26095);
or UO_2494 (O_2494,N_25195,N_29518);
and UO_2495 (O_2495,N_26303,N_25715);
and UO_2496 (O_2496,N_26745,N_26647);
nor UO_2497 (O_2497,N_26159,N_25322);
or UO_2498 (O_2498,N_25204,N_29858);
and UO_2499 (O_2499,N_28627,N_26543);
nand UO_2500 (O_2500,N_26029,N_29375);
nand UO_2501 (O_2501,N_27296,N_26347);
nor UO_2502 (O_2502,N_27476,N_25469);
nand UO_2503 (O_2503,N_28792,N_28506);
and UO_2504 (O_2504,N_29649,N_29755);
or UO_2505 (O_2505,N_25562,N_25020);
nor UO_2506 (O_2506,N_28335,N_28448);
or UO_2507 (O_2507,N_27179,N_29581);
or UO_2508 (O_2508,N_29308,N_28734);
nor UO_2509 (O_2509,N_25854,N_26823);
and UO_2510 (O_2510,N_29207,N_28379);
nor UO_2511 (O_2511,N_25523,N_29867);
and UO_2512 (O_2512,N_28811,N_27476);
or UO_2513 (O_2513,N_29872,N_29040);
and UO_2514 (O_2514,N_25299,N_25987);
nor UO_2515 (O_2515,N_26214,N_28276);
and UO_2516 (O_2516,N_25390,N_27400);
or UO_2517 (O_2517,N_29717,N_27493);
nor UO_2518 (O_2518,N_26410,N_28462);
nor UO_2519 (O_2519,N_28581,N_25914);
or UO_2520 (O_2520,N_26060,N_27099);
or UO_2521 (O_2521,N_25063,N_26236);
nand UO_2522 (O_2522,N_28254,N_29999);
and UO_2523 (O_2523,N_27774,N_29089);
nand UO_2524 (O_2524,N_27758,N_25942);
and UO_2525 (O_2525,N_25270,N_26694);
nor UO_2526 (O_2526,N_26528,N_29861);
nor UO_2527 (O_2527,N_25901,N_25383);
nand UO_2528 (O_2528,N_27342,N_29011);
or UO_2529 (O_2529,N_27335,N_26931);
and UO_2530 (O_2530,N_26689,N_28243);
and UO_2531 (O_2531,N_26831,N_26022);
and UO_2532 (O_2532,N_25890,N_28074);
or UO_2533 (O_2533,N_27591,N_28662);
nor UO_2534 (O_2534,N_27752,N_29262);
or UO_2535 (O_2535,N_28000,N_28475);
nor UO_2536 (O_2536,N_25899,N_28768);
and UO_2537 (O_2537,N_28243,N_26331);
or UO_2538 (O_2538,N_26447,N_27116);
or UO_2539 (O_2539,N_28392,N_26669);
nand UO_2540 (O_2540,N_29494,N_29054);
nor UO_2541 (O_2541,N_25290,N_27239);
nand UO_2542 (O_2542,N_26117,N_27804);
nor UO_2543 (O_2543,N_29773,N_26271);
and UO_2544 (O_2544,N_26839,N_28455);
nand UO_2545 (O_2545,N_25821,N_29100);
nand UO_2546 (O_2546,N_29632,N_28006);
and UO_2547 (O_2547,N_29403,N_29874);
or UO_2548 (O_2548,N_27434,N_27779);
nand UO_2549 (O_2549,N_29519,N_27813);
or UO_2550 (O_2550,N_29188,N_29988);
and UO_2551 (O_2551,N_27909,N_25302);
or UO_2552 (O_2552,N_27658,N_25386);
nor UO_2553 (O_2553,N_29586,N_29640);
or UO_2554 (O_2554,N_26351,N_27117);
nor UO_2555 (O_2555,N_25361,N_26889);
and UO_2556 (O_2556,N_26063,N_29488);
or UO_2557 (O_2557,N_28326,N_27638);
nor UO_2558 (O_2558,N_25377,N_26260);
or UO_2559 (O_2559,N_26477,N_26870);
or UO_2560 (O_2560,N_25695,N_29568);
nand UO_2561 (O_2561,N_26179,N_28178);
nand UO_2562 (O_2562,N_28068,N_27630);
or UO_2563 (O_2563,N_28139,N_29619);
nor UO_2564 (O_2564,N_25730,N_29025);
and UO_2565 (O_2565,N_29101,N_26641);
nor UO_2566 (O_2566,N_29377,N_28023);
and UO_2567 (O_2567,N_27945,N_27355);
and UO_2568 (O_2568,N_27900,N_28031);
or UO_2569 (O_2569,N_27006,N_25469);
nor UO_2570 (O_2570,N_29606,N_28980);
or UO_2571 (O_2571,N_29186,N_29980);
and UO_2572 (O_2572,N_27322,N_27512);
or UO_2573 (O_2573,N_28611,N_26882);
or UO_2574 (O_2574,N_29380,N_25812);
nor UO_2575 (O_2575,N_26048,N_27545);
nand UO_2576 (O_2576,N_27163,N_27778);
nor UO_2577 (O_2577,N_28654,N_26698);
or UO_2578 (O_2578,N_29153,N_27880);
nor UO_2579 (O_2579,N_28264,N_28045);
or UO_2580 (O_2580,N_25583,N_25567);
and UO_2581 (O_2581,N_27706,N_28225);
or UO_2582 (O_2582,N_28213,N_26666);
nand UO_2583 (O_2583,N_27468,N_28789);
nand UO_2584 (O_2584,N_26363,N_25403);
nand UO_2585 (O_2585,N_29373,N_26855);
and UO_2586 (O_2586,N_27067,N_27473);
nor UO_2587 (O_2587,N_27469,N_26105);
nand UO_2588 (O_2588,N_27814,N_29489);
nor UO_2589 (O_2589,N_28162,N_27603);
or UO_2590 (O_2590,N_28570,N_26398);
nand UO_2591 (O_2591,N_26252,N_29459);
and UO_2592 (O_2592,N_26638,N_27522);
nor UO_2593 (O_2593,N_29106,N_26004);
and UO_2594 (O_2594,N_26261,N_27923);
or UO_2595 (O_2595,N_29733,N_28639);
or UO_2596 (O_2596,N_27638,N_28962);
or UO_2597 (O_2597,N_28588,N_27872);
and UO_2598 (O_2598,N_29855,N_27619);
and UO_2599 (O_2599,N_28087,N_26338);
and UO_2600 (O_2600,N_29235,N_25595);
xnor UO_2601 (O_2601,N_25880,N_27912);
nor UO_2602 (O_2602,N_28216,N_29782);
nand UO_2603 (O_2603,N_26612,N_27642);
or UO_2604 (O_2604,N_25322,N_27923);
or UO_2605 (O_2605,N_28855,N_26297);
and UO_2606 (O_2606,N_27084,N_29061);
or UO_2607 (O_2607,N_26434,N_28968);
or UO_2608 (O_2608,N_26672,N_27852);
and UO_2609 (O_2609,N_28936,N_29622);
or UO_2610 (O_2610,N_28868,N_29507);
nor UO_2611 (O_2611,N_27580,N_27393);
or UO_2612 (O_2612,N_26210,N_29060);
and UO_2613 (O_2613,N_28442,N_27098);
nor UO_2614 (O_2614,N_29055,N_25521);
and UO_2615 (O_2615,N_28474,N_25691);
or UO_2616 (O_2616,N_29696,N_27986);
and UO_2617 (O_2617,N_29899,N_27542);
or UO_2618 (O_2618,N_28718,N_26858);
nand UO_2619 (O_2619,N_28781,N_25935);
or UO_2620 (O_2620,N_26181,N_29493);
nand UO_2621 (O_2621,N_27379,N_29562);
nand UO_2622 (O_2622,N_25047,N_26601);
nor UO_2623 (O_2623,N_25371,N_28878);
nand UO_2624 (O_2624,N_27474,N_27560);
nor UO_2625 (O_2625,N_26174,N_28672);
nand UO_2626 (O_2626,N_26209,N_26596);
nor UO_2627 (O_2627,N_29728,N_29639);
nand UO_2628 (O_2628,N_29291,N_28849);
nor UO_2629 (O_2629,N_27602,N_26876);
and UO_2630 (O_2630,N_26241,N_26337);
or UO_2631 (O_2631,N_27302,N_25676);
nor UO_2632 (O_2632,N_29195,N_25878);
or UO_2633 (O_2633,N_25429,N_28412);
nor UO_2634 (O_2634,N_27400,N_29149);
or UO_2635 (O_2635,N_26727,N_25807);
nor UO_2636 (O_2636,N_25996,N_27690);
xor UO_2637 (O_2637,N_29461,N_28599);
or UO_2638 (O_2638,N_25070,N_26455);
and UO_2639 (O_2639,N_29744,N_28180);
nor UO_2640 (O_2640,N_28138,N_28876);
nand UO_2641 (O_2641,N_25780,N_25673);
and UO_2642 (O_2642,N_27416,N_25140);
nand UO_2643 (O_2643,N_26982,N_29233);
nor UO_2644 (O_2644,N_26546,N_27826);
and UO_2645 (O_2645,N_28015,N_27332);
or UO_2646 (O_2646,N_28785,N_28498);
or UO_2647 (O_2647,N_25156,N_28109);
or UO_2648 (O_2648,N_29396,N_25334);
and UO_2649 (O_2649,N_27213,N_25463);
and UO_2650 (O_2650,N_28410,N_25727);
nor UO_2651 (O_2651,N_29936,N_25031);
and UO_2652 (O_2652,N_27080,N_26571);
nand UO_2653 (O_2653,N_28506,N_26143);
and UO_2654 (O_2654,N_27107,N_26610);
nor UO_2655 (O_2655,N_27842,N_25436);
and UO_2656 (O_2656,N_29110,N_27854);
and UO_2657 (O_2657,N_28289,N_28055);
or UO_2658 (O_2658,N_29454,N_28092);
or UO_2659 (O_2659,N_25212,N_29289);
nand UO_2660 (O_2660,N_25749,N_26184);
and UO_2661 (O_2661,N_25897,N_26517);
and UO_2662 (O_2662,N_28194,N_26937);
nor UO_2663 (O_2663,N_25396,N_26641);
and UO_2664 (O_2664,N_26244,N_26370);
and UO_2665 (O_2665,N_25431,N_29871);
or UO_2666 (O_2666,N_25133,N_29756);
nand UO_2667 (O_2667,N_28758,N_27637);
nor UO_2668 (O_2668,N_26673,N_27389);
nand UO_2669 (O_2669,N_28589,N_27265);
or UO_2670 (O_2670,N_27713,N_26269);
or UO_2671 (O_2671,N_25989,N_29179);
nand UO_2672 (O_2672,N_29866,N_26562);
nor UO_2673 (O_2673,N_26369,N_26699);
or UO_2674 (O_2674,N_27662,N_27220);
or UO_2675 (O_2675,N_26829,N_26532);
or UO_2676 (O_2676,N_25167,N_28779);
nor UO_2677 (O_2677,N_27025,N_29212);
or UO_2678 (O_2678,N_26874,N_25213);
or UO_2679 (O_2679,N_25405,N_26628);
nand UO_2680 (O_2680,N_27892,N_29235);
nor UO_2681 (O_2681,N_26918,N_29849);
and UO_2682 (O_2682,N_29253,N_27217);
or UO_2683 (O_2683,N_28674,N_29543);
and UO_2684 (O_2684,N_27729,N_25646);
nor UO_2685 (O_2685,N_26564,N_27803);
or UO_2686 (O_2686,N_25771,N_27786);
and UO_2687 (O_2687,N_27447,N_27162);
and UO_2688 (O_2688,N_26751,N_27389);
nand UO_2689 (O_2689,N_26511,N_29907);
nor UO_2690 (O_2690,N_29301,N_25210);
nand UO_2691 (O_2691,N_29046,N_29717);
nor UO_2692 (O_2692,N_25658,N_27043);
or UO_2693 (O_2693,N_28295,N_29758);
and UO_2694 (O_2694,N_28856,N_28711);
nand UO_2695 (O_2695,N_28080,N_28571);
or UO_2696 (O_2696,N_26720,N_26901);
nand UO_2697 (O_2697,N_27456,N_29773);
nand UO_2698 (O_2698,N_25801,N_29882);
and UO_2699 (O_2699,N_25953,N_27749);
and UO_2700 (O_2700,N_29897,N_25174);
or UO_2701 (O_2701,N_26440,N_29636);
xnor UO_2702 (O_2702,N_27609,N_29332);
nand UO_2703 (O_2703,N_29959,N_28420);
or UO_2704 (O_2704,N_29256,N_25392);
nand UO_2705 (O_2705,N_26906,N_28296);
and UO_2706 (O_2706,N_27390,N_25503);
and UO_2707 (O_2707,N_29712,N_28115);
and UO_2708 (O_2708,N_28164,N_28081);
nand UO_2709 (O_2709,N_29250,N_27412);
nand UO_2710 (O_2710,N_28683,N_27395);
and UO_2711 (O_2711,N_26334,N_26964);
and UO_2712 (O_2712,N_27212,N_25466);
nand UO_2713 (O_2713,N_29140,N_29739);
and UO_2714 (O_2714,N_26289,N_26739);
or UO_2715 (O_2715,N_29451,N_27381);
nor UO_2716 (O_2716,N_29040,N_27118);
nand UO_2717 (O_2717,N_29194,N_27331);
nand UO_2718 (O_2718,N_29346,N_29009);
nand UO_2719 (O_2719,N_28777,N_25175);
nand UO_2720 (O_2720,N_28335,N_25371);
nand UO_2721 (O_2721,N_25202,N_28517);
or UO_2722 (O_2722,N_27560,N_29030);
nand UO_2723 (O_2723,N_25138,N_27477);
and UO_2724 (O_2724,N_25624,N_28427);
or UO_2725 (O_2725,N_28381,N_28774);
and UO_2726 (O_2726,N_26991,N_26003);
nand UO_2727 (O_2727,N_28628,N_25301);
or UO_2728 (O_2728,N_28016,N_25965);
nand UO_2729 (O_2729,N_25376,N_29136);
nor UO_2730 (O_2730,N_29249,N_26471);
nor UO_2731 (O_2731,N_29383,N_27157);
and UO_2732 (O_2732,N_29867,N_28397);
or UO_2733 (O_2733,N_26704,N_26480);
nand UO_2734 (O_2734,N_28987,N_25348);
or UO_2735 (O_2735,N_26242,N_28970);
xnor UO_2736 (O_2736,N_25375,N_28999);
nor UO_2737 (O_2737,N_25655,N_28243);
and UO_2738 (O_2738,N_29073,N_27932);
nand UO_2739 (O_2739,N_27839,N_29961);
or UO_2740 (O_2740,N_27257,N_29415);
nand UO_2741 (O_2741,N_26851,N_29316);
nand UO_2742 (O_2742,N_25512,N_25283);
nor UO_2743 (O_2743,N_28545,N_25293);
nand UO_2744 (O_2744,N_27983,N_29141);
and UO_2745 (O_2745,N_29732,N_28303);
or UO_2746 (O_2746,N_29735,N_26834);
nor UO_2747 (O_2747,N_25924,N_26071);
nor UO_2748 (O_2748,N_29592,N_29560);
and UO_2749 (O_2749,N_25527,N_25368);
and UO_2750 (O_2750,N_29235,N_27088);
and UO_2751 (O_2751,N_29124,N_29424);
or UO_2752 (O_2752,N_29410,N_26938);
nand UO_2753 (O_2753,N_27071,N_29873);
nor UO_2754 (O_2754,N_29435,N_25033);
nand UO_2755 (O_2755,N_27219,N_27707);
or UO_2756 (O_2756,N_28143,N_28800);
nand UO_2757 (O_2757,N_29283,N_28791);
nor UO_2758 (O_2758,N_25017,N_26317);
and UO_2759 (O_2759,N_27801,N_27949);
nor UO_2760 (O_2760,N_27339,N_25737);
nand UO_2761 (O_2761,N_25359,N_28151);
nand UO_2762 (O_2762,N_25538,N_27445);
nand UO_2763 (O_2763,N_29734,N_25648);
nand UO_2764 (O_2764,N_28233,N_29502);
and UO_2765 (O_2765,N_29705,N_25751);
nor UO_2766 (O_2766,N_26385,N_27807);
nor UO_2767 (O_2767,N_29303,N_25925);
nand UO_2768 (O_2768,N_26079,N_27855);
and UO_2769 (O_2769,N_25219,N_29628);
nor UO_2770 (O_2770,N_28418,N_27989);
and UO_2771 (O_2771,N_28852,N_29415);
and UO_2772 (O_2772,N_29232,N_28142);
nor UO_2773 (O_2773,N_26761,N_29813);
nand UO_2774 (O_2774,N_25793,N_25317);
or UO_2775 (O_2775,N_26919,N_26265);
nand UO_2776 (O_2776,N_27273,N_26448);
or UO_2777 (O_2777,N_28741,N_26973);
or UO_2778 (O_2778,N_27956,N_27079);
or UO_2779 (O_2779,N_29535,N_25760);
nor UO_2780 (O_2780,N_29454,N_25076);
nor UO_2781 (O_2781,N_27364,N_25014);
nand UO_2782 (O_2782,N_26434,N_27057);
nor UO_2783 (O_2783,N_29220,N_27874);
and UO_2784 (O_2784,N_27282,N_27093);
or UO_2785 (O_2785,N_25361,N_27469);
nor UO_2786 (O_2786,N_28051,N_27252);
nand UO_2787 (O_2787,N_25167,N_25865);
or UO_2788 (O_2788,N_27212,N_25626);
nor UO_2789 (O_2789,N_27125,N_29761);
and UO_2790 (O_2790,N_28441,N_25311);
nor UO_2791 (O_2791,N_26318,N_28637);
nor UO_2792 (O_2792,N_25296,N_28965);
and UO_2793 (O_2793,N_26663,N_25181);
or UO_2794 (O_2794,N_28852,N_27643);
and UO_2795 (O_2795,N_28600,N_27890);
and UO_2796 (O_2796,N_28839,N_25824);
or UO_2797 (O_2797,N_29700,N_27832);
and UO_2798 (O_2798,N_29844,N_29526);
and UO_2799 (O_2799,N_27839,N_28202);
and UO_2800 (O_2800,N_29984,N_26530);
nand UO_2801 (O_2801,N_28972,N_25676);
or UO_2802 (O_2802,N_29404,N_29958);
or UO_2803 (O_2803,N_29186,N_28939);
nand UO_2804 (O_2804,N_27893,N_29942);
or UO_2805 (O_2805,N_28767,N_26163);
and UO_2806 (O_2806,N_28639,N_25723);
nor UO_2807 (O_2807,N_25207,N_26562);
and UO_2808 (O_2808,N_28654,N_25247);
xnor UO_2809 (O_2809,N_25600,N_28584);
and UO_2810 (O_2810,N_26930,N_27877);
nor UO_2811 (O_2811,N_28681,N_29933);
nor UO_2812 (O_2812,N_25845,N_26318);
nor UO_2813 (O_2813,N_25151,N_26035);
nand UO_2814 (O_2814,N_27678,N_29185);
nand UO_2815 (O_2815,N_28839,N_26188);
nand UO_2816 (O_2816,N_28763,N_27616);
nor UO_2817 (O_2817,N_26827,N_25400);
or UO_2818 (O_2818,N_25507,N_27547);
nor UO_2819 (O_2819,N_27059,N_27209);
nor UO_2820 (O_2820,N_25154,N_25918);
and UO_2821 (O_2821,N_25108,N_26179);
or UO_2822 (O_2822,N_26612,N_25502);
or UO_2823 (O_2823,N_26874,N_29140);
nor UO_2824 (O_2824,N_25139,N_28054);
nand UO_2825 (O_2825,N_28972,N_29397);
or UO_2826 (O_2826,N_29919,N_26526);
nor UO_2827 (O_2827,N_29074,N_28885);
nor UO_2828 (O_2828,N_27999,N_25298);
nor UO_2829 (O_2829,N_29179,N_28011);
nor UO_2830 (O_2830,N_28088,N_28653);
and UO_2831 (O_2831,N_28243,N_28574);
nor UO_2832 (O_2832,N_29771,N_26222);
and UO_2833 (O_2833,N_25029,N_26888);
nand UO_2834 (O_2834,N_27831,N_28029);
or UO_2835 (O_2835,N_26307,N_28616);
or UO_2836 (O_2836,N_27700,N_29268);
and UO_2837 (O_2837,N_29928,N_29240);
or UO_2838 (O_2838,N_27039,N_26611);
nand UO_2839 (O_2839,N_26368,N_29233);
nand UO_2840 (O_2840,N_29283,N_26142);
xor UO_2841 (O_2841,N_28100,N_27525);
xor UO_2842 (O_2842,N_25404,N_26522);
nor UO_2843 (O_2843,N_29290,N_25723);
and UO_2844 (O_2844,N_25017,N_25596);
nand UO_2845 (O_2845,N_27783,N_28574);
and UO_2846 (O_2846,N_25738,N_28627);
and UO_2847 (O_2847,N_29891,N_25424);
nand UO_2848 (O_2848,N_27848,N_27941);
nand UO_2849 (O_2849,N_26407,N_26263);
and UO_2850 (O_2850,N_26847,N_28184);
nor UO_2851 (O_2851,N_29709,N_25520);
nor UO_2852 (O_2852,N_27238,N_29090);
nor UO_2853 (O_2853,N_25216,N_26146);
and UO_2854 (O_2854,N_27549,N_26584);
and UO_2855 (O_2855,N_29350,N_29271);
or UO_2856 (O_2856,N_27658,N_25223);
nand UO_2857 (O_2857,N_29532,N_28737);
or UO_2858 (O_2858,N_25120,N_27805);
or UO_2859 (O_2859,N_26190,N_29894);
nor UO_2860 (O_2860,N_27317,N_28111);
and UO_2861 (O_2861,N_25482,N_26290);
nor UO_2862 (O_2862,N_25313,N_27398);
or UO_2863 (O_2863,N_25501,N_25584);
nor UO_2864 (O_2864,N_26598,N_28727);
nor UO_2865 (O_2865,N_26075,N_29286);
or UO_2866 (O_2866,N_26084,N_25281);
or UO_2867 (O_2867,N_27065,N_27663);
nand UO_2868 (O_2868,N_26296,N_28810);
and UO_2869 (O_2869,N_29308,N_27090);
nor UO_2870 (O_2870,N_27856,N_29254);
nand UO_2871 (O_2871,N_27933,N_29886);
nor UO_2872 (O_2872,N_27087,N_26176);
nor UO_2873 (O_2873,N_29723,N_27546);
nand UO_2874 (O_2874,N_26683,N_26634);
and UO_2875 (O_2875,N_29507,N_26947);
or UO_2876 (O_2876,N_25045,N_25876);
or UO_2877 (O_2877,N_28126,N_29626);
and UO_2878 (O_2878,N_27438,N_29552);
or UO_2879 (O_2879,N_26306,N_26382);
nand UO_2880 (O_2880,N_28483,N_28748);
nand UO_2881 (O_2881,N_29228,N_28281);
nor UO_2882 (O_2882,N_25535,N_26900);
and UO_2883 (O_2883,N_25944,N_27508);
and UO_2884 (O_2884,N_29568,N_26792);
xor UO_2885 (O_2885,N_29944,N_25050);
nand UO_2886 (O_2886,N_29164,N_25047);
and UO_2887 (O_2887,N_25125,N_27078);
or UO_2888 (O_2888,N_25162,N_28435);
nand UO_2889 (O_2889,N_28213,N_29077);
or UO_2890 (O_2890,N_29781,N_28577);
nor UO_2891 (O_2891,N_26319,N_29648);
nand UO_2892 (O_2892,N_26970,N_26861);
nand UO_2893 (O_2893,N_29504,N_29773);
nor UO_2894 (O_2894,N_26590,N_27457);
or UO_2895 (O_2895,N_26928,N_25654);
nor UO_2896 (O_2896,N_29569,N_26670);
and UO_2897 (O_2897,N_26304,N_28862);
or UO_2898 (O_2898,N_26634,N_26032);
nand UO_2899 (O_2899,N_26667,N_25324);
nand UO_2900 (O_2900,N_26722,N_26692);
nor UO_2901 (O_2901,N_26883,N_26784);
or UO_2902 (O_2902,N_27490,N_25783);
and UO_2903 (O_2903,N_28126,N_26542);
and UO_2904 (O_2904,N_28036,N_29094);
nand UO_2905 (O_2905,N_26690,N_25932);
or UO_2906 (O_2906,N_27294,N_26482);
or UO_2907 (O_2907,N_25120,N_27423);
and UO_2908 (O_2908,N_29779,N_26177);
nor UO_2909 (O_2909,N_29964,N_27647);
nand UO_2910 (O_2910,N_27418,N_26291);
nand UO_2911 (O_2911,N_25819,N_25658);
or UO_2912 (O_2912,N_28236,N_26275);
or UO_2913 (O_2913,N_27151,N_28456);
nand UO_2914 (O_2914,N_27875,N_26833);
nand UO_2915 (O_2915,N_28310,N_27915);
or UO_2916 (O_2916,N_28654,N_29243);
nor UO_2917 (O_2917,N_28191,N_27223);
and UO_2918 (O_2918,N_28771,N_27232);
and UO_2919 (O_2919,N_27014,N_26592);
or UO_2920 (O_2920,N_29640,N_25071);
nor UO_2921 (O_2921,N_29084,N_25989);
nand UO_2922 (O_2922,N_28956,N_27728);
and UO_2923 (O_2923,N_29932,N_26661);
and UO_2924 (O_2924,N_25033,N_25134);
or UO_2925 (O_2925,N_26797,N_25166);
or UO_2926 (O_2926,N_28464,N_27896);
xor UO_2927 (O_2927,N_26790,N_26089);
or UO_2928 (O_2928,N_29518,N_29271);
nand UO_2929 (O_2929,N_28422,N_26079);
nand UO_2930 (O_2930,N_25484,N_25593);
nand UO_2931 (O_2931,N_28735,N_25746);
and UO_2932 (O_2932,N_26569,N_25167);
or UO_2933 (O_2933,N_26904,N_27213);
and UO_2934 (O_2934,N_26421,N_25683);
or UO_2935 (O_2935,N_29570,N_25331);
or UO_2936 (O_2936,N_29045,N_27011);
or UO_2937 (O_2937,N_29481,N_29051);
and UO_2938 (O_2938,N_26055,N_25620);
and UO_2939 (O_2939,N_28779,N_29268);
and UO_2940 (O_2940,N_29516,N_28278);
xnor UO_2941 (O_2941,N_26145,N_28655);
nand UO_2942 (O_2942,N_25620,N_28444);
or UO_2943 (O_2943,N_28020,N_25564);
nor UO_2944 (O_2944,N_29971,N_29948);
nand UO_2945 (O_2945,N_27480,N_25503);
nor UO_2946 (O_2946,N_28366,N_26054);
or UO_2947 (O_2947,N_26753,N_29599);
xnor UO_2948 (O_2948,N_25735,N_25482);
and UO_2949 (O_2949,N_25243,N_28403);
and UO_2950 (O_2950,N_25975,N_27601);
nand UO_2951 (O_2951,N_28677,N_26696);
or UO_2952 (O_2952,N_26166,N_25975);
or UO_2953 (O_2953,N_27740,N_25176);
nand UO_2954 (O_2954,N_29395,N_28517);
nand UO_2955 (O_2955,N_27601,N_26986);
or UO_2956 (O_2956,N_27888,N_26189);
nor UO_2957 (O_2957,N_27473,N_26461);
nand UO_2958 (O_2958,N_26610,N_26428);
nand UO_2959 (O_2959,N_26570,N_28777);
nor UO_2960 (O_2960,N_29051,N_26391);
or UO_2961 (O_2961,N_29024,N_27672);
or UO_2962 (O_2962,N_29436,N_25182);
nor UO_2963 (O_2963,N_27630,N_28502);
or UO_2964 (O_2964,N_25576,N_28387);
nor UO_2965 (O_2965,N_26857,N_27921);
nand UO_2966 (O_2966,N_26711,N_26060);
or UO_2967 (O_2967,N_29708,N_25543);
nor UO_2968 (O_2968,N_26377,N_27546);
and UO_2969 (O_2969,N_29700,N_26873);
and UO_2970 (O_2970,N_29528,N_26383);
and UO_2971 (O_2971,N_27145,N_27666);
and UO_2972 (O_2972,N_26159,N_27421);
and UO_2973 (O_2973,N_25177,N_26854);
or UO_2974 (O_2974,N_26021,N_27995);
nor UO_2975 (O_2975,N_27965,N_27207);
and UO_2976 (O_2976,N_28274,N_26561);
and UO_2977 (O_2977,N_29415,N_29251);
nand UO_2978 (O_2978,N_26920,N_26012);
nand UO_2979 (O_2979,N_26427,N_27162);
and UO_2980 (O_2980,N_25192,N_25588);
and UO_2981 (O_2981,N_26327,N_25316);
nand UO_2982 (O_2982,N_29513,N_27427);
and UO_2983 (O_2983,N_28470,N_27622);
nor UO_2984 (O_2984,N_25046,N_29973);
or UO_2985 (O_2985,N_28278,N_28581);
nor UO_2986 (O_2986,N_25301,N_27996);
and UO_2987 (O_2987,N_29512,N_25048);
or UO_2988 (O_2988,N_25104,N_25545);
nand UO_2989 (O_2989,N_28419,N_27325);
and UO_2990 (O_2990,N_29216,N_27134);
or UO_2991 (O_2991,N_29683,N_26432);
nand UO_2992 (O_2992,N_27829,N_29978);
nor UO_2993 (O_2993,N_28902,N_27670);
or UO_2994 (O_2994,N_27200,N_27726);
nand UO_2995 (O_2995,N_26968,N_25707);
and UO_2996 (O_2996,N_29366,N_28310);
nand UO_2997 (O_2997,N_26237,N_29400);
and UO_2998 (O_2998,N_29108,N_26013);
nor UO_2999 (O_2999,N_28048,N_28456);
nor UO_3000 (O_3000,N_28005,N_29569);
nor UO_3001 (O_3001,N_29154,N_29275);
nor UO_3002 (O_3002,N_25067,N_27210);
or UO_3003 (O_3003,N_28473,N_29448);
or UO_3004 (O_3004,N_25409,N_25435);
and UO_3005 (O_3005,N_26422,N_28102);
nand UO_3006 (O_3006,N_28534,N_26385);
nand UO_3007 (O_3007,N_27405,N_26606);
nor UO_3008 (O_3008,N_25313,N_25464);
and UO_3009 (O_3009,N_29681,N_25283);
nand UO_3010 (O_3010,N_28635,N_27631);
or UO_3011 (O_3011,N_27222,N_27308);
or UO_3012 (O_3012,N_27196,N_26899);
xor UO_3013 (O_3013,N_27524,N_25595);
and UO_3014 (O_3014,N_27359,N_28176);
nor UO_3015 (O_3015,N_28753,N_28650);
nand UO_3016 (O_3016,N_27832,N_28437);
or UO_3017 (O_3017,N_25849,N_28916);
nor UO_3018 (O_3018,N_25443,N_27806);
or UO_3019 (O_3019,N_28816,N_29111);
or UO_3020 (O_3020,N_26942,N_26684);
and UO_3021 (O_3021,N_29980,N_26599);
and UO_3022 (O_3022,N_27394,N_29112);
or UO_3023 (O_3023,N_26472,N_29110);
nand UO_3024 (O_3024,N_26280,N_27376);
nor UO_3025 (O_3025,N_25019,N_26400);
and UO_3026 (O_3026,N_27223,N_27755);
nor UO_3027 (O_3027,N_26440,N_25491);
nor UO_3028 (O_3028,N_27458,N_27017);
and UO_3029 (O_3029,N_26398,N_26587);
nor UO_3030 (O_3030,N_29469,N_26740);
or UO_3031 (O_3031,N_28505,N_26749);
or UO_3032 (O_3032,N_29472,N_27074);
or UO_3033 (O_3033,N_29559,N_29000);
or UO_3034 (O_3034,N_29836,N_27742);
nand UO_3035 (O_3035,N_28502,N_26878);
and UO_3036 (O_3036,N_28761,N_26400);
and UO_3037 (O_3037,N_29984,N_26948);
and UO_3038 (O_3038,N_25761,N_28312);
and UO_3039 (O_3039,N_29811,N_27413);
nor UO_3040 (O_3040,N_27473,N_27319);
and UO_3041 (O_3041,N_29892,N_27690);
and UO_3042 (O_3042,N_27014,N_25913);
nand UO_3043 (O_3043,N_25739,N_25025);
and UO_3044 (O_3044,N_28213,N_25215);
and UO_3045 (O_3045,N_27801,N_25006);
nor UO_3046 (O_3046,N_28315,N_28146);
nand UO_3047 (O_3047,N_26473,N_25828);
nor UO_3048 (O_3048,N_29610,N_25387);
and UO_3049 (O_3049,N_28897,N_28857);
and UO_3050 (O_3050,N_28033,N_29508);
or UO_3051 (O_3051,N_27857,N_26661);
nand UO_3052 (O_3052,N_27753,N_27641);
nand UO_3053 (O_3053,N_27427,N_26981);
nand UO_3054 (O_3054,N_28712,N_27186);
and UO_3055 (O_3055,N_27733,N_29465);
or UO_3056 (O_3056,N_29689,N_29560);
nand UO_3057 (O_3057,N_28875,N_29565);
nor UO_3058 (O_3058,N_27619,N_29515);
and UO_3059 (O_3059,N_26052,N_25567);
and UO_3060 (O_3060,N_27521,N_25419);
nand UO_3061 (O_3061,N_27315,N_28140);
nand UO_3062 (O_3062,N_25833,N_26855);
nand UO_3063 (O_3063,N_29596,N_26992);
nor UO_3064 (O_3064,N_27869,N_25355);
nand UO_3065 (O_3065,N_27006,N_29595);
nand UO_3066 (O_3066,N_26215,N_25856);
or UO_3067 (O_3067,N_26632,N_29115);
or UO_3068 (O_3068,N_29561,N_26408);
and UO_3069 (O_3069,N_27938,N_25202);
nand UO_3070 (O_3070,N_26063,N_28861);
or UO_3071 (O_3071,N_27854,N_29179);
nor UO_3072 (O_3072,N_29712,N_29123);
nor UO_3073 (O_3073,N_26470,N_28777);
nand UO_3074 (O_3074,N_27772,N_29530);
nor UO_3075 (O_3075,N_27458,N_25995);
nand UO_3076 (O_3076,N_27543,N_27922);
nand UO_3077 (O_3077,N_29333,N_26014);
and UO_3078 (O_3078,N_28038,N_28843);
nor UO_3079 (O_3079,N_27286,N_28140);
nor UO_3080 (O_3080,N_26302,N_25334);
and UO_3081 (O_3081,N_25439,N_29780);
or UO_3082 (O_3082,N_26297,N_26301);
or UO_3083 (O_3083,N_27919,N_27848);
nor UO_3084 (O_3084,N_25974,N_29084);
or UO_3085 (O_3085,N_29974,N_28531);
nand UO_3086 (O_3086,N_27659,N_26851);
or UO_3087 (O_3087,N_26896,N_25755);
nor UO_3088 (O_3088,N_29514,N_29984);
nand UO_3089 (O_3089,N_27196,N_26727);
and UO_3090 (O_3090,N_28226,N_26995);
and UO_3091 (O_3091,N_27743,N_29645);
nand UO_3092 (O_3092,N_25778,N_25399);
nor UO_3093 (O_3093,N_26306,N_27435);
nand UO_3094 (O_3094,N_25211,N_28291);
or UO_3095 (O_3095,N_29860,N_28881);
and UO_3096 (O_3096,N_29539,N_27753);
or UO_3097 (O_3097,N_29694,N_29327);
or UO_3098 (O_3098,N_28579,N_25648);
nand UO_3099 (O_3099,N_26760,N_26342);
and UO_3100 (O_3100,N_29702,N_27030);
and UO_3101 (O_3101,N_26456,N_25883);
and UO_3102 (O_3102,N_28810,N_26637);
nand UO_3103 (O_3103,N_28106,N_29116);
and UO_3104 (O_3104,N_27841,N_29403);
nand UO_3105 (O_3105,N_26485,N_26949);
nor UO_3106 (O_3106,N_29966,N_27055);
or UO_3107 (O_3107,N_26580,N_26599);
nor UO_3108 (O_3108,N_27631,N_28204);
and UO_3109 (O_3109,N_25562,N_29378);
xor UO_3110 (O_3110,N_29616,N_28691);
or UO_3111 (O_3111,N_26000,N_29388);
nor UO_3112 (O_3112,N_29788,N_25451);
or UO_3113 (O_3113,N_27365,N_26484);
or UO_3114 (O_3114,N_28861,N_29285);
nor UO_3115 (O_3115,N_28587,N_26982);
nand UO_3116 (O_3116,N_29496,N_27413);
nand UO_3117 (O_3117,N_28280,N_28691);
nor UO_3118 (O_3118,N_27551,N_28416);
nand UO_3119 (O_3119,N_25733,N_27084);
or UO_3120 (O_3120,N_27084,N_26540);
xnor UO_3121 (O_3121,N_29093,N_27718);
or UO_3122 (O_3122,N_26951,N_27310);
and UO_3123 (O_3123,N_29392,N_27782);
or UO_3124 (O_3124,N_26207,N_27086);
or UO_3125 (O_3125,N_27418,N_28150);
nand UO_3126 (O_3126,N_28307,N_29998);
nand UO_3127 (O_3127,N_29265,N_27137);
nor UO_3128 (O_3128,N_27525,N_26091);
nor UO_3129 (O_3129,N_26431,N_27426);
and UO_3130 (O_3130,N_27111,N_29370);
or UO_3131 (O_3131,N_27677,N_27498);
nand UO_3132 (O_3132,N_28367,N_28764);
nor UO_3133 (O_3133,N_26121,N_28761);
nand UO_3134 (O_3134,N_25927,N_25574);
nand UO_3135 (O_3135,N_29625,N_27900);
nor UO_3136 (O_3136,N_27841,N_25085);
and UO_3137 (O_3137,N_25633,N_29849);
nand UO_3138 (O_3138,N_29200,N_26793);
nand UO_3139 (O_3139,N_27523,N_26450);
and UO_3140 (O_3140,N_25454,N_25822);
nor UO_3141 (O_3141,N_27841,N_27664);
nand UO_3142 (O_3142,N_26295,N_29792);
nand UO_3143 (O_3143,N_28839,N_29977);
nor UO_3144 (O_3144,N_26829,N_26109);
and UO_3145 (O_3145,N_26923,N_26143);
and UO_3146 (O_3146,N_27214,N_25193);
nor UO_3147 (O_3147,N_27776,N_25737);
nor UO_3148 (O_3148,N_28200,N_25594);
nand UO_3149 (O_3149,N_29427,N_29945);
or UO_3150 (O_3150,N_28383,N_26246);
nand UO_3151 (O_3151,N_29603,N_26405);
or UO_3152 (O_3152,N_28692,N_29315);
nand UO_3153 (O_3153,N_25408,N_29310);
or UO_3154 (O_3154,N_27321,N_29222);
nor UO_3155 (O_3155,N_28644,N_28218);
xor UO_3156 (O_3156,N_25872,N_28094);
nand UO_3157 (O_3157,N_27006,N_27289);
nand UO_3158 (O_3158,N_26077,N_25052);
and UO_3159 (O_3159,N_28153,N_29489);
or UO_3160 (O_3160,N_28418,N_26737);
and UO_3161 (O_3161,N_25397,N_28955);
nand UO_3162 (O_3162,N_29284,N_29731);
and UO_3163 (O_3163,N_27128,N_25069);
nand UO_3164 (O_3164,N_27754,N_27640);
nand UO_3165 (O_3165,N_29810,N_29683);
and UO_3166 (O_3166,N_28035,N_28637);
or UO_3167 (O_3167,N_25111,N_25777);
and UO_3168 (O_3168,N_25485,N_28550);
or UO_3169 (O_3169,N_29955,N_29196);
and UO_3170 (O_3170,N_29577,N_28521);
and UO_3171 (O_3171,N_29147,N_27942);
nand UO_3172 (O_3172,N_28907,N_25139);
nor UO_3173 (O_3173,N_26197,N_29753);
nor UO_3174 (O_3174,N_26818,N_27350);
or UO_3175 (O_3175,N_28232,N_27639);
nor UO_3176 (O_3176,N_29664,N_27843);
nand UO_3177 (O_3177,N_25745,N_29140);
nand UO_3178 (O_3178,N_28746,N_28084);
or UO_3179 (O_3179,N_27865,N_28311);
and UO_3180 (O_3180,N_25708,N_29621);
or UO_3181 (O_3181,N_27849,N_26777);
nor UO_3182 (O_3182,N_28872,N_29503);
and UO_3183 (O_3183,N_27936,N_28417);
nor UO_3184 (O_3184,N_27207,N_25064);
nor UO_3185 (O_3185,N_25486,N_25172);
nor UO_3186 (O_3186,N_27635,N_26095);
nor UO_3187 (O_3187,N_26332,N_26390);
and UO_3188 (O_3188,N_28656,N_27072);
and UO_3189 (O_3189,N_28891,N_28572);
or UO_3190 (O_3190,N_28284,N_27091);
or UO_3191 (O_3191,N_28071,N_28561);
nor UO_3192 (O_3192,N_27427,N_29666);
nand UO_3193 (O_3193,N_29184,N_28705);
nor UO_3194 (O_3194,N_28001,N_29022);
and UO_3195 (O_3195,N_28231,N_27711);
nor UO_3196 (O_3196,N_26154,N_27860);
nor UO_3197 (O_3197,N_29368,N_25700);
and UO_3198 (O_3198,N_28234,N_26972);
or UO_3199 (O_3199,N_26093,N_29592);
or UO_3200 (O_3200,N_27197,N_25512);
nor UO_3201 (O_3201,N_29292,N_28968);
and UO_3202 (O_3202,N_29976,N_29871);
or UO_3203 (O_3203,N_26482,N_27412);
nand UO_3204 (O_3204,N_29674,N_25035);
nor UO_3205 (O_3205,N_28900,N_27594);
nand UO_3206 (O_3206,N_29572,N_28156);
nand UO_3207 (O_3207,N_29181,N_28504);
nor UO_3208 (O_3208,N_29055,N_27088);
nand UO_3209 (O_3209,N_25120,N_26085);
nor UO_3210 (O_3210,N_25517,N_29275);
nor UO_3211 (O_3211,N_29798,N_27231);
or UO_3212 (O_3212,N_27747,N_29029);
and UO_3213 (O_3213,N_28356,N_25491);
nand UO_3214 (O_3214,N_25322,N_26603);
and UO_3215 (O_3215,N_25076,N_26150);
nor UO_3216 (O_3216,N_27068,N_27006);
and UO_3217 (O_3217,N_27808,N_26096);
nor UO_3218 (O_3218,N_26291,N_27928);
or UO_3219 (O_3219,N_29450,N_29554);
nor UO_3220 (O_3220,N_29060,N_25820);
or UO_3221 (O_3221,N_25098,N_28540);
nor UO_3222 (O_3222,N_26167,N_28055);
nor UO_3223 (O_3223,N_27720,N_25911);
nand UO_3224 (O_3224,N_29533,N_27687);
nand UO_3225 (O_3225,N_29614,N_25890);
and UO_3226 (O_3226,N_29165,N_26595);
and UO_3227 (O_3227,N_29653,N_29923);
nor UO_3228 (O_3228,N_29074,N_27731);
nor UO_3229 (O_3229,N_27108,N_27068);
nor UO_3230 (O_3230,N_25950,N_28845);
and UO_3231 (O_3231,N_25744,N_27851);
nand UO_3232 (O_3232,N_28168,N_28309);
nor UO_3233 (O_3233,N_25610,N_26171);
nand UO_3234 (O_3234,N_26661,N_27258);
nor UO_3235 (O_3235,N_25639,N_29529);
or UO_3236 (O_3236,N_26212,N_29461);
nor UO_3237 (O_3237,N_25495,N_25480);
nand UO_3238 (O_3238,N_28392,N_27027);
or UO_3239 (O_3239,N_29473,N_29041);
or UO_3240 (O_3240,N_28766,N_28637);
or UO_3241 (O_3241,N_27828,N_25821);
or UO_3242 (O_3242,N_29123,N_29916);
nor UO_3243 (O_3243,N_28542,N_28004);
nand UO_3244 (O_3244,N_27875,N_29893);
nor UO_3245 (O_3245,N_29300,N_29200);
or UO_3246 (O_3246,N_27333,N_29636);
and UO_3247 (O_3247,N_29440,N_28424);
or UO_3248 (O_3248,N_27045,N_26068);
nand UO_3249 (O_3249,N_26350,N_29899);
or UO_3250 (O_3250,N_29929,N_26143);
or UO_3251 (O_3251,N_27240,N_25133);
nand UO_3252 (O_3252,N_28928,N_28516);
or UO_3253 (O_3253,N_27355,N_28836);
xnor UO_3254 (O_3254,N_26734,N_25225);
or UO_3255 (O_3255,N_29702,N_27355);
and UO_3256 (O_3256,N_28045,N_28664);
nand UO_3257 (O_3257,N_27418,N_28811);
nor UO_3258 (O_3258,N_29869,N_28854);
nand UO_3259 (O_3259,N_26458,N_29488);
and UO_3260 (O_3260,N_29818,N_29457);
and UO_3261 (O_3261,N_29433,N_27208);
nand UO_3262 (O_3262,N_25317,N_25087);
or UO_3263 (O_3263,N_26905,N_29890);
and UO_3264 (O_3264,N_27576,N_29554);
and UO_3265 (O_3265,N_28430,N_28329);
nor UO_3266 (O_3266,N_26449,N_28526);
or UO_3267 (O_3267,N_26004,N_29820);
nand UO_3268 (O_3268,N_28956,N_27655);
nand UO_3269 (O_3269,N_28927,N_27001);
and UO_3270 (O_3270,N_26329,N_29870);
nand UO_3271 (O_3271,N_26078,N_26235);
nor UO_3272 (O_3272,N_25411,N_28475);
or UO_3273 (O_3273,N_27679,N_29045);
nand UO_3274 (O_3274,N_25047,N_25404);
or UO_3275 (O_3275,N_28360,N_26301);
nand UO_3276 (O_3276,N_26142,N_26912);
nand UO_3277 (O_3277,N_28125,N_26982);
and UO_3278 (O_3278,N_29029,N_25966);
nand UO_3279 (O_3279,N_26492,N_27960);
and UO_3280 (O_3280,N_25176,N_27489);
or UO_3281 (O_3281,N_29452,N_26228);
or UO_3282 (O_3282,N_26779,N_28428);
or UO_3283 (O_3283,N_26241,N_25953);
and UO_3284 (O_3284,N_25804,N_29798);
nor UO_3285 (O_3285,N_28000,N_29278);
nor UO_3286 (O_3286,N_28154,N_25348);
or UO_3287 (O_3287,N_27774,N_29743);
nand UO_3288 (O_3288,N_29812,N_28224);
and UO_3289 (O_3289,N_25796,N_25170);
and UO_3290 (O_3290,N_27467,N_27057);
nand UO_3291 (O_3291,N_26237,N_26714);
or UO_3292 (O_3292,N_29047,N_28106);
nor UO_3293 (O_3293,N_29727,N_29600);
or UO_3294 (O_3294,N_28392,N_28731);
nor UO_3295 (O_3295,N_25040,N_26546);
or UO_3296 (O_3296,N_29389,N_25819);
and UO_3297 (O_3297,N_28049,N_25955);
nand UO_3298 (O_3298,N_27646,N_27687);
nor UO_3299 (O_3299,N_29879,N_29296);
or UO_3300 (O_3300,N_26602,N_29839);
and UO_3301 (O_3301,N_25232,N_29022);
or UO_3302 (O_3302,N_27473,N_26627);
and UO_3303 (O_3303,N_26412,N_27274);
or UO_3304 (O_3304,N_27784,N_27073);
or UO_3305 (O_3305,N_28025,N_27548);
nand UO_3306 (O_3306,N_29814,N_25551);
nand UO_3307 (O_3307,N_27439,N_27828);
nor UO_3308 (O_3308,N_28415,N_29687);
and UO_3309 (O_3309,N_26774,N_29960);
and UO_3310 (O_3310,N_28715,N_26179);
nand UO_3311 (O_3311,N_29381,N_28624);
nor UO_3312 (O_3312,N_28480,N_27882);
or UO_3313 (O_3313,N_26564,N_25846);
and UO_3314 (O_3314,N_29840,N_25260);
and UO_3315 (O_3315,N_29205,N_29918);
or UO_3316 (O_3316,N_26202,N_26906);
nand UO_3317 (O_3317,N_26247,N_26656);
and UO_3318 (O_3318,N_29763,N_26953);
and UO_3319 (O_3319,N_26478,N_25639);
or UO_3320 (O_3320,N_25481,N_25799);
nor UO_3321 (O_3321,N_26846,N_29148);
nand UO_3322 (O_3322,N_28438,N_28729);
nor UO_3323 (O_3323,N_29553,N_26496);
and UO_3324 (O_3324,N_29284,N_27431);
nor UO_3325 (O_3325,N_25895,N_28026);
nor UO_3326 (O_3326,N_29668,N_28250);
nand UO_3327 (O_3327,N_26139,N_27029);
nand UO_3328 (O_3328,N_29841,N_29038);
nor UO_3329 (O_3329,N_27013,N_29452);
and UO_3330 (O_3330,N_26049,N_29531);
nor UO_3331 (O_3331,N_28775,N_27396);
or UO_3332 (O_3332,N_28886,N_29030);
or UO_3333 (O_3333,N_26549,N_25759);
and UO_3334 (O_3334,N_26581,N_26091);
nand UO_3335 (O_3335,N_28969,N_28441);
or UO_3336 (O_3336,N_28139,N_29093);
nand UO_3337 (O_3337,N_29637,N_28911);
nand UO_3338 (O_3338,N_28542,N_26390);
or UO_3339 (O_3339,N_29054,N_27060);
nand UO_3340 (O_3340,N_26175,N_25649);
or UO_3341 (O_3341,N_25354,N_25998);
and UO_3342 (O_3342,N_27773,N_28313);
nand UO_3343 (O_3343,N_26811,N_28367);
nor UO_3344 (O_3344,N_27451,N_27291);
nor UO_3345 (O_3345,N_28556,N_26144);
or UO_3346 (O_3346,N_28462,N_26024);
or UO_3347 (O_3347,N_26756,N_26598);
or UO_3348 (O_3348,N_25538,N_26690);
nand UO_3349 (O_3349,N_25498,N_27478);
and UO_3350 (O_3350,N_28884,N_26506);
nor UO_3351 (O_3351,N_26669,N_29871);
and UO_3352 (O_3352,N_27729,N_25886);
or UO_3353 (O_3353,N_27838,N_25553);
and UO_3354 (O_3354,N_26004,N_25074);
nor UO_3355 (O_3355,N_26697,N_25810);
and UO_3356 (O_3356,N_25102,N_28017);
nand UO_3357 (O_3357,N_29717,N_27492);
nor UO_3358 (O_3358,N_28967,N_25575);
nor UO_3359 (O_3359,N_29099,N_27234);
or UO_3360 (O_3360,N_25774,N_27986);
nand UO_3361 (O_3361,N_27894,N_27117);
or UO_3362 (O_3362,N_25073,N_25172);
nand UO_3363 (O_3363,N_29224,N_26384);
and UO_3364 (O_3364,N_26255,N_25940);
or UO_3365 (O_3365,N_27394,N_26882);
or UO_3366 (O_3366,N_28328,N_29272);
nand UO_3367 (O_3367,N_26539,N_29281);
or UO_3368 (O_3368,N_26552,N_25301);
nand UO_3369 (O_3369,N_26344,N_29868);
or UO_3370 (O_3370,N_28166,N_28024);
and UO_3371 (O_3371,N_25986,N_29586);
nand UO_3372 (O_3372,N_27924,N_28132);
or UO_3373 (O_3373,N_29591,N_28559);
and UO_3374 (O_3374,N_26291,N_26900);
or UO_3375 (O_3375,N_26193,N_28651);
nand UO_3376 (O_3376,N_25094,N_26406);
nor UO_3377 (O_3377,N_25187,N_29979);
nand UO_3378 (O_3378,N_27573,N_28585);
or UO_3379 (O_3379,N_26246,N_28508);
and UO_3380 (O_3380,N_26907,N_27964);
nand UO_3381 (O_3381,N_27643,N_25931);
nand UO_3382 (O_3382,N_26148,N_29686);
and UO_3383 (O_3383,N_29324,N_29677);
nor UO_3384 (O_3384,N_28151,N_26313);
nor UO_3385 (O_3385,N_26021,N_26055);
xnor UO_3386 (O_3386,N_29211,N_26263);
and UO_3387 (O_3387,N_29766,N_29800);
and UO_3388 (O_3388,N_27289,N_25391);
and UO_3389 (O_3389,N_25006,N_29539);
and UO_3390 (O_3390,N_26992,N_29312);
xnor UO_3391 (O_3391,N_26735,N_25729);
or UO_3392 (O_3392,N_26677,N_26492);
nor UO_3393 (O_3393,N_27302,N_26174);
nand UO_3394 (O_3394,N_28836,N_26749);
nand UO_3395 (O_3395,N_27796,N_29951);
or UO_3396 (O_3396,N_25787,N_29642);
and UO_3397 (O_3397,N_28233,N_27644);
and UO_3398 (O_3398,N_25598,N_25530);
nor UO_3399 (O_3399,N_28582,N_25915);
or UO_3400 (O_3400,N_26936,N_26548);
nor UO_3401 (O_3401,N_29009,N_27248);
nand UO_3402 (O_3402,N_27563,N_25793);
or UO_3403 (O_3403,N_28251,N_29922);
or UO_3404 (O_3404,N_28157,N_26505);
or UO_3405 (O_3405,N_29029,N_25699);
nand UO_3406 (O_3406,N_27673,N_29425);
nand UO_3407 (O_3407,N_28283,N_28259);
and UO_3408 (O_3408,N_29076,N_26709);
nand UO_3409 (O_3409,N_29943,N_29518);
nor UO_3410 (O_3410,N_28939,N_27608);
or UO_3411 (O_3411,N_26907,N_29047);
nand UO_3412 (O_3412,N_27444,N_29364);
nand UO_3413 (O_3413,N_29590,N_29020);
or UO_3414 (O_3414,N_26653,N_25274);
nand UO_3415 (O_3415,N_26904,N_28761);
nor UO_3416 (O_3416,N_27484,N_26569);
or UO_3417 (O_3417,N_28792,N_26328);
nand UO_3418 (O_3418,N_26274,N_27545);
nand UO_3419 (O_3419,N_27000,N_29342);
or UO_3420 (O_3420,N_27520,N_29228);
nor UO_3421 (O_3421,N_26636,N_27726);
or UO_3422 (O_3422,N_25832,N_27046);
and UO_3423 (O_3423,N_29198,N_26705);
and UO_3424 (O_3424,N_28623,N_26795);
nor UO_3425 (O_3425,N_29492,N_25998);
nor UO_3426 (O_3426,N_26305,N_29393);
or UO_3427 (O_3427,N_27151,N_28794);
and UO_3428 (O_3428,N_29217,N_26509);
and UO_3429 (O_3429,N_28998,N_27892);
nor UO_3430 (O_3430,N_29295,N_28501);
nand UO_3431 (O_3431,N_29140,N_28548);
nand UO_3432 (O_3432,N_28333,N_28234);
nand UO_3433 (O_3433,N_29099,N_26997);
nand UO_3434 (O_3434,N_25745,N_26059);
or UO_3435 (O_3435,N_29035,N_28873);
or UO_3436 (O_3436,N_25519,N_28201);
nand UO_3437 (O_3437,N_29973,N_29420);
and UO_3438 (O_3438,N_29420,N_28555);
nor UO_3439 (O_3439,N_26901,N_28630);
xor UO_3440 (O_3440,N_25156,N_29274);
or UO_3441 (O_3441,N_26041,N_28924);
nor UO_3442 (O_3442,N_25197,N_25150);
nand UO_3443 (O_3443,N_29972,N_25701);
nand UO_3444 (O_3444,N_25426,N_26634);
or UO_3445 (O_3445,N_25423,N_29980);
nor UO_3446 (O_3446,N_25655,N_25501);
nand UO_3447 (O_3447,N_25705,N_29559);
and UO_3448 (O_3448,N_26907,N_26153);
and UO_3449 (O_3449,N_28351,N_26066);
nand UO_3450 (O_3450,N_28079,N_29043);
and UO_3451 (O_3451,N_28704,N_26355);
and UO_3452 (O_3452,N_28090,N_25013);
nor UO_3453 (O_3453,N_28138,N_27401);
and UO_3454 (O_3454,N_26155,N_26434);
nand UO_3455 (O_3455,N_28088,N_25851);
nor UO_3456 (O_3456,N_27325,N_25362);
nor UO_3457 (O_3457,N_25332,N_26397);
or UO_3458 (O_3458,N_26409,N_26910);
or UO_3459 (O_3459,N_28876,N_29663);
nand UO_3460 (O_3460,N_28095,N_27597);
nor UO_3461 (O_3461,N_25759,N_29152);
and UO_3462 (O_3462,N_29722,N_25108);
or UO_3463 (O_3463,N_29595,N_27224);
nor UO_3464 (O_3464,N_26405,N_28895);
nand UO_3465 (O_3465,N_25699,N_29911);
xor UO_3466 (O_3466,N_25288,N_28211);
nor UO_3467 (O_3467,N_28209,N_25705);
and UO_3468 (O_3468,N_25737,N_25377);
nand UO_3469 (O_3469,N_26234,N_25510);
nor UO_3470 (O_3470,N_28498,N_26288);
nand UO_3471 (O_3471,N_26463,N_28740);
nand UO_3472 (O_3472,N_27644,N_25236);
or UO_3473 (O_3473,N_29303,N_28111);
and UO_3474 (O_3474,N_27210,N_28391);
and UO_3475 (O_3475,N_28353,N_29669);
nand UO_3476 (O_3476,N_29901,N_27003);
and UO_3477 (O_3477,N_25575,N_29505);
and UO_3478 (O_3478,N_28025,N_26573);
and UO_3479 (O_3479,N_27042,N_25291);
nor UO_3480 (O_3480,N_28578,N_25195);
and UO_3481 (O_3481,N_29604,N_27213);
or UO_3482 (O_3482,N_27429,N_25731);
nor UO_3483 (O_3483,N_28345,N_26160);
nor UO_3484 (O_3484,N_26005,N_25455);
nor UO_3485 (O_3485,N_27877,N_28419);
nor UO_3486 (O_3486,N_25002,N_25094);
nand UO_3487 (O_3487,N_28882,N_28477);
nand UO_3488 (O_3488,N_25268,N_29619);
or UO_3489 (O_3489,N_27915,N_29918);
and UO_3490 (O_3490,N_25646,N_29716);
nand UO_3491 (O_3491,N_28680,N_26345);
nand UO_3492 (O_3492,N_27467,N_25149);
nor UO_3493 (O_3493,N_28199,N_28712);
nand UO_3494 (O_3494,N_29602,N_28536);
nand UO_3495 (O_3495,N_28832,N_29322);
nor UO_3496 (O_3496,N_27012,N_28793);
nand UO_3497 (O_3497,N_28908,N_26479);
or UO_3498 (O_3498,N_29472,N_26929);
nand UO_3499 (O_3499,N_29143,N_25744);
endmodule