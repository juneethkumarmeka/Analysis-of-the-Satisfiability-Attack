module basic_500_3000_500_30_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_298,In_50);
or U1 (N_1,In_333,In_390);
and U2 (N_2,In_193,In_285);
nor U3 (N_3,In_138,In_228);
and U4 (N_4,In_55,In_168);
nor U5 (N_5,In_48,In_244);
nor U6 (N_6,In_195,In_347);
or U7 (N_7,In_352,In_305);
or U8 (N_8,In_99,In_259);
and U9 (N_9,In_145,In_426);
or U10 (N_10,In_136,In_419);
nand U11 (N_11,In_471,In_463);
nand U12 (N_12,In_179,In_234);
xor U13 (N_13,In_407,In_81);
or U14 (N_14,In_265,In_297);
or U15 (N_15,In_118,In_410);
nand U16 (N_16,In_78,In_393);
and U17 (N_17,In_467,In_233);
nand U18 (N_18,In_14,In_316);
and U19 (N_19,In_158,In_328);
and U20 (N_20,In_214,In_38);
and U21 (N_21,In_20,In_435);
xnor U22 (N_22,In_483,In_433);
xnor U23 (N_23,In_377,In_343);
and U24 (N_24,In_243,In_27);
and U25 (N_25,In_153,In_238);
nor U26 (N_26,In_330,In_446);
nand U27 (N_27,In_187,In_223);
nor U28 (N_28,In_424,In_92);
or U29 (N_29,In_415,In_348);
nand U30 (N_30,In_46,In_148);
nor U31 (N_31,In_7,In_459);
or U32 (N_32,In_462,In_40);
or U33 (N_33,In_411,In_263);
or U34 (N_34,In_277,In_339);
nor U35 (N_35,In_199,In_247);
or U36 (N_36,In_337,In_425);
nor U37 (N_37,In_60,In_432);
nand U38 (N_38,In_300,In_69);
and U39 (N_39,In_23,In_77);
nor U40 (N_40,In_438,In_366);
or U41 (N_41,In_96,In_254);
and U42 (N_42,In_437,In_37);
and U43 (N_43,In_113,In_342);
nor U44 (N_44,In_184,In_66);
nor U45 (N_45,In_353,In_323);
xnor U46 (N_46,In_98,In_196);
nand U47 (N_47,In_306,In_61);
xor U48 (N_48,In_452,In_135);
and U49 (N_49,In_255,In_279);
or U50 (N_50,In_192,In_268);
nand U51 (N_51,In_156,In_222);
and U52 (N_52,In_370,In_127);
or U53 (N_53,In_56,In_34);
or U54 (N_54,In_16,In_71);
nand U55 (N_55,In_320,In_22);
nand U56 (N_56,In_26,In_104);
or U57 (N_57,In_338,In_45);
xnor U58 (N_58,In_423,In_369);
nand U59 (N_59,In_232,In_210);
xor U60 (N_60,In_64,In_162);
nor U61 (N_61,In_224,In_35);
nor U62 (N_62,In_239,In_21);
and U63 (N_63,In_290,In_125);
nand U64 (N_64,In_44,In_481);
nand U65 (N_65,In_427,In_310);
nand U66 (N_66,In_129,In_190);
or U67 (N_67,In_384,In_264);
xor U68 (N_68,In_404,In_381);
and U69 (N_69,In_399,In_39);
nor U70 (N_70,In_387,In_451);
nand U71 (N_71,In_346,In_362);
nand U72 (N_72,In_165,In_495);
and U73 (N_73,In_147,In_47);
nor U74 (N_74,In_2,In_253);
nor U75 (N_75,In_314,In_349);
nor U76 (N_76,In_431,In_272);
nor U77 (N_77,In_496,In_294);
xnor U78 (N_78,In_336,In_230);
xnor U79 (N_79,In_17,In_31);
or U80 (N_80,In_422,In_477);
and U81 (N_81,In_140,In_183);
nor U82 (N_82,In_189,In_97);
and U83 (N_83,In_276,In_151);
and U84 (N_84,In_197,In_295);
nor U85 (N_85,In_200,In_345);
and U86 (N_86,In_59,In_360);
or U87 (N_87,In_315,In_332);
and U88 (N_88,In_486,In_269);
nor U89 (N_89,In_169,In_103);
nand U90 (N_90,In_335,In_174);
nor U91 (N_91,In_101,In_159);
or U92 (N_92,In_492,In_490);
and U93 (N_93,In_100,In_488);
or U94 (N_94,In_473,In_378);
nor U95 (N_95,In_363,In_464);
and U96 (N_96,In_304,In_24);
nor U97 (N_97,In_386,In_458);
nand U98 (N_98,In_341,In_376);
xnor U99 (N_99,In_57,In_73);
or U100 (N_100,In_429,In_167);
and U101 (N_101,In_442,In_211);
nand U102 (N_102,In_367,N_56);
nor U103 (N_103,In_131,In_216);
nand U104 (N_104,In_261,In_475);
and U105 (N_105,In_252,In_284);
xor U106 (N_106,N_21,N_19);
nand U107 (N_107,In_283,In_416);
xor U108 (N_108,In_188,In_219);
or U109 (N_109,In_89,In_389);
nand U110 (N_110,In_319,In_149);
nand U111 (N_111,In_357,In_240);
or U112 (N_112,In_445,N_17);
nor U113 (N_113,In_288,In_13);
nor U114 (N_114,N_0,N_35);
nor U115 (N_115,In_65,N_52);
nand U116 (N_116,In_373,In_182);
or U117 (N_117,In_198,In_251);
nor U118 (N_118,In_141,In_405);
nor U119 (N_119,In_291,In_355);
nand U120 (N_120,In_280,N_11);
nand U121 (N_121,In_146,In_201);
nor U122 (N_122,N_2,N_38);
xor U123 (N_123,In_241,In_220);
or U124 (N_124,In_217,In_249);
or U125 (N_125,In_160,N_95);
nor U126 (N_126,N_68,In_173);
nor U127 (N_127,In_105,In_106);
nor U128 (N_128,In_95,N_93);
or U129 (N_129,In_289,In_62);
and U130 (N_130,N_66,In_430);
nand U131 (N_131,In_41,N_57);
nor U132 (N_132,N_76,N_41);
nand U133 (N_133,In_235,In_309);
nor U134 (N_134,In_317,In_365);
nand U135 (N_135,In_397,In_443);
nand U136 (N_136,N_9,N_33);
or U137 (N_137,In_292,In_112);
nand U138 (N_138,N_96,In_177);
or U139 (N_139,In_266,In_63);
nand U140 (N_140,In_245,N_55);
and U141 (N_141,In_417,In_213);
xor U142 (N_142,In_440,N_44);
nor U143 (N_143,N_97,N_3);
nand U144 (N_144,In_364,In_42);
and U145 (N_145,In_83,N_16);
nor U146 (N_146,In_215,N_4);
xnor U147 (N_147,In_242,In_246);
nand U148 (N_148,N_70,N_13);
or U149 (N_149,In_406,In_9);
and U150 (N_150,In_128,N_45);
nor U151 (N_151,N_53,N_63);
or U152 (N_152,In_494,In_392);
nor U153 (N_153,In_258,N_89);
nand U154 (N_154,N_42,In_383);
or U155 (N_155,In_137,In_321);
or U156 (N_156,In_227,N_50);
or U157 (N_157,In_139,N_83);
nor U158 (N_158,In_303,In_191);
xnor U159 (N_159,In_88,In_30);
xnor U160 (N_160,N_77,In_461);
or U161 (N_161,In_311,N_99);
nand U162 (N_162,N_75,In_371);
or U163 (N_163,In_326,In_19);
nand U164 (N_164,In_409,In_385);
or U165 (N_165,In_122,N_28);
and U166 (N_166,In_395,In_194);
and U167 (N_167,In_221,In_93);
nor U168 (N_168,In_358,In_176);
or U169 (N_169,In_163,N_80);
nand U170 (N_170,In_5,In_267);
and U171 (N_171,N_37,In_344);
nand U172 (N_172,In_32,In_359);
or U173 (N_173,In_206,In_121);
nand U174 (N_174,In_324,In_157);
nor U175 (N_175,N_22,In_396);
nand U176 (N_176,In_49,In_79);
or U177 (N_177,In_448,In_497);
xnor U178 (N_178,In_109,In_447);
or U179 (N_179,In_456,N_49);
xnor U180 (N_180,In_408,In_286);
nand U181 (N_181,In_361,In_115);
nor U182 (N_182,In_453,In_0);
nand U183 (N_183,In_327,In_472);
nor U184 (N_184,In_282,In_166);
or U185 (N_185,N_8,In_480);
nand U186 (N_186,In_33,N_86);
nor U187 (N_187,In_296,In_351);
xnor U188 (N_188,In_1,N_7);
nor U189 (N_189,In_421,In_379);
nor U190 (N_190,In_51,In_82);
nor U191 (N_191,In_231,N_12);
nor U192 (N_192,In_8,N_84);
nand U193 (N_193,In_302,In_428);
nand U194 (N_194,In_53,In_150);
and U195 (N_195,In_52,In_76);
nor U196 (N_196,In_170,In_225);
nand U197 (N_197,In_491,N_36);
nor U198 (N_198,In_275,In_207);
or U199 (N_199,In_439,In_466);
nand U200 (N_200,In_18,N_193);
nand U201 (N_201,In_340,N_104);
nor U202 (N_202,In_256,N_136);
xnor U203 (N_203,In_154,In_400);
nand U204 (N_204,N_172,In_178);
or U205 (N_205,N_169,In_91);
nor U206 (N_206,In_229,In_420);
or U207 (N_207,N_30,N_102);
nor U208 (N_208,In_487,N_23);
nand U209 (N_209,In_15,In_274);
or U210 (N_210,In_72,N_118);
nand U211 (N_211,N_135,In_450);
and U212 (N_212,N_58,In_325);
nand U213 (N_213,N_62,In_331);
nand U214 (N_214,N_82,N_142);
nand U215 (N_215,In_68,In_54);
xor U216 (N_216,N_168,In_10);
or U217 (N_217,N_171,N_25);
or U218 (N_218,In_322,N_189);
nor U219 (N_219,In_354,N_188);
or U220 (N_220,N_127,N_54);
and U221 (N_221,N_129,N_147);
or U222 (N_222,N_59,N_1);
xnor U223 (N_223,N_115,N_153);
xor U224 (N_224,N_103,N_174);
nor U225 (N_225,N_29,N_90);
nand U226 (N_226,N_134,In_3);
nor U227 (N_227,In_380,In_454);
and U228 (N_228,N_109,N_27);
nor U229 (N_229,In_130,In_226);
or U230 (N_230,N_15,N_151);
nor U231 (N_231,N_114,In_143);
xor U232 (N_232,N_195,N_121);
and U233 (N_233,In_181,N_71);
xor U234 (N_234,In_126,N_156);
nor U235 (N_235,N_186,In_468);
and U236 (N_236,N_164,In_161);
nand U237 (N_237,In_312,In_485);
and U238 (N_238,N_5,In_12);
and U239 (N_239,In_270,In_208);
nand U240 (N_240,In_413,N_144);
or U241 (N_241,N_150,N_34);
nor U242 (N_242,N_73,N_170);
or U243 (N_243,N_74,N_111);
nand U244 (N_244,N_179,N_196);
and U245 (N_245,N_175,In_482);
and U246 (N_246,In_391,In_85);
xor U247 (N_247,N_110,N_119);
nand U248 (N_248,In_278,In_479);
nand U249 (N_249,In_436,N_100);
and U250 (N_250,N_137,N_10);
xnor U251 (N_251,In_368,N_32);
nor U252 (N_252,N_60,In_86);
and U253 (N_253,In_171,N_145);
or U254 (N_254,N_177,In_449);
nand U255 (N_255,N_180,N_126);
and U256 (N_256,N_46,N_141);
or U257 (N_257,N_154,N_187);
and U258 (N_258,In_388,In_152);
or U259 (N_259,In_382,N_183);
or U260 (N_260,N_140,In_202);
nor U261 (N_261,In_204,In_257);
or U262 (N_262,In_374,N_162);
and U263 (N_263,In_418,In_142);
nor U264 (N_264,In_25,In_444);
nor U265 (N_265,N_94,In_102);
xor U266 (N_266,N_143,In_28);
xor U267 (N_267,N_69,N_51);
nor U268 (N_268,In_111,N_47);
and U269 (N_269,N_199,N_107);
xnor U270 (N_270,In_180,In_356);
and U271 (N_271,N_160,In_403);
nand U272 (N_272,In_108,N_91);
nand U273 (N_273,In_299,In_402);
or U274 (N_274,N_85,N_113);
and U275 (N_275,In_209,In_414);
or U276 (N_276,In_205,N_166);
and U277 (N_277,In_110,In_273);
and U278 (N_278,In_29,N_178);
or U279 (N_279,In_329,N_197);
nor U280 (N_280,In_271,In_116);
or U281 (N_281,In_493,In_318);
and U282 (N_282,In_499,In_281);
or U283 (N_283,N_6,In_260);
nor U284 (N_284,N_65,N_176);
xor U285 (N_285,In_350,In_248);
and U286 (N_286,In_434,In_75);
and U287 (N_287,N_146,In_70);
nand U288 (N_288,In_489,N_67);
or U289 (N_289,N_185,In_123);
and U290 (N_290,In_455,N_31);
nor U291 (N_291,In_117,In_172);
nor U292 (N_292,In_87,In_58);
and U293 (N_293,In_457,N_81);
nand U294 (N_294,In_287,In_212);
nor U295 (N_295,In_474,N_182);
or U296 (N_296,In_484,In_262);
or U297 (N_297,In_185,In_186);
xnor U298 (N_298,N_92,N_192);
and U299 (N_299,In_398,N_130);
xnor U300 (N_300,N_184,In_114);
nor U301 (N_301,N_278,In_412);
or U302 (N_302,N_108,In_36);
nand U303 (N_303,In_460,In_175);
or U304 (N_304,N_206,N_223);
nand U305 (N_305,N_286,In_441);
nor U306 (N_306,In_90,N_273);
or U307 (N_307,In_134,N_64);
and U308 (N_308,N_282,N_230);
and U309 (N_309,In_465,N_98);
nor U310 (N_310,N_159,N_288);
and U311 (N_311,N_260,N_267);
nand U312 (N_312,In_11,N_117);
nand U313 (N_313,N_216,N_276);
xnor U314 (N_314,N_214,N_243);
and U315 (N_315,In_124,In_308);
nor U316 (N_316,N_148,N_266);
and U317 (N_317,N_43,In_498);
or U318 (N_318,N_190,N_39);
or U319 (N_319,N_18,In_144);
nand U320 (N_320,N_128,N_250);
or U321 (N_321,N_120,N_238);
nand U322 (N_322,N_256,N_283);
or U323 (N_323,N_122,N_163);
nor U324 (N_324,N_261,N_61);
and U325 (N_325,N_246,N_295);
nor U326 (N_326,N_268,N_251);
xor U327 (N_327,N_235,In_307);
and U328 (N_328,In_133,N_270);
xnor U329 (N_329,In_67,In_401);
nor U330 (N_330,N_158,N_293);
nor U331 (N_331,In_132,N_247);
xnor U332 (N_332,N_125,N_209);
nor U333 (N_333,N_269,N_285);
nand U334 (N_334,N_258,N_248);
nand U335 (N_335,N_289,N_133);
nand U336 (N_336,N_277,N_265);
or U337 (N_337,N_229,N_292);
and U338 (N_338,In_375,N_208);
or U339 (N_339,N_263,N_165);
or U340 (N_340,N_240,In_155);
nand U341 (N_341,N_217,N_106);
or U342 (N_342,N_225,N_255);
nor U343 (N_343,N_79,N_239);
nor U344 (N_344,N_101,N_284);
nor U345 (N_345,N_221,N_219);
nor U346 (N_346,N_234,N_299);
nor U347 (N_347,N_204,N_203);
xor U348 (N_348,N_233,N_257);
nand U349 (N_349,N_237,N_224);
nor U350 (N_350,N_259,N_241);
and U351 (N_351,N_167,N_26);
nor U352 (N_352,N_271,In_372);
or U353 (N_353,N_281,N_201);
nor U354 (N_354,N_152,In_470);
and U355 (N_355,N_191,N_231);
or U356 (N_356,N_40,In_236);
nor U357 (N_357,N_198,N_296);
nor U358 (N_358,N_88,In_218);
and U359 (N_359,In_164,N_274);
nand U360 (N_360,N_138,N_202);
nand U361 (N_361,In_476,N_210);
or U362 (N_362,In_334,N_161);
nor U363 (N_363,N_215,N_244);
or U364 (N_364,N_173,N_232);
or U365 (N_365,N_252,In_313);
and U366 (N_366,N_264,N_24);
and U367 (N_367,In_237,In_293);
nor U368 (N_368,In_478,In_394);
and U369 (N_369,N_132,N_279);
and U370 (N_370,N_213,N_194);
xnor U371 (N_371,N_220,N_228);
nor U372 (N_372,N_245,N_181);
nand U373 (N_373,In_119,In_107);
nand U374 (N_374,In_84,In_94);
nand U375 (N_375,In_120,N_14);
nor U376 (N_376,In_469,In_43);
and U377 (N_377,N_275,N_48);
nand U378 (N_378,N_226,N_297);
or U379 (N_379,N_253,N_272);
and U380 (N_380,N_139,N_157);
nor U381 (N_381,N_242,N_205);
and U382 (N_382,In_4,N_249);
or U383 (N_383,In_203,N_123);
and U384 (N_384,N_298,N_87);
or U385 (N_385,N_149,N_105);
and U386 (N_386,N_287,N_20);
nand U387 (N_387,In_250,N_262);
and U388 (N_388,N_212,N_254);
and U389 (N_389,N_290,N_280);
xnor U390 (N_390,N_207,N_294);
or U391 (N_391,N_112,In_74);
and U392 (N_392,N_227,N_155);
or U393 (N_393,N_116,In_6);
or U394 (N_394,N_78,N_222);
and U395 (N_395,N_124,N_211);
or U396 (N_396,N_131,In_80);
nor U397 (N_397,In_301,N_236);
xor U398 (N_398,N_72,N_200);
nor U399 (N_399,N_218,N_291);
nand U400 (N_400,N_337,N_386);
nor U401 (N_401,N_302,N_366);
nand U402 (N_402,N_398,N_340);
nand U403 (N_403,N_385,N_376);
or U404 (N_404,N_322,N_304);
xor U405 (N_405,N_362,N_348);
nand U406 (N_406,N_381,N_359);
and U407 (N_407,N_300,N_389);
nor U408 (N_408,N_368,N_338);
nor U409 (N_409,N_339,N_330);
nor U410 (N_410,N_328,N_383);
or U411 (N_411,N_341,N_352);
and U412 (N_412,N_369,N_346);
nand U413 (N_413,N_391,N_353);
nand U414 (N_414,N_344,N_354);
and U415 (N_415,N_397,N_335);
or U416 (N_416,N_367,N_313);
and U417 (N_417,N_351,N_311);
and U418 (N_418,N_331,N_342);
nor U419 (N_419,N_334,N_380);
nor U420 (N_420,N_306,N_303);
nor U421 (N_421,N_378,N_355);
nand U422 (N_422,N_357,N_319);
xor U423 (N_423,N_301,N_360);
and U424 (N_424,N_326,N_379);
xor U425 (N_425,N_307,N_375);
or U426 (N_426,N_324,N_382);
nor U427 (N_427,N_387,N_321);
and U428 (N_428,N_377,N_361);
nor U429 (N_429,N_388,N_316);
nor U430 (N_430,N_323,N_315);
and U431 (N_431,N_333,N_394);
and U432 (N_432,N_374,N_372);
nor U433 (N_433,N_371,N_325);
and U434 (N_434,N_309,N_358);
and U435 (N_435,N_347,N_308);
or U436 (N_436,N_317,N_392);
xnor U437 (N_437,N_350,N_332);
or U438 (N_438,N_336,N_393);
and U439 (N_439,N_314,N_390);
and U440 (N_440,N_305,N_370);
nand U441 (N_441,N_310,N_364);
or U442 (N_442,N_399,N_320);
nor U443 (N_443,N_329,N_343);
or U444 (N_444,N_365,N_312);
and U445 (N_445,N_373,N_349);
and U446 (N_446,N_363,N_384);
nor U447 (N_447,N_356,N_395);
nand U448 (N_448,N_318,N_327);
and U449 (N_449,N_345,N_396);
or U450 (N_450,N_320,N_377);
and U451 (N_451,N_305,N_325);
nand U452 (N_452,N_301,N_325);
nor U453 (N_453,N_315,N_376);
or U454 (N_454,N_340,N_374);
and U455 (N_455,N_391,N_379);
and U456 (N_456,N_357,N_327);
nor U457 (N_457,N_342,N_318);
or U458 (N_458,N_397,N_364);
or U459 (N_459,N_311,N_390);
nor U460 (N_460,N_381,N_317);
and U461 (N_461,N_379,N_389);
and U462 (N_462,N_397,N_372);
nand U463 (N_463,N_380,N_359);
nor U464 (N_464,N_322,N_312);
nand U465 (N_465,N_380,N_326);
nand U466 (N_466,N_313,N_396);
nand U467 (N_467,N_306,N_374);
or U468 (N_468,N_389,N_370);
nand U469 (N_469,N_397,N_373);
nor U470 (N_470,N_303,N_327);
nand U471 (N_471,N_301,N_365);
or U472 (N_472,N_334,N_336);
and U473 (N_473,N_393,N_337);
nand U474 (N_474,N_304,N_376);
and U475 (N_475,N_334,N_325);
and U476 (N_476,N_330,N_341);
and U477 (N_477,N_340,N_323);
or U478 (N_478,N_356,N_344);
xnor U479 (N_479,N_361,N_317);
nor U480 (N_480,N_378,N_309);
nand U481 (N_481,N_395,N_368);
or U482 (N_482,N_349,N_372);
nand U483 (N_483,N_373,N_353);
and U484 (N_484,N_364,N_328);
or U485 (N_485,N_386,N_338);
and U486 (N_486,N_302,N_340);
nand U487 (N_487,N_353,N_300);
xor U488 (N_488,N_345,N_355);
or U489 (N_489,N_337,N_334);
nand U490 (N_490,N_358,N_323);
nor U491 (N_491,N_314,N_312);
or U492 (N_492,N_326,N_368);
nand U493 (N_493,N_370,N_313);
or U494 (N_494,N_371,N_351);
nor U495 (N_495,N_370,N_316);
nand U496 (N_496,N_374,N_322);
nor U497 (N_497,N_312,N_338);
xnor U498 (N_498,N_387,N_319);
and U499 (N_499,N_310,N_352);
or U500 (N_500,N_416,N_421);
nor U501 (N_501,N_493,N_490);
or U502 (N_502,N_457,N_473);
nand U503 (N_503,N_417,N_412);
nor U504 (N_504,N_449,N_411);
or U505 (N_505,N_480,N_440);
nor U506 (N_506,N_443,N_483);
and U507 (N_507,N_409,N_407);
or U508 (N_508,N_438,N_430);
or U509 (N_509,N_460,N_425);
nand U510 (N_510,N_435,N_445);
or U511 (N_511,N_496,N_437);
nor U512 (N_512,N_414,N_424);
and U513 (N_513,N_419,N_422);
and U514 (N_514,N_415,N_406);
or U515 (N_515,N_461,N_476);
nor U516 (N_516,N_497,N_469);
nand U517 (N_517,N_441,N_475);
nor U518 (N_518,N_465,N_456);
nand U519 (N_519,N_439,N_484);
nor U520 (N_520,N_436,N_482);
xnor U521 (N_521,N_431,N_413);
nand U522 (N_522,N_472,N_471);
xnor U523 (N_523,N_454,N_481);
or U524 (N_524,N_494,N_492);
nand U525 (N_525,N_426,N_423);
and U526 (N_526,N_448,N_455);
and U527 (N_527,N_446,N_451);
or U528 (N_528,N_433,N_459);
or U529 (N_529,N_401,N_427);
or U530 (N_530,N_478,N_485);
nand U531 (N_531,N_467,N_402);
nor U532 (N_532,N_453,N_466);
and U533 (N_533,N_450,N_452);
and U534 (N_534,N_486,N_489);
nand U535 (N_535,N_434,N_404);
and U536 (N_536,N_420,N_491);
nor U537 (N_537,N_499,N_408);
or U538 (N_538,N_410,N_495);
nand U539 (N_539,N_463,N_470);
xnor U540 (N_540,N_458,N_428);
nor U541 (N_541,N_488,N_468);
nor U542 (N_542,N_498,N_462);
or U543 (N_543,N_447,N_464);
and U544 (N_544,N_400,N_405);
or U545 (N_545,N_444,N_432);
or U546 (N_546,N_418,N_479);
or U547 (N_547,N_442,N_477);
and U548 (N_548,N_487,N_474);
xor U549 (N_549,N_429,N_403);
or U550 (N_550,N_477,N_438);
nand U551 (N_551,N_478,N_421);
nand U552 (N_552,N_441,N_469);
nand U553 (N_553,N_481,N_475);
or U554 (N_554,N_422,N_416);
and U555 (N_555,N_408,N_439);
and U556 (N_556,N_427,N_456);
and U557 (N_557,N_449,N_448);
and U558 (N_558,N_484,N_453);
nor U559 (N_559,N_400,N_418);
or U560 (N_560,N_481,N_484);
nand U561 (N_561,N_492,N_470);
or U562 (N_562,N_431,N_434);
nor U563 (N_563,N_495,N_403);
and U564 (N_564,N_405,N_453);
nor U565 (N_565,N_482,N_416);
and U566 (N_566,N_430,N_496);
nand U567 (N_567,N_498,N_405);
or U568 (N_568,N_423,N_412);
or U569 (N_569,N_428,N_478);
xnor U570 (N_570,N_477,N_453);
or U571 (N_571,N_414,N_435);
and U572 (N_572,N_400,N_440);
nand U573 (N_573,N_445,N_461);
xnor U574 (N_574,N_469,N_468);
or U575 (N_575,N_431,N_455);
nor U576 (N_576,N_407,N_440);
xor U577 (N_577,N_479,N_441);
or U578 (N_578,N_494,N_470);
and U579 (N_579,N_436,N_457);
xor U580 (N_580,N_405,N_496);
nand U581 (N_581,N_495,N_416);
nor U582 (N_582,N_489,N_467);
or U583 (N_583,N_458,N_452);
xor U584 (N_584,N_424,N_448);
or U585 (N_585,N_433,N_403);
or U586 (N_586,N_456,N_499);
or U587 (N_587,N_439,N_444);
and U588 (N_588,N_477,N_411);
and U589 (N_589,N_432,N_408);
xnor U590 (N_590,N_401,N_467);
nor U591 (N_591,N_461,N_482);
and U592 (N_592,N_470,N_448);
nor U593 (N_593,N_427,N_485);
or U594 (N_594,N_435,N_449);
nand U595 (N_595,N_482,N_447);
nor U596 (N_596,N_489,N_457);
xor U597 (N_597,N_459,N_418);
nor U598 (N_598,N_491,N_490);
nor U599 (N_599,N_420,N_430);
and U600 (N_600,N_503,N_588);
and U601 (N_601,N_529,N_551);
or U602 (N_602,N_598,N_575);
and U603 (N_603,N_557,N_550);
nand U604 (N_604,N_591,N_534);
nor U605 (N_605,N_538,N_524);
nand U606 (N_606,N_585,N_543);
nor U607 (N_607,N_514,N_589);
nand U608 (N_608,N_577,N_531);
nand U609 (N_609,N_549,N_581);
or U610 (N_610,N_513,N_546);
nor U611 (N_611,N_592,N_528);
and U612 (N_612,N_521,N_535);
nor U613 (N_613,N_593,N_516);
and U614 (N_614,N_515,N_584);
nand U615 (N_615,N_530,N_556);
nand U616 (N_616,N_506,N_509);
nor U617 (N_617,N_502,N_560);
or U618 (N_618,N_508,N_523);
xnor U619 (N_619,N_568,N_547);
nor U620 (N_620,N_561,N_555);
or U621 (N_621,N_512,N_563);
or U622 (N_622,N_590,N_500);
and U623 (N_623,N_587,N_537);
or U624 (N_624,N_522,N_505);
nand U625 (N_625,N_595,N_596);
nor U626 (N_626,N_544,N_566);
nand U627 (N_627,N_541,N_526);
nand U628 (N_628,N_578,N_539);
nor U629 (N_629,N_507,N_552);
nor U630 (N_630,N_586,N_582);
nand U631 (N_631,N_519,N_510);
or U632 (N_632,N_583,N_517);
or U633 (N_633,N_569,N_574);
and U634 (N_634,N_518,N_548);
nor U635 (N_635,N_553,N_545);
nand U636 (N_636,N_536,N_562);
xnor U637 (N_637,N_597,N_511);
or U638 (N_638,N_501,N_564);
and U639 (N_639,N_599,N_565);
or U640 (N_640,N_504,N_542);
nand U641 (N_641,N_559,N_525);
and U642 (N_642,N_540,N_572);
xor U643 (N_643,N_554,N_558);
and U644 (N_644,N_520,N_594);
xnor U645 (N_645,N_573,N_571);
or U646 (N_646,N_532,N_579);
nor U647 (N_647,N_580,N_570);
nand U648 (N_648,N_576,N_527);
xor U649 (N_649,N_533,N_567);
nor U650 (N_650,N_560,N_551);
nand U651 (N_651,N_537,N_512);
nor U652 (N_652,N_560,N_596);
nand U653 (N_653,N_501,N_550);
or U654 (N_654,N_543,N_533);
nand U655 (N_655,N_518,N_574);
nand U656 (N_656,N_593,N_563);
xor U657 (N_657,N_591,N_533);
nand U658 (N_658,N_501,N_543);
nor U659 (N_659,N_531,N_515);
nor U660 (N_660,N_598,N_502);
nor U661 (N_661,N_544,N_551);
nor U662 (N_662,N_516,N_562);
nor U663 (N_663,N_544,N_543);
or U664 (N_664,N_599,N_549);
nand U665 (N_665,N_553,N_523);
xor U666 (N_666,N_580,N_514);
or U667 (N_667,N_510,N_505);
nand U668 (N_668,N_568,N_558);
and U669 (N_669,N_520,N_500);
nand U670 (N_670,N_569,N_553);
nand U671 (N_671,N_586,N_517);
and U672 (N_672,N_560,N_575);
or U673 (N_673,N_569,N_513);
and U674 (N_674,N_598,N_557);
xnor U675 (N_675,N_584,N_588);
nor U676 (N_676,N_539,N_590);
and U677 (N_677,N_578,N_536);
or U678 (N_678,N_510,N_541);
or U679 (N_679,N_568,N_575);
and U680 (N_680,N_595,N_502);
or U681 (N_681,N_535,N_572);
and U682 (N_682,N_514,N_537);
nor U683 (N_683,N_523,N_591);
nor U684 (N_684,N_518,N_565);
or U685 (N_685,N_584,N_560);
xor U686 (N_686,N_553,N_562);
and U687 (N_687,N_578,N_526);
nor U688 (N_688,N_599,N_531);
nand U689 (N_689,N_521,N_578);
or U690 (N_690,N_599,N_553);
nand U691 (N_691,N_526,N_581);
nor U692 (N_692,N_550,N_525);
and U693 (N_693,N_592,N_569);
nor U694 (N_694,N_583,N_553);
nor U695 (N_695,N_514,N_567);
nand U696 (N_696,N_564,N_516);
nand U697 (N_697,N_532,N_593);
or U698 (N_698,N_559,N_530);
and U699 (N_699,N_579,N_521);
nand U700 (N_700,N_682,N_678);
or U701 (N_701,N_631,N_694);
nor U702 (N_702,N_632,N_606);
and U703 (N_703,N_675,N_644);
nand U704 (N_704,N_600,N_635);
and U705 (N_705,N_671,N_690);
xnor U706 (N_706,N_610,N_612);
or U707 (N_707,N_699,N_611);
nor U708 (N_708,N_657,N_615);
nand U709 (N_709,N_654,N_687);
nor U710 (N_710,N_688,N_608);
and U711 (N_711,N_604,N_627);
nor U712 (N_712,N_695,N_652);
xnor U713 (N_713,N_693,N_669);
nand U714 (N_714,N_637,N_645);
nand U715 (N_715,N_666,N_689);
or U716 (N_716,N_629,N_665);
and U717 (N_717,N_619,N_674);
and U718 (N_718,N_681,N_642);
or U719 (N_719,N_684,N_698);
and U720 (N_720,N_651,N_685);
nor U721 (N_721,N_618,N_603);
nor U722 (N_722,N_686,N_659);
xor U723 (N_723,N_664,N_607);
or U724 (N_724,N_647,N_670);
nor U725 (N_725,N_653,N_672);
or U726 (N_726,N_683,N_648);
nand U727 (N_727,N_623,N_660);
nand U728 (N_728,N_677,N_697);
nand U729 (N_729,N_620,N_609);
nor U730 (N_730,N_668,N_667);
or U731 (N_731,N_601,N_602);
or U732 (N_732,N_673,N_630);
nor U733 (N_733,N_658,N_661);
and U734 (N_734,N_626,N_621);
and U735 (N_735,N_633,N_641);
nand U736 (N_736,N_656,N_616);
nor U737 (N_737,N_691,N_696);
or U738 (N_738,N_624,N_663);
or U739 (N_739,N_617,N_622);
nor U740 (N_740,N_662,N_649);
nor U741 (N_741,N_643,N_655);
and U742 (N_742,N_634,N_605);
nor U743 (N_743,N_650,N_640);
or U744 (N_744,N_614,N_628);
nand U745 (N_745,N_679,N_638);
nor U746 (N_746,N_676,N_680);
nor U747 (N_747,N_613,N_636);
and U748 (N_748,N_639,N_692);
or U749 (N_749,N_646,N_625);
nand U750 (N_750,N_674,N_656);
or U751 (N_751,N_662,N_617);
nor U752 (N_752,N_659,N_646);
nor U753 (N_753,N_692,N_632);
or U754 (N_754,N_606,N_646);
and U755 (N_755,N_691,N_609);
and U756 (N_756,N_697,N_601);
or U757 (N_757,N_658,N_698);
nor U758 (N_758,N_616,N_648);
or U759 (N_759,N_613,N_667);
nor U760 (N_760,N_669,N_664);
nand U761 (N_761,N_649,N_601);
or U762 (N_762,N_610,N_678);
or U763 (N_763,N_618,N_694);
nand U764 (N_764,N_665,N_679);
nand U765 (N_765,N_655,N_698);
or U766 (N_766,N_615,N_678);
nand U767 (N_767,N_661,N_641);
xor U768 (N_768,N_619,N_653);
or U769 (N_769,N_626,N_699);
nand U770 (N_770,N_616,N_659);
nand U771 (N_771,N_662,N_646);
or U772 (N_772,N_668,N_662);
nor U773 (N_773,N_677,N_633);
and U774 (N_774,N_618,N_620);
xor U775 (N_775,N_658,N_696);
and U776 (N_776,N_657,N_645);
nor U777 (N_777,N_682,N_631);
or U778 (N_778,N_695,N_640);
or U779 (N_779,N_664,N_662);
nand U780 (N_780,N_629,N_623);
or U781 (N_781,N_653,N_658);
nor U782 (N_782,N_679,N_600);
nand U783 (N_783,N_656,N_641);
or U784 (N_784,N_607,N_639);
nand U785 (N_785,N_685,N_693);
nand U786 (N_786,N_652,N_662);
nand U787 (N_787,N_679,N_690);
and U788 (N_788,N_689,N_643);
or U789 (N_789,N_601,N_655);
nor U790 (N_790,N_632,N_681);
nor U791 (N_791,N_690,N_657);
nor U792 (N_792,N_695,N_687);
and U793 (N_793,N_612,N_649);
xor U794 (N_794,N_629,N_637);
nand U795 (N_795,N_642,N_663);
or U796 (N_796,N_611,N_686);
and U797 (N_797,N_611,N_637);
xor U798 (N_798,N_601,N_613);
or U799 (N_799,N_616,N_638);
or U800 (N_800,N_775,N_700);
or U801 (N_801,N_759,N_762);
nand U802 (N_802,N_745,N_728);
nor U803 (N_803,N_704,N_743);
nor U804 (N_804,N_781,N_777);
xnor U805 (N_805,N_715,N_722);
xor U806 (N_806,N_731,N_721);
and U807 (N_807,N_784,N_751);
or U808 (N_808,N_770,N_787);
nor U809 (N_809,N_718,N_771);
and U810 (N_810,N_720,N_705);
nor U811 (N_811,N_779,N_795);
xnor U812 (N_812,N_736,N_729);
or U813 (N_813,N_707,N_740);
and U814 (N_814,N_794,N_766);
xor U815 (N_815,N_725,N_765);
xor U816 (N_816,N_796,N_789);
nor U817 (N_817,N_760,N_755);
nor U818 (N_818,N_733,N_747);
or U819 (N_819,N_746,N_773);
nand U820 (N_820,N_742,N_793);
or U821 (N_821,N_719,N_782);
nor U822 (N_822,N_769,N_726);
nor U823 (N_823,N_797,N_753);
or U824 (N_824,N_788,N_708);
and U825 (N_825,N_735,N_799);
nand U826 (N_826,N_774,N_709);
or U827 (N_827,N_778,N_786);
or U828 (N_828,N_752,N_717);
or U829 (N_829,N_714,N_750);
and U830 (N_830,N_702,N_744);
and U831 (N_831,N_757,N_772);
nor U832 (N_832,N_706,N_754);
and U833 (N_833,N_734,N_756);
xnor U834 (N_834,N_785,N_703);
nor U835 (N_835,N_780,N_701);
and U836 (N_836,N_723,N_791);
nand U837 (N_837,N_749,N_738);
or U838 (N_838,N_716,N_798);
nand U839 (N_839,N_712,N_748);
or U840 (N_840,N_724,N_730);
or U841 (N_841,N_713,N_739);
and U842 (N_842,N_758,N_732);
or U843 (N_843,N_727,N_737);
nand U844 (N_844,N_761,N_792);
and U845 (N_845,N_767,N_783);
and U846 (N_846,N_768,N_790);
nor U847 (N_847,N_764,N_776);
nand U848 (N_848,N_711,N_741);
and U849 (N_849,N_763,N_710);
and U850 (N_850,N_787,N_703);
and U851 (N_851,N_738,N_752);
nand U852 (N_852,N_727,N_703);
or U853 (N_853,N_798,N_735);
or U854 (N_854,N_767,N_745);
nand U855 (N_855,N_711,N_709);
and U856 (N_856,N_747,N_798);
nor U857 (N_857,N_750,N_732);
nor U858 (N_858,N_781,N_748);
and U859 (N_859,N_735,N_705);
xor U860 (N_860,N_747,N_706);
nand U861 (N_861,N_791,N_744);
nor U862 (N_862,N_731,N_730);
or U863 (N_863,N_788,N_737);
or U864 (N_864,N_720,N_789);
nor U865 (N_865,N_717,N_720);
and U866 (N_866,N_715,N_777);
nand U867 (N_867,N_714,N_791);
or U868 (N_868,N_747,N_758);
nor U869 (N_869,N_722,N_754);
and U870 (N_870,N_732,N_792);
or U871 (N_871,N_788,N_760);
or U872 (N_872,N_701,N_715);
and U873 (N_873,N_740,N_724);
or U874 (N_874,N_711,N_730);
nor U875 (N_875,N_785,N_750);
nand U876 (N_876,N_752,N_780);
xor U877 (N_877,N_778,N_726);
nand U878 (N_878,N_774,N_782);
and U879 (N_879,N_742,N_772);
xnor U880 (N_880,N_719,N_743);
nor U881 (N_881,N_727,N_740);
nand U882 (N_882,N_760,N_797);
and U883 (N_883,N_747,N_742);
nand U884 (N_884,N_770,N_767);
nand U885 (N_885,N_753,N_751);
and U886 (N_886,N_713,N_733);
nand U887 (N_887,N_701,N_750);
and U888 (N_888,N_761,N_726);
nand U889 (N_889,N_762,N_736);
xor U890 (N_890,N_773,N_705);
or U891 (N_891,N_720,N_777);
nor U892 (N_892,N_748,N_754);
nand U893 (N_893,N_730,N_773);
nand U894 (N_894,N_790,N_782);
or U895 (N_895,N_753,N_756);
nand U896 (N_896,N_776,N_772);
nor U897 (N_897,N_754,N_771);
nor U898 (N_898,N_713,N_756);
and U899 (N_899,N_794,N_733);
nor U900 (N_900,N_884,N_861);
nor U901 (N_901,N_857,N_818);
nand U902 (N_902,N_888,N_865);
nand U903 (N_903,N_826,N_845);
or U904 (N_904,N_870,N_854);
nand U905 (N_905,N_809,N_886);
and U906 (N_906,N_874,N_868);
xor U907 (N_907,N_820,N_898);
nand U908 (N_908,N_863,N_877);
and U909 (N_909,N_840,N_895);
nand U910 (N_910,N_838,N_890);
nand U911 (N_911,N_880,N_829);
and U912 (N_912,N_833,N_849);
and U913 (N_913,N_813,N_896);
or U914 (N_914,N_876,N_827);
and U915 (N_915,N_819,N_816);
or U916 (N_916,N_893,N_891);
xor U917 (N_917,N_843,N_897);
and U918 (N_918,N_878,N_839);
or U919 (N_919,N_814,N_872);
nand U920 (N_920,N_882,N_899);
and U921 (N_921,N_864,N_817);
nor U922 (N_922,N_873,N_851);
or U923 (N_923,N_804,N_837);
nor U924 (N_924,N_894,N_822);
nor U925 (N_925,N_834,N_889);
nand U926 (N_926,N_832,N_805);
nor U927 (N_927,N_831,N_847);
and U928 (N_928,N_836,N_811);
nand U929 (N_929,N_823,N_828);
and U930 (N_930,N_867,N_846);
and U931 (N_931,N_835,N_879);
nand U932 (N_932,N_800,N_860);
nor U933 (N_933,N_869,N_866);
or U934 (N_934,N_887,N_844);
xor U935 (N_935,N_808,N_815);
or U936 (N_936,N_802,N_853);
nand U937 (N_937,N_855,N_824);
or U938 (N_938,N_856,N_862);
or U939 (N_939,N_883,N_830);
or U940 (N_940,N_842,N_875);
or U941 (N_941,N_806,N_825);
and U942 (N_942,N_807,N_848);
nor U943 (N_943,N_810,N_812);
nor U944 (N_944,N_841,N_858);
nor U945 (N_945,N_852,N_801);
and U946 (N_946,N_871,N_892);
nand U947 (N_947,N_821,N_859);
nand U948 (N_948,N_850,N_885);
nor U949 (N_949,N_881,N_803);
and U950 (N_950,N_899,N_865);
or U951 (N_951,N_821,N_896);
nor U952 (N_952,N_894,N_875);
or U953 (N_953,N_855,N_801);
nand U954 (N_954,N_811,N_829);
or U955 (N_955,N_816,N_817);
and U956 (N_956,N_822,N_833);
nand U957 (N_957,N_852,N_822);
nand U958 (N_958,N_836,N_883);
nand U959 (N_959,N_849,N_834);
or U960 (N_960,N_827,N_854);
nand U961 (N_961,N_847,N_888);
nor U962 (N_962,N_859,N_869);
or U963 (N_963,N_892,N_836);
nand U964 (N_964,N_873,N_871);
nor U965 (N_965,N_864,N_859);
nor U966 (N_966,N_832,N_878);
and U967 (N_967,N_852,N_854);
nand U968 (N_968,N_860,N_833);
and U969 (N_969,N_858,N_880);
or U970 (N_970,N_843,N_873);
and U971 (N_971,N_860,N_842);
nor U972 (N_972,N_875,N_883);
nor U973 (N_973,N_807,N_861);
or U974 (N_974,N_862,N_806);
nand U975 (N_975,N_844,N_820);
nor U976 (N_976,N_888,N_816);
nand U977 (N_977,N_826,N_807);
and U978 (N_978,N_846,N_884);
nor U979 (N_979,N_832,N_807);
nor U980 (N_980,N_800,N_809);
nand U981 (N_981,N_879,N_807);
nand U982 (N_982,N_849,N_869);
or U983 (N_983,N_897,N_887);
nor U984 (N_984,N_826,N_828);
or U985 (N_985,N_839,N_888);
nor U986 (N_986,N_822,N_883);
nand U987 (N_987,N_838,N_893);
nand U988 (N_988,N_839,N_821);
or U989 (N_989,N_864,N_814);
nor U990 (N_990,N_888,N_836);
nand U991 (N_991,N_884,N_818);
nand U992 (N_992,N_803,N_897);
or U993 (N_993,N_899,N_831);
and U994 (N_994,N_832,N_829);
nand U995 (N_995,N_869,N_838);
or U996 (N_996,N_873,N_801);
or U997 (N_997,N_863,N_811);
and U998 (N_998,N_813,N_872);
nand U999 (N_999,N_811,N_850);
and U1000 (N_1000,N_980,N_905);
or U1001 (N_1001,N_940,N_929);
and U1002 (N_1002,N_908,N_914);
nand U1003 (N_1003,N_995,N_974);
nand U1004 (N_1004,N_987,N_966);
nor U1005 (N_1005,N_918,N_967);
or U1006 (N_1006,N_975,N_941);
nand U1007 (N_1007,N_931,N_973);
or U1008 (N_1008,N_962,N_997);
and U1009 (N_1009,N_937,N_935);
xnor U1010 (N_1010,N_994,N_954);
nand U1011 (N_1011,N_988,N_950);
nor U1012 (N_1012,N_989,N_923);
nand U1013 (N_1013,N_900,N_920);
and U1014 (N_1014,N_993,N_917);
or U1015 (N_1015,N_983,N_964);
nor U1016 (N_1016,N_985,N_965);
xor U1017 (N_1017,N_927,N_909);
or U1018 (N_1018,N_957,N_932);
nor U1019 (N_1019,N_960,N_919);
xnor U1020 (N_1020,N_952,N_991);
nor U1021 (N_1021,N_968,N_948);
or U1022 (N_1022,N_958,N_947);
xor U1023 (N_1023,N_970,N_911);
nor U1024 (N_1024,N_933,N_930);
and U1025 (N_1025,N_953,N_907);
nor U1026 (N_1026,N_976,N_972);
xnor U1027 (N_1027,N_934,N_912);
xor U1028 (N_1028,N_906,N_910);
or U1029 (N_1029,N_949,N_903);
nand U1030 (N_1030,N_926,N_943);
nand U1031 (N_1031,N_981,N_963);
and U1032 (N_1032,N_938,N_986);
nor U1033 (N_1033,N_925,N_915);
nand U1034 (N_1034,N_971,N_955);
nor U1035 (N_1035,N_902,N_921);
nand U1036 (N_1036,N_944,N_945);
nand U1037 (N_1037,N_942,N_951);
or U1038 (N_1038,N_924,N_984);
and U1039 (N_1039,N_999,N_946);
nand U1040 (N_1040,N_913,N_901);
and U1041 (N_1041,N_961,N_922);
nor U1042 (N_1042,N_969,N_977);
nand U1043 (N_1043,N_916,N_956);
nor U1044 (N_1044,N_928,N_936);
and U1045 (N_1045,N_996,N_982);
nor U1046 (N_1046,N_979,N_959);
nand U1047 (N_1047,N_904,N_998);
and U1048 (N_1048,N_992,N_978);
and U1049 (N_1049,N_990,N_939);
xnor U1050 (N_1050,N_976,N_951);
nand U1051 (N_1051,N_995,N_987);
nor U1052 (N_1052,N_984,N_985);
nand U1053 (N_1053,N_929,N_956);
or U1054 (N_1054,N_907,N_964);
or U1055 (N_1055,N_935,N_913);
nor U1056 (N_1056,N_998,N_926);
xnor U1057 (N_1057,N_945,N_961);
nand U1058 (N_1058,N_988,N_948);
or U1059 (N_1059,N_945,N_994);
and U1060 (N_1060,N_997,N_986);
or U1061 (N_1061,N_907,N_906);
nand U1062 (N_1062,N_974,N_964);
nor U1063 (N_1063,N_903,N_967);
nor U1064 (N_1064,N_900,N_978);
or U1065 (N_1065,N_997,N_991);
and U1066 (N_1066,N_961,N_973);
and U1067 (N_1067,N_924,N_949);
nor U1068 (N_1068,N_918,N_902);
nor U1069 (N_1069,N_963,N_923);
nand U1070 (N_1070,N_953,N_920);
and U1071 (N_1071,N_901,N_998);
or U1072 (N_1072,N_957,N_900);
nor U1073 (N_1073,N_990,N_993);
nand U1074 (N_1074,N_906,N_984);
nor U1075 (N_1075,N_955,N_993);
or U1076 (N_1076,N_914,N_946);
nor U1077 (N_1077,N_966,N_917);
or U1078 (N_1078,N_914,N_966);
xnor U1079 (N_1079,N_997,N_938);
and U1080 (N_1080,N_977,N_966);
xnor U1081 (N_1081,N_995,N_958);
or U1082 (N_1082,N_923,N_926);
nor U1083 (N_1083,N_972,N_984);
or U1084 (N_1084,N_910,N_970);
xor U1085 (N_1085,N_942,N_908);
xnor U1086 (N_1086,N_914,N_944);
or U1087 (N_1087,N_982,N_986);
nor U1088 (N_1088,N_961,N_996);
and U1089 (N_1089,N_953,N_952);
or U1090 (N_1090,N_982,N_944);
nand U1091 (N_1091,N_991,N_994);
and U1092 (N_1092,N_906,N_991);
and U1093 (N_1093,N_986,N_919);
and U1094 (N_1094,N_973,N_997);
or U1095 (N_1095,N_922,N_964);
or U1096 (N_1096,N_950,N_977);
nand U1097 (N_1097,N_989,N_955);
or U1098 (N_1098,N_979,N_918);
nor U1099 (N_1099,N_986,N_995);
nor U1100 (N_1100,N_1040,N_1056);
and U1101 (N_1101,N_1081,N_1048);
nor U1102 (N_1102,N_1030,N_1044);
nand U1103 (N_1103,N_1071,N_1046);
nor U1104 (N_1104,N_1074,N_1073);
nand U1105 (N_1105,N_1057,N_1014);
nor U1106 (N_1106,N_1031,N_1008);
or U1107 (N_1107,N_1036,N_1099);
nor U1108 (N_1108,N_1017,N_1035);
nand U1109 (N_1109,N_1019,N_1083);
nor U1110 (N_1110,N_1095,N_1025);
nand U1111 (N_1111,N_1018,N_1043);
or U1112 (N_1112,N_1050,N_1010);
nand U1113 (N_1113,N_1086,N_1005);
nand U1114 (N_1114,N_1091,N_1027);
xnor U1115 (N_1115,N_1075,N_1067);
and U1116 (N_1116,N_1082,N_1060);
xnor U1117 (N_1117,N_1013,N_1049);
nor U1118 (N_1118,N_1023,N_1066);
nand U1119 (N_1119,N_1011,N_1068);
nand U1120 (N_1120,N_1058,N_1047);
nand U1121 (N_1121,N_1098,N_1032);
and U1122 (N_1122,N_1000,N_1015);
xnor U1123 (N_1123,N_1088,N_1096);
nand U1124 (N_1124,N_1092,N_1079);
nand U1125 (N_1125,N_1080,N_1042);
and U1126 (N_1126,N_1020,N_1072);
nand U1127 (N_1127,N_1002,N_1087);
nor U1128 (N_1128,N_1097,N_1029);
nor U1129 (N_1129,N_1053,N_1028);
nor U1130 (N_1130,N_1012,N_1007);
nand U1131 (N_1131,N_1004,N_1009);
and U1132 (N_1132,N_1033,N_1089);
or U1133 (N_1133,N_1078,N_1061);
nand U1134 (N_1134,N_1038,N_1026);
and U1135 (N_1135,N_1055,N_1070);
nor U1136 (N_1136,N_1041,N_1085);
and U1137 (N_1137,N_1084,N_1065);
and U1138 (N_1138,N_1016,N_1024);
and U1139 (N_1139,N_1034,N_1045);
nand U1140 (N_1140,N_1052,N_1062);
nand U1141 (N_1141,N_1069,N_1064);
or U1142 (N_1142,N_1039,N_1001);
nand U1143 (N_1143,N_1094,N_1077);
nor U1144 (N_1144,N_1093,N_1003);
nand U1145 (N_1145,N_1006,N_1076);
and U1146 (N_1146,N_1054,N_1059);
nor U1147 (N_1147,N_1037,N_1090);
and U1148 (N_1148,N_1021,N_1051);
nor U1149 (N_1149,N_1022,N_1063);
xor U1150 (N_1150,N_1079,N_1089);
nand U1151 (N_1151,N_1036,N_1025);
nor U1152 (N_1152,N_1014,N_1003);
xor U1153 (N_1153,N_1051,N_1047);
nor U1154 (N_1154,N_1014,N_1024);
or U1155 (N_1155,N_1084,N_1012);
nor U1156 (N_1156,N_1099,N_1016);
and U1157 (N_1157,N_1077,N_1084);
xor U1158 (N_1158,N_1049,N_1080);
nand U1159 (N_1159,N_1000,N_1018);
and U1160 (N_1160,N_1012,N_1091);
or U1161 (N_1161,N_1097,N_1062);
nor U1162 (N_1162,N_1026,N_1053);
nand U1163 (N_1163,N_1038,N_1034);
or U1164 (N_1164,N_1022,N_1010);
nand U1165 (N_1165,N_1083,N_1059);
nand U1166 (N_1166,N_1037,N_1073);
and U1167 (N_1167,N_1045,N_1017);
and U1168 (N_1168,N_1008,N_1032);
or U1169 (N_1169,N_1060,N_1023);
and U1170 (N_1170,N_1030,N_1016);
and U1171 (N_1171,N_1054,N_1066);
xnor U1172 (N_1172,N_1085,N_1082);
nor U1173 (N_1173,N_1049,N_1053);
nor U1174 (N_1174,N_1014,N_1017);
and U1175 (N_1175,N_1004,N_1072);
nor U1176 (N_1176,N_1060,N_1065);
nand U1177 (N_1177,N_1026,N_1030);
or U1178 (N_1178,N_1058,N_1090);
or U1179 (N_1179,N_1011,N_1086);
or U1180 (N_1180,N_1090,N_1025);
and U1181 (N_1181,N_1026,N_1089);
and U1182 (N_1182,N_1041,N_1012);
nand U1183 (N_1183,N_1025,N_1011);
xnor U1184 (N_1184,N_1047,N_1099);
nor U1185 (N_1185,N_1056,N_1041);
and U1186 (N_1186,N_1020,N_1044);
or U1187 (N_1187,N_1062,N_1036);
and U1188 (N_1188,N_1032,N_1076);
nor U1189 (N_1189,N_1091,N_1057);
or U1190 (N_1190,N_1032,N_1041);
nand U1191 (N_1191,N_1002,N_1008);
nor U1192 (N_1192,N_1048,N_1029);
and U1193 (N_1193,N_1013,N_1051);
nor U1194 (N_1194,N_1085,N_1029);
nor U1195 (N_1195,N_1028,N_1033);
nor U1196 (N_1196,N_1005,N_1068);
or U1197 (N_1197,N_1013,N_1085);
or U1198 (N_1198,N_1048,N_1014);
xor U1199 (N_1199,N_1072,N_1081);
or U1200 (N_1200,N_1172,N_1173);
and U1201 (N_1201,N_1102,N_1132);
nand U1202 (N_1202,N_1196,N_1142);
nand U1203 (N_1203,N_1101,N_1189);
nand U1204 (N_1204,N_1143,N_1195);
nor U1205 (N_1205,N_1169,N_1138);
and U1206 (N_1206,N_1119,N_1116);
or U1207 (N_1207,N_1135,N_1147);
nor U1208 (N_1208,N_1158,N_1183);
nand U1209 (N_1209,N_1171,N_1144);
nor U1210 (N_1210,N_1178,N_1176);
and U1211 (N_1211,N_1168,N_1145);
nor U1212 (N_1212,N_1124,N_1128);
or U1213 (N_1213,N_1167,N_1100);
nor U1214 (N_1214,N_1141,N_1161);
or U1215 (N_1215,N_1164,N_1174);
or U1216 (N_1216,N_1146,N_1193);
nor U1217 (N_1217,N_1184,N_1156);
or U1218 (N_1218,N_1104,N_1190);
or U1219 (N_1219,N_1151,N_1160);
xor U1220 (N_1220,N_1118,N_1154);
or U1221 (N_1221,N_1134,N_1136);
or U1222 (N_1222,N_1149,N_1111);
and U1223 (N_1223,N_1108,N_1163);
nor U1224 (N_1224,N_1105,N_1112);
nor U1225 (N_1225,N_1122,N_1129);
and U1226 (N_1226,N_1179,N_1137);
and U1227 (N_1227,N_1170,N_1107);
and U1228 (N_1228,N_1115,N_1114);
nand U1229 (N_1229,N_1166,N_1152);
nor U1230 (N_1230,N_1109,N_1191);
or U1231 (N_1231,N_1106,N_1188);
nor U1232 (N_1232,N_1157,N_1182);
xnor U1233 (N_1233,N_1186,N_1180);
xor U1234 (N_1234,N_1125,N_1197);
nor U1235 (N_1235,N_1199,N_1148);
or U1236 (N_1236,N_1110,N_1133);
nand U1237 (N_1237,N_1131,N_1181);
or U1238 (N_1238,N_1103,N_1130);
nand U1239 (N_1239,N_1159,N_1127);
and U1240 (N_1240,N_1187,N_1155);
nand U1241 (N_1241,N_1117,N_1162);
and U1242 (N_1242,N_1194,N_1126);
and U1243 (N_1243,N_1153,N_1165);
and U1244 (N_1244,N_1192,N_1113);
nor U1245 (N_1245,N_1121,N_1150);
nand U1246 (N_1246,N_1177,N_1140);
or U1247 (N_1247,N_1120,N_1139);
nand U1248 (N_1248,N_1185,N_1123);
nor U1249 (N_1249,N_1198,N_1175);
or U1250 (N_1250,N_1166,N_1117);
nor U1251 (N_1251,N_1160,N_1169);
nand U1252 (N_1252,N_1158,N_1175);
and U1253 (N_1253,N_1123,N_1130);
or U1254 (N_1254,N_1120,N_1141);
nor U1255 (N_1255,N_1110,N_1193);
xnor U1256 (N_1256,N_1113,N_1171);
nor U1257 (N_1257,N_1121,N_1188);
nor U1258 (N_1258,N_1166,N_1163);
nand U1259 (N_1259,N_1137,N_1197);
nand U1260 (N_1260,N_1116,N_1175);
nor U1261 (N_1261,N_1140,N_1100);
or U1262 (N_1262,N_1129,N_1174);
nor U1263 (N_1263,N_1151,N_1171);
xnor U1264 (N_1264,N_1166,N_1100);
or U1265 (N_1265,N_1151,N_1187);
and U1266 (N_1266,N_1101,N_1157);
and U1267 (N_1267,N_1135,N_1109);
nor U1268 (N_1268,N_1103,N_1146);
and U1269 (N_1269,N_1132,N_1124);
nor U1270 (N_1270,N_1171,N_1169);
or U1271 (N_1271,N_1185,N_1167);
nor U1272 (N_1272,N_1118,N_1193);
nand U1273 (N_1273,N_1113,N_1148);
and U1274 (N_1274,N_1187,N_1180);
and U1275 (N_1275,N_1161,N_1197);
and U1276 (N_1276,N_1153,N_1160);
nand U1277 (N_1277,N_1108,N_1171);
nor U1278 (N_1278,N_1119,N_1117);
and U1279 (N_1279,N_1132,N_1157);
nor U1280 (N_1280,N_1152,N_1199);
nand U1281 (N_1281,N_1104,N_1183);
nand U1282 (N_1282,N_1188,N_1152);
nand U1283 (N_1283,N_1133,N_1109);
or U1284 (N_1284,N_1158,N_1151);
and U1285 (N_1285,N_1159,N_1183);
nand U1286 (N_1286,N_1186,N_1155);
xor U1287 (N_1287,N_1169,N_1148);
nand U1288 (N_1288,N_1160,N_1175);
nor U1289 (N_1289,N_1107,N_1167);
nor U1290 (N_1290,N_1112,N_1175);
nand U1291 (N_1291,N_1179,N_1187);
and U1292 (N_1292,N_1108,N_1157);
and U1293 (N_1293,N_1168,N_1161);
nand U1294 (N_1294,N_1117,N_1165);
or U1295 (N_1295,N_1117,N_1181);
and U1296 (N_1296,N_1184,N_1186);
nand U1297 (N_1297,N_1196,N_1182);
and U1298 (N_1298,N_1116,N_1161);
nand U1299 (N_1299,N_1187,N_1182);
or U1300 (N_1300,N_1266,N_1223);
or U1301 (N_1301,N_1280,N_1221);
or U1302 (N_1302,N_1297,N_1286);
or U1303 (N_1303,N_1231,N_1271);
nor U1304 (N_1304,N_1233,N_1253);
and U1305 (N_1305,N_1211,N_1298);
xor U1306 (N_1306,N_1261,N_1201);
nor U1307 (N_1307,N_1263,N_1282);
nor U1308 (N_1308,N_1299,N_1219);
nand U1309 (N_1309,N_1256,N_1290);
or U1310 (N_1310,N_1204,N_1259);
or U1311 (N_1311,N_1241,N_1200);
and U1312 (N_1312,N_1270,N_1262);
nand U1313 (N_1313,N_1206,N_1207);
nor U1314 (N_1314,N_1293,N_1274);
xor U1315 (N_1315,N_1240,N_1228);
nor U1316 (N_1316,N_1225,N_1284);
or U1317 (N_1317,N_1208,N_1287);
or U1318 (N_1318,N_1295,N_1278);
nand U1319 (N_1319,N_1215,N_1230);
or U1320 (N_1320,N_1243,N_1224);
and U1321 (N_1321,N_1214,N_1257);
or U1322 (N_1322,N_1247,N_1268);
nor U1323 (N_1323,N_1239,N_1269);
or U1324 (N_1324,N_1276,N_1249);
nor U1325 (N_1325,N_1213,N_1209);
xnor U1326 (N_1326,N_1234,N_1289);
xnor U1327 (N_1327,N_1216,N_1245);
nor U1328 (N_1328,N_1220,N_1248);
nand U1329 (N_1329,N_1279,N_1238);
or U1330 (N_1330,N_1217,N_1222);
nor U1331 (N_1331,N_1203,N_1255);
nor U1332 (N_1332,N_1232,N_1202);
nand U1333 (N_1333,N_1267,N_1205);
xor U1334 (N_1334,N_1291,N_1226);
nor U1335 (N_1335,N_1244,N_1210);
nand U1336 (N_1336,N_1283,N_1294);
or U1337 (N_1337,N_1252,N_1273);
nor U1338 (N_1338,N_1212,N_1242);
nand U1339 (N_1339,N_1237,N_1251);
and U1340 (N_1340,N_1246,N_1258);
or U1341 (N_1341,N_1288,N_1229);
or U1342 (N_1342,N_1235,N_1250);
nor U1343 (N_1343,N_1285,N_1265);
nor U1344 (N_1344,N_1281,N_1277);
nand U1345 (N_1345,N_1236,N_1254);
nor U1346 (N_1346,N_1296,N_1292);
nand U1347 (N_1347,N_1272,N_1260);
or U1348 (N_1348,N_1275,N_1218);
xnor U1349 (N_1349,N_1227,N_1264);
nor U1350 (N_1350,N_1262,N_1279);
and U1351 (N_1351,N_1262,N_1260);
xor U1352 (N_1352,N_1218,N_1238);
and U1353 (N_1353,N_1273,N_1237);
or U1354 (N_1354,N_1264,N_1272);
nor U1355 (N_1355,N_1270,N_1277);
nand U1356 (N_1356,N_1208,N_1275);
xor U1357 (N_1357,N_1265,N_1204);
nor U1358 (N_1358,N_1231,N_1260);
xnor U1359 (N_1359,N_1215,N_1266);
nor U1360 (N_1360,N_1235,N_1281);
nor U1361 (N_1361,N_1270,N_1253);
xnor U1362 (N_1362,N_1234,N_1294);
nand U1363 (N_1363,N_1269,N_1240);
xor U1364 (N_1364,N_1294,N_1222);
and U1365 (N_1365,N_1261,N_1283);
nand U1366 (N_1366,N_1212,N_1221);
nor U1367 (N_1367,N_1212,N_1289);
nor U1368 (N_1368,N_1299,N_1252);
and U1369 (N_1369,N_1255,N_1260);
or U1370 (N_1370,N_1223,N_1235);
xor U1371 (N_1371,N_1215,N_1292);
nor U1372 (N_1372,N_1298,N_1250);
and U1373 (N_1373,N_1271,N_1209);
or U1374 (N_1374,N_1227,N_1255);
nor U1375 (N_1375,N_1207,N_1250);
nor U1376 (N_1376,N_1271,N_1202);
nand U1377 (N_1377,N_1240,N_1280);
or U1378 (N_1378,N_1218,N_1295);
nor U1379 (N_1379,N_1299,N_1258);
nor U1380 (N_1380,N_1253,N_1298);
or U1381 (N_1381,N_1262,N_1272);
and U1382 (N_1382,N_1229,N_1262);
nand U1383 (N_1383,N_1271,N_1273);
nand U1384 (N_1384,N_1213,N_1204);
xnor U1385 (N_1385,N_1208,N_1249);
or U1386 (N_1386,N_1225,N_1209);
and U1387 (N_1387,N_1228,N_1235);
xnor U1388 (N_1388,N_1242,N_1226);
and U1389 (N_1389,N_1251,N_1207);
nor U1390 (N_1390,N_1245,N_1242);
or U1391 (N_1391,N_1259,N_1253);
xnor U1392 (N_1392,N_1268,N_1292);
nand U1393 (N_1393,N_1279,N_1276);
nand U1394 (N_1394,N_1229,N_1217);
or U1395 (N_1395,N_1211,N_1273);
or U1396 (N_1396,N_1277,N_1203);
or U1397 (N_1397,N_1256,N_1205);
and U1398 (N_1398,N_1266,N_1221);
and U1399 (N_1399,N_1283,N_1231);
nor U1400 (N_1400,N_1399,N_1358);
and U1401 (N_1401,N_1378,N_1337);
nor U1402 (N_1402,N_1306,N_1346);
nand U1403 (N_1403,N_1388,N_1330);
or U1404 (N_1404,N_1331,N_1348);
xnor U1405 (N_1405,N_1325,N_1315);
or U1406 (N_1406,N_1381,N_1321);
nand U1407 (N_1407,N_1304,N_1332);
and U1408 (N_1408,N_1309,N_1371);
nor U1409 (N_1409,N_1302,N_1336);
or U1410 (N_1410,N_1328,N_1350);
nand U1411 (N_1411,N_1366,N_1342);
and U1412 (N_1412,N_1339,N_1308);
nor U1413 (N_1413,N_1312,N_1357);
and U1414 (N_1414,N_1393,N_1323);
nand U1415 (N_1415,N_1314,N_1351);
nand U1416 (N_1416,N_1365,N_1380);
and U1417 (N_1417,N_1389,N_1318);
and U1418 (N_1418,N_1345,N_1320);
and U1419 (N_1419,N_1311,N_1395);
and U1420 (N_1420,N_1335,N_1322);
nand U1421 (N_1421,N_1386,N_1376);
and U1422 (N_1422,N_1374,N_1344);
and U1423 (N_1423,N_1372,N_1363);
nand U1424 (N_1424,N_1317,N_1390);
nand U1425 (N_1425,N_1398,N_1340);
xor U1426 (N_1426,N_1319,N_1397);
xor U1427 (N_1427,N_1373,N_1349);
nor U1428 (N_1428,N_1305,N_1361);
or U1429 (N_1429,N_1359,N_1334);
and U1430 (N_1430,N_1300,N_1324);
nor U1431 (N_1431,N_1391,N_1326);
and U1432 (N_1432,N_1384,N_1360);
nor U1433 (N_1433,N_1301,N_1338);
nor U1434 (N_1434,N_1382,N_1313);
or U1435 (N_1435,N_1367,N_1310);
nand U1436 (N_1436,N_1316,N_1356);
nand U1437 (N_1437,N_1354,N_1333);
and U1438 (N_1438,N_1383,N_1370);
xor U1439 (N_1439,N_1347,N_1362);
nor U1440 (N_1440,N_1394,N_1329);
or U1441 (N_1441,N_1364,N_1377);
and U1442 (N_1442,N_1375,N_1369);
or U1443 (N_1443,N_1327,N_1341);
nor U1444 (N_1444,N_1355,N_1353);
or U1445 (N_1445,N_1379,N_1392);
or U1446 (N_1446,N_1343,N_1307);
nor U1447 (N_1447,N_1352,N_1387);
nand U1448 (N_1448,N_1385,N_1368);
or U1449 (N_1449,N_1396,N_1303);
nor U1450 (N_1450,N_1306,N_1310);
nor U1451 (N_1451,N_1356,N_1338);
or U1452 (N_1452,N_1376,N_1373);
nor U1453 (N_1453,N_1312,N_1330);
nand U1454 (N_1454,N_1327,N_1339);
or U1455 (N_1455,N_1350,N_1387);
nor U1456 (N_1456,N_1300,N_1301);
nand U1457 (N_1457,N_1388,N_1336);
and U1458 (N_1458,N_1383,N_1345);
xor U1459 (N_1459,N_1360,N_1364);
nor U1460 (N_1460,N_1309,N_1374);
nor U1461 (N_1461,N_1397,N_1348);
nand U1462 (N_1462,N_1353,N_1367);
nand U1463 (N_1463,N_1386,N_1381);
nand U1464 (N_1464,N_1382,N_1331);
and U1465 (N_1465,N_1390,N_1352);
nand U1466 (N_1466,N_1384,N_1353);
nand U1467 (N_1467,N_1318,N_1398);
and U1468 (N_1468,N_1397,N_1342);
and U1469 (N_1469,N_1310,N_1376);
nor U1470 (N_1470,N_1397,N_1385);
and U1471 (N_1471,N_1315,N_1330);
nor U1472 (N_1472,N_1347,N_1381);
or U1473 (N_1473,N_1334,N_1355);
nor U1474 (N_1474,N_1381,N_1350);
and U1475 (N_1475,N_1310,N_1303);
or U1476 (N_1476,N_1361,N_1391);
nor U1477 (N_1477,N_1368,N_1399);
and U1478 (N_1478,N_1337,N_1349);
and U1479 (N_1479,N_1315,N_1387);
xnor U1480 (N_1480,N_1393,N_1348);
or U1481 (N_1481,N_1346,N_1340);
nand U1482 (N_1482,N_1352,N_1317);
or U1483 (N_1483,N_1329,N_1380);
nand U1484 (N_1484,N_1362,N_1335);
and U1485 (N_1485,N_1342,N_1378);
and U1486 (N_1486,N_1346,N_1391);
and U1487 (N_1487,N_1357,N_1309);
and U1488 (N_1488,N_1358,N_1363);
and U1489 (N_1489,N_1338,N_1306);
xnor U1490 (N_1490,N_1367,N_1387);
xor U1491 (N_1491,N_1397,N_1360);
and U1492 (N_1492,N_1389,N_1374);
or U1493 (N_1493,N_1315,N_1359);
and U1494 (N_1494,N_1360,N_1306);
or U1495 (N_1495,N_1305,N_1370);
nor U1496 (N_1496,N_1344,N_1314);
and U1497 (N_1497,N_1347,N_1357);
and U1498 (N_1498,N_1310,N_1329);
nand U1499 (N_1499,N_1349,N_1320);
and U1500 (N_1500,N_1422,N_1448);
nor U1501 (N_1501,N_1471,N_1469);
xor U1502 (N_1502,N_1411,N_1408);
nand U1503 (N_1503,N_1451,N_1476);
nand U1504 (N_1504,N_1414,N_1462);
and U1505 (N_1505,N_1467,N_1402);
and U1506 (N_1506,N_1423,N_1445);
or U1507 (N_1507,N_1418,N_1457);
and U1508 (N_1508,N_1403,N_1480);
or U1509 (N_1509,N_1413,N_1459);
xnor U1510 (N_1510,N_1401,N_1425);
xor U1511 (N_1511,N_1450,N_1482);
and U1512 (N_1512,N_1412,N_1405);
nand U1513 (N_1513,N_1416,N_1486);
nand U1514 (N_1514,N_1447,N_1433);
nor U1515 (N_1515,N_1434,N_1436);
nor U1516 (N_1516,N_1409,N_1454);
nor U1517 (N_1517,N_1494,N_1441);
nand U1518 (N_1518,N_1498,N_1446);
nor U1519 (N_1519,N_1435,N_1417);
nand U1520 (N_1520,N_1481,N_1439);
nor U1521 (N_1521,N_1493,N_1488);
or U1522 (N_1522,N_1489,N_1484);
or U1523 (N_1523,N_1453,N_1496);
nand U1524 (N_1524,N_1440,N_1410);
nor U1525 (N_1525,N_1490,N_1452);
nand U1526 (N_1526,N_1487,N_1415);
nand U1527 (N_1527,N_1466,N_1473);
or U1528 (N_1528,N_1479,N_1499);
and U1529 (N_1529,N_1464,N_1407);
xnor U1530 (N_1530,N_1400,N_1456);
nand U1531 (N_1531,N_1470,N_1485);
or U1532 (N_1532,N_1492,N_1475);
and U1533 (N_1533,N_1419,N_1495);
or U1534 (N_1534,N_1426,N_1421);
xnor U1535 (N_1535,N_1437,N_1429);
or U1536 (N_1536,N_1474,N_1444);
or U1537 (N_1537,N_1468,N_1404);
nor U1538 (N_1538,N_1491,N_1497);
or U1539 (N_1539,N_1478,N_1427);
and U1540 (N_1540,N_1483,N_1424);
nor U1541 (N_1541,N_1465,N_1449);
or U1542 (N_1542,N_1438,N_1406);
or U1543 (N_1543,N_1460,N_1443);
nor U1544 (N_1544,N_1432,N_1472);
and U1545 (N_1545,N_1420,N_1428);
xnor U1546 (N_1546,N_1463,N_1458);
xor U1547 (N_1547,N_1477,N_1442);
and U1548 (N_1548,N_1431,N_1455);
or U1549 (N_1549,N_1430,N_1461);
nor U1550 (N_1550,N_1452,N_1445);
and U1551 (N_1551,N_1438,N_1499);
and U1552 (N_1552,N_1468,N_1405);
nand U1553 (N_1553,N_1472,N_1436);
nand U1554 (N_1554,N_1472,N_1453);
and U1555 (N_1555,N_1478,N_1423);
or U1556 (N_1556,N_1478,N_1438);
and U1557 (N_1557,N_1467,N_1493);
and U1558 (N_1558,N_1479,N_1485);
nand U1559 (N_1559,N_1489,N_1461);
nand U1560 (N_1560,N_1410,N_1476);
and U1561 (N_1561,N_1455,N_1452);
or U1562 (N_1562,N_1403,N_1440);
and U1563 (N_1563,N_1435,N_1410);
xnor U1564 (N_1564,N_1403,N_1497);
nand U1565 (N_1565,N_1464,N_1436);
or U1566 (N_1566,N_1401,N_1478);
and U1567 (N_1567,N_1414,N_1455);
xnor U1568 (N_1568,N_1452,N_1435);
nand U1569 (N_1569,N_1484,N_1464);
nor U1570 (N_1570,N_1429,N_1475);
and U1571 (N_1571,N_1430,N_1468);
or U1572 (N_1572,N_1497,N_1479);
or U1573 (N_1573,N_1438,N_1493);
nor U1574 (N_1574,N_1432,N_1402);
nand U1575 (N_1575,N_1412,N_1479);
nand U1576 (N_1576,N_1487,N_1435);
or U1577 (N_1577,N_1492,N_1441);
or U1578 (N_1578,N_1403,N_1429);
nand U1579 (N_1579,N_1450,N_1498);
and U1580 (N_1580,N_1408,N_1409);
nor U1581 (N_1581,N_1431,N_1437);
nor U1582 (N_1582,N_1451,N_1493);
nand U1583 (N_1583,N_1466,N_1443);
nor U1584 (N_1584,N_1493,N_1479);
nand U1585 (N_1585,N_1454,N_1458);
nand U1586 (N_1586,N_1414,N_1446);
or U1587 (N_1587,N_1415,N_1450);
or U1588 (N_1588,N_1463,N_1416);
nor U1589 (N_1589,N_1435,N_1461);
or U1590 (N_1590,N_1450,N_1405);
xor U1591 (N_1591,N_1426,N_1451);
or U1592 (N_1592,N_1430,N_1497);
or U1593 (N_1593,N_1468,N_1439);
and U1594 (N_1594,N_1452,N_1448);
or U1595 (N_1595,N_1459,N_1495);
and U1596 (N_1596,N_1476,N_1478);
nand U1597 (N_1597,N_1455,N_1411);
xor U1598 (N_1598,N_1430,N_1438);
or U1599 (N_1599,N_1464,N_1475);
nor U1600 (N_1600,N_1534,N_1523);
nand U1601 (N_1601,N_1561,N_1501);
or U1602 (N_1602,N_1558,N_1554);
or U1603 (N_1603,N_1507,N_1551);
and U1604 (N_1604,N_1589,N_1515);
xnor U1605 (N_1605,N_1504,N_1541);
nor U1606 (N_1606,N_1560,N_1590);
and U1607 (N_1607,N_1574,N_1533);
or U1608 (N_1608,N_1584,N_1509);
and U1609 (N_1609,N_1569,N_1544);
and U1610 (N_1610,N_1527,N_1562);
nand U1611 (N_1611,N_1516,N_1546);
or U1612 (N_1612,N_1578,N_1545);
nand U1613 (N_1613,N_1548,N_1525);
nand U1614 (N_1614,N_1598,N_1587);
and U1615 (N_1615,N_1505,N_1595);
nor U1616 (N_1616,N_1512,N_1543);
or U1617 (N_1617,N_1599,N_1579);
xnor U1618 (N_1618,N_1529,N_1513);
nor U1619 (N_1619,N_1526,N_1594);
nand U1620 (N_1620,N_1550,N_1538);
and U1621 (N_1621,N_1592,N_1555);
and U1622 (N_1622,N_1542,N_1571);
xnor U1623 (N_1623,N_1506,N_1532);
nand U1624 (N_1624,N_1580,N_1518);
and U1625 (N_1625,N_1576,N_1522);
xnor U1626 (N_1626,N_1575,N_1552);
nor U1627 (N_1627,N_1524,N_1553);
nand U1628 (N_1628,N_1581,N_1517);
or U1629 (N_1629,N_1536,N_1559);
nor U1630 (N_1630,N_1539,N_1508);
or U1631 (N_1631,N_1514,N_1596);
and U1632 (N_1632,N_1570,N_1597);
nand U1633 (N_1633,N_1583,N_1503);
or U1634 (N_1634,N_1563,N_1521);
and U1635 (N_1635,N_1540,N_1588);
nor U1636 (N_1636,N_1511,N_1500);
and U1637 (N_1637,N_1591,N_1564);
nor U1638 (N_1638,N_1519,N_1585);
nand U1639 (N_1639,N_1537,N_1535);
nand U1640 (N_1640,N_1510,N_1573);
nor U1641 (N_1641,N_1528,N_1520);
or U1642 (N_1642,N_1572,N_1567);
or U1643 (N_1643,N_1566,N_1593);
xnor U1644 (N_1644,N_1586,N_1531);
and U1645 (N_1645,N_1577,N_1568);
nand U1646 (N_1646,N_1565,N_1502);
and U1647 (N_1647,N_1549,N_1530);
nand U1648 (N_1648,N_1582,N_1547);
or U1649 (N_1649,N_1556,N_1557);
nor U1650 (N_1650,N_1507,N_1526);
nor U1651 (N_1651,N_1598,N_1559);
xor U1652 (N_1652,N_1536,N_1549);
or U1653 (N_1653,N_1548,N_1586);
nor U1654 (N_1654,N_1556,N_1595);
nor U1655 (N_1655,N_1527,N_1598);
and U1656 (N_1656,N_1544,N_1509);
and U1657 (N_1657,N_1523,N_1572);
nand U1658 (N_1658,N_1562,N_1572);
nor U1659 (N_1659,N_1509,N_1591);
or U1660 (N_1660,N_1531,N_1543);
nor U1661 (N_1661,N_1515,N_1599);
nor U1662 (N_1662,N_1547,N_1550);
and U1663 (N_1663,N_1583,N_1529);
or U1664 (N_1664,N_1559,N_1568);
nor U1665 (N_1665,N_1589,N_1558);
nor U1666 (N_1666,N_1554,N_1508);
nor U1667 (N_1667,N_1528,N_1525);
nor U1668 (N_1668,N_1577,N_1519);
nand U1669 (N_1669,N_1511,N_1556);
xnor U1670 (N_1670,N_1520,N_1557);
nor U1671 (N_1671,N_1596,N_1550);
nor U1672 (N_1672,N_1579,N_1514);
nor U1673 (N_1673,N_1568,N_1510);
and U1674 (N_1674,N_1545,N_1571);
or U1675 (N_1675,N_1508,N_1580);
nand U1676 (N_1676,N_1583,N_1524);
or U1677 (N_1677,N_1573,N_1583);
nand U1678 (N_1678,N_1512,N_1570);
nor U1679 (N_1679,N_1540,N_1595);
or U1680 (N_1680,N_1545,N_1500);
and U1681 (N_1681,N_1562,N_1543);
or U1682 (N_1682,N_1508,N_1540);
xnor U1683 (N_1683,N_1571,N_1532);
xnor U1684 (N_1684,N_1503,N_1500);
and U1685 (N_1685,N_1550,N_1511);
and U1686 (N_1686,N_1506,N_1543);
or U1687 (N_1687,N_1565,N_1585);
nor U1688 (N_1688,N_1502,N_1509);
and U1689 (N_1689,N_1509,N_1507);
xnor U1690 (N_1690,N_1555,N_1530);
xor U1691 (N_1691,N_1562,N_1556);
or U1692 (N_1692,N_1510,N_1532);
or U1693 (N_1693,N_1556,N_1543);
or U1694 (N_1694,N_1548,N_1591);
or U1695 (N_1695,N_1559,N_1550);
nand U1696 (N_1696,N_1528,N_1542);
and U1697 (N_1697,N_1573,N_1547);
or U1698 (N_1698,N_1516,N_1573);
and U1699 (N_1699,N_1552,N_1544);
or U1700 (N_1700,N_1647,N_1605);
and U1701 (N_1701,N_1688,N_1668);
and U1702 (N_1702,N_1695,N_1694);
and U1703 (N_1703,N_1669,N_1649);
nor U1704 (N_1704,N_1628,N_1614);
nand U1705 (N_1705,N_1665,N_1673);
nor U1706 (N_1706,N_1661,N_1646);
and U1707 (N_1707,N_1693,N_1687);
nand U1708 (N_1708,N_1626,N_1641);
or U1709 (N_1709,N_1655,N_1659);
nor U1710 (N_1710,N_1631,N_1634);
nor U1711 (N_1711,N_1645,N_1638);
xnor U1712 (N_1712,N_1680,N_1632);
or U1713 (N_1713,N_1651,N_1689);
or U1714 (N_1714,N_1610,N_1624);
nand U1715 (N_1715,N_1636,N_1603);
nand U1716 (N_1716,N_1670,N_1675);
nand U1717 (N_1717,N_1686,N_1640);
or U1718 (N_1718,N_1676,N_1600);
nand U1719 (N_1719,N_1653,N_1621);
and U1720 (N_1720,N_1698,N_1616);
and U1721 (N_1721,N_1664,N_1667);
nand U1722 (N_1722,N_1611,N_1620);
and U1723 (N_1723,N_1643,N_1672);
or U1724 (N_1724,N_1613,N_1678);
nand U1725 (N_1725,N_1617,N_1642);
and U1726 (N_1726,N_1602,N_1635);
nor U1727 (N_1727,N_1684,N_1657);
and U1728 (N_1728,N_1682,N_1604);
or U1729 (N_1729,N_1696,N_1606);
and U1730 (N_1730,N_1677,N_1679);
xor U1731 (N_1731,N_1697,N_1690);
and U1732 (N_1732,N_1630,N_1658);
nand U1733 (N_1733,N_1652,N_1609);
xnor U1734 (N_1734,N_1662,N_1623);
nor U1735 (N_1735,N_1627,N_1663);
nand U1736 (N_1736,N_1601,N_1612);
xnor U1737 (N_1737,N_1691,N_1618);
or U1738 (N_1738,N_1615,N_1650);
or U1739 (N_1739,N_1644,N_1671);
or U1740 (N_1740,N_1683,N_1699);
nand U1741 (N_1741,N_1648,N_1681);
or U1742 (N_1742,N_1619,N_1666);
and U1743 (N_1743,N_1629,N_1660);
nand U1744 (N_1744,N_1637,N_1685);
or U1745 (N_1745,N_1674,N_1633);
or U1746 (N_1746,N_1654,N_1656);
nor U1747 (N_1747,N_1625,N_1607);
nand U1748 (N_1748,N_1622,N_1608);
or U1749 (N_1749,N_1639,N_1692);
and U1750 (N_1750,N_1690,N_1641);
nand U1751 (N_1751,N_1682,N_1635);
or U1752 (N_1752,N_1671,N_1665);
nand U1753 (N_1753,N_1629,N_1672);
and U1754 (N_1754,N_1669,N_1679);
and U1755 (N_1755,N_1608,N_1623);
or U1756 (N_1756,N_1645,N_1615);
xnor U1757 (N_1757,N_1638,N_1671);
or U1758 (N_1758,N_1676,N_1655);
nor U1759 (N_1759,N_1678,N_1649);
or U1760 (N_1760,N_1689,N_1661);
nand U1761 (N_1761,N_1616,N_1623);
nor U1762 (N_1762,N_1648,N_1643);
or U1763 (N_1763,N_1613,N_1674);
or U1764 (N_1764,N_1658,N_1621);
nand U1765 (N_1765,N_1611,N_1643);
nor U1766 (N_1766,N_1667,N_1601);
and U1767 (N_1767,N_1633,N_1666);
nand U1768 (N_1768,N_1606,N_1668);
and U1769 (N_1769,N_1616,N_1631);
and U1770 (N_1770,N_1632,N_1676);
xnor U1771 (N_1771,N_1661,N_1638);
or U1772 (N_1772,N_1695,N_1656);
nand U1773 (N_1773,N_1671,N_1689);
and U1774 (N_1774,N_1620,N_1653);
or U1775 (N_1775,N_1678,N_1690);
nor U1776 (N_1776,N_1618,N_1607);
and U1777 (N_1777,N_1605,N_1600);
and U1778 (N_1778,N_1673,N_1605);
and U1779 (N_1779,N_1626,N_1647);
or U1780 (N_1780,N_1613,N_1687);
and U1781 (N_1781,N_1687,N_1698);
and U1782 (N_1782,N_1635,N_1672);
and U1783 (N_1783,N_1699,N_1629);
and U1784 (N_1784,N_1686,N_1697);
and U1785 (N_1785,N_1665,N_1681);
nor U1786 (N_1786,N_1696,N_1678);
nor U1787 (N_1787,N_1653,N_1611);
and U1788 (N_1788,N_1601,N_1648);
or U1789 (N_1789,N_1650,N_1607);
and U1790 (N_1790,N_1642,N_1651);
xnor U1791 (N_1791,N_1660,N_1674);
nor U1792 (N_1792,N_1631,N_1684);
nand U1793 (N_1793,N_1603,N_1641);
or U1794 (N_1794,N_1615,N_1687);
xnor U1795 (N_1795,N_1677,N_1682);
nor U1796 (N_1796,N_1636,N_1653);
or U1797 (N_1797,N_1682,N_1672);
and U1798 (N_1798,N_1643,N_1665);
or U1799 (N_1799,N_1679,N_1629);
nand U1800 (N_1800,N_1728,N_1760);
nand U1801 (N_1801,N_1773,N_1711);
nor U1802 (N_1802,N_1798,N_1720);
nor U1803 (N_1803,N_1764,N_1724);
nor U1804 (N_1804,N_1781,N_1715);
nor U1805 (N_1805,N_1741,N_1784);
and U1806 (N_1806,N_1772,N_1752);
and U1807 (N_1807,N_1718,N_1717);
and U1808 (N_1808,N_1740,N_1786);
nor U1809 (N_1809,N_1769,N_1739);
or U1810 (N_1810,N_1761,N_1770);
nand U1811 (N_1811,N_1707,N_1756);
and U1812 (N_1812,N_1729,N_1731);
or U1813 (N_1813,N_1791,N_1721);
nand U1814 (N_1814,N_1792,N_1723);
nand U1815 (N_1815,N_1735,N_1754);
nor U1816 (N_1816,N_1771,N_1758);
and U1817 (N_1817,N_1779,N_1700);
and U1818 (N_1818,N_1710,N_1763);
nand U1819 (N_1819,N_1734,N_1757);
nor U1820 (N_1820,N_1749,N_1726);
nor U1821 (N_1821,N_1778,N_1790);
nand U1822 (N_1822,N_1799,N_1725);
nand U1823 (N_1823,N_1744,N_1796);
and U1824 (N_1824,N_1703,N_1795);
or U1825 (N_1825,N_1768,N_1742);
or U1826 (N_1826,N_1708,N_1701);
nand U1827 (N_1827,N_1746,N_1732);
or U1828 (N_1828,N_1712,N_1797);
or U1829 (N_1829,N_1762,N_1719);
nand U1830 (N_1830,N_1765,N_1727);
nor U1831 (N_1831,N_1737,N_1706);
nand U1832 (N_1832,N_1777,N_1702);
xor U1833 (N_1833,N_1767,N_1794);
xor U1834 (N_1834,N_1774,N_1775);
and U1835 (N_1835,N_1709,N_1716);
nor U1836 (N_1836,N_1751,N_1787);
and U1837 (N_1837,N_1748,N_1753);
nand U1838 (N_1838,N_1747,N_1713);
and U1839 (N_1839,N_1793,N_1730);
and U1840 (N_1840,N_1738,N_1782);
nor U1841 (N_1841,N_1789,N_1766);
nor U1842 (N_1842,N_1776,N_1736);
nand U1843 (N_1843,N_1714,N_1722);
nand U1844 (N_1844,N_1780,N_1733);
nand U1845 (N_1845,N_1788,N_1750);
and U1846 (N_1846,N_1704,N_1755);
or U1847 (N_1847,N_1783,N_1705);
and U1848 (N_1848,N_1759,N_1745);
nor U1849 (N_1849,N_1785,N_1743);
nor U1850 (N_1850,N_1708,N_1787);
nor U1851 (N_1851,N_1796,N_1707);
and U1852 (N_1852,N_1776,N_1726);
nor U1853 (N_1853,N_1750,N_1711);
nor U1854 (N_1854,N_1762,N_1794);
or U1855 (N_1855,N_1770,N_1700);
xor U1856 (N_1856,N_1765,N_1706);
nand U1857 (N_1857,N_1793,N_1794);
nand U1858 (N_1858,N_1771,N_1790);
nor U1859 (N_1859,N_1738,N_1759);
and U1860 (N_1860,N_1794,N_1764);
or U1861 (N_1861,N_1742,N_1770);
nor U1862 (N_1862,N_1735,N_1724);
nor U1863 (N_1863,N_1777,N_1791);
or U1864 (N_1864,N_1753,N_1794);
or U1865 (N_1865,N_1747,N_1785);
nor U1866 (N_1866,N_1792,N_1775);
xnor U1867 (N_1867,N_1717,N_1731);
and U1868 (N_1868,N_1777,N_1753);
nor U1869 (N_1869,N_1760,N_1716);
nor U1870 (N_1870,N_1701,N_1753);
or U1871 (N_1871,N_1760,N_1767);
nor U1872 (N_1872,N_1776,N_1710);
or U1873 (N_1873,N_1796,N_1766);
nor U1874 (N_1874,N_1756,N_1787);
and U1875 (N_1875,N_1729,N_1785);
nor U1876 (N_1876,N_1799,N_1722);
or U1877 (N_1877,N_1739,N_1750);
and U1878 (N_1878,N_1737,N_1732);
nor U1879 (N_1879,N_1786,N_1788);
nor U1880 (N_1880,N_1776,N_1768);
nor U1881 (N_1881,N_1723,N_1712);
and U1882 (N_1882,N_1720,N_1749);
or U1883 (N_1883,N_1710,N_1764);
nor U1884 (N_1884,N_1749,N_1778);
and U1885 (N_1885,N_1722,N_1778);
xor U1886 (N_1886,N_1728,N_1733);
nand U1887 (N_1887,N_1740,N_1792);
and U1888 (N_1888,N_1768,N_1718);
nor U1889 (N_1889,N_1754,N_1741);
or U1890 (N_1890,N_1751,N_1746);
nor U1891 (N_1891,N_1772,N_1749);
nor U1892 (N_1892,N_1757,N_1742);
or U1893 (N_1893,N_1785,N_1733);
nor U1894 (N_1894,N_1772,N_1775);
or U1895 (N_1895,N_1747,N_1765);
or U1896 (N_1896,N_1723,N_1735);
and U1897 (N_1897,N_1791,N_1784);
or U1898 (N_1898,N_1722,N_1720);
or U1899 (N_1899,N_1729,N_1750);
xnor U1900 (N_1900,N_1856,N_1861);
and U1901 (N_1901,N_1829,N_1809);
nand U1902 (N_1902,N_1837,N_1810);
or U1903 (N_1903,N_1873,N_1886);
and U1904 (N_1904,N_1899,N_1817);
or U1905 (N_1905,N_1881,N_1821);
and U1906 (N_1906,N_1845,N_1814);
nand U1907 (N_1907,N_1870,N_1868);
nor U1908 (N_1908,N_1812,N_1800);
and U1909 (N_1909,N_1889,N_1884);
or U1910 (N_1910,N_1848,N_1872);
nor U1911 (N_1911,N_1887,N_1807);
or U1912 (N_1912,N_1835,N_1855);
nor U1913 (N_1913,N_1895,N_1854);
or U1914 (N_1914,N_1871,N_1878);
and U1915 (N_1915,N_1828,N_1849);
xnor U1916 (N_1916,N_1816,N_1876);
nor U1917 (N_1917,N_1864,N_1825);
xor U1918 (N_1918,N_1827,N_1882);
nand U1919 (N_1919,N_1820,N_1883);
or U1920 (N_1920,N_1806,N_1838);
nand U1921 (N_1921,N_1865,N_1802);
xor U1922 (N_1922,N_1897,N_1808);
or U1923 (N_1923,N_1875,N_1859);
nor U1924 (N_1924,N_1804,N_1818);
and U1925 (N_1925,N_1880,N_1874);
and U1926 (N_1926,N_1847,N_1877);
xor U1927 (N_1927,N_1832,N_1836);
nand U1928 (N_1928,N_1863,N_1801);
and U1929 (N_1929,N_1840,N_1885);
or U1930 (N_1930,N_1893,N_1858);
nor U1931 (N_1931,N_1819,N_1857);
xnor U1932 (N_1932,N_1853,N_1830);
nand U1933 (N_1933,N_1892,N_1833);
or U1934 (N_1934,N_1803,N_1851);
nand U1935 (N_1935,N_1860,N_1890);
and U1936 (N_1936,N_1896,N_1888);
nor U1937 (N_1937,N_1834,N_1869);
nand U1938 (N_1938,N_1894,N_1862);
and U1939 (N_1939,N_1822,N_1824);
nor U1940 (N_1940,N_1842,N_1815);
xnor U1941 (N_1941,N_1841,N_1866);
or U1942 (N_1942,N_1826,N_1831);
nand U1943 (N_1943,N_1813,N_1879);
and U1944 (N_1944,N_1823,N_1811);
nand U1945 (N_1945,N_1843,N_1839);
and U1946 (N_1946,N_1852,N_1844);
or U1947 (N_1947,N_1846,N_1898);
or U1948 (N_1948,N_1805,N_1867);
xor U1949 (N_1949,N_1891,N_1850);
nand U1950 (N_1950,N_1817,N_1822);
nand U1951 (N_1951,N_1879,N_1891);
or U1952 (N_1952,N_1816,N_1883);
nor U1953 (N_1953,N_1812,N_1879);
nand U1954 (N_1954,N_1856,N_1832);
nand U1955 (N_1955,N_1831,N_1821);
nand U1956 (N_1956,N_1875,N_1805);
or U1957 (N_1957,N_1861,N_1812);
or U1958 (N_1958,N_1840,N_1826);
nand U1959 (N_1959,N_1817,N_1864);
or U1960 (N_1960,N_1893,N_1870);
or U1961 (N_1961,N_1898,N_1874);
or U1962 (N_1962,N_1840,N_1847);
and U1963 (N_1963,N_1870,N_1884);
nor U1964 (N_1964,N_1892,N_1808);
nor U1965 (N_1965,N_1850,N_1813);
nor U1966 (N_1966,N_1823,N_1880);
or U1967 (N_1967,N_1828,N_1870);
nor U1968 (N_1968,N_1844,N_1853);
nand U1969 (N_1969,N_1834,N_1824);
nor U1970 (N_1970,N_1802,N_1894);
nand U1971 (N_1971,N_1885,N_1888);
and U1972 (N_1972,N_1814,N_1827);
and U1973 (N_1973,N_1849,N_1877);
nor U1974 (N_1974,N_1818,N_1845);
nor U1975 (N_1975,N_1825,N_1816);
nand U1976 (N_1976,N_1872,N_1869);
xnor U1977 (N_1977,N_1827,N_1843);
or U1978 (N_1978,N_1804,N_1894);
nor U1979 (N_1979,N_1866,N_1864);
and U1980 (N_1980,N_1816,N_1897);
nor U1981 (N_1981,N_1864,N_1847);
and U1982 (N_1982,N_1851,N_1820);
and U1983 (N_1983,N_1899,N_1894);
nand U1984 (N_1984,N_1843,N_1890);
and U1985 (N_1985,N_1863,N_1885);
and U1986 (N_1986,N_1862,N_1824);
or U1987 (N_1987,N_1803,N_1841);
and U1988 (N_1988,N_1870,N_1812);
or U1989 (N_1989,N_1864,N_1813);
nor U1990 (N_1990,N_1838,N_1812);
nand U1991 (N_1991,N_1880,N_1820);
xor U1992 (N_1992,N_1845,N_1833);
nor U1993 (N_1993,N_1851,N_1862);
nor U1994 (N_1994,N_1859,N_1895);
or U1995 (N_1995,N_1868,N_1827);
nand U1996 (N_1996,N_1813,N_1806);
xor U1997 (N_1997,N_1803,N_1886);
or U1998 (N_1998,N_1836,N_1807);
xnor U1999 (N_1999,N_1816,N_1891);
or U2000 (N_2000,N_1973,N_1929);
and U2001 (N_2001,N_1982,N_1945);
nand U2002 (N_2002,N_1999,N_1951);
nand U2003 (N_2003,N_1972,N_1989);
nand U2004 (N_2004,N_1934,N_1948);
nor U2005 (N_2005,N_1907,N_1961);
nand U2006 (N_2006,N_1904,N_1966);
nand U2007 (N_2007,N_1921,N_1983);
nor U2008 (N_2008,N_1937,N_1985);
or U2009 (N_2009,N_1917,N_1991);
or U2010 (N_2010,N_1984,N_1970);
nand U2011 (N_2011,N_1969,N_1939);
nor U2012 (N_2012,N_1974,N_1909);
xnor U2013 (N_2013,N_1981,N_1931);
xnor U2014 (N_2014,N_1987,N_1975);
or U2015 (N_2015,N_1990,N_1986);
nand U2016 (N_2016,N_1968,N_1935);
and U2017 (N_2017,N_1952,N_1956);
nand U2018 (N_2018,N_1938,N_1903);
or U2019 (N_2019,N_1950,N_1927);
and U2020 (N_2020,N_1916,N_1905);
nor U2021 (N_2021,N_1944,N_1902);
nand U2022 (N_2022,N_1993,N_1913);
and U2023 (N_2023,N_1995,N_1915);
or U2024 (N_2024,N_1911,N_1958);
or U2025 (N_2025,N_1901,N_1971);
xnor U2026 (N_2026,N_1910,N_1919);
or U2027 (N_2027,N_1959,N_1930);
and U2028 (N_2028,N_1941,N_1960);
nor U2029 (N_2029,N_1908,N_1912);
and U2030 (N_2030,N_1967,N_1914);
xor U2031 (N_2031,N_1979,N_1978);
or U2032 (N_2032,N_1926,N_1918);
nand U2033 (N_2033,N_1906,N_1977);
and U2034 (N_2034,N_1936,N_1965);
xor U2035 (N_2035,N_1940,N_1954);
nand U2036 (N_2036,N_1980,N_1942);
nand U2037 (N_2037,N_1923,N_1946);
nor U2038 (N_2038,N_1922,N_1943);
nand U2039 (N_2039,N_1920,N_1933);
xor U2040 (N_2040,N_1957,N_1997);
and U2041 (N_2041,N_1932,N_1988);
nor U2042 (N_2042,N_1925,N_1955);
nor U2043 (N_2043,N_1949,N_1928);
and U2044 (N_2044,N_1998,N_1963);
or U2045 (N_2045,N_1900,N_1976);
and U2046 (N_2046,N_1994,N_1996);
nand U2047 (N_2047,N_1953,N_1964);
xor U2048 (N_2048,N_1924,N_1962);
nor U2049 (N_2049,N_1947,N_1992);
nor U2050 (N_2050,N_1918,N_1908);
nor U2051 (N_2051,N_1917,N_1961);
or U2052 (N_2052,N_1955,N_1938);
and U2053 (N_2053,N_1972,N_1954);
and U2054 (N_2054,N_1998,N_1971);
nor U2055 (N_2055,N_1995,N_1979);
nor U2056 (N_2056,N_1960,N_1932);
nor U2057 (N_2057,N_1932,N_1924);
nand U2058 (N_2058,N_1904,N_1950);
and U2059 (N_2059,N_1975,N_1981);
nor U2060 (N_2060,N_1998,N_1900);
nand U2061 (N_2061,N_1961,N_1998);
nor U2062 (N_2062,N_1914,N_1900);
or U2063 (N_2063,N_1994,N_1990);
or U2064 (N_2064,N_1964,N_1905);
nor U2065 (N_2065,N_1934,N_1935);
nand U2066 (N_2066,N_1901,N_1944);
or U2067 (N_2067,N_1940,N_1991);
or U2068 (N_2068,N_1962,N_1970);
and U2069 (N_2069,N_1957,N_1981);
and U2070 (N_2070,N_1993,N_1914);
or U2071 (N_2071,N_1962,N_1952);
nor U2072 (N_2072,N_1978,N_1939);
xor U2073 (N_2073,N_1977,N_1996);
or U2074 (N_2074,N_1903,N_1998);
or U2075 (N_2075,N_1903,N_1934);
nor U2076 (N_2076,N_1980,N_1977);
and U2077 (N_2077,N_1900,N_1906);
nor U2078 (N_2078,N_1999,N_1984);
or U2079 (N_2079,N_1964,N_1970);
nand U2080 (N_2080,N_1956,N_1967);
nor U2081 (N_2081,N_1973,N_1930);
nand U2082 (N_2082,N_1927,N_1995);
or U2083 (N_2083,N_1907,N_1977);
nand U2084 (N_2084,N_1973,N_1967);
and U2085 (N_2085,N_1966,N_1984);
and U2086 (N_2086,N_1940,N_1986);
xor U2087 (N_2087,N_1939,N_1920);
nand U2088 (N_2088,N_1923,N_1905);
nand U2089 (N_2089,N_1939,N_1909);
nand U2090 (N_2090,N_1952,N_1936);
and U2091 (N_2091,N_1921,N_1957);
or U2092 (N_2092,N_1985,N_1915);
and U2093 (N_2093,N_1993,N_1995);
nor U2094 (N_2094,N_1920,N_1973);
or U2095 (N_2095,N_1932,N_1926);
or U2096 (N_2096,N_1951,N_1909);
nand U2097 (N_2097,N_1922,N_1966);
nor U2098 (N_2098,N_1923,N_1944);
or U2099 (N_2099,N_1954,N_1999);
nor U2100 (N_2100,N_2051,N_2073);
nand U2101 (N_2101,N_2035,N_2005);
and U2102 (N_2102,N_2061,N_2003);
and U2103 (N_2103,N_2078,N_2008);
and U2104 (N_2104,N_2086,N_2033);
nor U2105 (N_2105,N_2026,N_2006);
xnor U2106 (N_2106,N_2012,N_2076);
or U2107 (N_2107,N_2010,N_2077);
and U2108 (N_2108,N_2065,N_2069);
nor U2109 (N_2109,N_2055,N_2017);
nor U2110 (N_2110,N_2080,N_2016);
or U2111 (N_2111,N_2060,N_2043);
nor U2112 (N_2112,N_2050,N_2067);
nand U2113 (N_2113,N_2087,N_2062);
and U2114 (N_2114,N_2015,N_2014);
nor U2115 (N_2115,N_2040,N_2023);
xor U2116 (N_2116,N_2011,N_2058);
and U2117 (N_2117,N_2022,N_2049);
nand U2118 (N_2118,N_2024,N_2041);
nor U2119 (N_2119,N_2059,N_2030);
or U2120 (N_2120,N_2052,N_2098);
or U2121 (N_2121,N_2085,N_2053);
nor U2122 (N_2122,N_2029,N_2096);
nand U2123 (N_2123,N_2032,N_2034);
or U2124 (N_2124,N_2063,N_2039);
nand U2125 (N_2125,N_2018,N_2054);
nor U2126 (N_2126,N_2013,N_2071);
nor U2127 (N_2127,N_2045,N_2019);
and U2128 (N_2128,N_2074,N_2082);
or U2129 (N_2129,N_2083,N_2097);
or U2130 (N_2130,N_2000,N_2070);
nor U2131 (N_2131,N_2092,N_2004);
or U2132 (N_2132,N_2081,N_2009);
nor U2133 (N_2133,N_2066,N_2028);
nor U2134 (N_2134,N_2037,N_2044);
nor U2135 (N_2135,N_2001,N_2091);
nor U2136 (N_2136,N_2093,N_2064);
xor U2137 (N_2137,N_2056,N_2046);
or U2138 (N_2138,N_2031,N_2036);
xor U2139 (N_2139,N_2038,N_2084);
and U2140 (N_2140,N_2021,N_2048);
or U2141 (N_2141,N_2089,N_2025);
nor U2142 (N_2142,N_2094,N_2042);
nand U2143 (N_2143,N_2057,N_2068);
nand U2144 (N_2144,N_2090,N_2099);
and U2145 (N_2145,N_2007,N_2002);
and U2146 (N_2146,N_2047,N_2020);
nor U2147 (N_2147,N_2088,N_2072);
nor U2148 (N_2148,N_2027,N_2075);
nor U2149 (N_2149,N_2079,N_2095);
or U2150 (N_2150,N_2063,N_2091);
nand U2151 (N_2151,N_2068,N_2060);
or U2152 (N_2152,N_2097,N_2000);
nor U2153 (N_2153,N_2093,N_2078);
nand U2154 (N_2154,N_2090,N_2051);
nand U2155 (N_2155,N_2029,N_2038);
nand U2156 (N_2156,N_2076,N_2023);
xor U2157 (N_2157,N_2024,N_2020);
nand U2158 (N_2158,N_2023,N_2024);
xnor U2159 (N_2159,N_2018,N_2061);
and U2160 (N_2160,N_2061,N_2073);
xnor U2161 (N_2161,N_2023,N_2008);
nor U2162 (N_2162,N_2060,N_2050);
or U2163 (N_2163,N_2052,N_2009);
nor U2164 (N_2164,N_2029,N_2006);
or U2165 (N_2165,N_2081,N_2080);
nand U2166 (N_2166,N_2009,N_2027);
and U2167 (N_2167,N_2038,N_2089);
or U2168 (N_2168,N_2081,N_2046);
nor U2169 (N_2169,N_2074,N_2071);
nand U2170 (N_2170,N_2077,N_2007);
nor U2171 (N_2171,N_2010,N_2034);
nor U2172 (N_2172,N_2019,N_2029);
nand U2173 (N_2173,N_2032,N_2029);
or U2174 (N_2174,N_2010,N_2072);
nand U2175 (N_2175,N_2085,N_2094);
and U2176 (N_2176,N_2094,N_2052);
nand U2177 (N_2177,N_2043,N_2014);
xnor U2178 (N_2178,N_2062,N_2078);
nand U2179 (N_2179,N_2055,N_2029);
nor U2180 (N_2180,N_2005,N_2058);
nor U2181 (N_2181,N_2067,N_2032);
or U2182 (N_2182,N_2050,N_2012);
nor U2183 (N_2183,N_2099,N_2020);
nand U2184 (N_2184,N_2089,N_2033);
or U2185 (N_2185,N_2017,N_2082);
and U2186 (N_2186,N_2044,N_2020);
nand U2187 (N_2187,N_2081,N_2059);
nand U2188 (N_2188,N_2029,N_2063);
and U2189 (N_2189,N_2013,N_2051);
nor U2190 (N_2190,N_2068,N_2007);
and U2191 (N_2191,N_2047,N_2045);
xor U2192 (N_2192,N_2033,N_2026);
and U2193 (N_2193,N_2022,N_2067);
nor U2194 (N_2194,N_2079,N_2024);
or U2195 (N_2195,N_2001,N_2053);
and U2196 (N_2196,N_2055,N_2008);
nand U2197 (N_2197,N_2073,N_2095);
and U2198 (N_2198,N_2053,N_2098);
nor U2199 (N_2199,N_2072,N_2059);
and U2200 (N_2200,N_2112,N_2160);
or U2201 (N_2201,N_2130,N_2111);
nand U2202 (N_2202,N_2119,N_2166);
or U2203 (N_2203,N_2141,N_2115);
nor U2204 (N_2204,N_2151,N_2176);
xnor U2205 (N_2205,N_2197,N_2173);
nor U2206 (N_2206,N_2164,N_2172);
or U2207 (N_2207,N_2168,N_2132);
nor U2208 (N_2208,N_2110,N_2105);
or U2209 (N_2209,N_2149,N_2179);
nand U2210 (N_2210,N_2185,N_2100);
nand U2211 (N_2211,N_2193,N_2125);
nand U2212 (N_2212,N_2142,N_2107);
or U2213 (N_2213,N_2195,N_2163);
nand U2214 (N_2214,N_2194,N_2187);
and U2215 (N_2215,N_2180,N_2131);
nand U2216 (N_2216,N_2157,N_2121);
or U2217 (N_2217,N_2184,N_2103);
or U2218 (N_2218,N_2108,N_2134);
or U2219 (N_2219,N_2147,N_2138);
nand U2220 (N_2220,N_2183,N_2153);
or U2221 (N_2221,N_2128,N_2175);
or U2222 (N_2222,N_2189,N_2135);
xor U2223 (N_2223,N_2122,N_2145);
nand U2224 (N_2224,N_2120,N_2192);
nor U2225 (N_2225,N_2113,N_2102);
and U2226 (N_2226,N_2199,N_2154);
nand U2227 (N_2227,N_2140,N_2104);
nor U2228 (N_2228,N_2170,N_2123);
and U2229 (N_2229,N_2169,N_2178);
nand U2230 (N_2230,N_2106,N_2159);
or U2231 (N_2231,N_2136,N_2191);
xor U2232 (N_2232,N_2198,N_2137);
or U2233 (N_2233,N_2188,N_2116);
xnor U2234 (N_2234,N_2118,N_2158);
or U2235 (N_2235,N_2165,N_2127);
or U2236 (N_2236,N_2152,N_2114);
and U2237 (N_2237,N_2133,N_2196);
nor U2238 (N_2238,N_2129,N_2177);
nand U2239 (N_2239,N_2171,N_2148);
or U2240 (N_2240,N_2146,N_2167);
nor U2241 (N_2241,N_2150,N_2162);
and U2242 (N_2242,N_2124,N_2186);
or U2243 (N_2243,N_2126,N_2117);
nand U2244 (N_2244,N_2156,N_2144);
or U2245 (N_2245,N_2174,N_2155);
and U2246 (N_2246,N_2109,N_2161);
or U2247 (N_2247,N_2101,N_2190);
and U2248 (N_2248,N_2143,N_2182);
nor U2249 (N_2249,N_2181,N_2139);
or U2250 (N_2250,N_2145,N_2182);
or U2251 (N_2251,N_2159,N_2175);
nand U2252 (N_2252,N_2164,N_2110);
nand U2253 (N_2253,N_2175,N_2142);
xor U2254 (N_2254,N_2191,N_2122);
or U2255 (N_2255,N_2157,N_2156);
or U2256 (N_2256,N_2148,N_2175);
nor U2257 (N_2257,N_2180,N_2183);
or U2258 (N_2258,N_2111,N_2121);
or U2259 (N_2259,N_2177,N_2146);
and U2260 (N_2260,N_2191,N_2186);
nor U2261 (N_2261,N_2185,N_2142);
nor U2262 (N_2262,N_2198,N_2123);
and U2263 (N_2263,N_2116,N_2187);
or U2264 (N_2264,N_2127,N_2169);
nand U2265 (N_2265,N_2114,N_2179);
xor U2266 (N_2266,N_2155,N_2165);
xnor U2267 (N_2267,N_2152,N_2118);
and U2268 (N_2268,N_2120,N_2158);
nor U2269 (N_2269,N_2152,N_2186);
or U2270 (N_2270,N_2177,N_2189);
xor U2271 (N_2271,N_2161,N_2137);
nand U2272 (N_2272,N_2154,N_2120);
xnor U2273 (N_2273,N_2133,N_2113);
nand U2274 (N_2274,N_2139,N_2159);
xnor U2275 (N_2275,N_2143,N_2119);
nor U2276 (N_2276,N_2136,N_2110);
or U2277 (N_2277,N_2100,N_2132);
nor U2278 (N_2278,N_2179,N_2190);
or U2279 (N_2279,N_2126,N_2110);
nor U2280 (N_2280,N_2169,N_2124);
and U2281 (N_2281,N_2189,N_2164);
or U2282 (N_2282,N_2133,N_2195);
and U2283 (N_2283,N_2185,N_2147);
nand U2284 (N_2284,N_2139,N_2193);
or U2285 (N_2285,N_2146,N_2110);
nand U2286 (N_2286,N_2109,N_2163);
and U2287 (N_2287,N_2184,N_2186);
xnor U2288 (N_2288,N_2140,N_2123);
nand U2289 (N_2289,N_2114,N_2113);
nor U2290 (N_2290,N_2110,N_2151);
or U2291 (N_2291,N_2114,N_2163);
and U2292 (N_2292,N_2199,N_2177);
and U2293 (N_2293,N_2142,N_2164);
or U2294 (N_2294,N_2111,N_2157);
nand U2295 (N_2295,N_2162,N_2128);
nand U2296 (N_2296,N_2191,N_2155);
nor U2297 (N_2297,N_2174,N_2154);
and U2298 (N_2298,N_2125,N_2103);
and U2299 (N_2299,N_2179,N_2163);
xnor U2300 (N_2300,N_2269,N_2228);
nand U2301 (N_2301,N_2284,N_2201);
nand U2302 (N_2302,N_2275,N_2247);
nand U2303 (N_2303,N_2261,N_2217);
nand U2304 (N_2304,N_2258,N_2251);
nand U2305 (N_2305,N_2286,N_2290);
xor U2306 (N_2306,N_2214,N_2219);
or U2307 (N_2307,N_2240,N_2202);
nor U2308 (N_2308,N_2280,N_2227);
xor U2309 (N_2309,N_2253,N_2243);
or U2310 (N_2310,N_2279,N_2216);
and U2311 (N_2311,N_2212,N_2271);
nor U2312 (N_2312,N_2274,N_2207);
nand U2313 (N_2313,N_2236,N_2297);
and U2314 (N_2314,N_2278,N_2241);
xnor U2315 (N_2315,N_2237,N_2200);
and U2316 (N_2316,N_2235,N_2206);
or U2317 (N_2317,N_2230,N_2267);
and U2318 (N_2318,N_2287,N_2204);
or U2319 (N_2319,N_2218,N_2282);
nor U2320 (N_2320,N_2210,N_2215);
or U2321 (N_2321,N_2221,N_2283);
xor U2322 (N_2322,N_2222,N_2294);
nand U2323 (N_2323,N_2260,N_2263);
nor U2324 (N_2324,N_2203,N_2223);
or U2325 (N_2325,N_2295,N_2213);
xor U2326 (N_2326,N_2245,N_2239);
nor U2327 (N_2327,N_2266,N_2248);
and U2328 (N_2328,N_2211,N_2256);
nand U2329 (N_2329,N_2259,N_2234);
nand U2330 (N_2330,N_2264,N_2257);
or U2331 (N_2331,N_2233,N_2232);
nand U2332 (N_2332,N_2250,N_2268);
nand U2333 (N_2333,N_2298,N_2209);
nor U2334 (N_2334,N_2277,N_2296);
and U2335 (N_2335,N_2293,N_2289);
nor U2336 (N_2336,N_2276,N_2238);
nand U2337 (N_2337,N_2231,N_2273);
or U2338 (N_2338,N_2299,N_2285);
and U2339 (N_2339,N_2225,N_2244);
and U2340 (N_2340,N_2224,N_2270);
nand U2341 (N_2341,N_2229,N_2255);
and U2342 (N_2342,N_2242,N_2246);
or U2343 (N_2343,N_2226,N_2220);
nor U2344 (N_2344,N_2254,N_2288);
or U2345 (N_2345,N_2265,N_2281);
xor U2346 (N_2346,N_2252,N_2205);
xor U2347 (N_2347,N_2249,N_2208);
nor U2348 (N_2348,N_2262,N_2292);
xnor U2349 (N_2349,N_2291,N_2272);
nor U2350 (N_2350,N_2288,N_2292);
xnor U2351 (N_2351,N_2215,N_2265);
xnor U2352 (N_2352,N_2219,N_2213);
nor U2353 (N_2353,N_2248,N_2281);
xor U2354 (N_2354,N_2271,N_2292);
and U2355 (N_2355,N_2211,N_2276);
nand U2356 (N_2356,N_2293,N_2201);
nor U2357 (N_2357,N_2298,N_2259);
xnor U2358 (N_2358,N_2265,N_2277);
xor U2359 (N_2359,N_2216,N_2224);
nand U2360 (N_2360,N_2229,N_2298);
nor U2361 (N_2361,N_2276,N_2233);
or U2362 (N_2362,N_2227,N_2221);
xor U2363 (N_2363,N_2285,N_2221);
nand U2364 (N_2364,N_2273,N_2277);
and U2365 (N_2365,N_2209,N_2206);
xnor U2366 (N_2366,N_2254,N_2217);
and U2367 (N_2367,N_2211,N_2299);
and U2368 (N_2368,N_2257,N_2262);
nand U2369 (N_2369,N_2219,N_2290);
or U2370 (N_2370,N_2210,N_2289);
nor U2371 (N_2371,N_2249,N_2238);
or U2372 (N_2372,N_2234,N_2246);
nor U2373 (N_2373,N_2276,N_2245);
nand U2374 (N_2374,N_2265,N_2275);
or U2375 (N_2375,N_2231,N_2240);
nor U2376 (N_2376,N_2255,N_2242);
and U2377 (N_2377,N_2204,N_2249);
nand U2378 (N_2378,N_2246,N_2248);
or U2379 (N_2379,N_2212,N_2256);
or U2380 (N_2380,N_2217,N_2267);
and U2381 (N_2381,N_2231,N_2214);
or U2382 (N_2382,N_2295,N_2242);
or U2383 (N_2383,N_2249,N_2274);
or U2384 (N_2384,N_2202,N_2297);
and U2385 (N_2385,N_2258,N_2213);
or U2386 (N_2386,N_2236,N_2205);
and U2387 (N_2387,N_2210,N_2235);
nor U2388 (N_2388,N_2260,N_2275);
or U2389 (N_2389,N_2263,N_2294);
xor U2390 (N_2390,N_2236,N_2221);
and U2391 (N_2391,N_2262,N_2272);
xor U2392 (N_2392,N_2299,N_2266);
or U2393 (N_2393,N_2282,N_2209);
and U2394 (N_2394,N_2221,N_2228);
xor U2395 (N_2395,N_2260,N_2292);
nand U2396 (N_2396,N_2244,N_2294);
or U2397 (N_2397,N_2220,N_2265);
nand U2398 (N_2398,N_2204,N_2233);
xnor U2399 (N_2399,N_2259,N_2284);
nor U2400 (N_2400,N_2344,N_2323);
or U2401 (N_2401,N_2358,N_2331);
nand U2402 (N_2402,N_2312,N_2318);
nand U2403 (N_2403,N_2302,N_2354);
nand U2404 (N_2404,N_2337,N_2316);
nand U2405 (N_2405,N_2367,N_2388);
or U2406 (N_2406,N_2369,N_2315);
or U2407 (N_2407,N_2324,N_2334);
nand U2408 (N_2408,N_2327,N_2368);
xnor U2409 (N_2409,N_2384,N_2362);
nor U2410 (N_2410,N_2342,N_2374);
nand U2411 (N_2411,N_2320,N_2329);
xor U2412 (N_2412,N_2310,N_2373);
nand U2413 (N_2413,N_2305,N_2325);
nor U2414 (N_2414,N_2371,N_2366);
nor U2415 (N_2415,N_2393,N_2338);
and U2416 (N_2416,N_2333,N_2356);
and U2417 (N_2417,N_2359,N_2313);
nand U2418 (N_2418,N_2386,N_2349);
nor U2419 (N_2419,N_2340,N_2357);
xor U2420 (N_2420,N_2332,N_2372);
and U2421 (N_2421,N_2319,N_2370);
nor U2422 (N_2422,N_2317,N_2381);
or U2423 (N_2423,N_2378,N_2387);
nand U2424 (N_2424,N_2391,N_2360);
xnor U2425 (N_2425,N_2343,N_2383);
or U2426 (N_2426,N_2361,N_2301);
nand U2427 (N_2427,N_2365,N_2335);
and U2428 (N_2428,N_2326,N_2321);
and U2429 (N_2429,N_2314,N_2339);
nor U2430 (N_2430,N_2399,N_2300);
or U2431 (N_2431,N_2328,N_2382);
xor U2432 (N_2432,N_2308,N_2380);
nor U2433 (N_2433,N_2396,N_2306);
and U2434 (N_2434,N_2379,N_2377);
nand U2435 (N_2435,N_2304,N_2395);
and U2436 (N_2436,N_2322,N_2347);
or U2437 (N_2437,N_2351,N_2398);
and U2438 (N_2438,N_2355,N_2353);
and U2439 (N_2439,N_2392,N_2363);
nor U2440 (N_2440,N_2352,N_2346);
nor U2441 (N_2441,N_2309,N_2311);
xnor U2442 (N_2442,N_2394,N_2307);
nand U2443 (N_2443,N_2350,N_2390);
nor U2444 (N_2444,N_2303,N_2385);
xor U2445 (N_2445,N_2345,N_2375);
nand U2446 (N_2446,N_2341,N_2389);
xnor U2447 (N_2447,N_2364,N_2336);
and U2448 (N_2448,N_2376,N_2397);
or U2449 (N_2449,N_2348,N_2330);
nor U2450 (N_2450,N_2318,N_2387);
or U2451 (N_2451,N_2316,N_2309);
and U2452 (N_2452,N_2355,N_2356);
nand U2453 (N_2453,N_2349,N_2304);
nand U2454 (N_2454,N_2342,N_2380);
nand U2455 (N_2455,N_2330,N_2370);
or U2456 (N_2456,N_2398,N_2363);
and U2457 (N_2457,N_2366,N_2379);
nand U2458 (N_2458,N_2356,N_2393);
nor U2459 (N_2459,N_2370,N_2389);
and U2460 (N_2460,N_2347,N_2345);
nor U2461 (N_2461,N_2341,N_2346);
nand U2462 (N_2462,N_2367,N_2300);
xor U2463 (N_2463,N_2381,N_2362);
and U2464 (N_2464,N_2361,N_2318);
nand U2465 (N_2465,N_2372,N_2320);
nor U2466 (N_2466,N_2335,N_2315);
xnor U2467 (N_2467,N_2328,N_2377);
nor U2468 (N_2468,N_2327,N_2300);
xor U2469 (N_2469,N_2378,N_2304);
xnor U2470 (N_2470,N_2345,N_2368);
and U2471 (N_2471,N_2337,N_2366);
or U2472 (N_2472,N_2325,N_2354);
nor U2473 (N_2473,N_2374,N_2309);
xor U2474 (N_2474,N_2366,N_2353);
or U2475 (N_2475,N_2373,N_2341);
nor U2476 (N_2476,N_2327,N_2369);
and U2477 (N_2477,N_2313,N_2355);
nand U2478 (N_2478,N_2332,N_2329);
nor U2479 (N_2479,N_2334,N_2384);
or U2480 (N_2480,N_2395,N_2370);
nand U2481 (N_2481,N_2327,N_2388);
nor U2482 (N_2482,N_2334,N_2342);
or U2483 (N_2483,N_2348,N_2316);
and U2484 (N_2484,N_2393,N_2334);
nor U2485 (N_2485,N_2376,N_2367);
nand U2486 (N_2486,N_2314,N_2363);
or U2487 (N_2487,N_2396,N_2360);
nand U2488 (N_2488,N_2337,N_2317);
nor U2489 (N_2489,N_2314,N_2313);
nor U2490 (N_2490,N_2387,N_2365);
and U2491 (N_2491,N_2366,N_2367);
and U2492 (N_2492,N_2319,N_2328);
and U2493 (N_2493,N_2325,N_2360);
or U2494 (N_2494,N_2305,N_2323);
nand U2495 (N_2495,N_2380,N_2333);
or U2496 (N_2496,N_2390,N_2336);
xnor U2497 (N_2497,N_2305,N_2327);
or U2498 (N_2498,N_2355,N_2325);
or U2499 (N_2499,N_2366,N_2374);
nand U2500 (N_2500,N_2433,N_2420);
nand U2501 (N_2501,N_2411,N_2463);
xnor U2502 (N_2502,N_2473,N_2405);
and U2503 (N_2503,N_2404,N_2446);
nor U2504 (N_2504,N_2493,N_2452);
or U2505 (N_2505,N_2441,N_2426);
nand U2506 (N_2506,N_2414,N_2478);
xor U2507 (N_2507,N_2460,N_2477);
and U2508 (N_2508,N_2412,N_2455);
and U2509 (N_2509,N_2410,N_2436);
nand U2510 (N_2510,N_2445,N_2431);
nand U2511 (N_2511,N_2415,N_2444);
and U2512 (N_2512,N_2403,N_2475);
xnor U2513 (N_2513,N_2497,N_2498);
and U2514 (N_2514,N_2494,N_2458);
and U2515 (N_2515,N_2491,N_2425);
xnor U2516 (N_2516,N_2489,N_2454);
nor U2517 (N_2517,N_2456,N_2439);
or U2518 (N_2518,N_2453,N_2464);
and U2519 (N_2519,N_2499,N_2479);
nor U2520 (N_2520,N_2407,N_2434);
xnor U2521 (N_2521,N_2484,N_2486);
xnor U2522 (N_2522,N_2416,N_2438);
nand U2523 (N_2523,N_2465,N_2481);
or U2524 (N_2524,N_2443,N_2450);
or U2525 (N_2525,N_2474,N_2440);
nand U2526 (N_2526,N_2409,N_2490);
nand U2527 (N_2527,N_2422,N_2429);
nor U2528 (N_2528,N_2451,N_2472);
and U2529 (N_2529,N_2496,N_2402);
nand U2530 (N_2530,N_2483,N_2448);
nand U2531 (N_2531,N_2480,N_2449);
nor U2532 (N_2532,N_2488,N_2432);
or U2533 (N_2533,N_2424,N_2468);
nand U2534 (N_2534,N_2428,N_2461);
nand U2535 (N_2535,N_2401,N_2482);
and U2536 (N_2536,N_2406,N_2469);
nor U2537 (N_2537,N_2430,N_2487);
or U2538 (N_2538,N_2447,N_2462);
and U2539 (N_2539,N_2413,N_2417);
or U2540 (N_2540,N_2485,N_2470);
or U2541 (N_2541,N_2442,N_2471);
nand U2542 (N_2542,N_2418,N_2459);
and U2543 (N_2543,N_2457,N_2466);
nor U2544 (N_2544,N_2435,N_2423);
nand U2545 (N_2545,N_2427,N_2421);
nor U2546 (N_2546,N_2408,N_2467);
and U2547 (N_2547,N_2476,N_2419);
or U2548 (N_2548,N_2400,N_2492);
or U2549 (N_2549,N_2495,N_2437);
nand U2550 (N_2550,N_2488,N_2459);
xnor U2551 (N_2551,N_2453,N_2452);
or U2552 (N_2552,N_2439,N_2468);
or U2553 (N_2553,N_2413,N_2401);
xor U2554 (N_2554,N_2418,N_2461);
nand U2555 (N_2555,N_2421,N_2440);
xor U2556 (N_2556,N_2430,N_2404);
nand U2557 (N_2557,N_2486,N_2499);
nand U2558 (N_2558,N_2448,N_2419);
xor U2559 (N_2559,N_2467,N_2400);
and U2560 (N_2560,N_2418,N_2456);
or U2561 (N_2561,N_2449,N_2431);
nor U2562 (N_2562,N_2415,N_2408);
nor U2563 (N_2563,N_2440,N_2413);
or U2564 (N_2564,N_2461,N_2457);
nor U2565 (N_2565,N_2495,N_2423);
nand U2566 (N_2566,N_2465,N_2434);
nand U2567 (N_2567,N_2411,N_2432);
and U2568 (N_2568,N_2415,N_2409);
and U2569 (N_2569,N_2406,N_2419);
nand U2570 (N_2570,N_2408,N_2477);
xnor U2571 (N_2571,N_2424,N_2426);
nand U2572 (N_2572,N_2461,N_2443);
or U2573 (N_2573,N_2406,N_2449);
or U2574 (N_2574,N_2482,N_2487);
nor U2575 (N_2575,N_2456,N_2489);
and U2576 (N_2576,N_2438,N_2442);
or U2577 (N_2577,N_2439,N_2464);
or U2578 (N_2578,N_2438,N_2424);
or U2579 (N_2579,N_2416,N_2403);
nand U2580 (N_2580,N_2482,N_2418);
nand U2581 (N_2581,N_2487,N_2446);
or U2582 (N_2582,N_2441,N_2465);
or U2583 (N_2583,N_2420,N_2415);
or U2584 (N_2584,N_2479,N_2472);
and U2585 (N_2585,N_2467,N_2479);
nand U2586 (N_2586,N_2457,N_2405);
nor U2587 (N_2587,N_2406,N_2473);
or U2588 (N_2588,N_2412,N_2418);
and U2589 (N_2589,N_2404,N_2492);
or U2590 (N_2590,N_2405,N_2440);
or U2591 (N_2591,N_2445,N_2436);
and U2592 (N_2592,N_2401,N_2418);
nor U2593 (N_2593,N_2419,N_2463);
and U2594 (N_2594,N_2402,N_2412);
or U2595 (N_2595,N_2470,N_2422);
nor U2596 (N_2596,N_2447,N_2482);
xnor U2597 (N_2597,N_2435,N_2425);
and U2598 (N_2598,N_2489,N_2471);
nor U2599 (N_2599,N_2485,N_2499);
and U2600 (N_2600,N_2519,N_2507);
nor U2601 (N_2601,N_2589,N_2500);
and U2602 (N_2602,N_2503,N_2599);
and U2603 (N_2603,N_2542,N_2540);
xor U2604 (N_2604,N_2593,N_2508);
xnor U2605 (N_2605,N_2578,N_2521);
and U2606 (N_2606,N_2547,N_2597);
or U2607 (N_2607,N_2553,N_2585);
nor U2608 (N_2608,N_2509,N_2517);
nand U2609 (N_2609,N_2526,N_2534);
and U2610 (N_2610,N_2587,N_2568);
or U2611 (N_2611,N_2551,N_2576);
nor U2612 (N_2612,N_2506,N_2504);
or U2613 (N_2613,N_2548,N_2567);
nand U2614 (N_2614,N_2592,N_2560);
nor U2615 (N_2615,N_2571,N_2586);
nand U2616 (N_2616,N_2535,N_2528);
and U2617 (N_2617,N_2596,N_2533);
nor U2618 (N_2618,N_2583,N_2538);
or U2619 (N_2619,N_2550,N_2524);
or U2620 (N_2620,N_2545,N_2544);
or U2621 (N_2621,N_2523,N_2570);
xor U2622 (N_2622,N_2565,N_2522);
xor U2623 (N_2623,N_2595,N_2525);
and U2624 (N_2624,N_2527,N_2543);
or U2625 (N_2625,N_2520,N_2588);
nor U2626 (N_2626,N_2505,N_2564);
nor U2627 (N_2627,N_2511,N_2584);
nand U2628 (N_2628,N_2552,N_2573);
or U2629 (N_2629,N_2502,N_2516);
or U2630 (N_2630,N_2537,N_2510);
nor U2631 (N_2631,N_2558,N_2577);
nor U2632 (N_2632,N_2514,N_2546);
nor U2633 (N_2633,N_2532,N_2572);
and U2634 (N_2634,N_2557,N_2559);
and U2635 (N_2635,N_2579,N_2562);
xnor U2636 (N_2636,N_2590,N_2575);
nand U2637 (N_2637,N_2536,N_2512);
nand U2638 (N_2638,N_2594,N_2582);
nand U2639 (N_2639,N_2539,N_2591);
nor U2640 (N_2640,N_2554,N_2529);
or U2641 (N_2641,N_2518,N_2549);
nor U2642 (N_2642,N_2574,N_2566);
xnor U2643 (N_2643,N_2555,N_2598);
nand U2644 (N_2644,N_2501,N_2581);
and U2645 (N_2645,N_2531,N_2580);
and U2646 (N_2646,N_2515,N_2563);
nor U2647 (N_2647,N_2513,N_2561);
and U2648 (N_2648,N_2556,N_2541);
nand U2649 (N_2649,N_2569,N_2530);
nand U2650 (N_2650,N_2543,N_2553);
and U2651 (N_2651,N_2579,N_2509);
nor U2652 (N_2652,N_2535,N_2594);
nor U2653 (N_2653,N_2592,N_2570);
nor U2654 (N_2654,N_2591,N_2538);
nor U2655 (N_2655,N_2563,N_2555);
nand U2656 (N_2656,N_2591,N_2515);
nor U2657 (N_2657,N_2527,N_2587);
and U2658 (N_2658,N_2587,N_2556);
nor U2659 (N_2659,N_2562,N_2599);
and U2660 (N_2660,N_2511,N_2510);
or U2661 (N_2661,N_2570,N_2557);
nor U2662 (N_2662,N_2542,N_2577);
nor U2663 (N_2663,N_2589,N_2520);
or U2664 (N_2664,N_2589,N_2596);
nor U2665 (N_2665,N_2550,N_2578);
or U2666 (N_2666,N_2562,N_2573);
and U2667 (N_2667,N_2550,N_2528);
nand U2668 (N_2668,N_2504,N_2568);
and U2669 (N_2669,N_2531,N_2570);
nor U2670 (N_2670,N_2572,N_2512);
nand U2671 (N_2671,N_2568,N_2541);
nand U2672 (N_2672,N_2569,N_2518);
nand U2673 (N_2673,N_2555,N_2519);
nand U2674 (N_2674,N_2520,N_2518);
and U2675 (N_2675,N_2574,N_2575);
nor U2676 (N_2676,N_2545,N_2550);
nand U2677 (N_2677,N_2555,N_2568);
nor U2678 (N_2678,N_2500,N_2575);
nor U2679 (N_2679,N_2540,N_2538);
and U2680 (N_2680,N_2522,N_2582);
nor U2681 (N_2681,N_2539,N_2567);
or U2682 (N_2682,N_2558,N_2501);
and U2683 (N_2683,N_2569,N_2563);
nand U2684 (N_2684,N_2545,N_2530);
and U2685 (N_2685,N_2541,N_2538);
or U2686 (N_2686,N_2594,N_2526);
nand U2687 (N_2687,N_2531,N_2507);
or U2688 (N_2688,N_2566,N_2547);
or U2689 (N_2689,N_2518,N_2536);
and U2690 (N_2690,N_2572,N_2527);
and U2691 (N_2691,N_2554,N_2566);
and U2692 (N_2692,N_2503,N_2570);
or U2693 (N_2693,N_2515,N_2541);
and U2694 (N_2694,N_2546,N_2556);
and U2695 (N_2695,N_2521,N_2546);
and U2696 (N_2696,N_2566,N_2596);
or U2697 (N_2697,N_2552,N_2544);
xor U2698 (N_2698,N_2565,N_2562);
nor U2699 (N_2699,N_2589,N_2592);
nor U2700 (N_2700,N_2627,N_2637);
or U2701 (N_2701,N_2669,N_2690);
and U2702 (N_2702,N_2611,N_2648);
nand U2703 (N_2703,N_2664,N_2677);
xnor U2704 (N_2704,N_2617,N_2675);
and U2705 (N_2705,N_2672,N_2624);
and U2706 (N_2706,N_2629,N_2695);
xnor U2707 (N_2707,N_2630,N_2612);
nand U2708 (N_2708,N_2623,N_2619);
or U2709 (N_2709,N_2602,N_2600);
or U2710 (N_2710,N_2625,N_2651);
or U2711 (N_2711,N_2604,N_2649);
nor U2712 (N_2712,N_2616,N_2621);
or U2713 (N_2713,N_2683,N_2653);
or U2714 (N_2714,N_2628,N_2606);
and U2715 (N_2715,N_2603,N_2681);
or U2716 (N_2716,N_2692,N_2697);
nor U2717 (N_2717,N_2643,N_2631);
and U2718 (N_2718,N_2635,N_2607);
or U2719 (N_2719,N_2679,N_2608);
nor U2720 (N_2720,N_2691,N_2696);
and U2721 (N_2721,N_2666,N_2626);
nor U2722 (N_2722,N_2640,N_2671);
nand U2723 (N_2723,N_2698,N_2661);
and U2724 (N_2724,N_2656,N_2674);
and U2725 (N_2725,N_2670,N_2610);
and U2726 (N_2726,N_2657,N_2614);
and U2727 (N_2727,N_2678,N_2658);
nand U2728 (N_2728,N_2673,N_2647);
and U2729 (N_2729,N_2699,N_2668);
nand U2730 (N_2730,N_2663,N_2613);
nor U2731 (N_2731,N_2667,N_2620);
and U2732 (N_2732,N_2636,N_2693);
nand U2733 (N_2733,N_2689,N_2644);
nor U2734 (N_2734,N_2684,N_2659);
and U2735 (N_2735,N_2660,N_2601);
nor U2736 (N_2736,N_2633,N_2687);
or U2737 (N_2737,N_2646,N_2682);
nor U2738 (N_2738,N_2680,N_2652);
nand U2739 (N_2739,N_2632,N_2676);
nand U2740 (N_2740,N_2654,N_2686);
or U2741 (N_2741,N_2665,N_2685);
nand U2742 (N_2742,N_2694,N_2639);
or U2743 (N_2743,N_2605,N_2650);
or U2744 (N_2744,N_2618,N_2622);
and U2745 (N_2745,N_2688,N_2642);
or U2746 (N_2746,N_2615,N_2609);
or U2747 (N_2747,N_2655,N_2641);
nand U2748 (N_2748,N_2645,N_2662);
or U2749 (N_2749,N_2638,N_2634);
or U2750 (N_2750,N_2630,N_2615);
xnor U2751 (N_2751,N_2693,N_2611);
and U2752 (N_2752,N_2613,N_2618);
nor U2753 (N_2753,N_2606,N_2659);
xnor U2754 (N_2754,N_2635,N_2636);
nor U2755 (N_2755,N_2690,N_2699);
or U2756 (N_2756,N_2673,N_2634);
nor U2757 (N_2757,N_2692,N_2672);
nand U2758 (N_2758,N_2651,N_2692);
or U2759 (N_2759,N_2638,N_2678);
xor U2760 (N_2760,N_2635,N_2646);
or U2761 (N_2761,N_2613,N_2668);
xnor U2762 (N_2762,N_2617,N_2614);
or U2763 (N_2763,N_2677,N_2699);
and U2764 (N_2764,N_2693,N_2647);
xnor U2765 (N_2765,N_2618,N_2663);
xnor U2766 (N_2766,N_2654,N_2649);
and U2767 (N_2767,N_2648,N_2699);
nand U2768 (N_2768,N_2602,N_2665);
and U2769 (N_2769,N_2629,N_2672);
nand U2770 (N_2770,N_2691,N_2683);
nor U2771 (N_2771,N_2683,N_2658);
nor U2772 (N_2772,N_2607,N_2655);
and U2773 (N_2773,N_2698,N_2684);
nand U2774 (N_2774,N_2623,N_2678);
nor U2775 (N_2775,N_2602,N_2697);
or U2776 (N_2776,N_2624,N_2692);
nor U2777 (N_2777,N_2659,N_2607);
or U2778 (N_2778,N_2676,N_2675);
nor U2779 (N_2779,N_2621,N_2618);
nand U2780 (N_2780,N_2622,N_2663);
nand U2781 (N_2781,N_2622,N_2645);
nand U2782 (N_2782,N_2689,N_2605);
and U2783 (N_2783,N_2603,N_2682);
and U2784 (N_2784,N_2668,N_2689);
or U2785 (N_2785,N_2682,N_2607);
and U2786 (N_2786,N_2618,N_2684);
xor U2787 (N_2787,N_2636,N_2631);
nor U2788 (N_2788,N_2651,N_2694);
nor U2789 (N_2789,N_2610,N_2661);
or U2790 (N_2790,N_2679,N_2694);
nand U2791 (N_2791,N_2640,N_2688);
nand U2792 (N_2792,N_2643,N_2674);
nor U2793 (N_2793,N_2681,N_2624);
nand U2794 (N_2794,N_2633,N_2683);
and U2795 (N_2795,N_2628,N_2674);
nand U2796 (N_2796,N_2615,N_2661);
xnor U2797 (N_2797,N_2631,N_2691);
or U2798 (N_2798,N_2602,N_2604);
nor U2799 (N_2799,N_2643,N_2626);
nor U2800 (N_2800,N_2738,N_2702);
nand U2801 (N_2801,N_2750,N_2701);
nand U2802 (N_2802,N_2770,N_2743);
nand U2803 (N_2803,N_2765,N_2709);
nand U2804 (N_2804,N_2749,N_2703);
xor U2805 (N_2805,N_2714,N_2780);
or U2806 (N_2806,N_2766,N_2754);
nor U2807 (N_2807,N_2700,N_2721);
and U2808 (N_2808,N_2711,N_2759);
or U2809 (N_2809,N_2725,N_2761);
nand U2810 (N_2810,N_2723,N_2758);
and U2811 (N_2811,N_2720,N_2742);
or U2812 (N_2812,N_2798,N_2708);
or U2813 (N_2813,N_2713,N_2799);
nor U2814 (N_2814,N_2793,N_2767);
and U2815 (N_2815,N_2707,N_2717);
nor U2816 (N_2816,N_2736,N_2737);
and U2817 (N_2817,N_2791,N_2771);
nor U2818 (N_2818,N_2739,N_2775);
and U2819 (N_2819,N_2779,N_2731);
and U2820 (N_2820,N_2728,N_2704);
nand U2821 (N_2821,N_2788,N_2747);
nor U2822 (N_2822,N_2716,N_2741);
or U2823 (N_2823,N_2794,N_2782);
nor U2824 (N_2824,N_2751,N_2727);
and U2825 (N_2825,N_2774,N_2730);
xnor U2826 (N_2826,N_2735,N_2789);
nor U2827 (N_2827,N_2769,N_2722);
nand U2828 (N_2828,N_2785,N_2796);
nand U2829 (N_2829,N_2724,N_2729);
and U2830 (N_2830,N_2712,N_2746);
and U2831 (N_2831,N_2792,N_2734);
or U2832 (N_2832,N_2763,N_2773);
or U2833 (N_2833,N_2760,N_2795);
and U2834 (N_2834,N_2744,N_2783);
nand U2835 (N_2835,N_2710,N_2784);
nand U2836 (N_2836,N_2733,N_2757);
nor U2837 (N_2837,N_2797,N_2776);
nand U2838 (N_2838,N_2755,N_2756);
or U2839 (N_2839,N_2752,N_2768);
and U2840 (N_2840,N_2762,N_2732);
nand U2841 (N_2841,N_2787,N_2777);
xnor U2842 (N_2842,N_2718,N_2740);
and U2843 (N_2843,N_2745,N_2778);
and U2844 (N_2844,N_2764,N_2706);
nor U2845 (N_2845,N_2748,N_2705);
or U2846 (N_2846,N_2781,N_2772);
or U2847 (N_2847,N_2786,N_2753);
and U2848 (N_2848,N_2715,N_2790);
nor U2849 (N_2849,N_2719,N_2726);
and U2850 (N_2850,N_2712,N_2797);
or U2851 (N_2851,N_2704,N_2761);
nand U2852 (N_2852,N_2799,N_2753);
nand U2853 (N_2853,N_2722,N_2700);
nand U2854 (N_2854,N_2764,N_2775);
xor U2855 (N_2855,N_2750,N_2765);
or U2856 (N_2856,N_2723,N_2700);
or U2857 (N_2857,N_2796,N_2734);
nor U2858 (N_2858,N_2794,N_2701);
or U2859 (N_2859,N_2720,N_2786);
or U2860 (N_2860,N_2732,N_2778);
nand U2861 (N_2861,N_2771,N_2702);
and U2862 (N_2862,N_2727,N_2784);
or U2863 (N_2863,N_2771,N_2709);
xor U2864 (N_2864,N_2776,N_2714);
xor U2865 (N_2865,N_2731,N_2715);
and U2866 (N_2866,N_2748,N_2788);
nor U2867 (N_2867,N_2709,N_2779);
or U2868 (N_2868,N_2769,N_2733);
or U2869 (N_2869,N_2780,N_2781);
and U2870 (N_2870,N_2724,N_2717);
nor U2871 (N_2871,N_2789,N_2788);
or U2872 (N_2872,N_2739,N_2756);
nor U2873 (N_2873,N_2736,N_2764);
nand U2874 (N_2874,N_2770,N_2752);
nor U2875 (N_2875,N_2737,N_2760);
nor U2876 (N_2876,N_2761,N_2706);
xnor U2877 (N_2877,N_2751,N_2739);
and U2878 (N_2878,N_2741,N_2765);
nor U2879 (N_2879,N_2762,N_2709);
or U2880 (N_2880,N_2704,N_2729);
or U2881 (N_2881,N_2753,N_2797);
nor U2882 (N_2882,N_2718,N_2754);
nand U2883 (N_2883,N_2721,N_2776);
xnor U2884 (N_2884,N_2734,N_2742);
and U2885 (N_2885,N_2742,N_2703);
and U2886 (N_2886,N_2704,N_2782);
nor U2887 (N_2887,N_2725,N_2709);
or U2888 (N_2888,N_2784,N_2733);
and U2889 (N_2889,N_2703,N_2712);
and U2890 (N_2890,N_2778,N_2742);
or U2891 (N_2891,N_2744,N_2702);
and U2892 (N_2892,N_2786,N_2768);
nor U2893 (N_2893,N_2719,N_2727);
nand U2894 (N_2894,N_2743,N_2704);
nand U2895 (N_2895,N_2754,N_2787);
nand U2896 (N_2896,N_2745,N_2729);
nor U2897 (N_2897,N_2703,N_2767);
or U2898 (N_2898,N_2792,N_2760);
nor U2899 (N_2899,N_2745,N_2705);
nor U2900 (N_2900,N_2858,N_2855);
xnor U2901 (N_2901,N_2893,N_2811);
and U2902 (N_2902,N_2806,N_2842);
nand U2903 (N_2903,N_2882,N_2853);
xor U2904 (N_2904,N_2833,N_2836);
and U2905 (N_2905,N_2895,N_2879);
or U2906 (N_2906,N_2897,N_2835);
nor U2907 (N_2907,N_2838,N_2816);
or U2908 (N_2908,N_2870,N_2880);
nand U2909 (N_2909,N_2875,N_2898);
nor U2910 (N_2910,N_2801,N_2844);
nor U2911 (N_2911,N_2871,N_2802);
xor U2912 (N_2912,N_2837,N_2843);
nand U2913 (N_2913,N_2864,N_2817);
nand U2914 (N_2914,N_2847,N_2877);
nor U2915 (N_2915,N_2803,N_2800);
nand U2916 (N_2916,N_2820,N_2881);
nand U2917 (N_2917,N_2830,N_2822);
or U2918 (N_2918,N_2831,N_2884);
xor U2919 (N_2919,N_2872,N_2899);
nor U2920 (N_2920,N_2805,N_2839);
nand U2921 (N_2921,N_2846,N_2865);
or U2922 (N_2922,N_2845,N_2825);
and U2923 (N_2923,N_2851,N_2834);
or U2924 (N_2924,N_2857,N_2890);
nand U2925 (N_2925,N_2894,N_2824);
nand U2926 (N_2926,N_2827,N_2814);
nand U2927 (N_2927,N_2863,N_2854);
nand U2928 (N_2928,N_2852,N_2892);
nor U2929 (N_2929,N_2873,N_2856);
and U2930 (N_2930,N_2886,N_2821);
xor U2931 (N_2931,N_2815,N_2818);
nor U2932 (N_2932,N_2887,N_2850);
nand U2933 (N_2933,N_2888,N_2859);
nor U2934 (N_2934,N_2826,N_2885);
and U2935 (N_2935,N_2849,N_2878);
and U2936 (N_2936,N_2808,N_2841);
or U2937 (N_2937,N_2861,N_2889);
and U2938 (N_2938,N_2868,N_2896);
nand U2939 (N_2939,N_2807,N_2876);
xnor U2940 (N_2940,N_2862,N_2869);
nand U2941 (N_2941,N_2867,N_2848);
or U2942 (N_2942,N_2832,N_2812);
nand U2943 (N_2943,N_2866,N_2860);
xor U2944 (N_2944,N_2891,N_2883);
nor U2945 (N_2945,N_2809,N_2819);
nor U2946 (N_2946,N_2840,N_2804);
and U2947 (N_2947,N_2810,N_2828);
nor U2948 (N_2948,N_2813,N_2823);
nand U2949 (N_2949,N_2829,N_2874);
and U2950 (N_2950,N_2894,N_2822);
nor U2951 (N_2951,N_2876,N_2824);
xnor U2952 (N_2952,N_2800,N_2842);
nor U2953 (N_2953,N_2877,N_2802);
xor U2954 (N_2954,N_2819,N_2889);
and U2955 (N_2955,N_2838,N_2886);
nor U2956 (N_2956,N_2849,N_2885);
nand U2957 (N_2957,N_2887,N_2839);
nand U2958 (N_2958,N_2831,N_2838);
nor U2959 (N_2959,N_2869,N_2839);
or U2960 (N_2960,N_2870,N_2851);
nand U2961 (N_2961,N_2800,N_2824);
nand U2962 (N_2962,N_2878,N_2832);
and U2963 (N_2963,N_2845,N_2862);
xor U2964 (N_2964,N_2874,N_2814);
and U2965 (N_2965,N_2885,N_2817);
nor U2966 (N_2966,N_2899,N_2826);
and U2967 (N_2967,N_2832,N_2862);
or U2968 (N_2968,N_2864,N_2836);
nand U2969 (N_2969,N_2802,N_2849);
nor U2970 (N_2970,N_2818,N_2810);
nor U2971 (N_2971,N_2818,N_2843);
or U2972 (N_2972,N_2873,N_2874);
nand U2973 (N_2973,N_2831,N_2851);
nand U2974 (N_2974,N_2827,N_2812);
nor U2975 (N_2975,N_2885,N_2813);
nand U2976 (N_2976,N_2895,N_2857);
nand U2977 (N_2977,N_2880,N_2835);
xnor U2978 (N_2978,N_2848,N_2845);
or U2979 (N_2979,N_2849,N_2898);
nor U2980 (N_2980,N_2860,N_2805);
and U2981 (N_2981,N_2829,N_2842);
and U2982 (N_2982,N_2809,N_2827);
or U2983 (N_2983,N_2854,N_2828);
nor U2984 (N_2984,N_2890,N_2847);
nor U2985 (N_2985,N_2828,N_2829);
and U2986 (N_2986,N_2810,N_2826);
and U2987 (N_2987,N_2808,N_2885);
or U2988 (N_2988,N_2828,N_2874);
or U2989 (N_2989,N_2864,N_2846);
or U2990 (N_2990,N_2843,N_2865);
xnor U2991 (N_2991,N_2846,N_2845);
xnor U2992 (N_2992,N_2888,N_2845);
nor U2993 (N_2993,N_2847,N_2821);
and U2994 (N_2994,N_2806,N_2896);
or U2995 (N_2995,N_2862,N_2898);
nor U2996 (N_2996,N_2836,N_2839);
nor U2997 (N_2997,N_2828,N_2891);
xnor U2998 (N_2998,N_2879,N_2813);
and U2999 (N_2999,N_2896,N_2818);
nand UO_0 (O_0,N_2916,N_2948);
nor UO_1 (O_1,N_2991,N_2951);
nor UO_2 (O_2,N_2925,N_2929);
nor UO_3 (O_3,N_2968,N_2955);
and UO_4 (O_4,N_2958,N_2939);
nand UO_5 (O_5,N_2972,N_2946);
or UO_6 (O_6,N_2982,N_2902);
nor UO_7 (O_7,N_2967,N_2927);
and UO_8 (O_8,N_2986,N_2910);
or UO_9 (O_9,N_2938,N_2957);
or UO_10 (O_10,N_2935,N_2974);
nor UO_11 (O_11,N_2942,N_2926);
and UO_12 (O_12,N_2922,N_2953);
nand UO_13 (O_13,N_2970,N_2941);
or UO_14 (O_14,N_2940,N_2990);
or UO_15 (O_15,N_2983,N_2900);
or UO_16 (O_16,N_2918,N_2949);
and UO_17 (O_17,N_2979,N_2901);
nor UO_18 (O_18,N_2952,N_2989);
or UO_19 (O_19,N_2903,N_2971);
and UO_20 (O_20,N_2965,N_2944);
or UO_21 (O_21,N_2998,N_2947);
nand UO_22 (O_22,N_2924,N_2907);
nor UO_23 (O_23,N_2912,N_2928);
nand UO_24 (O_24,N_2999,N_2936);
or UO_25 (O_25,N_2963,N_2913);
nand UO_26 (O_26,N_2937,N_2995);
or UO_27 (O_27,N_2993,N_2973);
nor UO_28 (O_28,N_2933,N_2976);
xor UO_29 (O_29,N_2988,N_2992);
nor UO_30 (O_30,N_2978,N_2956);
nand UO_31 (O_31,N_2985,N_2906);
nand UO_32 (O_32,N_2911,N_2969);
and UO_33 (O_33,N_2914,N_2934);
or UO_34 (O_34,N_2996,N_2962);
and UO_35 (O_35,N_2931,N_2921);
nand UO_36 (O_36,N_2960,N_2950);
and UO_37 (O_37,N_2977,N_2975);
nand UO_38 (O_38,N_2945,N_2930);
and UO_39 (O_39,N_2908,N_2917);
or UO_40 (O_40,N_2961,N_2915);
or UO_41 (O_41,N_2919,N_2966);
nor UO_42 (O_42,N_2904,N_2980);
nand UO_43 (O_43,N_2981,N_2905);
nor UO_44 (O_44,N_2923,N_2954);
or UO_45 (O_45,N_2964,N_2920);
or UO_46 (O_46,N_2987,N_2994);
and UO_47 (O_47,N_2932,N_2909);
nand UO_48 (O_48,N_2997,N_2943);
nor UO_49 (O_49,N_2984,N_2959);
and UO_50 (O_50,N_2956,N_2996);
or UO_51 (O_51,N_2946,N_2930);
xnor UO_52 (O_52,N_2944,N_2912);
nand UO_53 (O_53,N_2970,N_2909);
xnor UO_54 (O_54,N_2944,N_2940);
nand UO_55 (O_55,N_2983,N_2990);
or UO_56 (O_56,N_2935,N_2961);
or UO_57 (O_57,N_2991,N_2986);
nand UO_58 (O_58,N_2909,N_2960);
nor UO_59 (O_59,N_2916,N_2908);
nand UO_60 (O_60,N_2935,N_2952);
nor UO_61 (O_61,N_2920,N_2901);
nand UO_62 (O_62,N_2912,N_2915);
or UO_63 (O_63,N_2938,N_2981);
nor UO_64 (O_64,N_2988,N_2976);
or UO_65 (O_65,N_2961,N_2972);
or UO_66 (O_66,N_2915,N_2921);
or UO_67 (O_67,N_2994,N_2940);
xnor UO_68 (O_68,N_2913,N_2930);
nand UO_69 (O_69,N_2942,N_2978);
and UO_70 (O_70,N_2973,N_2946);
nand UO_71 (O_71,N_2919,N_2909);
or UO_72 (O_72,N_2987,N_2949);
nand UO_73 (O_73,N_2935,N_2950);
and UO_74 (O_74,N_2983,N_2951);
and UO_75 (O_75,N_2937,N_2956);
xor UO_76 (O_76,N_2903,N_2950);
nand UO_77 (O_77,N_2979,N_2987);
nor UO_78 (O_78,N_2940,N_2912);
nand UO_79 (O_79,N_2979,N_2923);
or UO_80 (O_80,N_2916,N_2974);
and UO_81 (O_81,N_2950,N_2991);
and UO_82 (O_82,N_2960,N_2985);
and UO_83 (O_83,N_2988,N_2987);
and UO_84 (O_84,N_2975,N_2952);
nor UO_85 (O_85,N_2966,N_2906);
nand UO_86 (O_86,N_2968,N_2906);
xor UO_87 (O_87,N_2931,N_2985);
nand UO_88 (O_88,N_2958,N_2988);
nand UO_89 (O_89,N_2946,N_2959);
nor UO_90 (O_90,N_2992,N_2916);
and UO_91 (O_91,N_2956,N_2967);
nor UO_92 (O_92,N_2904,N_2984);
and UO_93 (O_93,N_2911,N_2925);
or UO_94 (O_94,N_2961,N_2936);
nand UO_95 (O_95,N_2946,N_2933);
and UO_96 (O_96,N_2941,N_2913);
nand UO_97 (O_97,N_2996,N_2900);
or UO_98 (O_98,N_2902,N_2980);
nand UO_99 (O_99,N_2979,N_2971);
or UO_100 (O_100,N_2985,N_2913);
and UO_101 (O_101,N_2906,N_2991);
nor UO_102 (O_102,N_2971,N_2989);
or UO_103 (O_103,N_2966,N_2969);
and UO_104 (O_104,N_2976,N_2993);
nor UO_105 (O_105,N_2969,N_2917);
or UO_106 (O_106,N_2993,N_2949);
nand UO_107 (O_107,N_2941,N_2906);
nand UO_108 (O_108,N_2997,N_2924);
and UO_109 (O_109,N_2937,N_2989);
and UO_110 (O_110,N_2975,N_2982);
nand UO_111 (O_111,N_2913,N_2907);
nand UO_112 (O_112,N_2966,N_2936);
xnor UO_113 (O_113,N_2960,N_2901);
and UO_114 (O_114,N_2934,N_2916);
or UO_115 (O_115,N_2986,N_2965);
or UO_116 (O_116,N_2958,N_2968);
xnor UO_117 (O_117,N_2941,N_2954);
nor UO_118 (O_118,N_2965,N_2988);
nor UO_119 (O_119,N_2956,N_2909);
xnor UO_120 (O_120,N_2974,N_2962);
nor UO_121 (O_121,N_2969,N_2907);
or UO_122 (O_122,N_2913,N_2945);
nor UO_123 (O_123,N_2990,N_2972);
nor UO_124 (O_124,N_2944,N_2982);
nand UO_125 (O_125,N_2956,N_2999);
and UO_126 (O_126,N_2906,N_2926);
or UO_127 (O_127,N_2979,N_2937);
xnor UO_128 (O_128,N_2991,N_2949);
nor UO_129 (O_129,N_2920,N_2995);
and UO_130 (O_130,N_2973,N_2918);
nand UO_131 (O_131,N_2908,N_2966);
nand UO_132 (O_132,N_2977,N_2960);
nand UO_133 (O_133,N_2951,N_2975);
and UO_134 (O_134,N_2960,N_2900);
nor UO_135 (O_135,N_2992,N_2977);
xor UO_136 (O_136,N_2972,N_2969);
xor UO_137 (O_137,N_2937,N_2970);
or UO_138 (O_138,N_2931,N_2976);
and UO_139 (O_139,N_2941,N_2979);
or UO_140 (O_140,N_2995,N_2975);
nor UO_141 (O_141,N_2944,N_2995);
nor UO_142 (O_142,N_2995,N_2947);
nor UO_143 (O_143,N_2913,N_2928);
nor UO_144 (O_144,N_2906,N_2902);
nand UO_145 (O_145,N_2916,N_2962);
xnor UO_146 (O_146,N_2963,N_2971);
nand UO_147 (O_147,N_2970,N_2979);
nor UO_148 (O_148,N_2965,N_2992);
nand UO_149 (O_149,N_2980,N_2960);
nor UO_150 (O_150,N_2945,N_2909);
and UO_151 (O_151,N_2992,N_2907);
xor UO_152 (O_152,N_2957,N_2922);
nor UO_153 (O_153,N_2997,N_2909);
xor UO_154 (O_154,N_2955,N_2918);
or UO_155 (O_155,N_2992,N_2949);
and UO_156 (O_156,N_2971,N_2942);
xor UO_157 (O_157,N_2922,N_2919);
or UO_158 (O_158,N_2905,N_2907);
nor UO_159 (O_159,N_2915,N_2968);
nor UO_160 (O_160,N_2904,N_2907);
or UO_161 (O_161,N_2919,N_2965);
xor UO_162 (O_162,N_2974,N_2920);
nand UO_163 (O_163,N_2983,N_2962);
or UO_164 (O_164,N_2972,N_2922);
nand UO_165 (O_165,N_2913,N_2948);
or UO_166 (O_166,N_2905,N_2902);
and UO_167 (O_167,N_2922,N_2949);
or UO_168 (O_168,N_2985,N_2939);
nor UO_169 (O_169,N_2925,N_2948);
nand UO_170 (O_170,N_2985,N_2921);
nand UO_171 (O_171,N_2992,N_2917);
nor UO_172 (O_172,N_2959,N_2983);
and UO_173 (O_173,N_2944,N_2911);
or UO_174 (O_174,N_2903,N_2958);
or UO_175 (O_175,N_2922,N_2939);
nor UO_176 (O_176,N_2995,N_2909);
and UO_177 (O_177,N_2932,N_2964);
xnor UO_178 (O_178,N_2924,N_2939);
or UO_179 (O_179,N_2950,N_2955);
or UO_180 (O_180,N_2936,N_2916);
nor UO_181 (O_181,N_2943,N_2914);
and UO_182 (O_182,N_2914,N_2959);
nand UO_183 (O_183,N_2998,N_2942);
nand UO_184 (O_184,N_2959,N_2951);
nand UO_185 (O_185,N_2983,N_2938);
nor UO_186 (O_186,N_2909,N_2977);
or UO_187 (O_187,N_2991,N_2909);
xnor UO_188 (O_188,N_2991,N_2969);
nor UO_189 (O_189,N_2969,N_2990);
and UO_190 (O_190,N_2938,N_2973);
nor UO_191 (O_191,N_2905,N_2950);
or UO_192 (O_192,N_2902,N_2944);
nand UO_193 (O_193,N_2923,N_2961);
nand UO_194 (O_194,N_2950,N_2966);
and UO_195 (O_195,N_2974,N_2980);
xor UO_196 (O_196,N_2939,N_2943);
nor UO_197 (O_197,N_2982,N_2909);
nor UO_198 (O_198,N_2988,N_2933);
nor UO_199 (O_199,N_2988,N_2902);
nand UO_200 (O_200,N_2907,N_2902);
and UO_201 (O_201,N_2901,N_2912);
xor UO_202 (O_202,N_2920,N_2949);
nand UO_203 (O_203,N_2974,N_2919);
nor UO_204 (O_204,N_2948,N_2954);
or UO_205 (O_205,N_2973,N_2974);
or UO_206 (O_206,N_2954,N_2930);
xor UO_207 (O_207,N_2987,N_2970);
and UO_208 (O_208,N_2968,N_2923);
and UO_209 (O_209,N_2934,N_2932);
or UO_210 (O_210,N_2912,N_2905);
nand UO_211 (O_211,N_2935,N_2976);
and UO_212 (O_212,N_2920,N_2952);
or UO_213 (O_213,N_2915,N_2935);
nor UO_214 (O_214,N_2942,N_2946);
xor UO_215 (O_215,N_2948,N_2975);
xor UO_216 (O_216,N_2954,N_2916);
nand UO_217 (O_217,N_2904,N_2945);
or UO_218 (O_218,N_2904,N_2934);
xor UO_219 (O_219,N_2986,N_2923);
nor UO_220 (O_220,N_2968,N_2975);
nand UO_221 (O_221,N_2907,N_2974);
or UO_222 (O_222,N_2932,N_2986);
xor UO_223 (O_223,N_2976,N_2907);
nand UO_224 (O_224,N_2902,N_2972);
nand UO_225 (O_225,N_2928,N_2919);
and UO_226 (O_226,N_2943,N_2994);
and UO_227 (O_227,N_2924,N_2971);
nor UO_228 (O_228,N_2991,N_2959);
nor UO_229 (O_229,N_2987,N_2989);
nor UO_230 (O_230,N_2997,N_2953);
and UO_231 (O_231,N_2961,N_2980);
nand UO_232 (O_232,N_2930,N_2909);
nor UO_233 (O_233,N_2917,N_2981);
and UO_234 (O_234,N_2914,N_2991);
and UO_235 (O_235,N_2925,N_2991);
nor UO_236 (O_236,N_2955,N_2938);
nand UO_237 (O_237,N_2935,N_2991);
or UO_238 (O_238,N_2912,N_2963);
and UO_239 (O_239,N_2960,N_2916);
nand UO_240 (O_240,N_2962,N_2999);
or UO_241 (O_241,N_2982,N_2925);
and UO_242 (O_242,N_2950,N_2987);
or UO_243 (O_243,N_2954,N_2909);
and UO_244 (O_244,N_2973,N_2998);
nand UO_245 (O_245,N_2999,N_2938);
nand UO_246 (O_246,N_2981,N_2979);
and UO_247 (O_247,N_2971,N_2998);
or UO_248 (O_248,N_2976,N_2919);
nor UO_249 (O_249,N_2943,N_2956);
nand UO_250 (O_250,N_2923,N_2916);
nor UO_251 (O_251,N_2909,N_2934);
or UO_252 (O_252,N_2938,N_2948);
xnor UO_253 (O_253,N_2941,N_2903);
nand UO_254 (O_254,N_2966,N_2953);
nand UO_255 (O_255,N_2963,N_2952);
and UO_256 (O_256,N_2979,N_2984);
nand UO_257 (O_257,N_2923,N_2921);
nand UO_258 (O_258,N_2983,N_2914);
nor UO_259 (O_259,N_2929,N_2933);
and UO_260 (O_260,N_2900,N_2998);
nand UO_261 (O_261,N_2939,N_2946);
or UO_262 (O_262,N_2906,N_2907);
xor UO_263 (O_263,N_2971,N_2929);
or UO_264 (O_264,N_2922,N_2992);
xnor UO_265 (O_265,N_2908,N_2948);
nor UO_266 (O_266,N_2993,N_2967);
nor UO_267 (O_267,N_2936,N_2979);
or UO_268 (O_268,N_2997,N_2928);
nand UO_269 (O_269,N_2989,N_2911);
nand UO_270 (O_270,N_2953,N_2944);
xor UO_271 (O_271,N_2965,N_2995);
xnor UO_272 (O_272,N_2954,N_2980);
xor UO_273 (O_273,N_2918,N_2940);
nand UO_274 (O_274,N_2967,N_2955);
nand UO_275 (O_275,N_2909,N_2989);
nor UO_276 (O_276,N_2935,N_2949);
nand UO_277 (O_277,N_2945,N_2992);
or UO_278 (O_278,N_2998,N_2984);
nand UO_279 (O_279,N_2998,N_2916);
and UO_280 (O_280,N_2986,N_2989);
nor UO_281 (O_281,N_2913,N_2990);
or UO_282 (O_282,N_2966,N_2909);
nor UO_283 (O_283,N_2920,N_2987);
and UO_284 (O_284,N_2925,N_2906);
and UO_285 (O_285,N_2995,N_2967);
or UO_286 (O_286,N_2921,N_2936);
and UO_287 (O_287,N_2904,N_2949);
or UO_288 (O_288,N_2975,N_2981);
nor UO_289 (O_289,N_2938,N_2966);
and UO_290 (O_290,N_2907,N_2955);
nand UO_291 (O_291,N_2930,N_2928);
and UO_292 (O_292,N_2916,N_2976);
and UO_293 (O_293,N_2948,N_2984);
and UO_294 (O_294,N_2921,N_2994);
nor UO_295 (O_295,N_2987,N_2932);
nand UO_296 (O_296,N_2969,N_2971);
or UO_297 (O_297,N_2952,N_2992);
or UO_298 (O_298,N_2950,N_2975);
xnor UO_299 (O_299,N_2900,N_2920);
or UO_300 (O_300,N_2924,N_2916);
nand UO_301 (O_301,N_2955,N_2994);
and UO_302 (O_302,N_2974,N_2925);
nor UO_303 (O_303,N_2964,N_2958);
nand UO_304 (O_304,N_2956,N_2930);
xnor UO_305 (O_305,N_2905,N_2932);
nor UO_306 (O_306,N_2970,N_2927);
nor UO_307 (O_307,N_2907,N_2953);
xnor UO_308 (O_308,N_2971,N_2927);
nor UO_309 (O_309,N_2980,N_2953);
and UO_310 (O_310,N_2964,N_2934);
and UO_311 (O_311,N_2900,N_2953);
and UO_312 (O_312,N_2932,N_2996);
nor UO_313 (O_313,N_2941,N_2930);
nor UO_314 (O_314,N_2909,N_2981);
nand UO_315 (O_315,N_2919,N_2997);
nand UO_316 (O_316,N_2974,N_2926);
nor UO_317 (O_317,N_2907,N_2984);
nor UO_318 (O_318,N_2909,N_2908);
nor UO_319 (O_319,N_2926,N_2978);
or UO_320 (O_320,N_2921,N_2916);
xor UO_321 (O_321,N_2915,N_2943);
nor UO_322 (O_322,N_2990,N_2934);
or UO_323 (O_323,N_2975,N_2900);
and UO_324 (O_324,N_2904,N_2941);
nand UO_325 (O_325,N_2933,N_2973);
nor UO_326 (O_326,N_2981,N_2982);
nand UO_327 (O_327,N_2942,N_2956);
and UO_328 (O_328,N_2952,N_2909);
xor UO_329 (O_329,N_2955,N_2913);
and UO_330 (O_330,N_2988,N_2985);
nand UO_331 (O_331,N_2919,N_2907);
xnor UO_332 (O_332,N_2932,N_2940);
and UO_333 (O_333,N_2909,N_2992);
nor UO_334 (O_334,N_2921,N_2984);
xnor UO_335 (O_335,N_2970,N_2944);
or UO_336 (O_336,N_2956,N_2954);
and UO_337 (O_337,N_2914,N_2950);
nand UO_338 (O_338,N_2925,N_2976);
nand UO_339 (O_339,N_2958,N_2953);
and UO_340 (O_340,N_2924,N_2912);
nand UO_341 (O_341,N_2971,N_2977);
nand UO_342 (O_342,N_2936,N_2919);
xnor UO_343 (O_343,N_2919,N_2999);
or UO_344 (O_344,N_2962,N_2975);
nand UO_345 (O_345,N_2936,N_2906);
nor UO_346 (O_346,N_2919,N_2960);
and UO_347 (O_347,N_2946,N_2969);
or UO_348 (O_348,N_2906,N_2973);
xnor UO_349 (O_349,N_2900,N_2917);
nor UO_350 (O_350,N_2989,N_2992);
nand UO_351 (O_351,N_2926,N_2900);
and UO_352 (O_352,N_2975,N_2984);
and UO_353 (O_353,N_2902,N_2946);
and UO_354 (O_354,N_2985,N_2953);
and UO_355 (O_355,N_2955,N_2966);
and UO_356 (O_356,N_2938,N_2925);
or UO_357 (O_357,N_2943,N_2920);
or UO_358 (O_358,N_2988,N_2912);
nor UO_359 (O_359,N_2963,N_2987);
and UO_360 (O_360,N_2955,N_2965);
or UO_361 (O_361,N_2962,N_2935);
or UO_362 (O_362,N_2959,N_2979);
and UO_363 (O_363,N_2952,N_2987);
nand UO_364 (O_364,N_2994,N_2906);
xor UO_365 (O_365,N_2983,N_2924);
nor UO_366 (O_366,N_2917,N_2956);
nand UO_367 (O_367,N_2911,N_2987);
xor UO_368 (O_368,N_2930,N_2900);
and UO_369 (O_369,N_2925,N_2935);
or UO_370 (O_370,N_2961,N_2926);
nand UO_371 (O_371,N_2937,N_2976);
xor UO_372 (O_372,N_2936,N_2948);
nand UO_373 (O_373,N_2920,N_2951);
or UO_374 (O_374,N_2924,N_2902);
nand UO_375 (O_375,N_2948,N_2941);
nand UO_376 (O_376,N_2966,N_2903);
nand UO_377 (O_377,N_2963,N_2906);
xor UO_378 (O_378,N_2948,N_2919);
and UO_379 (O_379,N_2986,N_2938);
nor UO_380 (O_380,N_2982,N_2933);
and UO_381 (O_381,N_2929,N_2961);
and UO_382 (O_382,N_2913,N_2919);
or UO_383 (O_383,N_2901,N_2905);
nor UO_384 (O_384,N_2996,N_2919);
or UO_385 (O_385,N_2994,N_2989);
and UO_386 (O_386,N_2907,N_2918);
nor UO_387 (O_387,N_2901,N_2926);
or UO_388 (O_388,N_2931,N_2988);
and UO_389 (O_389,N_2937,N_2958);
nor UO_390 (O_390,N_2918,N_2958);
and UO_391 (O_391,N_2973,N_2930);
xor UO_392 (O_392,N_2927,N_2922);
nand UO_393 (O_393,N_2915,N_2947);
and UO_394 (O_394,N_2920,N_2912);
and UO_395 (O_395,N_2952,N_2993);
nand UO_396 (O_396,N_2953,N_2973);
nand UO_397 (O_397,N_2922,N_2986);
nor UO_398 (O_398,N_2961,N_2940);
nand UO_399 (O_399,N_2988,N_2951);
and UO_400 (O_400,N_2949,N_2972);
nand UO_401 (O_401,N_2933,N_2917);
nand UO_402 (O_402,N_2989,N_2963);
nand UO_403 (O_403,N_2932,N_2979);
and UO_404 (O_404,N_2983,N_2953);
nand UO_405 (O_405,N_2972,N_2941);
and UO_406 (O_406,N_2935,N_2977);
nand UO_407 (O_407,N_2964,N_2923);
nand UO_408 (O_408,N_2995,N_2953);
and UO_409 (O_409,N_2969,N_2978);
nand UO_410 (O_410,N_2901,N_2951);
or UO_411 (O_411,N_2949,N_2942);
and UO_412 (O_412,N_2942,N_2933);
nand UO_413 (O_413,N_2954,N_2914);
nand UO_414 (O_414,N_2929,N_2921);
nand UO_415 (O_415,N_2952,N_2927);
nand UO_416 (O_416,N_2922,N_2917);
nor UO_417 (O_417,N_2910,N_2913);
nand UO_418 (O_418,N_2923,N_2903);
nor UO_419 (O_419,N_2976,N_2982);
and UO_420 (O_420,N_2977,N_2957);
nand UO_421 (O_421,N_2953,N_2926);
nand UO_422 (O_422,N_2998,N_2980);
xor UO_423 (O_423,N_2983,N_2903);
or UO_424 (O_424,N_2943,N_2940);
or UO_425 (O_425,N_2905,N_2988);
or UO_426 (O_426,N_2910,N_2933);
nand UO_427 (O_427,N_2921,N_2950);
or UO_428 (O_428,N_2990,N_2915);
and UO_429 (O_429,N_2953,N_2933);
nor UO_430 (O_430,N_2945,N_2920);
nand UO_431 (O_431,N_2936,N_2960);
or UO_432 (O_432,N_2963,N_2946);
xnor UO_433 (O_433,N_2985,N_2925);
nor UO_434 (O_434,N_2937,N_2964);
or UO_435 (O_435,N_2943,N_2987);
and UO_436 (O_436,N_2985,N_2986);
and UO_437 (O_437,N_2945,N_2926);
nor UO_438 (O_438,N_2988,N_2927);
nand UO_439 (O_439,N_2952,N_2938);
xnor UO_440 (O_440,N_2935,N_2904);
nor UO_441 (O_441,N_2914,N_2909);
or UO_442 (O_442,N_2982,N_2905);
nor UO_443 (O_443,N_2974,N_2923);
or UO_444 (O_444,N_2900,N_2958);
nor UO_445 (O_445,N_2944,N_2963);
and UO_446 (O_446,N_2986,N_2921);
nand UO_447 (O_447,N_2900,N_2903);
nand UO_448 (O_448,N_2909,N_2979);
nor UO_449 (O_449,N_2940,N_2992);
or UO_450 (O_450,N_2991,N_2990);
and UO_451 (O_451,N_2980,N_2917);
nor UO_452 (O_452,N_2913,N_2906);
and UO_453 (O_453,N_2995,N_2984);
and UO_454 (O_454,N_2954,N_2952);
xor UO_455 (O_455,N_2960,N_2983);
nor UO_456 (O_456,N_2995,N_2966);
nor UO_457 (O_457,N_2964,N_2900);
and UO_458 (O_458,N_2961,N_2901);
or UO_459 (O_459,N_2997,N_2905);
or UO_460 (O_460,N_2998,N_2903);
and UO_461 (O_461,N_2995,N_2935);
and UO_462 (O_462,N_2956,N_2985);
nand UO_463 (O_463,N_2934,N_2991);
nor UO_464 (O_464,N_2983,N_2923);
or UO_465 (O_465,N_2926,N_2992);
and UO_466 (O_466,N_2906,N_2912);
nand UO_467 (O_467,N_2998,N_2902);
nor UO_468 (O_468,N_2941,N_2990);
or UO_469 (O_469,N_2924,N_2920);
and UO_470 (O_470,N_2949,N_2957);
and UO_471 (O_471,N_2951,N_2906);
and UO_472 (O_472,N_2929,N_2982);
nor UO_473 (O_473,N_2964,N_2903);
nand UO_474 (O_474,N_2987,N_2966);
xor UO_475 (O_475,N_2936,N_2969);
or UO_476 (O_476,N_2935,N_2901);
xnor UO_477 (O_477,N_2931,N_2939);
and UO_478 (O_478,N_2943,N_2938);
nor UO_479 (O_479,N_2931,N_2904);
xnor UO_480 (O_480,N_2910,N_2980);
nor UO_481 (O_481,N_2973,N_2920);
and UO_482 (O_482,N_2960,N_2968);
and UO_483 (O_483,N_2915,N_2977);
nand UO_484 (O_484,N_2948,N_2934);
nor UO_485 (O_485,N_2964,N_2916);
xnor UO_486 (O_486,N_2934,N_2910);
and UO_487 (O_487,N_2967,N_2987);
or UO_488 (O_488,N_2930,N_2915);
xnor UO_489 (O_489,N_2937,N_2922);
or UO_490 (O_490,N_2958,N_2929);
and UO_491 (O_491,N_2937,N_2954);
nand UO_492 (O_492,N_2982,N_2962);
nor UO_493 (O_493,N_2965,N_2917);
xor UO_494 (O_494,N_2955,N_2935);
nand UO_495 (O_495,N_2933,N_2995);
nor UO_496 (O_496,N_2901,N_2915);
nand UO_497 (O_497,N_2924,N_2937);
nand UO_498 (O_498,N_2905,N_2931);
nand UO_499 (O_499,N_2953,N_2952);
endmodule