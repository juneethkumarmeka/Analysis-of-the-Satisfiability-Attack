module basic_750_5000_1000_2_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2507,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2522,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2533,N_2534,N_2536,N_2537,N_2538,N_2539,N_2542,N_2543,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2554,N_2557,N_2558,N_2559,N_2560,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2611,N_2612,N_2613,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2623,N_2624,N_2625,N_2627,N_2628,N_2629,N_2630,N_2631,N_2633,N_2636,N_2637,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2648,N_2649,N_2650,N_2651,N_2653,N_2656,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2672,N_2674,N_2675,N_2676,N_2677,N_2678,N_2682,N_2683,N_2684,N_2687,N_2688,N_2690,N_2691,N_2693,N_2694,N_2696,N_2697,N_2698,N_2699,N_2700,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2760,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2804,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2824,N_2826,N_2827,N_2829,N_2830,N_2833,N_2834,N_2836,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2845,N_2846,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2857,N_2859,N_2860,N_2861,N_2862,N_2864,N_2866,N_2867,N_2869,N_2870,N_2871,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2891,N_2892,N_2893,N_2894,N_2896,N_2898,N_2900,N_2901,N_2903,N_2904,N_2905,N_2907,N_2908,N_2909,N_2911,N_2912,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2923,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2948,N_2949,N_2952,N_2953,N_2954,N_2956,N_2957,N_2958,N_2959,N_2962,N_2964,N_2965,N_2966,N_2967,N_2969,N_2970,N_2971,N_2976,N_2978,N_2979,N_2981,N_2983,N_2984,N_2985,N_2986,N_2987,N_2990,N_2991,N_2992,N_2994,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3018,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3038,N_3040,N_3041,N_3042,N_3043,N_3044,N_3046,N_3048,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3060,N_3061,N_3062,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3090,N_3091,N_3092,N_3093,N_3095,N_3096,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3170,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3196,N_3197,N_3199,N_3200,N_3201,N_3202,N_3203,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3214,N_3216,N_3217,N_3218,N_3219,N_3220,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3229,N_3230,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3239,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3260,N_3261,N_3263,N_3265,N_3266,N_3267,N_3269,N_3270,N_3272,N_3273,N_3274,N_3275,N_3277,N_3279,N_3281,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3301,N_3302,N_3303,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3319,N_3320,N_3321,N_3325,N_3327,N_3328,N_3329,N_3332,N_3333,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3343,N_3344,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3376,N_3377,N_3378,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3426,N_3427,N_3428,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3440,N_3441,N_3442,N_3444,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3453,N_3454,N_3455,N_3458,N_3459,N_3461,N_3462,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3487,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3498,N_3499,N_3500,N_3503,N_3504,N_3507,N_3511,N_3512,N_3514,N_3515,N_3516,N_3518,N_3519,N_3520,N_3521,N_3522,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3536,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3558,N_3559,N_3560,N_3561,N_3564,N_3566,N_3567,N_3568,N_3569,N_3571,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3582,N_3583,N_3584,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3604,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3613,N_3614,N_3616,N_3617,N_3618,N_3619,N_3620,N_3622,N_3623,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3632,N_3633,N_3636,N_3637,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3649,N_3650,N_3651,N_3653,N_3654,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3720,N_3722,N_3723,N_3726,N_3727,N_3728,N_3731,N_3732,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3777,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3803,N_3804,N_3805,N_3808,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3835,N_3836,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3869,N_3870,N_3871,N_3872,N_3874,N_3875,N_3877,N_3878,N_3879,N_3882,N_3883,N_3884,N_3885,N_3886,N_3888,N_3889,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3916,N_3917,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4010,N_4011,N_4014,N_4015,N_4017,N_4018,N_4019,N_4020,N_4021,N_4024,N_4026,N_4027,N_4028,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4055,N_4056,N_4058,N_4059,N_4060,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4076,N_4078,N_4079,N_4081,N_4082,N_4084,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4097,N_4098,N_4099,N_4100,N_4102,N_4104,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4121,N_4122,N_4124,N_4126,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4186,N_4187,N_4188,N_4190,N_4192,N_4193,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4220,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4241,N_4242,N_4243,N_4244,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4257,N_4259,N_4260,N_4261,N_4262,N_4266,N_4268,N_4269,N_4270,N_4272,N_4274,N_4275,N_4276,N_4277,N_4278,N_4281,N_4282,N_4283,N_4284,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4300,N_4301,N_4302,N_4304,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4326,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4335,N_4336,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4349,N_4351,N_4352,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4394,N_4395,N_4396,N_4397,N_4399,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4422,N_4423,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4438,N_4439,N_4440,N_4441,N_4443,N_4446,N_4447,N_4448,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4459,N_4460,N_4461,N_4463,N_4464,N_4465,N_4467,N_4468,N_4469,N_4470,N_4471,N_4473,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4496,N_4497,N_4500,N_4501,N_4502,N_4503,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4524,N_4526,N_4527,N_4528,N_4529,N_4530,N_4532,N_4533,N_4536,N_4537,N_4538,N_4541,N_4544,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4559,N_4560,N_4561,N_4562,N_4564,N_4565,N_4566,N_4567,N_4569,N_4570,N_4571,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4604,N_4605,N_4607,N_4608,N_4609,N_4610,N_4611,N_4614,N_4616,N_4617,N_4618,N_4620,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4632,N_4633,N_4634,N_4635,N_4636,N_4638,N_4639,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4649,N_4650,N_4652,N_4653,N_4654,N_4656,N_4657,N_4658,N_4659,N_4662,N_4663,N_4664,N_4665,N_4667,N_4668,N_4669,N_4672,N_4673,N_4676,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4699,N_4700,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4711,N_4715,N_4716,N_4717,N_4718,N_4719,N_4721,N_4722,N_4723,N_4724,N_4725,N_4727,N_4728,N_4729,N_4730,N_4731,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4754,N_4756,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4790,N_4792,N_4794,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4803,N_4805,N_4806,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4820,N_4821,N_4822,N_4823,N_4824,N_4826,N_4827,N_4829,N_4830,N_4831,N_4832,N_4836,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4856,N_4857,N_4858,N_4859,N_4860,N_4862,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4903,N_4904,N_4906,N_4908,N_4909,N_4910,N_4912,N_4913,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4924,N_4927,N_4928,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4945,N_4946,N_4948,N_4951,N_4953,N_4954,N_4956,N_4957,N_4958,N_4959,N_4960,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4979,N_4980,N_4981,N_4982,N_4985,N_4986,N_4987,N_4989,N_4990,N_4994,N_4995,N_4997,N_4998,N_4999;
nand U0 (N_0,In_267,In_409);
or U1 (N_1,In_611,In_631);
nand U2 (N_2,In_721,In_155);
nand U3 (N_3,In_254,In_501);
nor U4 (N_4,In_420,In_26);
or U5 (N_5,In_452,In_690);
nor U6 (N_6,In_192,In_327);
and U7 (N_7,In_536,In_310);
or U8 (N_8,In_285,In_625);
nor U9 (N_9,In_657,In_693);
nand U10 (N_10,In_340,In_649);
or U11 (N_11,In_707,In_390);
nor U12 (N_12,In_164,In_726);
nor U13 (N_13,In_470,In_547);
xor U14 (N_14,In_110,In_601);
nand U15 (N_15,In_0,In_580);
nand U16 (N_16,In_562,In_518);
and U17 (N_17,In_100,In_575);
and U18 (N_18,In_407,In_274);
or U19 (N_19,In_668,In_578);
and U20 (N_20,In_179,In_524);
nor U21 (N_21,In_720,In_665);
nand U22 (N_22,In_515,In_188);
or U23 (N_23,In_587,In_465);
nand U24 (N_24,In_156,In_508);
nand U25 (N_25,In_541,In_493);
nand U26 (N_26,In_667,In_102);
or U27 (N_27,In_451,In_216);
nor U28 (N_28,In_231,In_417);
nand U29 (N_29,In_727,In_299);
nand U30 (N_30,In_238,In_106);
nand U31 (N_31,In_256,In_675);
or U32 (N_32,In_653,In_467);
or U33 (N_33,In_641,In_77);
nor U34 (N_34,In_126,In_91);
and U35 (N_35,In_645,In_161);
or U36 (N_36,In_84,In_162);
or U37 (N_37,In_209,In_702);
or U38 (N_38,In_85,In_712);
or U39 (N_39,In_558,In_554);
and U40 (N_40,In_512,In_260);
or U41 (N_41,In_525,In_64);
or U42 (N_42,In_731,In_313);
xnor U43 (N_43,In_134,In_535);
or U44 (N_44,In_208,In_447);
or U45 (N_45,In_430,In_309);
nand U46 (N_46,In_288,In_70);
nor U47 (N_47,In_78,In_176);
nand U48 (N_48,In_98,In_442);
nand U49 (N_49,In_159,In_714);
nand U50 (N_50,In_343,In_549);
or U51 (N_51,In_568,In_503);
nand U52 (N_52,In_529,In_416);
or U53 (N_53,In_421,In_160);
nand U54 (N_54,In_369,In_199);
nor U55 (N_55,In_686,In_632);
nand U56 (N_56,In_249,In_300);
nor U57 (N_57,In_31,In_744);
and U58 (N_58,In_295,In_151);
and U59 (N_59,In_647,In_579);
nand U60 (N_60,In_545,In_698);
and U61 (N_61,In_172,In_105);
or U62 (N_62,In_688,In_328);
or U63 (N_63,In_373,In_356);
nor U64 (N_64,In_207,In_144);
and U65 (N_65,In_509,In_487);
nand U66 (N_66,In_415,In_259);
and U67 (N_67,In_537,In_92);
nor U68 (N_68,In_703,In_358);
nand U69 (N_69,In_643,In_431);
nor U70 (N_70,In_555,In_594);
nand U71 (N_71,In_227,In_150);
nor U72 (N_72,In_292,In_426);
xor U73 (N_73,In_165,In_119);
nor U74 (N_74,In_52,In_224);
nor U75 (N_75,In_93,In_315);
nor U76 (N_76,In_252,In_414);
or U77 (N_77,In_670,In_510);
nand U78 (N_78,In_71,In_200);
nand U79 (N_79,In_748,In_527);
nand U80 (N_80,In_571,In_459);
and U81 (N_81,In_174,In_616);
nand U82 (N_82,In_683,In_305);
nor U83 (N_83,In_226,In_335);
nor U84 (N_84,In_312,In_364);
nand U85 (N_85,In_29,In_76);
nand U86 (N_86,In_242,In_419);
and U87 (N_87,In_410,In_404);
nor U88 (N_88,In_41,In_546);
or U89 (N_89,In_652,In_177);
or U90 (N_90,In_507,In_63);
and U91 (N_91,In_214,In_290);
and U92 (N_92,In_21,In_379);
nand U93 (N_93,In_435,In_651);
or U94 (N_94,In_87,In_674);
nor U95 (N_95,In_719,In_143);
xnor U96 (N_96,In_514,In_573);
nand U97 (N_97,In_112,In_730);
nand U98 (N_98,In_736,In_169);
and U99 (N_99,In_363,In_293);
or U100 (N_100,In_307,In_598);
nor U101 (N_101,In_424,In_3);
and U102 (N_102,In_183,In_5);
and U103 (N_103,In_220,In_8);
nor U104 (N_104,In_572,In_83);
xor U105 (N_105,In_139,In_681);
xor U106 (N_106,In_23,In_137);
nand U107 (N_107,In_449,In_294);
and U108 (N_108,In_552,In_215);
and U109 (N_109,In_271,In_34);
and U110 (N_110,In_483,In_347);
nor U111 (N_111,In_154,In_479);
nand U112 (N_112,In_103,In_287);
nor U113 (N_113,In_197,In_732);
nor U114 (N_114,In_19,In_418);
nor U115 (N_115,In_478,In_619);
nand U116 (N_116,In_633,In_40);
and U117 (N_117,In_43,In_659);
nand U118 (N_118,In_733,In_704);
or U119 (N_119,In_116,In_436);
nand U120 (N_120,In_261,In_11);
or U121 (N_121,In_339,In_73);
nor U122 (N_122,In_49,In_157);
nand U123 (N_123,In_303,In_376);
nor U124 (N_124,In_301,In_740);
and U125 (N_125,In_357,In_79);
nor U126 (N_126,In_277,In_684);
nand U127 (N_127,In_669,In_565);
and U128 (N_128,In_69,In_253);
and U129 (N_129,In_716,In_354);
nand U130 (N_130,In_745,In_486);
or U131 (N_131,In_530,In_602);
nand U132 (N_132,In_236,In_316);
or U133 (N_133,In_570,In_735);
nor U134 (N_134,In_403,In_248);
or U135 (N_135,In_320,In_621);
nor U136 (N_136,In_60,In_246);
nand U137 (N_137,In_664,In_297);
and U138 (N_138,In_685,In_86);
or U139 (N_139,In_251,In_663);
nor U140 (N_140,In_279,In_24);
nand U141 (N_141,In_269,In_14);
or U142 (N_142,In_221,In_196);
and U143 (N_143,In_47,In_377);
xor U144 (N_144,In_202,In_463);
and U145 (N_145,In_175,In_229);
nand U146 (N_146,In_146,In_485);
nand U147 (N_147,In_427,In_694);
or U148 (N_148,In_710,In_550);
nor U149 (N_149,In_689,In_206);
nand U150 (N_150,In_495,In_350);
or U151 (N_151,In_286,In_506);
or U152 (N_152,In_630,In_408);
nand U153 (N_153,In_173,In_38);
and U154 (N_154,In_96,In_241);
nand U155 (N_155,In_386,In_687);
nand U156 (N_156,In_16,In_44);
nand U157 (N_157,In_20,In_266);
or U158 (N_158,In_351,In_245);
nor U159 (N_159,In_324,In_608);
and U160 (N_160,In_729,In_140);
nand U161 (N_161,In_658,In_39);
nand U162 (N_162,In_32,In_640);
nand U163 (N_163,In_272,In_444);
nand U164 (N_164,In_682,In_511);
nor U165 (N_165,In_713,In_603);
nor U166 (N_166,In_171,In_74);
nor U167 (N_167,In_233,In_184);
and U168 (N_168,In_66,In_636);
or U169 (N_169,In_393,In_380);
nor U170 (N_170,In_481,In_33);
nand U171 (N_171,In_326,In_135);
or U172 (N_172,In_428,In_461);
and U173 (N_173,In_378,In_265);
nor U174 (N_174,In_677,In_523);
nand U175 (N_175,In_268,In_255);
or U176 (N_176,In_217,In_434);
and U177 (N_177,In_388,In_212);
and U178 (N_178,In_498,In_634);
nor U179 (N_179,In_62,In_322);
nor U180 (N_180,In_345,In_708);
nand U181 (N_181,In_333,In_395);
xnor U182 (N_182,In_574,In_648);
and U183 (N_183,In_563,In_392);
xnor U184 (N_184,In_27,In_232);
or U185 (N_185,In_57,In_371);
nor U186 (N_186,In_168,In_747);
or U187 (N_187,In_400,In_230);
nor U188 (N_188,In_638,In_348);
nor U189 (N_189,In_482,In_423);
nor U190 (N_190,In_225,In_374);
nand U191 (N_191,In_411,In_4);
nor U192 (N_192,In_491,In_656);
and U193 (N_193,In_557,In_114);
or U194 (N_194,In_142,In_567);
or U195 (N_195,In_104,In_678);
nand U196 (N_196,In_178,In_422);
nor U197 (N_197,In_737,In_589);
nand U198 (N_198,In_739,In_50);
nand U199 (N_199,In_129,In_367);
nand U200 (N_200,In_127,In_560);
nor U201 (N_201,In_355,In_130);
nor U202 (N_202,In_239,In_584);
nor U203 (N_203,In_718,In_115);
nor U204 (N_204,In_15,In_58);
and U205 (N_205,In_605,In_457);
nor U206 (N_206,In_321,In_402);
nor U207 (N_207,In_592,In_551);
or U208 (N_208,In_472,In_650);
nor U209 (N_209,In_504,In_456);
or U210 (N_210,In_332,In_443);
or U211 (N_211,In_28,In_383);
xnor U212 (N_212,In_654,In_113);
and U213 (N_213,In_158,In_672);
and U214 (N_214,In_706,In_588);
or U215 (N_215,In_488,In_476);
or U216 (N_216,In_696,In_9);
or U217 (N_217,In_186,In_42);
nand U218 (N_218,In_412,In_240);
or U219 (N_219,In_724,In_539);
nor U220 (N_220,In_189,In_662);
or U221 (N_221,In_505,In_749);
and U222 (N_222,In_95,In_145);
nor U223 (N_223,In_89,In_325);
nor U224 (N_224,In_723,In_468);
nor U225 (N_225,In_247,In_540);
and U226 (N_226,In_553,In_695);
nand U227 (N_227,In_180,In_626);
nor U228 (N_228,In_118,In_170);
or U229 (N_229,In_368,In_341);
or U230 (N_230,In_25,In_500);
nand U231 (N_231,In_474,In_282);
and U232 (N_232,In_97,In_607);
or U233 (N_233,In_715,In_593);
or U234 (N_234,In_661,In_396);
or U235 (N_235,In_673,In_10);
nand U236 (N_236,In_17,In_148);
or U237 (N_237,In_627,In_599);
xor U238 (N_238,In_741,In_477);
nand U239 (N_239,In_205,In_384);
nand U240 (N_240,In_319,In_360);
or U241 (N_241,In_273,In_490);
nand U242 (N_242,In_136,In_211);
nor U243 (N_243,In_53,In_697);
nor U244 (N_244,In_306,In_51);
nor U245 (N_245,In_466,In_37);
nor U246 (N_246,In_615,In_464);
and U247 (N_247,In_556,In_701);
nand U248 (N_248,In_484,In_13);
nand U249 (N_249,In_352,In_166);
nor U250 (N_250,In_362,In_147);
nand U251 (N_251,In_639,In_646);
nor U252 (N_252,In_398,In_533);
nand U253 (N_253,In_65,In_577);
and U254 (N_254,In_88,In_121);
and U255 (N_255,In_679,In_612);
or U256 (N_256,In_289,In_124);
xnor U257 (N_257,In_391,In_746);
and U258 (N_258,In_521,In_542);
nand U259 (N_259,In_280,In_1);
nand U260 (N_260,In_446,In_6);
nor U261 (N_261,In_564,In_496);
nand U262 (N_262,In_725,In_604);
nor U263 (N_263,In_432,In_399);
nand U264 (N_264,In_582,In_263);
nor U265 (N_265,In_117,In_705);
nor U266 (N_266,In_437,In_433);
and U267 (N_267,In_331,In_480);
and U268 (N_268,In_330,In_344);
nor U269 (N_269,In_138,In_2);
and U270 (N_270,In_323,In_429);
or U271 (N_271,In_314,In_492);
and U272 (N_272,In_361,In_108);
or U273 (N_273,In_318,In_543);
nor U274 (N_274,In_458,In_342);
and U275 (N_275,In_338,In_450);
nor U276 (N_276,In_243,In_590);
nand U277 (N_277,In_445,In_284);
or U278 (N_278,In_276,In_691);
and U279 (N_279,In_614,In_489);
and U280 (N_280,In_462,In_591);
nor U281 (N_281,In_513,In_235);
nand U282 (N_282,In_548,In_149);
nand U283 (N_283,In_700,In_382);
nand U284 (N_284,In_475,In_296);
and U285 (N_285,In_181,In_516);
and U286 (N_286,In_365,In_620);
or U287 (N_287,In_128,In_244);
nand U288 (N_288,In_666,In_317);
nand U289 (N_289,In_68,In_734);
nand U290 (N_290,In_163,In_133);
nor U291 (N_291,In_576,In_618);
or U292 (N_292,In_204,In_370);
and U293 (N_293,In_48,In_660);
nand U294 (N_294,In_283,In_381);
nor U295 (N_295,In_45,In_499);
nor U296 (N_296,In_54,In_375);
or U297 (N_297,In_111,In_460);
or U298 (N_298,In_401,In_258);
or U299 (N_299,In_81,In_223);
nor U300 (N_300,In_635,In_519);
nand U301 (N_301,In_600,In_190);
and U302 (N_302,In_237,In_12);
nand U303 (N_303,In_191,In_583);
nand U304 (N_304,In_389,In_201);
nor U305 (N_305,In_7,In_406);
xnor U306 (N_306,In_99,In_107);
or U307 (N_307,In_439,In_262);
xnor U308 (N_308,In_61,In_728);
and U309 (N_309,In_152,In_438);
and U310 (N_310,In_655,In_22);
xor U311 (N_311,In_90,In_250);
or U312 (N_312,In_278,In_308);
and U313 (N_313,In_526,In_738);
nand U314 (N_314,In_531,In_67);
or U315 (N_315,In_585,In_743);
or U316 (N_316,In_132,In_80);
nor U317 (N_317,In_298,In_56);
or U318 (N_318,In_469,In_617);
nand U319 (N_319,In_302,In_94);
and U320 (N_320,In_629,In_610);
and U321 (N_321,In_534,In_336);
nor U322 (N_322,In_18,In_270);
or U323 (N_323,In_194,In_522);
nor U324 (N_324,In_372,In_613);
or U325 (N_325,In_385,In_454);
or U326 (N_326,In_120,In_257);
nor U327 (N_327,In_387,In_234);
nand U328 (N_328,In_72,In_131);
nor U329 (N_329,In_624,In_596);
and U330 (N_330,In_559,In_195);
nor U331 (N_331,In_671,In_544);
nand U332 (N_332,In_187,In_228);
or U333 (N_333,In_676,In_623);
and U334 (N_334,In_595,In_36);
nor U335 (N_335,In_425,In_538);
and U336 (N_336,In_55,In_502);
or U337 (N_337,In_349,In_334);
or U338 (N_338,In_193,In_141);
and U339 (N_339,In_346,In_35);
and U340 (N_340,In_440,In_167);
nand U341 (N_341,In_597,In_586);
and U342 (N_342,In_453,In_561);
or U343 (N_343,In_264,In_717);
nor U344 (N_344,In_637,In_218);
or U345 (N_345,In_59,In_359);
and U346 (N_346,In_275,In_153);
nand U347 (N_347,In_606,In_448);
nor U348 (N_348,In_30,In_75);
nand U349 (N_349,In_709,In_82);
xnor U350 (N_350,In_213,In_642);
or U351 (N_351,In_441,In_366);
and U352 (N_352,In_101,In_494);
or U353 (N_353,In_497,In_122);
nand U354 (N_354,In_471,In_198);
or U355 (N_355,In_413,In_210);
and U356 (N_356,In_353,In_517);
and U357 (N_357,In_609,In_394);
nand U358 (N_358,In_203,In_182);
nand U359 (N_359,In_125,In_532);
nor U360 (N_360,In_311,In_291);
nand U361 (N_361,In_528,In_566);
xor U362 (N_362,In_581,In_520);
or U363 (N_363,In_109,In_222);
nor U364 (N_364,In_692,In_569);
or U365 (N_365,In_628,In_680);
nor U366 (N_366,In_722,In_219);
or U367 (N_367,In_622,In_742);
or U368 (N_368,In_711,In_699);
nor U369 (N_369,In_644,In_304);
or U370 (N_370,In_123,In_46);
or U371 (N_371,In_185,In_281);
nor U372 (N_372,In_455,In_473);
nor U373 (N_373,In_337,In_397);
nor U374 (N_374,In_405,In_329);
and U375 (N_375,In_704,In_637);
nor U376 (N_376,In_15,In_494);
nor U377 (N_377,In_45,In_336);
or U378 (N_378,In_273,In_478);
nor U379 (N_379,In_66,In_171);
nand U380 (N_380,In_29,In_155);
or U381 (N_381,In_20,In_477);
and U382 (N_382,In_454,In_727);
nand U383 (N_383,In_686,In_584);
or U384 (N_384,In_520,In_530);
or U385 (N_385,In_62,In_36);
or U386 (N_386,In_67,In_208);
nor U387 (N_387,In_45,In_169);
nand U388 (N_388,In_367,In_114);
or U389 (N_389,In_169,In_407);
and U390 (N_390,In_77,In_58);
and U391 (N_391,In_259,In_732);
or U392 (N_392,In_748,In_41);
nor U393 (N_393,In_527,In_378);
or U394 (N_394,In_746,In_119);
nor U395 (N_395,In_674,In_80);
or U396 (N_396,In_82,In_316);
or U397 (N_397,In_559,In_107);
or U398 (N_398,In_393,In_79);
and U399 (N_399,In_263,In_30);
nand U400 (N_400,In_246,In_493);
or U401 (N_401,In_133,In_544);
nand U402 (N_402,In_354,In_62);
and U403 (N_403,In_681,In_425);
or U404 (N_404,In_246,In_167);
nand U405 (N_405,In_624,In_670);
nor U406 (N_406,In_327,In_448);
nor U407 (N_407,In_742,In_20);
and U408 (N_408,In_483,In_661);
and U409 (N_409,In_518,In_407);
and U410 (N_410,In_63,In_641);
nor U411 (N_411,In_268,In_466);
nor U412 (N_412,In_737,In_671);
or U413 (N_413,In_224,In_489);
nand U414 (N_414,In_114,In_540);
nand U415 (N_415,In_729,In_276);
and U416 (N_416,In_712,In_324);
nor U417 (N_417,In_244,In_295);
or U418 (N_418,In_379,In_166);
or U419 (N_419,In_419,In_594);
or U420 (N_420,In_645,In_239);
nand U421 (N_421,In_366,In_678);
nor U422 (N_422,In_599,In_721);
and U423 (N_423,In_570,In_153);
and U424 (N_424,In_578,In_346);
and U425 (N_425,In_439,In_424);
nand U426 (N_426,In_31,In_429);
nand U427 (N_427,In_462,In_627);
nand U428 (N_428,In_268,In_264);
or U429 (N_429,In_140,In_246);
nand U430 (N_430,In_166,In_204);
nor U431 (N_431,In_375,In_518);
nand U432 (N_432,In_733,In_684);
nor U433 (N_433,In_203,In_53);
nand U434 (N_434,In_4,In_414);
xnor U435 (N_435,In_576,In_2);
or U436 (N_436,In_500,In_44);
and U437 (N_437,In_595,In_628);
and U438 (N_438,In_328,In_606);
or U439 (N_439,In_131,In_720);
nand U440 (N_440,In_75,In_143);
nor U441 (N_441,In_602,In_194);
nand U442 (N_442,In_426,In_80);
nor U443 (N_443,In_468,In_731);
and U444 (N_444,In_665,In_365);
and U445 (N_445,In_277,In_415);
nor U446 (N_446,In_565,In_511);
or U447 (N_447,In_348,In_350);
nor U448 (N_448,In_72,In_0);
nor U449 (N_449,In_643,In_646);
or U450 (N_450,In_674,In_447);
or U451 (N_451,In_365,In_627);
and U452 (N_452,In_197,In_214);
or U453 (N_453,In_391,In_131);
nor U454 (N_454,In_316,In_376);
xor U455 (N_455,In_306,In_737);
nor U456 (N_456,In_685,In_466);
and U457 (N_457,In_24,In_554);
nand U458 (N_458,In_111,In_299);
nor U459 (N_459,In_563,In_8);
nand U460 (N_460,In_84,In_43);
nor U461 (N_461,In_268,In_157);
or U462 (N_462,In_458,In_656);
or U463 (N_463,In_68,In_176);
nand U464 (N_464,In_531,In_208);
or U465 (N_465,In_690,In_577);
nor U466 (N_466,In_746,In_280);
or U467 (N_467,In_20,In_286);
or U468 (N_468,In_53,In_588);
nor U469 (N_469,In_151,In_276);
nand U470 (N_470,In_25,In_361);
and U471 (N_471,In_199,In_494);
or U472 (N_472,In_628,In_418);
nor U473 (N_473,In_63,In_529);
nand U474 (N_474,In_286,In_301);
or U475 (N_475,In_51,In_433);
nor U476 (N_476,In_8,In_325);
nand U477 (N_477,In_158,In_726);
or U478 (N_478,In_126,In_407);
and U479 (N_479,In_294,In_594);
nor U480 (N_480,In_563,In_116);
nand U481 (N_481,In_632,In_237);
and U482 (N_482,In_32,In_646);
xor U483 (N_483,In_91,In_469);
or U484 (N_484,In_527,In_266);
and U485 (N_485,In_32,In_624);
or U486 (N_486,In_516,In_651);
and U487 (N_487,In_222,In_52);
nor U488 (N_488,In_82,In_347);
and U489 (N_489,In_361,In_405);
nor U490 (N_490,In_686,In_387);
or U491 (N_491,In_432,In_37);
nor U492 (N_492,In_78,In_16);
nand U493 (N_493,In_721,In_488);
or U494 (N_494,In_183,In_123);
nand U495 (N_495,In_251,In_168);
or U496 (N_496,In_726,In_202);
nor U497 (N_497,In_693,In_265);
nor U498 (N_498,In_106,In_204);
nor U499 (N_499,In_0,In_208);
nor U500 (N_500,In_483,In_160);
and U501 (N_501,In_553,In_210);
and U502 (N_502,In_60,In_89);
or U503 (N_503,In_32,In_507);
xor U504 (N_504,In_443,In_316);
and U505 (N_505,In_377,In_312);
nand U506 (N_506,In_323,In_517);
nor U507 (N_507,In_749,In_462);
and U508 (N_508,In_451,In_603);
or U509 (N_509,In_689,In_184);
nand U510 (N_510,In_167,In_117);
nand U511 (N_511,In_101,In_604);
or U512 (N_512,In_705,In_248);
nand U513 (N_513,In_448,In_384);
xor U514 (N_514,In_138,In_737);
and U515 (N_515,In_416,In_224);
and U516 (N_516,In_734,In_700);
or U517 (N_517,In_210,In_389);
nand U518 (N_518,In_5,In_239);
and U519 (N_519,In_87,In_72);
nor U520 (N_520,In_115,In_23);
nand U521 (N_521,In_532,In_19);
nand U522 (N_522,In_743,In_398);
and U523 (N_523,In_410,In_377);
nand U524 (N_524,In_87,In_201);
nor U525 (N_525,In_355,In_147);
xnor U526 (N_526,In_394,In_321);
nand U527 (N_527,In_213,In_710);
and U528 (N_528,In_608,In_344);
nand U529 (N_529,In_229,In_304);
nand U530 (N_530,In_247,In_228);
and U531 (N_531,In_112,In_506);
nor U532 (N_532,In_502,In_235);
nand U533 (N_533,In_520,In_432);
nand U534 (N_534,In_477,In_322);
nor U535 (N_535,In_545,In_629);
and U536 (N_536,In_217,In_105);
nor U537 (N_537,In_153,In_317);
nand U538 (N_538,In_209,In_580);
nand U539 (N_539,In_666,In_109);
or U540 (N_540,In_545,In_729);
and U541 (N_541,In_741,In_388);
or U542 (N_542,In_67,In_661);
and U543 (N_543,In_7,In_360);
or U544 (N_544,In_331,In_599);
or U545 (N_545,In_563,In_445);
or U546 (N_546,In_452,In_249);
nor U547 (N_547,In_643,In_507);
nand U548 (N_548,In_4,In_290);
nor U549 (N_549,In_698,In_132);
nor U550 (N_550,In_75,In_661);
and U551 (N_551,In_500,In_118);
or U552 (N_552,In_543,In_524);
and U553 (N_553,In_91,In_354);
or U554 (N_554,In_692,In_275);
nor U555 (N_555,In_185,In_494);
nand U556 (N_556,In_84,In_586);
nor U557 (N_557,In_64,In_488);
and U558 (N_558,In_614,In_611);
nand U559 (N_559,In_535,In_79);
or U560 (N_560,In_587,In_698);
nor U561 (N_561,In_635,In_280);
and U562 (N_562,In_332,In_25);
or U563 (N_563,In_214,In_507);
nand U564 (N_564,In_484,In_144);
nor U565 (N_565,In_212,In_606);
and U566 (N_566,In_412,In_409);
nor U567 (N_567,In_332,In_88);
and U568 (N_568,In_427,In_251);
or U569 (N_569,In_364,In_321);
or U570 (N_570,In_33,In_509);
nand U571 (N_571,In_100,In_311);
nand U572 (N_572,In_225,In_369);
or U573 (N_573,In_607,In_391);
nor U574 (N_574,In_390,In_652);
and U575 (N_575,In_320,In_469);
nor U576 (N_576,In_553,In_558);
nor U577 (N_577,In_311,In_244);
or U578 (N_578,In_707,In_551);
nor U579 (N_579,In_352,In_403);
nand U580 (N_580,In_611,In_601);
nand U581 (N_581,In_368,In_705);
and U582 (N_582,In_732,In_40);
nand U583 (N_583,In_373,In_310);
nand U584 (N_584,In_524,In_27);
nor U585 (N_585,In_66,In_576);
or U586 (N_586,In_287,In_20);
nand U587 (N_587,In_240,In_197);
nor U588 (N_588,In_139,In_123);
nor U589 (N_589,In_617,In_411);
or U590 (N_590,In_577,In_458);
nand U591 (N_591,In_532,In_180);
and U592 (N_592,In_118,In_128);
or U593 (N_593,In_591,In_625);
or U594 (N_594,In_427,In_589);
or U595 (N_595,In_169,In_464);
or U596 (N_596,In_585,In_450);
and U597 (N_597,In_607,In_542);
and U598 (N_598,In_361,In_163);
nand U599 (N_599,In_109,In_3);
xor U600 (N_600,In_95,In_285);
nand U601 (N_601,In_538,In_72);
and U602 (N_602,In_62,In_647);
and U603 (N_603,In_525,In_625);
or U604 (N_604,In_695,In_446);
or U605 (N_605,In_229,In_410);
or U606 (N_606,In_377,In_279);
or U607 (N_607,In_375,In_697);
or U608 (N_608,In_56,In_697);
and U609 (N_609,In_60,In_217);
nand U610 (N_610,In_498,In_91);
or U611 (N_611,In_595,In_539);
nor U612 (N_612,In_296,In_706);
and U613 (N_613,In_456,In_380);
or U614 (N_614,In_23,In_718);
and U615 (N_615,In_696,In_435);
or U616 (N_616,In_106,In_681);
or U617 (N_617,In_320,In_105);
and U618 (N_618,In_53,In_523);
nor U619 (N_619,In_149,In_243);
and U620 (N_620,In_551,In_452);
nor U621 (N_621,In_678,In_175);
or U622 (N_622,In_516,In_105);
nor U623 (N_623,In_54,In_199);
nand U624 (N_624,In_158,In_330);
and U625 (N_625,In_520,In_304);
and U626 (N_626,In_74,In_517);
nor U627 (N_627,In_57,In_668);
nor U628 (N_628,In_24,In_119);
nand U629 (N_629,In_417,In_290);
or U630 (N_630,In_150,In_575);
nand U631 (N_631,In_382,In_200);
nand U632 (N_632,In_357,In_533);
and U633 (N_633,In_592,In_735);
or U634 (N_634,In_81,In_490);
or U635 (N_635,In_202,In_218);
and U636 (N_636,In_100,In_77);
and U637 (N_637,In_259,In_192);
xor U638 (N_638,In_540,In_666);
nor U639 (N_639,In_546,In_482);
nor U640 (N_640,In_522,In_219);
nand U641 (N_641,In_583,In_514);
or U642 (N_642,In_652,In_691);
and U643 (N_643,In_4,In_668);
or U644 (N_644,In_488,In_154);
or U645 (N_645,In_714,In_691);
or U646 (N_646,In_682,In_57);
or U647 (N_647,In_603,In_727);
or U648 (N_648,In_610,In_745);
and U649 (N_649,In_9,In_525);
nor U650 (N_650,In_650,In_87);
or U651 (N_651,In_299,In_300);
and U652 (N_652,In_260,In_27);
or U653 (N_653,In_43,In_748);
nor U654 (N_654,In_50,In_254);
nor U655 (N_655,In_544,In_721);
and U656 (N_656,In_39,In_73);
and U657 (N_657,In_135,In_679);
nand U658 (N_658,In_336,In_527);
or U659 (N_659,In_253,In_290);
or U660 (N_660,In_394,In_462);
or U661 (N_661,In_513,In_590);
nand U662 (N_662,In_48,In_576);
or U663 (N_663,In_569,In_516);
and U664 (N_664,In_419,In_733);
or U665 (N_665,In_479,In_599);
and U666 (N_666,In_550,In_600);
nor U667 (N_667,In_691,In_387);
nand U668 (N_668,In_184,In_537);
nor U669 (N_669,In_558,In_97);
and U670 (N_670,In_593,In_166);
and U671 (N_671,In_208,In_216);
nor U672 (N_672,In_583,In_314);
xnor U673 (N_673,In_118,In_438);
and U674 (N_674,In_400,In_604);
nor U675 (N_675,In_189,In_514);
and U676 (N_676,In_348,In_428);
nor U677 (N_677,In_413,In_483);
nand U678 (N_678,In_139,In_173);
and U679 (N_679,In_663,In_558);
and U680 (N_680,In_111,In_648);
and U681 (N_681,In_71,In_46);
nand U682 (N_682,In_461,In_332);
nor U683 (N_683,In_89,In_646);
or U684 (N_684,In_625,In_21);
xor U685 (N_685,In_693,In_15);
or U686 (N_686,In_420,In_732);
nand U687 (N_687,In_112,In_585);
and U688 (N_688,In_686,In_546);
nor U689 (N_689,In_650,In_679);
xor U690 (N_690,In_47,In_551);
nand U691 (N_691,In_605,In_595);
and U692 (N_692,In_677,In_84);
or U693 (N_693,In_661,In_561);
nand U694 (N_694,In_278,In_11);
xnor U695 (N_695,In_261,In_184);
and U696 (N_696,In_503,In_549);
nor U697 (N_697,In_167,In_554);
and U698 (N_698,In_112,In_318);
and U699 (N_699,In_199,In_327);
or U700 (N_700,In_277,In_718);
nor U701 (N_701,In_37,In_531);
or U702 (N_702,In_461,In_47);
nand U703 (N_703,In_46,In_738);
nor U704 (N_704,In_160,In_153);
nand U705 (N_705,In_87,In_528);
or U706 (N_706,In_422,In_282);
nand U707 (N_707,In_747,In_484);
and U708 (N_708,In_10,In_484);
nor U709 (N_709,In_88,In_521);
and U710 (N_710,In_600,In_666);
and U711 (N_711,In_119,In_675);
or U712 (N_712,In_486,In_190);
or U713 (N_713,In_390,In_235);
or U714 (N_714,In_181,In_256);
and U715 (N_715,In_190,In_31);
nand U716 (N_716,In_66,In_25);
nor U717 (N_717,In_255,In_165);
nor U718 (N_718,In_629,In_707);
nor U719 (N_719,In_675,In_718);
and U720 (N_720,In_677,In_440);
nand U721 (N_721,In_370,In_559);
nor U722 (N_722,In_354,In_631);
or U723 (N_723,In_148,In_66);
or U724 (N_724,In_415,In_218);
nor U725 (N_725,In_432,In_735);
nand U726 (N_726,In_473,In_271);
and U727 (N_727,In_310,In_164);
nor U728 (N_728,In_172,In_398);
xnor U729 (N_729,In_47,In_106);
and U730 (N_730,In_3,In_597);
and U731 (N_731,In_561,In_278);
nor U732 (N_732,In_627,In_465);
nand U733 (N_733,In_121,In_655);
or U734 (N_734,In_747,In_641);
and U735 (N_735,In_263,In_321);
nor U736 (N_736,In_299,In_560);
nand U737 (N_737,In_93,In_412);
nand U738 (N_738,In_693,In_121);
nor U739 (N_739,In_606,In_503);
nand U740 (N_740,In_644,In_104);
or U741 (N_741,In_738,In_665);
nor U742 (N_742,In_540,In_582);
or U743 (N_743,In_620,In_651);
or U744 (N_744,In_512,In_160);
or U745 (N_745,In_548,In_108);
or U746 (N_746,In_523,In_236);
nand U747 (N_747,In_619,In_200);
and U748 (N_748,In_414,In_114);
and U749 (N_749,In_559,In_146);
nor U750 (N_750,In_596,In_474);
nor U751 (N_751,In_384,In_501);
xnor U752 (N_752,In_93,In_657);
nand U753 (N_753,In_38,In_563);
and U754 (N_754,In_39,In_174);
nand U755 (N_755,In_126,In_121);
nor U756 (N_756,In_327,In_715);
and U757 (N_757,In_330,In_31);
xnor U758 (N_758,In_7,In_387);
and U759 (N_759,In_195,In_95);
and U760 (N_760,In_462,In_150);
nor U761 (N_761,In_74,In_478);
and U762 (N_762,In_569,In_84);
nand U763 (N_763,In_624,In_683);
nor U764 (N_764,In_539,In_653);
nand U765 (N_765,In_4,In_213);
nor U766 (N_766,In_441,In_49);
and U767 (N_767,In_745,In_81);
nand U768 (N_768,In_293,In_525);
or U769 (N_769,In_117,In_267);
nor U770 (N_770,In_125,In_129);
or U771 (N_771,In_719,In_704);
or U772 (N_772,In_514,In_147);
and U773 (N_773,In_427,In_52);
and U774 (N_774,In_169,In_149);
nor U775 (N_775,In_221,In_576);
and U776 (N_776,In_58,In_544);
or U777 (N_777,In_499,In_562);
or U778 (N_778,In_665,In_676);
and U779 (N_779,In_187,In_272);
xor U780 (N_780,In_351,In_195);
and U781 (N_781,In_335,In_318);
nand U782 (N_782,In_232,In_312);
nor U783 (N_783,In_425,In_252);
and U784 (N_784,In_610,In_235);
or U785 (N_785,In_700,In_556);
and U786 (N_786,In_336,In_739);
or U787 (N_787,In_674,In_374);
nand U788 (N_788,In_621,In_315);
and U789 (N_789,In_17,In_319);
and U790 (N_790,In_170,In_609);
nand U791 (N_791,In_38,In_35);
xor U792 (N_792,In_668,In_530);
nor U793 (N_793,In_220,In_489);
nand U794 (N_794,In_713,In_623);
and U795 (N_795,In_482,In_367);
nor U796 (N_796,In_594,In_188);
nor U797 (N_797,In_365,In_166);
nor U798 (N_798,In_121,In_118);
and U799 (N_799,In_292,In_286);
nor U800 (N_800,In_17,In_358);
nand U801 (N_801,In_192,In_506);
nor U802 (N_802,In_658,In_327);
and U803 (N_803,In_206,In_238);
and U804 (N_804,In_634,In_445);
and U805 (N_805,In_726,In_511);
and U806 (N_806,In_19,In_602);
or U807 (N_807,In_57,In_34);
nand U808 (N_808,In_461,In_622);
or U809 (N_809,In_463,In_408);
or U810 (N_810,In_244,In_378);
nand U811 (N_811,In_547,In_643);
or U812 (N_812,In_16,In_413);
nor U813 (N_813,In_646,In_283);
and U814 (N_814,In_301,In_647);
and U815 (N_815,In_216,In_415);
or U816 (N_816,In_592,In_721);
and U817 (N_817,In_137,In_229);
and U818 (N_818,In_331,In_236);
nor U819 (N_819,In_272,In_63);
and U820 (N_820,In_251,In_262);
and U821 (N_821,In_528,In_53);
and U822 (N_822,In_222,In_476);
nand U823 (N_823,In_59,In_191);
nand U824 (N_824,In_458,In_457);
and U825 (N_825,In_422,In_721);
and U826 (N_826,In_546,In_423);
and U827 (N_827,In_642,In_558);
or U828 (N_828,In_169,In_277);
nand U829 (N_829,In_408,In_647);
nor U830 (N_830,In_474,In_449);
and U831 (N_831,In_681,In_169);
nand U832 (N_832,In_212,In_660);
and U833 (N_833,In_268,In_253);
and U834 (N_834,In_534,In_174);
or U835 (N_835,In_524,In_678);
and U836 (N_836,In_79,In_251);
or U837 (N_837,In_178,In_132);
nor U838 (N_838,In_137,In_699);
or U839 (N_839,In_125,In_19);
or U840 (N_840,In_415,In_572);
nor U841 (N_841,In_506,In_66);
nor U842 (N_842,In_712,In_142);
or U843 (N_843,In_328,In_276);
nand U844 (N_844,In_356,In_153);
nor U845 (N_845,In_398,In_744);
nand U846 (N_846,In_47,In_299);
or U847 (N_847,In_287,In_635);
nand U848 (N_848,In_591,In_590);
nor U849 (N_849,In_214,In_94);
or U850 (N_850,In_546,In_715);
or U851 (N_851,In_311,In_542);
and U852 (N_852,In_177,In_241);
nor U853 (N_853,In_14,In_537);
nor U854 (N_854,In_90,In_721);
or U855 (N_855,In_19,In_320);
nor U856 (N_856,In_554,In_639);
nor U857 (N_857,In_690,In_236);
or U858 (N_858,In_427,In_105);
and U859 (N_859,In_151,In_48);
nor U860 (N_860,In_167,In_483);
nand U861 (N_861,In_0,In_214);
nor U862 (N_862,In_479,In_0);
or U863 (N_863,In_218,In_599);
and U864 (N_864,In_478,In_156);
or U865 (N_865,In_190,In_513);
nor U866 (N_866,In_177,In_165);
or U867 (N_867,In_433,In_65);
and U868 (N_868,In_552,In_517);
nor U869 (N_869,In_208,In_311);
xnor U870 (N_870,In_705,In_460);
nand U871 (N_871,In_186,In_606);
or U872 (N_872,In_653,In_402);
nand U873 (N_873,In_52,In_21);
nor U874 (N_874,In_726,In_383);
nand U875 (N_875,In_619,In_268);
and U876 (N_876,In_114,In_493);
nor U877 (N_877,In_380,In_510);
nor U878 (N_878,In_694,In_673);
nor U879 (N_879,In_334,In_360);
nor U880 (N_880,In_52,In_301);
nor U881 (N_881,In_715,In_50);
nor U882 (N_882,In_402,In_278);
or U883 (N_883,In_200,In_46);
nand U884 (N_884,In_245,In_293);
and U885 (N_885,In_261,In_205);
nor U886 (N_886,In_697,In_454);
nand U887 (N_887,In_40,In_430);
and U888 (N_888,In_71,In_77);
nor U889 (N_889,In_57,In_480);
or U890 (N_890,In_371,In_715);
nor U891 (N_891,In_650,In_253);
nor U892 (N_892,In_116,In_431);
nand U893 (N_893,In_210,In_507);
nand U894 (N_894,In_7,In_178);
and U895 (N_895,In_640,In_199);
xnor U896 (N_896,In_193,In_602);
nand U897 (N_897,In_328,In_353);
or U898 (N_898,In_61,In_88);
or U899 (N_899,In_460,In_44);
and U900 (N_900,In_230,In_711);
nor U901 (N_901,In_453,In_494);
or U902 (N_902,In_559,In_116);
nor U903 (N_903,In_527,In_186);
and U904 (N_904,In_658,In_86);
and U905 (N_905,In_428,In_598);
and U906 (N_906,In_213,In_179);
nand U907 (N_907,In_499,In_519);
nor U908 (N_908,In_50,In_529);
nor U909 (N_909,In_55,In_56);
and U910 (N_910,In_630,In_672);
nor U911 (N_911,In_399,In_617);
and U912 (N_912,In_351,In_407);
nand U913 (N_913,In_636,In_131);
and U914 (N_914,In_595,In_122);
and U915 (N_915,In_749,In_281);
or U916 (N_916,In_71,In_352);
xor U917 (N_917,In_620,In_522);
and U918 (N_918,In_394,In_657);
nor U919 (N_919,In_547,In_65);
nand U920 (N_920,In_731,In_409);
and U921 (N_921,In_7,In_348);
or U922 (N_922,In_124,In_463);
xnor U923 (N_923,In_640,In_224);
or U924 (N_924,In_92,In_389);
or U925 (N_925,In_41,In_452);
nand U926 (N_926,In_191,In_6);
or U927 (N_927,In_281,In_723);
nor U928 (N_928,In_737,In_160);
or U929 (N_929,In_92,In_290);
and U930 (N_930,In_511,In_725);
and U931 (N_931,In_332,In_290);
and U932 (N_932,In_580,In_237);
nand U933 (N_933,In_314,In_31);
nand U934 (N_934,In_211,In_492);
or U935 (N_935,In_347,In_544);
and U936 (N_936,In_738,In_435);
nand U937 (N_937,In_589,In_326);
and U938 (N_938,In_709,In_84);
nor U939 (N_939,In_471,In_735);
and U940 (N_940,In_613,In_166);
and U941 (N_941,In_205,In_521);
nor U942 (N_942,In_1,In_2);
nand U943 (N_943,In_444,In_213);
and U944 (N_944,In_247,In_284);
and U945 (N_945,In_660,In_356);
or U946 (N_946,In_506,In_702);
nand U947 (N_947,In_684,In_557);
nor U948 (N_948,In_211,In_435);
and U949 (N_949,In_152,In_709);
nand U950 (N_950,In_41,In_22);
and U951 (N_951,In_579,In_402);
and U952 (N_952,In_630,In_128);
or U953 (N_953,In_726,In_561);
or U954 (N_954,In_575,In_252);
nor U955 (N_955,In_440,In_83);
nand U956 (N_956,In_505,In_153);
and U957 (N_957,In_154,In_636);
nor U958 (N_958,In_439,In_447);
nor U959 (N_959,In_462,In_263);
nand U960 (N_960,In_367,In_269);
and U961 (N_961,In_602,In_709);
nor U962 (N_962,In_131,In_93);
nor U963 (N_963,In_161,In_616);
or U964 (N_964,In_624,In_590);
or U965 (N_965,In_351,In_555);
or U966 (N_966,In_694,In_83);
nand U967 (N_967,In_279,In_38);
nand U968 (N_968,In_376,In_199);
and U969 (N_969,In_352,In_108);
nand U970 (N_970,In_705,In_482);
nor U971 (N_971,In_623,In_524);
nand U972 (N_972,In_334,In_303);
and U973 (N_973,In_358,In_366);
or U974 (N_974,In_408,In_710);
nand U975 (N_975,In_582,In_702);
xor U976 (N_976,In_224,In_470);
nor U977 (N_977,In_607,In_460);
or U978 (N_978,In_311,In_58);
or U979 (N_979,In_29,In_694);
xnor U980 (N_980,In_308,In_587);
nand U981 (N_981,In_514,In_385);
or U982 (N_982,In_48,In_667);
or U983 (N_983,In_732,In_422);
or U984 (N_984,In_629,In_386);
nand U985 (N_985,In_82,In_625);
nor U986 (N_986,In_16,In_334);
or U987 (N_987,In_425,In_0);
or U988 (N_988,In_273,In_532);
and U989 (N_989,In_452,In_5);
or U990 (N_990,In_437,In_630);
and U991 (N_991,In_591,In_728);
or U992 (N_992,In_671,In_44);
nand U993 (N_993,In_569,In_679);
and U994 (N_994,In_468,In_139);
nor U995 (N_995,In_474,In_625);
or U996 (N_996,In_111,In_531);
nand U997 (N_997,In_283,In_58);
or U998 (N_998,In_513,In_275);
nor U999 (N_999,In_664,In_224);
nand U1000 (N_1000,In_260,In_352);
and U1001 (N_1001,In_60,In_143);
nand U1002 (N_1002,In_68,In_270);
nor U1003 (N_1003,In_309,In_10);
nor U1004 (N_1004,In_66,In_541);
nand U1005 (N_1005,In_629,In_90);
nand U1006 (N_1006,In_425,In_520);
and U1007 (N_1007,In_51,In_409);
nor U1008 (N_1008,In_201,In_568);
nand U1009 (N_1009,In_325,In_272);
or U1010 (N_1010,In_627,In_201);
nor U1011 (N_1011,In_464,In_585);
xnor U1012 (N_1012,In_197,In_230);
and U1013 (N_1013,In_200,In_127);
nor U1014 (N_1014,In_47,In_493);
nor U1015 (N_1015,In_616,In_608);
nor U1016 (N_1016,In_343,In_743);
and U1017 (N_1017,In_286,In_719);
nor U1018 (N_1018,In_713,In_318);
or U1019 (N_1019,In_370,In_251);
and U1020 (N_1020,In_618,In_121);
or U1021 (N_1021,In_614,In_53);
and U1022 (N_1022,In_617,In_491);
or U1023 (N_1023,In_533,In_232);
or U1024 (N_1024,In_642,In_127);
or U1025 (N_1025,In_266,In_708);
and U1026 (N_1026,In_357,In_480);
or U1027 (N_1027,In_578,In_90);
or U1028 (N_1028,In_226,In_228);
and U1029 (N_1029,In_413,In_91);
and U1030 (N_1030,In_686,In_594);
nor U1031 (N_1031,In_570,In_144);
and U1032 (N_1032,In_178,In_118);
and U1033 (N_1033,In_396,In_720);
nand U1034 (N_1034,In_135,In_508);
nand U1035 (N_1035,In_570,In_562);
nor U1036 (N_1036,In_364,In_523);
and U1037 (N_1037,In_613,In_234);
or U1038 (N_1038,In_282,In_620);
or U1039 (N_1039,In_698,In_133);
or U1040 (N_1040,In_724,In_513);
nand U1041 (N_1041,In_612,In_197);
or U1042 (N_1042,In_161,In_193);
nand U1043 (N_1043,In_165,In_438);
nor U1044 (N_1044,In_591,In_45);
xnor U1045 (N_1045,In_247,In_362);
nand U1046 (N_1046,In_61,In_472);
nand U1047 (N_1047,In_671,In_115);
nor U1048 (N_1048,In_535,In_677);
nand U1049 (N_1049,In_435,In_598);
nor U1050 (N_1050,In_714,In_119);
or U1051 (N_1051,In_502,In_56);
nor U1052 (N_1052,In_42,In_554);
nor U1053 (N_1053,In_267,In_4);
and U1054 (N_1054,In_176,In_189);
nor U1055 (N_1055,In_508,In_350);
nand U1056 (N_1056,In_34,In_297);
xnor U1057 (N_1057,In_643,In_621);
nor U1058 (N_1058,In_313,In_139);
nand U1059 (N_1059,In_309,In_544);
nor U1060 (N_1060,In_478,In_416);
or U1061 (N_1061,In_48,In_544);
and U1062 (N_1062,In_464,In_603);
nor U1063 (N_1063,In_177,In_730);
and U1064 (N_1064,In_455,In_466);
nor U1065 (N_1065,In_432,In_367);
nand U1066 (N_1066,In_76,In_487);
nor U1067 (N_1067,In_236,In_198);
or U1068 (N_1068,In_696,In_245);
or U1069 (N_1069,In_136,In_472);
and U1070 (N_1070,In_248,In_400);
nor U1071 (N_1071,In_490,In_474);
nor U1072 (N_1072,In_729,In_141);
or U1073 (N_1073,In_693,In_35);
nand U1074 (N_1074,In_162,In_506);
or U1075 (N_1075,In_116,In_408);
nand U1076 (N_1076,In_422,In_681);
or U1077 (N_1077,In_631,In_458);
or U1078 (N_1078,In_166,In_305);
and U1079 (N_1079,In_339,In_419);
nand U1080 (N_1080,In_378,In_630);
xnor U1081 (N_1081,In_625,In_455);
nand U1082 (N_1082,In_206,In_552);
nand U1083 (N_1083,In_731,In_660);
nand U1084 (N_1084,In_497,In_234);
or U1085 (N_1085,In_737,In_286);
or U1086 (N_1086,In_564,In_739);
or U1087 (N_1087,In_443,In_411);
nand U1088 (N_1088,In_658,In_578);
nand U1089 (N_1089,In_406,In_167);
nor U1090 (N_1090,In_334,In_209);
xor U1091 (N_1091,In_540,In_200);
or U1092 (N_1092,In_57,In_424);
and U1093 (N_1093,In_44,In_0);
or U1094 (N_1094,In_667,In_519);
and U1095 (N_1095,In_252,In_368);
nand U1096 (N_1096,In_630,In_185);
and U1097 (N_1097,In_498,In_552);
and U1098 (N_1098,In_291,In_705);
and U1099 (N_1099,In_365,In_355);
nor U1100 (N_1100,In_591,In_209);
nand U1101 (N_1101,In_507,In_685);
nor U1102 (N_1102,In_242,In_372);
and U1103 (N_1103,In_460,In_186);
nand U1104 (N_1104,In_401,In_413);
nand U1105 (N_1105,In_690,In_510);
and U1106 (N_1106,In_116,In_465);
or U1107 (N_1107,In_89,In_43);
and U1108 (N_1108,In_226,In_516);
nor U1109 (N_1109,In_499,In_414);
nor U1110 (N_1110,In_413,In_256);
or U1111 (N_1111,In_71,In_81);
and U1112 (N_1112,In_305,In_652);
and U1113 (N_1113,In_689,In_6);
nor U1114 (N_1114,In_105,In_312);
and U1115 (N_1115,In_277,In_707);
nor U1116 (N_1116,In_471,In_517);
nand U1117 (N_1117,In_603,In_473);
nor U1118 (N_1118,In_631,In_193);
or U1119 (N_1119,In_320,In_125);
or U1120 (N_1120,In_604,In_220);
nor U1121 (N_1121,In_384,In_115);
and U1122 (N_1122,In_598,In_333);
or U1123 (N_1123,In_140,In_301);
or U1124 (N_1124,In_184,In_24);
or U1125 (N_1125,In_734,In_635);
nor U1126 (N_1126,In_499,In_688);
nor U1127 (N_1127,In_731,In_434);
nor U1128 (N_1128,In_407,In_18);
nand U1129 (N_1129,In_254,In_222);
and U1130 (N_1130,In_706,In_576);
and U1131 (N_1131,In_746,In_158);
or U1132 (N_1132,In_719,In_718);
nand U1133 (N_1133,In_703,In_732);
xnor U1134 (N_1134,In_543,In_686);
nand U1135 (N_1135,In_562,In_546);
nor U1136 (N_1136,In_646,In_406);
nand U1137 (N_1137,In_513,In_654);
or U1138 (N_1138,In_715,In_604);
and U1139 (N_1139,In_571,In_354);
or U1140 (N_1140,In_65,In_534);
nor U1141 (N_1141,In_437,In_413);
nor U1142 (N_1142,In_482,In_666);
nand U1143 (N_1143,In_545,In_336);
or U1144 (N_1144,In_372,In_667);
nor U1145 (N_1145,In_406,In_475);
and U1146 (N_1146,In_426,In_417);
and U1147 (N_1147,In_513,In_313);
nor U1148 (N_1148,In_76,In_482);
nand U1149 (N_1149,In_718,In_129);
and U1150 (N_1150,In_512,In_391);
and U1151 (N_1151,In_640,In_434);
or U1152 (N_1152,In_304,In_4);
or U1153 (N_1153,In_399,In_663);
and U1154 (N_1154,In_266,In_740);
and U1155 (N_1155,In_538,In_594);
or U1156 (N_1156,In_83,In_373);
or U1157 (N_1157,In_98,In_687);
nor U1158 (N_1158,In_354,In_537);
nor U1159 (N_1159,In_615,In_451);
nand U1160 (N_1160,In_294,In_483);
and U1161 (N_1161,In_201,In_275);
and U1162 (N_1162,In_421,In_456);
nor U1163 (N_1163,In_165,In_508);
and U1164 (N_1164,In_724,In_23);
and U1165 (N_1165,In_610,In_431);
nor U1166 (N_1166,In_195,In_277);
and U1167 (N_1167,In_295,In_665);
or U1168 (N_1168,In_515,In_366);
or U1169 (N_1169,In_192,In_176);
and U1170 (N_1170,In_384,In_0);
nor U1171 (N_1171,In_427,In_39);
or U1172 (N_1172,In_393,In_616);
xnor U1173 (N_1173,In_492,In_167);
or U1174 (N_1174,In_60,In_572);
or U1175 (N_1175,In_722,In_432);
nand U1176 (N_1176,In_511,In_529);
or U1177 (N_1177,In_414,In_290);
and U1178 (N_1178,In_129,In_541);
and U1179 (N_1179,In_437,In_318);
and U1180 (N_1180,In_565,In_393);
nand U1181 (N_1181,In_678,In_321);
or U1182 (N_1182,In_599,In_543);
and U1183 (N_1183,In_344,In_255);
nand U1184 (N_1184,In_104,In_330);
or U1185 (N_1185,In_150,In_609);
xor U1186 (N_1186,In_634,In_469);
and U1187 (N_1187,In_285,In_570);
or U1188 (N_1188,In_615,In_238);
or U1189 (N_1189,In_231,In_582);
nor U1190 (N_1190,In_617,In_207);
nor U1191 (N_1191,In_610,In_364);
or U1192 (N_1192,In_710,In_111);
nor U1193 (N_1193,In_614,In_189);
or U1194 (N_1194,In_406,In_8);
or U1195 (N_1195,In_520,In_199);
xor U1196 (N_1196,In_719,In_22);
or U1197 (N_1197,In_577,In_400);
nand U1198 (N_1198,In_392,In_736);
nand U1199 (N_1199,In_646,In_480);
xnor U1200 (N_1200,In_137,In_608);
or U1201 (N_1201,In_713,In_524);
nor U1202 (N_1202,In_308,In_288);
nor U1203 (N_1203,In_588,In_306);
nor U1204 (N_1204,In_62,In_408);
nor U1205 (N_1205,In_706,In_329);
or U1206 (N_1206,In_375,In_282);
and U1207 (N_1207,In_222,In_377);
and U1208 (N_1208,In_88,In_0);
or U1209 (N_1209,In_484,In_137);
nor U1210 (N_1210,In_623,In_426);
or U1211 (N_1211,In_426,In_658);
and U1212 (N_1212,In_662,In_364);
nand U1213 (N_1213,In_710,In_157);
or U1214 (N_1214,In_230,In_340);
or U1215 (N_1215,In_92,In_625);
nor U1216 (N_1216,In_577,In_498);
nor U1217 (N_1217,In_444,In_687);
xor U1218 (N_1218,In_208,In_164);
or U1219 (N_1219,In_389,In_577);
nand U1220 (N_1220,In_349,In_429);
nand U1221 (N_1221,In_748,In_114);
nor U1222 (N_1222,In_184,In_355);
nor U1223 (N_1223,In_40,In_3);
and U1224 (N_1224,In_134,In_172);
and U1225 (N_1225,In_24,In_243);
and U1226 (N_1226,In_344,In_130);
and U1227 (N_1227,In_47,In_705);
nor U1228 (N_1228,In_246,In_328);
nor U1229 (N_1229,In_86,In_363);
or U1230 (N_1230,In_489,In_162);
nor U1231 (N_1231,In_571,In_740);
nand U1232 (N_1232,In_203,In_163);
nand U1233 (N_1233,In_696,In_497);
nor U1234 (N_1234,In_86,In_98);
and U1235 (N_1235,In_423,In_716);
and U1236 (N_1236,In_684,In_351);
nor U1237 (N_1237,In_116,In_153);
nand U1238 (N_1238,In_653,In_265);
or U1239 (N_1239,In_158,In_506);
nand U1240 (N_1240,In_747,In_420);
nand U1241 (N_1241,In_59,In_533);
or U1242 (N_1242,In_181,In_55);
nor U1243 (N_1243,In_724,In_581);
and U1244 (N_1244,In_145,In_734);
and U1245 (N_1245,In_133,In_81);
or U1246 (N_1246,In_243,In_72);
nand U1247 (N_1247,In_269,In_295);
xnor U1248 (N_1248,In_335,In_706);
nor U1249 (N_1249,In_379,In_412);
or U1250 (N_1250,In_563,In_673);
or U1251 (N_1251,In_638,In_136);
nor U1252 (N_1252,In_149,In_172);
or U1253 (N_1253,In_546,In_221);
and U1254 (N_1254,In_181,In_455);
nor U1255 (N_1255,In_644,In_409);
nand U1256 (N_1256,In_705,In_149);
nor U1257 (N_1257,In_506,In_371);
nand U1258 (N_1258,In_348,In_261);
or U1259 (N_1259,In_180,In_577);
and U1260 (N_1260,In_707,In_591);
or U1261 (N_1261,In_217,In_429);
or U1262 (N_1262,In_670,In_265);
or U1263 (N_1263,In_550,In_274);
nor U1264 (N_1264,In_6,In_284);
or U1265 (N_1265,In_162,In_505);
nand U1266 (N_1266,In_440,In_309);
or U1267 (N_1267,In_164,In_616);
nand U1268 (N_1268,In_228,In_143);
nand U1269 (N_1269,In_506,In_27);
nor U1270 (N_1270,In_251,In_369);
nor U1271 (N_1271,In_49,In_29);
xor U1272 (N_1272,In_58,In_84);
or U1273 (N_1273,In_116,In_493);
or U1274 (N_1274,In_130,In_147);
nor U1275 (N_1275,In_31,In_417);
or U1276 (N_1276,In_411,In_303);
nand U1277 (N_1277,In_219,In_309);
nor U1278 (N_1278,In_186,In_634);
and U1279 (N_1279,In_527,In_628);
or U1280 (N_1280,In_330,In_346);
nand U1281 (N_1281,In_367,In_745);
nor U1282 (N_1282,In_12,In_220);
nor U1283 (N_1283,In_403,In_733);
nand U1284 (N_1284,In_321,In_605);
or U1285 (N_1285,In_626,In_134);
or U1286 (N_1286,In_226,In_528);
or U1287 (N_1287,In_149,In_379);
and U1288 (N_1288,In_519,In_355);
and U1289 (N_1289,In_722,In_598);
or U1290 (N_1290,In_382,In_673);
and U1291 (N_1291,In_604,In_189);
nor U1292 (N_1292,In_41,In_585);
and U1293 (N_1293,In_502,In_173);
and U1294 (N_1294,In_562,In_516);
nand U1295 (N_1295,In_700,In_233);
nor U1296 (N_1296,In_311,In_717);
or U1297 (N_1297,In_301,In_592);
nor U1298 (N_1298,In_492,In_114);
and U1299 (N_1299,In_325,In_630);
nand U1300 (N_1300,In_439,In_154);
nand U1301 (N_1301,In_741,In_410);
and U1302 (N_1302,In_318,In_88);
and U1303 (N_1303,In_252,In_348);
or U1304 (N_1304,In_680,In_468);
nand U1305 (N_1305,In_433,In_613);
nor U1306 (N_1306,In_393,In_373);
nor U1307 (N_1307,In_700,In_338);
xor U1308 (N_1308,In_339,In_455);
and U1309 (N_1309,In_106,In_726);
nand U1310 (N_1310,In_468,In_279);
or U1311 (N_1311,In_19,In_164);
and U1312 (N_1312,In_569,In_154);
nand U1313 (N_1313,In_332,In_44);
and U1314 (N_1314,In_167,In_37);
nand U1315 (N_1315,In_623,In_295);
or U1316 (N_1316,In_474,In_482);
nand U1317 (N_1317,In_201,In_308);
or U1318 (N_1318,In_425,In_591);
nand U1319 (N_1319,In_516,In_696);
nor U1320 (N_1320,In_145,In_650);
and U1321 (N_1321,In_139,In_243);
or U1322 (N_1322,In_326,In_542);
or U1323 (N_1323,In_301,In_366);
nor U1324 (N_1324,In_115,In_607);
nand U1325 (N_1325,In_741,In_518);
nand U1326 (N_1326,In_256,In_287);
nand U1327 (N_1327,In_577,In_433);
nor U1328 (N_1328,In_369,In_680);
nand U1329 (N_1329,In_713,In_322);
nor U1330 (N_1330,In_146,In_722);
and U1331 (N_1331,In_291,In_436);
or U1332 (N_1332,In_304,In_746);
nand U1333 (N_1333,In_394,In_519);
nand U1334 (N_1334,In_407,In_98);
and U1335 (N_1335,In_246,In_136);
or U1336 (N_1336,In_627,In_298);
and U1337 (N_1337,In_344,In_139);
nand U1338 (N_1338,In_497,In_12);
nand U1339 (N_1339,In_343,In_323);
or U1340 (N_1340,In_336,In_642);
or U1341 (N_1341,In_498,In_361);
nor U1342 (N_1342,In_440,In_566);
and U1343 (N_1343,In_209,In_97);
or U1344 (N_1344,In_527,In_605);
nand U1345 (N_1345,In_615,In_460);
and U1346 (N_1346,In_314,In_544);
and U1347 (N_1347,In_149,In_307);
and U1348 (N_1348,In_701,In_176);
or U1349 (N_1349,In_646,In_120);
nor U1350 (N_1350,In_334,In_438);
or U1351 (N_1351,In_48,In_374);
nor U1352 (N_1352,In_516,In_645);
and U1353 (N_1353,In_428,In_128);
and U1354 (N_1354,In_590,In_51);
and U1355 (N_1355,In_32,In_91);
nand U1356 (N_1356,In_477,In_5);
and U1357 (N_1357,In_691,In_636);
nor U1358 (N_1358,In_160,In_732);
nand U1359 (N_1359,In_246,In_125);
and U1360 (N_1360,In_498,In_468);
xnor U1361 (N_1361,In_555,In_112);
and U1362 (N_1362,In_67,In_276);
or U1363 (N_1363,In_717,In_589);
nand U1364 (N_1364,In_139,In_155);
nor U1365 (N_1365,In_567,In_745);
nor U1366 (N_1366,In_281,In_19);
or U1367 (N_1367,In_378,In_374);
nor U1368 (N_1368,In_441,In_670);
or U1369 (N_1369,In_285,In_469);
and U1370 (N_1370,In_459,In_702);
and U1371 (N_1371,In_624,In_75);
nor U1372 (N_1372,In_675,In_186);
nand U1373 (N_1373,In_488,In_367);
xnor U1374 (N_1374,In_308,In_628);
nor U1375 (N_1375,In_13,In_415);
nand U1376 (N_1376,In_367,In_272);
and U1377 (N_1377,In_463,In_180);
nand U1378 (N_1378,In_620,In_512);
nor U1379 (N_1379,In_308,In_119);
nor U1380 (N_1380,In_54,In_49);
and U1381 (N_1381,In_61,In_461);
and U1382 (N_1382,In_672,In_498);
or U1383 (N_1383,In_630,In_223);
nand U1384 (N_1384,In_118,In_14);
or U1385 (N_1385,In_131,In_298);
or U1386 (N_1386,In_238,In_67);
nand U1387 (N_1387,In_145,In_621);
nand U1388 (N_1388,In_41,In_334);
nor U1389 (N_1389,In_74,In_352);
nor U1390 (N_1390,In_525,In_314);
and U1391 (N_1391,In_256,In_541);
or U1392 (N_1392,In_252,In_327);
xor U1393 (N_1393,In_718,In_625);
and U1394 (N_1394,In_72,In_218);
nand U1395 (N_1395,In_83,In_642);
or U1396 (N_1396,In_144,In_388);
and U1397 (N_1397,In_353,In_52);
nand U1398 (N_1398,In_90,In_138);
or U1399 (N_1399,In_175,In_366);
nor U1400 (N_1400,In_191,In_739);
or U1401 (N_1401,In_575,In_169);
and U1402 (N_1402,In_736,In_73);
or U1403 (N_1403,In_300,In_732);
nor U1404 (N_1404,In_352,In_480);
nand U1405 (N_1405,In_397,In_711);
or U1406 (N_1406,In_325,In_594);
nor U1407 (N_1407,In_411,In_415);
or U1408 (N_1408,In_458,In_88);
and U1409 (N_1409,In_151,In_277);
nor U1410 (N_1410,In_412,In_110);
nor U1411 (N_1411,In_599,In_342);
nor U1412 (N_1412,In_640,In_278);
nor U1413 (N_1413,In_79,In_199);
or U1414 (N_1414,In_729,In_410);
and U1415 (N_1415,In_428,In_535);
or U1416 (N_1416,In_446,In_723);
nand U1417 (N_1417,In_114,In_449);
nor U1418 (N_1418,In_496,In_740);
nor U1419 (N_1419,In_710,In_425);
and U1420 (N_1420,In_205,In_102);
or U1421 (N_1421,In_461,In_725);
or U1422 (N_1422,In_524,In_268);
and U1423 (N_1423,In_301,In_467);
nand U1424 (N_1424,In_208,In_647);
nor U1425 (N_1425,In_82,In_439);
or U1426 (N_1426,In_276,In_52);
nor U1427 (N_1427,In_682,In_579);
nor U1428 (N_1428,In_640,In_235);
and U1429 (N_1429,In_667,In_451);
and U1430 (N_1430,In_310,In_433);
and U1431 (N_1431,In_467,In_448);
nor U1432 (N_1432,In_305,In_121);
xnor U1433 (N_1433,In_670,In_315);
and U1434 (N_1434,In_706,In_309);
or U1435 (N_1435,In_341,In_281);
or U1436 (N_1436,In_500,In_305);
and U1437 (N_1437,In_456,In_312);
and U1438 (N_1438,In_265,In_319);
nand U1439 (N_1439,In_713,In_139);
or U1440 (N_1440,In_438,In_332);
and U1441 (N_1441,In_399,In_27);
nor U1442 (N_1442,In_651,In_338);
nor U1443 (N_1443,In_381,In_615);
or U1444 (N_1444,In_585,In_634);
or U1445 (N_1445,In_247,In_29);
nand U1446 (N_1446,In_395,In_612);
and U1447 (N_1447,In_31,In_723);
and U1448 (N_1448,In_607,In_648);
and U1449 (N_1449,In_535,In_568);
nand U1450 (N_1450,In_665,In_17);
nand U1451 (N_1451,In_498,In_658);
nor U1452 (N_1452,In_69,In_618);
nand U1453 (N_1453,In_144,In_598);
and U1454 (N_1454,In_531,In_636);
nand U1455 (N_1455,In_649,In_655);
or U1456 (N_1456,In_224,In_242);
xnor U1457 (N_1457,In_530,In_423);
xor U1458 (N_1458,In_526,In_191);
and U1459 (N_1459,In_712,In_672);
and U1460 (N_1460,In_76,In_145);
or U1461 (N_1461,In_692,In_283);
nor U1462 (N_1462,In_155,In_639);
nand U1463 (N_1463,In_209,In_189);
and U1464 (N_1464,In_155,In_554);
or U1465 (N_1465,In_746,In_331);
or U1466 (N_1466,In_334,In_505);
nor U1467 (N_1467,In_578,In_30);
nand U1468 (N_1468,In_670,In_438);
nand U1469 (N_1469,In_79,In_1);
nand U1470 (N_1470,In_221,In_462);
nand U1471 (N_1471,In_727,In_122);
nand U1472 (N_1472,In_388,In_14);
and U1473 (N_1473,In_661,In_234);
nor U1474 (N_1474,In_126,In_568);
and U1475 (N_1475,In_602,In_383);
nand U1476 (N_1476,In_411,In_229);
and U1477 (N_1477,In_154,In_87);
nor U1478 (N_1478,In_285,In_663);
nor U1479 (N_1479,In_525,In_522);
xor U1480 (N_1480,In_206,In_63);
or U1481 (N_1481,In_236,In_25);
nor U1482 (N_1482,In_355,In_55);
nand U1483 (N_1483,In_391,In_312);
or U1484 (N_1484,In_585,In_347);
or U1485 (N_1485,In_11,In_427);
or U1486 (N_1486,In_119,In_274);
or U1487 (N_1487,In_1,In_321);
or U1488 (N_1488,In_198,In_616);
or U1489 (N_1489,In_319,In_440);
or U1490 (N_1490,In_144,In_139);
and U1491 (N_1491,In_461,In_7);
or U1492 (N_1492,In_330,In_151);
and U1493 (N_1493,In_713,In_480);
nand U1494 (N_1494,In_709,In_706);
nor U1495 (N_1495,In_610,In_301);
and U1496 (N_1496,In_251,In_119);
or U1497 (N_1497,In_688,In_230);
and U1498 (N_1498,In_282,In_107);
nor U1499 (N_1499,In_518,In_83);
xnor U1500 (N_1500,In_331,In_559);
nor U1501 (N_1501,In_172,In_496);
and U1502 (N_1502,In_250,In_50);
nor U1503 (N_1503,In_565,In_437);
nor U1504 (N_1504,In_395,In_457);
nor U1505 (N_1505,In_676,In_29);
and U1506 (N_1506,In_645,In_447);
and U1507 (N_1507,In_589,In_248);
and U1508 (N_1508,In_323,In_161);
or U1509 (N_1509,In_59,In_327);
nor U1510 (N_1510,In_256,In_555);
or U1511 (N_1511,In_109,In_147);
and U1512 (N_1512,In_389,In_444);
nand U1513 (N_1513,In_493,In_167);
or U1514 (N_1514,In_232,In_482);
nor U1515 (N_1515,In_315,In_369);
or U1516 (N_1516,In_586,In_507);
nor U1517 (N_1517,In_339,In_328);
nor U1518 (N_1518,In_101,In_718);
nor U1519 (N_1519,In_495,In_414);
or U1520 (N_1520,In_201,In_317);
nand U1521 (N_1521,In_145,In_193);
nor U1522 (N_1522,In_187,In_381);
nor U1523 (N_1523,In_480,In_578);
or U1524 (N_1524,In_114,In_22);
nor U1525 (N_1525,In_418,In_353);
or U1526 (N_1526,In_204,In_657);
or U1527 (N_1527,In_514,In_651);
nor U1528 (N_1528,In_499,In_642);
or U1529 (N_1529,In_157,In_716);
or U1530 (N_1530,In_525,In_178);
or U1531 (N_1531,In_320,In_267);
or U1532 (N_1532,In_92,In_430);
nor U1533 (N_1533,In_596,In_144);
and U1534 (N_1534,In_167,In_708);
nor U1535 (N_1535,In_275,In_523);
nor U1536 (N_1536,In_285,In_498);
nor U1537 (N_1537,In_426,In_339);
xnor U1538 (N_1538,In_314,In_637);
and U1539 (N_1539,In_163,In_159);
and U1540 (N_1540,In_312,In_310);
or U1541 (N_1541,In_107,In_483);
nand U1542 (N_1542,In_157,In_289);
nand U1543 (N_1543,In_198,In_549);
nand U1544 (N_1544,In_163,In_613);
nand U1545 (N_1545,In_398,In_34);
or U1546 (N_1546,In_280,In_317);
or U1547 (N_1547,In_370,In_120);
nor U1548 (N_1548,In_589,In_582);
and U1549 (N_1549,In_91,In_242);
and U1550 (N_1550,In_626,In_479);
nand U1551 (N_1551,In_115,In_182);
nor U1552 (N_1552,In_566,In_350);
and U1553 (N_1553,In_411,In_274);
or U1554 (N_1554,In_217,In_553);
nand U1555 (N_1555,In_676,In_141);
and U1556 (N_1556,In_68,In_417);
nor U1557 (N_1557,In_392,In_308);
nand U1558 (N_1558,In_490,In_155);
nor U1559 (N_1559,In_112,In_594);
nor U1560 (N_1560,In_159,In_643);
nor U1561 (N_1561,In_453,In_574);
nor U1562 (N_1562,In_253,In_54);
nand U1563 (N_1563,In_200,In_332);
or U1564 (N_1564,In_577,In_29);
nand U1565 (N_1565,In_229,In_477);
and U1566 (N_1566,In_222,In_22);
xor U1567 (N_1567,In_81,In_401);
nand U1568 (N_1568,In_111,In_88);
or U1569 (N_1569,In_265,In_334);
nor U1570 (N_1570,In_37,In_676);
nor U1571 (N_1571,In_328,In_676);
nand U1572 (N_1572,In_37,In_593);
nor U1573 (N_1573,In_44,In_399);
or U1574 (N_1574,In_693,In_549);
nor U1575 (N_1575,In_257,In_531);
xnor U1576 (N_1576,In_309,In_642);
or U1577 (N_1577,In_452,In_535);
or U1578 (N_1578,In_441,In_420);
nor U1579 (N_1579,In_223,In_369);
or U1580 (N_1580,In_605,In_406);
nor U1581 (N_1581,In_144,In_680);
nor U1582 (N_1582,In_93,In_653);
nand U1583 (N_1583,In_561,In_692);
nor U1584 (N_1584,In_114,In_433);
or U1585 (N_1585,In_746,In_434);
and U1586 (N_1586,In_292,In_237);
or U1587 (N_1587,In_441,In_353);
nor U1588 (N_1588,In_482,In_14);
nand U1589 (N_1589,In_550,In_308);
or U1590 (N_1590,In_695,In_457);
or U1591 (N_1591,In_511,In_569);
nand U1592 (N_1592,In_102,In_262);
nor U1593 (N_1593,In_122,In_534);
nor U1594 (N_1594,In_27,In_521);
nand U1595 (N_1595,In_568,In_630);
or U1596 (N_1596,In_347,In_297);
nand U1597 (N_1597,In_136,In_350);
nand U1598 (N_1598,In_454,In_503);
or U1599 (N_1599,In_732,In_628);
and U1600 (N_1600,In_301,In_635);
nand U1601 (N_1601,In_723,In_589);
nand U1602 (N_1602,In_179,In_188);
nand U1603 (N_1603,In_671,In_279);
and U1604 (N_1604,In_721,In_0);
nand U1605 (N_1605,In_446,In_435);
and U1606 (N_1606,In_393,In_199);
nor U1607 (N_1607,In_712,In_5);
nand U1608 (N_1608,In_415,In_539);
nand U1609 (N_1609,In_288,In_60);
nand U1610 (N_1610,In_47,In_448);
nor U1611 (N_1611,In_321,In_30);
or U1612 (N_1612,In_702,In_482);
or U1613 (N_1613,In_103,In_182);
nand U1614 (N_1614,In_46,In_341);
and U1615 (N_1615,In_724,In_580);
nand U1616 (N_1616,In_404,In_661);
nor U1617 (N_1617,In_246,In_586);
or U1618 (N_1618,In_313,In_23);
nor U1619 (N_1619,In_706,In_240);
nand U1620 (N_1620,In_487,In_235);
nand U1621 (N_1621,In_28,In_593);
and U1622 (N_1622,In_109,In_522);
nor U1623 (N_1623,In_116,In_654);
xor U1624 (N_1624,In_131,In_360);
or U1625 (N_1625,In_673,In_359);
nand U1626 (N_1626,In_451,In_643);
nand U1627 (N_1627,In_505,In_416);
nand U1628 (N_1628,In_417,In_513);
nand U1629 (N_1629,In_575,In_425);
or U1630 (N_1630,In_738,In_692);
or U1631 (N_1631,In_397,In_650);
nor U1632 (N_1632,In_533,In_37);
and U1633 (N_1633,In_740,In_409);
and U1634 (N_1634,In_81,In_569);
nand U1635 (N_1635,In_501,In_302);
and U1636 (N_1636,In_680,In_460);
nand U1637 (N_1637,In_344,In_157);
nor U1638 (N_1638,In_364,In_447);
or U1639 (N_1639,In_37,In_519);
or U1640 (N_1640,In_76,In_16);
nor U1641 (N_1641,In_4,In_92);
nor U1642 (N_1642,In_101,In_223);
nand U1643 (N_1643,In_598,In_389);
nand U1644 (N_1644,In_658,In_564);
nor U1645 (N_1645,In_426,In_200);
nor U1646 (N_1646,In_344,In_167);
and U1647 (N_1647,In_626,In_436);
nand U1648 (N_1648,In_527,In_501);
xnor U1649 (N_1649,In_646,In_447);
nand U1650 (N_1650,In_309,In_356);
xor U1651 (N_1651,In_534,In_202);
nor U1652 (N_1652,In_71,In_117);
and U1653 (N_1653,In_652,In_696);
nor U1654 (N_1654,In_285,In_60);
or U1655 (N_1655,In_393,In_68);
or U1656 (N_1656,In_731,In_529);
nor U1657 (N_1657,In_390,In_99);
nor U1658 (N_1658,In_525,In_453);
nor U1659 (N_1659,In_209,In_398);
or U1660 (N_1660,In_70,In_398);
and U1661 (N_1661,In_237,In_393);
nand U1662 (N_1662,In_153,In_402);
and U1663 (N_1663,In_176,In_88);
or U1664 (N_1664,In_564,In_300);
nor U1665 (N_1665,In_729,In_186);
nor U1666 (N_1666,In_317,In_307);
nor U1667 (N_1667,In_12,In_706);
nor U1668 (N_1668,In_19,In_286);
nand U1669 (N_1669,In_226,In_135);
xor U1670 (N_1670,In_635,In_633);
nand U1671 (N_1671,In_401,In_584);
nor U1672 (N_1672,In_154,In_521);
nand U1673 (N_1673,In_584,In_93);
nor U1674 (N_1674,In_206,In_202);
nor U1675 (N_1675,In_347,In_107);
nand U1676 (N_1676,In_472,In_12);
nand U1677 (N_1677,In_318,In_595);
and U1678 (N_1678,In_549,In_485);
and U1679 (N_1679,In_359,In_283);
nor U1680 (N_1680,In_95,In_102);
nor U1681 (N_1681,In_660,In_323);
xnor U1682 (N_1682,In_117,In_458);
nor U1683 (N_1683,In_154,In_73);
nor U1684 (N_1684,In_592,In_635);
or U1685 (N_1685,In_264,In_193);
nand U1686 (N_1686,In_315,In_148);
and U1687 (N_1687,In_50,In_218);
nand U1688 (N_1688,In_140,In_365);
and U1689 (N_1689,In_650,In_12);
nor U1690 (N_1690,In_205,In_343);
nand U1691 (N_1691,In_41,In_382);
nor U1692 (N_1692,In_736,In_1);
or U1693 (N_1693,In_620,In_131);
nand U1694 (N_1694,In_83,In_304);
and U1695 (N_1695,In_398,In_54);
and U1696 (N_1696,In_422,In_506);
and U1697 (N_1697,In_407,In_632);
or U1698 (N_1698,In_425,In_725);
nand U1699 (N_1699,In_149,In_582);
and U1700 (N_1700,In_696,In_234);
or U1701 (N_1701,In_496,In_635);
nor U1702 (N_1702,In_479,In_272);
or U1703 (N_1703,In_71,In_574);
nor U1704 (N_1704,In_161,In_651);
nor U1705 (N_1705,In_637,In_192);
and U1706 (N_1706,In_405,In_636);
or U1707 (N_1707,In_150,In_645);
nand U1708 (N_1708,In_694,In_724);
or U1709 (N_1709,In_510,In_140);
nor U1710 (N_1710,In_413,In_162);
nor U1711 (N_1711,In_9,In_472);
and U1712 (N_1712,In_111,In_617);
nand U1713 (N_1713,In_141,In_599);
or U1714 (N_1714,In_96,In_631);
and U1715 (N_1715,In_57,In_602);
or U1716 (N_1716,In_516,In_573);
nor U1717 (N_1717,In_375,In_152);
nand U1718 (N_1718,In_465,In_286);
nor U1719 (N_1719,In_452,In_274);
nand U1720 (N_1720,In_295,In_212);
or U1721 (N_1721,In_584,In_748);
xnor U1722 (N_1722,In_737,In_167);
nand U1723 (N_1723,In_594,In_190);
and U1724 (N_1724,In_152,In_724);
or U1725 (N_1725,In_265,In_631);
nand U1726 (N_1726,In_438,In_589);
nor U1727 (N_1727,In_458,In_41);
and U1728 (N_1728,In_741,In_342);
and U1729 (N_1729,In_551,In_623);
and U1730 (N_1730,In_708,In_532);
nand U1731 (N_1731,In_339,In_402);
and U1732 (N_1732,In_488,In_534);
and U1733 (N_1733,In_452,In_217);
or U1734 (N_1734,In_49,In_224);
and U1735 (N_1735,In_439,In_84);
nor U1736 (N_1736,In_238,In_429);
or U1737 (N_1737,In_270,In_201);
or U1738 (N_1738,In_696,In_328);
xor U1739 (N_1739,In_348,In_620);
nor U1740 (N_1740,In_455,In_157);
or U1741 (N_1741,In_229,In_306);
nand U1742 (N_1742,In_719,In_728);
or U1743 (N_1743,In_81,In_504);
nand U1744 (N_1744,In_571,In_735);
nor U1745 (N_1745,In_291,In_280);
and U1746 (N_1746,In_63,In_717);
and U1747 (N_1747,In_275,In_317);
or U1748 (N_1748,In_173,In_612);
nor U1749 (N_1749,In_65,In_474);
nor U1750 (N_1750,In_156,In_669);
nand U1751 (N_1751,In_276,In_521);
and U1752 (N_1752,In_705,In_527);
and U1753 (N_1753,In_171,In_456);
nor U1754 (N_1754,In_466,In_616);
or U1755 (N_1755,In_569,In_444);
and U1756 (N_1756,In_359,In_635);
nor U1757 (N_1757,In_563,In_629);
and U1758 (N_1758,In_211,In_475);
and U1759 (N_1759,In_259,In_561);
nor U1760 (N_1760,In_167,In_392);
and U1761 (N_1761,In_395,In_632);
and U1762 (N_1762,In_655,In_292);
nand U1763 (N_1763,In_218,In_443);
or U1764 (N_1764,In_609,In_400);
or U1765 (N_1765,In_212,In_642);
nand U1766 (N_1766,In_507,In_502);
nand U1767 (N_1767,In_357,In_214);
or U1768 (N_1768,In_14,In_379);
nand U1769 (N_1769,In_154,In_483);
or U1770 (N_1770,In_457,In_400);
nand U1771 (N_1771,In_112,In_279);
or U1772 (N_1772,In_128,In_723);
and U1773 (N_1773,In_553,In_485);
nand U1774 (N_1774,In_353,In_289);
and U1775 (N_1775,In_223,In_196);
or U1776 (N_1776,In_587,In_572);
nand U1777 (N_1777,In_60,In_360);
nand U1778 (N_1778,In_67,In_38);
nor U1779 (N_1779,In_733,In_332);
nand U1780 (N_1780,In_241,In_613);
or U1781 (N_1781,In_463,In_664);
nand U1782 (N_1782,In_150,In_492);
and U1783 (N_1783,In_618,In_451);
or U1784 (N_1784,In_703,In_683);
nor U1785 (N_1785,In_473,In_723);
and U1786 (N_1786,In_355,In_82);
nor U1787 (N_1787,In_708,In_387);
nand U1788 (N_1788,In_603,In_631);
nor U1789 (N_1789,In_94,In_697);
nand U1790 (N_1790,In_679,In_732);
and U1791 (N_1791,In_195,In_141);
or U1792 (N_1792,In_134,In_170);
nor U1793 (N_1793,In_39,In_205);
or U1794 (N_1794,In_120,In_724);
nand U1795 (N_1795,In_532,In_617);
nor U1796 (N_1796,In_156,In_17);
or U1797 (N_1797,In_11,In_104);
nor U1798 (N_1798,In_99,In_213);
and U1799 (N_1799,In_525,In_697);
and U1800 (N_1800,In_600,In_328);
nor U1801 (N_1801,In_402,In_593);
and U1802 (N_1802,In_369,In_583);
nand U1803 (N_1803,In_235,In_698);
nor U1804 (N_1804,In_613,In_715);
nor U1805 (N_1805,In_252,In_701);
or U1806 (N_1806,In_107,In_27);
nand U1807 (N_1807,In_445,In_142);
nor U1808 (N_1808,In_239,In_276);
and U1809 (N_1809,In_245,In_235);
or U1810 (N_1810,In_539,In_154);
nor U1811 (N_1811,In_521,In_732);
and U1812 (N_1812,In_588,In_56);
nand U1813 (N_1813,In_703,In_650);
nand U1814 (N_1814,In_74,In_556);
and U1815 (N_1815,In_103,In_11);
and U1816 (N_1816,In_588,In_727);
nor U1817 (N_1817,In_219,In_428);
nor U1818 (N_1818,In_701,In_512);
and U1819 (N_1819,In_581,In_56);
or U1820 (N_1820,In_90,In_27);
or U1821 (N_1821,In_42,In_256);
nand U1822 (N_1822,In_354,In_161);
nand U1823 (N_1823,In_412,In_459);
nor U1824 (N_1824,In_627,In_380);
and U1825 (N_1825,In_602,In_40);
and U1826 (N_1826,In_180,In_353);
nand U1827 (N_1827,In_424,In_706);
and U1828 (N_1828,In_543,In_104);
nor U1829 (N_1829,In_705,In_571);
and U1830 (N_1830,In_129,In_622);
or U1831 (N_1831,In_718,In_75);
and U1832 (N_1832,In_110,In_728);
or U1833 (N_1833,In_591,In_299);
nand U1834 (N_1834,In_196,In_147);
nor U1835 (N_1835,In_255,In_292);
nand U1836 (N_1836,In_632,In_76);
nor U1837 (N_1837,In_50,In_506);
and U1838 (N_1838,In_532,In_261);
or U1839 (N_1839,In_429,In_480);
or U1840 (N_1840,In_110,In_271);
nor U1841 (N_1841,In_332,In_114);
nand U1842 (N_1842,In_485,In_571);
and U1843 (N_1843,In_412,In_503);
or U1844 (N_1844,In_41,In_743);
nor U1845 (N_1845,In_429,In_99);
nand U1846 (N_1846,In_299,In_45);
and U1847 (N_1847,In_20,In_654);
and U1848 (N_1848,In_722,In_515);
or U1849 (N_1849,In_356,In_438);
and U1850 (N_1850,In_268,In_618);
nand U1851 (N_1851,In_530,In_115);
and U1852 (N_1852,In_743,In_175);
or U1853 (N_1853,In_517,In_103);
nand U1854 (N_1854,In_203,In_175);
and U1855 (N_1855,In_516,In_669);
or U1856 (N_1856,In_426,In_694);
or U1857 (N_1857,In_438,In_398);
and U1858 (N_1858,In_572,In_561);
or U1859 (N_1859,In_41,In_194);
or U1860 (N_1860,In_178,In_179);
nand U1861 (N_1861,In_302,In_323);
nand U1862 (N_1862,In_244,In_26);
nor U1863 (N_1863,In_700,In_46);
or U1864 (N_1864,In_603,In_595);
nand U1865 (N_1865,In_519,In_646);
nor U1866 (N_1866,In_733,In_334);
xor U1867 (N_1867,In_172,In_544);
xor U1868 (N_1868,In_250,In_528);
and U1869 (N_1869,In_603,In_591);
nor U1870 (N_1870,In_749,In_744);
nand U1871 (N_1871,In_524,In_22);
and U1872 (N_1872,In_282,In_509);
or U1873 (N_1873,In_145,In_388);
and U1874 (N_1874,In_304,In_636);
nand U1875 (N_1875,In_703,In_572);
nor U1876 (N_1876,In_389,In_601);
xor U1877 (N_1877,In_419,In_588);
or U1878 (N_1878,In_96,In_692);
or U1879 (N_1879,In_133,In_4);
or U1880 (N_1880,In_607,In_394);
and U1881 (N_1881,In_134,In_585);
and U1882 (N_1882,In_525,In_578);
and U1883 (N_1883,In_746,In_33);
and U1884 (N_1884,In_193,In_94);
xor U1885 (N_1885,In_318,In_407);
or U1886 (N_1886,In_332,In_336);
nor U1887 (N_1887,In_588,In_437);
or U1888 (N_1888,In_513,In_140);
or U1889 (N_1889,In_730,In_231);
nand U1890 (N_1890,In_66,In_588);
nand U1891 (N_1891,In_550,In_516);
nand U1892 (N_1892,In_714,In_483);
and U1893 (N_1893,In_633,In_441);
or U1894 (N_1894,In_627,In_238);
or U1895 (N_1895,In_270,In_126);
or U1896 (N_1896,In_247,In_617);
or U1897 (N_1897,In_54,In_81);
and U1898 (N_1898,In_344,In_722);
and U1899 (N_1899,In_170,In_537);
or U1900 (N_1900,In_691,In_745);
and U1901 (N_1901,In_589,In_220);
or U1902 (N_1902,In_521,In_92);
nor U1903 (N_1903,In_425,In_7);
nor U1904 (N_1904,In_259,In_89);
or U1905 (N_1905,In_668,In_488);
or U1906 (N_1906,In_612,In_438);
nand U1907 (N_1907,In_127,In_66);
nor U1908 (N_1908,In_748,In_463);
xor U1909 (N_1909,In_605,In_734);
nand U1910 (N_1910,In_418,In_309);
nand U1911 (N_1911,In_675,In_297);
and U1912 (N_1912,In_696,In_368);
and U1913 (N_1913,In_590,In_745);
or U1914 (N_1914,In_268,In_83);
and U1915 (N_1915,In_212,In_31);
or U1916 (N_1916,In_358,In_16);
nand U1917 (N_1917,In_700,In_687);
nor U1918 (N_1918,In_102,In_717);
nand U1919 (N_1919,In_567,In_113);
or U1920 (N_1920,In_441,In_392);
or U1921 (N_1921,In_584,In_741);
nor U1922 (N_1922,In_433,In_645);
or U1923 (N_1923,In_486,In_564);
and U1924 (N_1924,In_580,In_47);
or U1925 (N_1925,In_452,In_336);
nor U1926 (N_1926,In_72,In_556);
or U1927 (N_1927,In_28,In_349);
nand U1928 (N_1928,In_189,In_673);
and U1929 (N_1929,In_104,In_640);
nor U1930 (N_1930,In_449,In_105);
nand U1931 (N_1931,In_480,In_111);
xor U1932 (N_1932,In_495,In_275);
nor U1933 (N_1933,In_349,In_595);
nand U1934 (N_1934,In_282,In_577);
xnor U1935 (N_1935,In_506,In_686);
nand U1936 (N_1936,In_64,In_255);
or U1937 (N_1937,In_488,In_2);
and U1938 (N_1938,In_154,In_41);
or U1939 (N_1939,In_592,In_233);
nand U1940 (N_1940,In_25,In_639);
and U1941 (N_1941,In_726,In_44);
and U1942 (N_1942,In_426,In_190);
nor U1943 (N_1943,In_364,In_669);
nor U1944 (N_1944,In_145,In_19);
or U1945 (N_1945,In_180,In_412);
or U1946 (N_1946,In_416,In_617);
nand U1947 (N_1947,In_415,In_243);
nor U1948 (N_1948,In_51,In_339);
nand U1949 (N_1949,In_418,In_110);
nand U1950 (N_1950,In_536,In_4);
nand U1951 (N_1951,In_159,In_219);
nor U1952 (N_1952,In_245,In_443);
and U1953 (N_1953,In_66,In_31);
nand U1954 (N_1954,In_155,In_366);
and U1955 (N_1955,In_734,In_439);
or U1956 (N_1956,In_567,In_164);
and U1957 (N_1957,In_604,In_346);
nor U1958 (N_1958,In_138,In_489);
nand U1959 (N_1959,In_415,In_94);
and U1960 (N_1960,In_622,In_520);
nand U1961 (N_1961,In_345,In_726);
or U1962 (N_1962,In_77,In_447);
and U1963 (N_1963,In_298,In_422);
nor U1964 (N_1964,In_322,In_238);
and U1965 (N_1965,In_747,In_564);
xnor U1966 (N_1966,In_135,In_514);
xnor U1967 (N_1967,In_745,In_747);
or U1968 (N_1968,In_684,In_706);
or U1969 (N_1969,In_656,In_353);
nand U1970 (N_1970,In_599,In_70);
and U1971 (N_1971,In_515,In_654);
nand U1972 (N_1972,In_631,In_26);
xnor U1973 (N_1973,In_381,In_420);
or U1974 (N_1974,In_160,In_348);
nand U1975 (N_1975,In_265,In_82);
nor U1976 (N_1976,In_199,In_504);
or U1977 (N_1977,In_519,In_232);
and U1978 (N_1978,In_607,In_59);
or U1979 (N_1979,In_76,In_0);
nand U1980 (N_1980,In_625,In_137);
nand U1981 (N_1981,In_122,In_208);
nand U1982 (N_1982,In_422,In_203);
xor U1983 (N_1983,In_475,In_89);
or U1984 (N_1984,In_209,In_355);
nand U1985 (N_1985,In_165,In_141);
nand U1986 (N_1986,In_131,In_482);
and U1987 (N_1987,In_165,In_745);
nor U1988 (N_1988,In_401,In_588);
nand U1989 (N_1989,In_18,In_360);
and U1990 (N_1990,In_232,In_159);
nand U1991 (N_1991,In_10,In_712);
or U1992 (N_1992,In_703,In_489);
nand U1993 (N_1993,In_61,In_446);
or U1994 (N_1994,In_438,In_474);
and U1995 (N_1995,In_53,In_420);
nor U1996 (N_1996,In_290,In_361);
or U1997 (N_1997,In_154,In_114);
or U1998 (N_1998,In_97,In_217);
or U1999 (N_1999,In_214,In_175);
nand U2000 (N_2000,In_91,In_348);
or U2001 (N_2001,In_596,In_505);
nand U2002 (N_2002,In_90,In_697);
nand U2003 (N_2003,In_159,In_181);
and U2004 (N_2004,In_200,In_514);
or U2005 (N_2005,In_717,In_205);
or U2006 (N_2006,In_505,In_1);
nand U2007 (N_2007,In_227,In_163);
or U2008 (N_2008,In_349,In_61);
nor U2009 (N_2009,In_239,In_324);
or U2010 (N_2010,In_681,In_648);
nand U2011 (N_2011,In_447,In_91);
or U2012 (N_2012,In_441,In_728);
and U2013 (N_2013,In_472,In_463);
nor U2014 (N_2014,In_680,In_492);
or U2015 (N_2015,In_83,In_744);
and U2016 (N_2016,In_598,In_244);
and U2017 (N_2017,In_606,In_163);
nand U2018 (N_2018,In_378,In_218);
and U2019 (N_2019,In_588,In_291);
nor U2020 (N_2020,In_122,In_247);
and U2021 (N_2021,In_388,In_22);
or U2022 (N_2022,In_66,In_412);
nor U2023 (N_2023,In_77,In_416);
nor U2024 (N_2024,In_452,In_292);
and U2025 (N_2025,In_330,In_731);
xnor U2026 (N_2026,In_394,In_473);
and U2027 (N_2027,In_540,In_745);
or U2028 (N_2028,In_432,In_288);
and U2029 (N_2029,In_593,In_531);
and U2030 (N_2030,In_517,In_549);
nor U2031 (N_2031,In_568,In_84);
and U2032 (N_2032,In_576,In_439);
and U2033 (N_2033,In_582,In_98);
or U2034 (N_2034,In_622,In_183);
xor U2035 (N_2035,In_646,In_177);
nand U2036 (N_2036,In_714,In_171);
and U2037 (N_2037,In_644,In_735);
nor U2038 (N_2038,In_226,In_178);
nor U2039 (N_2039,In_702,In_102);
and U2040 (N_2040,In_303,In_725);
or U2041 (N_2041,In_683,In_431);
xor U2042 (N_2042,In_486,In_477);
nand U2043 (N_2043,In_264,In_277);
or U2044 (N_2044,In_742,In_407);
nand U2045 (N_2045,In_125,In_36);
nand U2046 (N_2046,In_219,In_356);
nand U2047 (N_2047,In_239,In_340);
or U2048 (N_2048,In_399,In_601);
nand U2049 (N_2049,In_201,In_723);
nor U2050 (N_2050,In_519,In_185);
and U2051 (N_2051,In_698,In_608);
and U2052 (N_2052,In_7,In_228);
nor U2053 (N_2053,In_680,In_129);
and U2054 (N_2054,In_206,In_700);
and U2055 (N_2055,In_678,In_481);
nor U2056 (N_2056,In_438,In_429);
nand U2057 (N_2057,In_429,In_698);
nor U2058 (N_2058,In_670,In_184);
nand U2059 (N_2059,In_234,In_736);
nand U2060 (N_2060,In_257,In_488);
xor U2061 (N_2061,In_619,In_44);
nor U2062 (N_2062,In_482,In_145);
and U2063 (N_2063,In_69,In_422);
nor U2064 (N_2064,In_315,In_637);
nand U2065 (N_2065,In_553,In_727);
or U2066 (N_2066,In_13,In_625);
or U2067 (N_2067,In_95,In_516);
and U2068 (N_2068,In_253,In_351);
or U2069 (N_2069,In_442,In_602);
nor U2070 (N_2070,In_20,In_139);
or U2071 (N_2071,In_97,In_568);
and U2072 (N_2072,In_319,In_270);
and U2073 (N_2073,In_106,In_164);
nand U2074 (N_2074,In_97,In_143);
xor U2075 (N_2075,In_167,In_27);
nand U2076 (N_2076,In_125,In_181);
and U2077 (N_2077,In_415,In_599);
nand U2078 (N_2078,In_223,In_668);
nand U2079 (N_2079,In_159,In_389);
or U2080 (N_2080,In_74,In_197);
and U2081 (N_2081,In_10,In_168);
nand U2082 (N_2082,In_613,In_529);
nand U2083 (N_2083,In_265,In_129);
and U2084 (N_2084,In_578,In_38);
and U2085 (N_2085,In_509,In_416);
and U2086 (N_2086,In_621,In_450);
or U2087 (N_2087,In_231,In_527);
nor U2088 (N_2088,In_498,In_692);
and U2089 (N_2089,In_340,In_684);
or U2090 (N_2090,In_498,In_130);
nand U2091 (N_2091,In_595,In_634);
and U2092 (N_2092,In_174,In_240);
and U2093 (N_2093,In_281,In_687);
and U2094 (N_2094,In_205,In_96);
or U2095 (N_2095,In_418,In_260);
nor U2096 (N_2096,In_73,In_157);
nand U2097 (N_2097,In_717,In_321);
nor U2098 (N_2098,In_91,In_143);
nand U2099 (N_2099,In_231,In_426);
nand U2100 (N_2100,In_626,In_293);
xor U2101 (N_2101,In_225,In_330);
or U2102 (N_2102,In_659,In_492);
and U2103 (N_2103,In_734,In_491);
nor U2104 (N_2104,In_8,In_402);
nor U2105 (N_2105,In_654,In_578);
or U2106 (N_2106,In_630,In_344);
and U2107 (N_2107,In_224,In_584);
and U2108 (N_2108,In_190,In_353);
xor U2109 (N_2109,In_582,In_597);
nor U2110 (N_2110,In_301,In_685);
and U2111 (N_2111,In_731,In_498);
or U2112 (N_2112,In_226,In_287);
xnor U2113 (N_2113,In_238,In_66);
or U2114 (N_2114,In_578,In_566);
nand U2115 (N_2115,In_338,In_693);
nor U2116 (N_2116,In_135,In_109);
nor U2117 (N_2117,In_471,In_338);
or U2118 (N_2118,In_602,In_619);
nor U2119 (N_2119,In_366,In_375);
nand U2120 (N_2120,In_680,In_90);
or U2121 (N_2121,In_470,In_735);
nor U2122 (N_2122,In_159,In_44);
nor U2123 (N_2123,In_270,In_170);
and U2124 (N_2124,In_589,In_397);
nand U2125 (N_2125,In_409,In_143);
nand U2126 (N_2126,In_232,In_246);
and U2127 (N_2127,In_677,In_48);
and U2128 (N_2128,In_738,In_342);
nor U2129 (N_2129,In_167,In_232);
nand U2130 (N_2130,In_526,In_210);
nand U2131 (N_2131,In_433,In_421);
or U2132 (N_2132,In_254,In_113);
or U2133 (N_2133,In_498,In_320);
nand U2134 (N_2134,In_393,In_257);
nand U2135 (N_2135,In_445,In_1);
and U2136 (N_2136,In_222,In_150);
and U2137 (N_2137,In_537,In_287);
nor U2138 (N_2138,In_409,In_311);
nor U2139 (N_2139,In_207,In_667);
or U2140 (N_2140,In_106,In_653);
or U2141 (N_2141,In_387,In_342);
and U2142 (N_2142,In_524,In_680);
or U2143 (N_2143,In_124,In_432);
or U2144 (N_2144,In_303,In_669);
nand U2145 (N_2145,In_350,In_665);
or U2146 (N_2146,In_669,In_204);
xnor U2147 (N_2147,In_469,In_611);
nand U2148 (N_2148,In_283,In_43);
nor U2149 (N_2149,In_704,In_326);
nand U2150 (N_2150,In_407,In_122);
nand U2151 (N_2151,In_86,In_481);
and U2152 (N_2152,In_526,In_430);
nand U2153 (N_2153,In_747,In_552);
or U2154 (N_2154,In_721,In_520);
nand U2155 (N_2155,In_144,In_76);
nand U2156 (N_2156,In_613,In_146);
xnor U2157 (N_2157,In_0,In_662);
nor U2158 (N_2158,In_648,In_576);
nor U2159 (N_2159,In_608,In_100);
nand U2160 (N_2160,In_41,In_435);
nor U2161 (N_2161,In_732,In_509);
and U2162 (N_2162,In_49,In_724);
or U2163 (N_2163,In_87,In_305);
xor U2164 (N_2164,In_694,In_654);
or U2165 (N_2165,In_600,In_698);
nand U2166 (N_2166,In_690,In_125);
nor U2167 (N_2167,In_467,In_359);
and U2168 (N_2168,In_297,In_133);
nor U2169 (N_2169,In_427,In_67);
or U2170 (N_2170,In_554,In_217);
and U2171 (N_2171,In_100,In_475);
nand U2172 (N_2172,In_324,In_556);
and U2173 (N_2173,In_121,In_378);
nand U2174 (N_2174,In_653,In_319);
nand U2175 (N_2175,In_350,In_87);
or U2176 (N_2176,In_188,In_92);
nor U2177 (N_2177,In_352,In_178);
nor U2178 (N_2178,In_655,In_564);
nand U2179 (N_2179,In_667,In_416);
and U2180 (N_2180,In_179,In_634);
and U2181 (N_2181,In_222,In_7);
or U2182 (N_2182,In_362,In_675);
nor U2183 (N_2183,In_212,In_728);
or U2184 (N_2184,In_27,In_568);
nor U2185 (N_2185,In_475,In_151);
nor U2186 (N_2186,In_421,In_15);
or U2187 (N_2187,In_100,In_209);
nor U2188 (N_2188,In_483,In_21);
nand U2189 (N_2189,In_604,In_313);
or U2190 (N_2190,In_301,In_34);
and U2191 (N_2191,In_351,In_454);
nand U2192 (N_2192,In_408,In_580);
and U2193 (N_2193,In_14,In_381);
nand U2194 (N_2194,In_389,In_671);
nor U2195 (N_2195,In_699,In_206);
or U2196 (N_2196,In_402,In_277);
and U2197 (N_2197,In_524,In_276);
nand U2198 (N_2198,In_256,In_4);
and U2199 (N_2199,In_737,In_565);
nor U2200 (N_2200,In_586,In_270);
or U2201 (N_2201,In_80,In_308);
and U2202 (N_2202,In_611,In_625);
or U2203 (N_2203,In_151,In_143);
nor U2204 (N_2204,In_166,In_62);
nor U2205 (N_2205,In_266,In_638);
or U2206 (N_2206,In_65,In_585);
and U2207 (N_2207,In_24,In_340);
and U2208 (N_2208,In_452,In_15);
nor U2209 (N_2209,In_558,In_621);
and U2210 (N_2210,In_470,In_221);
nor U2211 (N_2211,In_245,In_5);
nand U2212 (N_2212,In_29,In_646);
or U2213 (N_2213,In_146,In_44);
nand U2214 (N_2214,In_173,In_178);
and U2215 (N_2215,In_320,In_671);
or U2216 (N_2216,In_395,In_447);
nor U2217 (N_2217,In_456,In_217);
or U2218 (N_2218,In_190,In_595);
nor U2219 (N_2219,In_717,In_386);
nor U2220 (N_2220,In_410,In_19);
or U2221 (N_2221,In_211,In_511);
nor U2222 (N_2222,In_530,In_193);
or U2223 (N_2223,In_212,In_64);
or U2224 (N_2224,In_153,In_519);
nand U2225 (N_2225,In_193,In_703);
or U2226 (N_2226,In_75,In_2);
nor U2227 (N_2227,In_670,In_617);
nand U2228 (N_2228,In_207,In_257);
nand U2229 (N_2229,In_573,In_354);
and U2230 (N_2230,In_121,In_472);
nor U2231 (N_2231,In_614,In_103);
or U2232 (N_2232,In_518,In_544);
and U2233 (N_2233,In_571,In_681);
and U2234 (N_2234,In_371,In_510);
nor U2235 (N_2235,In_383,In_59);
or U2236 (N_2236,In_323,In_342);
and U2237 (N_2237,In_360,In_394);
and U2238 (N_2238,In_710,In_244);
nor U2239 (N_2239,In_164,In_456);
or U2240 (N_2240,In_417,In_718);
nand U2241 (N_2241,In_334,In_728);
and U2242 (N_2242,In_594,In_577);
nor U2243 (N_2243,In_551,In_665);
nand U2244 (N_2244,In_544,In_349);
or U2245 (N_2245,In_170,In_254);
nor U2246 (N_2246,In_144,In_687);
or U2247 (N_2247,In_703,In_254);
and U2248 (N_2248,In_43,In_729);
or U2249 (N_2249,In_696,In_140);
nand U2250 (N_2250,In_337,In_357);
and U2251 (N_2251,In_578,In_250);
and U2252 (N_2252,In_482,In_419);
and U2253 (N_2253,In_290,In_736);
or U2254 (N_2254,In_544,In_725);
or U2255 (N_2255,In_248,In_302);
and U2256 (N_2256,In_124,In_400);
and U2257 (N_2257,In_116,In_738);
nor U2258 (N_2258,In_8,In_686);
and U2259 (N_2259,In_245,In_431);
nor U2260 (N_2260,In_185,In_727);
nor U2261 (N_2261,In_168,In_395);
and U2262 (N_2262,In_376,In_160);
nor U2263 (N_2263,In_482,In_276);
and U2264 (N_2264,In_371,In_705);
nand U2265 (N_2265,In_294,In_41);
and U2266 (N_2266,In_489,In_588);
xnor U2267 (N_2267,In_698,In_428);
nor U2268 (N_2268,In_239,In_106);
and U2269 (N_2269,In_563,In_83);
nand U2270 (N_2270,In_618,In_643);
and U2271 (N_2271,In_131,In_592);
nor U2272 (N_2272,In_51,In_472);
xnor U2273 (N_2273,In_250,In_620);
nor U2274 (N_2274,In_423,In_306);
and U2275 (N_2275,In_588,In_516);
nor U2276 (N_2276,In_231,In_8);
and U2277 (N_2277,In_185,In_413);
nor U2278 (N_2278,In_717,In_190);
or U2279 (N_2279,In_262,In_125);
nand U2280 (N_2280,In_0,In_171);
or U2281 (N_2281,In_302,In_321);
nand U2282 (N_2282,In_575,In_125);
nand U2283 (N_2283,In_246,In_264);
or U2284 (N_2284,In_229,In_412);
nor U2285 (N_2285,In_553,In_308);
nand U2286 (N_2286,In_662,In_174);
and U2287 (N_2287,In_106,In_147);
or U2288 (N_2288,In_686,In_340);
and U2289 (N_2289,In_114,In_264);
xor U2290 (N_2290,In_534,In_402);
nand U2291 (N_2291,In_707,In_133);
and U2292 (N_2292,In_21,In_555);
and U2293 (N_2293,In_611,In_53);
or U2294 (N_2294,In_520,In_147);
nand U2295 (N_2295,In_259,In_738);
nor U2296 (N_2296,In_365,In_223);
nor U2297 (N_2297,In_676,In_43);
xnor U2298 (N_2298,In_735,In_311);
nor U2299 (N_2299,In_357,In_649);
nor U2300 (N_2300,In_721,In_668);
nand U2301 (N_2301,In_430,In_523);
nor U2302 (N_2302,In_402,In_276);
or U2303 (N_2303,In_128,In_611);
nor U2304 (N_2304,In_625,In_554);
nand U2305 (N_2305,In_16,In_305);
nand U2306 (N_2306,In_50,In_547);
nand U2307 (N_2307,In_564,In_505);
and U2308 (N_2308,In_95,In_363);
and U2309 (N_2309,In_257,In_506);
and U2310 (N_2310,In_295,In_79);
and U2311 (N_2311,In_554,In_159);
and U2312 (N_2312,In_480,In_7);
nor U2313 (N_2313,In_569,In_281);
nand U2314 (N_2314,In_663,In_570);
and U2315 (N_2315,In_289,In_438);
and U2316 (N_2316,In_708,In_524);
nor U2317 (N_2317,In_564,In_86);
or U2318 (N_2318,In_647,In_535);
and U2319 (N_2319,In_303,In_20);
nand U2320 (N_2320,In_357,In_264);
xnor U2321 (N_2321,In_36,In_516);
or U2322 (N_2322,In_213,In_681);
nor U2323 (N_2323,In_431,In_33);
nor U2324 (N_2324,In_235,In_179);
nor U2325 (N_2325,In_237,In_368);
or U2326 (N_2326,In_247,In_119);
nor U2327 (N_2327,In_426,In_695);
nor U2328 (N_2328,In_447,In_602);
nand U2329 (N_2329,In_724,In_626);
or U2330 (N_2330,In_41,In_9);
nand U2331 (N_2331,In_741,In_618);
or U2332 (N_2332,In_577,In_373);
or U2333 (N_2333,In_320,In_168);
and U2334 (N_2334,In_609,In_197);
nor U2335 (N_2335,In_425,In_385);
or U2336 (N_2336,In_242,In_560);
nand U2337 (N_2337,In_288,In_724);
and U2338 (N_2338,In_432,In_498);
or U2339 (N_2339,In_301,In_93);
or U2340 (N_2340,In_298,In_323);
nor U2341 (N_2341,In_508,In_162);
nor U2342 (N_2342,In_84,In_74);
or U2343 (N_2343,In_597,In_433);
nand U2344 (N_2344,In_485,In_677);
nand U2345 (N_2345,In_214,In_531);
nor U2346 (N_2346,In_269,In_730);
and U2347 (N_2347,In_421,In_243);
nor U2348 (N_2348,In_608,In_231);
or U2349 (N_2349,In_24,In_233);
nand U2350 (N_2350,In_499,In_515);
or U2351 (N_2351,In_411,In_691);
nor U2352 (N_2352,In_363,In_1);
or U2353 (N_2353,In_475,In_399);
and U2354 (N_2354,In_26,In_593);
nor U2355 (N_2355,In_452,In_159);
or U2356 (N_2356,In_743,In_222);
nand U2357 (N_2357,In_160,In_347);
or U2358 (N_2358,In_24,In_7);
and U2359 (N_2359,In_467,In_149);
nand U2360 (N_2360,In_519,In_299);
or U2361 (N_2361,In_326,In_717);
nand U2362 (N_2362,In_746,In_536);
nor U2363 (N_2363,In_710,In_28);
or U2364 (N_2364,In_624,In_396);
and U2365 (N_2365,In_12,In_178);
and U2366 (N_2366,In_56,In_163);
or U2367 (N_2367,In_643,In_469);
and U2368 (N_2368,In_250,In_530);
or U2369 (N_2369,In_689,In_622);
or U2370 (N_2370,In_451,In_732);
or U2371 (N_2371,In_134,In_368);
nor U2372 (N_2372,In_420,In_438);
nor U2373 (N_2373,In_288,In_405);
nor U2374 (N_2374,In_712,In_227);
or U2375 (N_2375,In_417,In_577);
nand U2376 (N_2376,In_277,In_229);
nor U2377 (N_2377,In_34,In_155);
nor U2378 (N_2378,In_375,In_743);
or U2379 (N_2379,In_183,In_246);
and U2380 (N_2380,In_26,In_455);
or U2381 (N_2381,In_213,In_586);
or U2382 (N_2382,In_154,In_141);
and U2383 (N_2383,In_284,In_718);
nor U2384 (N_2384,In_523,In_160);
and U2385 (N_2385,In_637,In_454);
or U2386 (N_2386,In_124,In_604);
nor U2387 (N_2387,In_649,In_371);
nor U2388 (N_2388,In_372,In_349);
or U2389 (N_2389,In_432,In_472);
or U2390 (N_2390,In_44,In_353);
and U2391 (N_2391,In_499,In_11);
nand U2392 (N_2392,In_175,In_636);
nor U2393 (N_2393,In_260,In_44);
and U2394 (N_2394,In_78,In_279);
or U2395 (N_2395,In_28,In_512);
or U2396 (N_2396,In_298,In_55);
nor U2397 (N_2397,In_636,In_262);
nor U2398 (N_2398,In_124,In_505);
nand U2399 (N_2399,In_557,In_298);
nor U2400 (N_2400,In_425,In_478);
or U2401 (N_2401,In_596,In_429);
nor U2402 (N_2402,In_239,In_310);
nand U2403 (N_2403,In_358,In_6);
nor U2404 (N_2404,In_268,In_121);
nand U2405 (N_2405,In_477,In_399);
nor U2406 (N_2406,In_626,In_537);
nor U2407 (N_2407,In_191,In_443);
and U2408 (N_2408,In_384,In_350);
and U2409 (N_2409,In_652,In_204);
nor U2410 (N_2410,In_401,In_329);
nand U2411 (N_2411,In_182,In_724);
nand U2412 (N_2412,In_192,In_718);
nor U2413 (N_2413,In_320,In_322);
and U2414 (N_2414,In_183,In_71);
nor U2415 (N_2415,In_103,In_588);
or U2416 (N_2416,In_512,In_274);
nand U2417 (N_2417,In_135,In_301);
nand U2418 (N_2418,In_644,In_395);
and U2419 (N_2419,In_226,In_411);
and U2420 (N_2420,In_139,In_434);
nand U2421 (N_2421,In_727,In_341);
and U2422 (N_2422,In_160,In_257);
and U2423 (N_2423,In_374,In_558);
nand U2424 (N_2424,In_178,In_216);
nor U2425 (N_2425,In_386,In_254);
nor U2426 (N_2426,In_71,In_285);
or U2427 (N_2427,In_180,In_671);
nor U2428 (N_2428,In_288,In_189);
and U2429 (N_2429,In_745,In_551);
or U2430 (N_2430,In_729,In_2);
nor U2431 (N_2431,In_407,In_214);
nor U2432 (N_2432,In_727,In_617);
xnor U2433 (N_2433,In_2,In_276);
and U2434 (N_2434,In_509,In_56);
nor U2435 (N_2435,In_157,In_703);
nand U2436 (N_2436,In_101,In_100);
xnor U2437 (N_2437,In_124,In_597);
and U2438 (N_2438,In_642,In_47);
nor U2439 (N_2439,In_386,In_642);
nor U2440 (N_2440,In_269,In_564);
and U2441 (N_2441,In_26,In_165);
and U2442 (N_2442,In_86,In_372);
and U2443 (N_2443,In_359,In_3);
nor U2444 (N_2444,In_415,In_665);
or U2445 (N_2445,In_30,In_81);
nor U2446 (N_2446,In_706,In_572);
nand U2447 (N_2447,In_198,In_148);
nand U2448 (N_2448,In_266,In_675);
or U2449 (N_2449,In_126,In_106);
nor U2450 (N_2450,In_611,In_253);
or U2451 (N_2451,In_360,In_214);
nand U2452 (N_2452,In_479,In_423);
xnor U2453 (N_2453,In_56,In_207);
and U2454 (N_2454,In_710,In_414);
and U2455 (N_2455,In_191,In_176);
or U2456 (N_2456,In_387,In_173);
and U2457 (N_2457,In_558,In_747);
nor U2458 (N_2458,In_600,In_521);
nor U2459 (N_2459,In_143,In_364);
nor U2460 (N_2460,In_0,In_569);
or U2461 (N_2461,In_360,In_484);
nand U2462 (N_2462,In_713,In_233);
nor U2463 (N_2463,In_238,In_667);
xnor U2464 (N_2464,In_189,In_501);
and U2465 (N_2465,In_547,In_566);
or U2466 (N_2466,In_19,In_584);
or U2467 (N_2467,In_406,In_47);
or U2468 (N_2468,In_141,In_48);
and U2469 (N_2469,In_227,In_233);
and U2470 (N_2470,In_225,In_456);
or U2471 (N_2471,In_6,In_550);
nor U2472 (N_2472,In_614,In_541);
and U2473 (N_2473,In_597,In_167);
nor U2474 (N_2474,In_699,In_238);
and U2475 (N_2475,In_359,In_41);
or U2476 (N_2476,In_261,In_576);
nand U2477 (N_2477,In_720,In_339);
or U2478 (N_2478,In_207,In_659);
and U2479 (N_2479,In_267,In_748);
nand U2480 (N_2480,In_604,In_596);
and U2481 (N_2481,In_9,In_241);
nand U2482 (N_2482,In_308,In_543);
and U2483 (N_2483,In_509,In_409);
and U2484 (N_2484,In_472,In_704);
nor U2485 (N_2485,In_48,In_493);
or U2486 (N_2486,In_80,In_393);
and U2487 (N_2487,In_693,In_122);
nor U2488 (N_2488,In_738,In_323);
nand U2489 (N_2489,In_715,In_491);
and U2490 (N_2490,In_161,In_605);
nand U2491 (N_2491,In_15,In_605);
nand U2492 (N_2492,In_392,In_440);
xnor U2493 (N_2493,In_437,In_477);
or U2494 (N_2494,In_54,In_486);
nand U2495 (N_2495,In_22,In_25);
and U2496 (N_2496,In_122,In_405);
nor U2497 (N_2497,In_181,In_346);
nand U2498 (N_2498,In_580,In_742);
or U2499 (N_2499,In_179,In_276);
or U2500 (N_2500,N_1835,N_2040);
or U2501 (N_2501,N_1467,N_1063);
nand U2502 (N_2502,N_777,N_351);
or U2503 (N_2503,N_677,N_2307);
nor U2504 (N_2504,N_1634,N_95);
or U2505 (N_2505,N_214,N_1828);
or U2506 (N_2506,N_115,N_103);
and U2507 (N_2507,N_2460,N_2100);
nand U2508 (N_2508,N_843,N_2137);
nand U2509 (N_2509,N_1559,N_528);
and U2510 (N_2510,N_1327,N_1888);
nor U2511 (N_2511,N_2171,N_1173);
nor U2512 (N_2512,N_489,N_1268);
nor U2513 (N_2513,N_2064,N_1245);
and U2514 (N_2514,N_2116,N_1961);
nor U2515 (N_2515,N_1930,N_1456);
nand U2516 (N_2516,N_189,N_405);
and U2517 (N_2517,N_1913,N_1366);
nand U2518 (N_2518,N_2183,N_1059);
nand U2519 (N_2519,N_1358,N_597);
and U2520 (N_2520,N_442,N_1717);
nor U2521 (N_2521,N_270,N_308);
or U2522 (N_2522,N_431,N_1161);
nand U2523 (N_2523,N_2120,N_1217);
and U2524 (N_2524,N_1962,N_290);
xor U2525 (N_2525,N_2434,N_1834);
and U2526 (N_2526,N_1931,N_666);
and U2527 (N_2527,N_465,N_1228);
and U2528 (N_2528,N_1738,N_2325);
and U2529 (N_2529,N_1874,N_2202);
xor U2530 (N_2530,N_482,N_1302);
or U2531 (N_2531,N_1723,N_1530);
nand U2532 (N_2532,N_965,N_1239);
and U2533 (N_2533,N_2396,N_1455);
nor U2534 (N_2534,N_163,N_538);
nand U2535 (N_2535,N_1957,N_704);
or U2536 (N_2536,N_1205,N_512);
nand U2537 (N_2537,N_640,N_1461);
or U2538 (N_2538,N_1504,N_1269);
nand U2539 (N_2539,N_1346,N_649);
or U2540 (N_2540,N_2005,N_1494);
and U2541 (N_2541,N_230,N_1544);
nor U2542 (N_2542,N_1785,N_1739);
nand U2543 (N_2543,N_1436,N_510);
and U2544 (N_2544,N_490,N_2132);
and U2545 (N_2545,N_4,N_746);
nor U2546 (N_2546,N_626,N_2170);
nor U2547 (N_2547,N_1534,N_2157);
and U2548 (N_2548,N_1577,N_1183);
nand U2549 (N_2549,N_1978,N_2442);
nor U2550 (N_2550,N_1103,N_132);
nor U2551 (N_2551,N_2255,N_121);
and U2552 (N_2552,N_893,N_585);
nor U2553 (N_2553,N_850,N_1630);
or U2554 (N_2554,N_1914,N_1378);
and U2555 (N_2555,N_552,N_1151);
nand U2556 (N_2556,N_225,N_1940);
or U2557 (N_2557,N_1043,N_1602);
nand U2558 (N_2558,N_1648,N_1411);
or U2559 (N_2559,N_1180,N_190);
and U2560 (N_2560,N_543,N_1772);
and U2561 (N_2561,N_2181,N_1793);
nor U2562 (N_2562,N_497,N_571);
nand U2563 (N_2563,N_1475,N_56);
or U2564 (N_2564,N_1365,N_178);
and U2565 (N_2565,N_999,N_355);
nor U2566 (N_2566,N_1748,N_1109);
nor U2567 (N_2567,N_200,N_2420);
nand U2568 (N_2568,N_1471,N_1274);
nand U2569 (N_2569,N_1572,N_940);
nand U2570 (N_2570,N_411,N_2451);
and U2571 (N_2571,N_1729,N_2191);
nand U2572 (N_2572,N_705,N_1995);
nor U2573 (N_2573,N_1097,N_1464);
or U2574 (N_2574,N_971,N_21);
or U2575 (N_2575,N_1155,N_1955);
nand U2576 (N_2576,N_984,N_2357);
xnor U2577 (N_2577,N_1380,N_1340);
nor U2578 (N_2578,N_244,N_1560);
and U2579 (N_2579,N_743,N_1871);
nor U2580 (N_2580,N_111,N_2187);
nor U2581 (N_2581,N_1580,N_2407);
nor U2582 (N_2582,N_2167,N_2054);
nand U2583 (N_2583,N_129,N_51);
xnor U2584 (N_2584,N_1112,N_1565);
and U2585 (N_2585,N_2402,N_1714);
or U2586 (N_2586,N_2382,N_550);
nor U2587 (N_2587,N_906,N_1053);
nor U2588 (N_2588,N_1869,N_384);
xor U2589 (N_2589,N_2465,N_20);
nor U2590 (N_2590,N_1332,N_622);
nand U2591 (N_2591,N_418,N_2152);
nor U2592 (N_2592,N_2343,N_172);
nor U2593 (N_2593,N_2332,N_32);
and U2594 (N_2594,N_540,N_2188);
xnor U2595 (N_2595,N_2318,N_2474);
nor U2596 (N_2596,N_1665,N_962);
or U2597 (N_2597,N_493,N_2436);
or U2598 (N_2598,N_616,N_1140);
and U2599 (N_2599,N_1562,N_495);
or U2600 (N_2600,N_1862,N_816);
nand U2601 (N_2601,N_881,N_2419);
nand U2602 (N_2602,N_1633,N_1604);
or U2603 (N_2603,N_900,N_2486);
xor U2604 (N_2604,N_1867,N_2021);
or U2605 (N_2605,N_1883,N_2240);
or U2606 (N_2606,N_2430,N_104);
and U2607 (N_2607,N_1376,N_1243);
nor U2608 (N_2608,N_2118,N_2374);
and U2609 (N_2609,N_1447,N_861);
and U2610 (N_2610,N_555,N_1042);
or U2611 (N_2611,N_557,N_1229);
nand U2612 (N_2612,N_695,N_2391);
and U2613 (N_2613,N_2192,N_263);
nor U2614 (N_2614,N_1550,N_633);
or U2615 (N_2615,N_224,N_109);
nor U2616 (N_2616,N_2409,N_358);
nor U2617 (N_2617,N_1400,N_1997);
nor U2618 (N_2618,N_2199,N_853);
nand U2619 (N_2619,N_1727,N_637);
and U2620 (N_2620,N_1600,N_83);
nand U2621 (N_2621,N_1527,N_381);
nor U2622 (N_2622,N_422,N_1209);
nand U2623 (N_2623,N_2003,N_1508);
and U2624 (N_2624,N_309,N_154);
nand U2625 (N_2625,N_1847,N_710);
or U2626 (N_2626,N_1429,N_302);
and U2627 (N_2627,N_1935,N_1421);
nor U2628 (N_2628,N_1003,N_272);
and U2629 (N_2629,N_1775,N_955);
or U2630 (N_2630,N_1419,N_92);
nand U2631 (N_2631,N_2186,N_1556);
and U2632 (N_2632,N_2421,N_1176);
or U2633 (N_2633,N_1282,N_1519);
nor U2634 (N_2634,N_797,N_1331);
and U2635 (N_2635,N_1982,N_213);
nor U2636 (N_2636,N_838,N_1959);
or U2637 (N_2637,N_602,N_2154);
or U2638 (N_2638,N_628,N_1902);
nand U2639 (N_2639,N_2111,N_1702);
or U2640 (N_2640,N_2238,N_2443);
or U2641 (N_2641,N_979,N_1855);
or U2642 (N_2642,N_236,N_1473);
nand U2643 (N_2643,N_1373,N_1732);
nand U2644 (N_2644,N_1683,N_278);
nand U2645 (N_2645,N_739,N_1949);
nand U2646 (N_2646,N_125,N_265);
nand U2647 (N_2647,N_2237,N_929);
nor U2648 (N_2648,N_1031,N_1258);
or U2649 (N_2649,N_678,N_76);
nor U2650 (N_2650,N_1334,N_1740);
nor U2651 (N_2651,N_2161,N_1706);
and U2652 (N_2652,N_854,N_417);
nor U2653 (N_2653,N_1001,N_983);
nor U2654 (N_2654,N_1184,N_399);
or U2655 (N_2655,N_232,N_2112);
nor U2656 (N_2656,N_1244,N_1008);
nor U2657 (N_2657,N_1768,N_2035);
nor U2658 (N_2658,N_261,N_2148);
and U2659 (N_2659,N_35,N_2057);
or U2660 (N_2660,N_359,N_1004);
nand U2661 (N_2661,N_2014,N_477);
and U2662 (N_2662,N_1975,N_392);
nor U2663 (N_2663,N_801,N_1110);
and U2664 (N_2664,N_744,N_1320);
nor U2665 (N_2665,N_305,N_541);
nand U2666 (N_2666,N_573,N_1388);
and U2667 (N_2667,N_108,N_463);
and U2668 (N_2668,N_1827,N_674);
and U2669 (N_2669,N_1589,N_1045);
nand U2670 (N_2670,N_1126,N_1082);
nor U2671 (N_2671,N_1623,N_480);
or U2672 (N_2672,N_539,N_349);
or U2673 (N_2673,N_294,N_1357);
and U2674 (N_2674,N_1535,N_2060);
or U2675 (N_2675,N_1284,N_1505);
and U2676 (N_2676,N_1197,N_694);
nand U2677 (N_2677,N_1312,N_395);
nand U2678 (N_2678,N_2252,N_909);
and U2679 (N_2679,N_269,N_2453);
and U2680 (N_2680,N_327,N_128);
or U2681 (N_2681,N_1105,N_2462);
or U2682 (N_2682,N_374,N_1277);
nand U2683 (N_2683,N_1104,N_2302);
nor U2684 (N_2684,N_394,N_2194);
nand U2685 (N_2685,N_255,N_2031);
nand U2686 (N_2686,N_2156,N_1860);
nand U2687 (N_2687,N_71,N_28);
and U2688 (N_2688,N_260,N_1487);
nand U2689 (N_2689,N_36,N_2445);
xnor U2690 (N_2690,N_2071,N_2044);
xnor U2691 (N_2691,N_1583,N_82);
or U2692 (N_2692,N_2455,N_918);
and U2693 (N_2693,N_846,N_855);
or U2694 (N_2694,N_1248,N_1543);
or U2695 (N_2695,N_1987,N_1697);
nand U2696 (N_2696,N_1756,N_329);
nand U2697 (N_2697,N_413,N_1742);
or U2698 (N_2698,N_2036,N_1313);
and U2699 (N_2699,N_1518,N_2018);
nand U2700 (N_2700,N_868,N_1669);
or U2701 (N_2701,N_375,N_1520);
nand U2702 (N_2702,N_2109,N_1865);
or U2703 (N_2703,N_2323,N_2398);
nor U2704 (N_2704,N_1611,N_2433);
nand U2705 (N_2705,N_1010,N_2211);
xor U2706 (N_2706,N_2053,N_1100);
and U2707 (N_2707,N_1442,N_949);
and U2708 (N_2708,N_670,N_741);
and U2709 (N_2709,N_581,N_1191);
nor U2710 (N_2710,N_2272,N_234);
and U2711 (N_2711,N_499,N_1722);
or U2712 (N_2712,N_1426,N_1310);
xnor U2713 (N_2713,N_13,N_2491);
or U2714 (N_2714,N_1350,N_1592);
nand U2715 (N_2715,N_858,N_1786);
and U2716 (N_2716,N_1657,N_85);
and U2717 (N_2717,N_523,N_1120);
or U2718 (N_2718,N_1726,N_66);
nand U2719 (N_2719,N_1292,N_453);
and U2720 (N_2720,N_1963,N_2178);
and U2721 (N_2721,N_1483,N_423);
nand U2722 (N_2722,N_2269,N_2144);
and U2723 (N_2723,N_1896,N_684);
nand U2724 (N_2724,N_1445,N_830);
nor U2725 (N_2725,N_231,N_867);
and U2726 (N_2726,N_1850,N_1776);
xnor U2727 (N_2727,N_1368,N_1208);
nor U2728 (N_2728,N_1540,N_937);
nor U2729 (N_2729,N_911,N_1462);
nor U2730 (N_2730,N_316,N_1230);
nor U2731 (N_2731,N_2114,N_1985);
nor U2732 (N_2732,N_1585,N_661);
nand U2733 (N_2733,N_2390,N_604);
nand U2734 (N_2734,N_2262,N_509);
or U2735 (N_2735,N_1782,N_880);
and U2736 (N_2736,N_724,N_1947);
and U2737 (N_2737,N_779,N_114);
or U2738 (N_2738,N_1492,N_587);
nand U2739 (N_2739,N_2025,N_412);
and U2740 (N_2740,N_1843,N_923);
or U2741 (N_2741,N_1907,N_1851);
nand U2742 (N_2742,N_1238,N_2131);
nand U2743 (N_2743,N_1127,N_1141);
nand U2744 (N_2744,N_1264,N_169);
nor U2745 (N_2745,N_2206,N_2038);
nand U2746 (N_2746,N_451,N_2280);
or U2747 (N_2747,N_414,N_2408);
nor U2748 (N_2748,N_1991,N_1122);
nand U2749 (N_2749,N_81,N_2329);
and U2750 (N_2750,N_2452,N_425);
xor U2751 (N_2751,N_69,N_1964);
or U2752 (N_2752,N_45,N_2427);
nor U2753 (N_2753,N_688,N_2082);
or U2754 (N_2754,N_781,N_242);
or U2755 (N_2755,N_2454,N_809);
and U2756 (N_2756,N_870,N_2239);
nand U2757 (N_2757,N_2356,N_648);
or U2758 (N_2758,N_565,N_470);
nor U2759 (N_2759,N_788,N_2022);
nand U2760 (N_2760,N_496,N_1397);
nand U2761 (N_2761,N_1747,N_1133);
nand U2762 (N_2762,N_542,N_426);
nand U2763 (N_2763,N_2294,N_2285);
xnor U2764 (N_2764,N_2130,N_787);
and U2765 (N_2765,N_2480,N_876);
or U2766 (N_2766,N_525,N_2028);
and U2767 (N_2767,N_2087,N_2043);
and U2768 (N_2768,N_1435,N_124);
nor U2769 (N_2769,N_450,N_1584);
or U2770 (N_2770,N_1646,N_1115);
nor U2771 (N_2771,N_1872,N_577);
nor U2772 (N_2772,N_348,N_2337);
nor U2773 (N_2773,N_837,N_1039);
or U2774 (N_2774,N_1878,N_2290);
and U2775 (N_2775,N_737,N_959);
nor U2776 (N_2776,N_2387,N_1825);
nand U2777 (N_2777,N_1130,N_530);
nor U2778 (N_2778,N_2000,N_2256);
nor U2779 (N_2779,N_2135,N_1612);
and U2780 (N_2780,N_1614,N_975);
or U2781 (N_2781,N_1143,N_1037);
nor U2782 (N_2782,N_352,N_2091);
nor U2783 (N_2783,N_1628,N_760);
nand U2784 (N_2784,N_895,N_734);
and U2785 (N_2785,N_296,N_2159);
or U2786 (N_2786,N_222,N_706);
and U2787 (N_2787,N_1317,N_1086);
nor U2788 (N_2788,N_2201,N_2483);
or U2789 (N_2789,N_141,N_1758);
and U2790 (N_2790,N_1676,N_1136);
or U2791 (N_2791,N_262,N_1725);
nand U2792 (N_2792,N_215,N_1062);
and U2793 (N_2793,N_102,N_806);
nor U2794 (N_2794,N_410,N_2142);
and U2795 (N_2795,N_1558,N_601);
and U2796 (N_2796,N_1568,N_2140);
nor U2797 (N_2797,N_2127,N_2316);
or U2798 (N_2798,N_1123,N_1236);
nor U2799 (N_2799,N_2342,N_576);
nor U2800 (N_2800,N_2386,N_562);
or U2801 (N_2801,N_928,N_350);
nand U2802 (N_2802,N_2089,N_1371);
nor U2803 (N_2803,N_815,N_1387);
and U2804 (N_2804,N_2271,N_729);
or U2805 (N_2805,N_745,N_170);
or U2806 (N_2806,N_1552,N_1099);
or U2807 (N_2807,N_2418,N_2414);
nor U2808 (N_2808,N_94,N_757);
nand U2809 (N_2809,N_1261,N_1305);
nand U2810 (N_2810,N_1453,N_2469);
nand U2811 (N_2811,N_1672,N_1621);
xor U2812 (N_2812,N_2383,N_844);
and U2813 (N_2813,N_2446,N_641);
and U2814 (N_2814,N_1854,N_651);
nand U2815 (N_2815,N_173,N_1249);
nand U2816 (N_2816,N_504,N_933);
and U2817 (N_2817,N_1641,N_1916);
and U2818 (N_2818,N_84,N_723);
and U2819 (N_2819,N_2079,N_1029);
or U2820 (N_2820,N_87,N_293);
or U2821 (N_2821,N_2253,N_2004);
nor U2822 (N_2822,N_1817,N_1574);
nor U2823 (N_2823,N_424,N_941);
nor U2824 (N_2824,N_357,N_1200);
and U2825 (N_2825,N_218,N_1790);
and U2826 (N_2826,N_123,N_1068);
and U2827 (N_2827,N_2248,N_1246);
and U2828 (N_2828,N_1255,N_2069);
or U2829 (N_2829,N_363,N_890);
nand U2830 (N_2830,N_653,N_795);
nor U2831 (N_2831,N_159,N_2174);
and U2832 (N_2832,N_1360,N_1076);
and U2833 (N_2833,N_1025,N_2432);
and U2834 (N_2834,N_2373,N_2169);
or U2835 (N_2835,N_954,N_511);
or U2836 (N_2836,N_2422,N_1212);
nor U2837 (N_2837,N_2412,N_1477);
nand U2838 (N_2838,N_995,N_464);
nand U2839 (N_2839,N_1868,N_391);
or U2840 (N_2840,N_663,N_2493);
nand U2841 (N_2841,N_1876,N_2065);
or U2842 (N_2842,N_238,N_1203);
nand U2843 (N_2843,N_2205,N_2377);
and U2844 (N_2844,N_2050,N_188);
nand U2845 (N_2845,N_1794,N_1698);
nand U2846 (N_2846,N_2284,N_1015);
xor U2847 (N_2847,N_687,N_1958);
or U2848 (N_2848,N_680,N_2458);
nand U2849 (N_2849,N_774,N_1194);
nor U2850 (N_2850,N_782,N_2384);
nor U2851 (N_2851,N_401,N_80);
or U2852 (N_2852,N_1681,N_1199);
and U2853 (N_2853,N_1791,N_2311);
nand U2854 (N_2854,N_513,N_2006);
xor U2855 (N_2855,N_1418,N_1899);
and U2856 (N_2856,N_501,N_1500);
and U2857 (N_2857,N_1448,N_47);
nand U2858 (N_2858,N_2499,N_1019);
nor U2859 (N_2859,N_1960,N_945);
or U2860 (N_2860,N_208,N_1085);
nand U2861 (N_2861,N_246,N_2180);
nor U2862 (N_2862,N_789,N_627);
and U2863 (N_2863,N_1348,N_1044);
and U2864 (N_2864,N_972,N_2415);
nor U2865 (N_2865,N_2228,N_2009);
nand U2866 (N_2866,N_676,N_2196);
nand U2867 (N_2867,N_268,N_1846);
nor U2868 (N_2868,N_2101,N_191);
and U2869 (N_2869,N_1829,N_55);
nand U2870 (N_2870,N_718,N_2244);
and U2871 (N_2871,N_829,N_52);
and U2872 (N_2872,N_1121,N_2147);
or U2873 (N_2873,N_1637,N_1128);
or U2874 (N_2874,N_1428,N_560);
and U2875 (N_2875,N_1384,N_1165);
nand U2876 (N_2876,N_408,N_2092);
and U2877 (N_2877,N_1146,N_1036);
and U2878 (N_2878,N_1303,N_393);
or U2879 (N_2879,N_2251,N_1444);
and U2880 (N_2880,N_767,N_2405);
or U2881 (N_2881,N_717,N_2163);
nor U2882 (N_2882,N_1569,N_40);
nor U2883 (N_2883,N_1158,N_235);
and U2884 (N_2884,N_494,N_2084);
nor U2885 (N_2885,N_1273,N_112);
nor U2886 (N_2886,N_652,N_491);
or U2887 (N_2887,N_2497,N_1406);
or U2888 (N_2888,N_2304,N_693);
nand U2889 (N_2889,N_754,N_946);
and U2890 (N_2890,N_775,N_2105);
nor U2891 (N_2891,N_1688,N_1414);
and U2892 (N_2892,N_1478,N_1342);
nand U2893 (N_2893,N_1318,N_1863);
and U2894 (N_2894,N_786,N_2371);
and U2895 (N_2895,N_1624,N_1286);
or U2896 (N_2896,N_1266,N_2441);
nand U2897 (N_2897,N_2472,N_1466);
or U2898 (N_2898,N_1830,N_1711);
xnor U2899 (N_2899,N_385,N_1150);
and U2900 (N_2900,N_313,N_1073);
or U2901 (N_2901,N_179,N_1117);
nor U2902 (N_2902,N_713,N_1696);
and U2903 (N_2903,N_2039,N_2265);
nand U2904 (N_2904,N_2254,N_889);
nor U2905 (N_2905,N_1710,N_593);
or U2906 (N_2906,N_939,N_1449);
and U2907 (N_2907,N_1667,N_1937);
or U2908 (N_2908,N_2347,N_1563);
nor U2909 (N_2909,N_306,N_1152);
nor U2910 (N_2910,N_756,N_368);
nand U2911 (N_2911,N_337,N_996);
nor U2912 (N_2912,N_1713,N_1898);
nand U2913 (N_2913,N_1207,N_1052);
and U2914 (N_2914,N_605,N_207);
nand U2915 (N_2915,N_2023,N_1503);
or U2916 (N_2916,N_379,N_1824);
nor U2917 (N_2917,N_460,N_182);
or U2918 (N_2918,N_2207,N_897);
and U2919 (N_2919,N_921,N_1906);
and U2920 (N_2920,N_1330,N_1700);
and U2921 (N_2921,N_387,N_2032);
nor U2922 (N_2922,N_17,N_1745);
nor U2923 (N_2923,N_898,N_582);
and U2924 (N_2924,N_143,N_2176);
and U2925 (N_2925,N_1581,N_1575);
nand U2926 (N_2926,N_2151,N_669);
nand U2927 (N_2927,N_1820,N_1061);
nand U2928 (N_2928,N_221,N_619);
or U2929 (N_2929,N_2463,N_1755);
nand U2930 (N_2930,N_551,N_1452);
nand U2931 (N_2931,N_2326,N_2479);
or U2932 (N_2932,N_273,N_570);
or U2933 (N_2933,N_1257,N_1285);
nand U2934 (N_2934,N_728,N_378);
nand U2935 (N_2935,N_1070,N_1853);
nand U2936 (N_2936,N_583,N_961);
or U2937 (N_2937,N_1805,N_1369);
and U2938 (N_2938,N_1027,N_1759);
or U2939 (N_2939,N_353,N_2155);
nor U2940 (N_2940,N_1016,N_982);
and U2941 (N_2941,N_1513,N_1107);
nor U2942 (N_2942,N_377,N_877);
or U2943 (N_2943,N_2321,N_1554);
and U2944 (N_2944,N_1389,N_287);
and U2945 (N_2945,N_2212,N_1567);
nor U2946 (N_2946,N_1712,N_1210);
nor U2947 (N_2947,N_1910,N_402);
and U2948 (N_2948,N_985,N_1803);
and U2949 (N_2949,N_742,N_991);
or U2950 (N_2950,N_1193,N_951);
nand U2951 (N_2951,N_434,N_160);
and U2952 (N_2952,N_2333,N_311);
nor U2953 (N_2953,N_333,N_1135);
nor U2954 (N_2954,N_968,N_318);
nand U2955 (N_2955,N_1415,N_1674);
or U2956 (N_2956,N_2428,N_635);
nand U2957 (N_2957,N_1101,N_2289);
or U2958 (N_2958,N_186,N_365);
and U2959 (N_2959,N_2426,N_2331);
or U2960 (N_2960,N_2413,N_46);
nor U2961 (N_2961,N_1892,N_1399);
or U2962 (N_2962,N_2217,N_1516);
and U2963 (N_2963,N_731,N_2278);
nor U2964 (N_2964,N_1139,N_2264);
or U2965 (N_2965,N_1716,N_1757);
nand U2966 (N_2966,N_1591,N_1861);
nor U2967 (N_2967,N_39,N_847);
or U2968 (N_2968,N_478,N_134);
or U2969 (N_2969,N_1922,N_343);
nand U2970 (N_2970,N_2073,N_1610);
nor U2971 (N_2971,N_1760,N_904);
nor U2972 (N_2972,N_1590,N_832);
nor U2973 (N_2973,N_233,N_664);
and U2974 (N_2974,N_53,N_1762);
nor U2975 (N_2975,N_2076,N_326);
and U2976 (N_2976,N_1643,N_671);
nor U2977 (N_2977,N_2083,N_1124);
nand U2978 (N_2978,N_1642,N_152);
nor U2979 (N_2979,N_2037,N_1116);
or U2980 (N_2980,N_1034,N_1555);
nor U2981 (N_2981,N_1576,N_771);
nor U2982 (N_2982,N_924,N_620);
nand U2983 (N_2983,N_1788,N_1687);
xor U2984 (N_2984,N_712,N_503);
nand U2985 (N_2985,N_1780,N_1531);
nand U2986 (N_2986,N_506,N_1055);
nand U2987 (N_2987,N_823,N_559);
nor U2988 (N_2988,N_2431,N_2358);
and U2989 (N_2989,N_989,N_416);
nand U2990 (N_2990,N_133,N_1904);
nand U2991 (N_2991,N_1054,N_1524);
or U2992 (N_2992,N_2214,N_698);
nand U2993 (N_2993,N_798,N_1915);
nand U2994 (N_2994,N_1557,N_2286);
nor U2995 (N_2995,N_280,N_1538);
nor U2996 (N_2996,N_324,N_1942);
or U2997 (N_2997,N_715,N_1608);
nor U2998 (N_2998,N_341,N_507);
and U2999 (N_2999,N_1781,N_2034);
or U3000 (N_3000,N_1849,N_1095);
and U3001 (N_3001,N_2496,N_1489);
and U3002 (N_3002,N_443,N_1118);
nor U3003 (N_3003,N_1020,N_2223);
and U3004 (N_3004,N_1684,N_1361);
or U3005 (N_3005,N_1398,N_15);
nor U3006 (N_3006,N_210,N_2138);
nor U3007 (N_3007,N_315,N_1166);
and U3008 (N_3008,N_404,N_2411);
and U3009 (N_3009,N_2494,N_122);
or U3010 (N_3010,N_660,N_812);
nand U3011 (N_3011,N_1689,N_2464);
nand U3012 (N_3012,N_1315,N_2344);
and U3013 (N_3013,N_749,N_119);
and U3014 (N_3014,N_2267,N_88);
nor U3015 (N_3015,N_732,N_1321);
and U3016 (N_3016,N_2010,N_2327);
and U3017 (N_3017,N_901,N_1986);
nor U3018 (N_3018,N_1751,N_1972);
or U3019 (N_3019,N_1265,N_987);
or U3020 (N_3020,N_415,N_1149);
nor U3021 (N_3021,N_2417,N_176);
nor U3022 (N_3022,N_2197,N_524);
or U3023 (N_3023,N_2008,N_2328);
nor U3024 (N_3024,N_701,N_1966);
and U3025 (N_3025,N_153,N_1067);
nor U3026 (N_3026,N_1901,N_1779);
nor U3027 (N_3027,N_2125,N_407);
nor U3028 (N_3028,N_1778,N_527);
nand U3029 (N_3029,N_813,N_865);
or U3030 (N_3030,N_2287,N_2380);
and U3031 (N_3031,N_2361,N_2222);
nand U3032 (N_3032,N_2393,N_646);
nor U3033 (N_3033,N_1952,N_1763);
or U3034 (N_3034,N_1511,N_2002);
nor U3035 (N_3035,N_1187,N_790);
nand U3036 (N_3036,N_271,N_1606);
or U3037 (N_3037,N_1064,N_1311);
or U3038 (N_3038,N_1647,N_1724);
nand U3039 (N_3039,N_859,N_1597);
and U3040 (N_3040,N_1324,N_396);
and U3041 (N_3041,N_2242,N_1227);
and U3042 (N_3042,N_607,N_1434);
or U3043 (N_3043,N_1336,N_520);
or U3044 (N_3044,N_796,N_1690);
or U3045 (N_3045,N_492,N_2438);
or U3046 (N_3046,N_1660,N_2338);
or U3047 (N_3047,N_1521,N_310);
xor U3048 (N_3048,N_515,N_852);
nand U3049 (N_3049,N_2158,N_1968);
or U3050 (N_3050,N_1102,N_2113);
and U3051 (N_3051,N_2012,N_38);
xnor U3052 (N_3052,N_2282,N_1894);
nor U3053 (N_3053,N_2047,N_1480);
or U3054 (N_3054,N_851,N_166);
nor U3055 (N_3055,N_1638,N_572);
or U3056 (N_3056,N_1806,N_610);
or U3057 (N_3057,N_2365,N_1733);
or U3058 (N_3058,N_1967,N_1743);
and U3059 (N_3059,N_2261,N_875);
nand U3060 (N_3060,N_455,N_2310);
and U3061 (N_3061,N_2208,N_30);
or U3062 (N_3062,N_1407,N_828);
and U3063 (N_3063,N_679,N_397);
nor U3064 (N_3064,N_783,N_2334);
and U3065 (N_3065,N_1186,N_1917);
nand U3066 (N_3066,N_2165,N_1394);
nand U3067 (N_3067,N_1201,N_508);
nor U3068 (N_3068,N_31,N_804);
and U3069 (N_3069,N_600,N_70);
or U3070 (N_3070,N_64,N_2103);
or U3071 (N_3071,N_1222,N_2243);
nor U3072 (N_3072,N_3,N_1948);
nand U3073 (N_3073,N_747,N_289);
nor U3074 (N_3074,N_1619,N_645);
nor U3075 (N_3075,N_300,N_93);
nand U3076 (N_3076,N_252,N_1490);
and U3077 (N_3077,N_2257,N_1114);
and U3078 (N_3078,N_773,N_1981);
or U3079 (N_3079,N_2185,N_1163);
nor U3080 (N_3080,N_1593,N_1432);
nor U3081 (N_3081,N_62,N_34);
or U3082 (N_3082,N_869,N_2094);
nor U3083 (N_3083,N_354,N_2179);
nor U3084 (N_3084,N_986,N_964);
and U3085 (N_3085,N_856,N_33);
nor U3086 (N_3086,N_636,N_1564);
or U3087 (N_3087,N_1771,N_1433);
nor U3088 (N_3088,N_1046,N_1164);
nand U3089 (N_3089,N_1137,N_2234);
and U3090 (N_3090,N_2226,N_1705);
nand U3091 (N_3091,N_1012,N_175);
nand U3092 (N_3092,N_866,N_445);
nand U3093 (N_3093,N_1300,N_12);
and U3094 (N_3094,N_483,N_2410);
or U3095 (N_3095,N_1682,N_1980);
nand U3096 (N_3096,N_2141,N_2070);
nand U3097 (N_3097,N_1486,N_2341);
or U3098 (N_3098,N_1801,N_2400);
nor U3099 (N_3099,N_922,N_1472);
nand U3100 (N_3100,N_1603,N_1658);
or U3101 (N_3101,N_194,N_696);
nor U3102 (N_3102,N_691,N_258);
nand U3103 (N_3103,N_1897,N_1219);
or U3104 (N_3104,N_1509,N_1024);
and U3105 (N_3105,N_871,N_992);
nand U3106 (N_3106,N_817,N_1145);
and U3107 (N_3107,N_361,N_217);
nand U3108 (N_3108,N_283,N_2198);
or U3109 (N_3109,N_130,N_27);
nor U3110 (N_3110,N_1457,N_1969);
nand U3111 (N_3111,N_662,N_1636);
nor U3112 (N_3112,N_91,N_9);
nand U3113 (N_3113,N_764,N_284);
and U3114 (N_3114,N_1218,N_325);
nor U3115 (N_3115,N_1525,N_2077);
or U3116 (N_3116,N_1328,N_997);
and U3117 (N_3117,N_629,N_177);
and U3118 (N_3118,N_1936,N_2231);
nor U3119 (N_3119,N_934,N_1167);
nor U3120 (N_3120,N_1233,N_2362);
nor U3121 (N_3121,N_19,N_2306);
nand U3122 (N_3122,N_1291,N_2061);
and U3123 (N_3123,N_948,N_1338);
or U3124 (N_3124,N_762,N_969);
nor U3125 (N_3125,N_1177,N_58);
nand U3126 (N_3126,N_2189,N_1996);
nand U3127 (N_3127,N_487,N_1664);
or U3128 (N_3128,N_1808,N_2444);
nor U3129 (N_3129,N_532,N_1905);
xnor U3130 (N_3130,N_1402,N_574);
nand U3131 (N_3131,N_526,N_421);
nand U3132 (N_3132,N_2297,N_2081);
or U3133 (N_3133,N_1770,N_803);
and U3134 (N_3134,N_1237,N_346);
nand U3135 (N_3135,N_110,N_1413);
or U3136 (N_3136,N_386,N_667);
or U3137 (N_3137,N_2015,N_903);
and U3138 (N_3138,N_266,N_248);
nand U3139 (N_3139,N_599,N_25);
nand U3140 (N_3140,N_466,N_1873);
nor U3141 (N_3141,N_2200,N_2193);
and U3142 (N_3142,N_759,N_2369);
or U3143 (N_3143,N_1491,N_1446);
nand U3144 (N_3144,N_2215,N_566);
and U3145 (N_3145,N_2182,N_1038);
nand U3146 (N_3146,N_1852,N_1777);
or U3147 (N_3147,N_1314,N_1810);
and U3148 (N_3148,N_1071,N_370);
nor U3149 (N_3149,N_2220,N_1065);
nand U3150 (N_3150,N_1088,N_1994);
and U3151 (N_3151,N_1501,N_1250);
nor U3152 (N_3152,N_167,N_547);
and U3153 (N_3153,N_2395,N_1926);
and U3154 (N_3154,N_1998,N_1571);
and U3155 (N_3155,N_264,N_1929);
xor U3156 (N_3156,N_1221,N_780);
and U3157 (N_3157,N_1276,N_1370);
and U3158 (N_3158,N_1322,N_1225);
xor U3159 (N_3159,N_29,N_887);
nand U3160 (N_3160,N_286,N_2150);
and U3161 (N_3161,N_59,N_1953);
or U3162 (N_3162,N_1256,N_281);
nand U3163 (N_3163,N_1325,N_2467);
nor U3164 (N_3164,N_947,N_2368);
or U3165 (N_3165,N_245,N_1297);
or U3166 (N_3166,N_1213,N_708);
and U3167 (N_3167,N_1355,N_2107);
or U3168 (N_3168,N_1172,N_206);
or U3169 (N_3169,N_1923,N_1058);
nand U3170 (N_3170,N_957,N_736);
or U3171 (N_3171,N_101,N_1427);
nand U3172 (N_3172,N_1841,N_1971);
or U3173 (N_3173,N_142,N_751);
and U3174 (N_3174,N_1579,N_882);
xnor U3175 (N_3175,N_2017,N_2330);
and U3176 (N_3176,N_533,N_1512);
nand U3177 (N_3177,N_468,N_1864);
and U3178 (N_3178,N_1170,N_500);
or U3179 (N_3179,N_1048,N_535);
or U3180 (N_3180,N_1481,N_403);
and U3181 (N_3181,N_720,N_943);
and U3182 (N_3182,N_1206,N_2074);
nor U3183 (N_3183,N_149,N_914);
nor U3184 (N_3184,N_1588,N_14);
nor U3185 (N_3185,N_138,N_1226);
nand U3186 (N_3186,N_86,N_126);
nand U3187 (N_3187,N_2301,N_1079);
and U3188 (N_3188,N_2128,N_1459);
nand U3189 (N_3189,N_274,N_634);
or U3190 (N_3190,N_400,N_1013);
nor U3191 (N_3191,N_1234,N_1840);
xnor U3192 (N_3192,N_709,N_2134);
nand U3193 (N_3193,N_2404,N_1005);
or U3194 (N_3194,N_2473,N_2363);
nand U3195 (N_3195,N_1032,N_784);
xor U3196 (N_3196,N_2489,N_611);
and U3197 (N_3197,N_1377,N_656);
xnor U3198 (N_3198,N_1323,N_1);
nand U3199 (N_3199,N_331,N_1586);
or U3200 (N_3200,N_1335,N_41);
nor U3201 (N_3201,N_1497,N_1653);
nor U3202 (N_3202,N_1741,N_1651);
and U3203 (N_3203,N_1083,N_1337);
and U3204 (N_3204,N_1075,N_2033);
and U3205 (N_3205,N_932,N_517);
or U3206 (N_3206,N_1950,N_107);
nor U3207 (N_3207,N_598,N_1347);
or U3208 (N_3208,N_298,N_1386);
nand U3209 (N_3209,N_1262,N_2423);
or U3210 (N_3210,N_998,N_146);
and U3211 (N_3211,N_1974,N_2121);
and U3212 (N_3212,N_339,N_591);
and U3213 (N_3213,N_2459,N_1422);
and U3214 (N_3214,N_1009,N_1595);
and U3215 (N_3215,N_2117,N_2317);
and U3216 (N_3216,N_1822,N_536);
nand U3217 (N_3217,N_2350,N_11);
nor U3218 (N_3218,N_1639,N_2221);
nand U3219 (N_3219,N_1789,N_1211);
and U3220 (N_3220,N_1106,N_1147);
nor U3221 (N_3221,N_740,N_1271);
nor U3222 (N_3222,N_437,N_192);
and U3223 (N_3223,N_807,N_907);
nand U3224 (N_3224,N_697,N_1656);
or U3225 (N_3225,N_267,N_1537);
nand U3226 (N_3226,N_772,N_1663);
or U3227 (N_3227,N_1528,N_1807);
nand U3228 (N_3228,N_1270,N_2249);
and U3229 (N_3229,N_1214,N_42);
nand U3230 (N_3230,N_199,N_488);
nor U3231 (N_3231,N_1485,N_1072);
nand U3232 (N_3232,N_1272,N_456);
or U3233 (N_3233,N_1440,N_2072);
nor U3234 (N_3234,N_554,N_1615);
or U3235 (N_3235,N_2230,N_2258);
and U3236 (N_3236,N_251,N_44);
or U3237 (N_3237,N_2204,N_345);
or U3238 (N_3238,N_1469,N_317);
nor U3239 (N_3239,N_505,N_2273);
or U3240 (N_3240,N_766,N_822);
and U3241 (N_3241,N_195,N_1450);
or U3242 (N_3242,N_1319,N_2055);
and U3243 (N_3243,N_758,N_105);
or U3244 (N_3244,N_320,N_2360);
and U3245 (N_3245,N_131,N_1216);
nand U3246 (N_3246,N_1918,N_171);
nand U3247 (N_3247,N_1938,N_2241);
nand U3248 (N_3248,N_1343,N_1267);
and U3249 (N_3249,N_89,N_1951);
xnor U3250 (N_3250,N_438,N_2013);
and U3251 (N_3251,N_1814,N_2312);
nand U3252 (N_3252,N_1030,N_516);
and U3253 (N_3253,N_484,N_156);
and U3254 (N_3254,N_174,N_1744);
or U3255 (N_3255,N_1160,N_606);
and U3256 (N_3256,N_841,N_322);
nand U3257 (N_3257,N_668,N_276);
and U3258 (N_3258,N_980,N_2145);
or U3259 (N_3259,N_1769,N_1192);
or U3260 (N_3260,N_818,N_596);
nand U3261 (N_3261,N_799,N_578);
or U3262 (N_3262,N_1515,N_256);
and U3263 (N_3263,N_2353,N_150);
nor U3264 (N_3264,N_1060,N_1157);
or U3265 (N_3265,N_1675,N_1650);
or U3266 (N_3266,N_575,N_219);
nor U3267 (N_3267,N_1553,N_26);
and U3268 (N_3268,N_467,N_2450);
or U3269 (N_3269,N_1352,N_1721);
nor U3270 (N_3270,N_78,N_896);
and U3271 (N_3271,N_1988,N_180);
xor U3272 (N_3272,N_2392,N_1691);
nand U3273 (N_3273,N_237,N_157);
nand U3274 (N_3274,N_2213,N_2364);
nor U3275 (N_3275,N_755,N_1220);
nand U3276 (N_3276,N_1412,N_1026);
xor U3277 (N_3277,N_814,N_1408);
nand U3278 (N_3278,N_1495,N_1661);
nor U3279 (N_3279,N_2119,N_840);
xor U3280 (N_3280,N_2281,N_1730);
xnor U3281 (N_3281,N_334,N_106);
or U3282 (N_3282,N_2274,N_1954);
or U3283 (N_3283,N_1006,N_1668);
or U3284 (N_3284,N_436,N_2319);
and U3285 (N_3285,N_835,N_623);
or U3286 (N_3286,N_2115,N_2300);
nor U3287 (N_3287,N_373,N_1903);
and U3288 (N_3288,N_730,N_1011);
nand U3289 (N_3289,N_1077,N_1279);
nand U3290 (N_3290,N_2293,N_727);
or U3291 (N_3291,N_1734,N_976);
nand U3292 (N_3292,N_1499,N_1460);
nand U3293 (N_3293,N_994,N_113);
nand U3294 (N_3294,N_568,N_380);
and U3295 (N_3295,N_820,N_862);
or U3296 (N_3296,N_1299,N_750);
and U3297 (N_3297,N_2283,N_257);
and U3298 (N_3298,N_1925,N_1699);
and U3299 (N_3299,N_1895,N_1609);
xnor U3300 (N_3300,N_1401,N_1125);
nor U3301 (N_3301,N_916,N_748);
or U3302 (N_3302,N_162,N_277);
xnor U3303 (N_3303,N_2184,N_884);
nor U3304 (N_3304,N_1728,N_249);
or U3305 (N_3305,N_1704,N_73);
nand U3306 (N_3306,N_1890,N_546);
nand U3307 (N_3307,N_978,N_1561);
and U3308 (N_3308,N_2093,N_1566);
or U3309 (N_3309,N_1804,N_1934);
nand U3310 (N_3310,N_1787,N_609);
or U3311 (N_3311,N_223,N_958);
or U3312 (N_3312,N_1047,N_1263);
or U3313 (N_3313,N_1670,N_1307);
nor U3314 (N_3314,N_2045,N_1241);
nor U3315 (N_3315,N_514,N_2487);
nor U3316 (N_3316,N_1198,N_1635);
nand U3317 (N_3317,N_2346,N_2397);
nand U3318 (N_3318,N_1353,N_1737);
nand U3319 (N_3319,N_1298,N_1659);
and U3320 (N_3320,N_1626,N_1232);
nor U3321 (N_3321,N_569,N_761);
nand U3322 (N_3322,N_860,N_1731);
nand U3323 (N_3323,N_1393,N_439);
or U3324 (N_3324,N_1629,N_1685);
nand U3325 (N_3325,N_1391,N_37);
xnor U3326 (N_3326,N_2457,N_1224);
or U3327 (N_3327,N_685,N_1842);
nand U3328 (N_3328,N_912,N_127);
or U3329 (N_3329,N_1977,N_2052);
or U3330 (N_3330,N_873,N_1468);
nand U3331 (N_3331,N_849,N_800);
nand U3332 (N_3332,N_50,N_1185);
and U3333 (N_3333,N_878,N_1367);
and U3334 (N_3334,N_2320,N_811);
nor U3335 (N_3335,N_2129,N_1767);
and U3336 (N_3336,N_2246,N_753);
nor U3337 (N_3337,N_1773,N_2498);
nor U3338 (N_3338,N_1488,N_462);
nor U3339 (N_3339,N_1306,N_1028);
nand U3340 (N_3340,N_1761,N_1231);
nand U3341 (N_3341,N_1812,N_960);
nand U3342 (N_3342,N_672,N_888);
nor U3343 (N_3343,N_1134,N_2437);
nand U3344 (N_3344,N_776,N_2247);
nor U3345 (N_3345,N_1764,N_1041);
and U3346 (N_3346,N_763,N_79);
and U3347 (N_3347,N_239,N_319);
nor U3348 (N_3348,N_1625,N_700);
and U3349 (N_3349,N_1215,N_1720);
or U3350 (N_3350,N_2435,N_6);
and U3351 (N_3351,N_498,N_2449);
nand U3352 (N_3352,N_1884,N_1479);
or U3353 (N_3353,N_2168,N_1976);
or U3354 (N_3354,N_977,N_1735);
or U3355 (N_3355,N_2016,N_632);
or U3356 (N_3356,N_625,N_944);
or U3357 (N_3357,N_1819,N_307);
and U3358 (N_3358,N_197,N_364);
or U3359 (N_3359,N_1911,N_2299);
nand U3360 (N_3360,N_1746,N_810);
nand U3361 (N_3361,N_2232,N_1578);
and U3362 (N_3362,N_63,N_1437);
nor U3363 (N_3363,N_1056,N_658);
and U3364 (N_3364,N_647,N_556);
and U3365 (N_3365,N_1909,N_1620);
nor U3366 (N_3366,N_433,N_1154);
and U3367 (N_3367,N_1605,N_2468);
or U3368 (N_3368,N_2088,N_711);
nor U3369 (N_3369,N_183,N_1750);
or U3370 (N_3370,N_2123,N_2026);
or U3371 (N_3371,N_2288,N_2416);
nor U3372 (N_3372,N_2440,N_1021);
nor U3373 (N_3373,N_165,N_2366);
or U3374 (N_3374,N_592,N_1885);
nor U3375 (N_3375,N_1857,N_1465);
nand U3376 (N_3376,N_792,N_2078);
xor U3377 (N_3377,N_707,N_2085);
nor U3378 (N_3378,N_1510,N_892);
nand U3379 (N_3379,N_457,N_2403);
or U3380 (N_3380,N_1845,N_872);
and U3381 (N_3381,N_432,N_137);
or U3382 (N_3382,N_920,N_389);
or U3383 (N_3383,N_2475,N_229);
nand U3384 (N_3384,N_1354,N_2104);
nand U3385 (N_3385,N_1993,N_205);
or U3386 (N_3386,N_1839,N_461);
nand U3387 (N_3387,N_1919,N_147);
nor U3388 (N_3388,N_1613,N_836);
nor U3389 (N_3389,N_1108,N_118);
and U3390 (N_3390,N_534,N_1341);
nand U3391 (N_3391,N_2352,N_2340);
nand U3392 (N_3392,N_1178,N_54);
and U3393 (N_3393,N_1431,N_2429);
nand U3394 (N_3394,N_673,N_1040);
nand U3395 (N_3395,N_689,N_1618);
nor U3396 (N_3396,N_2367,N_60);
and U3397 (N_3397,N_1113,N_2149);
nor U3398 (N_3398,N_1288,N_1990);
or U3399 (N_3399,N_2124,N_778);
or U3400 (N_3400,N_77,N_196);
nor U3401 (N_3401,N_1093,N_474);
nand U3402 (N_3402,N_303,N_1912);
or U3403 (N_3403,N_2090,N_1701);
nor U3404 (N_3404,N_563,N_5);
and U3405 (N_3405,N_1999,N_440);
or U3406 (N_3406,N_1622,N_1283);
and U3407 (N_3407,N_942,N_1551);
or U3408 (N_3408,N_927,N_473);
or U3409 (N_3409,N_1443,N_420);
nor U3410 (N_3410,N_1339,N_366);
or U3411 (N_3411,N_1533,N_1296);
nand U3412 (N_3412,N_2471,N_1920);
nor U3413 (N_3413,N_2348,N_521);
or U3414 (N_3414,N_1582,N_2295);
and U3415 (N_3415,N_1081,N_1686);
and U3416 (N_3416,N_2401,N_441);
and U3417 (N_3417,N_2315,N_198);
and U3418 (N_3418,N_1498,N_1132);
or U3419 (N_3419,N_1396,N_2099);
nand U3420 (N_3420,N_1640,N_938);
nor U3421 (N_3421,N_2388,N_2216);
nand U3422 (N_3422,N_144,N_1074);
and U3423 (N_3423,N_561,N_2291);
nor U3424 (N_3424,N_2219,N_1889);
nand U3425 (N_3425,N_458,N_2166);
nor U3426 (N_3426,N_1983,N_1138);
nor U3427 (N_3427,N_2122,N_2379);
nor U3428 (N_3428,N_1069,N_471);
xor U3429 (N_3429,N_2160,N_2110);
nand U3430 (N_3430,N_1718,N_553);
nand U3431 (N_3431,N_1753,N_454);
nand U3432 (N_3432,N_1496,N_1979);
or U3433 (N_3433,N_1098,N_139);
and U3434 (N_3434,N_1796,N_973);
xor U3435 (N_3435,N_211,N_518);
or U3436 (N_3436,N_1089,N_1529);
nand U3437 (N_3437,N_802,N_586);
or U3438 (N_3438,N_725,N_722);
nand U3439 (N_3439,N_1293,N_1666);
nand U3440 (N_3440,N_398,N_1363);
nand U3441 (N_3441,N_2098,N_590);
nor U3442 (N_3442,N_908,N_1900);
and U3443 (N_3443,N_842,N_2056);
or U3444 (N_3444,N_1736,N_1251);
and U3445 (N_3445,N_1018,N_2051);
and U3446 (N_3446,N_721,N_1792);
nand U3447 (N_3447,N_1784,N_1754);
or U3448 (N_3448,N_2355,N_544);
and U3449 (N_3449,N_2375,N_1813);
nor U3450 (N_3450,N_1956,N_899);
and U3451 (N_3451,N_1765,N_187);
nand U3452 (N_3452,N_891,N_2058);
nand U3453 (N_3453,N_2376,N_446);
or U3454 (N_3454,N_228,N_1441);
nor U3455 (N_3455,N_1719,N_1809);
and U3456 (N_3456,N_1189,N_1381);
or U3457 (N_3457,N_1144,N_1159);
or U3458 (N_3458,N_631,N_1438);
and U3459 (N_3459,N_2001,N_1252);
and U3460 (N_3460,N_589,N_449);
nand U3461 (N_3461,N_2218,N_1654);
nand U3462 (N_3462,N_699,N_2314);
and U3463 (N_3463,N_952,N_1289);
nand U3464 (N_3464,N_1356,N_485);
nor U3465 (N_3465,N_1502,N_321);
and U3466 (N_3466,N_963,N_567);
nand U3467 (N_3467,N_1815,N_2492);
nor U3468 (N_3468,N_936,N_2476);
and U3469 (N_3469,N_1891,N_1984);
nand U3470 (N_3470,N_967,N_2195);
nand U3471 (N_3471,N_1708,N_2309);
nand U3472 (N_3472,N_956,N_99);
nor U3473 (N_3473,N_970,N_148);
or U3474 (N_3474,N_1294,N_1927);
or U3475 (N_3475,N_1541,N_376);
nand U3476 (N_3476,N_22,N_1547);
and U3477 (N_3477,N_1417,N_1921);
or U3478 (N_3478,N_1546,N_43);
nor U3479 (N_3479,N_2378,N_549);
nor U3480 (N_3480,N_537,N_665);
and U3481 (N_3481,N_848,N_193);
nor U3482 (N_3482,N_382,N_1424);
nor U3483 (N_3483,N_1049,N_184);
nand U3484 (N_3484,N_226,N_1007);
or U3485 (N_3485,N_2024,N_1882);
and U3486 (N_3486,N_2482,N_819);
nand U3487 (N_3487,N_2162,N_1080);
or U3488 (N_3488,N_1941,N_966);
and U3489 (N_3489,N_2345,N_203);
or U3490 (N_3490,N_1678,N_1142);
and U3491 (N_3491,N_2349,N_1932);
and U3492 (N_3492,N_61,N_475);
or U3493 (N_3493,N_1119,N_1707);
or U3494 (N_3494,N_435,N_285);
nor U3495 (N_3495,N_1092,N_1390);
or U3496 (N_3496,N_2229,N_328);
and U3497 (N_3497,N_2322,N_1372);
or U3498 (N_3498,N_2063,N_2080);
nor U3499 (N_3499,N_558,N_1223);
or U3500 (N_3500,N_1287,N_347);
or U3501 (N_3501,N_168,N_1875);
nand U3502 (N_3502,N_1304,N_826);
nor U3503 (N_3503,N_614,N_2236);
nand U3504 (N_3504,N_2048,N_522);
nand U3505 (N_3505,N_2086,N_1451);
and U3506 (N_3506,N_794,N_2059);
or U3507 (N_3507,N_2394,N_1866);
xnor U3508 (N_3508,N_481,N_2224);
or U3509 (N_3509,N_1131,N_1404);
and U3510 (N_3510,N_2172,N_1182);
or U3511 (N_3511,N_1395,N_136);
nand U3512 (N_3512,N_1594,N_2470);
or U3513 (N_3513,N_2126,N_864);
or U3514 (N_3514,N_655,N_1174);
nor U3515 (N_3515,N_2336,N_1833);
xnor U3516 (N_3516,N_448,N_1195);
nor U3517 (N_3517,N_580,N_630);
xor U3518 (N_3518,N_624,N_643);
or U3519 (N_3519,N_1470,N_288);
nor U3520 (N_3520,N_340,N_295);
and U3521 (N_3521,N_1148,N_1887);
nor U3522 (N_3522,N_2381,N_1014);
nand U3523 (N_3523,N_915,N_1129);
or U3524 (N_3524,N_209,N_1522);
xor U3525 (N_3525,N_427,N_2029);
or U3526 (N_3526,N_406,N_67);
nor U3527 (N_3527,N_1474,N_1858);
nor U3528 (N_3528,N_0,N_1816);
or U3529 (N_3529,N_692,N_1715);
xnor U3530 (N_3530,N_1091,N_1308);
and U3531 (N_3531,N_1970,N_519);
xnor U3532 (N_3532,N_1797,N_827);
xor U3533 (N_3533,N_642,N_1933);
and U3534 (N_3534,N_312,N_1364);
or U3535 (N_3535,N_1482,N_48);
xnor U3536 (N_3536,N_371,N_1545);
nand U3537 (N_3537,N_548,N_1051);
nand U3538 (N_3538,N_2042,N_1416);
and U3539 (N_3539,N_2030,N_1881);
or U3540 (N_3540,N_2011,N_2478);
or U3541 (N_3541,N_833,N_1632);
or U3542 (N_3542,N_323,N_1410);
and U3543 (N_3543,N_863,N_332);
nand U3544 (N_3544,N_428,N_2490);
nor U3545 (N_3545,N_2210,N_360);
nor U3546 (N_3546,N_2351,N_1278);
nor U3547 (N_3547,N_1242,N_2477);
nor U3548 (N_3548,N_292,N_2175);
or U3549 (N_3549,N_2266,N_2385);
nand U3550 (N_3550,N_2041,N_1877);
and U3551 (N_3551,N_1945,N_770);
nor U3552 (N_3552,N_240,N_1507);
nand U3553 (N_3553,N_1022,N_2448);
xor U3554 (N_3554,N_726,N_2424);
and U3555 (N_3555,N_1476,N_657);
or U3556 (N_3556,N_545,N_1783);
xnor U3557 (N_3557,N_1458,N_2447);
nor U3558 (N_3558,N_1536,N_2102);
nor U3559 (N_3559,N_738,N_1153);
or U3560 (N_3560,N_1832,N_1939);
and U3561 (N_3561,N_618,N_1644);
or U3562 (N_3562,N_250,N_1084);
and U3563 (N_3563,N_1375,N_824);
and U3564 (N_3564,N_1382,N_974);
nor U3565 (N_3565,N_369,N_90);
nand U3566 (N_3566,N_388,N_1709);
or U3567 (N_3567,N_1326,N_1627);
nor U3568 (N_3568,N_1886,N_2292);
nor U3569 (N_3569,N_2439,N_1573);
and U3570 (N_3570,N_935,N_1673);
and U3571 (N_3571,N_216,N_1383);
nor U3572 (N_3572,N_993,N_452);
or U3573 (N_3573,N_579,N_2164);
nor U3574 (N_3574,N_1169,N_24);
and U3575 (N_3575,N_469,N_1908);
nor U3576 (N_3576,N_383,N_2027);
and U3577 (N_3577,N_1179,N_644);
or U3578 (N_3578,N_1196,N_603);
or U3579 (N_3579,N_1002,N_72);
or U3580 (N_3580,N_638,N_212);
or U3581 (N_3581,N_476,N_2177);
and U3582 (N_3582,N_2153,N_1235);
nand U3583 (N_3583,N_1989,N_839);
nand U3584 (N_3584,N_913,N_1652);
nor U3585 (N_3585,N_894,N_356);
nand U3586 (N_3586,N_1374,N_1463);
or U3587 (N_3587,N_1517,N_2296);
nand U3588 (N_3588,N_1992,N_1420);
and U3589 (N_3589,N_304,N_808);
or U3590 (N_3590,N_1617,N_2275);
or U3591 (N_3591,N_1774,N_1181);
or U3592 (N_3592,N_930,N_1280);
nor U3593 (N_3593,N_2372,N_120);
nor U3594 (N_3594,N_874,N_2143);
nor U3595 (N_3595,N_1677,N_910);
and U3596 (N_3596,N_1050,N_164);
xnor U3597 (N_3597,N_2461,N_390);
and U3598 (N_3598,N_2203,N_1548);
or U3599 (N_3599,N_1281,N_595);
nand U3600 (N_3600,N_1928,N_1240);
or U3601 (N_3601,N_2339,N_1259);
or U3602 (N_3602,N_2,N_805);
nor U3603 (N_3603,N_23,N_683);
and U3604 (N_3604,N_2227,N_531);
and U3605 (N_3605,N_1017,N_608);
or U3606 (N_3606,N_990,N_902);
and U3607 (N_3607,N_1345,N_613);
and U3608 (N_3608,N_1598,N_1430);
or U3609 (N_3609,N_1799,N_2209);
or U3610 (N_3610,N_821,N_241);
nor U3611 (N_3611,N_2259,N_2136);
nand U3612 (N_3612,N_2324,N_650);
and U3613 (N_3613,N_1856,N_158);
nand U3614 (N_3614,N_1859,N_690);
or U3615 (N_3615,N_2096,N_1973);
or U3616 (N_3616,N_161,N_2425);
or U3617 (N_3617,N_1893,N_1247);
nor U3618 (N_3618,N_1425,N_1351);
or U3619 (N_3619,N_1587,N_529);
nand U3620 (N_3620,N_1096,N_682);
or U3621 (N_3621,N_686,N_675);
nor U3622 (N_3622,N_1924,N_1752);
and U3623 (N_3623,N_2263,N_1826);
and U3624 (N_3624,N_1879,N_714);
nor U3625 (N_3625,N_1649,N_617);
or U3626 (N_3626,N_831,N_301);
nor U3627 (N_3627,N_2133,N_2019);
and U3628 (N_3628,N_2146,N_2066);
and U3629 (N_3629,N_1823,N_1671);
and U3630 (N_3630,N_2485,N_259);
nand U3631 (N_3631,N_201,N_2007);
nand U3632 (N_3632,N_220,N_883);
or U3633 (N_3633,N_227,N_885);
nand U3634 (N_3634,N_68,N_1253);
or U3635 (N_3635,N_275,N_857);
and U3636 (N_3636,N_1695,N_1766);
and U3637 (N_3637,N_2049,N_1880);
and U3638 (N_3638,N_1693,N_100);
nand U3639 (N_3639,N_588,N_1631);
nand U3640 (N_3640,N_486,N_1811);
or U3641 (N_3641,N_1333,N_716);
nor U3642 (N_3642,N_594,N_2406);
nor U3643 (N_3643,N_845,N_735);
or U3644 (N_3644,N_2095,N_409);
or U3645 (N_3645,N_2062,N_2277);
nor U3646 (N_3646,N_1795,N_1000);
and U3647 (N_3647,N_8,N_135);
nand U3648 (N_3648,N_1204,N_1078);
nor U3649 (N_3649,N_926,N_344);
nor U3650 (N_3650,N_1838,N_1570);
and U3651 (N_3651,N_1066,N_1692);
nor U3652 (N_3652,N_1094,N_2305);
nor U3653 (N_3653,N_1836,N_2389);
and U3654 (N_3654,N_2399,N_988);
or U3655 (N_3655,N_444,N_1679);
and U3656 (N_3656,N_917,N_1749);
nand U3657 (N_3657,N_1362,N_447);
or U3658 (N_3658,N_1542,N_1344);
nor U3659 (N_3659,N_1802,N_18);
or U3660 (N_3660,N_2190,N_1616);
nand U3661 (N_3661,N_1295,N_733);
nor U3662 (N_3662,N_584,N_1680);
and U3663 (N_3663,N_1549,N_1694);
nor U3664 (N_3664,N_1848,N_1493);
or U3665 (N_3665,N_291,N_338);
and U3666 (N_3666,N_2067,N_1439);
nor U3667 (N_3667,N_2313,N_2108);
nand U3668 (N_3668,N_204,N_1254);
nand U3669 (N_3669,N_1514,N_2370);
nand U3670 (N_3670,N_2276,N_116);
or U3671 (N_3671,N_243,N_10);
nor U3672 (N_3672,N_791,N_2075);
and U3673 (N_3673,N_362,N_659);
or U3674 (N_3674,N_825,N_2298);
or U3675 (N_3675,N_834,N_1596);
nor U3676 (N_3676,N_65,N_253);
nor U3677 (N_3677,N_1111,N_1607);
nor U3678 (N_3678,N_2097,N_2308);
or U3679 (N_3679,N_7,N_1943);
nand U3680 (N_3680,N_1655,N_430);
nand U3681 (N_3681,N_1965,N_925);
nor U3682 (N_3682,N_2484,N_372);
nand U3683 (N_3683,N_2173,N_145);
nand U3684 (N_3684,N_2245,N_472);
and U3685 (N_3685,N_1202,N_75);
or U3686 (N_3686,N_2068,N_703);
and U3687 (N_3687,N_1662,N_2225);
or U3688 (N_3688,N_953,N_1090);
nor U3689 (N_3689,N_1423,N_97);
or U3690 (N_3690,N_765,N_479);
nor U3691 (N_3691,N_879,N_1831);
and U3692 (N_3692,N_2233,N_612);
nor U3693 (N_3693,N_1844,N_1645);
nand U3694 (N_3694,N_151,N_314);
nand U3695 (N_3695,N_1162,N_2466);
nand U3696 (N_3696,N_1316,N_1526);
and U3697 (N_3697,N_1379,N_1035);
or U3698 (N_3698,N_2335,N_335);
nand U3699 (N_3699,N_1946,N_1539);
nand U3700 (N_3700,N_57,N_2250);
nor U3701 (N_3701,N_639,N_1506);
or U3702 (N_3702,N_1385,N_1403);
nand U3703 (N_3703,N_2106,N_140);
and U3704 (N_3704,N_297,N_2456);
or U3705 (N_3705,N_654,N_342);
or U3706 (N_3706,N_181,N_1523);
and U3707 (N_3707,N_299,N_1870);
nor U3708 (N_3708,N_1818,N_768);
and U3709 (N_3709,N_1057,N_769);
or U3710 (N_3710,N_1409,N_981);
nand U3711 (N_3711,N_2303,N_2139);
nand U3712 (N_3712,N_752,N_1800);
nand U3713 (N_3713,N_1087,N_1171);
and U3714 (N_3714,N_2495,N_681);
and U3715 (N_3715,N_1601,N_2481);
and U3716 (N_3716,N_2270,N_1033);
nor U3717 (N_3717,N_1301,N_2354);
nor U3718 (N_3718,N_254,N_502);
nand U3719 (N_3719,N_615,N_621);
nand U3720 (N_3720,N_793,N_905);
or U3721 (N_3721,N_2235,N_2046);
and U3722 (N_3722,N_1290,N_702);
nand U3723 (N_3723,N_950,N_459);
nor U3724 (N_3724,N_279,N_1349);
nand U3725 (N_3725,N_1405,N_1392);
and U3726 (N_3726,N_1190,N_2260);
nand U3727 (N_3727,N_336,N_1260);
nor U3728 (N_3728,N_49,N_931);
or U3729 (N_3729,N_2020,N_785);
or U3730 (N_3730,N_419,N_1821);
nand U3731 (N_3731,N_1837,N_919);
or U3732 (N_3732,N_1329,N_719);
or U3733 (N_3733,N_1798,N_202);
or U3734 (N_3734,N_117,N_1023);
or U3735 (N_3735,N_16,N_367);
and U3736 (N_3736,N_429,N_1188);
nand U3737 (N_3737,N_1156,N_247);
and U3738 (N_3738,N_74,N_886);
nor U3739 (N_3739,N_98,N_1484);
and U3740 (N_3740,N_1599,N_564);
or U3741 (N_3741,N_96,N_1359);
nand U3742 (N_3742,N_2488,N_185);
nand U3743 (N_3743,N_1168,N_2279);
nor U3744 (N_3744,N_2268,N_1175);
and U3745 (N_3745,N_330,N_1309);
nor U3746 (N_3746,N_282,N_155);
nand U3747 (N_3747,N_1532,N_1454);
or U3748 (N_3748,N_1944,N_2359);
or U3749 (N_3749,N_1703,N_1275);
and U3750 (N_3750,N_262,N_1854);
nand U3751 (N_3751,N_887,N_826);
nand U3752 (N_3752,N_911,N_1968);
and U3753 (N_3753,N_663,N_1625);
nand U3754 (N_3754,N_261,N_981);
and U3755 (N_3755,N_1911,N_1295);
nand U3756 (N_3756,N_1557,N_1072);
or U3757 (N_3757,N_1825,N_1128);
or U3758 (N_3758,N_60,N_2304);
nor U3759 (N_3759,N_1042,N_796);
or U3760 (N_3760,N_1397,N_1811);
nand U3761 (N_3761,N_1598,N_1496);
and U3762 (N_3762,N_2437,N_1798);
nand U3763 (N_3763,N_2485,N_2477);
and U3764 (N_3764,N_480,N_352);
or U3765 (N_3765,N_897,N_692);
nand U3766 (N_3766,N_1914,N_2248);
and U3767 (N_3767,N_2076,N_2361);
and U3768 (N_3768,N_1934,N_38);
and U3769 (N_3769,N_926,N_601);
nand U3770 (N_3770,N_1902,N_752);
nand U3771 (N_3771,N_1064,N_2365);
or U3772 (N_3772,N_731,N_649);
nor U3773 (N_3773,N_515,N_274);
and U3774 (N_3774,N_1602,N_592);
nor U3775 (N_3775,N_2059,N_1393);
nand U3776 (N_3776,N_370,N_826);
xor U3777 (N_3777,N_2207,N_303);
nor U3778 (N_3778,N_2242,N_755);
and U3779 (N_3779,N_511,N_72);
and U3780 (N_3780,N_1683,N_507);
nand U3781 (N_3781,N_281,N_898);
nand U3782 (N_3782,N_1027,N_954);
nand U3783 (N_3783,N_2,N_791);
nand U3784 (N_3784,N_733,N_1183);
nand U3785 (N_3785,N_1108,N_1724);
and U3786 (N_3786,N_38,N_54);
or U3787 (N_3787,N_948,N_253);
and U3788 (N_3788,N_2000,N_1313);
nor U3789 (N_3789,N_1535,N_359);
nor U3790 (N_3790,N_1129,N_437);
nor U3791 (N_3791,N_2314,N_210);
nand U3792 (N_3792,N_746,N_697);
nand U3793 (N_3793,N_64,N_2396);
nand U3794 (N_3794,N_1276,N_291);
and U3795 (N_3795,N_438,N_337);
or U3796 (N_3796,N_34,N_1877);
nor U3797 (N_3797,N_527,N_2045);
or U3798 (N_3798,N_702,N_1849);
or U3799 (N_3799,N_1136,N_1826);
nand U3800 (N_3800,N_1043,N_303);
and U3801 (N_3801,N_997,N_1023);
nor U3802 (N_3802,N_1935,N_1406);
or U3803 (N_3803,N_469,N_588);
nand U3804 (N_3804,N_2334,N_1849);
and U3805 (N_3805,N_2455,N_1735);
nor U3806 (N_3806,N_1505,N_568);
nor U3807 (N_3807,N_2106,N_293);
nand U3808 (N_3808,N_570,N_1007);
nor U3809 (N_3809,N_237,N_2139);
nor U3810 (N_3810,N_114,N_1190);
and U3811 (N_3811,N_1563,N_1050);
nor U3812 (N_3812,N_1750,N_489);
and U3813 (N_3813,N_481,N_2386);
nor U3814 (N_3814,N_1075,N_1251);
nor U3815 (N_3815,N_1381,N_1528);
and U3816 (N_3816,N_897,N_771);
or U3817 (N_3817,N_396,N_536);
or U3818 (N_3818,N_633,N_1241);
nand U3819 (N_3819,N_2472,N_2101);
and U3820 (N_3820,N_76,N_982);
nand U3821 (N_3821,N_2224,N_274);
nand U3822 (N_3822,N_1974,N_1302);
nand U3823 (N_3823,N_1362,N_2070);
nand U3824 (N_3824,N_548,N_903);
nand U3825 (N_3825,N_248,N_2122);
and U3826 (N_3826,N_1607,N_1917);
and U3827 (N_3827,N_2105,N_2367);
and U3828 (N_3828,N_1898,N_1932);
or U3829 (N_3829,N_1911,N_1454);
nand U3830 (N_3830,N_1499,N_807);
or U3831 (N_3831,N_662,N_2212);
and U3832 (N_3832,N_2103,N_2309);
nor U3833 (N_3833,N_649,N_37);
nand U3834 (N_3834,N_2376,N_2070);
and U3835 (N_3835,N_1657,N_1429);
and U3836 (N_3836,N_249,N_1143);
and U3837 (N_3837,N_33,N_1702);
or U3838 (N_3838,N_2127,N_1573);
nand U3839 (N_3839,N_722,N_639);
nor U3840 (N_3840,N_2387,N_576);
and U3841 (N_3841,N_332,N_1805);
or U3842 (N_3842,N_1403,N_1769);
and U3843 (N_3843,N_221,N_1425);
nor U3844 (N_3844,N_958,N_644);
nand U3845 (N_3845,N_2256,N_2213);
xnor U3846 (N_3846,N_1535,N_1152);
nor U3847 (N_3847,N_2039,N_2030);
nand U3848 (N_3848,N_1191,N_540);
or U3849 (N_3849,N_830,N_948);
nor U3850 (N_3850,N_1280,N_1769);
or U3851 (N_3851,N_561,N_2035);
and U3852 (N_3852,N_2418,N_2474);
nor U3853 (N_3853,N_1520,N_474);
and U3854 (N_3854,N_365,N_1);
nand U3855 (N_3855,N_998,N_1919);
or U3856 (N_3856,N_1391,N_161);
nor U3857 (N_3857,N_2197,N_633);
or U3858 (N_3858,N_777,N_2125);
and U3859 (N_3859,N_603,N_123);
nor U3860 (N_3860,N_595,N_1128);
nand U3861 (N_3861,N_2269,N_2080);
and U3862 (N_3862,N_1845,N_2356);
nor U3863 (N_3863,N_1846,N_1977);
or U3864 (N_3864,N_1061,N_1789);
nor U3865 (N_3865,N_2304,N_2204);
nand U3866 (N_3866,N_1948,N_1553);
nand U3867 (N_3867,N_1162,N_782);
or U3868 (N_3868,N_1023,N_1689);
nor U3869 (N_3869,N_865,N_1575);
nand U3870 (N_3870,N_2123,N_1779);
or U3871 (N_3871,N_2053,N_816);
nand U3872 (N_3872,N_1212,N_286);
and U3873 (N_3873,N_295,N_424);
nor U3874 (N_3874,N_458,N_619);
nand U3875 (N_3875,N_2434,N_1965);
nand U3876 (N_3876,N_988,N_859);
and U3877 (N_3877,N_1414,N_1974);
nor U3878 (N_3878,N_1640,N_1721);
or U3879 (N_3879,N_965,N_245);
and U3880 (N_3880,N_1132,N_2192);
or U3881 (N_3881,N_367,N_214);
nor U3882 (N_3882,N_963,N_1458);
xor U3883 (N_3883,N_1553,N_278);
and U3884 (N_3884,N_371,N_397);
nor U3885 (N_3885,N_1036,N_1490);
and U3886 (N_3886,N_357,N_623);
nor U3887 (N_3887,N_1969,N_1098);
nand U3888 (N_3888,N_834,N_248);
nor U3889 (N_3889,N_2139,N_352);
and U3890 (N_3890,N_1808,N_700);
and U3891 (N_3891,N_1690,N_1642);
nor U3892 (N_3892,N_1753,N_1836);
nand U3893 (N_3893,N_1894,N_2392);
and U3894 (N_3894,N_1800,N_303);
nor U3895 (N_3895,N_1543,N_1276);
nor U3896 (N_3896,N_743,N_595);
nand U3897 (N_3897,N_1069,N_2183);
and U3898 (N_3898,N_1268,N_2136);
nor U3899 (N_3899,N_66,N_1027);
and U3900 (N_3900,N_1181,N_1304);
xnor U3901 (N_3901,N_2440,N_2401);
or U3902 (N_3902,N_905,N_1953);
xor U3903 (N_3903,N_795,N_2161);
nor U3904 (N_3904,N_946,N_1885);
or U3905 (N_3905,N_2174,N_282);
or U3906 (N_3906,N_2358,N_2054);
or U3907 (N_3907,N_548,N_1241);
nor U3908 (N_3908,N_328,N_13);
and U3909 (N_3909,N_1269,N_594);
nand U3910 (N_3910,N_1381,N_1897);
and U3911 (N_3911,N_1363,N_828);
or U3912 (N_3912,N_1817,N_2067);
and U3913 (N_3913,N_1104,N_2210);
or U3914 (N_3914,N_446,N_2419);
xor U3915 (N_3915,N_423,N_747);
xor U3916 (N_3916,N_1616,N_2408);
and U3917 (N_3917,N_7,N_493);
nand U3918 (N_3918,N_1190,N_1389);
and U3919 (N_3919,N_2458,N_1093);
and U3920 (N_3920,N_2362,N_1211);
and U3921 (N_3921,N_1763,N_839);
and U3922 (N_3922,N_1332,N_1975);
nand U3923 (N_3923,N_1418,N_2271);
or U3924 (N_3924,N_1909,N_2461);
nor U3925 (N_3925,N_2421,N_1876);
or U3926 (N_3926,N_967,N_1079);
and U3927 (N_3927,N_2000,N_108);
nor U3928 (N_3928,N_2318,N_1322);
and U3929 (N_3929,N_1529,N_645);
and U3930 (N_3930,N_1419,N_131);
or U3931 (N_3931,N_1981,N_1066);
xnor U3932 (N_3932,N_763,N_1350);
or U3933 (N_3933,N_1344,N_59);
or U3934 (N_3934,N_429,N_486);
xor U3935 (N_3935,N_480,N_385);
or U3936 (N_3936,N_635,N_631);
and U3937 (N_3937,N_2383,N_464);
nand U3938 (N_3938,N_509,N_783);
or U3939 (N_3939,N_1092,N_205);
or U3940 (N_3940,N_475,N_1257);
or U3941 (N_3941,N_19,N_2480);
and U3942 (N_3942,N_691,N_96);
and U3943 (N_3943,N_700,N_761);
or U3944 (N_3944,N_1044,N_139);
nor U3945 (N_3945,N_1993,N_1067);
nor U3946 (N_3946,N_1344,N_1838);
nor U3947 (N_3947,N_196,N_512);
nand U3948 (N_3948,N_881,N_1203);
and U3949 (N_3949,N_1421,N_879);
nand U3950 (N_3950,N_868,N_2416);
and U3951 (N_3951,N_1265,N_1588);
or U3952 (N_3952,N_462,N_1429);
and U3953 (N_3953,N_989,N_337);
nand U3954 (N_3954,N_255,N_2219);
nand U3955 (N_3955,N_1300,N_2362);
and U3956 (N_3956,N_2258,N_2121);
or U3957 (N_3957,N_2348,N_695);
nand U3958 (N_3958,N_750,N_67);
or U3959 (N_3959,N_1163,N_353);
or U3960 (N_3960,N_1720,N_93);
and U3961 (N_3961,N_1514,N_2068);
or U3962 (N_3962,N_1883,N_992);
nor U3963 (N_3963,N_2029,N_2250);
or U3964 (N_3964,N_673,N_2112);
nand U3965 (N_3965,N_506,N_571);
and U3966 (N_3966,N_867,N_2140);
or U3967 (N_3967,N_109,N_163);
nand U3968 (N_3968,N_2074,N_689);
nor U3969 (N_3969,N_914,N_1987);
nor U3970 (N_3970,N_1429,N_2296);
or U3971 (N_3971,N_1538,N_1469);
nand U3972 (N_3972,N_2151,N_1186);
nor U3973 (N_3973,N_1847,N_1809);
and U3974 (N_3974,N_391,N_483);
or U3975 (N_3975,N_1854,N_2398);
nor U3976 (N_3976,N_1235,N_548);
nand U3977 (N_3977,N_2486,N_2423);
and U3978 (N_3978,N_1515,N_1593);
nand U3979 (N_3979,N_610,N_2461);
nand U3980 (N_3980,N_1668,N_2156);
and U3981 (N_3981,N_1837,N_1627);
and U3982 (N_3982,N_1233,N_2491);
nor U3983 (N_3983,N_2193,N_2332);
or U3984 (N_3984,N_944,N_2012);
or U3985 (N_3985,N_518,N_101);
or U3986 (N_3986,N_826,N_2434);
or U3987 (N_3987,N_109,N_1105);
or U3988 (N_3988,N_153,N_1696);
or U3989 (N_3989,N_1866,N_1279);
and U3990 (N_3990,N_1365,N_1708);
and U3991 (N_3991,N_1788,N_450);
and U3992 (N_3992,N_160,N_1759);
nor U3993 (N_3993,N_1298,N_1859);
or U3994 (N_3994,N_1148,N_2333);
and U3995 (N_3995,N_1246,N_1235);
or U3996 (N_3996,N_355,N_1586);
or U3997 (N_3997,N_196,N_541);
or U3998 (N_3998,N_1681,N_1314);
or U3999 (N_3999,N_987,N_1702);
nand U4000 (N_4000,N_873,N_1974);
nor U4001 (N_4001,N_1701,N_2204);
nor U4002 (N_4002,N_1425,N_288);
or U4003 (N_4003,N_345,N_1313);
nor U4004 (N_4004,N_2095,N_1037);
nor U4005 (N_4005,N_2219,N_380);
or U4006 (N_4006,N_1852,N_1678);
nor U4007 (N_4007,N_2429,N_2473);
or U4008 (N_4008,N_850,N_1223);
nand U4009 (N_4009,N_1461,N_438);
and U4010 (N_4010,N_1823,N_1794);
and U4011 (N_4011,N_468,N_186);
nor U4012 (N_4012,N_2229,N_879);
and U4013 (N_4013,N_453,N_907);
nand U4014 (N_4014,N_1156,N_2081);
nor U4015 (N_4015,N_174,N_1241);
nor U4016 (N_4016,N_702,N_2401);
and U4017 (N_4017,N_580,N_2301);
nand U4018 (N_4018,N_1600,N_2057);
nand U4019 (N_4019,N_637,N_230);
nor U4020 (N_4020,N_1768,N_399);
or U4021 (N_4021,N_1343,N_1296);
or U4022 (N_4022,N_1441,N_757);
and U4023 (N_4023,N_23,N_1114);
or U4024 (N_4024,N_2100,N_2051);
and U4025 (N_4025,N_208,N_590);
nand U4026 (N_4026,N_330,N_308);
and U4027 (N_4027,N_1931,N_882);
or U4028 (N_4028,N_2021,N_1363);
nand U4029 (N_4029,N_422,N_1183);
and U4030 (N_4030,N_1633,N_985);
and U4031 (N_4031,N_1051,N_323);
and U4032 (N_4032,N_666,N_1761);
or U4033 (N_4033,N_724,N_2179);
or U4034 (N_4034,N_2493,N_1871);
or U4035 (N_4035,N_1212,N_1462);
and U4036 (N_4036,N_551,N_2377);
nor U4037 (N_4037,N_1739,N_201);
or U4038 (N_4038,N_1518,N_600);
and U4039 (N_4039,N_0,N_1563);
or U4040 (N_4040,N_128,N_1320);
nand U4041 (N_4041,N_724,N_90);
nand U4042 (N_4042,N_133,N_1134);
and U4043 (N_4043,N_1495,N_469);
or U4044 (N_4044,N_1900,N_1865);
nor U4045 (N_4045,N_855,N_84);
xnor U4046 (N_4046,N_663,N_738);
nor U4047 (N_4047,N_1358,N_2490);
nor U4048 (N_4048,N_1802,N_1937);
nor U4049 (N_4049,N_436,N_2300);
and U4050 (N_4050,N_402,N_801);
xnor U4051 (N_4051,N_1520,N_1407);
and U4052 (N_4052,N_523,N_662);
nand U4053 (N_4053,N_1014,N_212);
nor U4054 (N_4054,N_1056,N_1811);
and U4055 (N_4055,N_2019,N_950);
nor U4056 (N_4056,N_1276,N_1215);
or U4057 (N_4057,N_2428,N_1124);
nor U4058 (N_4058,N_311,N_2385);
and U4059 (N_4059,N_1524,N_404);
nor U4060 (N_4060,N_2432,N_226);
nor U4061 (N_4061,N_114,N_1546);
nor U4062 (N_4062,N_674,N_1382);
and U4063 (N_4063,N_2109,N_179);
and U4064 (N_4064,N_2052,N_1765);
nor U4065 (N_4065,N_2213,N_815);
and U4066 (N_4066,N_654,N_1412);
xnor U4067 (N_4067,N_1202,N_2037);
or U4068 (N_4068,N_448,N_2447);
and U4069 (N_4069,N_1809,N_2484);
or U4070 (N_4070,N_2120,N_2231);
and U4071 (N_4071,N_38,N_1824);
nand U4072 (N_4072,N_109,N_1998);
nor U4073 (N_4073,N_1051,N_1022);
nand U4074 (N_4074,N_470,N_624);
xor U4075 (N_4075,N_1246,N_2489);
or U4076 (N_4076,N_264,N_223);
nand U4077 (N_4077,N_519,N_1071);
and U4078 (N_4078,N_2173,N_128);
or U4079 (N_4079,N_76,N_1243);
nand U4080 (N_4080,N_2390,N_2427);
nor U4081 (N_4081,N_1941,N_2094);
or U4082 (N_4082,N_479,N_1881);
nor U4083 (N_4083,N_1373,N_1493);
nor U4084 (N_4084,N_2283,N_2227);
or U4085 (N_4085,N_1812,N_917);
and U4086 (N_4086,N_349,N_2496);
nor U4087 (N_4087,N_1141,N_79);
nor U4088 (N_4088,N_953,N_1644);
nand U4089 (N_4089,N_674,N_489);
nor U4090 (N_4090,N_1791,N_1900);
nand U4091 (N_4091,N_919,N_1889);
and U4092 (N_4092,N_2101,N_371);
nand U4093 (N_4093,N_727,N_1859);
and U4094 (N_4094,N_1375,N_1593);
xnor U4095 (N_4095,N_1619,N_268);
nor U4096 (N_4096,N_2437,N_625);
and U4097 (N_4097,N_496,N_1068);
and U4098 (N_4098,N_873,N_1507);
nand U4099 (N_4099,N_486,N_1838);
xor U4100 (N_4100,N_2062,N_417);
nor U4101 (N_4101,N_2306,N_1808);
nor U4102 (N_4102,N_1016,N_1911);
nand U4103 (N_4103,N_2327,N_46);
nand U4104 (N_4104,N_72,N_1092);
or U4105 (N_4105,N_1447,N_585);
and U4106 (N_4106,N_323,N_1774);
and U4107 (N_4107,N_1343,N_2297);
or U4108 (N_4108,N_1615,N_1704);
and U4109 (N_4109,N_833,N_1787);
and U4110 (N_4110,N_1353,N_2162);
and U4111 (N_4111,N_349,N_146);
nor U4112 (N_4112,N_1287,N_345);
nand U4113 (N_4113,N_607,N_1193);
nor U4114 (N_4114,N_352,N_2085);
or U4115 (N_4115,N_1183,N_352);
or U4116 (N_4116,N_1048,N_1547);
and U4117 (N_4117,N_705,N_1211);
nand U4118 (N_4118,N_1536,N_1508);
and U4119 (N_4119,N_875,N_2100);
or U4120 (N_4120,N_1777,N_477);
or U4121 (N_4121,N_1797,N_184);
nand U4122 (N_4122,N_2089,N_1860);
xor U4123 (N_4123,N_1248,N_1226);
or U4124 (N_4124,N_2267,N_1493);
and U4125 (N_4125,N_2021,N_1762);
and U4126 (N_4126,N_2352,N_495);
nand U4127 (N_4127,N_1297,N_120);
and U4128 (N_4128,N_2453,N_751);
nor U4129 (N_4129,N_501,N_1876);
or U4130 (N_4130,N_2319,N_2487);
or U4131 (N_4131,N_862,N_1725);
xnor U4132 (N_4132,N_2289,N_2279);
and U4133 (N_4133,N_1804,N_1524);
and U4134 (N_4134,N_2382,N_1382);
and U4135 (N_4135,N_1468,N_780);
and U4136 (N_4136,N_594,N_226);
nor U4137 (N_4137,N_1110,N_1414);
and U4138 (N_4138,N_303,N_111);
xnor U4139 (N_4139,N_1740,N_1297);
and U4140 (N_4140,N_2176,N_2380);
or U4141 (N_4141,N_2408,N_2216);
nor U4142 (N_4142,N_136,N_41);
and U4143 (N_4143,N_193,N_710);
nand U4144 (N_4144,N_410,N_1795);
nor U4145 (N_4145,N_1513,N_1488);
nand U4146 (N_4146,N_1207,N_896);
nor U4147 (N_4147,N_1271,N_1678);
and U4148 (N_4148,N_1157,N_173);
nand U4149 (N_4149,N_572,N_120);
or U4150 (N_4150,N_45,N_525);
nand U4151 (N_4151,N_1013,N_1505);
or U4152 (N_4152,N_1030,N_258);
nand U4153 (N_4153,N_1550,N_1570);
and U4154 (N_4154,N_1264,N_133);
and U4155 (N_4155,N_404,N_546);
nor U4156 (N_4156,N_469,N_2429);
or U4157 (N_4157,N_219,N_1142);
nor U4158 (N_4158,N_2294,N_1042);
and U4159 (N_4159,N_932,N_290);
nand U4160 (N_4160,N_576,N_1760);
or U4161 (N_4161,N_140,N_796);
xnor U4162 (N_4162,N_985,N_459);
nand U4163 (N_4163,N_588,N_1184);
or U4164 (N_4164,N_126,N_2393);
and U4165 (N_4165,N_1121,N_690);
nand U4166 (N_4166,N_1564,N_802);
nor U4167 (N_4167,N_1106,N_820);
or U4168 (N_4168,N_1016,N_931);
xnor U4169 (N_4169,N_285,N_778);
nor U4170 (N_4170,N_505,N_968);
nand U4171 (N_4171,N_2486,N_1084);
or U4172 (N_4172,N_202,N_455);
nand U4173 (N_4173,N_445,N_1152);
nand U4174 (N_4174,N_2181,N_527);
nor U4175 (N_4175,N_2429,N_2193);
nand U4176 (N_4176,N_1073,N_8);
and U4177 (N_4177,N_31,N_148);
and U4178 (N_4178,N_339,N_962);
nor U4179 (N_4179,N_832,N_496);
nor U4180 (N_4180,N_1775,N_480);
and U4181 (N_4181,N_2132,N_348);
or U4182 (N_4182,N_147,N_907);
nand U4183 (N_4183,N_448,N_423);
nor U4184 (N_4184,N_1119,N_2261);
or U4185 (N_4185,N_557,N_890);
nand U4186 (N_4186,N_1279,N_1285);
or U4187 (N_4187,N_89,N_1248);
nor U4188 (N_4188,N_1534,N_2259);
and U4189 (N_4189,N_1238,N_167);
nand U4190 (N_4190,N_1381,N_2201);
or U4191 (N_4191,N_532,N_1645);
or U4192 (N_4192,N_377,N_1632);
or U4193 (N_4193,N_135,N_65);
or U4194 (N_4194,N_313,N_463);
nor U4195 (N_4195,N_767,N_1723);
nor U4196 (N_4196,N_1965,N_1200);
nor U4197 (N_4197,N_701,N_2182);
nand U4198 (N_4198,N_1884,N_1473);
and U4199 (N_4199,N_725,N_2215);
or U4200 (N_4200,N_1510,N_924);
or U4201 (N_4201,N_1464,N_482);
xnor U4202 (N_4202,N_1950,N_2048);
or U4203 (N_4203,N_1898,N_62);
nor U4204 (N_4204,N_94,N_1132);
or U4205 (N_4205,N_542,N_1927);
or U4206 (N_4206,N_1662,N_1763);
or U4207 (N_4207,N_510,N_962);
nor U4208 (N_4208,N_342,N_1328);
or U4209 (N_4209,N_1849,N_2312);
and U4210 (N_4210,N_2206,N_128);
nand U4211 (N_4211,N_1759,N_820);
nor U4212 (N_4212,N_1580,N_2187);
and U4213 (N_4213,N_1135,N_759);
or U4214 (N_4214,N_1303,N_714);
or U4215 (N_4215,N_2424,N_2166);
and U4216 (N_4216,N_2023,N_995);
and U4217 (N_4217,N_369,N_1323);
nand U4218 (N_4218,N_275,N_441);
nand U4219 (N_4219,N_331,N_230);
nand U4220 (N_4220,N_1295,N_2094);
nand U4221 (N_4221,N_1368,N_2488);
and U4222 (N_4222,N_921,N_1424);
or U4223 (N_4223,N_2379,N_378);
and U4224 (N_4224,N_1933,N_386);
xnor U4225 (N_4225,N_1305,N_1222);
and U4226 (N_4226,N_1743,N_191);
xnor U4227 (N_4227,N_2245,N_2449);
nand U4228 (N_4228,N_150,N_2131);
nor U4229 (N_4229,N_2052,N_1357);
nand U4230 (N_4230,N_2014,N_1857);
or U4231 (N_4231,N_1053,N_2373);
nor U4232 (N_4232,N_484,N_2095);
nor U4233 (N_4233,N_639,N_1092);
or U4234 (N_4234,N_360,N_1702);
nand U4235 (N_4235,N_2451,N_979);
nor U4236 (N_4236,N_1849,N_239);
and U4237 (N_4237,N_1165,N_2462);
and U4238 (N_4238,N_81,N_1148);
or U4239 (N_4239,N_209,N_2175);
and U4240 (N_4240,N_2146,N_2249);
or U4241 (N_4241,N_1417,N_809);
nand U4242 (N_4242,N_1499,N_2379);
nor U4243 (N_4243,N_2184,N_109);
and U4244 (N_4244,N_399,N_2085);
or U4245 (N_4245,N_1083,N_740);
nand U4246 (N_4246,N_2124,N_543);
and U4247 (N_4247,N_136,N_1371);
nor U4248 (N_4248,N_1109,N_410);
and U4249 (N_4249,N_1038,N_1234);
and U4250 (N_4250,N_2278,N_356);
or U4251 (N_4251,N_1112,N_2350);
and U4252 (N_4252,N_2312,N_1002);
nand U4253 (N_4253,N_1256,N_1400);
or U4254 (N_4254,N_2146,N_1053);
nor U4255 (N_4255,N_1779,N_1872);
nand U4256 (N_4256,N_1861,N_1137);
or U4257 (N_4257,N_2292,N_1540);
nor U4258 (N_4258,N_1822,N_1901);
and U4259 (N_4259,N_1728,N_1732);
or U4260 (N_4260,N_19,N_1373);
or U4261 (N_4261,N_1588,N_1522);
nor U4262 (N_4262,N_365,N_203);
nor U4263 (N_4263,N_726,N_994);
nand U4264 (N_4264,N_1013,N_428);
nor U4265 (N_4265,N_1521,N_1473);
nand U4266 (N_4266,N_2309,N_1713);
and U4267 (N_4267,N_800,N_437);
and U4268 (N_4268,N_2168,N_322);
nand U4269 (N_4269,N_1314,N_2036);
or U4270 (N_4270,N_1198,N_682);
nor U4271 (N_4271,N_43,N_1249);
and U4272 (N_4272,N_1191,N_970);
or U4273 (N_4273,N_703,N_1762);
nand U4274 (N_4274,N_2111,N_1197);
nor U4275 (N_4275,N_1052,N_853);
or U4276 (N_4276,N_1760,N_1203);
nor U4277 (N_4277,N_1609,N_994);
nand U4278 (N_4278,N_304,N_1048);
nand U4279 (N_4279,N_649,N_986);
or U4280 (N_4280,N_954,N_1142);
and U4281 (N_4281,N_1008,N_2374);
nor U4282 (N_4282,N_138,N_1632);
nand U4283 (N_4283,N_1813,N_1374);
and U4284 (N_4284,N_1081,N_1492);
and U4285 (N_4285,N_678,N_1644);
or U4286 (N_4286,N_930,N_570);
and U4287 (N_4287,N_2263,N_1331);
or U4288 (N_4288,N_2384,N_2377);
nor U4289 (N_4289,N_386,N_2358);
and U4290 (N_4290,N_1389,N_612);
or U4291 (N_4291,N_1873,N_1290);
nor U4292 (N_4292,N_1833,N_2224);
or U4293 (N_4293,N_1089,N_1677);
or U4294 (N_4294,N_1818,N_711);
nand U4295 (N_4295,N_2399,N_1253);
xnor U4296 (N_4296,N_1831,N_1209);
nand U4297 (N_4297,N_1709,N_636);
and U4298 (N_4298,N_2423,N_1383);
xnor U4299 (N_4299,N_557,N_1058);
and U4300 (N_4300,N_321,N_311);
or U4301 (N_4301,N_1604,N_158);
and U4302 (N_4302,N_1941,N_235);
and U4303 (N_4303,N_933,N_1096);
or U4304 (N_4304,N_1596,N_998);
and U4305 (N_4305,N_1320,N_2403);
nand U4306 (N_4306,N_187,N_1997);
and U4307 (N_4307,N_1639,N_1155);
and U4308 (N_4308,N_152,N_1892);
nor U4309 (N_4309,N_531,N_1777);
xnor U4310 (N_4310,N_1665,N_1849);
nand U4311 (N_4311,N_1397,N_76);
and U4312 (N_4312,N_613,N_1020);
and U4313 (N_4313,N_41,N_1505);
or U4314 (N_4314,N_2179,N_1436);
nand U4315 (N_4315,N_984,N_2106);
nor U4316 (N_4316,N_923,N_2300);
nor U4317 (N_4317,N_1067,N_1550);
and U4318 (N_4318,N_1191,N_1047);
nand U4319 (N_4319,N_153,N_1771);
nor U4320 (N_4320,N_991,N_1826);
nor U4321 (N_4321,N_2389,N_2053);
nand U4322 (N_4322,N_1101,N_2383);
nand U4323 (N_4323,N_1157,N_1521);
nor U4324 (N_4324,N_2070,N_24);
or U4325 (N_4325,N_1011,N_253);
or U4326 (N_4326,N_2489,N_99);
nor U4327 (N_4327,N_1144,N_1616);
and U4328 (N_4328,N_1318,N_115);
or U4329 (N_4329,N_2369,N_2002);
nor U4330 (N_4330,N_493,N_1044);
nor U4331 (N_4331,N_883,N_218);
nand U4332 (N_4332,N_232,N_890);
nor U4333 (N_4333,N_1912,N_926);
nand U4334 (N_4334,N_2398,N_788);
or U4335 (N_4335,N_1738,N_2390);
or U4336 (N_4336,N_1168,N_1680);
or U4337 (N_4337,N_528,N_535);
nand U4338 (N_4338,N_1233,N_1073);
nand U4339 (N_4339,N_1564,N_1504);
nor U4340 (N_4340,N_1157,N_755);
and U4341 (N_4341,N_994,N_157);
nor U4342 (N_4342,N_2040,N_871);
and U4343 (N_4343,N_740,N_1579);
nor U4344 (N_4344,N_1607,N_1894);
or U4345 (N_4345,N_704,N_591);
nor U4346 (N_4346,N_654,N_2053);
nor U4347 (N_4347,N_435,N_431);
nand U4348 (N_4348,N_1624,N_1338);
nor U4349 (N_4349,N_526,N_1102);
nand U4350 (N_4350,N_1605,N_2234);
nand U4351 (N_4351,N_2246,N_1008);
nor U4352 (N_4352,N_939,N_167);
and U4353 (N_4353,N_425,N_695);
nor U4354 (N_4354,N_2448,N_254);
nor U4355 (N_4355,N_1342,N_405);
nor U4356 (N_4356,N_458,N_2474);
or U4357 (N_4357,N_1338,N_1431);
nand U4358 (N_4358,N_2162,N_1859);
nor U4359 (N_4359,N_2121,N_2110);
and U4360 (N_4360,N_2335,N_959);
nor U4361 (N_4361,N_344,N_1961);
or U4362 (N_4362,N_1562,N_1090);
nor U4363 (N_4363,N_1369,N_2075);
nor U4364 (N_4364,N_2110,N_2292);
nand U4365 (N_4365,N_1031,N_2426);
or U4366 (N_4366,N_2463,N_1341);
nor U4367 (N_4367,N_2397,N_793);
or U4368 (N_4368,N_2250,N_1968);
nand U4369 (N_4369,N_1130,N_1506);
or U4370 (N_4370,N_2209,N_1722);
or U4371 (N_4371,N_2362,N_262);
and U4372 (N_4372,N_304,N_1695);
nand U4373 (N_4373,N_2280,N_1216);
nand U4374 (N_4374,N_1862,N_160);
nor U4375 (N_4375,N_2078,N_2335);
or U4376 (N_4376,N_807,N_1217);
xor U4377 (N_4377,N_874,N_903);
nor U4378 (N_4378,N_2021,N_2156);
or U4379 (N_4379,N_2341,N_302);
and U4380 (N_4380,N_402,N_341);
nand U4381 (N_4381,N_743,N_1102);
and U4382 (N_4382,N_804,N_1050);
nand U4383 (N_4383,N_820,N_1601);
nor U4384 (N_4384,N_1310,N_2017);
or U4385 (N_4385,N_802,N_284);
or U4386 (N_4386,N_1197,N_540);
and U4387 (N_4387,N_1609,N_1718);
or U4388 (N_4388,N_556,N_2023);
nand U4389 (N_4389,N_627,N_688);
or U4390 (N_4390,N_1253,N_1572);
or U4391 (N_4391,N_963,N_1813);
and U4392 (N_4392,N_2482,N_2289);
or U4393 (N_4393,N_536,N_680);
or U4394 (N_4394,N_1456,N_448);
nor U4395 (N_4395,N_1509,N_2126);
nor U4396 (N_4396,N_786,N_2358);
nor U4397 (N_4397,N_14,N_735);
or U4398 (N_4398,N_50,N_90);
nand U4399 (N_4399,N_1297,N_1239);
nand U4400 (N_4400,N_1361,N_520);
nand U4401 (N_4401,N_1602,N_2322);
xor U4402 (N_4402,N_1223,N_1696);
nor U4403 (N_4403,N_2173,N_1438);
nor U4404 (N_4404,N_699,N_2324);
or U4405 (N_4405,N_2122,N_1205);
nor U4406 (N_4406,N_2039,N_499);
nor U4407 (N_4407,N_1847,N_1364);
or U4408 (N_4408,N_1679,N_2072);
and U4409 (N_4409,N_1213,N_2411);
or U4410 (N_4410,N_2000,N_2060);
nor U4411 (N_4411,N_36,N_2234);
or U4412 (N_4412,N_1103,N_2310);
and U4413 (N_4413,N_2094,N_626);
nand U4414 (N_4414,N_911,N_2150);
nand U4415 (N_4415,N_2401,N_630);
or U4416 (N_4416,N_352,N_476);
or U4417 (N_4417,N_784,N_2353);
or U4418 (N_4418,N_2381,N_2049);
nor U4419 (N_4419,N_240,N_7);
nor U4420 (N_4420,N_2473,N_993);
or U4421 (N_4421,N_1420,N_1516);
and U4422 (N_4422,N_2467,N_1841);
or U4423 (N_4423,N_782,N_2354);
and U4424 (N_4424,N_372,N_1737);
xnor U4425 (N_4425,N_1124,N_1818);
or U4426 (N_4426,N_2393,N_933);
or U4427 (N_4427,N_1993,N_750);
and U4428 (N_4428,N_1436,N_1983);
nand U4429 (N_4429,N_598,N_2461);
and U4430 (N_4430,N_1168,N_536);
or U4431 (N_4431,N_117,N_80);
and U4432 (N_4432,N_2273,N_1689);
xnor U4433 (N_4433,N_1671,N_1494);
and U4434 (N_4434,N_1097,N_1664);
and U4435 (N_4435,N_1049,N_2067);
xnor U4436 (N_4436,N_1255,N_1963);
or U4437 (N_4437,N_1488,N_2246);
nand U4438 (N_4438,N_1794,N_1571);
nor U4439 (N_4439,N_892,N_2101);
nor U4440 (N_4440,N_2171,N_297);
and U4441 (N_4441,N_2039,N_1758);
and U4442 (N_4442,N_2472,N_834);
nor U4443 (N_4443,N_1901,N_894);
and U4444 (N_4444,N_1926,N_1883);
and U4445 (N_4445,N_1232,N_236);
or U4446 (N_4446,N_2073,N_1448);
and U4447 (N_4447,N_2039,N_1676);
nand U4448 (N_4448,N_1225,N_1937);
or U4449 (N_4449,N_526,N_1126);
nor U4450 (N_4450,N_1528,N_1997);
and U4451 (N_4451,N_156,N_603);
nor U4452 (N_4452,N_2281,N_60);
or U4453 (N_4453,N_933,N_1431);
or U4454 (N_4454,N_2399,N_285);
and U4455 (N_4455,N_1221,N_595);
or U4456 (N_4456,N_316,N_1579);
and U4457 (N_4457,N_1936,N_1252);
and U4458 (N_4458,N_2015,N_1940);
and U4459 (N_4459,N_1565,N_764);
xor U4460 (N_4460,N_902,N_772);
and U4461 (N_4461,N_1192,N_1365);
nor U4462 (N_4462,N_1851,N_1698);
nand U4463 (N_4463,N_1339,N_945);
nor U4464 (N_4464,N_1797,N_2399);
xor U4465 (N_4465,N_1415,N_1108);
nor U4466 (N_4466,N_1048,N_754);
and U4467 (N_4467,N_2472,N_727);
or U4468 (N_4468,N_1002,N_2408);
nor U4469 (N_4469,N_255,N_1040);
nand U4470 (N_4470,N_2059,N_1368);
nand U4471 (N_4471,N_820,N_984);
and U4472 (N_4472,N_557,N_2234);
nor U4473 (N_4473,N_638,N_421);
and U4474 (N_4474,N_1402,N_886);
and U4475 (N_4475,N_694,N_1981);
and U4476 (N_4476,N_214,N_232);
nor U4477 (N_4477,N_819,N_2232);
nand U4478 (N_4478,N_890,N_2317);
or U4479 (N_4479,N_1807,N_283);
or U4480 (N_4480,N_2489,N_2165);
and U4481 (N_4481,N_2106,N_292);
and U4482 (N_4482,N_615,N_2056);
nor U4483 (N_4483,N_1623,N_2328);
nor U4484 (N_4484,N_2327,N_446);
and U4485 (N_4485,N_588,N_2355);
nand U4486 (N_4486,N_1495,N_955);
or U4487 (N_4487,N_2436,N_99);
nor U4488 (N_4488,N_871,N_1118);
and U4489 (N_4489,N_2471,N_2447);
and U4490 (N_4490,N_598,N_1892);
or U4491 (N_4491,N_1135,N_2275);
nand U4492 (N_4492,N_608,N_1544);
and U4493 (N_4493,N_1688,N_501);
or U4494 (N_4494,N_0,N_1231);
or U4495 (N_4495,N_320,N_1935);
or U4496 (N_4496,N_710,N_335);
and U4497 (N_4497,N_1142,N_89);
nor U4498 (N_4498,N_170,N_2412);
nand U4499 (N_4499,N_138,N_1333);
nand U4500 (N_4500,N_939,N_2204);
nor U4501 (N_4501,N_2424,N_298);
or U4502 (N_4502,N_398,N_765);
or U4503 (N_4503,N_2415,N_2306);
nor U4504 (N_4504,N_1811,N_1526);
or U4505 (N_4505,N_499,N_568);
and U4506 (N_4506,N_2082,N_1314);
or U4507 (N_4507,N_2482,N_1338);
xor U4508 (N_4508,N_1265,N_1116);
nand U4509 (N_4509,N_583,N_128);
nand U4510 (N_4510,N_1788,N_1904);
nor U4511 (N_4511,N_1668,N_370);
nand U4512 (N_4512,N_489,N_1369);
or U4513 (N_4513,N_378,N_6);
and U4514 (N_4514,N_1675,N_1439);
nand U4515 (N_4515,N_2222,N_96);
or U4516 (N_4516,N_2038,N_1683);
and U4517 (N_4517,N_2205,N_2211);
or U4518 (N_4518,N_1269,N_1130);
and U4519 (N_4519,N_1391,N_1009);
or U4520 (N_4520,N_2389,N_1746);
and U4521 (N_4521,N_2246,N_1961);
nand U4522 (N_4522,N_1796,N_318);
nand U4523 (N_4523,N_1486,N_2413);
or U4524 (N_4524,N_509,N_2149);
or U4525 (N_4525,N_1570,N_82);
nor U4526 (N_4526,N_2352,N_656);
nor U4527 (N_4527,N_1877,N_24);
or U4528 (N_4528,N_1935,N_2240);
nor U4529 (N_4529,N_947,N_779);
and U4530 (N_4530,N_2017,N_1613);
or U4531 (N_4531,N_1922,N_2293);
or U4532 (N_4532,N_660,N_1456);
or U4533 (N_4533,N_296,N_367);
nor U4534 (N_4534,N_563,N_98);
nor U4535 (N_4535,N_1486,N_2084);
or U4536 (N_4536,N_2045,N_712);
or U4537 (N_4537,N_497,N_1671);
nand U4538 (N_4538,N_1369,N_871);
nor U4539 (N_4539,N_2192,N_379);
nand U4540 (N_4540,N_2244,N_716);
nor U4541 (N_4541,N_1252,N_1771);
nor U4542 (N_4542,N_1527,N_2410);
nor U4543 (N_4543,N_863,N_975);
nand U4544 (N_4544,N_358,N_1693);
or U4545 (N_4545,N_2446,N_430);
nor U4546 (N_4546,N_2386,N_1820);
and U4547 (N_4547,N_2253,N_482);
or U4548 (N_4548,N_1549,N_234);
or U4549 (N_4549,N_701,N_426);
nor U4550 (N_4550,N_399,N_1461);
and U4551 (N_4551,N_1933,N_1764);
and U4552 (N_4552,N_1918,N_1604);
and U4553 (N_4553,N_507,N_270);
or U4554 (N_4554,N_929,N_1393);
or U4555 (N_4555,N_1822,N_708);
nand U4556 (N_4556,N_2362,N_382);
and U4557 (N_4557,N_1115,N_996);
and U4558 (N_4558,N_353,N_2319);
or U4559 (N_4559,N_622,N_1372);
and U4560 (N_4560,N_1793,N_1247);
nor U4561 (N_4561,N_214,N_633);
or U4562 (N_4562,N_2277,N_2182);
and U4563 (N_4563,N_972,N_794);
nor U4564 (N_4564,N_1844,N_1410);
and U4565 (N_4565,N_1471,N_743);
or U4566 (N_4566,N_2011,N_945);
and U4567 (N_4567,N_2211,N_740);
or U4568 (N_4568,N_1576,N_474);
and U4569 (N_4569,N_36,N_1820);
nand U4570 (N_4570,N_2194,N_2303);
and U4571 (N_4571,N_333,N_1172);
or U4572 (N_4572,N_240,N_1377);
nand U4573 (N_4573,N_1787,N_1018);
nor U4574 (N_4574,N_761,N_1520);
nand U4575 (N_4575,N_2334,N_997);
and U4576 (N_4576,N_1307,N_1844);
or U4577 (N_4577,N_1529,N_1534);
nor U4578 (N_4578,N_440,N_817);
and U4579 (N_4579,N_503,N_604);
nor U4580 (N_4580,N_200,N_1070);
nand U4581 (N_4581,N_214,N_412);
and U4582 (N_4582,N_1337,N_524);
or U4583 (N_4583,N_211,N_1853);
and U4584 (N_4584,N_1366,N_681);
nand U4585 (N_4585,N_588,N_335);
nor U4586 (N_4586,N_2079,N_1643);
or U4587 (N_4587,N_2150,N_364);
nor U4588 (N_4588,N_1465,N_1582);
or U4589 (N_4589,N_1832,N_2463);
and U4590 (N_4590,N_49,N_820);
or U4591 (N_4591,N_397,N_1814);
nor U4592 (N_4592,N_867,N_1076);
nand U4593 (N_4593,N_917,N_1483);
and U4594 (N_4594,N_842,N_2103);
and U4595 (N_4595,N_442,N_629);
and U4596 (N_4596,N_638,N_957);
or U4597 (N_4597,N_919,N_1332);
nor U4598 (N_4598,N_1868,N_1396);
or U4599 (N_4599,N_1919,N_183);
nor U4600 (N_4600,N_2004,N_1667);
nand U4601 (N_4601,N_1931,N_148);
nor U4602 (N_4602,N_197,N_484);
nor U4603 (N_4603,N_1274,N_1710);
nor U4604 (N_4604,N_809,N_1375);
or U4605 (N_4605,N_1683,N_1658);
or U4606 (N_4606,N_1677,N_894);
and U4607 (N_4607,N_858,N_1009);
xnor U4608 (N_4608,N_967,N_438);
and U4609 (N_4609,N_648,N_765);
or U4610 (N_4610,N_482,N_1249);
nor U4611 (N_4611,N_48,N_214);
and U4612 (N_4612,N_2431,N_2045);
and U4613 (N_4613,N_1158,N_202);
nor U4614 (N_4614,N_2317,N_888);
and U4615 (N_4615,N_467,N_2210);
or U4616 (N_4616,N_2145,N_2349);
nand U4617 (N_4617,N_2453,N_920);
nand U4618 (N_4618,N_144,N_1506);
and U4619 (N_4619,N_1340,N_677);
nor U4620 (N_4620,N_1284,N_939);
nand U4621 (N_4621,N_216,N_1252);
and U4622 (N_4622,N_2462,N_2227);
nor U4623 (N_4623,N_2101,N_1280);
or U4624 (N_4624,N_454,N_2272);
nor U4625 (N_4625,N_1688,N_2032);
nand U4626 (N_4626,N_865,N_2377);
nor U4627 (N_4627,N_317,N_1722);
and U4628 (N_4628,N_2013,N_1222);
xor U4629 (N_4629,N_2135,N_1084);
or U4630 (N_4630,N_2342,N_9);
nor U4631 (N_4631,N_677,N_974);
nand U4632 (N_4632,N_1717,N_2189);
or U4633 (N_4633,N_1306,N_1276);
nor U4634 (N_4634,N_869,N_1495);
nor U4635 (N_4635,N_1681,N_1634);
nor U4636 (N_4636,N_625,N_1111);
or U4637 (N_4637,N_751,N_2126);
nand U4638 (N_4638,N_676,N_1908);
or U4639 (N_4639,N_2094,N_1060);
or U4640 (N_4640,N_374,N_2334);
nand U4641 (N_4641,N_847,N_1659);
nand U4642 (N_4642,N_243,N_1309);
or U4643 (N_4643,N_506,N_86);
or U4644 (N_4644,N_448,N_1282);
nand U4645 (N_4645,N_2323,N_1880);
xnor U4646 (N_4646,N_1430,N_1588);
or U4647 (N_4647,N_1771,N_369);
nor U4648 (N_4648,N_2485,N_1909);
or U4649 (N_4649,N_1564,N_136);
and U4650 (N_4650,N_1005,N_534);
or U4651 (N_4651,N_365,N_568);
or U4652 (N_4652,N_152,N_900);
or U4653 (N_4653,N_1859,N_642);
and U4654 (N_4654,N_84,N_1828);
and U4655 (N_4655,N_2484,N_1313);
nor U4656 (N_4656,N_599,N_1332);
or U4657 (N_4657,N_1278,N_1135);
or U4658 (N_4658,N_671,N_1209);
and U4659 (N_4659,N_903,N_1771);
nor U4660 (N_4660,N_2318,N_950);
nor U4661 (N_4661,N_1779,N_2434);
nand U4662 (N_4662,N_2086,N_699);
xnor U4663 (N_4663,N_1231,N_876);
nor U4664 (N_4664,N_1606,N_431);
and U4665 (N_4665,N_130,N_1996);
nand U4666 (N_4666,N_1018,N_2480);
nand U4667 (N_4667,N_1232,N_1603);
or U4668 (N_4668,N_705,N_2252);
nor U4669 (N_4669,N_1782,N_488);
nor U4670 (N_4670,N_1660,N_856);
or U4671 (N_4671,N_1596,N_508);
nor U4672 (N_4672,N_806,N_1044);
nor U4673 (N_4673,N_866,N_434);
and U4674 (N_4674,N_1023,N_1623);
nor U4675 (N_4675,N_227,N_1515);
or U4676 (N_4676,N_2236,N_1090);
nand U4677 (N_4677,N_1653,N_2305);
nand U4678 (N_4678,N_1826,N_1852);
or U4679 (N_4679,N_1986,N_551);
or U4680 (N_4680,N_2420,N_653);
nor U4681 (N_4681,N_415,N_2353);
nor U4682 (N_4682,N_503,N_84);
nor U4683 (N_4683,N_1394,N_320);
or U4684 (N_4684,N_1432,N_2396);
and U4685 (N_4685,N_2395,N_1319);
nand U4686 (N_4686,N_450,N_353);
or U4687 (N_4687,N_1799,N_1045);
xnor U4688 (N_4688,N_1353,N_1707);
nor U4689 (N_4689,N_751,N_1143);
nand U4690 (N_4690,N_924,N_371);
nand U4691 (N_4691,N_2326,N_1016);
nor U4692 (N_4692,N_88,N_1665);
and U4693 (N_4693,N_267,N_1216);
nand U4694 (N_4694,N_1942,N_1228);
nand U4695 (N_4695,N_1304,N_1349);
and U4696 (N_4696,N_1222,N_356);
xor U4697 (N_4697,N_184,N_6);
or U4698 (N_4698,N_548,N_2429);
nor U4699 (N_4699,N_244,N_901);
nand U4700 (N_4700,N_1529,N_1614);
xor U4701 (N_4701,N_1581,N_1499);
xor U4702 (N_4702,N_1161,N_1157);
or U4703 (N_4703,N_803,N_1176);
nand U4704 (N_4704,N_78,N_2050);
or U4705 (N_4705,N_1348,N_2244);
nand U4706 (N_4706,N_1943,N_369);
and U4707 (N_4707,N_623,N_278);
nor U4708 (N_4708,N_914,N_1167);
or U4709 (N_4709,N_199,N_885);
and U4710 (N_4710,N_1079,N_722);
and U4711 (N_4711,N_2143,N_1070);
nor U4712 (N_4712,N_2405,N_2352);
nor U4713 (N_4713,N_1591,N_1131);
or U4714 (N_4714,N_2382,N_1978);
or U4715 (N_4715,N_1146,N_1085);
nand U4716 (N_4716,N_681,N_929);
nor U4717 (N_4717,N_590,N_2418);
and U4718 (N_4718,N_1568,N_164);
nor U4719 (N_4719,N_309,N_816);
or U4720 (N_4720,N_1339,N_661);
nor U4721 (N_4721,N_2455,N_1394);
nand U4722 (N_4722,N_2362,N_820);
nand U4723 (N_4723,N_1971,N_915);
nand U4724 (N_4724,N_2136,N_377);
nand U4725 (N_4725,N_2066,N_376);
nor U4726 (N_4726,N_2417,N_1359);
nand U4727 (N_4727,N_1458,N_1136);
nor U4728 (N_4728,N_2274,N_1381);
and U4729 (N_4729,N_485,N_900);
nand U4730 (N_4730,N_1970,N_2462);
or U4731 (N_4731,N_443,N_2202);
or U4732 (N_4732,N_2352,N_1570);
and U4733 (N_4733,N_814,N_1101);
nor U4734 (N_4734,N_1290,N_306);
or U4735 (N_4735,N_2395,N_2497);
xnor U4736 (N_4736,N_347,N_1948);
nor U4737 (N_4737,N_949,N_216);
nand U4738 (N_4738,N_250,N_1584);
and U4739 (N_4739,N_2100,N_2140);
and U4740 (N_4740,N_1408,N_1655);
nand U4741 (N_4741,N_920,N_141);
nand U4742 (N_4742,N_1489,N_179);
and U4743 (N_4743,N_1917,N_1374);
or U4744 (N_4744,N_1453,N_321);
and U4745 (N_4745,N_4,N_1495);
and U4746 (N_4746,N_1198,N_809);
nor U4747 (N_4747,N_1186,N_88);
or U4748 (N_4748,N_1066,N_1430);
nand U4749 (N_4749,N_2491,N_1247);
nor U4750 (N_4750,N_351,N_2143);
and U4751 (N_4751,N_366,N_349);
and U4752 (N_4752,N_568,N_2482);
nor U4753 (N_4753,N_1622,N_2127);
or U4754 (N_4754,N_673,N_1549);
nand U4755 (N_4755,N_426,N_1866);
and U4756 (N_4756,N_1194,N_381);
nand U4757 (N_4757,N_170,N_1790);
nor U4758 (N_4758,N_380,N_465);
or U4759 (N_4759,N_583,N_1502);
or U4760 (N_4760,N_334,N_203);
and U4761 (N_4761,N_291,N_2080);
and U4762 (N_4762,N_1869,N_1091);
and U4763 (N_4763,N_365,N_1087);
and U4764 (N_4764,N_1320,N_1580);
nor U4765 (N_4765,N_632,N_620);
and U4766 (N_4766,N_1616,N_434);
xor U4767 (N_4767,N_335,N_985);
or U4768 (N_4768,N_618,N_72);
nand U4769 (N_4769,N_2177,N_2028);
nor U4770 (N_4770,N_1134,N_2211);
or U4771 (N_4771,N_428,N_954);
xor U4772 (N_4772,N_1234,N_1814);
nor U4773 (N_4773,N_2235,N_1978);
nand U4774 (N_4774,N_1959,N_604);
or U4775 (N_4775,N_788,N_632);
and U4776 (N_4776,N_2105,N_1102);
nor U4777 (N_4777,N_1382,N_1357);
nand U4778 (N_4778,N_1841,N_2103);
nor U4779 (N_4779,N_1265,N_680);
and U4780 (N_4780,N_1697,N_967);
or U4781 (N_4781,N_251,N_901);
nand U4782 (N_4782,N_1923,N_2421);
nor U4783 (N_4783,N_806,N_1607);
and U4784 (N_4784,N_389,N_584);
or U4785 (N_4785,N_1165,N_1300);
nor U4786 (N_4786,N_87,N_2022);
or U4787 (N_4787,N_1093,N_2102);
and U4788 (N_4788,N_1538,N_1021);
xnor U4789 (N_4789,N_379,N_2302);
nand U4790 (N_4790,N_1289,N_1545);
nor U4791 (N_4791,N_382,N_1777);
nor U4792 (N_4792,N_462,N_1013);
nand U4793 (N_4793,N_961,N_2387);
or U4794 (N_4794,N_2276,N_2237);
nor U4795 (N_4795,N_2126,N_569);
nand U4796 (N_4796,N_2142,N_2345);
and U4797 (N_4797,N_462,N_1585);
or U4798 (N_4798,N_974,N_2091);
nor U4799 (N_4799,N_2078,N_1475);
nand U4800 (N_4800,N_1448,N_815);
and U4801 (N_4801,N_209,N_572);
nor U4802 (N_4802,N_2269,N_2290);
and U4803 (N_4803,N_1631,N_775);
or U4804 (N_4804,N_2498,N_1010);
nor U4805 (N_4805,N_2135,N_1915);
nor U4806 (N_4806,N_1808,N_2094);
nand U4807 (N_4807,N_1108,N_404);
and U4808 (N_4808,N_2077,N_557);
nor U4809 (N_4809,N_1228,N_835);
or U4810 (N_4810,N_1129,N_1126);
nand U4811 (N_4811,N_1530,N_100);
or U4812 (N_4812,N_2170,N_242);
and U4813 (N_4813,N_1899,N_1005);
nand U4814 (N_4814,N_1684,N_1133);
and U4815 (N_4815,N_1477,N_381);
nand U4816 (N_4816,N_1634,N_1961);
and U4817 (N_4817,N_1049,N_2199);
and U4818 (N_4818,N_300,N_1307);
or U4819 (N_4819,N_2006,N_408);
nor U4820 (N_4820,N_1160,N_1234);
nand U4821 (N_4821,N_1168,N_847);
nand U4822 (N_4822,N_1435,N_1248);
xor U4823 (N_4823,N_1386,N_1943);
nor U4824 (N_4824,N_2239,N_2451);
nand U4825 (N_4825,N_2265,N_2095);
nor U4826 (N_4826,N_315,N_8);
nor U4827 (N_4827,N_2107,N_1707);
nor U4828 (N_4828,N_1260,N_1860);
nor U4829 (N_4829,N_2406,N_308);
nand U4830 (N_4830,N_2122,N_688);
xnor U4831 (N_4831,N_804,N_1637);
or U4832 (N_4832,N_1981,N_553);
or U4833 (N_4833,N_737,N_2210);
nor U4834 (N_4834,N_2003,N_984);
nor U4835 (N_4835,N_273,N_2436);
nand U4836 (N_4836,N_1897,N_253);
or U4837 (N_4837,N_881,N_2407);
nand U4838 (N_4838,N_1265,N_2077);
or U4839 (N_4839,N_1497,N_118);
nand U4840 (N_4840,N_782,N_2112);
and U4841 (N_4841,N_1674,N_977);
nand U4842 (N_4842,N_2456,N_1931);
and U4843 (N_4843,N_1934,N_1602);
and U4844 (N_4844,N_730,N_1820);
and U4845 (N_4845,N_1799,N_1691);
and U4846 (N_4846,N_1438,N_1208);
or U4847 (N_4847,N_914,N_2171);
nand U4848 (N_4848,N_1270,N_1244);
or U4849 (N_4849,N_1333,N_2226);
or U4850 (N_4850,N_1950,N_2451);
nand U4851 (N_4851,N_1896,N_336);
and U4852 (N_4852,N_1495,N_1197);
or U4853 (N_4853,N_1512,N_97);
or U4854 (N_4854,N_778,N_2033);
or U4855 (N_4855,N_53,N_10);
nor U4856 (N_4856,N_135,N_733);
nor U4857 (N_4857,N_549,N_1844);
and U4858 (N_4858,N_2087,N_1297);
or U4859 (N_4859,N_1467,N_988);
nand U4860 (N_4860,N_854,N_228);
xnor U4861 (N_4861,N_2131,N_1377);
nand U4862 (N_4862,N_587,N_2112);
nor U4863 (N_4863,N_1933,N_1467);
or U4864 (N_4864,N_2247,N_246);
nand U4865 (N_4865,N_2042,N_2178);
and U4866 (N_4866,N_1323,N_1224);
or U4867 (N_4867,N_106,N_2234);
nand U4868 (N_4868,N_1294,N_883);
and U4869 (N_4869,N_1542,N_1228);
nor U4870 (N_4870,N_1344,N_2330);
nor U4871 (N_4871,N_889,N_656);
nor U4872 (N_4872,N_691,N_91);
and U4873 (N_4873,N_1755,N_104);
nand U4874 (N_4874,N_834,N_1222);
or U4875 (N_4875,N_2294,N_1502);
or U4876 (N_4876,N_301,N_1159);
and U4877 (N_4877,N_1753,N_2135);
xor U4878 (N_4878,N_1272,N_351);
nand U4879 (N_4879,N_141,N_2280);
or U4880 (N_4880,N_136,N_1050);
and U4881 (N_4881,N_2198,N_290);
or U4882 (N_4882,N_1524,N_1346);
nand U4883 (N_4883,N_1484,N_442);
nor U4884 (N_4884,N_150,N_953);
and U4885 (N_4885,N_865,N_350);
and U4886 (N_4886,N_433,N_1178);
nand U4887 (N_4887,N_1975,N_178);
nand U4888 (N_4888,N_776,N_1203);
nand U4889 (N_4889,N_471,N_2322);
nand U4890 (N_4890,N_983,N_918);
or U4891 (N_4891,N_308,N_411);
nor U4892 (N_4892,N_376,N_2347);
nor U4893 (N_4893,N_2477,N_1677);
nand U4894 (N_4894,N_2261,N_1612);
or U4895 (N_4895,N_912,N_1558);
or U4896 (N_4896,N_2308,N_2291);
nand U4897 (N_4897,N_2261,N_1434);
and U4898 (N_4898,N_1551,N_1608);
nand U4899 (N_4899,N_2324,N_2448);
or U4900 (N_4900,N_1023,N_239);
and U4901 (N_4901,N_811,N_1805);
and U4902 (N_4902,N_1678,N_1010);
or U4903 (N_4903,N_2251,N_1175);
and U4904 (N_4904,N_947,N_2271);
nor U4905 (N_4905,N_315,N_498);
or U4906 (N_4906,N_1388,N_1078);
xnor U4907 (N_4907,N_2065,N_103);
or U4908 (N_4908,N_845,N_610);
xnor U4909 (N_4909,N_395,N_1861);
and U4910 (N_4910,N_1392,N_719);
nor U4911 (N_4911,N_587,N_2350);
xor U4912 (N_4912,N_2191,N_634);
or U4913 (N_4913,N_1662,N_2162);
nor U4914 (N_4914,N_1660,N_2130);
nor U4915 (N_4915,N_1270,N_910);
or U4916 (N_4916,N_40,N_2273);
xnor U4917 (N_4917,N_801,N_1111);
nand U4918 (N_4918,N_479,N_2319);
and U4919 (N_4919,N_1675,N_317);
or U4920 (N_4920,N_1479,N_1344);
and U4921 (N_4921,N_1730,N_1469);
xnor U4922 (N_4922,N_834,N_1067);
xor U4923 (N_4923,N_1948,N_350);
or U4924 (N_4924,N_846,N_2262);
nor U4925 (N_4925,N_2398,N_1340);
and U4926 (N_4926,N_2222,N_1833);
or U4927 (N_4927,N_415,N_2356);
nor U4928 (N_4928,N_1724,N_1481);
nand U4929 (N_4929,N_1138,N_539);
nor U4930 (N_4930,N_37,N_1032);
nor U4931 (N_4931,N_37,N_98);
nor U4932 (N_4932,N_1747,N_978);
nand U4933 (N_4933,N_1497,N_865);
and U4934 (N_4934,N_1982,N_1626);
nand U4935 (N_4935,N_2025,N_102);
nand U4936 (N_4936,N_285,N_1595);
and U4937 (N_4937,N_309,N_241);
or U4938 (N_4938,N_1533,N_458);
nand U4939 (N_4939,N_457,N_1779);
nor U4940 (N_4940,N_812,N_445);
and U4941 (N_4941,N_2460,N_248);
nand U4942 (N_4942,N_2001,N_244);
or U4943 (N_4943,N_1216,N_382);
and U4944 (N_4944,N_2397,N_302);
nand U4945 (N_4945,N_906,N_1058);
or U4946 (N_4946,N_1508,N_117);
and U4947 (N_4947,N_76,N_746);
or U4948 (N_4948,N_499,N_771);
and U4949 (N_4949,N_5,N_840);
or U4950 (N_4950,N_1602,N_1229);
and U4951 (N_4951,N_203,N_196);
nand U4952 (N_4952,N_785,N_1041);
nor U4953 (N_4953,N_1015,N_528);
nand U4954 (N_4954,N_1642,N_1105);
nor U4955 (N_4955,N_2278,N_1534);
nor U4956 (N_4956,N_1972,N_688);
nor U4957 (N_4957,N_1478,N_2277);
nor U4958 (N_4958,N_844,N_450);
nor U4959 (N_4959,N_651,N_1838);
or U4960 (N_4960,N_797,N_182);
and U4961 (N_4961,N_2248,N_1510);
nor U4962 (N_4962,N_1248,N_1752);
nor U4963 (N_4963,N_1165,N_810);
and U4964 (N_4964,N_137,N_1939);
nor U4965 (N_4965,N_1436,N_740);
nor U4966 (N_4966,N_2054,N_1351);
and U4967 (N_4967,N_182,N_1664);
nand U4968 (N_4968,N_929,N_2163);
and U4969 (N_4969,N_480,N_872);
or U4970 (N_4970,N_141,N_2042);
or U4971 (N_4971,N_2055,N_1507);
nor U4972 (N_4972,N_939,N_424);
or U4973 (N_4973,N_356,N_1167);
or U4974 (N_4974,N_684,N_489);
and U4975 (N_4975,N_1346,N_1858);
nor U4976 (N_4976,N_200,N_1595);
and U4977 (N_4977,N_200,N_103);
and U4978 (N_4978,N_378,N_298);
xor U4979 (N_4979,N_532,N_3);
nor U4980 (N_4980,N_1568,N_1012);
nor U4981 (N_4981,N_2354,N_1701);
nor U4982 (N_4982,N_429,N_1815);
nor U4983 (N_4983,N_554,N_2451);
nor U4984 (N_4984,N_22,N_1213);
and U4985 (N_4985,N_1686,N_1960);
or U4986 (N_4986,N_1664,N_1887);
and U4987 (N_4987,N_2350,N_323);
nand U4988 (N_4988,N_2135,N_1342);
or U4989 (N_4989,N_1469,N_1149);
nand U4990 (N_4990,N_1264,N_947);
nor U4991 (N_4991,N_2355,N_1503);
nand U4992 (N_4992,N_1636,N_347);
or U4993 (N_4993,N_2330,N_1648);
or U4994 (N_4994,N_316,N_1791);
or U4995 (N_4995,N_935,N_2037);
nor U4996 (N_4996,N_1095,N_974);
nor U4997 (N_4997,N_1943,N_1147);
or U4998 (N_4998,N_1487,N_2181);
nand U4999 (N_4999,N_2023,N_2431);
or UO_0 (O_0,N_3209,N_4842);
or UO_1 (O_1,N_3256,N_2700);
nand UO_2 (O_2,N_3383,N_4500);
nand UO_3 (O_3,N_4824,N_4529);
and UO_4 (O_4,N_3299,N_4817);
nand UO_5 (O_5,N_3432,N_2760);
nand UO_6 (O_6,N_4343,N_2514);
and UO_7 (O_7,N_2604,N_2814);
nor UO_8 (O_8,N_3986,N_4252);
or UO_9 (O_9,N_4627,N_4598);
nand UO_10 (O_10,N_3886,N_3021);
nand UO_11 (O_11,N_2569,N_3970);
or UO_12 (O_12,N_3277,N_2703);
or UO_13 (O_13,N_3902,N_3611);
nor UO_14 (O_14,N_2948,N_4528);
or UO_15 (O_15,N_4808,N_3113);
xor UO_16 (O_16,N_3315,N_4359);
nor UO_17 (O_17,N_3932,N_4238);
and UO_18 (O_18,N_4155,N_2534);
nor UO_19 (O_19,N_3723,N_4411);
nor UO_20 (O_20,N_3001,N_3384);
nand UO_21 (O_21,N_4632,N_3865);
and UO_22 (O_22,N_3956,N_3910);
or UO_23 (O_23,N_2682,N_3199);
nor UO_24 (O_24,N_4163,N_2780);
or UO_25 (O_25,N_4957,N_4869);
nor UO_26 (O_26,N_4414,N_3559);
and UO_27 (O_27,N_4172,N_3118);
and UO_28 (O_28,N_3202,N_4699);
nor UO_29 (O_29,N_4118,N_4653);
nand UO_30 (O_30,N_4625,N_3893);
or UO_31 (O_31,N_4294,N_4487);
xor UO_32 (O_32,N_2594,N_4066);
nand UO_33 (O_33,N_2723,N_3575);
nor UO_34 (O_34,N_2676,N_4484);
or UO_35 (O_35,N_4917,N_4948);
and UO_36 (O_36,N_4042,N_3187);
nand UO_37 (O_37,N_2694,N_3549);
nand UO_38 (O_38,N_4436,N_4904);
nor UO_39 (O_39,N_4090,N_3177);
nand UO_40 (O_40,N_4406,N_3396);
and UO_41 (O_41,N_4051,N_2727);
xor UO_42 (O_42,N_2848,N_4490);
nand UO_43 (O_43,N_3352,N_2699);
and UO_44 (O_44,N_2605,N_3905);
or UO_45 (O_45,N_4469,N_4805);
nor UO_46 (O_46,N_3420,N_2769);
and UO_47 (O_47,N_3258,N_4746);
nor UO_48 (O_48,N_3316,N_3564);
nand UO_49 (O_49,N_2807,N_2909);
and UO_50 (O_50,N_4320,N_3616);
and UO_51 (O_51,N_3321,N_3601);
and UO_52 (O_52,N_4459,N_2667);
and UO_53 (O_53,N_3988,N_4416);
nand UO_54 (O_54,N_2901,N_2571);
nand UO_55 (O_55,N_3608,N_4939);
and UO_56 (O_56,N_4872,N_4765);
nand UO_57 (O_57,N_4680,N_4697);
nor UO_58 (O_58,N_4547,N_2643);
or UO_59 (O_59,N_4046,N_4179);
or UO_60 (O_60,N_3448,N_3617);
nor UO_61 (O_61,N_4870,N_3598);
and UO_62 (O_62,N_4236,N_3968);
nand UO_63 (O_63,N_4700,N_4464);
nor UO_64 (O_64,N_4731,N_4479);
or UO_65 (O_65,N_2566,N_4912);
nand UO_66 (O_66,N_4387,N_3569);
nand UO_67 (O_67,N_2639,N_2949);
or UO_68 (O_68,N_2838,N_2874);
or UO_69 (O_69,N_2911,N_3785);
nand UO_70 (O_70,N_4705,N_4609);
xnor UO_71 (O_71,N_2952,N_3119);
nand UO_72 (O_72,N_3057,N_2653);
and UO_73 (O_73,N_4723,N_3389);
nor UO_74 (O_74,N_3832,N_4199);
or UO_75 (O_75,N_3023,N_4181);
xor UO_76 (O_76,N_4794,N_3010);
nor UO_77 (O_77,N_2711,N_3969);
and UO_78 (O_78,N_3718,N_3711);
nor UO_79 (O_79,N_3732,N_3132);
nor UO_80 (O_80,N_4292,N_3154);
or UO_81 (O_81,N_2775,N_2702);
and UO_82 (O_82,N_4112,N_2763);
or UO_83 (O_83,N_3766,N_2597);
nand UO_84 (O_84,N_4345,N_4425);
nand UO_85 (O_85,N_4076,N_4220);
or UO_86 (O_86,N_4867,N_4065);
nand UO_87 (O_87,N_4122,N_3955);
and UO_88 (O_88,N_3137,N_2628);
nand UO_89 (O_89,N_4933,N_2512);
nand UO_90 (O_90,N_4839,N_2520);
or UO_91 (O_91,N_4169,N_3930);
or UO_92 (O_92,N_2784,N_3659);
or UO_93 (O_93,N_3896,N_4761);
nor UO_94 (O_94,N_3771,N_4207);
nor UO_95 (O_95,N_2560,N_3128);
nor UO_96 (O_96,N_3176,N_4716);
or UO_97 (O_97,N_3715,N_4778);
and UO_98 (O_98,N_3249,N_3740);
or UO_99 (O_99,N_2985,N_3116);
nand UO_100 (O_100,N_4015,N_3760);
nor UO_101 (O_101,N_3962,N_3752);
nor UO_102 (O_102,N_2946,N_3989);
and UO_103 (O_103,N_2659,N_3470);
nor UO_104 (O_104,N_4428,N_2636);
nand UO_105 (O_105,N_4634,N_4200);
and UO_106 (O_106,N_3139,N_2929);
nor UO_107 (O_107,N_3933,N_2777);
and UO_108 (O_108,N_3793,N_4764);
nor UO_109 (O_109,N_3579,N_4696);
and UO_110 (O_110,N_3336,N_4044);
or UO_111 (O_111,N_3141,N_2774);
xor UO_112 (O_112,N_4116,N_2559);
and UO_113 (O_113,N_4970,N_3427);
nand UO_114 (O_114,N_3779,N_4098);
nor UO_115 (O_115,N_3269,N_3061);
and UO_116 (O_116,N_4519,N_3040);
nor UO_117 (O_117,N_2545,N_3800);
nor UO_118 (O_118,N_2741,N_2778);
and UO_119 (O_119,N_3223,N_4813);
and UO_120 (O_120,N_2794,N_2817);
nand UO_121 (O_121,N_2797,N_4936);
nor UO_122 (O_122,N_4997,N_4141);
nor UO_123 (O_123,N_4043,N_4149);
nand UO_124 (O_124,N_3816,N_3756);
nand UO_125 (O_125,N_4126,N_4893);
nor UO_126 (O_126,N_2564,N_3033);
or UO_127 (O_127,N_4018,N_4173);
and UO_128 (O_128,N_4014,N_3541);
and UO_129 (O_129,N_4877,N_4121);
and UO_130 (O_130,N_2841,N_3327);
nor UO_131 (O_131,N_3295,N_4084);
xnor UO_132 (O_132,N_2772,N_2502);
and UO_133 (O_133,N_4689,N_4439);
xnor UO_134 (O_134,N_4158,N_3422);
nor UO_135 (O_135,N_4366,N_3878);
nand UO_136 (O_136,N_4575,N_2984);
nor UO_137 (O_137,N_4706,N_4017);
nor UO_138 (O_138,N_2930,N_3644);
and UO_139 (O_139,N_4100,N_4771);
or UO_140 (O_140,N_4559,N_3346);
and UO_141 (O_141,N_4287,N_4190);
nor UO_142 (O_142,N_3812,N_4368);
and UO_143 (O_143,N_2548,N_3387);
nor UO_144 (O_144,N_3849,N_3670);
or UO_145 (O_145,N_4463,N_3610);
nand UO_146 (O_146,N_3882,N_3158);
or UO_147 (O_147,N_2630,N_3998);
and UO_148 (O_148,N_4719,N_3028);
xnor UO_149 (O_149,N_3866,N_3762);
or UO_150 (O_150,N_4119,N_4692);
nor UO_151 (O_151,N_4070,N_3085);
and UO_152 (O_152,N_4526,N_2710);
nor UO_153 (O_153,N_2611,N_3841);
nand UO_154 (O_154,N_2799,N_3909);
nand UO_155 (O_155,N_3661,N_4483);
or UO_156 (O_156,N_3114,N_4311);
nand UO_157 (O_157,N_4989,N_3586);
or UO_158 (O_158,N_3412,N_4924);
and UO_159 (O_159,N_3250,N_3254);
or UO_160 (O_160,N_4064,N_2743);
or UO_161 (O_161,N_3538,N_3043);
nand UO_162 (O_162,N_4478,N_3105);
nand UO_163 (O_163,N_2875,N_3046);
or UO_164 (O_164,N_4342,N_3613);
nor UO_165 (O_165,N_4391,N_3546);
or UO_166 (O_166,N_4777,N_3960);
or UO_167 (O_167,N_3974,N_4021);
nor UO_168 (O_168,N_4423,N_3870);
nand UO_169 (O_169,N_3386,N_3927);
or UO_170 (O_170,N_2978,N_3237);
nand UO_171 (O_171,N_4148,N_3438);
and UO_172 (O_172,N_3366,N_3683);
nand UO_173 (O_173,N_4170,N_3797);
nor UO_174 (O_174,N_3248,N_3984);
xor UO_175 (O_175,N_4377,N_3576);
or UO_176 (O_176,N_4916,N_2937);
or UO_177 (O_177,N_3775,N_3458);
or UO_178 (O_178,N_3338,N_3399);
nand UO_179 (O_179,N_4274,N_2585);
and UO_180 (O_180,N_3450,N_3496);
nand UO_181 (O_181,N_3794,N_4328);
nor UO_182 (O_182,N_4730,N_4056);
and UO_183 (O_183,N_4748,N_2574);
nor UO_184 (O_184,N_3645,N_3398);
nand UO_185 (O_185,N_3709,N_4131);
nor UO_186 (O_186,N_2675,N_3138);
or UO_187 (O_187,N_2558,N_3983);
nand UO_188 (O_188,N_4826,N_4000);
and UO_189 (O_189,N_2668,N_3946);
nor UO_190 (O_190,N_3349,N_3703);
nand UO_191 (O_191,N_4427,N_3551);
and UO_192 (O_192,N_2579,N_2608);
nor UO_193 (O_193,N_4544,N_3431);
nor UO_194 (O_194,N_2693,N_3791);
nand UO_195 (O_195,N_2537,N_3308);
or UO_196 (O_196,N_4074,N_4347);
nand UO_197 (O_197,N_3235,N_2891);
or UO_198 (O_198,N_3846,N_4433);
or UO_199 (O_199,N_4117,N_3646);
and UO_200 (O_200,N_4344,N_4928);
or UO_201 (O_201,N_2598,N_4758);
and UO_202 (O_202,N_3894,N_4979);
and UO_203 (O_203,N_3951,N_4790);
and UO_204 (O_204,N_2733,N_4623);
nand UO_205 (O_205,N_3919,N_2565);
or UO_206 (O_206,N_4410,N_4862);
nor UO_207 (O_207,N_3035,N_3351);
and UO_208 (O_208,N_2629,N_4266);
nor UO_209 (O_209,N_4192,N_4228);
and UO_210 (O_210,N_4278,N_4454);
and UO_211 (O_211,N_3149,N_4509);
or UO_212 (O_212,N_3633,N_3436);
and UO_213 (O_213,N_3978,N_3699);
nor UO_214 (O_214,N_2886,N_3086);
nand UO_215 (O_215,N_2958,N_4740);
and UO_216 (O_216,N_2570,N_3531);
or UO_217 (O_217,N_2928,N_3397);
and UO_218 (O_218,N_2589,N_3708);
nor UO_219 (O_219,N_3244,N_4766);
and UO_220 (O_220,N_4827,N_4203);
nor UO_221 (O_221,N_3217,N_4154);
nand UO_222 (O_222,N_4966,N_3133);
nor UO_223 (O_223,N_2821,N_4330);
nor UO_224 (O_224,N_4047,N_3411);
nand UO_225 (O_225,N_3545,N_4739);
nand UO_226 (O_226,N_3678,N_3941);
nor UO_227 (O_227,N_4269,N_3243);
or UO_228 (O_228,N_4360,N_4830);
and UO_229 (O_229,N_3260,N_3591);
and UO_230 (O_230,N_3424,N_3247);
and UO_231 (O_231,N_2756,N_3685);
nand UO_232 (O_232,N_3582,N_2873);
and UO_233 (O_233,N_3554,N_3289);
nand UO_234 (O_234,N_4213,N_3925);
or UO_235 (O_235,N_3305,N_3500);
nand UO_236 (O_236,N_4089,N_3662);
nor UO_237 (O_237,N_3855,N_4524);
nand UO_238 (O_238,N_3804,N_3754);
and UO_239 (O_239,N_4222,N_2987);
nand UO_240 (O_240,N_3587,N_2536);
nor UO_241 (O_241,N_4803,N_3290);
nor UO_242 (O_242,N_3126,N_3637);
and UO_243 (O_243,N_4115,N_3639);
and UO_244 (O_244,N_2590,N_3167);
and UO_245 (O_245,N_2744,N_4334);
nor UO_246 (O_246,N_4372,N_4136);
nor UO_247 (O_247,N_3129,N_3150);
nor UO_248 (O_248,N_2941,N_2840);
nor UO_249 (O_249,N_4254,N_4340);
nor UO_250 (O_250,N_3102,N_4897);
nor UO_251 (O_251,N_4965,N_3810);
or UO_252 (O_252,N_4068,N_2730);
or UO_253 (O_253,N_3056,N_4844);
and UO_254 (O_254,N_4822,N_3859);
nand UO_255 (O_255,N_3328,N_3985);
nor UO_256 (O_256,N_3274,N_2642);
nor UO_257 (O_257,N_2896,N_2738);
nand UO_258 (O_258,N_3442,N_4140);
nor UO_259 (O_259,N_4773,N_4921);
or UO_260 (O_260,N_4556,N_2795);
xnor UO_261 (O_261,N_4289,N_2851);
nand UO_262 (O_262,N_2584,N_4592);
or UO_263 (O_263,N_3618,N_2940);
nor UO_264 (O_264,N_4071,N_3967);
nand UO_265 (O_265,N_4704,N_4364);
or UO_266 (O_266,N_2871,N_3702);
nand UO_267 (O_267,N_3823,N_4810);
or UO_268 (O_268,N_3065,N_4395);
nor UO_269 (O_269,N_4027,N_4058);
nor UO_270 (O_270,N_3272,N_4506);
xnor UO_271 (O_271,N_4501,N_4574);
nand UO_272 (O_272,N_4549,N_3484);
nand UO_273 (O_273,N_4168,N_2981);
nand UO_274 (O_274,N_3515,N_3140);
nand UO_275 (O_275,N_3924,N_4889);
nand UO_276 (O_276,N_3296,N_3811);
and UO_277 (O_277,N_4841,N_2706);
or UO_278 (O_278,N_2877,N_4796);
nand UO_279 (O_279,N_2971,N_3799);
nor UO_280 (O_280,N_2934,N_2866);
or UO_281 (O_281,N_4201,N_3142);
and UO_282 (O_282,N_2712,N_4657);
and UO_283 (O_283,N_4217,N_2771);
or UO_284 (O_284,N_4262,N_2964);
xor UO_285 (O_285,N_4494,N_3098);
or UO_286 (O_286,N_2804,N_2829);
nand UO_287 (O_287,N_3405,N_3401);
and UO_288 (O_288,N_3495,N_4847);
or UO_289 (O_289,N_3344,N_4031);
and UO_290 (O_290,N_4049,N_2510);
or UO_291 (O_291,N_2539,N_2845);
or UO_292 (O_292,N_4888,N_2677);
nor UO_293 (O_293,N_4045,N_3625);
or UO_294 (O_294,N_3883,N_3162);
or UO_295 (O_295,N_4283,N_4527);
or UO_296 (O_296,N_4521,N_3578);
nand UO_297 (O_297,N_3293,N_3285);
or UO_298 (O_298,N_4781,N_4910);
xnor UO_299 (O_299,N_2783,N_4750);
nor UO_300 (O_300,N_2623,N_3940);
xor UO_301 (O_301,N_2592,N_2811);
or UO_302 (O_302,N_3547,N_3337);
or UO_303 (O_303,N_2983,N_2547);
and UO_304 (O_304,N_2820,N_2870);
nand UO_305 (O_305,N_3310,N_3034);
nand UO_306 (O_306,N_4276,N_3440);
xor UO_307 (O_307,N_3751,N_2962);
or UO_308 (O_308,N_4272,N_4645);
nor UO_309 (O_309,N_4493,N_3392);
and UO_310 (O_310,N_4488,N_3125);
and UO_311 (O_311,N_4963,N_4130);
or UO_312 (O_312,N_4313,N_3556);
nand UO_313 (O_313,N_3444,N_4435);
or UO_314 (O_314,N_4404,N_3172);
and UO_315 (O_315,N_2939,N_3630);
nand UO_316 (O_316,N_4390,N_3688);
nor UO_317 (O_317,N_3789,N_3068);
and UO_318 (O_318,N_3897,N_4134);
nor UO_319 (O_319,N_3627,N_2790);
nand UO_320 (O_320,N_3560,N_3343);
and UO_321 (O_321,N_3170,N_2853);
nor UO_322 (O_322,N_3101,N_3183);
nand UO_323 (O_323,N_4747,N_3777);
nand UO_324 (O_324,N_3080,N_3211);
nand UO_325 (O_325,N_3558,N_4980);
or UO_326 (O_326,N_3311,N_4431);
nor UO_327 (O_327,N_4838,N_4094);
or UO_328 (O_328,N_4848,N_4854);
nor UO_329 (O_329,N_3548,N_3692);
and UO_330 (O_330,N_4073,N_3091);
nor UO_331 (O_331,N_2809,N_3148);
nand UO_332 (O_332,N_3568,N_4636);
nor UO_333 (O_333,N_3938,N_4477);
nor UO_334 (O_334,N_4284,N_4260);
and UO_335 (O_335,N_3748,N_3522);
or UO_336 (O_336,N_2836,N_3075);
nand UO_337 (O_337,N_2640,N_3070);
nor UO_338 (O_338,N_2852,N_3246);
nor UO_339 (O_339,N_3038,N_4566);
or UO_340 (O_340,N_3850,N_3469);
xor UO_341 (O_341,N_3270,N_4452);
or UO_342 (O_342,N_3773,N_4422);
nor UO_343 (O_343,N_3332,N_4310);
nor UO_344 (O_344,N_2543,N_3219);
or UO_345 (O_345,N_4316,N_3212);
nor UO_346 (O_346,N_3543,N_4297);
nor UO_347 (O_347,N_3020,N_3782);
or UO_348 (O_348,N_3421,N_3255);
or UO_349 (O_349,N_4481,N_4184);
nand UO_350 (O_350,N_4654,N_2942);
nand UO_351 (O_351,N_4307,N_3901);
nor UO_352 (O_352,N_3441,N_3370);
and UO_353 (O_353,N_3130,N_2997);
nand UO_354 (O_354,N_4441,N_4296);
and UO_355 (O_355,N_3889,N_4954);
or UO_356 (O_356,N_2862,N_3996);
nor UO_357 (O_357,N_3404,N_3284);
and UO_358 (O_358,N_3206,N_4879);
or UO_359 (O_359,N_4124,N_2861);
or UO_360 (O_360,N_3503,N_3561);
and UO_361 (O_361,N_3261,N_3191);
or UO_362 (O_362,N_4577,N_3914);
and UO_363 (O_363,N_4235,N_3487);
nor UO_364 (O_364,N_4261,N_4554);
and UO_365 (O_365,N_3577,N_3192);
nor UO_366 (O_366,N_2600,N_4920);
nand UO_367 (O_367,N_4964,N_4934);
nand UO_368 (O_368,N_2705,N_2707);
or UO_369 (O_369,N_3006,N_4985);
and UO_370 (O_370,N_2669,N_4202);
or UO_371 (O_371,N_3697,N_2526);
nand UO_372 (O_372,N_3626,N_2854);
nand UO_373 (O_373,N_3977,N_3048);
or UO_374 (O_374,N_3829,N_4432);
or UO_375 (O_375,N_3391,N_2721);
nor UO_376 (O_376,N_4756,N_2519);
or UO_377 (O_377,N_3761,N_2620);
nor UO_378 (O_378,N_4639,N_4323);
or UO_379 (O_379,N_2660,N_4762);
nor UO_380 (O_380,N_4718,N_3210);
and UO_381 (O_381,N_3072,N_3066);
nand UO_382 (O_382,N_3847,N_4512);
nand UO_383 (O_383,N_3372,N_4288);
or UO_384 (O_384,N_3701,N_2552);
nor UO_385 (O_385,N_4511,N_2954);
and UO_386 (O_386,N_4153,N_4570);
nand UO_387 (O_387,N_3093,N_4754);
and UO_388 (O_388,N_3224,N_3347);
nand UO_389 (O_389,N_4470,N_3529);
nand UO_390 (O_390,N_4429,N_2793);
and UO_391 (O_391,N_4249,N_4550);
or UO_392 (O_392,N_4702,N_4557);
nor UO_393 (O_393,N_3062,N_3651);
or UO_394 (O_394,N_3030,N_3667);
or UO_395 (O_395,N_4744,N_3875);
nor UO_396 (O_396,N_4711,N_3051);
and UO_397 (O_397,N_4453,N_3871);
nor UO_398 (O_398,N_3840,N_4319);
nor UO_399 (O_399,N_3417,N_3749);
nand UO_400 (O_400,N_2745,N_4461);
nor UO_401 (O_401,N_2750,N_4157);
or UO_402 (O_402,N_3200,N_4874);
and UO_403 (O_403,N_3201,N_3121);
or UO_404 (O_404,N_3884,N_4197);
nor UO_405 (O_405,N_3359,N_2881);
or UO_406 (O_406,N_3781,N_4152);
and UO_407 (O_407,N_3599,N_2834);
or UO_408 (O_408,N_2747,N_3472);
nor UO_409 (O_409,N_2791,N_3981);
nand UO_410 (O_410,N_2782,N_4767);
and UO_411 (O_411,N_4003,N_3302);
or UO_412 (O_412,N_4769,N_4722);
nand UO_413 (O_413,N_4402,N_4104);
nand UO_414 (O_414,N_4851,N_2806);
and UO_415 (O_415,N_4975,N_3205);
nor UO_416 (O_416,N_3253,N_2562);
nor UO_417 (O_417,N_3032,N_4816);
and UO_418 (O_418,N_3573,N_4178);
nor UO_419 (O_419,N_2524,N_4476);
or UO_420 (O_420,N_2500,N_3265);
nor UO_421 (O_421,N_4129,N_3948);
nor UO_422 (O_422,N_3297,N_3013);
nor UO_423 (O_423,N_4388,N_4514);
nand UO_424 (O_424,N_3227,N_3473);
nor UO_425 (O_425,N_3959,N_2991);
and UO_426 (O_426,N_3844,N_3720);
nand UO_427 (O_427,N_4397,N_4187);
nand UO_428 (O_428,N_4026,N_2732);
and UO_429 (O_429,N_4362,N_4298);
or UO_430 (O_430,N_2554,N_3159);
nand UO_431 (O_431,N_4434,N_3004);
and UO_432 (O_432,N_4150,N_3593);
or UO_433 (O_433,N_3188,N_2625);
nand UO_434 (O_434,N_3929,N_4335);
nand UO_435 (O_435,N_3251,N_3609);
or UO_436 (O_436,N_4931,N_4091);
nand UO_437 (O_437,N_4729,N_3658);
and UO_438 (O_438,N_4629,N_4166);
nor UO_439 (O_439,N_3232,N_3208);
and UO_440 (O_440,N_4788,N_2779);
nand UO_441 (O_441,N_4537,N_2754);
or UO_442 (O_442,N_3679,N_3220);
nor UO_443 (O_443,N_4502,N_4690);
and UO_444 (O_444,N_4852,N_3835);
and UO_445 (O_445,N_3942,N_3742);
and UO_446 (O_446,N_2905,N_3462);
nand UO_447 (O_447,N_4160,N_3413);
nor UO_448 (O_448,N_3478,N_4635);
nor UO_449 (O_449,N_3197,N_4321);
and UO_450 (O_450,N_2992,N_4038);
or UO_451 (O_451,N_3012,N_3737);
and UO_452 (O_452,N_3673,N_3203);
nor UO_453 (O_453,N_3447,N_3257);
and UO_454 (O_454,N_2781,N_2726);
nor UO_455 (O_455,N_4571,N_2900);
or UO_456 (O_456,N_2551,N_4415);
nand UO_457 (O_457,N_2926,N_4595);
nor UO_458 (O_458,N_3433,N_3088);
nor UO_459 (O_459,N_2801,N_2748);
nand UO_460 (O_460,N_4322,N_3923);
nor UO_461 (O_461,N_3163,N_2931);
and UO_462 (O_462,N_3428,N_4915);
and UO_463 (O_463,N_4976,N_4780);
nor UO_464 (O_464,N_3229,N_3060);
or UO_465 (O_465,N_4438,N_4505);
xor UO_466 (O_466,N_3348,N_3241);
nor UO_467 (O_467,N_4608,N_4779);
nand UO_468 (O_468,N_4688,N_4006);
or UO_469 (O_469,N_3475,N_3382);
or UO_470 (O_470,N_4681,N_4620);
or UO_471 (O_471,N_3081,N_4137);
and UO_472 (O_472,N_2802,N_3367);
nand UO_473 (O_473,N_4396,N_2557);
or UO_474 (O_474,N_3283,N_2785);
nand UO_475 (O_475,N_4102,N_3731);
nor UO_476 (O_476,N_2691,N_4687);
nand UO_477 (O_477,N_4455,N_2595);
nand UO_478 (O_478,N_3222,N_4182);
and UO_479 (O_479,N_3406,N_2812);
and UO_480 (O_480,N_2616,N_2768);
nand UO_481 (O_481,N_4683,N_4111);
nand UO_482 (O_482,N_2957,N_3824);
or UO_483 (O_483,N_4010,N_4811);
or UO_484 (O_484,N_2767,N_2815);
nand UO_485 (O_485,N_4389,N_3964);
or UO_486 (O_486,N_3054,N_2507);
or UO_487 (O_487,N_4774,N_3533);
or UO_488 (O_488,N_3600,N_2522);
or UO_489 (O_489,N_2567,N_3763);
nand UO_490 (O_490,N_4244,N_4108);
or UO_491 (O_491,N_3542,N_4281);
and UO_492 (O_492,N_4290,N_3641);
or UO_493 (O_493,N_2907,N_3860);
nor UO_494 (O_494,N_2830,N_3803);
or UO_495 (O_495,N_3862,N_3485);
and UO_496 (O_496,N_4485,N_4309);
and UO_497 (O_497,N_2665,N_4370);
nand UO_498 (O_498,N_4365,N_4231);
nand UO_499 (O_499,N_4473,N_2530);
nand UO_500 (O_500,N_4881,N_3186);
and UO_501 (O_501,N_4326,N_2880);
nand UO_502 (O_502,N_3378,N_4471);
and UO_503 (O_503,N_3912,N_2683);
and UO_504 (O_504,N_4792,N_2920);
and UO_505 (O_505,N_3566,N_4600);
or UO_506 (O_506,N_3079,N_2864);
nor UO_507 (O_507,N_3373,N_4306);
nor UO_508 (O_508,N_4301,N_2687);
nor UO_509 (O_509,N_4241,N_4599);
nor UO_510 (O_510,N_2725,N_3796);
and UO_511 (O_511,N_4234,N_2662);
nor UO_512 (O_512,N_2986,N_2935);
or UO_513 (O_513,N_3103,N_4617);
and UO_514 (O_514,N_3466,N_2722);
nor UO_515 (O_515,N_4355,N_3848);
or UO_516 (O_516,N_4945,N_2527);
or UO_517 (O_517,N_4646,N_4403);
or UO_518 (O_518,N_3022,N_3371);
nand UO_519 (O_519,N_3459,N_3745);
or UO_520 (O_520,N_2843,N_4019);
and UO_521 (O_521,N_3122,N_2916);
and UO_522 (O_522,N_3917,N_4812);
nor UO_523 (O_523,N_2601,N_3242);
nand UO_524 (O_524,N_4357,N_4315);
nor UO_525 (O_525,N_3842,N_4772);
or UO_526 (O_526,N_2739,N_4725);
nand UO_527 (O_527,N_4417,N_3614);
nand UO_528 (O_528,N_3306,N_4226);
nor UO_529 (O_529,N_3317,N_3672);
nand UO_530 (O_530,N_2813,N_3082);
nor UO_531 (O_531,N_4616,N_4998);
and UO_532 (O_532,N_3288,N_4132);
nor UO_533 (O_533,N_4383,N_3368);
nand UO_534 (O_534,N_4679,N_2619);
or UO_535 (O_535,N_3628,N_2919);
nor UO_536 (O_536,N_3997,N_3668);
nor UO_537 (O_537,N_3069,N_3120);
nand UO_538 (O_538,N_4958,N_4578);
and UO_539 (O_539,N_4607,N_3590);
and UO_540 (O_540,N_3820,N_4906);
nor UO_541 (O_541,N_3390,N_2859);
or UO_542 (O_542,N_4709,N_3580);
nand UO_543 (O_543,N_4551,N_4806);
and UO_544 (O_544,N_4703,N_3234);
and UO_545 (O_545,N_4626,N_4938);
nor UO_546 (O_546,N_4969,N_3706);
and UO_547 (O_547,N_2827,N_4176);
xnor UO_548 (O_548,N_4759,N_4894);
or UO_549 (O_549,N_3528,N_4033);
nor UO_550 (O_550,N_4749,N_4062);
nand UO_551 (O_551,N_2690,N_2918);
nand UO_552 (O_552,N_4624,N_3843);
and UO_553 (O_553,N_4594,N_2513);
nor UO_554 (O_554,N_2789,N_3899);
and UO_555 (O_555,N_3095,N_2511);
nand UO_556 (O_556,N_3156,N_4333);
nand UO_557 (O_557,N_4138,N_3402);
or UO_558 (O_558,N_4242,N_4250);
or UO_559 (O_559,N_4257,N_4214);
nand UO_560 (O_560,N_4291,N_4093);
xnor UO_561 (O_561,N_4799,N_3263);
or UO_562 (O_562,N_4375,N_2888);
or UO_563 (O_563,N_2599,N_3521);
nand UO_564 (O_564,N_4167,N_3913);
nand UO_565 (O_565,N_4533,N_3772);
or UO_566 (O_566,N_3110,N_3482);
nand UO_567 (O_567,N_4081,N_3467);
nand UO_568 (O_568,N_2751,N_4516);
nand UO_569 (O_569,N_2621,N_4815);
nor UO_570 (O_570,N_4159,N_3728);
nor UO_571 (O_571,N_3408,N_4282);
or UO_572 (O_572,N_3014,N_4486);
nor UO_573 (O_573,N_4591,N_2766);
nand UO_574 (O_574,N_4468,N_3184);
nand UO_575 (O_575,N_3018,N_2914);
nand UO_576 (O_576,N_4060,N_3869);
nor UO_577 (O_577,N_4656,N_3656);
nor UO_578 (O_578,N_4663,N_2648);
or UO_579 (O_579,N_3160,N_4072);
nor UO_580 (O_580,N_2580,N_3980);
and UO_581 (O_581,N_4216,N_2740);
or UO_582 (O_582,N_3966,N_3275);
or UO_583 (O_583,N_3596,N_2704);
and UO_584 (O_584,N_4562,N_4561);
or UO_585 (O_585,N_3157,N_3155);
nand UO_586 (O_586,N_3594,N_3055);
or UO_587 (O_587,N_2518,N_4246);
and UO_588 (O_588,N_4899,N_3965);
nand UO_589 (O_589,N_4768,N_3695);
or UO_590 (O_590,N_3836,N_4918);
nor UO_591 (O_591,N_4082,N_4088);
and UO_592 (O_592,N_2967,N_2698);
nor UO_593 (O_593,N_4460,N_4650);
nand UO_594 (O_594,N_3892,N_4275);
nand UO_595 (O_595,N_2878,N_4001);
nor UO_596 (O_596,N_2810,N_4041);
nand UO_597 (O_597,N_4146,N_3524);
nand UO_598 (O_598,N_4614,N_4034);
nand UO_599 (O_599,N_2800,N_3340);
nand UO_600 (O_600,N_2637,N_3813);
nor UO_601 (O_601,N_4579,N_4503);
and UO_602 (O_602,N_4891,N_3815);
nor UO_603 (O_603,N_3117,N_3294);
and UO_604 (O_604,N_3588,N_3863);
or UO_605 (O_605,N_4227,N_3825);
and UO_606 (O_606,N_3822,N_3790);
and UO_607 (O_607,N_4564,N_4973);
and UO_608 (O_608,N_4413,N_3982);
and UO_609 (O_609,N_3783,N_3632);
nor UO_610 (O_610,N_4215,N_2735);
nor UO_611 (O_611,N_3174,N_2893);
nor UO_612 (O_612,N_2656,N_2923);
nand UO_613 (O_613,N_3355,N_4358);
and UO_614 (O_614,N_4785,N_3147);
nand UO_615 (O_615,N_4367,N_3044);
and UO_616 (O_616,N_2883,N_3451);
or UO_617 (O_617,N_4248,N_3726);
nand UO_618 (O_618,N_2572,N_2885);
or UO_619 (O_619,N_4145,N_4035);
or UO_620 (O_620,N_4007,N_3325);
nand UO_621 (O_621,N_3354,N_4336);
and UO_622 (O_622,N_4673,N_4450);
and UO_623 (O_623,N_3693,N_4886);
or UO_624 (O_624,N_4951,N_2609);
nand UO_625 (O_625,N_4801,N_4277);
nand UO_626 (O_626,N_3686,N_3979);
or UO_627 (O_627,N_4995,N_4724);
or UO_628 (O_628,N_3852,N_4560);
or UO_629 (O_629,N_2728,N_4585);
nand UO_630 (O_630,N_3700,N_3606);
nor UO_631 (O_631,N_4647,N_4050);
or UO_632 (O_632,N_4642,N_4004);
nand UO_633 (O_633,N_3073,N_3698);
or UO_634 (O_634,N_4223,N_4849);
and UO_635 (O_635,N_3314,N_4225);
and UO_636 (O_636,N_4786,N_4230);
and UO_637 (O_637,N_2752,N_3477);
and UO_638 (O_638,N_2649,N_4032);
nor UO_639 (O_639,N_4139,N_4295);
nor UO_640 (O_640,N_4871,N_4821);
nand UO_641 (O_641,N_3705,N_4092);
or UO_642 (O_642,N_4878,N_2959);
or UO_643 (O_643,N_2627,N_3526);
nand UO_644 (O_644,N_3602,N_3765);
nor UO_645 (O_645,N_3904,N_2542);
nor UO_646 (O_646,N_3589,N_3976);
nor UO_647 (O_647,N_4865,N_2792);
nand UO_648 (O_648,N_4829,N_2582);
nor UO_649 (O_649,N_3143,N_3874);
or UO_650 (O_650,N_4078,N_3845);
and UO_651 (O_651,N_3015,N_4467);
or UO_652 (O_652,N_3024,N_4508);
nor UO_653 (O_653,N_4604,N_3109);
nand UO_654 (O_654,N_4818,N_2624);
or UO_655 (O_655,N_4892,N_3854);
or UO_656 (O_656,N_4312,N_3654);
nor UO_657 (O_657,N_4622,N_4037);
or UO_658 (O_658,N_4346,N_4727);
nand UO_659 (O_659,N_2717,N_4224);
nand UO_660 (O_660,N_3453,N_2894);
nand UO_661 (O_661,N_3319,N_3361);
nor UO_662 (O_662,N_4820,N_2583);
or UO_663 (O_663,N_2719,N_4351);
and UO_664 (O_664,N_4555,N_3104);
nand UO_665 (O_665,N_4919,N_4188);
nand UO_666 (O_666,N_4186,N_3784);
nor UO_667 (O_667,N_3374,N_3136);
and UO_668 (O_668,N_3301,N_3795);
nor UO_669 (O_669,N_2591,N_4532);
or UO_670 (O_670,N_4451,N_2764);
nand UO_671 (O_671,N_2903,N_3629);
or UO_672 (O_672,N_2593,N_4990);
nor UO_673 (O_673,N_3218,N_4008);
xnor UO_674 (O_674,N_4742,N_3971);
nand UO_675 (O_675,N_4836,N_2650);
or UO_676 (O_676,N_4143,N_3226);
nand UO_677 (O_677,N_4430,N_4496);
or UO_678 (O_678,N_2945,N_3916);
and UO_679 (O_679,N_3494,N_2713);
and UO_680 (O_680,N_4354,N_3950);
nor UO_681 (O_681,N_3691,N_4941);
nand UO_682 (O_682,N_2684,N_3076);
or UO_683 (O_683,N_4959,N_3360);
nor UO_684 (O_684,N_4317,N_4510);
nand UO_685 (O_685,N_4678,N_3753);
nor UO_686 (O_686,N_4412,N_3050);
nor UO_687 (O_687,N_2915,N_3660);
and UO_688 (O_688,N_3002,N_3520);
nor UO_689 (O_689,N_3992,N_2924);
or UO_690 (O_690,N_4180,N_4734);
and UO_691 (O_691,N_4760,N_4751);
nor UO_692 (O_692,N_3945,N_4233);
nand UO_693 (O_693,N_2979,N_3671);
nor UO_694 (O_694,N_3507,N_4024);
or UO_695 (O_695,N_2708,N_4890);
and UO_696 (O_696,N_2994,N_2575);
nor UO_697 (O_697,N_2846,N_4541);
nor UO_698 (O_698,N_3622,N_3991);
xor UO_699 (O_699,N_3491,N_4356);
and UO_700 (O_700,N_2798,N_4694);
nor UO_701 (O_701,N_2976,N_2969);
nor UO_702 (O_702,N_4304,N_4097);
nor UO_703 (O_703,N_2612,N_3911);
xor UO_704 (O_704,N_3499,N_4831);
nand UO_705 (O_705,N_4569,N_3898);
nand UO_706 (O_706,N_2731,N_3555);
or UO_707 (O_707,N_4887,N_3353);
or UO_708 (O_708,N_4229,N_4491);
nand UO_709 (O_709,N_2879,N_2678);
or UO_710 (O_710,N_3099,N_2816);
or UO_711 (O_711,N_2714,N_4232);
nand UO_712 (O_712,N_3903,N_4286);
nor UO_713 (O_713,N_2661,N_3127);
and UO_714 (O_714,N_3233,N_2857);
and UO_715 (O_715,N_3516,N_4162);
xor UO_716 (O_716,N_3064,N_3410);
or UO_717 (O_717,N_3583,N_4206);
or UO_718 (O_718,N_2528,N_2882);
and UO_719 (O_719,N_3636,N_3741);
and UO_720 (O_720,N_3312,N_2990);
nand UO_721 (O_721,N_3446,N_3144);
nand UO_722 (O_722,N_2631,N_4610);
nor UO_723 (O_723,N_4652,N_3937);
nand UO_724 (O_724,N_3430,N_3817);
nor UO_725 (O_725,N_3145,N_3245);
xor UO_726 (O_726,N_3005,N_4212);
and UO_727 (O_727,N_3757,N_2670);
nand UO_728 (O_728,N_4040,N_2746);
or UO_729 (O_729,N_4518,N_3365);
nor UO_730 (O_730,N_3743,N_3958);
nand UO_731 (O_731,N_4728,N_3298);
and UO_732 (O_732,N_3710,N_2765);
nand UO_733 (O_733,N_4913,N_4538);
nand UO_734 (O_734,N_4530,N_2887);
and UO_735 (O_735,N_3527,N_3175);
and UO_736 (O_736,N_2808,N_2515);
or UO_737 (O_737,N_4783,N_4385);
and UO_738 (O_738,N_3664,N_2618);
nor UO_739 (O_739,N_4937,N_4982);
nor UO_740 (O_740,N_4161,N_4401);
nor UO_741 (O_741,N_3134,N_3990);
nor UO_742 (O_742,N_3650,N_4858);
nor UO_743 (O_743,N_4628,N_3744);
nand UO_744 (O_744,N_3435,N_4972);
nand UO_745 (O_745,N_4373,N_4633);
nand UO_746 (O_746,N_4576,N_4597);
nor UO_747 (O_747,N_4341,N_3414);
xnor UO_748 (O_748,N_3216,N_4999);
or UO_749 (O_749,N_4002,N_4581);
nor UO_750 (O_750,N_2892,N_3550);
and UO_751 (O_751,N_4596,N_3999);
or UO_752 (O_752,N_3376,N_2833);
or UO_753 (O_753,N_3957,N_4850);
and UO_754 (O_754,N_3042,N_4586);
nor UO_755 (O_755,N_3900,N_4644);
nor UO_756 (O_756,N_3770,N_3827);
or UO_757 (O_757,N_4376,N_3833);
and UO_758 (O_758,N_2956,N_4618);
nor UO_759 (O_759,N_3567,N_3619);
xor UO_760 (O_760,N_3071,N_4956);
or UO_761 (O_761,N_4517,N_3041);
nand UO_762 (O_762,N_4981,N_2842);
nand UO_763 (O_763,N_4968,N_4776);
and UO_764 (O_764,N_3681,N_4418);
and UO_765 (O_765,N_3339,N_2607);
nor UO_766 (O_766,N_3479,N_4659);
or UO_767 (O_767,N_4268,N_3025);
nand UO_768 (O_768,N_4109,N_4967);
nand UO_769 (O_769,N_4440,N_4695);
or UO_770 (O_770,N_2596,N_4883);
nor UO_771 (O_771,N_4590,N_4643);
nand UO_772 (O_772,N_2613,N_4548);
xnor UO_773 (O_773,N_4482,N_4715);
nor UO_774 (O_774,N_3722,N_3830);
and UO_775 (O_775,N_3419,N_2736);
and UO_776 (O_776,N_2581,N_4409);
and UO_777 (O_777,N_4922,N_4308);
and UO_778 (O_778,N_3519,N_3831);
or UO_779 (O_779,N_4552,N_4204);
and UO_780 (O_780,N_4394,N_4205);
and UO_781 (O_781,N_3395,N_4193);
or UO_782 (O_782,N_3657,N_3313);
and UO_783 (O_783,N_3096,N_3111);
or UO_784 (O_784,N_3856,N_2672);
nor UO_785 (O_785,N_4055,N_4270);
nand UO_786 (O_786,N_3267,N_4738);
nor UO_787 (O_787,N_2876,N_4873);
and UO_788 (O_788,N_4113,N_3694);
nor UO_789 (O_789,N_3078,N_3712);
and UO_790 (O_790,N_4974,N_3798);
or UO_791 (O_791,N_3480,N_3704);
nor UO_792 (O_792,N_4611,N_2819);
and UO_793 (O_793,N_3669,N_4672);
or UO_794 (O_794,N_3239,N_3190);
and UO_795 (O_795,N_3943,N_2839);
or UO_796 (O_796,N_3895,N_4960);
nor UO_797 (O_797,N_3112,N_4593);
or UO_798 (O_798,N_2904,N_3525);
nand UO_799 (O_799,N_3858,N_3476);
nand UO_800 (O_800,N_3369,N_4589);
or UO_801 (O_801,N_4927,N_3266);
or UO_802 (O_802,N_4876,N_3604);
and UO_803 (O_803,N_3738,N_2633);
or UO_804 (O_804,N_4638,N_2788);
nand UO_805 (O_805,N_2932,N_4086);
and UO_806 (O_806,N_2755,N_4507);
or UO_807 (O_807,N_4171,N_3571);
nor UO_808 (O_808,N_3814,N_3536);
nor UO_809 (O_809,N_3885,N_4565);
or UO_810 (O_810,N_2697,N_3461);
nor UO_811 (O_811,N_4741,N_4465);
or UO_812 (O_812,N_3292,N_4946);
nor UO_813 (O_813,N_4522,N_2826);
or UO_814 (O_814,N_4665,N_3949);
xnor UO_815 (O_815,N_4664,N_3423);
and UO_816 (O_816,N_3483,N_2742);
nand UO_817 (O_817,N_4497,N_3926);
nor UO_818 (O_818,N_3713,N_4067);
and UO_819 (O_819,N_4685,N_4407);
nor UO_820 (O_820,N_4063,N_3921);
and UO_821 (O_821,N_4668,N_3303);
nor UO_822 (O_822,N_4896,N_4845);
nand UO_823 (O_823,N_4832,N_2867);
and UO_824 (O_824,N_3993,N_2525);
nand UO_825 (O_825,N_3867,N_4457);
nor UO_826 (O_826,N_3975,N_3821);
nand UO_827 (O_827,N_4901,N_2776);
or UO_828 (O_828,N_3727,N_3307);
nand UO_829 (O_829,N_2869,N_3838);
nand UO_830 (O_830,N_2921,N_4721);
and UO_831 (O_831,N_3236,N_2996);
nand UO_832 (O_832,N_4856,N_3879);
nor UO_833 (O_833,N_2509,N_2644);
and UO_834 (O_834,N_3788,N_3663);
xor UO_835 (O_835,N_4798,N_3385);
nor UO_836 (O_836,N_3717,N_2546);
and UO_837 (O_837,N_4164,N_4219);
or UO_838 (O_838,N_4880,N_4809);
nor UO_839 (O_839,N_4662,N_3329);
and UO_840 (O_840,N_3287,N_3439);
or UO_841 (O_841,N_4859,N_4151);
nand UO_842 (O_842,N_4745,N_2944);
and UO_843 (O_843,N_4361,N_3252);
nor UO_844 (O_844,N_3388,N_3682);
nor UO_845 (O_845,N_4682,N_3750);
and UO_846 (O_846,N_2550,N_3077);
nor UO_847 (O_847,N_2533,N_3468);
xor UO_848 (O_848,N_3922,N_2517);
nand UO_849 (O_849,N_3714,N_3394);
nor UO_850 (O_850,N_2666,N_4605);
or UO_851 (O_851,N_2818,N_3107);
or UO_852 (O_852,N_2787,N_3716);
or UO_853 (O_853,N_4020,N_4737);
nand UO_854 (O_854,N_4448,N_2617);
nor UO_855 (O_855,N_3934,N_3350);
nand UO_856 (O_856,N_3888,N_3649);
or UO_857 (O_857,N_3185,N_4676);
nor UO_858 (O_858,N_2663,N_4743);
nand UO_859 (O_859,N_3400,N_2965);
and UO_860 (O_860,N_3273,N_3225);
nor UO_861 (O_861,N_4332,N_2938);
and UO_862 (O_862,N_4567,N_3647);
or UO_863 (O_863,N_4237,N_4584);
nor UO_864 (O_864,N_3736,N_3333);
nand UO_865 (O_865,N_2664,N_3828);
or UO_866 (O_866,N_3166,N_4005);
nand UO_867 (O_867,N_2998,N_3115);
or UO_868 (O_868,N_3434,N_3952);
or UO_869 (O_869,N_3449,N_4546);
nand UO_870 (O_870,N_4480,N_4399);
and UO_871 (O_871,N_4846,N_2749);
nand UO_872 (O_872,N_3607,N_3009);
nand UO_873 (O_873,N_3418,N_4814);
xnor UO_874 (O_874,N_3377,N_2674);
and UO_875 (O_875,N_3592,N_3214);
nor UO_876 (O_876,N_3623,N_3481);
or UO_877 (O_877,N_4300,N_4030);
and UO_878 (O_878,N_2758,N_4898);
or UO_879 (O_879,N_4039,N_2970);
xor UO_880 (O_880,N_3416,N_4860);
nor UO_881 (O_881,N_2516,N_3090);
nor UO_882 (O_882,N_3877,N_4583);
or UO_883 (O_883,N_2943,N_2529);
nor UO_884 (O_884,N_4686,N_2770);
or UO_885 (O_885,N_3027,N_4302);
and UO_886 (O_886,N_4784,N_4369);
or UO_887 (O_887,N_4787,N_4553);
nand UO_888 (O_888,N_3011,N_2718);
nand UO_889 (O_889,N_4339,N_3552);
and UO_890 (O_890,N_3936,N_3690);
and UO_891 (O_891,N_4352,N_2884);
nor UO_892 (O_892,N_3053,N_3677);
nand UO_893 (O_893,N_2860,N_3584);
or UO_894 (O_894,N_3931,N_4381);
nor UO_895 (O_895,N_2724,N_3908);
and UO_896 (O_896,N_4935,N_3474);
nor UO_897 (O_897,N_4198,N_3182);
or UO_898 (O_898,N_4183,N_4099);
and UO_899 (O_899,N_4843,N_3083);
xnor UO_900 (O_900,N_4667,N_3684);
nor UO_901 (O_901,N_3123,N_2912);
nor UO_902 (O_902,N_3492,N_3642);
or UO_903 (O_903,N_3961,N_3928);
nand UO_904 (O_904,N_4382,N_2538);
nor UO_905 (O_905,N_2573,N_4408);
and UO_906 (O_906,N_2615,N_4209);
nand UO_907 (O_907,N_4243,N_3872);
or UO_908 (O_908,N_4987,N_2577);
and UO_909 (O_909,N_4324,N_3851);
nor UO_910 (O_910,N_4492,N_3465);
and UO_911 (O_911,N_3944,N_4864);
xor UO_912 (O_912,N_3512,N_4386);
or UO_913 (O_913,N_4900,N_3036);
nand UO_914 (O_914,N_4443,N_4329);
and UO_915 (O_915,N_4971,N_3362);
nor UO_916 (O_916,N_4693,N_3518);
and UO_917 (O_917,N_2850,N_3808);
nand UO_918 (O_918,N_4259,N_4736);
nand UO_919 (O_919,N_4107,N_3857);
nor UO_920 (O_920,N_4426,N_4106);
nor UO_921 (O_921,N_4253,N_4371);
nor UO_922 (O_922,N_3920,N_4011);
and UO_923 (O_923,N_4909,N_4110);
nor UO_924 (O_924,N_4707,N_2651);
and UO_925 (O_925,N_2503,N_3792);
or UO_926 (O_926,N_4658,N_4293);
nand UO_927 (O_927,N_2715,N_3100);
nand UO_928 (O_928,N_3687,N_4142);
and UO_929 (O_929,N_4247,N_3052);
nand UO_930 (O_930,N_4174,N_2641);
and UO_931 (O_931,N_2568,N_3092);
or UO_932 (O_932,N_4908,N_3805);
or UO_933 (O_933,N_3739,N_2720);
xnor UO_934 (O_934,N_4405,N_3067);
nor UO_935 (O_935,N_4588,N_2576);
and UO_936 (O_936,N_2757,N_2908);
or UO_937 (O_937,N_3207,N_3680);
nor UO_938 (O_938,N_2753,N_4797);
or UO_939 (O_939,N_4536,N_3553);
nor UO_940 (O_940,N_4903,N_4446);
nand UO_941 (O_941,N_3758,N_3026);
or UO_942 (O_942,N_3674,N_2729);
and UO_943 (O_943,N_3574,N_3124);
nor UO_944 (O_944,N_2563,N_3643);
or UO_945 (O_945,N_3963,N_3178);
or UO_946 (O_946,N_3504,N_3407);
nand UO_947 (O_947,N_2898,N_3907);
nor UO_948 (O_948,N_3358,N_3058);
and UO_949 (O_949,N_2953,N_3539);
nor UO_950 (O_950,N_2606,N_4318);
and UO_951 (O_951,N_2824,N_3514);
and UO_952 (O_952,N_4853,N_3454);
and UO_953 (O_953,N_4986,N_3764);
nand UO_954 (O_954,N_4735,N_4380);
and UO_955 (O_955,N_3135,N_4582);
nand UO_956 (O_956,N_3146,N_3335);
or UO_957 (O_957,N_2966,N_3164);
or UO_958 (O_958,N_4349,N_4520);
or UO_959 (O_959,N_4649,N_4379);
or UO_960 (O_960,N_3131,N_3540);
and UO_961 (O_961,N_4866,N_3403);
or UO_962 (O_962,N_4177,N_3189);
and UO_963 (O_963,N_3087,N_4048);
nand UO_964 (O_964,N_4208,N_3653);
or UO_965 (O_965,N_3320,N_3279);
and UO_966 (O_966,N_4884,N_3409);
nand UO_967 (O_967,N_4669,N_2737);
nand UO_968 (O_968,N_4374,N_3498);
and UO_969 (O_969,N_2999,N_3179);
or UO_970 (O_970,N_3196,N_4800);
xnor UO_971 (O_971,N_4447,N_2917);
xor UO_972 (O_972,N_3530,N_4717);
xnor UO_973 (O_973,N_3161,N_3173);
and UO_974 (O_974,N_3774,N_3620);
or UO_975 (O_975,N_3947,N_4059);
nor UO_976 (O_976,N_4069,N_4953);
nand UO_977 (O_977,N_4823,N_3003);
and UO_978 (O_978,N_3780,N_2658);
nor UO_979 (O_979,N_3995,N_4932);
and UO_980 (O_980,N_4994,N_3864);
nor UO_981 (O_981,N_3973,N_4133);
nor UO_982 (O_982,N_3640,N_3464);
and UO_983 (O_983,N_4752,N_3532);
nand UO_984 (O_984,N_3786,N_4079);
nand UO_985 (O_985,N_3084,N_2936);
and UO_986 (O_986,N_3000,N_2696);
or UO_987 (O_987,N_4251,N_4885);
or UO_988 (O_988,N_3675,N_3511);
and UO_989 (O_989,N_4515,N_3426);
or UO_990 (O_990,N_3031,N_4868);
nor UO_991 (O_991,N_3493,N_3230);
nor UO_992 (O_992,N_4456,N_4028);
nor UO_993 (O_993,N_3281,N_2688);
or UO_994 (O_994,N_4641,N_4940);
nand UO_995 (O_995,N_3939,N_2549);
nor UO_996 (O_996,N_3363,N_3309);
nand UO_997 (O_997,N_4857,N_3165);
nor UO_998 (O_998,N_4363,N_4840);
nand UO_999 (O_999,N_3455,N_4770);
endmodule