module basic_2000_20000_2500_100_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_333,In_1199);
nor U1 (N_1,In_951,In_138);
or U2 (N_2,In_375,In_941);
and U3 (N_3,In_1858,In_1702);
and U4 (N_4,In_757,In_1500);
nand U5 (N_5,In_560,In_1045);
and U6 (N_6,In_632,In_1448);
or U7 (N_7,In_1397,In_249);
or U8 (N_8,In_491,In_82);
nor U9 (N_9,In_1118,In_403);
and U10 (N_10,In_164,In_1785);
nand U11 (N_11,In_1881,In_199);
and U12 (N_12,In_953,In_112);
or U13 (N_13,In_270,In_1366);
or U14 (N_14,In_704,In_1803);
nand U15 (N_15,In_257,In_1699);
or U16 (N_16,In_1498,In_1750);
and U17 (N_17,In_501,In_582);
and U18 (N_18,In_216,In_519);
and U19 (N_19,In_700,In_636);
and U20 (N_20,In_1868,In_1684);
or U21 (N_21,In_1010,In_534);
or U22 (N_22,In_1845,In_324);
nor U23 (N_23,In_931,In_1067);
nand U24 (N_24,In_273,In_424);
nand U25 (N_25,In_1023,In_1089);
nand U26 (N_26,In_597,In_261);
and U27 (N_27,In_398,In_1435);
or U28 (N_28,In_1114,In_1959);
nor U29 (N_29,In_1449,In_1661);
or U30 (N_30,In_774,In_1124);
and U31 (N_31,In_1692,In_1063);
or U32 (N_32,In_127,In_485);
and U33 (N_33,In_605,In_1044);
or U34 (N_34,In_1130,In_940);
and U35 (N_35,In_392,In_440);
or U36 (N_36,In_51,In_1161);
nand U37 (N_37,In_1564,In_6);
and U38 (N_38,In_552,In_1052);
nand U39 (N_39,In_1530,In_1589);
nand U40 (N_40,In_1962,In_1687);
nor U41 (N_41,In_1210,In_1024);
nor U42 (N_42,In_1372,In_1882);
nor U43 (N_43,In_1489,In_683);
nor U44 (N_44,In_1377,In_22);
nand U45 (N_45,In_1009,In_1127);
nand U46 (N_46,In_1221,In_1720);
nor U47 (N_47,In_389,In_1808);
nor U48 (N_48,In_669,In_541);
nand U49 (N_49,In_1745,In_452);
or U50 (N_50,In_1952,In_1918);
or U51 (N_51,In_1636,In_1375);
nand U52 (N_52,In_1618,In_698);
and U53 (N_53,In_83,In_1125);
nand U54 (N_54,In_1176,In_1732);
and U55 (N_55,In_513,In_765);
nand U56 (N_56,In_1439,In_1832);
or U57 (N_57,In_472,In_684);
or U58 (N_58,In_1735,In_1443);
and U59 (N_59,In_1778,In_1656);
and U60 (N_60,In_1517,In_1227);
nand U61 (N_61,In_1809,In_677);
nor U62 (N_62,In_1425,In_337);
or U63 (N_63,In_1966,In_11);
nor U64 (N_64,In_1653,In_1911);
nand U65 (N_65,In_760,In_1115);
nand U66 (N_66,In_1837,In_884);
nor U67 (N_67,In_30,In_253);
and U68 (N_68,In_116,In_1603);
nand U69 (N_69,In_44,In_1463);
and U70 (N_70,In_1766,In_1037);
nor U71 (N_71,In_1050,In_368);
or U72 (N_72,In_807,In_203);
or U73 (N_73,In_500,In_1558);
nand U74 (N_74,In_1036,In_438);
nand U75 (N_75,In_1825,In_716);
nand U76 (N_76,In_359,In_1880);
and U77 (N_77,In_997,In_1040);
nand U78 (N_78,In_497,In_890);
nand U79 (N_79,In_1250,In_531);
nor U80 (N_80,In_746,In_896);
nor U81 (N_81,In_1658,In_1901);
and U82 (N_82,In_1129,In_834);
nor U83 (N_83,In_393,In_153);
and U84 (N_84,In_1597,In_1126);
or U85 (N_85,In_451,In_1823);
nand U86 (N_86,In_955,In_628);
nand U87 (N_87,In_61,In_1925);
and U88 (N_88,In_518,In_1897);
nand U89 (N_89,In_207,In_275);
and U90 (N_90,In_1613,In_1200);
nor U91 (N_91,In_1865,In_1566);
xnor U92 (N_92,In_95,In_178);
or U93 (N_93,In_1693,In_307);
nor U94 (N_94,In_788,In_1524);
or U95 (N_95,In_544,In_606);
or U96 (N_96,In_1312,In_37);
nand U97 (N_97,In_1593,In_1864);
or U98 (N_98,In_1514,In_868);
or U99 (N_99,In_1828,In_35);
or U100 (N_100,In_991,In_150);
xnor U101 (N_101,In_1098,In_664);
nand U102 (N_102,In_1112,In_1947);
and U103 (N_103,In_295,In_1359);
nand U104 (N_104,In_883,In_1565);
nor U105 (N_105,In_1331,In_526);
nor U106 (N_106,In_866,In_121);
and U107 (N_107,In_1777,In_355);
and U108 (N_108,In_743,In_803);
or U109 (N_109,In_1348,In_292);
and U110 (N_110,In_1384,In_961);
nand U111 (N_111,In_1921,In_1937);
or U112 (N_112,In_1756,In_1602);
nor U113 (N_113,In_197,In_291);
nand U114 (N_114,In_1401,In_33);
nor U115 (N_115,In_1343,In_1800);
nand U116 (N_116,In_1427,In_434);
nor U117 (N_117,In_901,In_902);
or U118 (N_118,In_1839,In_1477);
and U119 (N_119,In_1159,In_1493);
nor U120 (N_120,In_767,In_137);
and U121 (N_121,In_1540,In_1434);
and U122 (N_122,In_367,In_420);
nor U123 (N_123,In_120,In_283);
nor U124 (N_124,In_1400,In_742);
and U125 (N_125,In_692,In_65);
and U126 (N_126,In_512,In_19);
and U127 (N_127,In_1726,In_0);
or U128 (N_128,In_1334,In_1932);
or U129 (N_129,In_565,In_1383);
nand U130 (N_130,In_694,In_1926);
nand U131 (N_131,In_1406,In_1108);
nor U132 (N_132,In_332,In_924);
and U133 (N_133,In_483,In_1103);
nor U134 (N_134,In_448,In_668);
nor U135 (N_135,In_272,In_1177);
nor U136 (N_136,In_1607,In_509);
or U137 (N_137,In_1629,In_528);
or U138 (N_138,In_1355,In_461);
or U139 (N_139,In_111,In_894);
nor U140 (N_140,In_1347,In_613);
or U141 (N_141,In_1888,In_658);
or U142 (N_142,In_1578,In_561);
or U143 (N_143,In_1550,In_857);
and U144 (N_144,In_1190,In_973);
nor U145 (N_145,In_262,In_506);
nor U146 (N_146,In_1934,In_1549);
and U147 (N_147,In_487,In_980);
nor U148 (N_148,In_564,In_1122);
nand U149 (N_149,In_627,In_263);
or U150 (N_150,In_1584,In_917);
nand U151 (N_151,In_809,In_622);
and U152 (N_152,In_520,In_1806);
and U153 (N_153,In_1277,In_688);
and U154 (N_154,In_1396,In_614);
nor U155 (N_155,In_1614,In_192);
nand U156 (N_156,In_1665,In_66);
nand U157 (N_157,In_1407,In_749);
or U158 (N_158,In_1132,In_831);
or U159 (N_159,In_390,In_816);
and U160 (N_160,In_828,In_871);
or U161 (N_161,In_149,In_899);
and U162 (N_162,In_1314,In_1993);
xnor U163 (N_163,In_1510,In_984);
nor U164 (N_164,In_1626,In_1963);
and U165 (N_165,In_405,In_869);
or U166 (N_166,In_504,In_1622);
and U167 (N_167,In_1026,In_388);
nor U168 (N_168,In_486,In_195);
and U169 (N_169,In_130,In_629);
nor U170 (N_170,In_1446,In_673);
or U171 (N_171,In_1090,In_251);
or U172 (N_172,In_932,In_1546);
and U173 (N_173,In_1150,In_570);
nand U174 (N_174,In_1499,In_57);
nor U175 (N_175,In_576,In_1928);
and U176 (N_176,In_959,In_2);
nand U177 (N_177,In_719,In_1513);
nand U178 (N_178,In_1765,In_758);
nand U179 (N_179,In_267,In_1541);
nand U180 (N_180,In_260,In_342);
and U181 (N_181,In_670,In_1297);
nor U182 (N_182,In_1672,In_1251);
and U183 (N_183,In_769,In_1450);
or U184 (N_184,In_558,In_1066);
nor U185 (N_185,In_667,In_569);
nand U186 (N_186,In_1344,In_1688);
or U187 (N_187,In_1955,In_986);
nand U188 (N_188,In_1013,In_235);
or U189 (N_189,In_588,In_770);
nor U190 (N_190,In_1011,In_1872);
nand U191 (N_191,In_1571,In_1781);
nand U192 (N_192,In_1568,In_551);
and U193 (N_193,In_94,In_995);
or U194 (N_194,In_1902,In_1751);
and U195 (N_195,In_312,In_649);
nand U196 (N_196,In_289,In_939);
or U197 (N_197,In_1907,In_4);
nand U198 (N_198,In_43,In_876);
nand U199 (N_199,In_563,In_1031);
and U200 (N_200,In_1264,In_1491);
nor U201 (N_201,In_1748,In_1582);
or U202 (N_202,In_1877,In_641);
or U203 (N_203,In_1790,In_1943);
nand U204 (N_204,In_258,In_1674);
nand U205 (N_205,In_354,In_1849);
nand U206 (N_206,In_254,In_1638);
or U207 (N_207,In_1906,In_971);
or U208 (N_208,In_1392,In_1095);
nor U209 (N_209,N_14,In_1245);
nand U210 (N_210,In_1810,In_1904);
nor U211 (N_211,In_1410,In_1753);
or U212 (N_212,N_44,In_1285);
and U213 (N_213,N_73,In_993);
and U214 (N_214,In_1276,In_453);
or U215 (N_215,In_812,In_1157);
nor U216 (N_216,In_1739,In_1058);
and U217 (N_217,In_233,In_888);
nand U218 (N_218,In_1552,In_1172);
nand U219 (N_219,In_1079,N_56);
nand U220 (N_220,In_287,In_1005);
nor U221 (N_221,In_234,In_1447);
nand U222 (N_222,In_717,In_1283);
and U223 (N_223,In_1681,In_1795);
nor U224 (N_224,In_274,In_1194);
nand U225 (N_225,In_1203,In_1000);
or U226 (N_226,In_341,N_196);
nand U227 (N_227,N_67,In_1957);
or U228 (N_228,In_416,N_30);
nand U229 (N_229,In_1497,N_178);
nor U230 (N_230,In_1246,In_557);
and U231 (N_231,In_413,In_1835);
and U232 (N_232,In_1639,In_193);
nor U233 (N_233,In_248,In_1935);
nand U234 (N_234,In_1265,In_180);
nand U235 (N_235,In_1861,In_1744);
nor U236 (N_236,In_376,In_1544);
and U237 (N_237,In_994,In_5);
or U238 (N_238,In_1296,In_1700);
nand U239 (N_239,In_1951,In_1398);
and U240 (N_240,In_1923,In_598);
xor U241 (N_241,N_93,In_52);
and U242 (N_242,In_278,In_71);
nand U243 (N_243,In_1254,In_929);
nand U244 (N_244,In_173,In_678);
and U245 (N_245,In_1949,N_89);
nor U246 (N_246,In_567,In_826);
and U247 (N_247,In_1174,In_323);
xor U248 (N_248,In_977,N_177);
nor U249 (N_249,In_1082,In_1273);
nor U250 (N_250,In_800,In_1426);
or U251 (N_251,In_1736,In_962);
nand U252 (N_252,In_439,In_425);
nand U253 (N_253,In_1402,In_517);
and U254 (N_254,In_1168,N_39);
nor U255 (N_255,In_1848,In_615);
or U256 (N_256,In_1721,In_877);
nand U257 (N_257,N_22,In_860);
and U258 (N_258,In_837,In_1152);
nand U259 (N_259,In_1887,In_1535);
nand U260 (N_260,In_1110,In_1038);
nand U261 (N_261,In_1624,In_1315);
nand U262 (N_262,In_881,In_1752);
nand U263 (N_263,In_1562,In_802);
and U264 (N_264,In_1631,In_1214);
and U265 (N_265,In_1671,In_1080);
and U266 (N_266,In_1743,In_1512);
and U267 (N_267,In_1836,N_87);
nand U268 (N_268,In_1056,In_1831);
nand U269 (N_269,In_1116,In_456);
nor U270 (N_270,In_1337,In_643);
nor U271 (N_271,In_352,In_446);
nor U272 (N_272,In_490,In_737);
and U273 (N_273,In_1465,N_20);
nand U274 (N_274,N_48,In_10);
and U275 (N_275,In_417,In_714);
nand U276 (N_276,In_726,In_1370);
and U277 (N_277,In_177,In_470);
or U278 (N_278,In_1418,In_620);
nand U279 (N_279,In_1290,In_1456);
nor U280 (N_280,In_194,In_1302);
and U281 (N_281,In_1764,In_1061);
or U282 (N_282,In_780,In_387);
or U283 (N_283,In_469,In_1300);
nand U284 (N_284,In_591,In_475);
xnor U285 (N_285,In_1776,In_1780);
or U286 (N_286,In_1812,In_1249);
and U287 (N_287,In_1455,In_804);
or U288 (N_288,In_1642,In_1022);
nor U289 (N_289,In_524,In_176);
nand U290 (N_290,N_122,In_1087);
nand U291 (N_291,In_1155,In_1076);
nand U292 (N_292,In_1797,In_623);
nand U293 (N_293,In_841,In_1595);
nor U294 (N_294,In_1704,In_1912);
and U295 (N_295,In_1452,In_1395);
nand U296 (N_296,In_1802,In_1521);
nor U297 (N_297,In_1259,In_872);
or U298 (N_298,In_1649,N_144);
or U299 (N_299,In_1824,In_1468);
and U300 (N_300,In_886,In_1223);
nand U301 (N_301,In_1071,In_1545);
nor U302 (N_302,In_1866,In_1917);
nand U303 (N_303,In_1585,In_155);
or U304 (N_304,N_140,In_1444);
nand U305 (N_305,In_166,In_695);
and U306 (N_306,In_1680,In_648);
and U307 (N_307,In_706,In_1092);
or U308 (N_308,In_157,In_383);
nand U309 (N_309,In_970,N_86);
nor U310 (N_310,In_708,In_402);
nand U311 (N_311,In_1445,In_1184);
nand U312 (N_312,In_1519,In_1754);
or U313 (N_313,In_230,N_54);
nand U314 (N_314,In_1569,N_98);
nand U315 (N_315,In_436,N_24);
and U316 (N_316,In_1718,In_1160);
and U317 (N_317,In_1588,In_482);
and U318 (N_318,In_1958,In_795);
nand U319 (N_319,In_1403,In_1027);
nor U320 (N_320,In_1035,In_1784);
nor U321 (N_321,N_129,N_37);
or U322 (N_322,In_1263,In_619);
nand U323 (N_323,In_1454,N_92);
nand U324 (N_324,In_599,In_1244);
nand U325 (N_325,In_1387,In_404);
and U326 (N_326,In_1113,In_1716);
or U327 (N_327,In_1804,In_1710);
or U328 (N_328,In_1728,In_1580);
nand U329 (N_329,In_947,In_1218);
and U330 (N_330,In_93,In_1529);
or U331 (N_331,In_1528,In_1637);
nand U332 (N_332,In_522,In_1205);
nor U333 (N_333,In_589,In_1581);
or U334 (N_334,In_607,In_1978);
nor U335 (N_335,In_555,In_573);
or U336 (N_336,In_912,In_186);
and U337 (N_337,In_1025,In_1526);
and U338 (N_338,N_4,In_170);
or U339 (N_339,In_386,In_593);
or U340 (N_340,In_1977,In_1303);
nor U341 (N_341,N_104,In_1775);
xnor U342 (N_342,In_1441,In_1652);
nor U343 (N_343,In_709,In_1749);
nor U344 (N_344,N_99,N_74);
or U345 (N_345,In_992,In_1431);
nand U346 (N_346,In_271,In_748);
or U347 (N_347,In_546,In_185);
nand U348 (N_348,In_679,In_1274);
nand U349 (N_349,In_1635,In_1191);
or U350 (N_350,In_1999,In_999);
and U351 (N_351,In_1729,In_1247);
nor U352 (N_352,N_29,N_31);
nor U353 (N_353,In_514,In_210);
and U354 (N_354,In_1480,In_1028);
or U355 (N_355,In_1818,In_1979);
or U356 (N_356,In_1326,In_447);
or U357 (N_357,In_1253,In_1292);
nand U358 (N_358,In_1148,In_934);
nor U359 (N_359,In_844,In_987);
and U360 (N_360,In_1547,In_1320);
nand U361 (N_361,In_1863,In_1207);
nor U362 (N_362,In_1890,In_712);
nor U363 (N_363,In_479,In_204);
nor U364 (N_364,In_823,In_922);
and U365 (N_365,In_73,In_601);
nor U366 (N_366,In_1504,In_60);
nand U367 (N_367,In_460,In_1922);
nor U368 (N_368,In_846,In_152);
xnor U369 (N_369,N_84,In_1120);
nor U370 (N_370,In_1295,In_1442);
and U371 (N_371,In_321,In_1985);
nand U372 (N_372,In_630,In_1936);
nor U373 (N_373,In_1717,In_554);
nand U374 (N_374,In_406,In_1596);
nor U375 (N_375,In_1733,In_330);
or U376 (N_376,In_1536,In_960);
nand U377 (N_377,In_175,In_445);
nand U378 (N_378,In_1931,In_384);
nand U379 (N_379,In_1057,In_1807);
nand U380 (N_380,In_1991,In_63);
and U381 (N_381,In_412,In_699);
nand U382 (N_382,In_887,In_721);
nand U383 (N_383,In_1423,In_1826);
nand U384 (N_384,In_1843,In_1942);
or U385 (N_385,In_1206,In_1876);
or U386 (N_386,In_820,In_768);
nand U387 (N_387,N_28,N_157);
or U388 (N_388,In_1859,In_553);
and U389 (N_389,In_167,In_1121);
nor U390 (N_390,In_243,In_28);
nor U391 (N_391,In_1829,In_42);
and U392 (N_392,N_168,In_1424);
or U393 (N_393,In_227,In_676);
xnor U394 (N_394,N_158,In_935);
nor U395 (N_395,In_1678,In_1973);
and U396 (N_396,In_1053,In_1185);
nor U397 (N_397,N_132,In_1019);
and U398 (N_398,In_783,In_1870);
nor U399 (N_399,In_1988,In_133);
nor U400 (N_400,In_15,In_1644);
nand U401 (N_401,N_221,In_1034);
or U402 (N_402,N_125,In_1106);
or U403 (N_403,In_895,In_1457);
or U404 (N_404,In_1123,In_603);
or U405 (N_405,In_1175,In_981);
nor U406 (N_406,N_330,In_1767);
and U407 (N_407,In_1987,In_818);
or U408 (N_408,In_313,In_1511);
nor U409 (N_409,In_1919,In_728);
or U410 (N_410,In_1712,N_23);
or U411 (N_411,In_1760,In_1628);
or U412 (N_412,In_331,In_1078);
and U413 (N_413,In_1871,In_550);
and U414 (N_414,In_715,In_1081);
and U415 (N_415,In_1892,N_10);
nor U416 (N_416,In_1553,In_1724);
nor U417 (N_417,In_801,N_96);
and U418 (N_418,In_646,In_1946);
nand U419 (N_419,In_1586,In_724);
or U420 (N_420,In_602,In_31);
and U421 (N_421,N_166,In_1139);
or U422 (N_422,N_211,In_55);
and U423 (N_423,In_1388,In_642);
nor U424 (N_424,In_1968,N_11);
and U425 (N_425,N_199,In_224);
or U426 (N_426,N_66,In_870);
or U427 (N_427,In_755,In_1091);
nand U428 (N_428,In_104,N_113);
or U429 (N_429,In_725,N_285);
or U430 (N_430,N_343,N_128);
or U431 (N_431,In_179,In_1771);
nor U432 (N_432,In_824,In_798);
nand U433 (N_433,In_335,In_781);
and U434 (N_434,In_741,N_234);
nor U435 (N_435,In_1611,In_282);
nand U436 (N_436,In_1117,N_250);
nand U437 (N_437,In_1660,In_1181);
or U438 (N_438,In_1576,In_1021);
and U439 (N_439,N_161,N_272);
or U440 (N_440,In_1014,In_1233);
nand U441 (N_441,N_218,In_653);
nor U442 (N_442,N_340,N_154);
and U443 (N_443,In_893,In_577);
or U444 (N_444,In_1099,In_1989);
nand U445 (N_445,In_1186,In_1670);
nor U446 (N_446,N_85,N_7);
nand U447 (N_447,In_1311,In_488);
nor U448 (N_448,In_1041,In_911);
or U449 (N_449,In_85,In_1408);
nand U450 (N_450,In_1619,In_1088);
nand U451 (N_451,N_38,In_650);
nand U452 (N_452,In_1703,In_586);
nor U453 (N_453,In_1758,In_1983);
nand U454 (N_454,In_508,N_282);
or U455 (N_455,In_1248,In_1339);
nand U456 (N_456,In_139,In_1953);
and U457 (N_457,N_296,In_20);
or U458 (N_458,N_136,In_399);
nand U459 (N_459,In_891,In_1503);
nand U460 (N_460,In_1630,N_325);
nand U461 (N_461,In_115,N_299);
nor U462 (N_462,In_505,In_422);
and U463 (N_463,N_171,N_249);
or U464 (N_464,In_1533,In_495);
nand U465 (N_465,N_246,In_1055);
nor U466 (N_466,N_328,In_744);
nand U467 (N_467,In_1062,In_381);
or U468 (N_468,In_240,N_215);
nand U469 (N_469,In_1461,N_97);
nor U470 (N_470,In_1460,N_333);
nand U471 (N_471,In_494,In_1834);
xnor U472 (N_472,In_172,In_808);
nor U473 (N_473,In_151,In_53);
nor U474 (N_474,In_1505,In_753);
or U475 (N_475,N_5,In_1008);
nor U476 (N_476,In_1616,In_1365);
and U477 (N_477,In_1275,In_183);
or U478 (N_478,In_229,N_180);
and U479 (N_479,In_1234,In_759);
nand U480 (N_480,In_1830,N_124);
nor U481 (N_481,In_621,In_1084);
or U482 (N_482,In_1811,In_1896);
nand U483 (N_483,In_1501,In_815);
nor U484 (N_484,In_228,In_898);
nor U485 (N_485,N_191,In_1663);
nor U486 (N_486,In_1015,In_735);
nor U487 (N_487,N_256,In_366);
nand U488 (N_488,In_1484,In_1255);
nor U489 (N_489,In_1697,N_317);
nand U490 (N_490,In_1142,In_503);
nand U491 (N_491,In_635,In_372);
nand U492 (N_492,In_1770,N_137);
nand U493 (N_493,In_640,In_1662);
or U494 (N_494,N_220,In_255);
nor U495 (N_495,In_435,In_400);
nand U496 (N_496,In_574,In_1235);
nand U497 (N_497,In_1007,In_1490);
nand U498 (N_498,In_1419,In_382);
and U499 (N_499,In_1039,In_819);
nand U500 (N_500,N_78,In_1133);
or U501 (N_501,N_352,In_1945);
and U502 (N_502,In_1371,In_222);
nor U503 (N_503,In_1154,In_1385);
nor U504 (N_504,In_1363,In_1908);
nor U505 (N_505,In_1137,In_410);
nand U506 (N_506,In_1669,In_1451);
or U507 (N_507,In_1787,In_1166);
nand U508 (N_508,N_135,In_1518);
nand U509 (N_509,N_279,N_393);
nand U510 (N_510,In_1197,In_1100);
nor U511 (N_511,N_359,In_1675);
and U512 (N_512,N_72,In_1494);
nor U513 (N_513,In_429,In_1466);
nand U514 (N_514,In_739,In_1412);
nor U515 (N_515,In_1373,In_976);
and U516 (N_516,In_548,N_287);
or U517 (N_517,In_1969,In_459);
and U518 (N_518,N_155,N_310);
and U519 (N_519,In_1594,In_1379);
nand U520 (N_520,In_880,N_43);
nor U521 (N_521,In_566,In_1575);
or U522 (N_522,In_590,N_3);
nand U523 (N_523,In_1266,In_1085);
nor U524 (N_524,N_71,N_255);
or U525 (N_525,In_785,In_101);
or U526 (N_526,In_1163,In_122);
and U527 (N_527,In_1689,In_1180);
nor U528 (N_528,In_1643,In_1543);
and U529 (N_529,N_120,In_849);
or U530 (N_530,N_207,In_200);
nand U531 (N_531,In_225,In_533);
nor U532 (N_532,In_62,In_1984);
nand U533 (N_533,In_1722,In_1228);
or U534 (N_534,In_421,In_1042);
nand U535 (N_535,In_191,In_1668);
or U536 (N_536,N_281,N_275);
nand U537 (N_537,In_1289,In_297);
and U538 (N_538,In_1757,In_1573);
and U539 (N_539,N_36,N_311);
or U540 (N_540,In_786,In_1413);
nor U541 (N_541,In_102,N_111);
nand U542 (N_542,N_134,N_312);
or U543 (N_543,In_1996,In_1920);
and U544 (N_544,N_286,In_90);
nor U545 (N_545,In_845,In_1539);
or U546 (N_546,In_49,In_587);
or U547 (N_547,In_99,In_691);
nor U548 (N_548,N_379,In_545);
nand U549 (N_549,In_266,In_1299);
nor U550 (N_550,N_60,In_928);
or U551 (N_551,In_1216,In_1182);
and U552 (N_552,In_762,In_1915);
nand U553 (N_553,In_1714,N_100);
or U554 (N_554,In_697,In_1682);
nand U555 (N_555,In_1734,In_1131);
nand U556 (N_556,In_1691,In_693);
nand U557 (N_557,In_1873,In_827);
nand U558 (N_558,In_1428,N_110);
and U559 (N_559,In_1349,In_515);
nor U560 (N_560,In_308,N_19);
or U561 (N_561,In_1939,In_779);
or U562 (N_562,In_415,In_1261);
and U563 (N_563,In_465,In_1475);
nand U564 (N_564,In_1236,N_318);
nand U565 (N_565,In_680,N_50);
or U566 (N_566,In_426,In_1229);
nor U567 (N_567,N_105,In_1507);
nor U568 (N_568,In_1138,In_1531);
nand U569 (N_569,N_130,N_169);
and U570 (N_570,In_1833,In_131);
nand U571 (N_571,In_147,In_219);
and U572 (N_572,N_175,In_723);
or U573 (N_573,N_152,In_954);
and U574 (N_574,In_1532,N_308);
or U575 (N_575,In_364,In_361);
nor U576 (N_576,In_1226,In_408);
or U577 (N_577,In_1791,In_764);
or U578 (N_578,In_75,In_1621);
nand U579 (N_579,N_387,N_61);
or U580 (N_580,In_1762,In_580);
or U581 (N_581,In_978,In_832);
and U582 (N_582,In_540,N_159);
nand U583 (N_583,In_1209,In_536);
or U584 (N_584,In_362,N_248);
nand U585 (N_585,N_254,In_1198);
xor U586 (N_586,In_1559,N_226);
nor U587 (N_587,In_279,In_1313);
and U588 (N_588,In_1632,N_358);
nor U589 (N_589,In_281,In_1794);
nor U590 (N_590,In_1128,In_858);
and U591 (N_591,N_264,In_821);
nor U592 (N_592,N_244,In_1213);
and U593 (N_593,In_1525,In_1633);
or U594 (N_594,In_80,In_686);
or U595 (N_595,In_1738,In_437);
or U596 (N_596,In_68,In_610);
nor U597 (N_597,In_326,In_1354);
nor U598 (N_598,In_936,In_238);
nand U599 (N_599,In_156,In_1459);
and U600 (N_600,In_1048,In_455);
or U601 (N_601,In_1980,N_415);
and U602 (N_602,In_1792,In_162);
and U603 (N_603,In_209,In_1879);
nor U604 (N_604,In_276,In_12);
and U605 (N_605,N_294,In_1686);
nor U606 (N_606,N_228,N_460);
or U607 (N_607,N_153,In_146);
and U608 (N_608,In_395,In_198);
nor U609 (N_609,In_752,In_750);
or U610 (N_610,N_320,N_504);
and U611 (N_611,N_142,N_107);
and U612 (N_612,In_67,In_1258);
and U613 (N_613,In_659,In_1737);
nor U614 (N_614,In_579,In_1335);
or U615 (N_615,In_1913,N_499);
or U616 (N_616,In_1093,In_696);
and U617 (N_617,In_1353,In_1308);
nand U618 (N_618,In_612,In_662);
or U619 (N_619,N_362,In_1158);
nor U620 (N_620,In_1886,N_558);
or U621 (N_621,In_1620,N_344);
xnor U622 (N_622,N_204,In_1232);
nand U623 (N_623,In_1974,In_96);
nor U624 (N_624,N_446,In_1740);
or U625 (N_625,In_637,In_609);
xor U626 (N_626,In_107,In_1288);
nor U627 (N_627,In_1970,N_420);
nor U628 (N_628,N_469,N_465);
or U629 (N_629,In_805,In_378);
or U630 (N_630,In_983,In_882);
nand U631 (N_631,N_165,In_1574);
and U632 (N_632,In_731,In_1927);
nor U633 (N_633,In_908,N_569);
or U634 (N_634,N_193,In_1195);
or U635 (N_635,In_1215,N_592);
or U636 (N_636,N_350,In_1485);
nand U637 (N_637,In_474,In_1995);
or U638 (N_638,In_1690,N_298);
nand U639 (N_639,In_41,In_1317);
nor U640 (N_640,In_1583,N_450);
nor U641 (N_641,N_265,In_740);
and U642 (N_642,In_1471,N_598);
nor U643 (N_643,N_581,In_1875);
and U644 (N_644,N_75,In_1143);
nand U645 (N_645,N_479,In_1998);
or U646 (N_646,In_915,N_173);
xnor U647 (N_647,N_35,In_290);
nor U648 (N_648,In_1905,N_188);
nand U649 (N_649,In_1075,N_160);
or U650 (N_650,N_554,In_559);
and U651 (N_651,In_47,N_456);
nand U652 (N_652,In_1242,In_318);
nand U653 (N_653,N_561,In_427);
nor U654 (N_654,In_1914,In_1074);
nor U655 (N_655,In_604,In_1049);
nor U656 (N_656,In_879,N_412);
or U657 (N_657,In_1679,In_710);
and U658 (N_658,In_431,In_1072);
or U659 (N_659,In_373,In_1298);
or U660 (N_660,N_502,N_363);
or U661 (N_661,In_1965,N_490);
or U662 (N_662,In_856,N_295);
and U663 (N_663,In_1202,In_1358);
nand U664 (N_664,In_1789,In_797);
nand U665 (N_665,In_863,N_46);
nand U666 (N_666,N_52,N_183);
nor U667 (N_667,N_300,In_791);
nand U668 (N_668,In_206,In_300);
or U669 (N_669,N_205,In_1083);
nor U670 (N_670,In_409,In_1241);
nor U671 (N_671,In_159,In_892);
nand U672 (N_672,In_288,N_427);
or U673 (N_673,In_223,In_1600);
and U674 (N_674,In_631,N_94);
nand U675 (N_675,N_219,In_1319);
nand U676 (N_676,N_476,In_1432);
nand U677 (N_677,In_910,In_1924);
and U678 (N_678,N_148,In_1799);
or U679 (N_679,N_366,In_1271);
and U680 (N_680,N_506,N_432);
and U681 (N_681,In_655,In_813);
nor U682 (N_682,In_1369,In_45);
and U683 (N_683,N_579,In_1956);
nor U684 (N_684,In_1004,In_493);
nand U685 (N_685,In_1715,In_867);
nand U686 (N_686,N_8,In_1891);
or U687 (N_687,In_163,In_1307);
or U688 (N_688,In_1102,In_796);
and U689 (N_689,N_192,N_95);
nand U690 (N_690,In_1860,N_118);
nand U691 (N_691,In_1192,N_372);
nand U692 (N_692,In_69,In_143);
and U693 (N_693,N_497,In_1851);
or U694 (N_694,N_437,In_507);
nor U695 (N_695,In_299,In_1393);
or U696 (N_696,N_331,N_356);
or U697 (N_697,In_1262,In_1814);
nand U698 (N_698,N_537,In_701);
nand U699 (N_699,In_428,In_1646);
nor U700 (N_700,In_345,In_990);
nand U701 (N_701,In_1857,N_1);
or U702 (N_702,N_464,In_1606);
and U703 (N_703,N_408,In_1030);
and U704 (N_704,N_447,In_718);
or U705 (N_705,In_161,In_916);
nand U706 (N_706,In_411,In_1847);
nand U707 (N_707,N_538,In_773);
or U708 (N_708,In_1170,In_889);
and U709 (N_709,N_334,In_1793);
and U710 (N_710,N_293,N_319);
and U711 (N_711,In_571,In_1479);
nor U712 (N_712,In_1960,In_184);
nor U713 (N_713,N_543,In_1361);
nor U714 (N_714,N_505,In_734);
nand U715 (N_715,N_131,N_401);
nor U716 (N_716,In_556,N_58);
or U717 (N_717,N_351,In_148);
nor U718 (N_718,N_461,In_1779);
or U719 (N_719,In_242,In_141);
nand U720 (N_720,In_454,In_705);
nand U721 (N_721,In_1537,N_562);
nor U722 (N_722,N_565,N_512);
or U723 (N_723,In_963,In_1805);
or U724 (N_724,N_174,In_100);
nor U725 (N_725,N_227,In_1788);
nor U726 (N_726,N_108,In_322);
nor U727 (N_727,In_284,In_918);
nor U728 (N_728,In_1367,N_315);
and U729 (N_729,In_1323,In_1405);
or U730 (N_730,In_106,N_283);
and U731 (N_731,In_1601,N_487);
xor U732 (N_732,In_124,In_1225);
or U733 (N_733,N_515,In_1201);
and U734 (N_734,In_1217,In_77);
nor U735 (N_735,N_377,In_1554);
or U736 (N_736,In_1755,In_1874);
and U737 (N_737,N_466,N_594);
nor U738 (N_738,N_449,In_369);
or U739 (N_739,N_45,In_268);
nand U740 (N_740,In_1436,In_1212);
and U741 (N_741,N_590,In_511);
xor U742 (N_742,In_656,In_989);
or U743 (N_743,N_302,In_674);
nor U744 (N_744,In_1430,In_1272);
nand U745 (N_745,In_1827,In_72);
nor U746 (N_746,In_1815,N_585);
or U747 (N_747,In_1104,In_29);
nand U748 (N_748,N_151,N_489);
nor U749 (N_749,N_518,In_1321);
nand U750 (N_750,N_326,N_455);
nor U751 (N_751,N_309,In_498);
nor U752 (N_752,N_521,In_1086);
nor U753 (N_753,N_520,In_394);
or U754 (N_754,In_1654,In_904);
nor U755 (N_755,In_861,In_938);
or U756 (N_756,In_958,N_445);
and U757 (N_757,In_158,In_1409);
or U758 (N_758,In_1774,N_259);
nor U759 (N_759,In_1193,N_402);
or U760 (N_760,In_532,N_540);
nand U761 (N_761,In_651,N_493);
or U762 (N_762,N_414,In_1281);
or U763 (N_763,In_317,In_1310);
or U764 (N_764,In_1096,In_232);
or U765 (N_765,N_77,N_482);
and U766 (N_766,In_1470,N_17);
nor U767 (N_767,In_923,In_97);
nand U768 (N_768,In_160,In_1356);
nand U769 (N_769,In_1474,In_720);
nand U770 (N_770,In_1910,In_1153);
and U771 (N_771,N_430,N_365);
and U772 (N_772,N_307,In_481);
nand U773 (N_773,N_398,In_523);
or U774 (N_774,In_21,In_1869);
nor U775 (N_775,In_1659,In_663);
or U776 (N_776,In_423,In_1059);
nor U777 (N_777,N_212,In_771);
and U778 (N_778,In_1741,N_405);
and U779 (N_779,N_470,In_854);
and U780 (N_780,In_1898,In_660);
or U781 (N_781,N_202,In_1136);
nand U782 (N_782,In_1842,In_1577);
nand U783 (N_783,In_1464,In_169);
or U784 (N_784,In_873,N_322);
nand U785 (N_785,In_118,In_7);
nor U786 (N_786,In_933,In_1240);
and U787 (N_787,N_306,N_532);
nor U788 (N_788,In_1768,In_325);
and U789 (N_789,N_480,N_399);
or U790 (N_790,N_103,In_205);
nor U791 (N_791,N_556,N_478);
nand U792 (N_792,In_638,In_259);
nand U793 (N_793,In_1472,In_967);
nor U794 (N_794,N_568,In_754);
nor U795 (N_795,In_356,N_203);
and U796 (N_796,In_449,In_154);
and U797 (N_797,N_126,In_126);
or U798 (N_798,In_92,In_778);
and U799 (N_799,N_115,In_1421);
or U800 (N_800,In_624,N_752);
and U801 (N_801,In_626,N_225);
and U802 (N_802,N_624,N_34);
or U803 (N_803,In_294,In_1516);
and U804 (N_804,In_1486,In_365);
nor U805 (N_805,N_785,In_982);
nand U806 (N_806,In_1330,In_952);
and U807 (N_807,N_467,In_329);
nor U808 (N_808,N_503,N_648);
nor U809 (N_809,N_342,In_1012);
and U810 (N_810,In_1390,N_566);
nand U811 (N_811,In_314,N_548);
or U812 (N_812,N_726,N_324);
nor U813 (N_813,In_442,N_637);
or U814 (N_814,N_245,N_457);
nor U815 (N_815,In_231,In_91);
nor U816 (N_816,N_440,In_23);
and U817 (N_817,In_1961,In_123);
or U818 (N_818,In_1382,In_1481);
and U819 (N_819,N_710,N_507);
or U820 (N_820,N_172,N_607);
nand U821 (N_821,In_1708,In_1929);
nand U822 (N_822,In_1967,In_1705);
or U823 (N_823,In_1840,In_1551);
or U824 (N_824,N_49,N_787);
nand U825 (N_825,N_410,In_864);
and U826 (N_826,In_202,In_966);
or U827 (N_827,N_719,N_263);
nor U828 (N_828,In_1817,In_969);
nand U829 (N_829,In_1077,In_1651);
nor U830 (N_830,In_1,In_1701);
and U831 (N_831,N_236,In_657);
and U832 (N_832,In_909,In_110);
nor U833 (N_833,In_379,N_145);
or U834 (N_834,In_444,In_1677);
and U835 (N_835,N_614,N_680);
and U836 (N_836,In_1336,In_132);
nand U837 (N_837,N_723,In_64);
nand U838 (N_838,In_1930,N_691);
and U839 (N_839,In_747,In_1523);
and U840 (N_840,N_628,In_529);
and U841 (N_841,In_585,In_1054);
nand U842 (N_842,N_741,In_666);
nor U843 (N_843,In_525,N_747);
nand U844 (N_844,In_348,N_80);
or U845 (N_845,N_795,N_355);
nand U846 (N_846,In_956,In_1982);
or U847 (N_847,N_732,In_1433);
and U848 (N_848,N_448,N_65);
nand U849 (N_849,N_632,In_1342);
xor U850 (N_850,N_280,N_584);
or U851 (N_851,N_123,In_135);
or U852 (N_852,In_634,In_1854);
xor U853 (N_853,N_114,N_224);
and U854 (N_854,In_1634,In_1570);
and U855 (N_855,In_1696,In_722);
nor U856 (N_856,In_441,N_421);
nand U857 (N_857,N_411,In_1164);
or U858 (N_858,N_396,N_636);
and U859 (N_859,In_3,In_480);
nand U860 (N_860,In_792,N_79);
nor U861 (N_861,In_17,In_1786);
nand U862 (N_862,N_761,In_1243);
nand U863 (N_863,N_277,N_409);
and U864 (N_864,N_243,In_729);
nand U865 (N_865,In_196,In_957);
or U866 (N_866,In_1997,In_377);
and U867 (N_867,N_535,In_1462);
nor U868 (N_868,N_289,In_1727);
nand U869 (N_869,N_619,In_689);
nand U870 (N_870,In_1189,N_587);
and U871 (N_871,In_98,In_1415);
or U872 (N_872,In_468,N_627);
and U873 (N_873,In_247,N_709);
nor U874 (N_874,N_698,In_1515);
nor U875 (N_875,N_618,N_267);
and U876 (N_876,N_381,In_380);
nand U877 (N_877,N_539,In_396);
nor U878 (N_878,N_545,In_972);
or U879 (N_879,In_244,In_302);
or U880 (N_880,N_658,N_76);
nor U881 (N_881,In_1414,In_286);
or U882 (N_882,N_564,In_1885);
and U883 (N_883,In_1453,N_443);
nor U884 (N_884,In_357,N_758);
and U885 (N_885,N_553,In_1579);
nand U886 (N_886,In_1196,In_562);
and U887 (N_887,N_776,N_357);
nor U888 (N_888,N_163,N_742);
nor U889 (N_889,N_746,N_766);
nand U890 (N_890,N_395,In_241);
and U891 (N_891,In_1605,In_1506);
or U892 (N_892,N_663,N_270);
and U893 (N_893,N_697,In_1222);
and U894 (N_894,N_711,N_774);
and U895 (N_895,In_1469,In_1948);
nand U896 (N_896,N_797,In_391);
and U897 (N_897,In_1648,In_732);
nor U898 (N_898,N_329,N_721);
nand U899 (N_899,In_1473,N_784);
nand U900 (N_900,In_1950,N_271);
or U901 (N_901,In_1178,In_900);
or U902 (N_902,N_400,In_1645);
or U903 (N_903,In_644,In_1309);
nor U904 (N_904,In_547,In_1156);
nor U905 (N_905,N_424,In_702);
and U906 (N_906,N_323,N_15);
or U907 (N_907,N_109,In_784);
nor U908 (N_908,In_1002,N_16);
nand U909 (N_909,N_672,In_305);
or U910 (N_910,N_276,N_660);
nand U911 (N_911,In_1496,In_264);
and U912 (N_912,N_771,N_26);
and U913 (N_913,N_9,In_463);
or U914 (N_914,In_713,N_391);
nor U915 (N_915,N_494,In_129);
and U916 (N_916,In_109,N_511);
nand U917 (N_917,In_600,In_280);
nor U918 (N_918,In_836,N_523);
nor U919 (N_919,N_791,In_113);
or U920 (N_920,N_338,In_1941);
nor U921 (N_921,N_394,In_584);
nand U922 (N_922,N_417,N_452);
and U923 (N_923,In_1889,In_1169);
and U924 (N_924,N_459,N_534);
or U925 (N_925,In_1141,N_413);
nand U926 (N_926,In_1394,N_757);
nand U927 (N_927,In_26,In_1417);
and U928 (N_928,N_288,In_927);
nor U929 (N_929,N_150,N_679);
and U930 (N_930,In_304,In_476);
and U931 (N_931,In_1992,In_140);
nor U932 (N_932,In_1821,N_524);
nand U933 (N_933,N_631,N_682);
nand U934 (N_934,In_489,In_703);
nor U935 (N_935,N_222,N_760);
or U936 (N_936,In_1280,In_1146);
or U937 (N_937,In_1237,In_1483);
and U938 (N_938,N_609,In_418);
nor U939 (N_939,In_201,N_208);
or U940 (N_940,N_346,N_403);
nand U941 (N_941,N_576,In_690);
or U942 (N_942,In_1940,In_1422);
nor U943 (N_943,In_1328,In_1666);
nand U944 (N_944,In_1017,In_1655);
and U945 (N_945,In_1647,N_336);
nand U946 (N_946,In_687,In_1850);
or U947 (N_947,In_921,N_528);
nor U948 (N_948,N_704,N_522);
and U949 (N_949,N_588,N_740);
and U950 (N_950,In_611,N_656);
and U951 (N_951,N_273,In_430);
or U952 (N_952,In_1852,In_1855);
nand U953 (N_953,In_568,N_673);
or U954 (N_954,In_1338,N_670);
nor U955 (N_955,In_675,In_772);
or U956 (N_956,In_1590,In_1020);
or U957 (N_957,In_1252,N_703);
or U958 (N_958,N_451,In_538);
or U959 (N_959,N_139,N_737);
nor U960 (N_960,N_274,N_69);
nand U961 (N_961,In_1509,In_625);
nor U962 (N_962,In_1032,In_1346);
and U963 (N_963,N_788,In_833);
nor U964 (N_964,N_674,In_1916);
nand U965 (N_965,In_128,N_718);
nand U966 (N_966,N_373,In_919);
and U967 (N_967,In_188,In_450);
and U968 (N_968,N_601,In_1105);
or U969 (N_969,N_570,N_778);
xor U970 (N_970,In_334,In_1219);
nor U971 (N_971,In_1016,In_790);
or U972 (N_972,N_27,N_792);
nor U973 (N_973,N_55,N_708);
nor U974 (N_974,N_644,In_855);
nand U975 (N_975,N_495,In_89);
or U976 (N_976,In_25,In_1165);
and U977 (N_977,In_1838,N_418);
and U978 (N_978,N_782,In_1046);
or U979 (N_979,In_948,In_814);
or U980 (N_980,In_1609,In_214);
nand U981 (N_981,In_1846,In_217);
nor U982 (N_982,In_1615,N_580);
nand U983 (N_983,In_136,In_1332);
and U984 (N_984,In_1986,In_1065);
and U985 (N_985,In_835,In_1801);
and U986 (N_986,In_1664,In_1119);
nor U987 (N_987,In_949,N_655);
and U988 (N_988,In_1429,N_368);
nand U989 (N_989,In_1325,In_925);
and U990 (N_990,In_466,In_1555);
or U991 (N_991,N_364,In_298);
xor U992 (N_992,In_838,N_527);
nor U993 (N_993,N_297,N_608);
nor U994 (N_994,In_189,In_39);
or U995 (N_995,In_1527,N_444);
and U996 (N_996,In_652,N_529);
xnor U997 (N_997,N_375,In_1747);
nand U998 (N_998,In_521,N_141);
nand U999 (N_999,N_337,N_374);
nand U1000 (N_1000,In_914,N_303);
and U1001 (N_1001,In_502,In_1640);
nand U1002 (N_1002,N_915,N_794);
nand U1003 (N_1003,N_577,N_814);
nand U1004 (N_1004,N_491,N_32);
xor U1005 (N_1005,In_419,N_811);
nor U1006 (N_1006,In_530,In_401);
nor U1007 (N_1007,In_549,N_47);
or U1008 (N_1008,N_416,In_343);
nand U1009 (N_1009,N_617,In_187);
nor U1010 (N_1010,N_536,In_761);
nor U1011 (N_1011,In_1975,In_1047);
or U1012 (N_1012,In_1599,N_813);
and U1013 (N_1013,N_90,N_638);
nor U1014 (N_1014,N_821,N_385);
and U1015 (N_1015,In_1368,N_903);
and U1016 (N_1016,In_79,N_837);
or U1017 (N_1017,N_278,In_1380);
nand U1018 (N_1018,In_1673,N_383);
or U1019 (N_1019,N_981,N_885);
and U1020 (N_1020,N_877,N_629);
and U1021 (N_1021,N_756,In_1761);
or U1022 (N_1022,In_751,In_220);
nand U1023 (N_1023,N_769,In_1909);
or U1024 (N_1024,N_389,In_338);
nand U1025 (N_1025,N_751,In_1306);
nor U1026 (N_1026,N_753,N_57);
nor U1027 (N_1027,N_845,In_1188);
xnor U1028 (N_1028,In_59,In_885);
or U1029 (N_1029,N_693,In_344);
or U1030 (N_1030,N_176,N_21);
and U1031 (N_1031,In_527,N_855);
nand U1032 (N_1032,N_825,In_477);
nand U1033 (N_1033,In_766,In_336);
nand U1034 (N_1034,In_226,In_315);
nand U1035 (N_1035,In_1709,N_994);
or U1036 (N_1036,In_1482,N_349);
nor U1037 (N_1037,N_937,N_863);
nor U1038 (N_1038,In_1878,N_533);
nand U1039 (N_1039,In_671,In_174);
nand U1040 (N_1040,In_432,N_369);
and U1041 (N_1041,N_625,In_374);
nor U1042 (N_1042,N_731,N_705);
or U1043 (N_1043,N_611,In_1211);
or U1044 (N_1044,In_1101,N_40);
or U1045 (N_1045,In_86,N_967);
nor U1046 (N_1046,N_314,In_1294);
nor U1047 (N_1047,N_935,N_210);
nand U1048 (N_1048,In_36,In_913);
and U1049 (N_1049,N_68,In_745);
or U1050 (N_1050,In_806,In_647);
or U1051 (N_1051,In_84,N_292);
or U1052 (N_1052,N_969,N_591);
and U1053 (N_1053,In_777,In_464);
or U1054 (N_1054,N_121,N_439);
nand U1055 (N_1055,N_934,In_385);
and U1056 (N_1056,In_1437,In_114);
or U1057 (N_1057,In_1685,In_1707);
and U1058 (N_1058,N_962,N_82);
or U1059 (N_1059,N_951,In_1627);
or U1060 (N_1060,In_1324,N_733);
or U1061 (N_1061,N_454,N_559);
and U1062 (N_1062,N_258,In_108);
nand U1063 (N_1063,N_809,N_198);
or U1064 (N_1064,N_815,In_211);
nor U1065 (N_1065,In_1151,In_347);
nor U1066 (N_1066,N_472,N_906);
and U1067 (N_1067,N_397,In_1316);
or U1068 (N_1068,N_835,N_2);
nand U1069 (N_1069,In_842,In_349);
nor U1070 (N_1070,N_685,In_117);
or U1071 (N_1071,In_1695,N_147);
or U1072 (N_1072,N_635,N_908);
and U1073 (N_1073,N_668,N_964);
and U1074 (N_1074,N_404,N_713);
and U1075 (N_1075,In_1411,N_650);
nand U1076 (N_1076,N_361,N_127);
or U1077 (N_1077,In_682,In_1893);
nor U1078 (N_1078,N_902,N_930);
and U1079 (N_1079,In_1650,N_957);
nand U1080 (N_1080,N_442,N_305);
or U1081 (N_1081,In_358,N_850);
nor U1082 (N_1082,In_351,In_38);
nand U1083 (N_1083,N_392,In_27);
and U1084 (N_1084,N_840,N_887);
and U1085 (N_1085,N_112,In_996);
and U1086 (N_1086,N_531,In_839);
nor U1087 (N_1087,N_956,In_1301);
nand U1088 (N_1088,N_770,N_370);
or U1089 (N_1089,In_1796,In_1183);
nand U1090 (N_1090,In_1204,N_574);
nand U1091 (N_1091,In_1284,In_1140);
or U1092 (N_1092,In_1043,N_143);
nand U1093 (N_1093,In_81,N_816);
nor U1094 (N_1094,N_223,N_268);
nand U1095 (N_1095,N_729,In_1097);
nor U1096 (N_1096,In_499,In_218);
nor U1097 (N_1097,N_453,N_805);
or U1098 (N_1098,N_242,N_671);
or U1099 (N_1099,In_851,N_940);
nand U1100 (N_1100,In_787,In_817);
and U1101 (N_1101,In_975,In_998);
or U1102 (N_1102,In_1990,N_960);
and U1103 (N_1103,N_918,N_572);
nor U1104 (N_1104,In_1376,In_825);
and U1105 (N_1105,In_1587,N_762);
nand U1106 (N_1106,In_974,N_474);
and U1107 (N_1107,In_319,N_200);
nor U1108 (N_1108,In_1286,In_1841);
nand U1109 (N_1109,In_862,In_58);
or U1110 (N_1110,N_707,N_738);
or U1111 (N_1111,N_768,N_231);
or U1112 (N_1112,In_736,In_874);
or U1113 (N_1113,N_301,In_707);
or U1114 (N_1114,In_1287,In_840);
or U1115 (N_1115,N_779,In_1899);
nor U1116 (N_1116,N_804,In_618);
and U1117 (N_1117,N_904,In_1520);
and U1118 (N_1118,N_763,N_692);
nor U1119 (N_1119,N_968,N_744);
and U1120 (N_1120,In_14,N_700);
nor U1121 (N_1121,N_806,In_830);
nor U1122 (N_1122,N_890,N_388);
and U1123 (N_1123,In_617,N_313);
or U1124 (N_1124,N_613,N_879);
nor U1125 (N_1125,N_911,In_462);
nor U1126 (N_1126,N_945,In_1994);
and U1127 (N_1127,In_985,N_284);
and U1128 (N_1128,N_916,N_914);
and U1129 (N_1129,In_645,In_1068);
nand U1130 (N_1130,N_253,In_1604);
xnor U1131 (N_1131,In_457,In_811);
and U1132 (N_1132,N_724,In_1548);
nor U1133 (N_1133,N_861,N_201);
or U1134 (N_1134,In_1746,N_818);
nand U1135 (N_1135,In_1822,In_245);
nand U1136 (N_1136,N_972,In_1257);
and U1137 (N_1137,N_560,N_810);
nand U1138 (N_1138,N_378,N_376);
nand U1139 (N_1139,N_606,In_1560);
and U1140 (N_1140,N_894,In_1187);
nor U1141 (N_1141,N_232,N_335);
and U1142 (N_1142,N_367,N_830);
nor U1143 (N_1143,N_247,In_56);
nor U1144 (N_1144,N_973,In_1563);
nor U1145 (N_1145,In_1894,N_59);
nand U1146 (N_1146,N_720,In_1329);
nor U1147 (N_1147,N_101,In_18);
nand U1148 (N_1148,N_843,N_836);
or U1149 (N_1149,In_54,In_142);
or U1150 (N_1150,In_1933,In_1759);
nor U1151 (N_1151,N_853,In_847);
nand U1152 (N_1152,N_997,N_488);
nand U1153 (N_1153,N_290,In_1001);
nand U1154 (N_1154,N_513,In_105);
nor U1155 (N_1155,N_715,N_944);
and U1156 (N_1156,N_922,N_995);
nand U1157 (N_1157,In_988,In_8);
nand U1158 (N_1158,In_1220,In_16);
nor U1159 (N_1159,In_1171,N_390);
nor U1160 (N_1160,In_265,N_353);
or U1161 (N_1161,N_645,N_800);
and U1162 (N_1162,In_1698,N_91);
nor U1163 (N_1163,N_347,N_434);
xor U1164 (N_1164,In_40,N_828);
or U1165 (N_1165,N_194,N_921);
nand U1166 (N_1166,In_1731,In_829);
or U1167 (N_1167,N_851,In_1657);
and U1168 (N_1168,N_988,N_947);
nand U1169 (N_1169,N_749,In_1900);
and U1170 (N_1170,In_1782,In_256);
and U1171 (N_1171,In_633,N_354);
or U1172 (N_1172,N_544,N_829);
nor U1173 (N_1173,In_1006,N_952);
or U1174 (N_1174,N_839,N_654);
or U1175 (N_1175,In_859,N_978);
nor U1176 (N_1176,N_233,N_786);
and U1177 (N_1177,In_1173,N_589);
or U1178 (N_1178,N_599,N_714);
and U1179 (N_1179,In_537,In_654);
and U1180 (N_1180,N_895,In_1557);
and U1181 (N_1181,In_782,N_604);
nand U1182 (N_1182,N_717,N_881);
nor U1183 (N_1183,In_1230,In_738);
nand U1184 (N_1184,N_873,N_684);
nand U1185 (N_1185,N_304,In_794);
nand U1186 (N_1186,In_1162,N_950);
or U1187 (N_1187,N_976,In_1293);
nor U1188 (N_1188,In_1625,In_145);
nand U1189 (N_1189,N_681,N_239);
nor U1190 (N_1190,N_869,In_339);
or U1191 (N_1191,N_189,N_185);
nand U1192 (N_1192,In_1719,N_739);
or U1193 (N_1193,In_1060,N_683);
and U1194 (N_1194,N_240,N_360);
nor U1195 (N_1195,N_217,N_983);
nand U1196 (N_1196,In_1676,In_964);
nor U1197 (N_1197,N_481,N_25);
or U1198 (N_1198,N_898,In_1572);
nor U1199 (N_1199,In_168,N_687);
nor U1200 (N_1200,N_1157,N_1008);
xnor U1201 (N_1201,In_70,In_1341);
xnor U1202 (N_1202,N_790,N_701);
or U1203 (N_1203,In_1069,In_1608);
or U1204 (N_1204,In_221,In_1134);
nor U1205 (N_1205,N_1021,N_1162);
or U1206 (N_1206,In_1351,N_555);
nand U1207 (N_1207,N_184,N_823);
nand U1208 (N_1208,In_1964,N_1158);
nand U1209 (N_1209,In_311,In_1352);
nor U1210 (N_1210,N_1142,In_119);
nand U1211 (N_1211,N_1189,N_827);
nand U1212 (N_1212,N_1078,N_1187);
nand U1213 (N_1213,In_1305,N_824);
and U1214 (N_1214,In_897,In_303);
or U1215 (N_1215,N_664,N_1023);
nor U1216 (N_1216,In_539,N_796);
or U1217 (N_1217,N_1135,N_907);
and U1218 (N_1218,In_1350,N_675);
or U1219 (N_1219,In_756,N_924);
or U1220 (N_1220,In_473,N_1014);
and U1221 (N_1221,N_214,N_195);
or U1222 (N_1222,N_563,N_857);
nand U1223 (N_1223,In_578,In_1389);
nor U1224 (N_1224,N_261,N_1098);
nand U1225 (N_1225,N_260,In_250);
nor U1226 (N_1226,In_1522,In_1813);
and U1227 (N_1227,In_1478,N_436);
or U1228 (N_1228,N_1017,N_514);
xnor U1229 (N_1229,In_1723,N_1059);
or U1230 (N_1230,N_530,In_616);
nand U1231 (N_1231,In_1884,N_1146);
nand U1232 (N_1232,N_1068,N_959);
and U1233 (N_1233,In_920,In_1360);
or U1234 (N_1234,N_525,In_1333);
or U1235 (N_1235,N_886,N_789);
and U1236 (N_1236,In_878,In_48);
or U1237 (N_1237,N_1055,In_1070);
or U1238 (N_1238,In_328,In_1107);
or U1239 (N_1239,N_1160,N_1010);
nor U1240 (N_1240,N_1025,N_498);
and U1241 (N_1241,N_605,In_1591);
or U1242 (N_1242,N_1026,In_1003);
and U1243 (N_1243,N_547,In_496);
nand U1244 (N_1244,N_897,N_998);
nand U1245 (N_1245,N_519,N_557);
nor U1246 (N_1246,N_1198,In_46);
nand U1247 (N_1247,N_931,N_876);
and U1248 (N_1248,In_1179,In_853);
nand U1249 (N_1249,N_1195,N_820);
nand U1250 (N_1250,N_339,In_1404);
and U1251 (N_1251,In_583,In_1239);
or U1252 (N_1252,In_171,In_443);
nand U1253 (N_1253,N_595,N_996);
nor U1254 (N_1254,In_1534,N_41);
nor U1255 (N_1255,N_316,N_958);
or U1256 (N_1256,N_1067,In_510);
nand U1257 (N_1257,In_433,N_1114);
or U1258 (N_1258,N_641,In_950);
nand U1259 (N_1259,N_775,N_912);
nor U1260 (N_1260,N_1169,N_991);
nor U1261 (N_1261,In_1238,N_269);
nand U1262 (N_1262,N_798,N_759);
or U1263 (N_1263,In_850,In_848);
or U1264 (N_1264,N_116,N_600);
and U1265 (N_1265,In_946,In_212);
nor U1266 (N_1266,N_549,N_646);
and U1267 (N_1267,In_74,In_1364);
nor U1268 (N_1268,In_1357,In_875);
nand U1269 (N_1269,N_992,N_1153);
and U1270 (N_1270,N_986,N_748);
or U1271 (N_1271,N_1137,N_1086);
or U1272 (N_1272,N_1046,In_277);
nand U1273 (N_1273,In_592,N_722);
or U1274 (N_1274,In_76,N_1105);
nor U1275 (N_1275,N_1173,In_979);
nor U1276 (N_1276,In_346,N_164);
nand U1277 (N_1277,In_865,In_581);
or U1278 (N_1278,N_1176,N_1020);
nand U1279 (N_1279,N_1053,N_1106);
and U1280 (N_1280,N_892,N_878);
nor U1281 (N_1281,N_826,In_1769);
or U1282 (N_1282,N_927,In_1282);
or U1283 (N_1283,N_651,N_1031);
nand U1284 (N_1284,N_665,N_974);
nor U1285 (N_1285,N_1143,In_252);
nand U1286 (N_1286,N_716,N_486);
nor U1287 (N_1287,N_807,N_750);
nor U1288 (N_1288,N_1000,In_535);
and U1289 (N_1289,N_1154,N_1118);
nand U1290 (N_1290,N_517,N_871);
or U1291 (N_1291,In_236,N_1085);
and U1292 (N_1292,In_799,N_963);
nor U1293 (N_1293,In_1208,In_639);
and U1294 (N_1294,N_846,N_933);
nand U1295 (N_1295,In_1270,N_1168);
nand U1296 (N_1296,N_883,N_610);
nand U1297 (N_1297,N_117,N_634);
nand U1298 (N_1298,N_510,N_1185);
and U1299 (N_1299,N_1072,In_968);
or U1300 (N_1300,In_1862,N_1050);
nand U1301 (N_1301,N_12,N_925);
or U1302 (N_1302,In_1641,N_859);
or U1303 (N_1303,N_954,In_930);
and U1304 (N_1304,In_353,N_484);
and U1305 (N_1305,In_1938,N_1033);
and U1306 (N_1306,N_18,In_1386);
nand U1307 (N_1307,N_838,N_428);
nand U1308 (N_1308,N_623,N_777);
nand U1309 (N_1309,N_1012,N_321);
and U1310 (N_1310,In_309,N_596);
and U1311 (N_1311,N_229,N_1179);
nand U1312 (N_1312,In_310,N_689);
nor U1313 (N_1313,N_438,In_1224);
or U1314 (N_1314,N_942,N_230);
or U1315 (N_1315,N_88,N_1049);
and U1316 (N_1316,N_1035,In_1972);
nor U1317 (N_1317,N_327,N_1058);
nor U1318 (N_1318,N_1140,N_1038);
nor U1319 (N_1319,In_1598,N_1104);
and U1320 (N_1320,N_345,N_647);
nand U1321 (N_1321,N_197,In_1094);
or U1322 (N_1322,N_582,N_667);
and U1323 (N_1323,N_889,In_1730);
and U1324 (N_1324,N_186,N_341);
or U1325 (N_1325,N_662,N_842);
or U1326 (N_1326,In_1711,N_987);
or U1327 (N_1327,In_1391,N_586);
nand U1328 (N_1328,N_970,In_516);
nor U1329 (N_1329,In_1051,In_293);
nand U1330 (N_1330,N_1199,N_462);
or U1331 (N_1331,In_285,In_301);
or U1332 (N_1332,N_407,N_696);
nand U1333 (N_1333,N_888,N_1184);
and U1334 (N_1334,N_1109,In_1345);
or U1335 (N_1335,In_371,N_946);
and U1336 (N_1336,In_685,N_616);
and U1337 (N_1337,N_1004,N_251);
nand U1338 (N_1338,N_583,N_546);
or U1339 (N_1339,N_734,In_1256);
nor U1340 (N_1340,In_1362,N_896);
or U1341 (N_1341,N_1099,In_1853);
and U1342 (N_1342,N_917,In_1064);
or U1343 (N_1343,N_541,N_780);
and U1344 (N_1344,N_1164,In_246);
or U1345 (N_1345,N_899,In_926);
nor U1346 (N_1346,N_1051,N_977);
nand U1347 (N_1347,N_929,N_858);
and U1348 (N_1348,N_872,In_458);
or U1349 (N_1349,In_78,N_1172);
nand U1350 (N_1350,N_875,In_1883);
and U1351 (N_1351,In_661,N_1065);
or U1352 (N_1352,N_657,N_900);
and U1353 (N_1353,N_980,N_252);
nand U1354 (N_1354,N_1054,N_803);
nand U1355 (N_1355,In_1291,In_906);
nand U1356 (N_1356,N_81,N_1037);
nor U1357 (N_1357,N_1069,N_53);
nand U1358 (N_1358,N_291,In_1438);
nor U1359 (N_1359,N_727,N_1003);
nand U1360 (N_1360,N_477,N_1115);
nand U1361 (N_1361,N_1092,N_1174);
and U1362 (N_1362,N_743,N_1071);
or U1363 (N_1363,N_433,In_1816);
nor U1364 (N_1364,In_1033,N_425);
nor U1365 (N_1365,N_961,N_867);
nand U1366 (N_1366,N_593,N_985);
nand U1367 (N_1367,In_1567,N_702);
nor U1368 (N_1368,N_695,In_1895);
and U1369 (N_1369,N_181,N_1063);
nand U1370 (N_1370,In_1742,In_1167);
and U1371 (N_1371,In_50,N_686);
nand U1372 (N_1372,N_630,In_478);
and U1373 (N_1373,N_216,In_1495);
or U1374 (N_1374,N_483,N_182);
or U1375 (N_1375,N_1163,N_1116);
nand U1376 (N_1376,In_269,N_1007);
or U1377 (N_1377,N_949,In_905);
and U1378 (N_1378,In_350,N_1133);
nand U1379 (N_1379,N_841,N_819);
and U1380 (N_1380,N_468,N_1113);
or U1381 (N_1381,In_320,In_414);
and U1382 (N_1382,N_621,N_1111);
or U1383 (N_1383,N_209,N_639);
or U1384 (N_1384,In_1713,In_1561);
nand U1385 (N_1385,In_1416,N_1080);
or U1386 (N_1386,N_783,N_659);
or U1387 (N_1387,N_1048,N_426);
and U1388 (N_1388,N_473,N_1156);
or U1389 (N_1389,N_1047,N_688);
nand U1390 (N_1390,In_190,N_1039);
xor U1391 (N_1391,In_1612,N_138);
nor U1392 (N_1392,N_1122,In_907);
nand U1393 (N_1393,N_979,N_1128);
xor U1394 (N_1394,N_832,N_975);
nand U1395 (N_1395,N_652,N_1027);
nor U1396 (N_1396,N_735,N_1193);
and U1397 (N_1397,N_1130,In_1508);
nand U1398 (N_1398,N_508,N_953);
nor U1399 (N_1399,In_1773,N_1108);
and U1400 (N_1400,N_781,In_1029);
nor U1401 (N_1401,N_910,N_1323);
nor U1402 (N_1402,In_852,In_1278);
nand U1403 (N_1403,N_755,N_1255);
and U1404 (N_1404,N_848,In_665);
and U1405 (N_1405,In_1340,N_1226);
nor U1406 (N_1406,N_162,In_1502);
and U1407 (N_1407,N_1028,N_1204);
nor U1408 (N_1408,N_1212,N_1147);
nor U1409 (N_1409,N_913,N_575);
nor U1410 (N_1410,N_1265,N_955);
or U1411 (N_1411,N_1299,N_1346);
nor U1412 (N_1412,N_1359,N_939);
and U1413 (N_1413,N_1167,In_945);
nor U1414 (N_1414,In_542,N_1388);
nand U1415 (N_1415,N_990,In_34);
or U1416 (N_1416,In_103,N_812);
nand U1417 (N_1417,N_578,N_1018);
and U1418 (N_1418,N_1317,N_1365);
or U1419 (N_1419,N_1150,N_1084);
nand U1420 (N_1420,N_1387,In_1772);
nand U1421 (N_1421,N_1015,N_874);
and U1422 (N_1422,N_571,N_1375);
nand U1423 (N_1423,N_1197,N_1235);
nand U1424 (N_1424,In_9,N_1029);
and U1425 (N_1425,N_1340,N_1088);
or U1426 (N_1426,In_1476,N_1367);
or U1427 (N_1427,N_880,In_789);
or U1428 (N_1428,N_603,N_206);
nand U1429 (N_1429,In_1231,N_1330);
nor U1430 (N_1430,N_63,N_567);
nand U1431 (N_1431,In_1487,N_1206);
and U1432 (N_1432,N_551,N_1370);
and U1433 (N_1433,N_1392,N_1041);
nor U1434 (N_1434,In_208,N_1350);
nor U1435 (N_1435,In_1267,N_1188);
and U1436 (N_1436,N_1070,N_865);
and U1437 (N_1437,N_1207,N_1279);
and U1438 (N_1438,N_1342,In_1844);
nor U1439 (N_1439,N_1309,N_1182);
nor U1440 (N_1440,N_83,N_380);
or U1441 (N_1441,N_1148,N_1374);
or U1442 (N_1442,N_1343,N_1295);
and U1443 (N_1443,N_1259,N_1227);
or U1444 (N_1444,N_745,N_241);
xnor U1445 (N_1445,N_965,In_727);
nand U1446 (N_1446,N_1262,In_543);
and U1447 (N_1447,N_802,In_340);
nor U1448 (N_1448,N_1332,N_1381);
nor U1449 (N_1449,N_699,N_1009);
nor U1450 (N_1450,N_458,In_943);
or U1451 (N_1451,N_33,N_706);
and U1452 (N_1452,N_1045,N_526);
or U1453 (N_1453,N_1382,In_595);
xor U1454 (N_1454,N_1327,N_1305);
nand U1455 (N_1455,In_134,N_1242);
nand U1456 (N_1456,In_1856,N_496);
or U1457 (N_1457,N_884,N_1244);
or U1458 (N_1458,N_573,N_1149);
or U1459 (N_1459,N_167,N_844);
and U1460 (N_1460,In_572,N_854);
nor U1461 (N_1461,N_901,N_371);
or U1462 (N_1462,N_1138,N_640);
or U1463 (N_1463,N_1361,In_1542);
nand U1464 (N_1464,N_1251,N_1228);
and U1465 (N_1465,N_1139,In_575);
and U1466 (N_1466,N_1257,In_1279);
nor U1467 (N_1467,In_1694,N_170);
and U1468 (N_1468,N_1186,N_1083);
nor U1469 (N_1469,In_1488,N_1205);
nor U1470 (N_1470,N_1032,N_1284);
and U1471 (N_1471,N_849,In_492);
or U1472 (N_1472,In_775,N_1229);
or U1473 (N_1473,N_1165,N_262);
nor U1474 (N_1474,N_1013,In_181);
nand U1475 (N_1475,N_1268,N_1094);
nor U1476 (N_1476,N_948,N_834);
or U1477 (N_1477,N_1089,N_187);
nor U1478 (N_1478,N_676,N_1379);
nand U1479 (N_1479,N_1101,In_1592);
nor U1480 (N_1480,N_238,N_1183);
or U1481 (N_1481,N_891,N_1219);
and U1482 (N_1482,N_982,In_822);
nand U1483 (N_1483,In_1763,N_1125);
and U1484 (N_1484,N_1132,N_1040);
nor U1485 (N_1485,N_213,N_1254);
nand U1486 (N_1486,N_1286,In_1820);
nor U1487 (N_1487,N_1353,N_42);
nor U1488 (N_1488,N_1221,N_257);
or U1489 (N_1489,N_1360,N_669);
or U1490 (N_1490,N_1329,N_643);
nand U1491 (N_1491,N_1249,N_133);
or U1492 (N_1492,N_1356,In_316);
nor U1493 (N_1493,N_633,In_239);
nor U1494 (N_1494,N_1398,N_920);
or U1495 (N_1495,N_1246,N_1238);
nand U1496 (N_1496,N_1311,N_1399);
nor U1497 (N_1497,N_754,In_810);
nand U1498 (N_1498,N_463,N_1395);
or U1499 (N_1499,N_1349,N_266);
nor U1500 (N_1500,N_1191,N_905);
and U1501 (N_1501,N_190,N_1151);
nand U1502 (N_1502,In_1378,In_407);
or U1503 (N_1503,N_1261,N_1260);
and U1504 (N_1504,N_1044,N_597);
nor U1505 (N_1505,N_1081,N_384);
or U1506 (N_1506,N_1036,In_1667);
or U1507 (N_1507,N_1326,N_772);
nand U1508 (N_1508,N_441,N_1074);
and U1509 (N_1509,N_1200,N_615);
nor U1510 (N_1510,N_1266,N_429);
nor U1511 (N_1511,N_552,N_1178);
nor U1512 (N_1512,N_1331,In_370);
nand U1513 (N_1513,In_1944,N_1090);
or U1514 (N_1514,N_1123,In_1623);
nor U1515 (N_1515,In_1318,N_1136);
nor U1516 (N_1516,N_1214,N_1344);
and U1517 (N_1517,N_1384,N_1364);
nand U1518 (N_1518,N_1371,N_70);
nor U1519 (N_1519,N_1333,In_793);
nor U1520 (N_1520,N_1222,N_1348);
nand U1521 (N_1521,In_32,N_1376);
nand U1522 (N_1522,N_909,N_106);
or U1523 (N_1523,N_1369,N_386);
nand U1524 (N_1524,N_1285,N_1296);
and U1525 (N_1525,N_941,In_327);
or U1526 (N_1526,N_926,N_1224);
or U1527 (N_1527,N_1120,N_1250);
and U1528 (N_1528,N_612,N_730);
nand U1529 (N_1529,In_594,N_1231);
or U1530 (N_1530,N_435,N_882);
and U1531 (N_1531,N_1302,N_1216);
xnor U1532 (N_1532,In_397,N_1103);
xnor U1533 (N_1533,N_864,N_1303);
nor U1534 (N_1534,In_182,N_1192);
nor U1535 (N_1535,N_1241,N_1247);
nand U1536 (N_1536,N_1306,In_608);
nand U1537 (N_1537,In_1399,N_237);
and U1538 (N_1538,In_1458,In_484);
or U1539 (N_1539,N_1263,In_1683);
nor U1540 (N_1540,In_1144,In_596);
nand U1541 (N_1541,N_1210,In_1556);
nand U1542 (N_1542,N_1145,N_1289);
nand U1543 (N_1543,N_6,In_213);
and U1544 (N_1544,N_1271,N_179);
nand U1545 (N_1545,N_1310,In_1111);
nand U1546 (N_1546,N_1062,N_1218);
nor U1547 (N_1547,N_1393,N_1079);
and U1548 (N_1548,N_1372,N_1270);
nand U1549 (N_1549,In_1617,N_51);
nand U1550 (N_1550,N_1391,N_1322);
or U1551 (N_1551,N_1308,N_1121);
or U1552 (N_1552,N_642,N_1082);
and U1553 (N_1553,N_501,In_672);
nand U1554 (N_1554,N_736,In_1147);
and U1555 (N_1555,N_1290,N_1358);
nand U1556 (N_1556,In_843,N_928);
and U1557 (N_1557,N_1386,N_1141);
nand U1558 (N_1558,N_1066,N_1223);
and U1559 (N_1559,N_1294,N_1338);
nand U1560 (N_1560,N_1256,N_984);
nor U1561 (N_1561,N_764,N_1177);
nand U1562 (N_1562,N_1276,In_1145);
and U1563 (N_1563,N_1129,N_1313);
nor U1564 (N_1564,N_1196,N_1274);
xnor U1565 (N_1565,In_1610,In_1327);
nor U1566 (N_1566,N_1076,N_1234);
nor U1567 (N_1567,N_1321,N_1315);
nand U1568 (N_1568,N_936,N_1144);
nor U1569 (N_1569,In_1135,N_1339);
and U1570 (N_1570,N_1264,In_1268);
and U1571 (N_1571,N_1380,N_661);
and U1572 (N_1572,N_509,N_847);
nand U1573 (N_1573,N_119,N_1159);
or U1574 (N_1574,N_1005,N_1016);
nor U1575 (N_1575,N_1283,N_1267);
nor U1576 (N_1576,In_471,N_1233);
nand U1577 (N_1577,N_626,N_1287);
and U1578 (N_1578,In_467,N_1181);
or U1579 (N_1579,N_1383,N_919);
and U1580 (N_1580,N_870,N_1239);
or U1581 (N_1581,N_893,N_1307);
nand U1582 (N_1582,N_1354,N_149);
or U1583 (N_1583,N_1275,N_1152);
and U1584 (N_1584,In_1867,N_1282);
or U1585 (N_1585,In_1783,In_1819);
or U1586 (N_1586,In_681,N_1312);
nor U1587 (N_1587,N_1240,N_1180);
and U1588 (N_1588,N_1237,N_678);
nand U1589 (N_1589,N_1253,N_550);
nor U1590 (N_1590,N_1258,In_1981);
nor U1591 (N_1591,N_694,N_1119);
or U1592 (N_1592,N_712,N_1112);
nor U1593 (N_1593,N_1345,In_763);
and U1594 (N_1594,N_1097,N_13);
nor U1595 (N_1595,N_1341,In_13);
or U1596 (N_1596,In_88,N_423);
or U1597 (N_1597,N_1245,N_1293);
or U1598 (N_1598,In_1538,N_822);
nand U1599 (N_1599,N_1209,N_765);
nor U1600 (N_1600,N_1520,In_87);
and U1601 (N_1601,N_1413,N_1194);
nor U1602 (N_1602,N_1458,N_1537);
and U1603 (N_1603,N_1019,N_1463);
nand U1604 (N_1604,N_852,N_1161);
nor U1605 (N_1605,N_1420,N_1175);
or U1606 (N_1606,In_711,N_1454);
nor U1607 (N_1607,N_1061,N_1538);
and U1608 (N_1608,N_1403,N_0);
nand U1609 (N_1609,N_767,In_237);
nand U1610 (N_1610,N_1496,In_306);
nor U1611 (N_1611,N_1217,N_1368);
and U1612 (N_1612,N_1489,N_1402);
and U1613 (N_1613,N_1437,N_1549);
nor U1614 (N_1614,N_1208,N_1573);
nor U1615 (N_1615,N_1414,N_653);
nand U1616 (N_1616,N_1378,N_1546);
nor U1617 (N_1617,N_1318,N_1495);
and U1618 (N_1618,N_1587,N_1459);
or U1619 (N_1619,N_799,N_1225);
nor U1620 (N_1620,N_348,N_1441);
nor U1621 (N_1621,N_1211,N_993);
and U1622 (N_1622,N_1569,N_475);
and U1623 (N_1623,N_1406,In_1269);
nor U1624 (N_1624,N_1423,N_1377);
nor U1625 (N_1625,N_801,N_1487);
and U1626 (N_1626,N_649,N_1100);
or U1627 (N_1627,N_1482,N_1336);
and U1628 (N_1628,In_360,N_1510);
nand U1629 (N_1629,N_1591,N_419);
nor U1630 (N_1630,N_1567,N_1316);
nand U1631 (N_1631,N_1529,In_125);
or U1632 (N_1632,N_1431,N_1478);
and U1633 (N_1633,N_1304,In_363);
nand U1634 (N_1634,N_1102,In_1304);
and U1635 (N_1635,N_1220,N_1508);
nor U1636 (N_1636,N_1001,In_1903);
nor U1637 (N_1637,N_1445,N_1554);
nand U1638 (N_1638,N_1483,N_1297);
or U1639 (N_1639,N_1213,N_1473);
nor U1640 (N_1640,N_1434,In_937);
or U1641 (N_1641,N_1556,N_1464);
nor U1642 (N_1642,N_1410,N_1586);
nor U1643 (N_1643,N_1486,N_1401);
or U1644 (N_1644,N_1439,N_471);
and U1645 (N_1645,N_382,In_730);
nor U1646 (N_1646,N_1301,N_1077);
nor U1647 (N_1647,N_728,N_1551);
nand U1648 (N_1648,N_1530,N_1492);
or U1649 (N_1649,N_516,In_1149);
nand U1650 (N_1650,N_966,N_1057);
or U1651 (N_1651,N_1540,N_1570);
nor U1652 (N_1652,In_733,N_1389);
and U1653 (N_1653,N_1230,N_1467);
or U1654 (N_1654,N_860,N_1056);
or U1655 (N_1655,N_1424,N_1568);
and U1656 (N_1656,N_1451,N_1170);
and U1657 (N_1657,N_1291,N_1599);
nand U1658 (N_1658,In_1322,N_923);
nand U1659 (N_1659,N_1485,N_1288);
nor U1660 (N_1660,N_817,N_1096);
nand U1661 (N_1661,N_1559,N_1416);
and U1662 (N_1662,N_1272,In_1954);
nor U1663 (N_1663,N_1390,In_1374);
or U1664 (N_1664,N_64,N_1584);
and U1665 (N_1665,N_1590,N_622);
or U1666 (N_1666,In_165,N_725);
nand U1667 (N_1667,N_1564,In_1467);
and U1668 (N_1668,N_1542,N_862);
and U1669 (N_1669,N_1002,N_1448);
or U1670 (N_1670,N_1512,N_1517);
nand U1671 (N_1671,N_1576,N_1432);
nor U1672 (N_1672,N_485,In_1260);
nand U1673 (N_1673,N_1427,N_1166);
and U1674 (N_1674,N_1442,N_1248);
and U1675 (N_1675,N_146,N_1455);
nor U1676 (N_1676,N_1475,N_1465);
or U1677 (N_1677,N_1471,N_1417);
nor U1678 (N_1678,In_965,N_1407);
or U1679 (N_1679,In_1381,N_1553);
nand U1680 (N_1680,In_1492,N_1503);
and U1681 (N_1681,N_1351,N_1460);
nor U1682 (N_1682,In_1976,N_1190);
or U1683 (N_1683,N_1506,N_1444);
xor U1684 (N_1684,N_1042,N_1446);
nor U1685 (N_1685,N_1052,N_1469);
or U1686 (N_1686,N_1024,N_406);
nor U1687 (N_1687,N_1127,N_1522);
or U1688 (N_1688,N_856,N_1594);
nor U1689 (N_1689,N_620,N_1515);
or U1690 (N_1690,N_1548,N_1531);
and U1691 (N_1691,N_1335,N_1494);
and U1692 (N_1692,N_1596,N_1415);
or U1693 (N_1693,N_1425,In_1420);
or U1694 (N_1694,N_1528,N_1588);
nor U1695 (N_1695,N_1527,N_1043);
and U1696 (N_1696,N_542,N_1366);
nand U1697 (N_1697,N_1215,N_1479);
nand U1698 (N_1698,N_1545,In_1725);
nor U1699 (N_1699,N_1334,N_1509);
nor U1700 (N_1700,N_1095,In_215);
or U1701 (N_1701,N_1452,N_1578);
nand U1702 (N_1702,N_1273,N_1555);
xnor U1703 (N_1703,N_1589,N_1450);
nand U1704 (N_1704,N_1087,N_1502);
or U1705 (N_1705,N_1126,N_868);
and U1706 (N_1706,N_1474,N_1011);
and U1707 (N_1707,N_1281,N_1034);
nand U1708 (N_1708,N_1203,N_1557);
nor U1709 (N_1709,N_1466,N_1438);
nor U1710 (N_1710,N_1565,N_156);
nor U1711 (N_1711,N_1535,N_1405);
nand U1712 (N_1712,N_1435,N_1488);
and U1713 (N_1713,N_1064,N_1500);
nand U1714 (N_1714,N_1408,N_1443);
and U1715 (N_1715,N_1575,N_1499);
or U1716 (N_1716,N_1582,In_776);
nor U1717 (N_1717,N_1533,N_1550);
and U1718 (N_1718,N_1481,N_1447);
or U1719 (N_1719,N_1397,N_1547);
nor U1720 (N_1720,N_1337,N_1552);
nand U1721 (N_1721,N_1525,N_1558);
nor U1722 (N_1722,N_1357,N_1155);
or U1723 (N_1723,N_431,N_1498);
nand U1724 (N_1724,N_1472,N_1511);
nand U1725 (N_1725,N_1532,N_1091);
nand U1726 (N_1726,In_1798,In_1018);
or U1727 (N_1727,N_1544,In_942);
and U1728 (N_1728,N_1277,N_1453);
and U1729 (N_1729,N_1404,N_332);
nor U1730 (N_1730,N_1314,N_1476);
nor U1731 (N_1731,N_1574,In_1706);
nand U1732 (N_1732,N_1430,N_1560);
and U1733 (N_1733,N_1394,In_1440);
and U1734 (N_1734,N_793,N_1428);
and U1735 (N_1735,N_602,N_1524);
and U1736 (N_1736,N_1363,N_1480);
or U1737 (N_1737,N_943,N_1592);
nor U1738 (N_1738,N_1563,N_1490);
or U1739 (N_1739,N_1513,N_1519);
and U1740 (N_1740,N_690,N_1117);
nand U1741 (N_1741,N_1298,N_1504);
and U1742 (N_1742,In_144,N_1236);
nand U1743 (N_1743,N_1598,N_1457);
nor U1744 (N_1744,N_1426,N_1419);
or U1745 (N_1745,N_1534,N_989);
and U1746 (N_1746,N_1536,N_1543);
nand U1747 (N_1747,N_1493,N_422);
nand U1748 (N_1748,N_666,N_999);
or U1749 (N_1749,N_1541,N_1400);
and U1750 (N_1750,N_1412,N_1006);
nor U1751 (N_1751,In_903,N_1597);
nor U1752 (N_1752,N_1232,N_1022);
or U1753 (N_1753,N_1583,N_971);
nor U1754 (N_1754,N_1468,N_1577);
and U1755 (N_1755,N_1385,N_1396);
nor U1756 (N_1756,N_1585,N_1324);
nand U1757 (N_1757,N_1516,N_1521);
nand U1758 (N_1758,In_296,N_1501);
nor U1759 (N_1759,N_833,N_1202);
and U1760 (N_1760,N_1462,N_1075);
nor U1761 (N_1761,N_1562,N_492);
or U1762 (N_1762,N_1252,N_1107);
nand U1763 (N_1763,N_1373,N_102);
or U1764 (N_1764,N_1523,N_1595);
xnor U1765 (N_1765,N_1073,N_1300);
or U1766 (N_1766,N_1477,In_24);
or U1767 (N_1767,N_1134,N_1319);
nor U1768 (N_1768,N_866,N_1355);
nand U1769 (N_1769,N_1456,N_1328);
nor U1770 (N_1770,N_1418,N_1409);
or U1771 (N_1771,N_1436,N_1422);
and U1772 (N_1772,N_1171,In_1971);
and U1773 (N_1773,N_1093,N_1561);
nand U1774 (N_1774,N_1461,N_235);
and U1775 (N_1775,N_1505,N_1580);
and U1776 (N_1776,N_1320,N_1347);
or U1777 (N_1777,In_1109,N_1449);
nand U1778 (N_1778,N_1497,N_1325);
and U1779 (N_1779,N_1362,N_1243);
or U1780 (N_1780,N_677,N_1411);
nand U1781 (N_1781,N_1539,N_1110);
nand U1782 (N_1782,N_1514,N_1201);
and U1783 (N_1783,N_1280,N_1269);
nor U1784 (N_1784,N_1484,N_1440);
nor U1785 (N_1785,N_62,In_1073);
and U1786 (N_1786,N_1352,N_1571);
xnor U1787 (N_1787,N_1491,In_944);
and U1788 (N_1788,N_1470,N_500);
nor U1789 (N_1789,N_1518,N_1581);
nand U1790 (N_1790,N_808,N_773);
nor U1791 (N_1791,N_1507,N_1433);
nand U1792 (N_1792,N_1421,N_1593);
or U1793 (N_1793,N_1572,N_1429);
nand U1794 (N_1794,N_1030,N_1060);
and U1795 (N_1795,N_831,N_932);
and U1796 (N_1796,N_1131,N_1278);
or U1797 (N_1797,N_1579,N_1566);
and U1798 (N_1798,N_1292,N_1124);
nor U1799 (N_1799,N_938,N_1526);
or U1800 (N_1800,N_1714,N_1650);
and U1801 (N_1801,N_1603,N_1711);
nor U1802 (N_1802,N_1640,N_1700);
nor U1803 (N_1803,N_1605,N_1668);
xor U1804 (N_1804,N_1658,N_1713);
or U1805 (N_1805,N_1725,N_1673);
nor U1806 (N_1806,N_1695,N_1619);
and U1807 (N_1807,N_1751,N_1698);
nor U1808 (N_1808,N_1697,N_1622);
nor U1809 (N_1809,N_1652,N_1749);
nor U1810 (N_1810,N_1703,N_1674);
nor U1811 (N_1811,N_1748,N_1781);
nand U1812 (N_1812,N_1790,N_1638);
nand U1813 (N_1813,N_1601,N_1761);
nand U1814 (N_1814,N_1712,N_1688);
and U1815 (N_1815,N_1689,N_1607);
nand U1816 (N_1816,N_1710,N_1686);
nand U1817 (N_1817,N_1647,N_1609);
nand U1818 (N_1818,N_1798,N_1777);
or U1819 (N_1819,N_1610,N_1677);
or U1820 (N_1820,N_1796,N_1758);
and U1821 (N_1821,N_1735,N_1684);
and U1822 (N_1822,N_1683,N_1726);
or U1823 (N_1823,N_1627,N_1661);
xnor U1824 (N_1824,N_1694,N_1727);
nor U1825 (N_1825,N_1653,N_1679);
nand U1826 (N_1826,N_1680,N_1624);
nand U1827 (N_1827,N_1718,N_1730);
nor U1828 (N_1828,N_1728,N_1693);
nand U1829 (N_1829,N_1626,N_1656);
nor U1830 (N_1830,N_1696,N_1769);
or U1831 (N_1831,N_1768,N_1691);
nand U1832 (N_1832,N_1669,N_1705);
or U1833 (N_1833,N_1775,N_1614);
and U1834 (N_1834,N_1739,N_1715);
and U1835 (N_1835,N_1742,N_1745);
nor U1836 (N_1836,N_1618,N_1651);
nand U1837 (N_1837,N_1762,N_1682);
nor U1838 (N_1838,N_1717,N_1702);
nor U1839 (N_1839,N_1662,N_1719);
or U1840 (N_1840,N_1635,N_1690);
and U1841 (N_1841,N_1724,N_1630);
and U1842 (N_1842,N_1634,N_1741);
nor U1843 (N_1843,N_1763,N_1699);
or U1844 (N_1844,N_1667,N_1789);
or U1845 (N_1845,N_1657,N_1760);
or U1846 (N_1846,N_1767,N_1786);
nor U1847 (N_1847,N_1687,N_1746);
or U1848 (N_1848,N_1615,N_1799);
nand U1849 (N_1849,N_1752,N_1738);
or U1850 (N_1850,N_1780,N_1685);
or U1851 (N_1851,N_1797,N_1787);
and U1852 (N_1852,N_1766,N_1611);
nor U1853 (N_1853,N_1747,N_1663);
or U1854 (N_1854,N_1707,N_1732);
or U1855 (N_1855,N_1733,N_1637);
nand U1856 (N_1856,N_1720,N_1666);
and U1857 (N_1857,N_1782,N_1729);
nand U1858 (N_1858,N_1606,N_1623);
nand U1859 (N_1859,N_1743,N_1704);
or U1860 (N_1860,N_1791,N_1788);
nor U1861 (N_1861,N_1636,N_1676);
or U1862 (N_1862,N_1716,N_1757);
nor U1863 (N_1863,N_1648,N_1646);
nand U1864 (N_1864,N_1617,N_1731);
and U1865 (N_1865,N_1645,N_1621);
nand U1866 (N_1866,N_1773,N_1753);
and U1867 (N_1867,N_1671,N_1783);
or U1868 (N_1868,N_1654,N_1600);
nor U1869 (N_1869,N_1723,N_1756);
nand U1870 (N_1870,N_1759,N_1664);
nand U1871 (N_1871,N_1672,N_1659);
nor U1872 (N_1872,N_1616,N_1706);
nor U1873 (N_1873,N_1744,N_1774);
and U1874 (N_1874,N_1631,N_1793);
or U1875 (N_1875,N_1701,N_1770);
nor U1876 (N_1876,N_1678,N_1629);
and U1877 (N_1877,N_1660,N_1675);
and U1878 (N_1878,N_1644,N_1625);
nand U1879 (N_1879,N_1620,N_1771);
xor U1880 (N_1880,N_1602,N_1632);
nor U1881 (N_1881,N_1772,N_1778);
or U1882 (N_1882,N_1649,N_1604);
nand U1883 (N_1883,N_1792,N_1692);
and U1884 (N_1884,N_1776,N_1708);
or U1885 (N_1885,N_1764,N_1765);
nor U1886 (N_1886,N_1795,N_1740);
or U1887 (N_1887,N_1670,N_1665);
or U1888 (N_1888,N_1613,N_1784);
or U1889 (N_1889,N_1709,N_1721);
nor U1890 (N_1890,N_1754,N_1642);
and U1891 (N_1891,N_1681,N_1779);
nand U1892 (N_1892,N_1785,N_1734);
nor U1893 (N_1893,N_1755,N_1722);
and U1894 (N_1894,N_1794,N_1641);
or U1895 (N_1895,N_1643,N_1750);
and U1896 (N_1896,N_1628,N_1655);
nor U1897 (N_1897,N_1608,N_1639);
nand U1898 (N_1898,N_1612,N_1737);
or U1899 (N_1899,N_1736,N_1633);
and U1900 (N_1900,N_1622,N_1612);
or U1901 (N_1901,N_1647,N_1765);
nand U1902 (N_1902,N_1797,N_1702);
and U1903 (N_1903,N_1706,N_1608);
and U1904 (N_1904,N_1707,N_1735);
or U1905 (N_1905,N_1613,N_1691);
xnor U1906 (N_1906,N_1788,N_1750);
and U1907 (N_1907,N_1728,N_1765);
or U1908 (N_1908,N_1652,N_1748);
nor U1909 (N_1909,N_1652,N_1710);
or U1910 (N_1910,N_1757,N_1666);
or U1911 (N_1911,N_1734,N_1602);
nor U1912 (N_1912,N_1645,N_1681);
nor U1913 (N_1913,N_1713,N_1721);
nor U1914 (N_1914,N_1696,N_1738);
nand U1915 (N_1915,N_1610,N_1761);
and U1916 (N_1916,N_1751,N_1622);
and U1917 (N_1917,N_1799,N_1684);
nand U1918 (N_1918,N_1629,N_1681);
or U1919 (N_1919,N_1762,N_1779);
nor U1920 (N_1920,N_1746,N_1632);
or U1921 (N_1921,N_1690,N_1758);
or U1922 (N_1922,N_1772,N_1612);
and U1923 (N_1923,N_1653,N_1754);
nor U1924 (N_1924,N_1730,N_1763);
or U1925 (N_1925,N_1638,N_1693);
or U1926 (N_1926,N_1732,N_1731);
and U1927 (N_1927,N_1713,N_1678);
and U1928 (N_1928,N_1756,N_1783);
or U1929 (N_1929,N_1763,N_1744);
nand U1930 (N_1930,N_1742,N_1702);
nand U1931 (N_1931,N_1628,N_1657);
and U1932 (N_1932,N_1778,N_1711);
nand U1933 (N_1933,N_1600,N_1682);
nor U1934 (N_1934,N_1666,N_1628);
or U1935 (N_1935,N_1611,N_1734);
nand U1936 (N_1936,N_1713,N_1700);
nor U1937 (N_1937,N_1728,N_1616);
or U1938 (N_1938,N_1702,N_1638);
nor U1939 (N_1939,N_1791,N_1746);
or U1940 (N_1940,N_1768,N_1736);
or U1941 (N_1941,N_1642,N_1720);
nand U1942 (N_1942,N_1653,N_1641);
nor U1943 (N_1943,N_1634,N_1621);
and U1944 (N_1944,N_1760,N_1622);
nor U1945 (N_1945,N_1739,N_1617);
nand U1946 (N_1946,N_1626,N_1642);
and U1947 (N_1947,N_1761,N_1696);
nand U1948 (N_1948,N_1791,N_1608);
or U1949 (N_1949,N_1611,N_1704);
or U1950 (N_1950,N_1649,N_1616);
nor U1951 (N_1951,N_1729,N_1742);
nor U1952 (N_1952,N_1646,N_1757);
and U1953 (N_1953,N_1623,N_1748);
nor U1954 (N_1954,N_1634,N_1639);
and U1955 (N_1955,N_1729,N_1733);
nand U1956 (N_1956,N_1651,N_1659);
or U1957 (N_1957,N_1798,N_1687);
nor U1958 (N_1958,N_1626,N_1691);
nand U1959 (N_1959,N_1667,N_1703);
nand U1960 (N_1960,N_1777,N_1678);
nor U1961 (N_1961,N_1793,N_1686);
or U1962 (N_1962,N_1600,N_1613);
nand U1963 (N_1963,N_1725,N_1687);
and U1964 (N_1964,N_1794,N_1617);
nor U1965 (N_1965,N_1741,N_1636);
or U1966 (N_1966,N_1657,N_1741);
nor U1967 (N_1967,N_1760,N_1632);
nand U1968 (N_1968,N_1787,N_1727);
and U1969 (N_1969,N_1785,N_1783);
nand U1970 (N_1970,N_1769,N_1788);
and U1971 (N_1971,N_1709,N_1666);
nand U1972 (N_1972,N_1690,N_1701);
nand U1973 (N_1973,N_1618,N_1649);
nand U1974 (N_1974,N_1763,N_1666);
xnor U1975 (N_1975,N_1730,N_1631);
nor U1976 (N_1976,N_1614,N_1761);
and U1977 (N_1977,N_1704,N_1719);
nand U1978 (N_1978,N_1799,N_1662);
xnor U1979 (N_1979,N_1613,N_1655);
nand U1980 (N_1980,N_1671,N_1644);
nor U1981 (N_1981,N_1664,N_1607);
nor U1982 (N_1982,N_1733,N_1728);
nor U1983 (N_1983,N_1618,N_1783);
or U1984 (N_1984,N_1751,N_1753);
nand U1985 (N_1985,N_1689,N_1776);
xor U1986 (N_1986,N_1624,N_1738);
nand U1987 (N_1987,N_1792,N_1738);
and U1988 (N_1988,N_1610,N_1725);
nand U1989 (N_1989,N_1698,N_1654);
or U1990 (N_1990,N_1610,N_1679);
and U1991 (N_1991,N_1713,N_1655);
and U1992 (N_1992,N_1656,N_1680);
or U1993 (N_1993,N_1719,N_1604);
nor U1994 (N_1994,N_1696,N_1603);
nand U1995 (N_1995,N_1771,N_1730);
or U1996 (N_1996,N_1658,N_1692);
nand U1997 (N_1997,N_1674,N_1621);
or U1998 (N_1998,N_1649,N_1753);
and U1999 (N_1999,N_1689,N_1681);
nor U2000 (N_2000,N_1939,N_1801);
and U2001 (N_2001,N_1905,N_1819);
and U2002 (N_2002,N_1874,N_1812);
nand U2003 (N_2003,N_1871,N_1860);
or U2004 (N_2004,N_1805,N_1880);
nor U2005 (N_2005,N_1859,N_1892);
nand U2006 (N_2006,N_1800,N_1932);
nand U2007 (N_2007,N_1869,N_1864);
nand U2008 (N_2008,N_1913,N_1988);
or U2009 (N_2009,N_1921,N_1978);
nand U2010 (N_2010,N_1893,N_1803);
or U2011 (N_2011,N_1862,N_1907);
or U2012 (N_2012,N_1854,N_1968);
and U2013 (N_2013,N_1828,N_1998);
nor U2014 (N_2014,N_1851,N_1951);
and U2015 (N_2015,N_1936,N_1933);
nand U2016 (N_2016,N_1982,N_1802);
nand U2017 (N_2017,N_1983,N_1993);
and U2018 (N_2018,N_1891,N_1996);
or U2019 (N_2019,N_1945,N_1957);
nand U2020 (N_2020,N_1840,N_1818);
or U2021 (N_2021,N_1898,N_1847);
nor U2022 (N_2022,N_1931,N_1959);
nand U2023 (N_2023,N_1810,N_1916);
nand U2024 (N_2024,N_1811,N_1920);
and U2025 (N_2025,N_1943,N_1886);
nand U2026 (N_2026,N_1873,N_1947);
nand U2027 (N_2027,N_1888,N_1855);
and U2028 (N_2028,N_1879,N_1868);
and U2029 (N_2029,N_1836,N_1877);
nand U2030 (N_2030,N_1815,N_1875);
or U2031 (N_2031,N_1928,N_1992);
and U2032 (N_2032,N_1838,N_1857);
and U2033 (N_2033,N_1915,N_1963);
or U2034 (N_2034,N_1911,N_1935);
or U2035 (N_2035,N_1927,N_1849);
or U2036 (N_2036,N_1882,N_1865);
nor U2037 (N_2037,N_1834,N_1899);
nand U2038 (N_2038,N_1926,N_1843);
or U2039 (N_2039,N_1853,N_1930);
xnor U2040 (N_2040,N_1906,N_1835);
or U2041 (N_2041,N_1842,N_1953);
or U2042 (N_2042,N_1950,N_1946);
nand U2043 (N_2043,N_1971,N_1841);
nand U2044 (N_2044,N_1856,N_1914);
or U2045 (N_2045,N_1977,N_1833);
nor U2046 (N_2046,N_1894,N_1948);
nand U2047 (N_2047,N_1878,N_1850);
or U2048 (N_2048,N_1955,N_1962);
and U2049 (N_2049,N_1852,N_1901);
or U2050 (N_2050,N_1980,N_1897);
or U2051 (N_2051,N_1986,N_1997);
and U2052 (N_2052,N_1960,N_1966);
nor U2053 (N_2053,N_1956,N_1823);
and U2054 (N_2054,N_1895,N_1990);
or U2055 (N_2055,N_1970,N_1813);
nand U2056 (N_2056,N_1985,N_1903);
or U2057 (N_2057,N_1807,N_1937);
or U2058 (N_2058,N_1964,N_1979);
nor U2059 (N_2059,N_1919,N_1984);
nand U2060 (N_2060,N_1909,N_1923);
nor U2061 (N_2061,N_1885,N_1973);
nand U2062 (N_2062,N_1830,N_1845);
nor U2063 (N_2063,N_1981,N_1822);
nor U2064 (N_2064,N_1816,N_1902);
nor U2065 (N_2065,N_1863,N_1858);
nand U2066 (N_2066,N_1804,N_1952);
nor U2067 (N_2067,N_1866,N_1876);
or U2068 (N_2068,N_1900,N_1994);
nand U2069 (N_2069,N_1825,N_1975);
or U2070 (N_2070,N_1890,N_1958);
nor U2071 (N_2071,N_1976,N_1965);
nand U2072 (N_2072,N_1809,N_1820);
nor U2073 (N_2073,N_1938,N_1829);
nand U2074 (N_2074,N_1814,N_1999);
or U2075 (N_2075,N_1969,N_1883);
nand U2076 (N_2076,N_1908,N_1941);
nand U2077 (N_2077,N_1910,N_1817);
and U2078 (N_2078,N_1806,N_1826);
or U2079 (N_2079,N_1904,N_1940);
or U2080 (N_2080,N_1944,N_1861);
nor U2081 (N_2081,N_1912,N_1848);
nor U2082 (N_2082,N_1991,N_1974);
nand U2083 (N_2083,N_1844,N_1821);
nand U2084 (N_2084,N_1924,N_1925);
nor U2085 (N_2085,N_1896,N_1867);
nor U2086 (N_2086,N_1887,N_1918);
nand U2087 (N_2087,N_1954,N_1881);
nor U2088 (N_2088,N_1934,N_1808);
or U2089 (N_2089,N_1870,N_1889);
nor U2090 (N_2090,N_1967,N_1832);
and U2091 (N_2091,N_1831,N_1987);
or U2092 (N_2092,N_1839,N_1989);
nor U2093 (N_2093,N_1922,N_1824);
nor U2094 (N_2094,N_1961,N_1884);
or U2095 (N_2095,N_1942,N_1827);
nand U2096 (N_2096,N_1949,N_1872);
nand U2097 (N_2097,N_1846,N_1995);
nor U2098 (N_2098,N_1929,N_1972);
nand U2099 (N_2099,N_1917,N_1837);
and U2100 (N_2100,N_1920,N_1939);
nand U2101 (N_2101,N_1885,N_1800);
or U2102 (N_2102,N_1811,N_1973);
nor U2103 (N_2103,N_1841,N_1956);
nand U2104 (N_2104,N_1959,N_1805);
nand U2105 (N_2105,N_1882,N_1928);
nand U2106 (N_2106,N_1982,N_1812);
or U2107 (N_2107,N_1969,N_1943);
or U2108 (N_2108,N_1950,N_1885);
nor U2109 (N_2109,N_1877,N_1986);
nand U2110 (N_2110,N_1864,N_1895);
nand U2111 (N_2111,N_1957,N_1844);
nor U2112 (N_2112,N_1928,N_1824);
nor U2113 (N_2113,N_1882,N_1843);
nand U2114 (N_2114,N_1903,N_1811);
nor U2115 (N_2115,N_1993,N_1823);
nand U2116 (N_2116,N_1847,N_1945);
and U2117 (N_2117,N_1926,N_1816);
nor U2118 (N_2118,N_1978,N_1882);
and U2119 (N_2119,N_1877,N_1805);
and U2120 (N_2120,N_1806,N_1976);
nand U2121 (N_2121,N_1927,N_1857);
and U2122 (N_2122,N_1855,N_1804);
and U2123 (N_2123,N_1801,N_1947);
nand U2124 (N_2124,N_1902,N_1918);
nor U2125 (N_2125,N_1988,N_1815);
or U2126 (N_2126,N_1908,N_1923);
and U2127 (N_2127,N_1933,N_1929);
nand U2128 (N_2128,N_1891,N_1890);
or U2129 (N_2129,N_1999,N_1939);
nand U2130 (N_2130,N_1964,N_1968);
nor U2131 (N_2131,N_1890,N_1889);
and U2132 (N_2132,N_1815,N_1963);
or U2133 (N_2133,N_1927,N_1827);
nand U2134 (N_2134,N_1925,N_1833);
nor U2135 (N_2135,N_1958,N_1853);
nand U2136 (N_2136,N_1941,N_1983);
or U2137 (N_2137,N_1891,N_1819);
and U2138 (N_2138,N_1871,N_1911);
or U2139 (N_2139,N_1981,N_1858);
nor U2140 (N_2140,N_1940,N_1842);
or U2141 (N_2141,N_1868,N_1877);
nand U2142 (N_2142,N_1971,N_1845);
or U2143 (N_2143,N_1829,N_1820);
nor U2144 (N_2144,N_1938,N_1978);
nand U2145 (N_2145,N_1989,N_1948);
nand U2146 (N_2146,N_1923,N_1925);
nand U2147 (N_2147,N_1820,N_1981);
and U2148 (N_2148,N_1848,N_1906);
nor U2149 (N_2149,N_1993,N_1999);
nand U2150 (N_2150,N_1835,N_1825);
nor U2151 (N_2151,N_1951,N_1836);
and U2152 (N_2152,N_1864,N_1988);
nand U2153 (N_2153,N_1855,N_1864);
nor U2154 (N_2154,N_1968,N_1884);
and U2155 (N_2155,N_1979,N_1841);
nor U2156 (N_2156,N_1801,N_1946);
nand U2157 (N_2157,N_1908,N_1931);
nor U2158 (N_2158,N_1964,N_1952);
nor U2159 (N_2159,N_1971,N_1816);
or U2160 (N_2160,N_1880,N_1822);
or U2161 (N_2161,N_1878,N_1871);
or U2162 (N_2162,N_1861,N_1864);
nand U2163 (N_2163,N_1928,N_1851);
and U2164 (N_2164,N_1839,N_1997);
nor U2165 (N_2165,N_1901,N_1990);
and U2166 (N_2166,N_1806,N_1906);
and U2167 (N_2167,N_1801,N_1948);
and U2168 (N_2168,N_1937,N_1893);
nor U2169 (N_2169,N_1851,N_1898);
nand U2170 (N_2170,N_1943,N_1910);
nand U2171 (N_2171,N_1981,N_1880);
nor U2172 (N_2172,N_1804,N_1842);
nand U2173 (N_2173,N_1894,N_1886);
and U2174 (N_2174,N_1862,N_1883);
nor U2175 (N_2175,N_1969,N_1835);
and U2176 (N_2176,N_1844,N_1890);
nor U2177 (N_2177,N_1928,N_1804);
nor U2178 (N_2178,N_1924,N_1942);
nand U2179 (N_2179,N_1898,N_1880);
nor U2180 (N_2180,N_1924,N_1963);
and U2181 (N_2181,N_1901,N_1937);
nor U2182 (N_2182,N_1889,N_1921);
nor U2183 (N_2183,N_1800,N_1832);
or U2184 (N_2184,N_1906,N_1938);
or U2185 (N_2185,N_1848,N_1860);
and U2186 (N_2186,N_1889,N_1976);
or U2187 (N_2187,N_1880,N_1997);
and U2188 (N_2188,N_1872,N_1892);
nand U2189 (N_2189,N_1989,N_1913);
and U2190 (N_2190,N_1870,N_1974);
or U2191 (N_2191,N_1980,N_1927);
or U2192 (N_2192,N_1907,N_1843);
nor U2193 (N_2193,N_1973,N_1880);
nand U2194 (N_2194,N_1857,N_1864);
nor U2195 (N_2195,N_1986,N_1898);
nand U2196 (N_2196,N_1834,N_1877);
or U2197 (N_2197,N_1854,N_1839);
nand U2198 (N_2198,N_1988,N_1868);
and U2199 (N_2199,N_1844,N_1927);
nor U2200 (N_2200,N_2177,N_2143);
nor U2201 (N_2201,N_2170,N_2138);
nor U2202 (N_2202,N_2041,N_2183);
nor U2203 (N_2203,N_2169,N_2115);
nor U2204 (N_2204,N_2055,N_2108);
nand U2205 (N_2205,N_2069,N_2196);
and U2206 (N_2206,N_2072,N_2151);
and U2207 (N_2207,N_2189,N_2077);
nand U2208 (N_2208,N_2101,N_2057);
nand U2209 (N_2209,N_2134,N_2104);
and U2210 (N_2210,N_2049,N_2197);
nor U2211 (N_2211,N_2199,N_2109);
and U2212 (N_2212,N_2064,N_2027);
or U2213 (N_2213,N_2154,N_2085);
nor U2214 (N_2214,N_2149,N_2082);
and U2215 (N_2215,N_2067,N_2174);
or U2216 (N_2216,N_2022,N_2025);
or U2217 (N_2217,N_2031,N_2146);
or U2218 (N_2218,N_2137,N_2176);
or U2219 (N_2219,N_2139,N_2142);
nand U2220 (N_2220,N_2158,N_2020);
nor U2221 (N_2221,N_2033,N_2047);
or U2222 (N_2222,N_2186,N_2079);
nor U2223 (N_2223,N_2181,N_2075);
nand U2224 (N_2224,N_2087,N_2097);
nand U2225 (N_2225,N_2026,N_2175);
nand U2226 (N_2226,N_2013,N_2122);
nor U2227 (N_2227,N_2102,N_2001);
or U2228 (N_2228,N_2081,N_2110);
and U2229 (N_2229,N_2065,N_2187);
and U2230 (N_2230,N_2179,N_2121);
nor U2231 (N_2231,N_2019,N_2116);
or U2232 (N_2232,N_2126,N_2074);
nand U2233 (N_2233,N_2078,N_2192);
and U2234 (N_2234,N_2073,N_2166);
nand U2235 (N_2235,N_2002,N_2129);
or U2236 (N_2236,N_2059,N_2058);
nand U2237 (N_2237,N_2091,N_2061);
nor U2238 (N_2238,N_2015,N_2133);
nor U2239 (N_2239,N_2178,N_2105);
nor U2240 (N_2240,N_2119,N_2161);
and U2241 (N_2241,N_2157,N_2172);
nor U2242 (N_2242,N_2114,N_2023);
or U2243 (N_2243,N_2046,N_2052);
or U2244 (N_2244,N_2009,N_2090);
nor U2245 (N_2245,N_2053,N_2063);
and U2246 (N_2246,N_2185,N_2144);
and U2247 (N_2247,N_2044,N_2092);
nor U2248 (N_2248,N_2029,N_2120);
or U2249 (N_2249,N_2050,N_2048);
or U2250 (N_2250,N_2088,N_2123);
or U2251 (N_2251,N_2008,N_2124);
nor U2252 (N_2252,N_2167,N_2099);
nand U2253 (N_2253,N_2117,N_2014);
and U2254 (N_2254,N_2024,N_2100);
and U2255 (N_2255,N_2113,N_2000);
nor U2256 (N_2256,N_2035,N_2125);
nand U2257 (N_2257,N_2068,N_2007);
nand U2258 (N_2258,N_2165,N_2136);
and U2259 (N_2259,N_2162,N_2037);
and U2260 (N_2260,N_2004,N_2159);
or U2261 (N_2261,N_2017,N_2148);
nor U2262 (N_2262,N_2152,N_2171);
nand U2263 (N_2263,N_2089,N_2191);
nor U2264 (N_2264,N_2111,N_2150);
nand U2265 (N_2265,N_2054,N_2128);
and U2266 (N_2266,N_2080,N_2094);
and U2267 (N_2267,N_2042,N_2010);
nand U2268 (N_2268,N_2011,N_2006);
nand U2269 (N_2269,N_2147,N_2182);
or U2270 (N_2270,N_2012,N_2032);
nand U2271 (N_2271,N_2135,N_2039);
and U2272 (N_2272,N_2036,N_2130);
nor U2273 (N_2273,N_2005,N_2038);
nand U2274 (N_2274,N_2131,N_2016);
xnor U2275 (N_2275,N_2107,N_2030);
and U2276 (N_2276,N_2003,N_2021);
or U2277 (N_2277,N_2066,N_2034);
or U2278 (N_2278,N_2188,N_2062);
or U2279 (N_2279,N_2194,N_2095);
or U2280 (N_2280,N_2190,N_2193);
and U2281 (N_2281,N_2070,N_2173);
and U2282 (N_2282,N_2140,N_2112);
nand U2283 (N_2283,N_2106,N_2083);
or U2284 (N_2284,N_2093,N_2103);
nand U2285 (N_2285,N_2060,N_2156);
or U2286 (N_2286,N_2184,N_2155);
or U2287 (N_2287,N_2096,N_2043);
nand U2288 (N_2288,N_2076,N_2071);
nor U2289 (N_2289,N_2098,N_2180);
nor U2290 (N_2290,N_2127,N_2045);
or U2291 (N_2291,N_2084,N_2056);
or U2292 (N_2292,N_2028,N_2168);
xnor U2293 (N_2293,N_2195,N_2164);
and U2294 (N_2294,N_2160,N_2118);
and U2295 (N_2295,N_2086,N_2153);
nand U2296 (N_2296,N_2051,N_2141);
and U2297 (N_2297,N_2145,N_2163);
or U2298 (N_2298,N_2040,N_2132);
nor U2299 (N_2299,N_2198,N_2018);
or U2300 (N_2300,N_2082,N_2094);
or U2301 (N_2301,N_2078,N_2154);
nand U2302 (N_2302,N_2082,N_2073);
and U2303 (N_2303,N_2188,N_2160);
nand U2304 (N_2304,N_2006,N_2023);
and U2305 (N_2305,N_2037,N_2169);
and U2306 (N_2306,N_2144,N_2134);
nand U2307 (N_2307,N_2166,N_2033);
or U2308 (N_2308,N_2045,N_2198);
and U2309 (N_2309,N_2000,N_2037);
nor U2310 (N_2310,N_2076,N_2113);
and U2311 (N_2311,N_2018,N_2037);
nand U2312 (N_2312,N_2025,N_2056);
and U2313 (N_2313,N_2002,N_2039);
nor U2314 (N_2314,N_2146,N_2056);
and U2315 (N_2315,N_2049,N_2198);
or U2316 (N_2316,N_2185,N_2062);
nand U2317 (N_2317,N_2162,N_2187);
nor U2318 (N_2318,N_2039,N_2164);
or U2319 (N_2319,N_2136,N_2152);
nor U2320 (N_2320,N_2012,N_2194);
nor U2321 (N_2321,N_2104,N_2154);
nand U2322 (N_2322,N_2015,N_2120);
nand U2323 (N_2323,N_2181,N_2046);
nor U2324 (N_2324,N_2151,N_2003);
or U2325 (N_2325,N_2055,N_2162);
or U2326 (N_2326,N_2022,N_2009);
and U2327 (N_2327,N_2139,N_2045);
nor U2328 (N_2328,N_2161,N_2170);
or U2329 (N_2329,N_2109,N_2063);
nor U2330 (N_2330,N_2146,N_2127);
or U2331 (N_2331,N_2199,N_2106);
and U2332 (N_2332,N_2037,N_2051);
and U2333 (N_2333,N_2179,N_2029);
and U2334 (N_2334,N_2018,N_2169);
or U2335 (N_2335,N_2155,N_2151);
nand U2336 (N_2336,N_2180,N_2007);
and U2337 (N_2337,N_2038,N_2169);
or U2338 (N_2338,N_2021,N_2037);
nand U2339 (N_2339,N_2150,N_2186);
nor U2340 (N_2340,N_2022,N_2108);
nand U2341 (N_2341,N_2122,N_2148);
nand U2342 (N_2342,N_2003,N_2121);
nor U2343 (N_2343,N_2172,N_2151);
nor U2344 (N_2344,N_2185,N_2045);
and U2345 (N_2345,N_2024,N_2129);
or U2346 (N_2346,N_2108,N_2063);
and U2347 (N_2347,N_2064,N_2092);
nand U2348 (N_2348,N_2021,N_2027);
or U2349 (N_2349,N_2186,N_2078);
nand U2350 (N_2350,N_2160,N_2184);
or U2351 (N_2351,N_2015,N_2156);
or U2352 (N_2352,N_2071,N_2139);
nor U2353 (N_2353,N_2114,N_2188);
and U2354 (N_2354,N_2001,N_2077);
nand U2355 (N_2355,N_2062,N_2002);
nor U2356 (N_2356,N_2067,N_2045);
nor U2357 (N_2357,N_2164,N_2128);
nor U2358 (N_2358,N_2065,N_2093);
nand U2359 (N_2359,N_2198,N_2027);
and U2360 (N_2360,N_2066,N_2069);
or U2361 (N_2361,N_2078,N_2027);
or U2362 (N_2362,N_2091,N_2129);
nor U2363 (N_2363,N_2101,N_2187);
nand U2364 (N_2364,N_2125,N_2049);
or U2365 (N_2365,N_2054,N_2141);
or U2366 (N_2366,N_2093,N_2194);
nand U2367 (N_2367,N_2012,N_2168);
nand U2368 (N_2368,N_2060,N_2095);
nor U2369 (N_2369,N_2078,N_2056);
nand U2370 (N_2370,N_2070,N_2035);
nand U2371 (N_2371,N_2180,N_2063);
nor U2372 (N_2372,N_2070,N_2020);
nand U2373 (N_2373,N_2189,N_2157);
or U2374 (N_2374,N_2148,N_2177);
xnor U2375 (N_2375,N_2186,N_2053);
nor U2376 (N_2376,N_2153,N_2022);
and U2377 (N_2377,N_2102,N_2176);
and U2378 (N_2378,N_2026,N_2087);
nor U2379 (N_2379,N_2167,N_2132);
nand U2380 (N_2380,N_2089,N_2195);
nand U2381 (N_2381,N_2004,N_2081);
or U2382 (N_2382,N_2140,N_2159);
and U2383 (N_2383,N_2062,N_2182);
and U2384 (N_2384,N_2134,N_2090);
nand U2385 (N_2385,N_2012,N_2052);
or U2386 (N_2386,N_2021,N_2080);
nand U2387 (N_2387,N_2124,N_2142);
and U2388 (N_2388,N_2052,N_2023);
or U2389 (N_2389,N_2193,N_2120);
or U2390 (N_2390,N_2196,N_2068);
xnor U2391 (N_2391,N_2107,N_2092);
and U2392 (N_2392,N_2176,N_2127);
and U2393 (N_2393,N_2172,N_2060);
and U2394 (N_2394,N_2033,N_2089);
nor U2395 (N_2395,N_2115,N_2130);
nand U2396 (N_2396,N_2077,N_2103);
and U2397 (N_2397,N_2010,N_2166);
nor U2398 (N_2398,N_2001,N_2166);
and U2399 (N_2399,N_2049,N_2012);
nor U2400 (N_2400,N_2296,N_2293);
nand U2401 (N_2401,N_2329,N_2206);
or U2402 (N_2402,N_2342,N_2333);
nand U2403 (N_2403,N_2301,N_2389);
nor U2404 (N_2404,N_2377,N_2357);
nor U2405 (N_2405,N_2273,N_2394);
and U2406 (N_2406,N_2303,N_2224);
or U2407 (N_2407,N_2276,N_2290);
or U2408 (N_2408,N_2381,N_2317);
or U2409 (N_2409,N_2239,N_2243);
or U2410 (N_2410,N_2348,N_2203);
nor U2411 (N_2411,N_2305,N_2252);
nand U2412 (N_2412,N_2214,N_2275);
and U2413 (N_2413,N_2259,N_2398);
and U2414 (N_2414,N_2332,N_2284);
or U2415 (N_2415,N_2265,N_2231);
nand U2416 (N_2416,N_2356,N_2360);
nor U2417 (N_2417,N_2248,N_2218);
or U2418 (N_2418,N_2285,N_2247);
and U2419 (N_2419,N_2277,N_2253);
nand U2420 (N_2420,N_2320,N_2223);
nor U2421 (N_2421,N_2232,N_2226);
nand U2422 (N_2422,N_2324,N_2220);
nor U2423 (N_2423,N_2246,N_2309);
or U2424 (N_2424,N_2399,N_2294);
or U2425 (N_2425,N_2291,N_2280);
or U2426 (N_2426,N_2233,N_2311);
or U2427 (N_2427,N_2271,N_2352);
or U2428 (N_2428,N_2374,N_2228);
nor U2429 (N_2429,N_2205,N_2328);
nand U2430 (N_2430,N_2359,N_2221);
nand U2431 (N_2431,N_2281,N_2336);
nor U2432 (N_2432,N_2347,N_2380);
or U2433 (N_2433,N_2297,N_2346);
nor U2434 (N_2434,N_2326,N_2373);
and U2435 (N_2435,N_2319,N_2264);
and U2436 (N_2436,N_2242,N_2244);
and U2437 (N_2437,N_2210,N_2371);
nand U2438 (N_2438,N_2379,N_2364);
nor U2439 (N_2439,N_2331,N_2261);
nand U2440 (N_2440,N_2208,N_2200);
or U2441 (N_2441,N_2327,N_2338);
or U2442 (N_2442,N_2213,N_2256);
nor U2443 (N_2443,N_2304,N_2386);
nand U2444 (N_2444,N_2260,N_2362);
nand U2445 (N_2445,N_2295,N_2351);
nor U2446 (N_2446,N_2343,N_2245);
nand U2447 (N_2447,N_2300,N_2368);
and U2448 (N_2448,N_2278,N_2251);
and U2449 (N_2449,N_2370,N_2255);
nand U2450 (N_2450,N_2202,N_2369);
nand U2451 (N_2451,N_2289,N_2257);
and U2452 (N_2452,N_2286,N_2314);
or U2453 (N_2453,N_2227,N_2395);
and U2454 (N_2454,N_2313,N_2238);
or U2455 (N_2455,N_2263,N_2321);
nor U2456 (N_2456,N_2358,N_2375);
and U2457 (N_2457,N_2225,N_2204);
and U2458 (N_2458,N_2287,N_2310);
nor U2459 (N_2459,N_2383,N_2353);
nor U2460 (N_2460,N_2298,N_2272);
and U2461 (N_2461,N_2241,N_2268);
nor U2462 (N_2462,N_2349,N_2397);
nand U2463 (N_2463,N_2288,N_2384);
or U2464 (N_2464,N_2299,N_2361);
nor U2465 (N_2465,N_2222,N_2234);
nand U2466 (N_2466,N_2316,N_2267);
and U2467 (N_2467,N_2388,N_2396);
and U2468 (N_2468,N_2254,N_2211);
or U2469 (N_2469,N_2236,N_2308);
nand U2470 (N_2470,N_2282,N_2217);
nand U2471 (N_2471,N_2270,N_2212);
nand U2472 (N_2472,N_2330,N_2325);
nand U2473 (N_2473,N_2207,N_2382);
nand U2474 (N_2474,N_2279,N_2323);
and U2475 (N_2475,N_2337,N_2315);
nor U2476 (N_2476,N_2240,N_2366);
or U2477 (N_2477,N_2391,N_2339);
and U2478 (N_2478,N_2219,N_2306);
nor U2479 (N_2479,N_2354,N_2262);
and U2480 (N_2480,N_2344,N_2269);
xnor U2481 (N_2481,N_2390,N_2292);
nand U2482 (N_2482,N_2302,N_2367);
or U2483 (N_2483,N_2274,N_2392);
nor U2484 (N_2484,N_2363,N_2335);
or U2485 (N_2485,N_2350,N_2230);
nor U2486 (N_2486,N_2340,N_2322);
or U2487 (N_2487,N_2387,N_2365);
and U2488 (N_2488,N_2318,N_2235);
and U2489 (N_2489,N_2250,N_2258);
nor U2490 (N_2490,N_2249,N_2372);
nand U2491 (N_2491,N_2216,N_2345);
nand U2492 (N_2492,N_2237,N_2266);
nand U2493 (N_2493,N_2378,N_2355);
and U2494 (N_2494,N_2209,N_2334);
nand U2495 (N_2495,N_2393,N_2283);
and U2496 (N_2496,N_2341,N_2312);
nor U2497 (N_2497,N_2201,N_2215);
or U2498 (N_2498,N_2376,N_2385);
or U2499 (N_2499,N_2307,N_2229);
nor U2500 (N_2500,N_2377,N_2394);
nor U2501 (N_2501,N_2375,N_2208);
or U2502 (N_2502,N_2303,N_2293);
or U2503 (N_2503,N_2397,N_2222);
nor U2504 (N_2504,N_2223,N_2319);
xnor U2505 (N_2505,N_2316,N_2387);
and U2506 (N_2506,N_2216,N_2316);
or U2507 (N_2507,N_2353,N_2200);
nor U2508 (N_2508,N_2282,N_2319);
and U2509 (N_2509,N_2386,N_2396);
nor U2510 (N_2510,N_2219,N_2361);
or U2511 (N_2511,N_2214,N_2364);
or U2512 (N_2512,N_2219,N_2340);
nor U2513 (N_2513,N_2281,N_2204);
nor U2514 (N_2514,N_2273,N_2312);
and U2515 (N_2515,N_2288,N_2390);
nor U2516 (N_2516,N_2346,N_2399);
and U2517 (N_2517,N_2221,N_2229);
and U2518 (N_2518,N_2333,N_2361);
or U2519 (N_2519,N_2336,N_2345);
and U2520 (N_2520,N_2280,N_2260);
and U2521 (N_2521,N_2274,N_2327);
nand U2522 (N_2522,N_2283,N_2208);
or U2523 (N_2523,N_2263,N_2377);
nor U2524 (N_2524,N_2266,N_2218);
nand U2525 (N_2525,N_2232,N_2267);
nand U2526 (N_2526,N_2278,N_2207);
or U2527 (N_2527,N_2399,N_2327);
or U2528 (N_2528,N_2280,N_2325);
nor U2529 (N_2529,N_2211,N_2360);
or U2530 (N_2530,N_2280,N_2220);
or U2531 (N_2531,N_2297,N_2344);
or U2532 (N_2532,N_2336,N_2235);
or U2533 (N_2533,N_2394,N_2266);
nor U2534 (N_2534,N_2327,N_2364);
nor U2535 (N_2535,N_2249,N_2318);
nand U2536 (N_2536,N_2294,N_2347);
and U2537 (N_2537,N_2234,N_2236);
and U2538 (N_2538,N_2230,N_2367);
or U2539 (N_2539,N_2339,N_2214);
or U2540 (N_2540,N_2240,N_2264);
nor U2541 (N_2541,N_2343,N_2224);
and U2542 (N_2542,N_2256,N_2375);
and U2543 (N_2543,N_2344,N_2256);
nor U2544 (N_2544,N_2344,N_2324);
nor U2545 (N_2545,N_2210,N_2279);
or U2546 (N_2546,N_2289,N_2297);
nand U2547 (N_2547,N_2299,N_2309);
or U2548 (N_2548,N_2383,N_2314);
or U2549 (N_2549,N_2205,N_2363);
or U2550 (N_2550,N_2216,N_2224);
nand U2551 (N_2551,N_2284,N_2393);
or U2552 (N_2552,N_2350,N_2357);
nor U2553 (N_2553,N_2258,N_2353);
nor U2554 (N_2554,N_2325,N_2316);
or U2555 (N_2555,N_2312,N_2316);
or U2556 (N_2556,N_2383,N_2266);
nand U2557 (N_2557,N_2399,N_2209);
or U2558 (N_2558,N_2247,N_2294);
nor U2559 (N_2559,N_2322,N_2279);
nor U2560 (N_2560,N_2388,N_2258);
nor U2561 (N_2561,N_2223,N_2274);
nor U2562 (N_2562,N_2276,N_2372);
and U2563 (N_2563,N_2211,N_2275);
nor U2564 (N_2564,N_2340,N_2244);
nor U2565 (N_2565,N_2239,N_2209);
or U2566 (N_2566,N_2240,N_2364);
nor U2567 (N_2567,N_2244,N_2260);
or U2568 (N_2568,N_2343,N_2232);
and U2569 (N_2569,N_2316,N_2224);
nand U2570 (N_2570,N_2335,N_2399);
and U2571 (N_2571,N_2208,N_2322);
or U2572 (N_2572,N_2266,N_2294);
or U2573 (N_2573,N_2272,N_2366);
nand U2574 (N_2574,N_2231,N_2257);
nor U2575 (N_2575,N_2250,N_2338);
nand U2576 (N_2576,N_2219,N_2260);
nor U2577 (N_2577,N_2304,N_2292);
and U2578 (N_2578,N_2386,N_2215);
and U2579 (N_2579,N_2314,N_2337);
or U2580 (N_2580,N_2362,N_2391);
or U2581 (N_2581,N_2397,N_2334);
and U2582 (N_2582,N_2354,N_2342);
nor U2583 (N_2583,N_2262,N_2367);
nor U2584 (N_2584,N_2343,N_2257);
xnor U2585 (N_2585,N_2286,N_2313);
and U2586 (N_2586,N_2305,N_2312);
nor U2587 (N_2587,N_2378,N_2329);
or U2588 (N_2588,N_2384,N_2242);
or U2589 (N_2589,N_2377,N_2238);
and U2590 (N_2590,N_2369,N_2318);
nor U2591 (N_2591,N_2315,N_2371);
and U2592 (N_2592,N_2217,N_2296);
or U2593 (N_2593,N_2390,N_2375);
or U2594 (N_2594,N_2316,N_2339);
nor U2595 (N_2595,N_2293,N_2289);
nor U2596 (N_2596,N_2214,N_2309);
and U2597 (N_2597,N_2279,N_2282);
or U2598 (N_2598,N_2313,N_2362);
or U2599 (N_2599,N_2276,N_2393);
nand U2600 (N_2600,N_2474,N_2413);
or U2601 (N_2601,N_2552,N_2458);
nor U2602 (N_2602,N_2476,N_2566);
nand U2603 (N_2603,N_2526,N_2439);
or U2604 (N_2604,N_2466,N_2497);
nor U2605 (N_2605,N_2480,N_2455);
and U2606 (N_2606,N_2522,N_2503);
or U2607 (N_2607,N_2578,N_2479);
or U2608 (N_2608,N_2547,N_2470);
and U2609 (N_2609,N_2471,N_2440);
or U2610 (N_2610,N_2417,N_2537);
and U2611 (N_2611,N_2530,N_2441);
and U2612 (N_2612,N_2478,N_2412);
nand U2613 (N_2613,N_2505,N_2502);
or U2614 (N_2614,N_2434,N_2457);
or U2615 (N_2615,N_2475,N_2557);
or U2616 (N_2616,N_2533,N_2499);
xor U2617 (N_2617,N_2542,N_2546);
nand U2618 (N_2618,N_2524,N_2583);
nand U2619 (N_2619,N_2482,N_2445);
or U2620 (N_2620,N_2550,N_2421);
nand U2621 (N_2621,N_2536,N_2450);
or U2622 (N_2622,N_2477,N_2443);
and U2623 (N_2623,N_2428,N_2459);
nor U2624 (N_2624,N_2405,N_2464);
or U2625 (N_2625,N_2461,N_2563);
and U2626 (N_2626,N_2518,N_2535);
nand U2627 (N_2627,N_2565,N_2548);
or U2628 (N_2628,N_2506,N_2594);
or U2629 (N_2629,N_2574,N_2510);
nor U2630 (N_2630,N_2593,N_2473);
nand U2631 (N_2631,N_2415,N_2483);
or U2632 (N_2632,N_2467,N_2418);
and U2633 (N_2633,N_2597,N_2484);
or U2634 (N_2634,N_2519,N_2579);
nand U2635 (N_2635,N_2512,N_2487);
or U2636 (N_2636,N_2521,N_2433);
and U2637 (N_2637,N_2426,N_2488);
nand U2638 (N_2638,N_2504,N_2481);
or U2639 (N_2639,N_2493,N_2581);
or U2640 (N_2640,N_2584,N_2465);
nand U2641 (N_2641,N_2525,N_2419);
or U2642 (N_2642,N_2402,N_2486);
or U2643 (N_2643,N_2490,N_2437);
nor U2644 (N_2644,N_2589,N_2453);
nor U2645 (N_2645,N_2569,N_2575);
nand U2646 (N_2646,N_2553,N_2400);
or U2647 (N_2647,N_2409,N_2407);
nor U2648 (N_2648,N_2410,N_2534);
or U2649 (N_2649,N_2401,N_2411);
and U2650 (N_2650,N_2585,N_2501);
or U2651 (N_2651,N_2564,N_2436);
xor U2652 (N_2652,N_2424,N_2496);
or U2653 (N_2653,N_2460,N_2591);
nand U2654 (N_2654,N_2442,N_2554);
and U2655 (N_2655,N_2427,N_2572);
nor U2656 (N_2656,N_2551,N_2447);
or U2657 (N_2657,N_2529,N_2491);
and U2658 (N_2658,N_2543,N_2446);
or U2659 (N_2659,N_2549,N_2573);
nor U2660 (N_2660,N_2500,N_2562);
or U2661 (N_2661,N_2570,N_2580);
xor U2662 (N_2662,N_2590,N_2523);
nor U2663 (N_2663,N_2539,N_2598);
nand U2664 (N_2664,N_2452,N_2462);
nor U2665 (N_2665,N_2599,N_2485);
nand U2666 (N_2666,N_2469,N_2438);
nand U2667 (N_2667,N_2408,N_2404);
nor U2668 (N_2668,N_2596,N_2507);
nand U2669 (N_2669,N_2527,N_2449);
and U2670 (N_2670,N_2406,N_2444);
or U2671 (N_2671,N_2516,N_2538);
nand U2672 (N_2672,N_2513,N_2498);
or U2673 (N_2673,N_2448,N_2414);
or U2674 (N_2674,N_2511,N_2541);
or U2675 (N_2675,N_2425,N_2432);
and U2676 (N_2676,N_2514,N_2508);
and U2677 (N_2677,N_2472,N_2509);
or U2678 (N_2678,N_2588,N_2545);
or U2679 (N_2679,N_2528,N_2451);
nor U2680 (N_2680,N_2456,N_2463);
nor U2681 (N_2681,N_2423,N_2586);
nor U2682 (N_2682,N_2592,N_2515);
or U2683 (N_2683,N_2544,N_2422);
nand U2684 (N_2684,N_2489,N_2559);
nor U2685 (N_2685,N_2435,N_2420);
or U2686 (N_2686,N_2561,N_2556);
and U2687 (N_2687,N_2532,N_2431);
nand U2688 (N_2688,N_2454,N_2571);
and U2689 (N_2689,N_2595,N_2568);
nand U2690 (N_2690,N_2517,N_2582);
nor U2691 (N_2691,N_2587,N_2576);
nor U2692 (N_2692,N_2577,N_2494);
and U2693 (N_2693,N_2540,N_2430);
nor U2694 (N_2694,N_2558,N_2520);
nand U2695 (N_2695,N_2429,N_2468);
nor U2696 (N_2696,N_2560,N_2531);
xnor U2697 (N_2697,N_2555,N_2403);
or U2698 (N_2698,N_2495,N_2492);
and U2699 (N_2699,N_2416,N_2567);
and U2700 (N_2700,N_2572,N_2574);
nand U2701 (N_2701,N_2423,N_2402);
nand U2702 (N_2702,N_2537,N_2560);
nand U2703 (N_2703,N_2587,N_2509);
and U2704 (N_2704,N_2564,N_2550);
nor U2705 (N_2705,N_2593,N_2426);
nand U2706 (N_2706,N_2509,N_2481);
and U2707 (N_2707,N_2402,N_2584);
and U2708 (N_2708,N_2435,N_2561);
and U2709 (N_2709,N_2462,N_2598);
and U2710 (N_2710,N_2563,N_2569);
or U2711 (N_2711,N_2598,N_2538);
nor U2712 (N_2712,N_2578,N_2433);
and U2713 (N_2713,N_2526,N_2555);
nand U2714 (N_2714,N_2588,N_2597);
nand U2715 (N_2715,N_2431,N_2424);
nand U2716 (N_2716,N_2538,N_2557);
and U2717 (N_2717,N_2588,N_2563);
nor U2718 (N_2718,N_2574,N_2550);
nor U2719 (N_2719,N_2565,N_2421);
and U2720 (N_2720,N_2512,N_2428);
nand U2721 (N_2721,N_2436,N_2539);
or U2722 (N_2722,N_2569,N_2520);
nand U2723 (N_2723,N_2441,N_2560);
nor U2724 (N_2724,N_2570,N_2583);
or U2725 (N_2725,N_2566,N_2434);
nor U2726 (N_2726,N_2457,N_2516);
nor U2727 (N_2727,N_2534,N_2472);
or U2728 (N_2728,N_2568,N_2579);
or U2729 (N_2729,N_2498,N_2575);
or U2730 (N_2730,N_2480,N_2477);
nor U2731 (N_2731,N_2474,N_2489);
nand U2732 (N_2732,N_2458,N_2482);
and U2733 (N_2733,N_2557,N_2417);
nor U2734 (N_2734,N_2446,N_2539);
nor U2735 (N_2735,N_2428,N_2418);
and U2736 (N_2736,N_2433,N_2575);
nor U2737 (N_2737,N_2507,N_2514);
nand U2738 (N_2738,N_2566,N_2454);
nand U2739 (N_2739,N_2569,N_2537);
nand U2740 (N_2740,N_2475,N_2542);
or U2741 (N_2741,N_2422,N_2402);
nor U2742 (N_2742,N_2541,N_2509);
or U2743 (N_2743,N_2495,N_2481);
nand U2744 (N_2744,N_2590,N_2516);
nand U2745 (N_2745,N_2575,N_2528);
nor U2746 (N_2746,N_2445,N_2532);
nor U2747 (N_2747,N_2512,N_2468);
or U2748 (N_2748,N_2459,N_2434);
nand U2749 (N_2749,N_2465,N_2493);
and U2750 (N_2750,N_2516,N_2439);
nor U2751 (N_2751,N_2468,N_2443);
or U2752 (N_2752,N_2546,N_2488);
and U2753 (N_2753,N_2430,N_2574);
and U2754 (N_2754,N_2580,N_2450);
or U2755 (N_2755,N_2438,N_2499);
and U2756 (N_2756,N_2455,N_2436);
nor U2757 (N_2757,N_2490,N_2403);
or U2758 (N_2758,N_2519,N_2415);
or U2759 (N_2759,N_2480,N_2501);
or U2760 (N_2760,N_2597,N_2413);
nand U2761 (N_2761,N_2466,N_2553);
or U2762 (N_2762,N_2484,N_2422);
nor U2763 (N_2763,N_2468,N_2527);
or U2764 (N_2764,N_2406,N_2452);
nand U2765 (N_2765,N_2537,N_2585);
nor U2766 (N_2766,N_2543,N_2463);
or U2767 (N_2767,N_2552,N_2541);
and U2768 (N_2768,N_2417,N_2435);
nand U2769 (N_2769,N_2543,N_2483);
or U2770 (N_2770,N_2472,N_2491);
nor U2771 (N_2771,N_2510,N_2543);
or U2772 (N_2772,N_2496,N_2578);
or U2773 (N_2773,N_2420,N_2491);
or U2774 (N_2774,N_2599,N_2577);
and U2775 (N_2775,N_2435,N_2530);
nand U2776 (N_2776,N_2522,N_2484);
nor U2777 (N_2777,N_2582,N_2400);
or U2778 (N_2778,N_2508,N_2405);
or U2779 (N_2779,N_2511,N_2596);
or U2780 (N_2780,N_2467,N_2469);
and U2781 (N_2781,N_2526,N_2456);
nand U2782 (N_2782,N_2526,N_2451);
nor U2783 (N_2783,N_2561,N_2465);
or U2784 (N_2784,N_2548,N_2409);
nor U2785 (N_2785,N_2460,N_2506);
nand U2786 (N_2786,N_2465,N_2553);
or U2787 (N_2787,N_2552,N_2481);
or U2788 (N_2788,N_2557,N_2434);
nand U2789 (N_2789,N_2483,N_2508);
nor U2790 (N_2790,N_2443,N_2486);
and U2791 (N_2791,N_2533,N_2569);
nand U2792 (N_2792,N_2502,N_2433);
xor U2793 (N_2793,N_2566,N_2577);
or U2794 (N_2794,N_2454,N_2434);
nor U2795 (N_2795,N_2478,N_2527);
xor U2796 (N_2796,N_2460,N_2540);
nor U2797 (N_2797,N_2488,N_2584);
or U2798 (N_2798,N_2476,N_2591);
and U2799 (N_2799,N_2464,N_2449);
nand U2800 (N_2800,N_2626,N_2756);
nor U2801 (N_2801,N_2737,N_2632);
and U2802 (N_2802,N_2783,N_2667);
nor U2803 (N_2803,N_2779,N_2746);
nor U2804 (N_2804,N_2727,N_2630);
or U2805 (N_2805,N_2760,N_2795);
or U2806 (N_2806,N_2697,N_2798);
nand U2807 (N_2807,N_2695,N_2644);
or U2808 (N_2808,N_2732,N_2600);
or U2809 (N_2809,N_2722,N_2637);
nor U2810 (N_2810,N_2750,N_2622);
or U2811 (N_2811,N_2789,N_2650);
or U2812 (N_2812,N_2742,N_2743);
or U2813 (N_2813,N_2683,N_2786);
nand U2814 (N_2814,N_2726,N_2645);
nor U2815 (N_2815,N_2604,N_2755);
nor U2816 (N_2816,N_2734,N_2671);
nor U2817 (N_2817,N_2649,N_2691);
or U2818 (N_2818,N_2670,N_2723);
nor U2819 (N_2819,N_2762,N_2716);
nand U2820 (N_2820,N_2784,N_2769);
and U2821 (N_2821,N_2654,N_2617);
or U2822 (N_2822,N_2793,N_2614);
nor U2823 (N_2823,N_2694,N_2741);
or U2824 (N_2824,N_2688,N_2763);
nand U2825 (N_2825,N_2752,N_2773);
or U2826 (N_2826,N_2736,N_2674);
nor U2827 (N_2827,N_2663,N_2747);
or U2828 (N_2828,N_2796,N_2687);
nand U2829 (N_2829,N_2635,N_2680);
xnor U2830 (N_2830,N_2767,N_2609);
or U2831 (N_2831,N_2788,N_2754);
nor U2832 (N_2832,N_2704,N_2682);
nor U2833 (N_2833,N_2745,N_2730);
nor U2834 (N_2834,N_2708,N_2748);
and U2835 (N_2835,N_2728,N_2690);
nand U2836 (N_2836,N_2603,N_2761);
nor U2837 (N_2837,N_2648,N_2764);
nor U2838 (N_2838,N_2666,N_2628);
nor U2839 (N_2839,N_2780,N_2735);
nor U2840 (N_2840,N_2787,N_2612);
or U2841 (N_2841,N_2725,N_2794);
nor U2842 (N_2842,N_2608,N_2660);
nand U2843 (N_2843,N_2719,N_2673);
nand U2844 (N_2844,N_2738,N_2729);
and U2845 (N_2845,N_2665,N_2661);
nand U2846 (N_2846,N_2634,N_2631);
nand U2847 (N_2847,N_2679,N_2705);
nor U2848 (N_2848,N_2618,N_2621);
or U2849 (N_2849,N_2771,N_2712);
or U2850 (N_2850,N_2655,N_2790);
nor U2851 (N_2851,N_2636,N_2768);
or U2852 (N_2852,N_2669,N_2781);
nand U2853 (N_2853,N_2785,N_2616);
nor U2854 (N_2854,N_2696,N_2624);
and U2855 (N_2855,N_2757,N_2642);
and U2856 (N_2856,N_2689,N_2797);
nand U2857 (N_2857,N_2611,N_2646);
nor U2858 (N_2858,N_2692,N_2676);
or U2859 (N_2859,N_2700,N_2657);
or U2860 (N_2860,N_2721,N_2610);
or U2861 (N_2861,N_2638,N_2629);
nand U2862 (N_2862,N_2792,N_2703);
nor U2863 (N_2863,N_2759,N_2765);
nor U2864 (N_2864,N_2711,N_2739);
xnor U2865 (N_2865,N_2684,N_2772);
nor U2866 (N_2866,N_2633,N_2685);
or U2867 (N_2867,N_2686,N_2625);
or U2868 (N_2868,N_2643,N_2623);
nand U2869 (N_2869,N_2799,N_2620);
nor U2870 (N_2870,N_2702,N_2774);
nor U2871 (N_2871,N_2777,N_2677);
nor U2872 (N_2872,N_2652,N_2775);
and U2873 (N_2873,N_2653,N_2641);
nand U2874 (N_2874,N_2602,N_2718);
nand U2875 (N_2875,N_2675,N_2601);
and U2876 (N_2876,N_2707,N_2693);
nand U2877 (N_2877,N_2651,N_2672);
and U2878 (N_2878,N_2751,N_2758);
nor U2879 (N_2879,N_2766,N_2782);
nand U2880 (N_2880,N_2659,N_2744);
nand U2881 (N_2881,N_2713,N_2733);
or U2882 (N_2882,N_2619,N_2605);
nor U2883 (N_2883,N_2668,N_2778);
or U2884 (N_2884,N_2640,N_2740);
and U2885 (N_2885,N_2699,N_2749);
nand U2886 (N_2886,N_2715,N_2698);
and U2887 (N_2887,N_2658,N_2613);
nor U2888 (N_2888,N_2606,N_2681);
and U2889 (N_2889,N_2615,N_2717);
nand U2890 (N_2890,N_2753,N_2664);
nand U2891 (N_2891,N_2709,N_2776);
nand U2892 (N_2892,N_2701,N_2710);
or U2893 (N_2893,N_2706,N_2607);
and U2894 (N_2894,N_2724,N_2770);
nor U2895 (N_2895,N_2647,N_2791);
and U2896 (N_2896,N_2720,N_2627);
nand U2897 (N_2897,N_2656,N_2731);
nand U2898 (N_2898,N_2639,N_2678);
and U2899 (N_2899,N_2662,N_2714);
or U2900 (N_2900,N_2600,N_2770);
or U2901 (N_2901,N_2755,N_2743);
and U2902 (N_2902,N_2765,N_2643);
nor U2903 (N_2903,N_2734,N_2602);
and U2904 (N_2904,N_2792,N_2649);
or U2905 (N_2905,N_2644,N_2765);
nand U2906 (N_2906,N_2699,N_2797);
or U2907 (N_2907,N_2670,N_2660);
and U2908 (N_2908,N_2784,N_2620);
nor U2909 (N_2909,N_2741,N_2742);
nand U2910 (N_2910,N_2727,N_2617);
nand U2911 (N_2911,N_2617,N_2793);
nand U2912 (N_2912,N_2622,N_2717);
or U2913 (N_2913,N_2733,N_2710);
and U2914 (N_2914,N_2715,N_2712);
or U2915 (N_2915,N_2605,N_2775);
and U2916 (N_2916,N_2798,N_2646);
nor U2917 (N_2917,N_2717,N_2796);
or U2918 (N_2918,N_2765,N_2748);
nor U2919 (N_2919,N_2766,N_2694);
or U2920 (N_2920,N_2622,N_2742);
and U2921 (N_2921,N_2706,N_2721);
nand U2922 (N_2922,N_2660,N_2728);
and U2923 (N_2923,N_2749,N_2736);
nor U2924 (N_2924,N_2755,N_2710);
nand U2925 (N_2925,N_2636,N_2717);
or U2926 (N_2926,N_2703,N_2659);
nor U2927 (N_2927,N_2772,N_2721);
or U2928 (N_2928,N_2781,N_2711);
and U2929 (N_2929,N_2687,N_2600);
nor U2930 (N_2930,N_2620,N_2733);
or U2931 (N_2931,N_2797,N_2633);
or U2932 (N_2932,N_2697,N_2762);
nand U2933 (N_2933,N_2690,N_2618);
nor U2934 (N_2934,N_2628,N_2710);
nor U2935 (N_2935,N_2615,N_2651);
and U2936 (N_2936,N_2700,N_2774);
nand U2937 (N_2937,N_2736,N_2765);
or U2938 (N_2938,N_2744,N_2610);
and U2939 (N_2939,N_2659,N_2740);
or U2940 (N_2940,N_2660,N_2720);
nand U2941 (N_2941,N_2658,N_2639);
nand U2942 (N_2942,N_2600,N_2787);
nor U2943 (N_2943,N_2707,N_2746);
nor U2944 (N_2944,N_2725,N_2610);
or U2945 (N_2945,N_2667,N_2618);
nor U2946 (N_2946,N_2759,N_2716);
or U2947 (N_2947,N_2798,N_2608);
nand U2948 (N_2948,N_2777,N_2714);
nor U2949 (N_2949,N_2678,N_2636);
or U2950 (N_2950,N_2652,N_2797);
and U2951 (N_2951,N_2719,N_2660);
or U2952 (N_2952,N_2715,N_2667);
nor U2953 (N_2953,N_2760,N_2711);
nor U2954 (N_2954,N_2622,N_2674);
or U2955 (N_2955,N_2688,N_2615);
nand U2956 (N_2956,N_2615,N_2687);
and U2957 (N_2957,N_2756,N_2707);
nor U2958 (N_2958,N_2716,N_2681);
nand U2959 (N_2959,N_2714,N_2667);
or U2960 (N_2960,N_2723,N_2640);
or U2961 (N_2961,N_2767,N_2754);
nor U2962 (N_2962,N_2679,N_2720);
and U2963 (N_2963,N_2647,N_2728);
and U2964 (N_2964,N_2799,N_2723);
or U2965 (N_2965,N_2794,N_2690);
and U2966 (N_2966,N_2611,N_2661);
nor U2967 (N_2967,N_2761,N_2776);
nand U2968 (N_2968,N_2616,N_2726);
nand U2969 (N_2969,N_2676,N_2698);
and U2970 (N_2970,N_2639,N_2724);
or U2971 (N_2971,N_2713,N_2695);
or U2972 (N_2972,N_2632,N_2726);
nand U2973 (N_2973,N_2669,N_2654);
or U2974 (N_2974,N_2763,N_2744);
nor U2975 (N_2975,N_2720,N_2656);
nand U2976 (N_2976,N_2721,N_2692);
and U2977 (N_2977,N_2652,N_2767);
or U2978 (N_2978,N_2743,N_2731);
or U2979 (N_2979,N_2730,N_2771);
nor U2980 (N_2980,N_2781,N_2720);
nor U2981 (N_2981,N_2652,N_2600);
and U2982 (N_2982,N_2749,N_2632);
nand U2983 (N_2983,N_2633,N_2753);
nor U2984 (N_2984,N_2630,N_2789);
nand U2985 (N_2985,N_2765,N_2792);
nand U2986 (N_2986,N_2753,N_2623);
and U2987 (N_2987,N_2695,N_2770);
or U2988 (N_2988,N_2666,N_2768);
or U2989 (N_2989,N_2782,N_2742);
or U2990 (N_2990,N_2657,N_2787);
nand U2991 (N_2991,N_2748,N_2614);
nor U2992 (N_2992,N_2788,N_2616);
or U2993 (N_2993,N_2748,N_2652);
and U2994 (N_2994,N_2625,N_2684);
nor U2995 (N_2995,N_2779,N_2693);
and U2996 (N_2996,N_2615,N_2654);
nor U2997 (N_2997,N_2724,N_2650);
or U2998 (N_2998,N_2649,N_2739);
or U2999 (N_2999,N_2737,N_2668);
nand U3000 (N_3000,N_2996,N_2823);
and U3001 (N_3001,N_2840,N_2859);
xor U3002 (N_3002,N_2941,N_2848);
or U3003 (N_3003,N_2993,N_2808);
nor U3004 (N_3004,N_2990,N_2952);
and U3005 (N_3005,N_2901,N_2869);
or U3006 (N_3006,N_2915,N_2992);
nor U3007 (N_3007,N_2893,N_2944);
nand U3008 (N_3008,N_2966,N_2889);
and U3009 (N_3009,N_2972,N_2853);
or U3010 (N_3010,N_2846,N_2958);
nor U3011 (N_3011,N_2877,N_2898);
nor U3012 (N_3012,N_2805,N_2986);
and U3013 (N_3013,N_2912,N_2997);
and U3014 (N_3014,N_2994,N_2922);
or U3015 (N_3015,N_2890,N_2904);
or U3016 (N_3016,N_2902,N_2978);
or U3017 (N_3017,N_2943,N_2973);
or U3018 (N_3018,N_2892,N_2850);
or U3019 (N_3019,N_2878,N_2903);
and U3020 (N_3020,N_2825,N_2933);
xnor U3021 (N_3021,N_2905,N_2935);
or U3022 (N_3022,N_2842,N_2959);
xor U3023 (N_3023,N_2860,N_2862);
or U3024 (N_3024,N_2880,N_2955);
nor U3025 (N_3025,N_2951,N_2866);
nand U3026 (N_3026,N_2836,N_2907);
or U3027 (N_3027,N_2995,N_2984);
nand U3028 (N_3028,N_2855,N_2948);
nand U3029 (N_3029,N_2830,N_2826);
and U3030 (N_3030,N_2977,N_2974);
nor U3031 (N_3031,N_2954,N_2945);
and U3032 (N_3032,N_2926,N_2818);
and U3033 (N_3033,N_2932,N_2835);
nor U3034 (N_3034,N_2983,N_2810);
nand U3035 (N_3035,N_2987,N_2950);
or U3036 (N_3036,N_2806,N_2828);
nand U3037 (N_3037,N_2916,N_2971);
or U3038 (N_3038,N_2815,N_2968);
and U3039 (N_3039,N_2949,N_2947);
and U3040 (N_3040,N_2938,N_2852);
nor U3041 (N_3041,N_2851,N_2864);
and U3042 (N_3042,N_2969,N_2875);
or U3043 (N_3043,N_2980,N_2876);
and U3044 (N_3044,N_2834,N_2849);
and U3045 (N_3045,N_2942,N_2865);
nand U3046 (N_3046,N_2924,N_2881);
xnor U3047 (N_3047,N_2988,N_2920);
nand U3048 (N_3048,N_2991,N_2923);
nor U3049 (N_3049,N_2837,N_2801);
nand U3050 (N_3050,N_2970,N_2913);
nand U3051 (N_3051,N_2940,N_2857);
or U3052 (N_3052,N_2804,N_2999);
and U3053 (N_3053,N_2900,N_2819);
nand U3054 (N_3054,N_2975,N_2817);
nand U3055 (N_3055,N_2831,N_2931);
or U3056 (N_3056,N_2939,N_2946);
and U3057 (N_3057,N_2976,N_2800);
and U3058 (N_3058,N_2919,N_2824);
or U3059 (N_3059,N_2909,N_2841);
and U3060 (N_3060,N_2989,N_2921);
or U3061 (N_3061,N_2927,N_2872);
or U3062 (N_3062,N_2809,N_2807);
nor U3063 (N_3063,N_2908,N_2888);
nand U3064 (N_3064,N_2879,N_2873);
nor U3065 (N_3065,N_2930,N_2833);
nor U3066 (N_3066,N_2967,N_2963);
nand U3067 (N_3067,N_2979,N_2937);
and U3068 (N_3068,N_2917,N_2839);
nand U3069 (N_3069,N_2925,N_2936);
nand U3070 (N_3070,N_2914,N_2934);
or U3071 (N_3071,N_2845,N_2812);
and U3072 (N_3072,N_2802,N_2961);
or U3073 (N_3073,N_2870,N_2957);
and U3074 (N_3074,N_2962,N_2832);
nand U3075 (N_3075,N_2897,N_2882);
nor U3076 (N_3076,N_2891,N_2803);
nand U3077 (N_3077,N_2953,N_2811);
nand U3078 (N_3078,N_2887,N_2985);
nor U3079 (N_3079,N_2854,N_2816);
or U3080 (N_3080,N_2960,N_2827);
nand U3081 (N_3081,N_2883,N_2910);
nand U3082 (N_3082,N_2884,N_2886);
or U3083 (N_3083,N_2894,N_2929);
or U3084 (N_3084,N_2928,N_2822);
nand U3085 (N_3085,N_2868,N_2965);
or U3086 (N_3086,N_2896,N_2885);
nand U3087 (N_3087,N_2844,N_2871);
nand U3088 (N_3088,N_2847,N_2956);
nand U3089 (N_3089,N_2998,N_2820);
nor U3090 (N_3090,N_2829,N_2821);
and U3091 (N_3091,N_2856,N_2843);
nor U3092 (N_3092,N_2838,N_2906);
and U3093 (N_3093,N_2981,N_2918);
nand U3094 (N_3094,N_2858,N_2911);
nor U3095 (N_3095,N_2964,N_2861);
and U3096 (N_3096,N_2813,N_2895);
nor U3097 (N_3097,N_2814,N_2899);
or U3098 (N_3098,N_2867,N_2863);
nand U3099 (N_3099,N_2874,N_2982);
nor U3100 (N_3100,N_2877,N_2830);
nor U3101 (N_3101,N_2870,N_2807);
nor U3102 (N_3102,N_2874,N_2887);
nor U3103 (N_3103,N_2902,N_2873);
and U3104 (N_3104,N_2918,N_2877);
xor U3105 (N_3105,N_2810,N_2957);
nor U3106 (N_3106,N_2933,N_2987);
nand U3107 (N_3107,N_2995,N_2862);
nand U3108 (N_3108,N_2871,N_2901);
nor U3109 (N_3109,N_2820,N_2876);
nor U3110 (N_3110,N_2934,N_2966);
and U3111 (N_3111,N_2948,N_2845);
nand U3112 (N_3112,N_2824,N_2923);
and U3113 (N_3113,N_2844,N_2812);
nand U3114 (N_3114,N_2952,N_2837);
or U3115 (N_3115,N_2966,N_2841);
nor U3116 (N_3116,N_2830,N_2855);
or U3117 (N_3117,N_2823,N_2861);
nand U3118 (N_3118,N_2932,N_2955);
or U3119 (N_3119,N_2923,N_2987);
nand U3120 (N_3120,N_2917,N_2971);
and U3121 (N_3121,N_2855,N_2961);
or U3122 (N_3122,N_2935,N_2849);
and U3123 (N_3123,N_2864,N_2923);
or U3124 (N_3124,N_2837,N_2922);
nor U3125 (N_3125,N_2925,N_2849);
nand U3126 (N_3126,N_2985,N_2914);
nor U3127 (N_3127,N_2995,N_2857);
xor U3128 (N_3128,N_2867,N_2902);
nor U3129 (N_3129,N_2832,N_2910);
nand U3130 (N_3130,N_2868,N_2827);
or U3131 (N_3131,N_2957,N_2925);
nor U3132 (N_3132,N_2849,N_2807);
nand U3133 (N_3133,N_2846,N_2849);
nand U3134 (N_3134,N_2870,N_2851);
nand U3135 (N_3135,N_2891,N_2882);
or U3136 (N_3136,N_2986,N_2947);
nand U3137 (N_3137,N_2992,N_2960);
or U3138 (N_3138,N_2828,N_2958);
or U3139 (N_3139,N_2808,N_2824);
nor U3140 (N_3140,N_2976,N_2957);
nand U3141 (N_3141,N_2801,N_2807);
or U3142 (N_3142,N_2914,N_2831);
and U3143 (N_3143,N_2803,N_2824);
or U3144 (N_3144,N_2978,N_2841);
nand U3145 (N_3145,N_2996,N_2864);
or U3146 (N_3146,N_2906,N_2948);
and U3147 (N_3147,N_2810,N_2803);
or U3148 (N_3148,N_2825,N_2972);
nor U3149 (N_3149,N_2920,N_2944);
nor U3150 (N_3150,N_2908,N_2900);
nand U3151 (N_3151,N_2925,N_2864);
and U3152 (N_3152,N_2860,N_2815);
nor U3153 (N_3153,N_2812,N_2879);
and U3154 (N_3154,N_2847,N_2890);
or U3155 (N_3155,N_2863,N_2946);
or U3156 (N_3156,N_2962,N_2972);
nor U3157 (N_3157,N_2931,N_2850);
or U3158 (N_3158,N_2887,N_2814);
nand U3159 (N_3159,N_2941,N_2983);
nand U3160 (N_3160,N_2981,N_2895);
nor U3161 (N_3161,N_2864,N_2891);
and U3162 (N_3162,N_2914,N_2999);
nor U3163 (N_3163,N_2956,N_2867);
nand U3164 (N_3164,N_2943,N_2900);
nor U3165 (N_3165,N_2902,N_2897);
nor U3166 (N_3166,N_2922,N_2972);
xnor U3167 (N_3167,N_2820,N_2930);
nand U3168 (N_3168,N_2883,N_2879);
nor U3169 (N_3169,N_2897,N_2861);
nor U3170 (N_3170,N_2887,N_2998);
and U3171 (N_3171,N_2825,N_2877);
or U3172 (N_3172,N_2892,N_2813);
nand U3173 (N_3173,N_2990,N_2825);
and U3174 (N_3174,N_2980,N_2842);
nor U3175 (N_3175,N_2899,N_2848);
nand U3176 (N_3176,N_2932,N_2875);
nor U3177 (N_3177,N_2984,N_2915);
nand U3178 (N_3178,N_2935,N_2917);
nor U3179 (N_3179,N_2895,N_2850);
and U3180 (N_3180,N_2857,N_2890);
or U3181 (N_3181,N_2820,N_2978);
or U3182 (N_3182,N_2917,N_2953);
or U3183 (N_3183,N_2927,N_2909);
and U3184 (N_3184,N_2889,N_2859);
nor U3185 (N_3185,N_2970,N_2951);
or U3186 (N_3186,N_2820,N_2814);
nor U3187 (N_3187,N_2827,N_2977);
and U3188 (N_3188,N_2849,N_2907);
nand U3189 (N_3189,N_2988,N_2933);
or U3190 (N_3190,N_2859,N_2863);
nand U3191 (N_3191,N_2939,N_2916);
or U3192 (N_3192,N_2893,N_2835);
or U3193 (N_3193,N_2909,N_2903);
or U3194 (N_3194,N_2872,N_2841);
or U3195 (N_3195,N_2896,N_2807);
or U3196 (N_3196,N_2934,N_2832);
nor U3197 (N_3197,N_2830,N_2990);
nand U3198 (N_3198,N_2858,N_2928);
nor U3199 (N_3199,N_2922,N_2970);
nor U3200 (N_3200,N_3150,N_3166);
nand U3201 (N_3201,N_3039,N_3007);
nor U3202 (N_3202,N_3187,N_3096);
nor U3203 (N_3203,N_3000,N_3161);
nand U3204 (N_3204,N_3192,N_3031);
nor U3205 (N_3205,N_3181,N_3127);
or U3206 (N_3206,N_3160,N_3151);
or U3207 (N_3207,N_3041,N_3020);
or U3208 (N_3208,N_3018,N_3042);
and U3209 (N_3209,N_3143,N_3063);
nor U3210 (N_3210,N_3112,N_3065);
or U3211 (N_3211,N_3129,N_3074);
nor U3212 (N_3212,N_3009,N_3076);
nor U3213 (N_3213,N_3088,N_3109);
and U3214 (N_3214,N_3064,N_3040);
nand U3215 (N_3215,N_3106,N_3053);
nand U3216 (N_3216,N_3101,N_3177);
nor U3217 (N_3217,N_3061,N_3144);
or U3218 (N_3218,N_3196,N_3117);
nand U3219 (N_3219,N_3170,N_3059);
nand U3220 (N_3220,N_3026,N_3176);
nor U3221 (N_3221,N_3068,N_3149);
nor U3222 (N_3222,N_3029,N_3189);
nand U3223 (N_3223,N_3111,N_3071);
nor U3224 (N_3224,N_3054,N_3139);
nand U3225 (N_3225,N_3125,N_3008);
and U3226 (N_3226,N_3168,N_3001);
or U3227 (N_3227,N_3186,N_3121);
and U3228 (N_3228,N_3102,N_3021);
nor U3229 (N_3229,N_3091,N_3138);
or U3230 (N_3230,N_3037,N_3077);
nor U3231 (N_3231,N_3157,N_3052);
and U3232 (N_3232,N_3123,N_3055);
nand U3233 (N_3233,N_3067,N_3045);
and U3234 (N_3234,N_3162,N_3058);
and U3235 (N_3235,N_3056,N_3155);
nor U3236 (N_3236,N_3093,N_3128);
nand U3237 (N_3237,N_3173,N_3167);
and U3238 (N_3238,N_3133,N_3132);
or U3239 (N_3239,N_3080,N_3022);
nor U3240 (N_3240,N_3158,N_3087);
nand U3241 (N_3241,N_3083,N_3113);
or U3242 (N_3242,N_3038,N_3108);
and U3243 (N_3243,N_3194,N_3156);
nand U3244 (N_3244,N_3146,N_3104);
or U3245 (N_3245,N_3030,N_3005);
nand U3246 (N_3246,N_3193,N_3153);
nor U3247 (N_3247,N_3179,N_3180);
or U3248 (N_3248,N_3062,N_3050);
nor U3249 (N_3249,N_3024,N_3118);
and U3250 (N_3250,N_3142,N_3174);
nand U3251 (N_3251,N_3140,N_3100);
nand U3252 (N_3252,N_3191,N_3164);
nor U3253 (N_3253,N_3044,N_3015);
nor U3254 (N_3254,N_3197,N_3035);
nor U3255 (N_3255,N_3199,N_3122);
nor U3256 (N_3256,N_3114,N_3175);
or U3257 (N_3257,N_3136,N_3027);
nor U3258 (N_3258,N_3060,N_3078);
nand U3259 (N_3259,N_3016,N_3012);
or U3260 (N_3260,N_3032,N_3019);
nand U3261 (N_3261,N_3047,N_3137);
nand U3262 (N_3262,N_3082,N_3002);
and U3263 (N_3263,N_3036,N_3165);
or U3264 (N_3264,N_3075,N_3190);
nor U3265 (N_3265,N_3073,N_3089);
nor U3266 (N_3266,N_3049,N_3171);
nand U3267 (N_3267,N_3198,N_3023);
nand U3268 (N_3268,N_3184,N_3145);
nand U3269 (N_3269,N_3069,N_3110);
nor U3270 (N_3270,N_3195,N_3135);
or U3271 (N_3271,N_3126,N_3163);
or U3272 (N_3272,N_3051,N_3043);
nand U3273 (N_3273,N_3057,N_3034);
and U3274 (N_3274,N_3006,N_3081);
or U3275 (N_3275,N_3033,N_3086);
nand U3276 (N_3276,N_3103,N_3141);
nor U3277 (N_3277,N_3028,N_3154);
and U3278 (N_3278,N_3084,N_3079);
nand U3279 (N_3279,N_3014,N_3119);
and U3280 (N_3280,N_3159,N_3172);
nor U3281 (N_3281,N_3124,N_3099);
nor U3282 (N_3282,N_3120,N_3098);
or U3283 (N_3283,N_3169,N_3066);
or U3284 (N_3284,N_3090,N_3134);
or U3285 (N_3285,N_3010,N_3048);
or U3286 (N_3286,N_3085,N_3152);
or U3287 (N_3287,N_3131,N_3011);
or U3288 (N_3288,N_3046,N_3178);
nand U3289 (N_3289,N_3092,N_3116);
or U3290 (N_3290,N_3095,N_3185);
nand U3291 (N_3291,N_3107,N_3182);
or U3292 (N_3292,N_3183,N_3097);
or U3293 (N_3293,N_3188,N_3072);
xor U3294 (N_3294,N_3094,N_3013);
nand U3295 (N_3295,N_3105,N_3003);
or U3296 (N_3296,N_3115,N_3025);
nor U3297 (N_3297,N_3148,N_3004);
xor U3298 (N_3298,N_3147,N_3070);
nand U3299 (N_3299,N_3017,N_3130);
and U3300 (N_3300,N_3167,N_3075);
and U3301 (N_3301,N_3148,N_3121);
nand U3302 (N_3302,N_3076,N_3058);
nor U3303 (N_3303,N_3113,N_3064);
nand U3304 (N_3304,N_3019,N_3011);
nand U3305 (N_3305,N_3161,N_3172);
and U3306 (N_3306,N_3162,N_3077);
nand U3307 (N_3307,N_3111,N_3040);
or U3308 (N_3308,N_3051,N_3012);
nor U3309 (N_3309,N_3020,N_3097);
nor U3310 (N_3310,N_3074,N_3139);
and U3311 (N_3311,N_3078,N_3191);
nor U3312 (N_3312,N_3160,N_3133);
and U3313 (N_3313,N_3133,N_3076);
or U3314 (N_3314,N_3116,N_3097);
and U3315 (N_3315,N_3037,N_3108);
nand U3316 (N_3316,N_3078,N_3020);
or U3317 (N_3317,N_3003,N_3139);
nand U3318 (N_3318,N_3004,N_3020);
nand U3319 (N_3319,N_3172,N_3083);
or U3320 (N_3320,N_3185,N_3133);
or U3321 (N_3321,N_3176,N_3154);
and U3322 (N_3322,N_3143,N_3107);
nor U3323 (N_3323,N_3096,N_3052);
nand U3324 (N_3324,N_3164,N_3131);
or U3325 (N_3325,N_3097,N_3031);
and U3326 (N_3326,N_3199,N_3175);
and U3327 (N_3327,N_3105,N_3074);
nor U3328 (N_3328,N_3039,N_3167);
and U3329 (N_3329,N_3123,N_3192);
nand U3330 (N_3330,N_3147,N_3031);
nand U3331 (N_3331,N_3174,N_3053);
nand U3332 (N_3332,N_3105,N_3071);
and U3333 (N_3333,N_3093,N_3048);
nand U3334 (N_3334,N_3008,N_3004);
nor U3335 (N_3335,N_3129,N_3022);
nand U3336 (N_3336,N_3076,N_3039);
nor U3337 (N_3337,N_3062,N_3170);
nand U3338 (N_3338,N_3071,N_3077);
or U3339 (N_3339,N_3172,N_3147);
nand U3340 (N_3340,N_3066,N_3007);
nand U3341 (N_3341,N_3104,N_3172);
and U3342 (N_3342,N_3125,N_3016);
and U3343 (N_3343,N_3154,N_3066);
nor U3344 (N_3344,N_3081,N_3166);
or U3345 (N_3345,N_3179,N_3198);
and U3346 (N_3346,N_3074,N_3112);
or U3347 (N_3347,N_3085,N_3173);
nand U3348 (N_3348,N_3186,N_3065);
and U3349 (N_3349,N_3022,N_3072);
nor U3350 (N_3350,N_3007,N_3080);
and U3351 (N_3351,N_3029,N_3052);
nand U3352 (N_3352,N_3163,N_3004);
xor U3353 (N_3353,N_3027,N_3068);
nor U3354 (N_3354,N_3126,N_3169);
nand U3355 (N_3355,N_3067,N_3032);
nand U3356 (N_3356,N_3130,N_3075);
or U3357 (N_3357,N_3190,N_3123);
or U3358 (N_3358,N_3135,N_3173);
nor U3359 (N_3359,N_3076,N_3103);
nor U3360 (N_3360,N_3063,N_3131);
nand U3361 (N_3361,N_3197,N_3128);
nand U3362 (N_3362,N_3161,N_3110);
and U3363 (N_3363,N_3023,N_3063);
or U3364 (N_3364,N_3009,N_3074);
and U3365 (N_3365,N_3158,N_3044);
and U3366 (N_3366,N_3031,N_3189);
nor U3367 (N_3367,N_3158,N_3071);
and U3368 (N_3368,N_3105,N_3130);
or U3369 (N_3369,N_3141,N_3073);
nor U3370 (N_3370,N_3189,N_3081);
or U3371 (N_3371,N_3056,N_3013);
or U3372 (N_3372,N_3090,N_3136);
and U3373 (N_3373,N_3192,N_3054);
nor U3374 (N_3374,N_3043,N_3192);
or U3375 (N_3375,N_3101,N_3041);
nor U3376 (N_3376,N_3183,N_3161);
nand U3377 (N_3377,N_3135,N_3023);
nor U3378 (N_3378,N_3057,N_3161);
nor U3379 (N_3379,N_3017,N_3049);
nand U3380 (N_3380,N_3096,N_3160);
or U3381 (N_3381,N_3167,N_3193);
and U3382 (N_3382,N_3195,N_3082);
nand U3383 (N_3383,N_3085,N_3136);
or U3384 (N_3384,N_3090,N_3152);
nor U3385 (N_3385,N_3084,N_3001);
nor U3386 (N_3386,N_3149,N_3006);
nor U3387 (N_3387,N_3048,N_3193);
nand U3388 (N_3388,N_3199,N_3058);
or U3389 (N_3389,N_3005,N_3032);
nand U3390 (N_3390,N_3077,N_3055);
nor U3391 (N_3391,N_3058,N_3178);
nand U3392 (N_3392,N_3046,N_3042);
and U3393 (N_3393,N_3146,N_3016);
nor U3394 (N_3394,N_3122,N_3191);
nor U3395 (N_3395,N_3087,N_3148);
nor U3396 (N_3396,N_3138,N_3003);
nand U3397 (N_3397,N_3033,N_3197);
nor U3398 (N_3398,N_3165,N_3110);
nand U3399 (N_3399,N_3123,N_3156);
or U3400 (N_3400,N_3255,N_3264);
and U3401 (N_3401,N_3318,N_3238);
and U3402 (N_3402,N_3258,N_3299);
and U3403 (N_3403,N_3208,N_3274);
or U3404 (N_3404,N_3213,N_3362);
and U3405 (N_3405,N_3314,N_3350);
or U3406 (N_3406,N_3239,N_3306);
or U3407 (N_3407,N_3374,N_3376);
nor U3408 (N_3408,N_3226,N_3300);
nor U3409 (N_3409,N_3364,N_3331);
or U3410 (N_3410,N_3246,N_3220);
nor U3411 (N_3411,N_3349,N_3269);
and U3412 (N_3412,N_3295,N_3293);
nor U3413 (N_3413,N_3320,N_3347);
nand U3414 (N_3414,N_3273,N_3242);
and U3415 (N_3415,N_3275,N_3359);
nand U3416 (N_3416,N_3330,N_3270);
nor U3417 (N_3417,N_3252,N_3217);
and U3418 (N_3418,N_3250,N_3379);
nor U3419 (N_3419,N_3286,N_3309);
or U3420 (N_3420,N_3276,N_3263);
or U3421 (N_3421,N_3310,N_3385);
nand U3422 (N_3422,N_3381,N_3343);
and U3423 (N_3423,N_3341,N_3233);
or U3424 (N_3424,N_3215,N_3249);
nor U3425 (N_3425,N_3296,N_3329);
and U3426 (N_3426,N_3334,N_3390);
nor U3427 (N_3427,N_3287,N_3353);
or U3428 (N_3428,N_3387,N_3257);
nand U3429 (N_3429,N_3277,N_3312);
nand U3430 (N_3430,N_3308,N_3365);
nor U3431 (N_3431,N_3377,N_3280);
xnor U3432 (N_3432,N_3209,N_3243);
or U3433 (N_3433,N_3214,N_3327);
nand U3434 (N_3434,N_3348,N_3323);
or U3435 (N_3435,N_3304,N_3292);
or U3436 (N_3436,N_3301,N_3302);
nor U3437 (N_3437,N_3216,N_3360);
nand U3438 (N_3438,N_3333,N_3394);
and U3439 (N_3439,N_3279,N_3352);
or U3440 (N_3440,N_3241,N_3399);
or U3441 (N_3441,N_3319,N_3338);
and U3442 (N_3442,N_3383,N_3201);
nand U3443 (N_3443,N_3211,N_3342);
or U3444 (N_3444,N_3262,N_3363);
nand U3445 (N_3445,N_3378,N_3397);
or U3446 (N_3446,N_3210,N_3235);
or U3447 (N_3447,N_3265,N_3278);
and U3448 (N_3448,N_3290,N_3245);
and U3449 (N_3449,N_3373,N_3236);
nor U3450 (N_3450,N_3336,N_3355);
nand U3451 (N_3451,N_3326,N_3253);
nand U3452 (N_3452,N_3354,N_3204);
and U3453 (N_3453,N_3389,N_3247);
nor U3454 (N_3454,N_3256,N_3337);
nor U3455 (N_3455,N_3366,N_3282);
nand U3456 (N_3456,N_3324,N_3224);
nand U3457 (N_3457,N_3391,N_3221);
nand U3458 (N_3458,N_3315,N_3266);
nand U3459 (N_3459,N_3340,N_3294);
nor U3460 (N_3460,N_3322,N_3356);
or U3461 (N_3461,N_3313,N_3218);
or U3462 (N_3462,N_3254,N_3358);
or U3463 (N_3463,N_3212,N_3231);
or U3464 (N_3464,N_3200,N_3248);
nand U3465 (N_3465,N_3283,N_3369);
xor U3466 (N_3466,N_3344,N_3361);
nand U3467 (N_3467,N_3368,N_3321);
or U3468 (N_3468,N_3203,N_3392);
nand U3469 (N_3469,N_3345,N_3375);
or U3470 (N_3470,N_3384,N_3234);
or U3471 (N_3471,N_3305,N_3251);
nand U3472 (N_3472,N_3284,N_3298);
nor U3473 (N_3473,N_3259,N_3240);
and U3474 (N_3474,N_3223,N_3388);
and U3475 (N_3475,N_3380,N_3328);
and U3476 (N_3476,N_3281,N_3244);
and U3477 (N_3477,N_3261,N_3232);
and U3478 (N_3478,N_3371,N_3222);
nor U3479 (N_3479,N_3288,N_3303);
and U3480 (N_3480,N_3370,N_3386);
and U3481 (N_3481,N_3202,N_3260);
nor U3482 (N_3482,N_3382,N_3351);
and U3483 (N_3483,N_3332,N_3289);
and U3484 (N_3484,N_3307,N_3396);
nor U3485 (N_3485,N_3272,N_3206);
nor U3486 (N_3486,N_3357,N_3285);
nor U3487 (N_3487,N_3227,N_3267);
or U3488 (N_3488,N_3316,N_3225);
or U3489 (N_3489,N_3237,N_3317);
and U3490 (N_3490,N_3339,N_3372);
or U3491 (N_3491,N_3346,N_3367);
nor U3492 (N_3492,N_3229,N_3297);
or U3493 (N_3493,N_3311,N_3393);
and U3494 (N_3494,N_3205,N_3335);
nand U3495 (N_3495,N_3395,N_3219);
nand U3496 (N_3496,N_3325,N_3228);
nand U3497 (N_3497,N_3271,N_3268);
nor U3498 (N_3498,N_3398,N_3291);
nor U3499 (N_3499,N_3207,N_3230);
nor U3500 (N_3500,N_3296,N_3352);
nor U3501 (N_3501,N_3370,N_3351);
and U3502 (N_3502,N_3381,N_3248);
nor U3503 (N_3503,N_3341,N_3204);
nand U3504 (N_3504,N_3338,N_3300);
and U3505 (N_3505,N_3227,N_3259);
and U3506 (N_3506,N_3205,N_3310);
nor U3507 (N_3507,N_3341,N_3372);
or U3508 (N_3508,N_3364,N_3363);
or U3509 (N_3509,N_3203,N_3356);
or U3510 (N_3510,N_3279,N_3220);
or U3511 (N_3511,N_3314,N_3262);
and U3512 (N_3512,N_3259,N_3301);
nor U3513 (N_3513,N_3213,N_3389);
and U3514 (N_3514,N_3264,N_3224);
and U3515 (N_3515,N_3367,N_3339);
and U3516 (N_3516,N_3389,N_3302);
or U3517 (N_3517,N_3334,N_3351);
or U3518 (N_3518,N_3362,N_3393);
or U3519 (N_3519,N_3329,N_3280);
nand U3520 (N_3520,N_3261,N_3284);
nand U3521 (N_3521,N_3215,N_3325);
nand U3522 (N_3522,N_3304,N_3325);
nand U3523 (N_3523,N_3370,N_3279);
or U3524 (N_3524,N_3398,N_3321);
nand U3525 (N_3525,N_3315,N_3276);
nand U3526 (N_3526,N_3294,N_3371);
or U3527 (N_3527,N_3359,N_3240);
nand U3528 (N_3528,N_3217,N_3292);
and U3529 (N_3529,N_3221,N_3258);
xor U3530 (N_3530,N_3325,N_3376);
nor U3531 (N_3531,N_3347,N_3322);
or U3532 (N_3532,N_3334,N_3298);
and U3533 (N_3533,N_3301,N_3344);
and U3534 (N_3534,N_3282,N_3322);
or U3535 (N_3535,N_3365,N_3304);
and U3536 (N_3536,N_3285,N_3374);
nor U3537 (N_3537,N_3269,N_3201);
or U3538 (N_3538,N_3248,N_3341);
nor U3539 (N_3539,N_3308,N_3357);
or U3540 (N_3540,N_3201,N_3339);
and U3541 (N_3541,N_3271,N_3210);
nor U3542 (N_3542,N_3239,N_3279);
and U3543 (N_3543,N_3361,N_3286);
and U3544 (N_3544,N_3368,N_3338);
or U3545 (N_3545,N_3334,N_3226);
and U3546 (N_3546,N_3340,N_3391);
nand U3547 (N_3547,N_3390,N_3295);
or U3548 (N_3548,N_3308,N_3204);
nand U3549 (N_3549,N_3314,N_3211);
and U3550 (N_3550,N_3300,N_3330);
or U3551 (N_3551,N_3369,N_3250);
nor U3552 (N_3552,N_3225,N_3269);
or U3553 (N_3553,N_3275,N_3393);
and U3554 (N_3554,N_3396,N_3200);
and U3555 (N_3555,N_3349,N_3232);
nor U3556 (N_3556,N_3379,N_3268);
or U3557 (N_3557,N_3310,N_3334);
and U3558 (N_3558,N_3312,N_3390);
xnor U3559 (N_3559,N_3279,N_3309);
nand U3560 (N_3560,N_3339,N_3214);
and U3561 (N_3561,N_3334,N_3227);
nand U3562 (N_3562,N_3355,N_3207);
nand U3563 (N_3563,N_3257,N_3383);
or U3564 (N_3564,N_3217,N_3361);
or U3565 (N_3565,N_3344,N_3375);
nor U3566 (N_3566,N_3337,N_3324);
and U3567 (N_3567,N_3250,N_3224);
or U3568 (N_3568,N_3272,N_3280);
or U3569 (N_3569,N_3276,N_3256);
nand U3570 (N_3570,N_3285,N_3260);
or U3571 (N_3571,N_3323,N_3346);
nand U3572 (N_3572,N_3375,N_3301);
nand U3573 (N_3573,N_3272,N_3316);
or U3574 (N_3574,N_3233,N_3345);
or U3575 (N_3575,N_3260,N_3387);
nor U3576 (N_3576,N_3200,N_3226);
and U3577 (N_3577,N_3231,N_3249);
and U3578 (N_3578,N_3258,N_3220);
nand U3579 (N_3579,N_3345,N_3262);
and U3580 (N_3580,N_3226,N_3203);
or U3581 (N_3581,N_3276,N_3224);
or U3582 (N_3582,N_3320,N_3228);
nor U3583 (N_3583,N_3234,N_3293);
or U3584 (N_3584,N_3270,N_3309);
and U3585 (N_3585,N_3302,N_3294);
and U3586 (N_3586,N_3293,N_3252);
nand U3587 (N_3587,N_3222,N_3389);
and U3588 (N_3588,N_3285,N_3290);
nand U3589 (N_3589,N_3338,N_3253);
and U3590 (N_3590,N_3320,N_3202);
nor U3591 (N_3591,N_3364,N_3225);
and U3592 (N_3592,N_3250,N_3376);
or U3593 (N_3593,N_3231,N_3221);
or U3594 (N_3594,N_3303,N_3278);
and U3595 (N_3595,N_3352,N_3336);
nor U3596 (N_3596,N_3227,N_3207);
nand U3597 (N_3597,N_3389,N_3305);
nor U3598 (N_3598,N_3240,N_3341);
and U3599 (N_3599,N_3258,N_3262);
nand U3600 (N_3600,N_3457,N_3456);
nor U3601 (N_3601,N_3535,N_3500);
and U3602 (N_3602,N_3419,N_3403);
xnor U3603 (N_3603,N_3481,N_3566);
nand U3604 (N_3604,N_3517,N_3507);
or U3605 (N_3605,N_3436,N_3561);
nand U3606 (N_3606,N_3474,N_3422);
nor U3607 (N_3607,N_3478,N_3448);
nor U3608 (N_3608,N_3534,N_3524);
or U3609 (N_3609,N_3511,N_3529);
nand U3610 (N_3610,N_3551,N_3408);
or U3611 (N_3611,N_3485,N_3458);
nand U3612 (N_3612,N_3495,N_3514);
or U3613 (N_3613,N_3475,N_3538);
and U3614 (N_3614,N_3581,N_3586);
nand U3615 (N_3615,N_3413,N_3564);
nand U3616 (N_3616,N_3546,N_3560);
nor U3617 (N_3617,N_3497,N_3559);
or U3618 (N_3618,N_3579,N_3552);
nor U3619 (N_3619,N_3589,N_3400);
or U3620 (N_3620,N_3569,N_3558);
nor U3621 (N_3621,N_3466,N_3577);
or U3622 (N_3622,N_3482,N_3424);
xor U3623 (N_3623,N_3440,N_3426);
and U3624 (N_3624,N_3556,N_3463);
and U3625 (N_3625,N_3469,N_3404);
or U3626 (N_3626,N_3471,N_3575);
nand U3627 (N_3627,N_3541,N_3460);
nor U3628 (N_3628,N_3487,N_3416);
nor U3629 (N_3629,N_3493,N_3515);
or U3630 (N_3630,N_3486,N_3519);
nand U3631 (N_3631,N_3582,N_3498);
nand U3632 (N_3632,N_3578,N_3451);
nand U3633 (N_3633,N_3407,N_3585);
xor U3634 (N_3634,N_3472,N_3583);
nor U3635 (N_3635,N_3429,N_3414);
and U3636 (N_3636,N_3473,N_3438);
or U3637 (N_3637,N_3433,N_3480);
or U3638 (N_3638,N_3434,N_3593);
nand U3639 (N_3639,N_3431,N_3592);
nor U3640 (N_3640,N_3570,N_3542);
nor U3641 (N_3641,N_3402,N_3450);
and U3642 (N_3642,N_3439,N_3557);
nor U3643 (N_3643,N_3447,N_3454);
nor U3644 (N_3644,N_3553,N_3547);
nand U3645 (N_3645,N_3572,N_3533);
or U3646 (N_3646,N_3548,N_3568);
and U3647 (N_3647,N_3509,N_3405);
nand U3648 (N_3648,N_3415,N_3502);
and U3649 (N_3649,N_3468,N_3488);
nand U3650 (N_3650,N_3544,N_3432);
nor U3651 (N_3651,N_3573,N_3567);
nor U3652 (N_3652,N_3597,N_3499);
or U3653 (N_3653,N_3441,N_3508);
or U3654 (N_3654,N_3512,N_3503);
xnor U3655 (N_3655,N_3489,N_3521);
or U3656 (N_3656,N_3555,N_3598);
nand U3657 (N_3657,N_3562,N_3412);
or U3658 (N_3658,N_3494,N_3563);
nand U3659 (N_3659,N_3423,N_3516);
nor U3660 (N_3660,N_3513,N_3574);
or U3661 (N_3661,N_3470,N_3442);
nand U3662 (N_3662,N_3504,N_3554);
and U3663 (N_3663,N_3591,N_3540);
nand U3664 (N_3664,N_3490,N_3537);
nand U3665 (N_3665,N_3427,N_3417);
and U3666 (N_3666,N_3501,N_3444);
or U3667 (N_3667,N_3527,N_3421);
nor U3668 (N_3668,N_3459,N_3420);
nand U3669 (N_3669,N_3571,N_3506);
nand U3670 (N_3670,N_3435,N_3476);
nand U3671 (N_3671,N_3549,N_3599);
nand U3672 (N_3672,N_3443,N_3409);
nor U3673 (N_3673,N_3425,N_3526);
nor U3674 (N_3674,N_3532,N_3543);
or U3675 (N_3675,N_3455,N_3483);
nor U3676 (N_3676,N_3464,N_3580);
nand U3677 (N_3677,N_3406,N_3461);
nor U3678 (N_3678,N_3545,N_3445);
and U3679 (N_3679,N_3587,N_3411);
nand U3680 (N_3680,N_3530,N_3492);
or U3681 (N_3681,N_3452,N_3477);
nand U3682 (N_3682,N_3496,N_3479);
or U3683 (N_3683,N_3523,N_3437);
nor U3684 (N_3684,N_3428,N_3449);
or U3685 (N_3685,N_3510,N_3539);
and U3686 (N_3686,N_3531,N_3453);
nor U3687 (N_3687,N_3525,N_3484);
nand U3688 (N_3688,N_3410,N_3588);
and U3689 (N_3689,N_3595,N_3522);
nor U3690 (N_3690,N_3418,N_3565);
or U3691 (N_3691,N_3528,N_3584);
nand U3692 (N_3692,N_3401,N_3550);
nor U3693 (N_3693,N_3462,N_3590);
nor U3694 (N_3694,N_3446,N_3465);
nand U3695 (N_3695,N_3467,N_3520);
or U3696 (N_3696,N_3596,N_3518);
or U3697 (N_3697,N_3430,N_3505);
or U3698 (N_3698,N_3491,N_3536);
or U3699 (N_3699,N_3594,N_3576);
or U3700 (N_3700,N_3443,N_3504);
nor U3701 (N_3701,N_3516,N_3419);
and U3702 (N_3702,N_3532,N_3479);
or U3703 (N_3703,N_3459,N_3576);
and U3704 (N_3704,N_3506,N_3441);
and U3705 (N_3705,N_3506,N_3475);
nand U3706 (N_3706,N_3499,N_3404);
and U3707 (N_3707,N_3471,N_3428);
and U3708 (N_3708,N_3446,N_3421);
nand U3709 (N_3709,N_3488,N_3567);
or U3710 (N_3710,N_3404,N_3422);
or U3711 (N_3711,N_3567,N_3548);
and U3712 (N_3712,N_3439,N_3486);
xor U3713 (N_3713,N_3513,N_3514);
or U3714 (N_3714,N_3410,N_3415);
nor U3715 (N_3715,N_3591,N_3411);
nor U3716 (N_3716,N_3505,N_3501);
nor U3717 (N_3717,N_3563,N_3440);
nor U3718 (N_3718,N_3515,N_3565);
nor U3719 (N_3719,N_3412,N_3430);
nor U3720 (N_3720,N_3444,N_3545);
nand U3721 (N_3721,N_3532,N_3433);
and U3722 (N_3722,N_3414,N_3501);
and U3723 (N_3723,N_3441,N_3521);
or U3724 (N_3724,N_3547,N_3520);
or U3725 (N_3725,N_3522,N_3427);
or U3726 (N_3726,N_3577,N_3462);
or U3727 (N_3727,N_3442,N_3588);
nor U3728 (N_3728,N_3431,N_3476);
nor U3729 (N_3729,N_3410,N_3528);
and U3730 (N_3730,N_3422,N_3557);
and U3731 (N_3731,N_3419,N_3452);
or U3732 (N_3732,N_3509,N_3541);
or U3733 (N_3733,N_3414,N_3485);
or U3734 (N_3734,N_3503,N_3529);
and U3735 (N_3735,N_3520,N_3518);
or U3736 (N_3736,N_3463,N_3522);
and U3737 (N_3737,N_3459,N_3583);
nor U3738 (N_3738,N_3436,N_3421);
or U3739 (N_3739,N_3470,N_3417);
nand U3740 (N_3740,N_3555,N_3408);
and U3741 (N_3741,N_3499,N_3509);
or U3742 (N_3742,N_3420,N_3573);
nand U3743 (N_3743,N_3472,N_3591);
nor U3744 (N_3744,N_3480,N_3517);
nand U3745 (N_3745,N_3542,N_3407);
nand U3746 (N_3746,N_3433,N_3528);
nor U3747 (N_3747,N_3570,N_3476);
and U3748 (N_3748,N_3403,N_3524);
nor U3749 (N_3749,N_3516,N_3583);
and U3750 (N_3750,N_3563,N_3428);
and U3751 (N_3751,N_3447,N_3561);
nor U3752 (N_3752,N_3553,N_3417);
and U3753 (N_3753,N_3413,N_3594);
nand U3754 (N_3754,N_3508,N_3515);
and U3755 (N_3755,N_3502,N_3483);
nor U3756 (N_3756,N_3560,N_3586);
nor U3757 (N_3757,N_3539,N_3418);
and U3758 (N_3758,N_3470,N_3591);
nand U3759 (N_3759,N_3512,N_3437);
and U3760 (N_3760,N_3584,N_3555);
nor U3761 (N_3761,N_3414,N_3507);
or U3762 (N_3762,N_3465,N_3599);
or U3763 (N_3763,N_3579,N_3435);
and U3764 (N_3764,N_3572,N_3455);
and U3765 (N_3765,N_3520,N_3512);
nor U3766 (N_3766,N_3453,N_3522);
and U3767 (N_3767,N_3443,N_3487);
and U3768 (N_3768,N_3512,N_3491);
nand U3769 (N_3769,N_3489,N_3549);
or U3770 (N_3770,N_3594,N_3457);
nand U3771 (N_3771,N_3411,N_3463);
and U3772 (N_3772,N_3473,N_3510);
or U3773 (N_3773,N_3497,N_3572);
and U3774 (N_3774,N_3591,N_3560);
and U3775 (N_3775,N_3557,N_3509);
nand U3776 (N_3776,N_3575,N_3465);
nor U3777 (N_3777,N_3523,N_3557);
or U3778 (N_3778,N_3520,N_3510);
or U3779 (N_3779,N_3411,N_3505);
and U3780 (N_3780,N_3496,N_3591);
nand U3781 (N_3781,N_3592,N_3458);
nand U3782 (N_3782,N_3573,N_3593);
nor U3783 (N_3783,N_3592,N_3419);
or U3784 (N_3784,N_3584,N_3599);
nand U3785 (N_3785,N_3555,N_3469);
or U3786 (N_3786,N_3435,N_3487);
nand U3787 (N_3787,N_3497,N_3502);
nor U3788 (N_3788,N_3434,N_3568);
or U3789 (N_3789,N_3401,N_3492);
nand U3790 (N_3790,N_3512,N_3575);
or U3791 (N_3791,N_3513,N_3402);
and U3792 (N_3792,N_3575,N_3534);
nor U3793 (N_3793,N_3442,N_3465);
nor U3794 (N_3794,N_3519,N_3507);
or U3795 (N_3795,N_3433,N_3567);
nand U3796 (N_3796,N_3475,N_3544);
or U3797 (N_3797,N_3535,N_3408);
nand U3798 (N_3798,N_3513,N_3420);
nand U3799 (N_3799,N_3597,N_3522);
or U3800 (N_3800,N_3705,N_3648);
and U3801 (N_3801,N_3737,N_3745);
nand U3802 (N_3802,N_3791,N_3731);
nand U3803 (N_3803,N_3613,N_3688);
nor U3804 (N_3804,N_3796,N_3704);
nand U3805 (N_3805,N_3733,N_3607);
or U3806 (N_3806,N_3794,N_3681);
nand U3807 (N_3807,N_3717,N_3721);
nor U3808 (N_3808,N_3798,N_3734);
nand U3809 (N_3809,N_3647,N_3771);
nor U3810 (N_3810,N_3679,N_3610);
nand U3811 (N_3811,N_3746,N_3626);
nor U3812 (N_3812,N_3664,N_3697);
and U3813 (N_3813,N_3602,N_3718);
or U3814 (N_3814,N_3793,N_3789);
and U3815 (N_3815,N_3722,N_3735);
and U3816 (N_3816,N_3684,N_3689);
nand U3817 (N_3817,N_3636,N_3692);
and U3818 (N_3818,N_3642,N_3658);
nand U3819 (N_3819,N_3795,N_3677);
xnor U3820 (N_3820,N_3787,N_3779);
or U3821 (N_3821,N_3605,N_3749);
or U3822 (N_3822,N_3790,N_3674);
nor U3823 (N_3823,N_3799,N_3615);
nand U3824 (N_3824,N_3606,N_3661);
and U3825 (N_3825,N_3725,N_3616);
nor U3826 (N_3826,N_3634,N_3769);
nand U3827 (N_3827,N_3676,N_3707);
and U3828 (N_3828,N_3776,N_3719);
nor U3829 (N_3829,N_3627,N_3739);
or U3830 (N_3830,N_3780,N_3750);
nand U3831 (N_3831,N_3638,N_3713);
and U3832 (N_3832,N_3690,N_3736);
nand U3833 (N_3833,N_3762,N_3632);
and U3834 (N_3834,N_3673,N_3714);
nor U3835 (N_3835,N_3773,N_3728);
or U3836 (N_3836,N_3641,N_3631);
nor U3837 (N_3837,N_3645,N_3720);
nor U3838 (N_3838,N_3782,N_3743);
or U3839 (N_3839,N_3608,N_3604);
nor U3840 (N_3840,N_3633,N_3612);
and U3841 (N_3841,N_3700,N_3660);
nand U3842 (N_3842,N_3603,N_3662);
or U3843 (N_3843,N_3706,N_3772);
and U3844 (N_3844,N_3619,N_3715);
nor U3845 (N_3845,N_3748,N_3770);
and U3846 (N_3846,N_3781,N_3672);
nand U3847 (N_3847,N_3764,N_3614);
and U3848 (N_3848,N_3628,N_3695);
nor U3849 (N_3849,N_3797,N_3792);
nand U3850 (N_3850,N_3784,N_3687);
and U3851 (N_3851,N_3653,N_3759);
nor U3852 (N_3852,N_3708,N_3699);
nand U3853 (N_3853,N_3624,N_3761);
xnor U3854 (N_3854,N_3757,N_3785);
and U3855 (N_3855,N_3741,N_3670);
and U3856 (N_3856,N_3709,N_3742);
nand U3857 (N_3857,N_3702,N_3740);
nand U3858 (N_3858,N_3755,N_3665);
or U3859 (N_3859,N_3703,N_3635);
nor U3860 (N_3860,N_3685,N_3650);
nand U3861 (N_3861,N_3767,N_3629);
or U3862 (N_3862,N_3763,N_3783);
and U3863 (N_3863,N_3753,N_3617);
nand U3864 (N_3864,N_3710,N_3774);
and U3865 (N_3865,N_3694,N_3758);
nand U3866 (N_3866,N_3752,N_3659);
or U3867 (N_3867,N_3640,N_3651);
or U3868 (N_3868,N_3738,N_3751);
nand U3869 (N_3869,N_3671,N_3643);
nor U3870 (N_3870,N_3729,N_3678);
nand U3871 (N_3871,N_3726,N_3778);
and U3872 (N_3872,N_3744,N_3663);
or U3873 (N_3873,N_3657,N_3654);
or U3874 (N_3874,N_3655,N_3630);
and U3875 (N_3875,N_3682,N_3701);
xor U3876 (N_3876,N_3668,N_3646);
and U3877 (N_3877,N_3724,N_3727);
and U3878 (N_3878,N_3623,N_3712);
nand U3879 (N_3879,N_3622,N_3621);
nor U3880 (N_3880,N_3656,N_3768);
or U3881 (N_3881,N_3639,N_3667);
nand U3882 (N_3882,N_3680,N_3618);
or U3883 (N_3883,N_3716,N_3747);
nor U3884 (N_3884,N_3620,N_3696);
or U3885 (N_3885,N_3711,N_3649);
and U3886 (N_3886,N_3732,N_3601);
nand U3887 (N_3887,N_3637,N_3754);
and U3888 (N_3888,N_3600,N_3756);
or U3889 (N_3889,N_3723,N_3686);
or U3890 (N_3890,N_3786,N_3683);
and U3891 (N_3891,N_3652,N_3693);
nand U3892 (N_3892,N_3625,N_3609);
and U3893 (N_3893,N_3669,N_3777);
and U3894 (N_3894,N_3644,N_3788);
nand U3895 (N_3895,N_3760,N_3766);
nand U3896 (N_3896,N_3666,N_3611);
nand U3897 (N_3897,N_3698,N_3675);
nor U3898 (N_3898,N_3775,N_3730);
xnor U3899 (N_3899,N_3765,N_3691);
xnor U3900 (N_3900,N_3664,N_3676);
and U3901 (N_3901,N_3620,N_3610);
nor U3902 (N_3902,N_3680,N_3706);
and U3903 (N_3903,N_3722,N_3648);
or U3904 (N_3904,N_3791,N_3772);
nand U3905 (N_3905,N_3764,N_3762);
nor U3906 (N_3906,N_3753,N_3758);
and U3907 (N_3907,N_3746,N_3774);
or U3908 (N_3908,N_3757,N_3692);
nor U3909 (N_3909,N_3745,N_3721);
and U3910 (N_3910,N_3687,N_3619);
and U3911 (N_3911,N_3764,N_3752);
and U3912 (N_3912,N_3647,N_3697);
or U3913 (N_3913,N_3722,N_3631);
nor U3914 (N_3914,N_3686,N_3756);
nand U3915 (N_3915,N_3668,N_3717);
or U3916 (N_3916,N_3765,N_3752);
and U3917 (N_3917,N_3787,N_3641);
or U3918 (N_3918,N_3645,N_3687);
and U3919 (N_3919,N_3660,N_3782);
nand U3920 (N_3920,N_3702,N_3669);
and U3921 (N_3921,N_3643,N_3712);
or U3922 (N_3922,N_3764,N_3782);
or U3923 (N_3923,N_3639,N_3676);
and U3924 (N_3924,N_3799,N_3741);
and U3925 (N_3925,N_3672,N_3798);
and U3926 (N_3926,N_3773,N_3713);
nand U3927 (N_3927,N_3614,N_3715);
or U3928 (N_3928,N_3664,N_3603);
and U3929 (N_3929,N_3710,N_3631);
and U3930 (N_3930,N_3694,N_3646);
nand U3931 (N_3931,N_3739,N_3732);
nand U3932 (N_3932,N_3637,N_3751);
or U3933 (N_3933,N_3784,N_3679);
nor U3934 (N_3934,N_3753,N_3791);
nand U3935 (N_3935,N_3773,N_3790);
and U3936 (N_3936,N_3676,N_3666);
and U3937 (N_3937,N_3701,N_3745);
nor U3938 (N_3938,N_3720,N_3644);
and U3939 (N_3939,N_3707,N_3607);
and U3940 (N_3940,N_3749,N_3641);
nand U3941 (N_3941,N_3684,N_3742);
nor U3942 (N_3942,N_3728,N_3771);
and U3943 (N_3943,N_3727,N_3774);
nand U3944 (N_3944,N_3732,N_3695);
and U3945 (N_3945,N_3702,N_3786);
nand U3946 (N_3946,N_3710,N_3715);
or U3947 (N_3947,N_3759,N_3738);
and U3948 (N_3948,N_3669,N_3765);
nand U3949 (N_3949,N_3732,N_3706);
and U3950 (N_3950,N_3745,N_3757);
or U3951 (N_3951,N_3664,N_3600);
nor U3952 (N_3952,N_3622,N_3678);
or U3953 (N_3953,N_3799,N_3742);
or U3954 (N_3954,N_3645,N_3669);
nor U3955 (N_3955,N_3604,N_3704);
nor U3956 (N_3956,N_3759,N_3608);
nor U3957 (N_3957,N_3642,N_3616);
and U3958 (N_3958,N_3703,N_3792);
nor U3959 (N_3959,N_3688,N_3619);
and U3960 (N_3960,N_3614,N_3747);
and U3961 (N_3961,N_3604,N_3638);
and U3962 (N_3962,N_3650,N_3721);
nand U3963 (N_3963,N_3660,N_3711);
and U3964 (N_3964,N_3717,N_3732);
nand U3965 (N_3965,N_3779,N_3711);
nand U3966 (N_3966,N_3730,N_3624);
and U3967 (N_3967,N_3778,N_3771);
or U3968 (N_3968,N_3629,N_3717);
and U3969 (N_3969,N_3642,N_3676);
nor U3970 (N_3970,N_3795,N_3738);
or U3971 (N_3971,N_3711,N_3604);
and U3972 (N_3972,N_3671,N_3607);
nor U3973 (N_3973,N_3634,N_3649);
nand U3974 (N_3974,N_3719,N_3723);
nand U3975 (N_3975,N_3604,N_3706);
nand U3976 (N_3976,N_3671,N_3717);
and U3977 (N_3977,N_3645,N_3652);
nor U3978 (N_3978,N_3637,N_3629);
nand U3979 (N_3979,N_3665,N_3654);
nand U3980 (N_3980,N_3697,N_3773);
nor U3981 (N_3981,N_3633,N_3680);
nand U3982 (N_3982,N_3672,N_3716);
nor U3983 (N_3983,N_3620,N_3724);
nand U3984 (N_3984,N_3710,N_3600);
and U3985 (N_3985,N_3606,N_3656);
and U3986 (N_3986,N_3700,N_3633);
nand U3987 (N_3987,N_3763,N_3792);
nor U3988 (N_3988,N_3748,N_3619);
nor U3989 (N_3989,N_3615,N_3684);
or U3990 (N_3990,N_3734,N_3606);
nand U3991 (N_3991,N_3699,N_3646);
nand U3992 (N_3992,N_3642,N_3663);
and U3993 (N_3993,N_3604,N_3750);
nor U3994 (N_3994,N_3619,N_3637);
and U3995 (N_3995,N_3674,N_3779);
nand U3996 (N_3996,N_3712,N_3672);
nand U3997 (N_3997,N_3778,N_3627);
or U3998 (N_3998,N_3656,N_3761);
nor U3999 (N_3999,N_3729,N_3796);
or U4000 (N_4000,N_3876,N_3965);
xor U4001 (N_4001,N_3892,N_3810);
and U4002 (N_4002,N_3886,N_3845);
nor U4003 (N_4003,N_3922,N_3873);
or U4004 (N_4004,N_3879,N_3935);
and U4005 (N_4005,N_3909,N_3809);
nor U4006 (N_4006,N_3803,N_3833);
or U4007 (N_4007,N_3991,N_3866);
nor U4008 (N_4008,N_3881,N_3942);
and U4009 (N_4009,N_3952,N_3808);
and U4010 (N_4010,N_3917,N_3924);
and U4011 (N_4011,N_3934,N_3925);
or U4012 (N_4012,N_3901,N_3926);
nand U4013 (N_4013,N_3896,N_3825);
nand U4014 (N_4014,N_3945,N_3911);
or U4015 (N_4015,N_3899,N_3827);
and U4016 (N_4016,N_3969,N_3981);
or U4017 (N_4017,N_3861,N_3872);
or U4018 (N_4018,N_3943,N_3839);
or U4019 (N_4019,N_3995,N_3954);
nor U4020 (N_4020,N_3947,N_3992);
nor U4021 (N_4021,N_3936,N_3802);
nand U4022 (N_4022,N_3951,N_3842);
and U4023 (N_4023,N_3850,N_3915);
or U4024 (N_4024,N_3914,N_3955);
and U4025 (N_4025,N_3890,N_3804);
or U4026 (N_4026,N_3964,N_3865);
nand U4027 (N_4027,N_3843,N_3993);
nand U4028 (N_4028,N_3805,N_3877);
or U4029 (N_4029,N_3836,N_3972);
nor U4030 (N_4030,N_3921,N_3832);
nand U4031 (N_4031,N_3869,N_3916);
nor U4032 (N_4032,N_3834,N_3961);
or U4033 (N_4033,N_3870,N_3871);
nor U4034 (N_4034,N_3887,N_3801);
and U4035 (N_4035,N_3851,N_3800);
or U4036 (N_4036,N_3852,N_3996);
or U4037 (N_4037,N_3897,N_3889);
nor U4038 (N_4038,N_3908,N_3819);
nor U4039 (N_4039,N_3953,N_3944);
nand U4040 (N_4040,N_3874,N_3841);
and U4041 (N_4041,N_3878,N_3813);
nor U4042 (N_4042,N_3923,N_3855);
nor U4043 (N_4043,N_3975,N_3958);
or U4044 (N_4044,N_3971,N_3941);
nand U4045 (N_4045,N_3929,N_3902);
and U4046 (N_4046,N_3824,N_3977);
and U4047 (N_4047,N_3918,N_3905);
nand U4048 (N_4048,N_3847,N_3970);
and U4049 (N_4049,N_3898,N_3820);
nand U4050 (N_4050,N_3986,N_3864);
and U4051 (N_4051,N_3967,N_3831);
or U4052 (N_4052,N_3997,N_3867);
nor U4053 (N_4053,N_3907,N_3959);
or U4054 (N_4054,N_3999,N_3960);
nor U4055 (N_4055,N_3868,N_3933);
nor U4056 (N_4056,N_3837,N_3816);
and U4057 (N_4057,N_3856,N_3957);
or U4058 (N_4058,N_3859,N_3930);
or U4059 (N_4059,N_3882,N_3912);
nor U4060 (N_4060,N_3829,N_3956);
and U4061 (N_4061,N_3963,N_3811);
nand U4062 (N_4062,N_3913,N_3939);
or U4063 (N_4063,N_3822,N_3910);
and U4064 (N_4064,N_3826,N_3814);
nor U4065 (N_4065,N_3974,N_3883);
and U4066 (N_4066,N_3835,N_3906);
or U4067 (N_4067,N_3860,N_3968);
nand U4068 (N_4068,N_3976,N_3919);
nand U4069 (N_4069,N_3818,N_3880);
nor U4070 (N_4070,N_3940,N_3979);
and U4071 (N_4071,N_3982,N_3844);
and U4072 (N_4072,N_3985,N_3962);
or U4073 (N_4073,N_3848,N_3830);
nand U4074 (N_4074,N_3863,N_3904);
nand U4075 (N_4075,N_3990,N_3875);
nand U4076 (N_4076,N_3948,N_3987);
nand U4077 (N_4077,N_3900,N_3853);
and U4078 (N_4078,N_3821,N_3884);
nand U4079 (N_4079,N_3928,N_3949);
nand U4080 (N_4080,N_3849,N_3903);
nor U4081 (N_4081,N_3885,N_3857);
or U4082 (N_4082,N_3920,N_3938);
or U4083 (N_4083,N_3806,N_3854);
xnor U4084 (N_4084,N_3894,N_3978);
and U4085 (N_4085,N_3807,N_3812);
and U4086 (N_4086,N_3823,N_3846);
nand U4087 (N_4087,N_3891,N_3983);
nand U4088 (N_4088,N_3989,N_3840);
nor U4089 (N_4089,N_3988,N_3998);
and U4090 (N_4090,N_3862,N_3893);
nand U4091 (N_4091,N_3828,N_3927);
or U4092 (N_4092,N_3980,N_3888);
or U4093 (N_4093,N_3815,N_3966);
nor U4094 (N_4094,N_3932,N_3984);
nand U4095 (N_4095,N_3994,N_3931);
nand U4096 (N_4096,N_3838,N_3817);
nor U4097 (N_4097,N_3895,N_3946);
or U4098 (N_4098,N_3973,N_3950);
nand U4099 (N_4099,N_3858,N_3937);
nand U4100 (N_4100,N_3870,N_3834);
or U4101 (N_4101,N_3971,N_3934);
or U4102 (N_4102,N_3869,N_3874);
xnor U4103 (N_4103,N_3855,N_3987);
nor U4104 (N_4104,N_3919,N_3985);
nand U4105 (N_4105,N_3903,N_3803);
and U4106 (N_4106,N_3810,N_3943);
nand U4107 (N_4107,N_3932,N_3823);
and U4108 (N_4108,N_3985,N_3805);
and U4109 (N_4109,N_3840,N_3892);
and U4110 (N_4110,N_3890,N_3918);
nor U4111 (N_4111,N_3863,N_3934);
or U4112 (N_4112,N_3878,N_3883);
nand U4113 (N_4113,N_3953,N_3800);
and U4114 (N_4114,N_3848,N_3843);
or U4115 (N_4115,N_3932,N_3802);
nor U4116 (N_4116,N_3834,N_3958);
nor U4117 (N_4117,N_3850,N_3970);
nand U4118 (N_4118,N_3870,N_3986);
and U4119 (N_4119,N_3821,N_3829);
nand U4120 (N_4120,N_3910,N_3906);
and U4121 (N_4121,N_3923,N_3936);
nor U4122 (N_4122,N_3926,N_3968);
or U4123 (N_4123,N_3969,N_3968);
nand U4124 (N_4124,N_3967,N_3951);
nand U4125 (N_4125,N_3957,N_3980);
nor U4126 (N_4126,N_3805,N_3885);
nand U4127 (N_4127,N_3870,N_3897);
nand U4128 (N_4128,N_3884,N_3829);
nand U4129 (N_4129,N_3997,N_3955);
nor U4130 (N_4130,N_3865,N_3903);
nor U4131 (N_4131,N_3909,N_3923);
nor U4132 (N_4132,N_3913,N_3982);
nor U4133 (N_4133,N_3910,N_3844);
and U4134 (N_4134,N_3931,N_3948);
nand U4135 (N_4135,N_3801,N_3812);
nand U4136 (N_4136,N_3802,N_3874);
or U4137 (N_4137,N_3907,N_3942);
nor U4138 (N_4138,N_3846,N_3871);
and U4139 (N_4139,N_3956,N_3862);
and U4140 (N_4140,N_3838,N_3839);
or U4141 (N_4141,N_3986,N_3888);
xnor U4142 (N_4142,N_3842,N_3906);
nand U4143 (N_4143,N_3971,N_3868);
nand U4144 (N_4144,N_3965,N_3906);
or U4145 (N_4145,N_3869,N_3802);
and U4146 (N_4146,N_3985,N_3840);
nor U4147 (N_4147,N_3917,N_3886);
nor U4148 (N_4148,N_3982,N_3966);
or U4149 (N_4149,N_3829,N_3938);
and U4150 (N_4150,N_3857,N_3869);
nor U4151 (N_4151,N_3807,N_3945);
nor U4152 (N_4152,N_3964,N_3844);
and U4153 (N_4153,N_3833,N_3905);
nor U4154 (N_4154,N_3996,N_3817);
nor U4155 (N_4155,N_3924,N_3995);
and U4156 (N_4156,N_3921,N_3971);
nand U4157 (N_4157,N_3948,N_3968);
nand U4158 (N_4158,N_3867,N_3853);
nor U4159 (N_4159,N_3987,N_3818);
nor U4160 (N_4160,N_3804,N_3915);
or U4161 (N_4161,N_3871,N_3938);
or U4162 (N_4162,N_3862,N_3821);
or U4163 (N_4163,N_3958,N_3974);
nor U4164 (N_4164,N_3890,N_3885);
or U4165 (N_4165,N_3985,N_3865);
or U4166 (N_4166,N_3954,N_3920);
and U4167 (N_4167,N_3811,N_3808);
nand U4168 (N_4168,N_3973,N_3975);
xnor U4169 (N_4169,N_3913,N_3835);
nor U4170 (N_4170,N_3852,N_3952);
or U4171 (N_4171,N_3833,N_3964);
nand U4172 (N_4172,N_3966,N_3865);
and U4173 (N_4173,N_3868,N_3875);
nand U4174 (N_4174,N_3951,N_3830);
or U4175 (N_4175,N_3962,N_3864);
and U4176 (N_4176,N_3900,N_3985);
or U4177 (N_4177,N_3970,N_3961);
and U4178 (N_4178,N_3904,N_3829);
nor U4179 (N_4179,N_3863,N_3829);
nand U4180 (N_4180,N_3811,N_3947);
nor U4181 (N_4181,N_3986,N_3945);
nand U4182 (N_4182,N_3863,N_3989);
and U4183 (N_4183,N_3997,N_3909);
nand U4184 (N_4184,N_3836,N_3959);
nor U4185 (N_4185,N_3932,N_3967);
nor U4186 (N_4186,N_3968,N_3936);
nor U4187 (N_4187,N_3926,N_3990);
nor U4188 (N_4188,N_3890,N_3979);
or U4189 (N_4189,N_3889,N_3898);
nand U4190 (N_4190,N_3814,N_3853);
nand U4191 (N_4191,N_3945,N_3924);
xnor U4192 (N_4192,N_3823,N_3825);
nor U4193 (N_4193,N_3846,N_3955);
nor U4194 (N_4194,N_3867,N_3830);
nor U4195 (N_4195,N_3935,N_3868);
or U4196 (N_4196,N_3877,N_3888);
and U4197 (N_4197,N_3862,N_3878);
nor U4198 (N_4198,N_3990,N_3911);
nor U4199 (N_4199,N_3835,N_3936);
nor U4200 (N_4200,N_4176,N_4050);
nor U4201 (N_4201,N_4118,N_4123);
nor U4202 (N_4202,N_4020,N_4004);
nand U4203 (N_4203,N_4150,N_4141);
and U4204 (N_4204,N_4132,N_4171);
and U4205 (N_4205,N_4192,N_4175);
or U4206 (N_4206,N_4094,N_4145);
nor U4207 (N_4207,N_4166,N_4080);
nand U4208 (N_4208,N_4000,N_4098);
or U4209 (N_4209,N_4158,N_4074);
nor U4210 (N_4210,N_4173,N_4052);
nor U4211 (N_4211,N_4023,N_4042);
nand U4212 (N_4212,N_4193,N_4129);
nor U4213 (N_4213,N_4085,N_4009);
or U4214 (N_4214,N_4057,N_4165);
nor U4215 (N_4215,N_4177,N_4126);
and U4216 (N_4216,N_4078,N_4186);
or U4217 (N_4217,N_4063,N_4014);
nand U4218 (N_4218,N_4086,N_4021);
nand U4219 (N_4219,N_4089,N_4161);
nor U4220 (N_4220,N_4127,N_4025);
or U4221 (N_4221,N_4134,N_4071);
nor U4222 (N_4222,N_4148,N_4077);
or U4223 (N_4223,N_4054,N_4181);
nand U4224 (N_4224,N_4033,N_4082);
or U4225 (N_4225,N_4075,N_4007);
and U4226 (N_4226,N_4169,N_4001);
and U4227 (N_4227,N_4027,N_4048);
nand U4228 (N_4228,N_4065,N_4041);
nor U4229 (N_4229,N_4062,N_4051);
xor U4230 (N_4230,N_4101,N_4157);
nor U4231 (N_4231,N_4115,N_4011);
nand U4232 (N_4232,N_4045,N_4144);
xnor U4233 (N_4233,N_4090,N_4138);
or U4234 (N_4234,N_4196,N_4188);
nor U4235 (N_4235,N_4174,N_4106);
nand U4236 (N_4236,N_4010,N_4109);
and U4237 (N_4237,N_4055,N_4093);
or U4238 (N_4238,N_4122,N_4038);
nand U4239 (N_4239,N_4187,N_4066);
nand U4240 (N_4240,N_4018,N_4028);
xnor U4241 (N_4241,N_4029,N_4131);
nand U4242 (N_4242,N_4114,N_4003);
and U4243 (N_4243,N_4095,N_4111);
and U4244 (N_4244,N_4043,N_4079);
nor U4245 (N_4245,N_4163,N_4053);
and U4246 (N_4246,N_4191,N_4155);
or U4247 (N_4247,N_4160,N_4137);
and U4248 (N_4248,N_4184,N_4081);
and U4249 (N_4249,N_4046,N_4013);
and U4250 (N_4250,N_4006,N_4049);
xor U4251 (N_4251,N_4100,N_4092);
nor U4252 (N_4252,N_4142,N_4084);
nor U4253 (N_4253,N_4154,N_4149);
nor U4254 (N_4254,N_4199,N_4058);
and U4255 (N_4255,N_4147,N_4113);
or U4256 (N_4256,N_4087,N_4039);
nand U4257 (N_4257,N_4022,N_4030);
or U4258 (N_4258,N_4040,N_4197);
xor U4259 (N_4259,N_4107,N_4056);
nand U4260 (N_4260,N_4124,N_4152);
and U4261 (N_4261,N_4128,N_4036);
and U4262 (N_4262,N_4015,N_4099);
or U4263 (N_4263,N_4153,N_4120);
nand U4264 (N_4264,N_4088,N_4140);
and U4265 (N_4265,N_4143,N_4083);
nor U4266 (N_4266,N_4178,N_4139);
and U4267 (N_4267,N_4130,N_4104);
and U4268 (N_4268,N_4185,N_4002);
or U4269 (N_4269,N_4194,N_4195);
nand U4270 (N_4270,N_4156,N_4103);
and U4271 (N_4271,N_4164,N_4135);
and U4272 (N_4272,N_4168,N_4179);
nor U4273 (N_4273,N_4182,N_4097);
or U4274 (N_4274,N_4110,N_4016);
nand U4275 (N_4275,N_4067,N_4167);
or U4276 (N_4276,N_4112,N_4012);
nor U4277 (N_4277,N_4096,N_4072);
and U4278 (N_4278,N_4091,N_4190);
and U4279 (N_4279,N_4073,N_4136);
or U4280 (N_4280,N_4044,N_4170);
nor U4281 (N_4281,N_4076,N_4064);
nor U4282 (N_4282,N_4159,N_4105);
nand U4283 (N_4283,N_4108,N_4151);
nand U4284 (N_4284,N_4068,N_4017);
or U4285 (N_4285,N_4162,N_4172);
nor U4286 (N_4286,N_4180,N_4024);
nand U4287 (N_4287,N_4189,N_4069);
nor U4288 (N_4288,N_4102,N_4146);
and U4289 (N_4289,N_4035,N_4060);
nand U4290 (N_4290,N_4026,N_4183);
or U4291 (N_4291,N_4047,N_4005);
nand U4292 (N_4292,N_4133,N_4125);
or U4293 (N_4293,N_4119,N_4117);
or U4294 (N_4294,N_4034,N_4008);
nand U4295 (N_4295,N_4019,N_4059);
nand U4296 (N_4296,N_4032,N_4031);
and U4297 (N_4297,N_4121,N_4037);
nand U4298 (N_4298,N_4061,N_4198);
nand U4299 (N_4299,N_4116,N_4070);
or U4300 (N_4300,N_4143,N_4059);
or U4301 (N_4301,N_4097,N_4166);
and U4302 (N_4302,N_4017,N_4056);
nor U4303 (N_4303,N_4009,N_4153);
nor U4304 (N_4304,N_4085,N_4108);
nand U4305 (N_4305,N_4045,N_4036);
or U4306 (N_4306,N_4095,N_4155);
and U4307 (N_4307,N_4165,N_4047);
nor U4308 (N_4308,N_4000,N_4158);
and U4309 (N_4309,N_4031,N_4195);
or U4310 (N_4310,N_4174,N_4176);
nand U4311 (N_4311,N_4150,N_4065);
or U4312 (N_4312,N_4076,N_4169);
or U4313 (N_4313,N_4138,N_4092);
nand U4314 (N_4314,N_4145,N_4096);
nor U4315 (N_4315,N_4120,N_4137);
or U4316 (N_4316,N_4114,N_4198);
or U4317 (N_4317,N_4192,N_4080);
and U4318 (N_4318,N_4145,N_4105);
nand U4319 (N_4319,N_4058,N_4180);
nand U4320 (N_4320,N_4036,N_4088);
or U4321 (N_4321,N_4054,N_4164);
nor U4322 (N_4322,N_4152,N_4131);
nor U4323 (N_4323,N_4075,N_4170);
or U4324 (N_4324,N_4171,N_4033);
or U4325 (N_4325,N_4199,N_4105);
nor U4326 (N_4326,N_4082,N_4018);
nor U4327 (N_4327,N_4062,N_4019);
xnor U4328 (N_4328,N_4101,N_4137);
xor U4329 (N_4329,N_4121,N_4115);
and U4330 (N_4330,N_4137,N_4105);
nand U4331 (N_4331,N_4151,N_4021);
nor U4332 (N_4332,N_4021,N_4050);
and U4333 (N_4333,N_4106,N_4098);
or U4334 (N_4334,N_4059,N_4013);
and U4335 (N_4335,N_4102,N_4048);
nand U4336 (N_4336,N_4198,N_4105);
and U4337 (N_4337,N_4002,N_4000);
or U4338 (N_4338,N_4172,N_4093);
nor U4339 (N_4339,N_4005,N_4196);
and U4340 (N_4340,N_4123,N_4188);
nor U4341 (N_4341,N_4180,N_4044);
or U4342 (N_4342,N_4005,N_4088);
nor U4343 (N_4343,N_4044,N_4056);
or U4344 (N_4344,N_4068,N_4085);
or U4345 (N_4345,N_4120,N_4028);
or U4346 (N_4346,N_4048,N_4016);
nor U4347 (N_4347,N_4182,N_4112);
and U4348 (N_4348,N_4076,N_4044);
nand U4349 (N_4349,N_4103,N_4087);
or U4350 (N_4350,N_4079,N_4153);
nand U4351 (N_4351,N_4001,N_4071);
nor U4352 (N_4352,N_4099,N_4120);
or U4353 (N_4353,N_4061,N_4100);
nor U4354 (N_4354,N_4124,N_4100);
and U4355 (N_4355,N_4100,N_4073);
nor U4356 (N_4356,N_4085,N_4183);
nand U4357 (N_4357,N_4006,N_4046);
nand U4358 (N_4358,N_4132,N_4166);
nand U4359 (N_4359,N_4102,N_4014);
nand U4360 (N_4360,N_4034,N_4119);
and U4361 (N_4361,N_4022,N_4177);
nor U4362 (N_4362,N_4168,N_4081);
or U4363 (N_4363,N_4042,N_4001);
or U4364 (N_4364,N_4039,N_4024);
or U4365 (N_4365,N_4159,N_4015);
or U4366 (N_4366,N_4157,N_4142);
nor U4367 (N_4367,N_4023,N_4006);
and U4368 (N_4368,N_4194,N_4043);
or U4369 (N_4369,N_4179,N_4169);
or U4370 (N_4370,N_4042,N_4100);
nand U4371 (N_4371,N_4061,N_4125);
nand U4372 (N_4372,N_4130,N_4105);
or U4373 (N_4373,N_4184,N_4069);
or U4374 (N_4374,N_4132,N_4001);
and U4375 (N_4375,N_4119,N_4171);
nand U4376 (N_4376,N_4167,N_4096);
xor U4377 (N_4377,N_4149,N_4055);
and U4378 (N_4378,N_4144,N_4086);
nand U4379 (N_4379,N_4007,N_4133);
and U4380 (N_4380,N_4108,N_4115);
and U4381 (N_4381,N_4081,N_4037);
and U4382 (N_4382,N_4157,N_4130);
nor U4383 (N_4383,N_4094,N_4116);
nand U4384 (N_4384,N_4026,N_4129);
or U4385 (N_4385,N_4108,N_4011);
and U4386 (N_4386,N_4109,N_4113);
or U4387 (N_4387,N_4145,N_4098);
or U4388 (N_4388,N_4107,N_4006);
or U4389 (N_4389,N_4014,N_4057);
nand U4390 (N_4390,N_4181,N_4140);
nand U4391 (N_4391,N_4191,N_4067);
nor U4392 (N_4392,N_4124,N_4128);
and U4393 (N_4393,N_4147,N_4140);
or U4394 (N_4394,N_4139,N_4040);
nor U4395 (N_4395,N_4034,N_4189);
or U4396 (N_4396,N_4150,N_4184);
nand U4397 (N_4397,N_4034,N_4079);
nor U4398 (N_4398,N_4094,N_4118);
nand U4399 (N_4399,N_4035,N_4021);
nand U4400 (N_4400,N_4364,N_4331);
and U4401 (N_4401,N_4270,N_4300);
and U4402 (N_4402,N_4310,N_4268);
and U4403 (N_4403,N_4200,N_4255);
nand U4404 (N_4404,N_4336,N_4271);
or U4405 (N_4405,N_4269,N_4395);
nand U4406 (N_4406,N_4386,N_4347);
nand U4407 (N_4407,N_4321,N_4213);
and U4408 (N_4408,N_4334,N_4311);
xnor U4409 (N_4409,N_4263,N_4216);
nand U4410 (N_4410,N_4383,N_4391);
and U4411 (N_4411,N_4218,N_4252);
and U4412 (N_4412,N_4377,N_4384);
xnor U4413 (N_4413,N_4276,N_4204);
and U4414 (N_4414,N_4394,N_4344);
or U4415 (N_4415,N_4235,N_4380);
or U4416 (N_4416,N_4365,N_4289);
nand U4417 (N_4417,N_4370,N_4237);
nor U4418 (N_4418,N_4284,N_4322);
and U4419 (N_4419,N_4378,N_4264);
or U4420 (N_4420,N_4242,N_4317);
nand U4421 (N_4421,N_4371,N_4257);
nand U4422 (N_4422,N_4375,N_4222);
and U4423 (N_4423,N_4369,N_4228);
nand U4424 (N_4424,N_4313,N_4307);
nor U4425 (N_4425,N_4265,N_4214);
or U4426 (N_4426,N_4261,N_4248);
or U4427 (N_4427,N_4354,N_4387);
nand U4428 (N_4428,N_4324,N_4330);
nor U4429 (N_4429,N_4254,N_4298);
nor U4430 (N_4430,N_4390,N_4202);
nand U4431 (N_4431,N_4227,N_4294);
or U4432 (N_4432,N_4340,N_4337);
nand U4433 (N_4433,N_4362,N_4350);
nor U4434 (N_4434,N_4397,N_4296);
nor U4435 (N_4435,N_4238,N_4262);
and U4436 (N_4436,N_4389,N_4287);
nor U4437 (N_4437,N_4385,N_4291);
nor U4438 (N_4438,N_4224,N_4256);
and U4439 (N_4439,N_4244,N_4356);
nand U4440 (N_4440,N_4372,N_4320);
nand U4441 (N_4441,N_4209,N_4292);
and U4442 (N_4442,N_4220,N_4274);
nor U4443 (N_4443,N_4381,N_4273);
nor U4444 (N_4444,N_4328,N_4308);
or U4445 (N_4445,N_4203,N_4280);
nand U4446 (N_4446,N_4339,N_4286);
nor U4447 (N_4447,N_4205,N_4314);
nor U4448 (N_4448,N_4323,N_4223);
nor U4449 (N_4449,N_4379,N_4283);
nand U4450 (N_4450,N_4253,N_4278);
nand U4451 (N_4451,N_4388,N_4333);
nor U4452 (N_4452,N_4368,N_4246);
and U4453 (N_4453,N_4250,N_4366);
or U4454 (N_4454,N_4306,N_4319);
and U4455 (N_4455,N_4303,N_4293);
nand U4456 (N_4456,N_4382,N_4367);
and U4457 (N_4457,N_4239,N_4206);
and U4458 (N_4458,N_4399,N_4201);
or U4459 (N_4459,N_4297,N_4285);
nand U4460 (N_4460,N_4258,N_4376);
nand U4461 (N_4461,N_4290,N_4211);
nand U4462 (N_4462,N_4353,N_4355);
and U4463 (N_4463,N_4312,N_4327);
nand U4464 (N_4464,N_4358,N_4342);
nand U4465 (N_4465,N_4325,N_4245);
nor U4466 (N_4466,N_4338,N_4221);
or U4467 (N_4467,N_4281,N_4335);
or U4468 (N_4468,N_4233,N_4361);
and U4469 (N_4469,N_4215,N_4225);
nor U4470 (N_4470,N_4295,N_4341);
nor U4471 (N_4471,N_4247,N_4240);
nand U4472 (N_4472,N_4212,N_4234);
and U4473 (N_4473,N_4315,N_4230);
or U4474 (N_4474,N_4357,N_4267);
nor U4475 (N_4475,N_4329,N_4345);
and U4476 (N_4476,N_4302,N_4249);
nand U4477 (N_4477,N_4210,N_4351);
and U4478 (N_4478,N_4208,N_4266);
and U4479 (N_4479,N_4243,N_4251);
nand U4480 (N_4480,N_4241,N_4359);
nor U4481 (N_4481,N_4232,N_4318);
nand U4482 (N_4482,N_4374,N_4396);
nor U4483 (N_4483,N_4343,N_4217);
and U4484 (N_4484,N_4219,N_4299);
nor U4485 (N_4485,N_4277,N_4229);
nand U4486 (N_4486,N_4304,N_4260);
nand U4487 (N_4487,N_4316,N_4226);
or U4488 (N_4488,N_4236,N_4275);
nand U4489 (N_4489,N_4348,N_4231);
nand U4490 (N_4490,N_4393,N_4360);
or U4491 (N_4491,N_4301,N_4309);
nand U4492 (N_4492,N_4363,N_4349);
or U4493 (N_4493,N_4352,N_4207);
nand U4494 (N_4494,N_4392,N_4272);
nand U4495 (N_4495,N_4282,N_4279);
or U4496 (N_4496,N_4259,N_4346);
and U4497 (N_4497,N_4373,N_4398);
and U4498 (N_4498,N_4288,N_4326);
nand U4499 (N_4499,N_4305,N_4332);
nor U4500 (N_4500,N_4379,N_4276);
nand U4501 (N_4501,N_4335,N_4350);
xnor U4502 (N_4502,N_4306,N_4271);
and U4503 (N_4503,N_4387,N_4218);
nor U4504 (N_4504,N_4353,N_4282);
nand U4505 (N_4505,N_4213,N_4231);
nor U4506 (N_4506,N_4247,N_4292);
or U4507 (N_4507,N_4282,N_4267);
nand U4508 (N_4508,N_4241,N_4270);
or U4509 (N_4509,N_4394,N_4364);
nor U4510 (N_4510,N_4309,N_4206);
nor U4511 (N_4511,N_4326,N_4263);
nor U4512 (N_4512,N_4327,N_4209);
nand U4513 (N_4513,N_4254,N_4252);
or U4514 (N_4514,N_4390,N_4326);
nand U4515 (N_4515,N_4225,N_4231);
and U4516 (N_4516,N_4217,N_4385);
nand U4517 (N_4517,N_4324,N_4220);
and U4518 (N_4518,N_4370,N_4312);
nor U4519 (N_4519,N_4231,N_4268);
and U4520 (N_4520,N_4241,N_4224);
and U4521 (N_4521,N_4318,N_4308);
nor U4522 (N_4522,N_4239,N_4337);
and U4523 (N_4523,N_4296,N_4251);
nand U4524 (N_4524,N_4202,N_4382);
or U4525 (N_4525,N_4316,N_4222);
and U4526 (N_4526,N_4351,N_4208);
and U4527 (N_4527,N_4255,N_4386);
nand U4528 (N_4528,N_4252,N_4238);
or U4529 (N_4529,N_4345,N_4353);
and U4530 (N_4530,N_4263,N_4253);
nand U4531 (N_4531,N_4212,N_4241);
nor U4532 (N_4532,N_4237,N_4246);
nor U4533 (N_4533,N_4222,N_4207);
or U4534 (N_4534,N_4361,N_4376);
nor U4535 (N_4535,N_4270,N_4278);
nand U4536 (N_4536,N_4398,N_4342);
and U4537 (N_4537,N_4227,N_4248);
nor U4538 (N_4538,N_4243,N_4385);
nor U4539 (N_4539,N_4273,N_4217);
and U4540 (N_4540,N_4350,N_4265);
and U4541 (N_4541,N_4219,N_4213);
nor U4542 (N_4542,N_4276,N_4259);
nand U4543 (N_4543,N_4385,N_4209);
xnor U4544 (N_4544,N_4339,N_4399);
or U4545 (N_4545,N_4317,N_4343);
or U4546 (N_4546,N_4206,N_4258);
and U4547 (N_4547,N_4270,N_4248);
nand U4548 (N_4548,N_4310,N_4303);
nand U4549 (N_4549,N_4273,N_4223);
and U4550 (N_4550,N_4269,N_4357);
nor U4551 (N_4551,N_4324,N_4332);
or U4552 (N_4552,N_4275,N_4284);
or U4553 (N_4553,N_4275,N_4207);
or U4554 (N_4554,N_4273,N_4385);
nand U4555 (N_4555,N_4302,N_4317);
nand U4556 (N_4556,N_4337,N_4377);
and U4557 (N_4557,N_4384,N_4263);
and U4558 (N_4558,N_4340,N_4319);
or U4559 (N_4559,N_4258,N_4306);
nand U4560 (N_4560,N_4254,N_4292);
and U4561 (N_4561,N_4388,N_4342);
and U4562 (N_4562,N_4209,N_4359);
nand U4563 (N_4563,N_4256,N_4269);
or U4564 (N_4564,N_4381,N_4201);
nor U4565 (N_4565,N_4228,N_4233);
and U4566 (N_4566,N_4314,N_4369);
or U4567 (N_4567,N_4240,N_4336);
or U4568 (N_4568,N_4390,N_4334);
nor U4569 (N_4569,N_4202,N_4273);
or U4570 (N_4570,N_4314,N_4201);
or U4571 (N_4571,N_4219,N_4210);
or U4572 (N_4572,N_4366,N_4298);
nor U4573 (N_4573,N_4256,N_4218);
or U4574 (N_4574,N_4398,N_4213);
nor U4575 (N_4575,N_4246,N_4281);
or U4576 (N_4576,N_4283,N_4219);
nor U4577 (N_4577,N_4228,N_4342);
nand U4578 (N_4578,N_4297,N_4303);
nand U4579 (N_4579,N_4248,N_4273);
nand U4580 (N_4580,N_4331,N_4362);
nor U4581 (N_4581,N_4231,N_4249);
nand U4582 (N_4582,N_4387,N_4374);
nand U4583 (N_4583,N_4391,N_4264);
nand U4584 (N_4584,N_4290,N_4240);
nand U4585 (N_4585,N_4206,N_4333);
nor U4586 (N_4586,N_4354,N_4253);
or U4587 (N_4587,N_4290,N_4305);
and U4588 (N_4588,N_4216,N_4310);
and U4589 (N_4589,N_4314,N_4325);
nor U4590 (N_4590,N_4349,N_4315);
or U4591 (N_4591,N_4354,N_4372);
nor U4592 (N_4592,N_4353,N_4284);
nand U4593 (N_4593,N_4294,N_4394);
or U4594 (N_4594,N_4350,N_4242);
nor U4595 (N_4595,N_4230,N_4393);
and U4596 (N_4596,N_4352,N_4371);
nand U4597 (N_4597,N_4308,N_4310);
and U4598 (N_4598,N_4218,N_4335);
nor U4599 (N_4599,N_4269,N_4371);
nor U4600 (N_4600,N_4571,N_4575);
or U4601 (N_4601,N_4471,N_4449);
and U4602 (N_4602,N_4567,N_4443);
and U4603 (N_4603,N_4402,N_4572);
nor U4604 (N_4604,N_4502,N_4569);
or U4605 (N_4605,N_4577,N_4465);
nor U4606 (N_4606,N_4462,N_4562);
nand U4607 (N_4607,N_4512,N_4532);
nand U4608 (N_4608,N_4403,N_4422);
nand U4609 (N_4609,N_4404,N_4435);
nand U4610 (N_4610,N_4540,N_4506);
and U4611 (N_4611,N_4416,N_4491);
nand U4612 (N_4612,N_4494,N_4530);
nor U4613 (N_4613,N_4542,N_4480);
and U4614 (N_4614,N_4438,N_4584);
and U4615 (N_4615,N_4489,N_4406);
nor U4616 (N_4616,N_4568,N_4486);
nand U4617 (N_4617,N_4466,N_4588);
nand U4618 (N_4618,N_4495,N_4536);
or U4619 (N_4619,N_4440,N_4523);
nor U4620 (N_4620,N_4457,N_4436);
nand U4621 (N_4621,N_4556,N_4483);
nor U4622 (N_4622,N_4586,N_4549);
and U4623 (N_4623,N_4504,N_4488);
or U4624 (N_4624,N_4533,N_4413);
or U4625 (N_4625,N_4596,N_4551);
nand U4626 (N_4626,N_4529,N_4427);
and U4627 (N_4627,N_4447,N_4524);
and U4628 (N_4628,N_4554,N_4493);
or U4629 (N_4629,N_4446,N_4415);
nor U4630 (N_4630,N_4583,N_4552);
and U4631 (N_4631,N_4428,N_4579);
and U4632 (N_4632,N_4505,N_4570);
and U4633 (N_4633,N_4564,N_4520);
or U4634 (N_4634,N_4478,N_4459);
nor U4635 (N_4635,N_4418,N_4558);
and U4636 (N_4636,N_4414,N_4469);
nand U4637 (N_4637,N_4578,N_4590);
nor U4638 (N_4638,N_4409,N_4464);
and U4639 (N_4639,N_4425,N_4509);
and U4640 (N_4640,N_4525,N_4455);
and U4641 (N_4641,N_4454,N_4501);
or U4642 (N_4642,N_4595,N_4429);
or U4643 (N_4643,N_4482,N_4473);
and U4644 (N_4644,N_4432,N_4510);
or U4645 (N_4645,N_4574,N_4516);
nand U4646 (N_4646,N_4497,N_4582);
nand U4647 (N_4647,N_4592,N_4534);
xor U4648 (N_4648,N_4557,N_4405);
and U4649 (N_4649,N_4518,N_4531);
and U4650 (N_4650,N_4426,N_4500);
nor U4651 (N_4651,N_4423,N_4594);
nor U4652 (N_4652,N_4522,N_4492);
and U4653 (N_4653,N_4521,N_4580);
nor U4654 (N_4654,N_4546,N_4585);
and U4655 (N_4655,N_4400,N_4496);
nand U4656 (N_4656,N_4545,N_4484);
nor U4657 (N_4657,N_4442,N_4566);
and U4658 (N_4658,N_4470,N_4424);
and U4659 (N_4659,N_4412,N_4417);
nand U4660 (N_4660,N_4553,N_4448);
nand U4661 (N_4661,N_4503,N_4517);
nor U4662 (N_4662,N_4421,N_4410);
nor U4663 (N_4663,N_4481,N_4451);
nor U4664 (N_4664,N_4431,N_4419);
or U4665 (N_4665,N_4541,N_4548);
and U4666 (N_4666,N_4561,N_4441);
and U4667 (N_4667,N_4434,N_4444);
nor U4668 (N_4668,N_4499,N_4576);
nand U4669 (N_4669,N_4513,N_4445);
or U4670 (N_4670,N_4490,N_4463);
or U4671 (N_4671,N_4589,N_4535);
nand U4672 (N_4672,N_4526,N_4539);
nand U4673 (N_4673,N_4485,N_4597);
and U4674 (N_4674,N_4474,N_4507);
and U4675 (N_4675,N_4511,N_4476);
or U4676 (N_4676,N_4547,N_4461);
nand U4677 (N_4677,N_4528,N_4475);
nor U4678 (N_4678,N_4487,N_4420);
and U4679 (N_4679,N_4514,N_4565);
nor U4680 (N_4680,N_4555,N_4593);
nor U4681 (N_4681,N_4587,N_4439);
and U4682 (N_4682,N_4527,N_4401);
nor U4683 (N_4683,N_4538,N_4598);
or U4684 (N_4684,N_4453,N_4479);
nor U4685 (N_4685,N_4437,N_4559);
or U4686 (N_4686,N_4519,N_4543);
and U4687 (N_4687,N_4477,N_4460);
and U4688 (N_4688,N_4450,N_4498);
nor U4689 (N_4689,N_4515,N_4472);
nand U4690 (N_4690,N_4544,N_4411);
or U4691 (N_4691,N_4563,N_4456);
or U4692 (N_4692,N_4430,N_4573);
and U4693 (N_4693,N_4560,N_4407);
or U4694 (N_4694,N_4458,N_4537);
nor U4695 (N_4695,N_4599,N_4452);
and U4696 (N_4696,N_4581,N_4433);
or U4697 (N_4697,N_4550,N_4468);
nand U4698 (N_4698,N_4467,N_4591);
nand U4699 (N_4699,N_4408,N_4508);
or U4700 (N_4700,N_4593,N_4409);
nand U4701 (N_4701,N_4553,N_4497);
nand U4702 (N_4702,N_4486,N_4403);
and U4703 (N_4703,N_4475,N_4495);
or U4704 (N_4704,N_4473,N_4567);
and U4705 (N_4705,N_4403,N_4595);
and U4706 (N_4706,N_4574,N_4554);
or U4707 (N_4707,N_4579,N_4557);
nor U4708 (N_4708,N_4561,N_4544);
or U4709 (N_4709,N_4402,N_4477);
or U4710 (N_4710,N_4468,N_4406);
nor U4711 (N_4711,N_4441,N_4419);
and U4712 (N_4712,N_4525,N_4524);
nor U4713 (N_4713,N_4542,N_4493);
or U4714 (N_4714,N_4579,N_4418);
and U4715 (N_4715,N_4438,N_4441);
or U4716 (N_4716,N_4597,N_4405);
and U4717 (N_4717,N_4548,N_4510);
nor U4718 (N_4718,N_4506,N_4492);
nand U4719 (N_4719,N_4589,N_4416);
and U4720 (N_4720,N_4488,N_4575);
or U4721 (N_4721,N_4423,N_4587);
nand U4722 (N_4722,N_4476,N_4472);
nor U4723 (N_4723,N_4529,N_4538);
or U4724 (N_4724,N_4468,N_4590);
nor U4725 (N_4725,N_4530,N_4434);
or U4726 (N_4726,N_4591,N_4557);
nand U4727 (N_4727,N_4566,N_4525);
or U4728 (N_4728,N_4404,N_4453);
nor U4729 (N_4729,N_4463,N_4447);
nand U4730 (N_4730,N_4468,N_4570);
and U4731 (N_4731,N_4567,N_4426);
and U4732 (N_4732,N_4509,N_4415);
and U4733 (N_4733,N_4405,N_4473);
and U4734 (N_4734,N_4489,N_4593);
and U4735 (N_4735,N_4443,N_4468);
nand U4736 (N_4736,N_4582,N_4503);
and U4737 (N_4737,N_4533,N_4412);
and U4738 (N_4738,N_4482,N_4546);
nor U4739 (N_4739,N_4416,N_4585);
nand U4740 (N_4740,N_4489,N_4591);
and U4741 (N_4741,N_4565,N_4410);
and U4742 (N_4742,N_4527,N_4511);
or U4743 (N_4743,N_4527,N_4411);
or U4744 (N_4744,N_4584,N_4440);
or U4745 (N_4745,N_4568,N_4502);
or U4746 (N_4746,N_4494,N_4566);
or U4747 (N_4747,N_4424,N_4573);
nand U4748 (N_4748,N_4544,N_4577);
or U4749 (N_4749,N_4566,N_4449);
or U4750 (N_4750,N_4565,N_4541);
nor U4751 (N_4751,N_4431,N_4541);
or U4752 (N_4752,N_4452,N_4420);
nor U4753 (N_4753,N_4498,N_4415);
or U4754 (N_4754,N_4486,N_4561);
or U4755 (N_4755,N_4436,N_4425);
or U4756 (N_4756,N_4468,N_4551);
nor U4757 (N_4757,N_4516,N_4481);
nand U4758 (N_4758,N_4575,N_4433);
and U4759 (N_4759,N_4470,N_4504);
nor U4760 (N_4760,N_4473,N_4459);
nand U4761 (N_4761,N_4495,N_4532);
or U4762 (N_4762,N_4577,N_4471);
and U4763 (N_4763,N_4455,N_4519);
nor U4764 (N_4764,N_4544,N_4529);
or U4765 (N_4765,N_4474,N_4589);
and U4766 (N_4766,N_4575,N_4565);
or U4767 (N_4767,N_4541,N_4508);
nand U4768 (N_4768,N_4451,N_4596);
or U4769 (N_4769,N_4507,N_4544);
nand U4770 (N_4770,N_4544,N_4452);
nor U4771 (N_4771,N_4523,N_4422);
nor U4772 (N_4772,N_4400,N_4503);
and U4773 (N_4773,N_4506,N_4468);
and U4774 (N_4774,N_4495,N_4575);
nand U4775 (N_4775,N_4524,N_4552);
and U4776 (N_4776,N_4521,N_4512);
and U4777 (N_4777,N_4542,N_4536);
nor U4778 (N_4778,N_4441,N_4596);
nor U4779 (N_4779,N_4432,N_4557);
and U4780 (N_4780,N_4498,N_4497);
nand U4781 (N_4781,N_4501,N_4588);
or U4782 (N_4782,N_4479,N_4439);
and U4783 (N_4783,N_4536,N_4409);
and U4784 (N_4784,N_4579,N_4581);
nand U4785 (N_4785,N_4569,N_4556);
and U4786 (N_4786,N_4465,N_4409);
nand U4787 (N_4787,N_4568,N_4588);
nand U4788 (N_4788,N_4429,N_4400);
xor U4789 (N_4789,N_4546,N_4516);
or U4790 (N_4790,N_4422,N_4418);
and U4791 (N_4791,N_4411,N_4476);
nor U4792 (N_4792,N_4545,N_4438);
or U4793 (N_4793,N_4549,N_4444);
and U4794 (N_4794,N_4594,N_4533);
and U4795 (N_4795,N_4470,N_4560);
nor U4796 (N_4796,N_4460,N_4466);
or U4797 (N_4797,N_4488,N_4466);
nand U4798 (N_4798,N_4441,N_4521);
and U4799 (N_4799,N_4408,N_4588);
or U4800 (N_4800,N_4696,N_4769);
nor U4801 (N_4801,N_4600,N_4785);
nand U4802 (N_4802,N_4715,N_4615);
and U4803 (N_4803,N_4736,N_4705);
and U4804 (N_4804,N_4759,N_4761);
or U4805 (N_4805,N_4729,N_4716);
nor U4806 (N_4806,N_4687,N_4651);
or U4807 (N_4807,N_4668,N_4797);
xnor U4808 (N_4808,N_4799,N_4674);
or U4809 (N_4809,N_4607,N_4790);
or U4810 (N_4810,N_4760,N_4734);
or U4811 (N_4811,N_4731,N_4695);
nand U4812 (N_4812,N_4739,N_4634);
and U4813 (N_4813,N_4644,N_4743);
or U4814 (N_4814,N_4603,N_4633);
nand U4815 (N_4815,N_4707,N_4602);
nand U4816 (N_4816,N_4704,N_4624);
nand U4817 (N_4817,N_4654,N_4689);
nor U4818 (N_4818,N_4749,N_4718);
nor U4819 (N_4819,N_4642,N_4610);
nor U4820 (N_4820,N_4616,N_4669);
and U4821 (N_4821,N_4751,N_4636);
nand U4822 (N_4822,N_4673,N_4675);
nor U4823 (N_4823,N_4667,N_4775);
nor U4824 (N_4824,N_4764,N_4782);
and U4825 (N_4825,N_4640,N_4697);
nand U4826 (N_4826,N_4774,N_4781);
or U4827 (N_4827,N_4795,N_4720);
nor U4828 (N_4828,N_4740,N_4620);
or U4829 (N_4829,N_4737,N_4618);
nand U4830 (N_4830,N_4710,N_4784);
or U4831 (N_4831,N_4730,N_4728);
and U4832 (N_4832,N_4681,N_4738);
and U4833 (N_4833,N_4641,N_4701);
nand U4834 (N_4834,N_4676,N_4794);
or U4835 (N_4835,N_4745,N_4611);
or U4836 (N_4836,N_4711,N_4635);
and U4837 (N_4837,N_4639,N_4721);
and U4838 (N_4838,N_4645,N_4629);
or U4839 (N_4839,N_4765,N_4755);
nor U4840 (N_4840,N_4766,N_4780);
or U4841 (N_4841,N_4677,N_4714);
nor U4842 (N_4842,N_4778,N_4698);
or U4843 (N_4843,N_4692,N_4763);
nand U4844 (N_4844,N_4694,N_4750);
or U4845 (N_4845,N_4631,N_4757);
nor U4846 (N_4846,N_4670,N_4742);
nand U4847 (N_4847,N_4684,N_4638);
nand U4848 (N_4848,N_4617,N_4762);
or U4849 (N_4849,N_4657,N_4659);
xnor U4850 (N_4850,N_4726,N_4693);
and U4851 (N_4851,N_4612,N_4619);
nor U4852 (N_4852,N_4748,N_4604);
nor U4853 (N_4853,N_4756,N_4625);
and U4854 (N_4854,N_4699,N_4767);
nor U4855 (N_4855,N_4605,N_4777);
or U4856 (N_4856,N_4725,N_4702);
and U4857 (N_4857,N_4768,N_4746);
xor U4858 (N_4858,N_4723,N_4691);
nor U4859 (N_4859,N_4621,N_4666);
or U4860 (N_4860,N_4680,N_4626);
and U4861 (N_4861,N_4628,N_4792);
nor U4862 (N_4862,N_4796,N_4632);
nand U4863 (N_4863,N_4608,N_4647);
and U4864 (N_4864,N_4601,N_4708);
and U4865 (N_4865,N_4735,N_4671);
and U4866 (N_4866,N_4719,N_4706);
nor U4867 (N_4867,N_4685,N_4623);
nor U4868 (N_4868,N_4649,N_4788);
nand U4869 (N_4869,N_4773,N_4650);
nand U4870 (N_4870,N_4682,N_4653);
nand U4871 (N_4871,N_4664,N_4732);
and U4872 (N_4872,N_4643,N_4789);
and U4873 (N_4873,N_4747,N_4700);
nand U4874 (N_4874,N_4614,N_4663);
or U4875 (N_4875,N_4772,N_4793);
and U4876 (N_4876,N_4662,N_4672);
or U4877 (N_4877,N_4646,N_4786);
and U4878 (N_4878,N_4648,N_4713);
and U4879 (N_4879,N_4660,N_4679);
or U4880 (N_4880,N_4683,N_4758);
or U4881 (N_4881,N_4656,N_4630);
and U4882 (N_4882,N_4690,N_4703);
nand U4883 (N_4883,N_4724,N_4709);
or U4884 (N_4884,N_4661,N_4686);
or U4885 (N_4885,N_4658,N_4609);
nand U4886 (N_4886,N_4606,N_4783);
nor U4887 (N_4887,N_4752,N_4727);
and U4888 (N_4888,N_4688,N_4787);
nor U4889 (N_4889,N_4779,N_4712);
or U4890 (N_4890,N_4678,N_4741);
nor U4891 (N_4891,N_4776,N_4655);
and U4892 (N_4892,N_4613,N_4770);
nor U4893 (N_4893,N_4627,N_4753);
nand U4894 (N_4894,N_4665,N_4744);
and U4895 (N_4895,N_4722,N_4622);
nand U4896 (N_4896,N_4637,N_4733);
or U4897 (N_4897,N_4754,N_4652);
or U4898 (N_4898,N_4791,N_4798);
nand U4899 (N_4899,N_4771,N_4717);
and U4900 (N_4900,N_4650,N_4697);
nor U4901 (N_4901,N_4695,N_4772);
nand U4902 (N_4902,N_4753,N_4621);
nand U4903 (N_4903,N_4609,N_4601);
or U4904 (N_4904,N_4720,N_4662);
nand U4905 (N_4905,N_4660,N_4653);
and U4906 (N_4906,N_4699,N_4620);
or U4907 (N_4907,N_4722,N_4711);
or U4908 (N_4908,N_4762,N_4693);
or U4909 (N_4909,N_4728,N_4717);
or U4910 (N_4910,N_4729,N_4608);
and U4911 (N_4911,N_4793,N_4671);
and U4912 (N_4912,N_4712,N_4615);
or U4913 (N_4913,N_4673,N_4638);
nand U4914 (N_4914,N_4720,N_4676);
and U4915 (N_4915,N_4614,N_4683);
and U4916 (N_4916,N_4621,N_4710);
and U4917 (N_4917,N_4633,N_4668);
nand U4918 (N_4918,N_4787,N_4683);
nand U4919 (N_4919,N_4734,N_4788);
nand U4920 (N_4920,N_4758,N_4779);
nand U4921 (N_4921,N_4730,N_4645);
nand U4922 (N_4922,N_4775,N_4674);
and U4923 (N_4923,N_4632,N_4777);
nand U4924 (N_4924,N_4701,N_4715);
nand U4925 (N_4925,N_4659,N_4624);
nor U4926 (N_4926,N_4692,N_4735);
nand U4927 (N_4927,N_4754,N_4778);
and U4928 (N_4928,N_4709,N_4601);
and U4929 (N_4929,N_4740,N_4709);
or U4930 (N_4930,N_4656,N_4711);
and U4931 (N_4931,N_4726,N_4722);
or U4932 (N_4932,N_4706,N_4787);
and U4933 (N_4933,N_4604,N_4674);
nand U4934 (N_4934,N_4766,N_4679);
and U4935 (N_4935,N_4733,N_4773);
nand U4936 (N_4936,N_4612,N_4765);
nor U4937 (N_4937,N_4629,N_4718);
nand U4938 (N_4938,N_4607,N_4740);
or U4939 (N_4939,N_4765,N_4742);
and U4940 (N_4940,N_4747,N_4607);
nor U4941 (N_4941,N_4712,N_4601);
nor U4942 (N_4942,N_4798,N_4765);
nand U4943 (N_4943,N_4617,N_4770);
nor U4944 (N_4944,N_4641,N_4771);
or U4945 (N_4945,N_4659,N_4694);
nor U4946 (N_4946,N_4723,N_4638);
and U4947 (N_4947,N_4715,N_4671);
and U4948 (N_4948,N_4706,N_4649);
nor U4949 (N_4949,N_4796,N_4744);
xor U4950 (N_4950,N_4611,N_4642);
or U4951 (N_4951,N_4635,N_4764);
or U4952 (N_4952,N_4743,N_4712);
nand U4953 (N_4953,N_4709,N_4674);
nor U4954 (N_4954,N_4608,N_4798);
nor U4955 (N_4955,N_4676,N_4657);
and U4956 (N_4956,N_4704,N_4767);
and U4957 (N_4957,N_4648,N_4711);
or U4958 (N_4958,N_4737,N_4719);
nand U4959 (N_4959,N_4699,N_4659);
nand U4960 (N_4960,N_4659,N_4794);
and U4961 (N_4961,N_4703,N_4630);
nor U4962 (N_4962,N_4630,N_4610);
nor U4963 (N_4963,N_4726,N_4701);
nand U4964 (N_4964,N_4716,N_4702);
or U4965 (N_4965,N_4673,N_4608);
or U4966 (N_4966,N_4692,N_4647);
nor U4967 (N_4967,N_4767,N_4650);
or U4968 (N_4968,N_4742,N_4799);
nand U4969 (N_4969,N_4697,N_4707);
or U4970 (N_4970,N_4715,N_4748);
and U4971 (N_4971,N_4672,N_4737);
or U4972 (N_4972,N_4696,N_4684);
nand U4973 (N_4973,N_4703,N_4656);
and U4974 (N_4974,N_4639,N_4781);
and U4975 (N_4975,N_4706,N_4623);
nor U4976 (N_4976,N_4741,N_4783);
nand U4977 (N_4977,N_4758,N_4628);
nor U4978 (N_4978,N_4605,N_4697);
nor U4979 (N_4979,N_4649,N_4735);
and U4980 (N_4980,N_4681,N_4759);
nor U4981 (N_4981,N_4711,N_4684);
nand U4982 (N_4982,N_4749,N_4645);
and U4983 (N_4983,N_4785,N_4623);
and U4984 (N_4984,N_4724,N_4666);
nand U4985 (N_4985,N_4754,N_4706);
or U4986 (N_4986,N_4626,N_4782);
nor U4987 (N_4987,N_4778,N_4639);
nor U4988 (N_4988,N_4690,N_4665);
nor U4989 (N_4989,N_4667,N_4755);
nand U4990 (N_4990,N_4793,N_4694);
nor U4991 (N_4991,N_4605,N_4664);
or U4992 (N_4992,N_4660,N_4780);
nand U4993 (N_4993,N_4784,N_4783);
or U4994 (N_4994,N_4798,N_4737);
nand U4995 (N_4995,N_4706,N_4675);
nand U4996 (N_4996,N_4709,N_4671);
nand U4997 (N_4997,N_4630,N_4662);
and U4998 (N_4998,N_4656,N_4747);
and U4999 (N_4999,N_4669,N_4632);
and U5000 (N_5000,N_4849,N_4947);
and U5001 (N_5001,N_4960,N_4950);
nor U5002 (N_5002,N_4821,N_4842);
and U5003 (N_5003,N_4844,N_4990);
or U5004 (N_5004,N_4853,N_4926);
and U5005 (N_5005,N_4931,N_4877);
or U5006 (N_5006,N_4965,N_4891);
or U5007 (N_5007,N_4837,N_4971);
nor U5008 (N_5008,N_4973,N_4813);
and U5009 (N_5009,N_4864,N_4991);
nand U5010 (N_5010,N_4803,N_4952);
nor U5011 (N_5011,N_4957,N_4880);
and U5012 (N_5012,N_4805,N_4898);
and U5013 (N_5013,N_4881,N_4862);
and U5014 (N_5014,N_4863,N_4997);
nor U5015 (N_5015,N_4937,N_4944);
nor U5016 (N_5016,N_4954,N_4963);
and U5017 (N_5017,N_4988,N_4866);
nor U5018 (N_5018,N_4940,N_4928);
nor U5019 (N_5019,N_4999,N_4946);
nor U5020 (N_5020,N_4984,N_4834);
or U5021 (N_5021,N_4967,N_4911);
or U5022 (N_5022,N_4904,N_4979);
and U5023 (N_5023,N_4978,N_4943);
nor U5024 (N_5024,N_4976,N_4901);
nor U5025 (N_5025,N_4802,N_4932);
or U5026 (N_5026,N_4888,N_4817);
nor U5027 (N_5027,N_4884,N_4808);
nand U5028 (N_5028,N_4876,N_4839);
nor U5029 (N_5029,N_4989,N_4882);
or U5030 (N_5030,N_4879,N_4917);
and U5031 (N_5031,N_4861,N_4910);
nand U5032 (N_5032,N_4942,N_4833);
nand U5033 (N_5033,N_4987,N_4915);
and U5034 (N_5034,N_4945,N_4820);
nand U5035 (N_5035,N_4930,N_4852);
nand U5036 (N_5036,N_4860,N_4812);
or U5037 (N_5037,N_4993,N_4892);
and U5038 (N_5038,N_4994,N_4953);
nand U5039 (N_5039,N_4800,N_4832);
nor U5040 (N_5040,N_4948,N_4830);
nor U5041 (N_5041,N_4824,N_4806);
nand U5042 (N_5042,N_4835,N_4903);
and U5043 (N_5043,N_4956,N_4872);
and U5044 (N_5044,N_4935,N_4889);
or U5045 (N_5045,N_4894,N_4924);
xnor U5046 (N_5046,N_4909,N_4958);
or U5047 (N_5047,N_4907,N_4847);
or U5048 (N_5048,N_4809,N_4887);
or U5049 (N_5049,N_4814,N_4906);
or U5050 (N_5050,N_4949,N_4843);
and U5051 (N_5051,N_4941,N_4900);
nor U5052 (N_5052,N_4962,N_4826);
xnor U5053 (N_5053,N_4983,N_4846);
nor U5054 (N_5054,N_4896,N_4961);
nor U5055 (N_5055,N_4873,N_4905);
or U5056 (N_5056,N_4922,N_4977);
and U5057 (N_5057,N_4825,N_4831);
or U5058 (N_5058,N_4874,N_4854);
nor U5059 (N_5059,N_4850,N_4859);
and U5060 (N_5060,N_4810,N_4823);
nor U5061 (N_5061,N_4893,N_4841);
nand U5062 (N_5062,N_4939,N_4972);
or U5063 (N_5063,N_4938,N_4913);
nand U5064 (N_5064,N_4836,N_4918);
or U5065 (N_5065,N_4811,N_4920);
or U5066 (N_5066,N_4878,N_4919);
or U5067 (N_5067,N_4801,N_4966);
nand U5068 (N_5068,N_4916,N_4964);
nand U5069 (N_5069,N_4996,N_4921);
or U5070 (N_5070,N_4970,N_4927);
nor U5071 (N_5071,N_4815,N_4851);
or U5072 (N_5072,N_4968,N_4897);
nand U5073 (N_5073,N_4982,N_4867);
and U5074 (N_5074,N_4840,N_4980);
or U5075 (N_5075,N_4865,N_4858);
nor U5076 (N_5076,N_4827,N_4816);
nand U5077 (N_5077,N_4829,N_4828);
and U5078 (N_5078,N_4934,N_4848);
nand U5079 (N_5079,N_4998,N_4871);
nand U5080 (N_5080,N_4807,N_4929);
nor U5081 (N_5081,N_4899,N_4870);
and U5082 (N_5082,N_4895,N_4933);
and U5083 (N_5083,N_4908,N_4857);
nor U5084 (N_5084,N_4819,N_4822);
nor U5085 (N_5085,N_4986,N_4902);
or U5086 (N_5086,N_4875,N_4868);
and U5087 (N_5087,N_4818,N_4975);
and U5088 (N_5088,N_4804,N_4951);
nor U5089 (N_5089,N_4955,N_4838);
or U5090 (N_5090,N_4914,N_4885);
and U5091 (N_5091,N_4869,N_4959);
and U5092 (N_5092,N_4845,N_4890);
nand U5093 (N_5093,N_4974,N_4936);
and U5094 (N_5094,N_4925,N_4995);
xor U5095 (N_5095,N_4912,N_4856);
nor U5096 (N_5096,N_4969,N_4985);
nand U5097 (N_5097,N_4981,N_4855);
and U5098 (N_5098,N_4883,N_4923);
and U5099 (N_5099,N_4992,N_4886);
or U5100 (N_5100,N_4871,N_4831);
or U5101 (N_5101,N_4936,N_4988);
nand U5102 (N_5102,N_4832,N_4914);
and U5103 (N_5103,N_4854,N_4897);
nand U5104 (N_5104,N_4855,N_4907);
nor U5105 (N_5105,N_4895,N_4879);
nor U5106 (N_5106,N_4801,N_4809);
or U5107 (N_5107,N_4923,N_4838);
or U5108 (N_5108,N_4988,N_4874);
nand U5109 (N_5109,N_4835,N_4837);
nor U5110 (N_5110,N_4996,N_4955);
nor U5111 (N_5111,N_4987,N_4844);
or U5112 (N_5112,N_4998,N_4874);
nand U5113 (N_5113,N_4930,N_4846);
and U5114 (N_5114,N_4952,N_4939);
or U5115 (N_5115,N_4912,N_4818);
and U5116 (N_5116,N_4919,N_4910);
and U5117 (N_5117,N_4835,N_4984);
and U5118 (N_5118,N_4968,N_4818);
and U5119 (N_5119,N_4819,N_4904);
nand U5120 (N_5120,N_4910,N_4874);
and U5121 (N_5121,N_4995,N_4972);
and U5122 (N_5122,N_4945,N_4946);
or U5123 (N_5123,N_4895,N_4811);
nand U5124 (N_5124,N_4956,N_4858);
nor U5125 (N_5125,N_4807,N_4969);
nand U5126 (N_5126,N_4818,N_4955);
or U5127 (N_5127,N_4928,N_4836);
and U5128 (N_5128,N_4929,N_4951);
nand U5129 (N_5129,N_4942,N_4986);
or U5130 (N_5130,N_4806,N_4999);
and U5131 (N_5131,N_4883,N_4857);
nand U5132 (N_5132,N_4803,N_4898);
nand U5133 (N_5133,N_4829,N_4919);
nor U5134 (N_5134,N_4949,N_4985);
xor U5135 (N_5135,N_4899,N_4987);
nor U5136 (N_5136,N_4961,N_4804);
nor U5137 (N_5137,N_4804,N_4944);
and U5138 (N_5138,N_4841,N_4831);
or U5139 (N_5139,N_4905,N_4924);
nand U5140 (N_5140,N_4959,N_4809);
or U5141 (N_5141,N_4952,N_4978);
and U5142 (N_5142,N_4828,N_4970);
nor U5143 (N_5143,N_4839,N_4825);
or U5144 (N_5144,N_4997,N_4873);
nor U5145 (N_5145,N_4967,N_4910);
xor U5146 (N_5146,N_4976,N_4820);
nand U5147 (N_5147,N_4978,N_4896);
and U5148 (N_5148,N_4888,N_4956);
and U5149 (N_5149,N_4964,N_4967);
nand U5150 (N_5150,N_4936,N_4931);
or U5151 (N_5151,N_4944,N_4988);
and U5152 (N_5152,N_4932,N_4893);
or U5153 (N_5153,N_4869,N_4828);
or U5154 (N_5154,N_4833,N_4857);
and U5155 (N_5155,N_4890,N_4898);
nor U5156 (N_5156,N_4839,N_4999);
and U5157 (N_5157,N_4847,N_4916);
and U5158 (N_5158,N_4893,N_4970);
or U5159 (N_5159,N_4853,N_4948);
nand U5160 (N_5160,N_4946,N_4833);
and U5161 (N_5161,N_4814,N_4988);
nand U5162 (N_5162,N_4907,N_4974);
nand U5163 (N_5163,N_4990,N_4924);
nor U5164 (N_5164,N_4917,N_4899);
nor U5165 (N_5165,N_4961,N_4840);
xor U5166 (N_5166,N_4900,N_4882);
or U5167 (N_5167,N_4899,N_4869);
or U5168 (N_5168,N_4959,N_4977);
and U5169 (N_5169,N_4998,N_4824);
nor U5170 (N_5170,N_4873,N_4872);
or U5171 (N_5171,N_4943,N_4959);
nor U5172 (N_5172,N_4815,N_4958);
or U5173 (N_5173,N_4868,N_4986);
and U5174 (N_5174,N_4840,N_4903);
or U5175 (N_5175,N_4846,N_4965);
or U5176 (N_5176,N_4905,N_4995);
or U5177 (N_5177,N_4907,N_4931);
or U5178 (N_5178,N_4885,N_4979);
or U5179 (N_5179,N_4806,N_4988);
nand U5180 (N_5180,N_4872,N_4891);
nand U5181 (N_5181,N_4837,N_4915);
nor U5182 (N_5182,N_4930,N_4921);
nor U5183 (N_5183,N_4943,N_4866);
or U5184 (N_5184,N_4815,N_4952);
nor U5185 (N_5185,N_4916,N_4968);
and U5186 (N_5186,N_4905,N_4939);
nand U5187 (N_5187,N_4877,N_4814);
and U5188 (N_5188,N_4991,N_4885);
nand U5189 (N_5189,N_4956,N_4896);
nor U5190 (N_5190,N_4931,N_4887);
nand U5191 (N_5191,N_4983,N_4867);
and U5192 (N_5192,N_4853,N_4818);
and U5193 (N_5193,N_4874,N_4806);
or U5194 (N_5194,N_4952,N_4862);
nand U5195 (N_5195,N_4854,N_4917);
or U5196 (N_5196,N_4895,N_4860);
or U5197 (N_5197,N_4952,N_4990);
nor U5198 (N_5198,N_4835,N_4930);
nand U5199 (N_5199,N_4868,N_4883);
or U5200 (N_5200,N_5119,N_5154);
and U5201 (N_5201,N_5051,N_5055);
and U5202 (N_5202,N_5149,N_5019);
or U5203 (N_5203,N_5027,N_5124);
and U5204 (N_5204,N_5180,N_5071);
nor U5205 (N_5205,N_5063,N_5098);
and U5206 (N_5206,N_5128,N_5144);
and U5207 (N_5207,N_5042,N_5168);
and U5208 (N_5208,N_5061,N_5093);
nor U5209 (N_5209,N_5029,N_5038);
and U5210 (N_5210,N_5165,N_5131);
and U5211 (N_5211,N_5049,N_5178);
nand U5212 (N_5212,N_5028,N_5053);
or U5213 (N_5213,N_5037,N_5075);
or U5214 (N_5214,N_5187,N_5040);
nor U5215 (N_5215,N_5155,N_5169);
nand U5216 (N_5216,N_5020,N_5186);
and U5217 (N_5217,N_5068,N_5036);
nand U5218 (N_5218,N_5003,N_5190);
or U5219 (N_5219,N_5185,N_5088);
or U5220 (N_5220,N_5084,N_5145);
xnor U5221 (N_5221,N_5066,N_5010);
nand U5222 (N_5222,N_5160,N_5070);
or U5223 (N_5223,N_5085,N_5167);
nand U5224 (N_5224,N_5123,N_5058);
or U5225 (N_5225,N_5059,N_5089);
or U5226 (N_5226,N_5140,N_5114);
nor U5227 (N_5227,N_5033,N_5166);
or U5228 (N_5228,N_5146,N_5159);
nor U5229 (N_5229,N_5013,N_5151);
or U5230 (N_5230,N_5090,N_5017);
nand U5231 (N_5231,N_5138,N_5104);
nand U5232 (N_5232,N_5095,N_5176);
or U5233 (N_5233,N_5039,N_5106);
nand U5234 (N_5234,N_5122,N_5082);
and U5235 (N_5235,N_5035,N_5173);
nor U5236 (N_5236,N_5179,N_5044);
nor U5237 (N_5237,N_5094,N_5023);
or U5238 (N_5238,N_5134,N_5076);
nor U5239 (N_5239,N_5164,N_5143);
or U5240 (N_5240,N_5148,N_5195);
or U5241 (N_5241,N_5030,N_5047);
nor U5242 (N_5242,N_5198,N_5133);
or U5243 (N_5243,N_5183,N_5009);
and U5244 (N_5244,N_5118,N_5054);
or U5245 (N_5245,N_5005,N_5142);
nor U5246 (N_5246,N_5115,N_5056);
and U5247 (N_5247,N_5110,N_5153);
or U5248 (N_5248,N_5021,N_5116);
or U5249 (N_5249,N_5012,N_5163);
nand U5250 (N_5250,N_5136,N_5034);
nor U5251 (N_5251,N_5091,N_5080);
nand U5252 (N_5252,N_5126,N_5018);
nor U5253 (N_5253,N_5192,N_5135);
nand U5254 (N_5254,N_5177,N_5196);
nand U5255 (N_5255,N_5026,N_5015);
or U5256 (N_5256,N_5007,N_5087);
or U5257 (N_5257,N_5031,N_5107);
nand U5258 (N_5258,N_5162,N_5139);
and U5259 (N_5259,N_5150,N_5057);
nand U5260 (N_5260,N_5147,N_5022);
nand U5261 (N_5261,N_5172,N_5000);
nor U5262 (N_5262,N_5103,N_5156);
nor U5263 (N_5263,N_5092,N_5004);
and U5264 (N_5264,N_5043,N_5006);
nand U5265 (N_5265,N_5062,N_5045);
or U5266 (N_5266,N_5041,N_5060);
or U5267 (N_5267,N_5002,N_5109);
or U5268 (N_5268,N_5072,N_5079);
and U5269 (N_5269,N_5137,N_5102);
nor U5270 (N_5270,N_5032,N_5181);
nand U5271 (N_5271,N_5074,N_5008);
and U5272 (N_5272,N_5048,N_5184);
nand U5273 (N_5273,N_5129,N_5199);
or U5274 (N_5274,N_5193,N_5065);
nor U5275 (N_5275,N_5001,N_5161);
and U5276 (N_5276,N_5067,N_5120);
nand U5277 (N_5277,N_5069,N_5083);
and U5278 (N_5278,N_5157,N_5111);
nand U5279 (N_5279,N_5046,N_5050);
nor U5280 (N_5280,N_5108,N_5174);
nand U5281 (N_5281,N_5170,N_5152);
and U5282 (N_5282,N_5064,N_5141);
nor U5283 (N_5283,N_5171,N_5016);
nor U5284 (N_5284,N_5096,N_5086);
nand U5285 (N_5285,N_5125,N_5097);
and U5286 (N_5286,N_5189,N_5158);
or U5287 (N_5287,N_5052,N_5132);
or U5288 (N_5288,N_5100,N_5101);
and U5289 (N_5289,N_5077,N_5188);
or U5290 (N_5290,N_5117,N_5024);
or U5291 (N_5291,N_5025,N_5197);
or U5292 (N_5292,N_5099,N_5175);
nand U5293 (N_5293,N_5121,N_5081);
nand U5294 (N_5294,N_5078,N_5014);
nand U5295 (N_5295,N_5182,N_5191);
nand U5296 (N_5296,N_5194,N_5112);
nand U5297 (N_5297,N_5073,N_5011);
nor U5298 (N_5298,N_5127,N_5130);
or U5299 (N_5299,N_5113,N_5105);
or U5300 (N_5300,N_5146,N_5161);
nand U5301 (N_5301,N_5032,N_5107);
and U5302 (N_5302,N_5129,N_5193);
nor U5303 (N_5303,N_5194,N_5166);
nor U5304 (N_5304,N_5093,N_5154);
xor U5305 (N_5305,N_5007,N_5059);
or U5306 (N_5306,N_5195,N_5166);
nor U5307 (N_5307,N_5059,N_5111);
or U5308 (N_5308,N_5043,N_5000);
and U5309 (N_5309,N_5175,N_5027);
nor U5310 (N_5310,N_5178,N_5086);
nor U5311 (N_5311,N_5157,N_5174);
nor U5312 (N_5312,N_5084,N_5085);
nand U5313 (N_5313,N_5008,N_5093);
and U5314 (N_5314,N_5140,N_5195);
or U5315 (N_5315,N_5108,N_5091);
and U5316 (N_5316,N_5108,N_5100);
or U5317 (N_5317,N_5037,N_5172);
or U5318 (N_5318,N_5139,N_5135);
or U5319 (N_5319,N_5030,N_5043);
nand U5320 (N_5320,N_5039,N_5120);
nor U5321 (N_5321,N_5073,N_5177);
nor U5322 (N_5322,N_5042,N_5171);
and U5323 (N_5323,N_5021,N_5054);
or U5324 (N_5324,N_5022,N_5068);
and U5325 (N_5325,N_5149,N_5122);
nor U5326 (N_5326,N_5132,N_5135);
and U5327 (N_5327,N_5125,N_5012);
or U5328 (N_5328,N_5013,N_5145);
nor U5329 (N_5329,N_5106,N_5088);
and U5330 (N_5330,N_5133,N_5127);
nand U5331 (N_5331,N_5071,N_5081);
nand U5332 (N_5332,N_5013,N_5088);
nor U5333 (N_5333,N_5197,N_5031);
or U5334 (N_5334,N_5004,N_5039);
and U5335 (N_5335,N_5018,N_5144);
nand U5336 (N_5336,N_5191,N_5033);
nand U5337 (N_5337,N_5019,N_5165);
and U5338 (N_5338,N_5115,N_5108);
or U5339 (N_5339,N_5152,N_5026);
nor U5340 (N_5340,N_5191,N_5066);
nand U5341 (N_5341,N_5064,N_5110);
or U5342 (N_5342,N_5145,N_5001);
nor U5343 (N_5343,N_5020,N_5032);
or U5344 (N_5344,N_5032,N_5076);
nand U5345 (N_5345,N_5122,N_5086);
nand U5346 (N_5346,N_5043,N_5176);
nand U5347 (N_5347,N_5079,N_5143);
nand U5348 (N_5348,N_5146,N_5030);
and U5349 (N_5349,N_5025,N_5103);
nor U5350 (N_5350,N_5045,N_5057);
nand U5351 (N_5351,N_5030,N_5076);
and U5352 (N_5352,N_5074,N_5023);
nor U5353 (N_5353,N_5198,N_5077);
and U5354 (N_5354,N_5118,N_5199);
or U5355 (N_5355,N_5112,N_5114);
nand U5356 (N_5356,N_5080,N_5010);
nand U5357 (N_5357,N_5177,N_5022);
and U5358 (N_5358,N_5110,N_5156);
or U5359 (N_5359,N_5140,N_5013);
nand U5360 (N_5360,N_5064,N_5023);
or U5361 (N_5361,N_5035,N_5153);
and U5362 (N_5362,N_5013,N_5195);
and U5363 (N_5363,N_5177,N_5027);
or U5364 (N_5364,N_5008,N_5031);
and U5365 (N_5365,N_5080,N_5191);
nor U5366 (N_5366,N_5074,N_5174);
nand U5367 (N_5367,N_5146,N_5100);
nand U5368 (N_5368,N_5160,N_5018);
nand U5369 (N_5369,N_5037,N_5144);
and U5370 (N_5370,N_5159,N_5009);
nor U5371 (N_5371,N_5058,N_5018);
and U5372 (N_5372,N_5108,N_5004);
and U5373 (N_5373,N_5080,N_5106);
or U5374 (N_5374,N_5090,N_5064);
or U5375 (N_5375,N_5042,N_5021);
or U5376 (N_5376,N_5191,N_5058);
nand U5377 (N_5377,N_5188,N_5194);
nand U5378 (N_5378,N_5157,N_5029);
or U5379 (N_5379,N_5038,N_5176);
nor U5380 (N_5380,N_5173,N_5017);
nand U5381 (N_5381,N_5003,N_5097);
nor U5382 (N_5382,N_5023,N_5181);
or U5383 (N_5383,N_5036,N_5072);
or U5384 (N_5384,N_5000,N_5182);
nand U5385 (N_5385,N_5006,N_5121);
nor U5386 (N_5386,N_5022,N_5087);
nand U5387 (N_5387,N_5194,N_5146);
nand U5388 (N_5388,N_5193,N_5133);
nor U5389 (N_5389,N_5138,N_5175);
nor U5390 (N_5390,N_5118,N_5027);
or U5391 (N_5391,N_5148,N_5011);
nand U5392 (N_5392,N_5051,N_5158);
or U5393 (N_5393,N_5187,N_5137);
or U5394 (N_5394,N_5189,N_5063);
and U5395 (N_5395,N_5161,N_5059);
or U5396 (N_5396,N_5092,N_5185);
nand U5397 (N_5397,N_5034,N_5075);
and U5398 (N_5398,N_5174,N_5173);
nand U5399 (N_5399,N_5102,N_5121);
or U5400 (N_5400,N_5363,N_5200);
or U5401 (N_5401,N_5352,N_5260);
nand U5402 (N_5402,N_5388,N_5203);
and U5403 (N_5403,N_5245,N_5279);
xnor U5404 (N_5404,N_5362,N_5310);
nor U5405 (N_5405,N_5379,N_5269);
nor U5406 (N_5406,N_5394,N_5205);
nor U5407 (N_5407,N_5303,N_5300);
and U5408 (N_5408,N_5317,N_5386);
nor U5409 (N_5409,N_5393,N_5270);
nand U5410 (N_5410,N_5206,N_5396);
nor U5411 (N_5411,N_5373,N_5258);
or U5412 (N_5412,N_5228,N_5313);
and U5413 (N_5413,N_5225,N_5268);
or U5414 (N_5414,N_5332,N_5283);
nand U5415 (N_5415,N_5399,N_5368);
and U5416 (N_5416,N_5380,N_5309);
or U5417 (N_5417,N_5390,N_5219);
and U5418 (N_5418,N_5359,N_5339);
and U5419 (N_5419,N_5361,N_5285);
nor U5420 (N_5420,N_5244,N_5257);
and U5421 (N_5421,N_5289,N_5253);
and U5422 (N_5422,N_5273,N_5202);
nor U5423 (N_5423,N_5311,N_5249);
nand U5424 (N_5424,N_5385,N_5345);
or U5425 (N_5425,N_5357,N_5375);
and U5426 (N_5426,N_5207,N_5237);
or U5427 (N_5427,N_5217,N_5224);
or U5428 (N_5428,N_5328,N_5354);
nor U5429 (N_5429,N_5251,N_5227);
or U5430 (N_5430,N_5292,N_5241);
nor U5431 (N_5431,N_5376,N_5383);
or U5432 (N_5432,N_5341,N_5204);
and U5433 (N_5433,N_5274,N_5236);
nand U5434 (N_5434,N_5329,N_5323);
and U5435 (N_5435,N_5367,N_5264);
nor U5436 (N_5436,N_5247,N_5299);
and U5437 (N_5437,N_5389,N_5226);
nand U5438 (N_5438,N_5302,N_5278);
or U5439 (N_5439,N_5201,N_5209);
nand U5440 (N_5440,N_5377,N_5340);
nor U5441 (N_5441,N_5261,N_5333);
and U5442 (N_5442,N_5344,N_5398);
or U5443 (N_5443,N_5304,N_5334);
xnor U5444 (N_5444,N_5238,N_5240);
nor U5445 (N_5445,N_5369,N_5305);
nor U5446 (N_5446,N_5239,N_5277);
nor U5447 (N_5447,N_5231,N_5208);
and U5448 (N_5448,N_5378,N_5347);
or U5449 (N_5449,N_5322,N_5214);
nand U5450 (N_5450,N_5335,N_5229);
nor U5451 (N_5451,N_5348,N_5280);
nor U5452 (N_5452,N_5391,N_5256);
nand U5453 (N_5453,N_5321,N_5265);
nor U5454 (N_5454,N_5291,N_5315);
nand U5455 (N_5455,N_5326,N_5223);
or U5456 (N_5456,N_5282,N_5293);
nor U5457 (N_5457,N_5301,N_5222);
nor U5458 (N_5458,N_5212,N_5397);
and U5459 (N_5459,N_5370,N_5364);
or U5460 (N_5460,N_5215,N_5365);
nor U5461 (N_5461,N_5213,N_5342);
nand U5462 (N_5462,N_5330,N_5297);
or U5463 (N_5463,N_5248,N_5250);
nand U5464 (N_5464,N_5320,N_5308);
and U5465 (N_5465,N_5210,N_5294);
or U5466 (N_5466,N_5254,N_5392);
nor U5467 (N_5467,N_5360,N_5371);
nand U5468 (N_5468,N_5284,N_5349);
nand U5469 (N_5469,N_5287,N_5255);
nand U5470 (N_5470,N_5318,N_5276);
or U5471 (N_5471,N_5271,N_5382);
nor U5472 (N_5472,N_5366,N_5346);
nor U5473 (N_5473,N_5312,N_5350);
nand U5474 (N_5474,N_5314,N_5286);
nand U5475 (N_5475,N_5381,N_5331);
or U5476 (N_5476,N_5307,N_5211);
or U5477 (N_5477,N_5296,N_5235);
and U5478 (N_5478,N_5262,N_5384);
and U5479 (N_5479,N_5252,N_5246);
or U5480 (N_5480,N_5336,N_5387);
or U5481 (N_5481,N_5306,N_5267);
or U5482 (N_5482,N_5266,N_5232);
nand U5483 (N_5483,N_5243,N_5233);
nand U5484 (N_5484,N_5242,N_5338);
nand U5485 (N_5485,N_5216,N_5372);
nand U5486 (N_5486,N_5343,N_5358);
xnor U5487 (N_5487,N_5319,N_5272);
or U5488 (N_5488,N_5325,N_5374);
nand U5489 (N_5489,N_5327,N_5355);
or U5490 (N_5490,N_5351,N_5316);
nand U5491 (N_5491,N_5395,N_5220);
and U5492 (N_5492,N_5298,N_5324);
nor U5493 (N_5493,N_5353,N_5259);
nand U5494 (N_5494,N_5275,N_5337);
nor U5495 (N_5495,N_5281,N_5290);
and U5496 (N_5496,N_5218,N_5230);
nor U5497 (N_5497,N_5221,N_5234);
nand U5498 (N_5498,N_5295,N_5356);
and U5499 (N_5499,N_5263,N_5288);
nand U5500 (N_5500,N_5378,N_5286);
or U5501 (N_5501,N_5226,N_5398);
or U5502 (N_5502,N_5308,N_5249);
nand U5503 (N_5503,N_5234,N_5378);
and U5504 (N_5504,N_5297,N_5248);
nand U5505 (N_5505,N_5230,N_5217);
nand U5506 (N_5506,N_5300,N_5266);
nor U5507 (N_5507,N_5356,N_5270);
or U5508 (N_5508,N_5333,N_5207);
and U5509 (N_5509,N_5289,N_5250);
nand U5510 (N_5510,N_5219,N_5237);
and U5511 (N_5511,N_5388,N_5301);
nand U5512 (N_5512,N_5383,N_5333);
or U5513 (N_5513,N_5236,N_5336);
or U5514 (N_5514,N_5357,N_5252);
nor U5515 (N_5515,N_5398,N_5395);
or U5516 (N_5516,N_5215,N_5205);
or U5517 (N_5517,N_5358,N_5251);
nor U5518 (N_5518,N_5226,N_5296);
nand U5519 (N_5519,N_5345,N_5236);
or U5520 (N_5520,N_5317,N_5328);
nor U5521 (N_5521,N_5297,N_5359);
nand U5522 (N_5522,N_5218,N_5347);
nand U5523 (N_5523,N_5387,N_5287);
nor U5524 (N_5524,N_5323,N_5377);
and U5525 (N_5525,N_5238,N_5276);
nand U5526 (N_5526,N_5301,N_5201);
nand U5527 (N_5527,N_5282,N_5255);
nand U5528 (N_5528,N_5382,N_5246);
and U5529 (N_5529,N_5369,N_5365);
nor U5530 (N_5530,N_5209,N_5315);
and U5531 (N_5531,N_5211,N_5254);
nand U5532 (N_5532,N_5272,N_5366);
or U5533 (N_5533,N_5201,N_5259);
or U5534 (N_5534,N_5354,N_5379);
or U5535 (N_5535,N_5267,N_5213);
or U5536 (N_5536,N_5339,N_5329);
or U5537 (N_5537,N_5260,N_5292);
or U5538 (N_5538,N_5365,N_5278);
nor U5539 (N_5539,N_5310,N_5235);
or U5540 (N_5540,N_5371,N_5346);
nand U5541 (N_5541,N_5240,N_5250);
and U5542 (N_5542,N_5362,N_5259);
xor U5543 (N_5543,N_5312,N_5280);
and U5544 (N_5544,N_5351,N_5238);
and U5545 (N_5545,N_5312,N_5277);
and U5546 (N_5546,N_5301,N_5290);
or U5547 (N_5547,N_5399,N_5378);
nor U5548 (N_5548,N_5316,N_5308);
nand U5549 (N_5549,N_5284,N_5297);
and U5550 (N_5550,N_5380,N_5397);
xnor U5551 (N_5551,N_5273,N_5343);
nand U5552 (N_5552,N_5302,N_5252);
nor U5553 (N_5553,N_5395,N_5368);
and U5554 (N_5554,N_5254,N_5393);
or U5555 (N_5555,N_5354,N_5304);
or U5556 (N_5556,N_5219,N_5358);
nand U5557 (N_5557,N_5356,N_5301);
and U5558 (N_5558,N_5203,N_5319);
or U5559 (N_5559,N_5218,N_5224);
nor U5560 (N_5560,N_5248,N_5388);
nand U5561 (N_5561,N_5307,N_5201);
nand U5562 (N_5562,N_5260,N_5264);
and U5563 (N_5563,N_5241,N_5219);
and U5564 (N_5564,N_5378,N_5203);
nand U5565 (N_5565,N_5210,N_5268);
nand U5566 (N_5566,N_5237,N_5354);
or U5567 (N_5567,N_5237,N_5320);
nor U5568 (N_5568,N_5247,N_5203);
or U5569 (N_5569,N_5398,N_5356);
nand U5570 (N_5570,N_5338,N_5274);
nor U5571 (N_5571,N_5253,N_5287);
and U5572 (N_5572,N_5366,N_5218);
xor U5573 (N_5573,N_5289,N_5238);
nand U5574 (N_5574,N_5381,N_5201);
nor U5575 (N_5575,N_5360,N_5356);
nor U5576 (N_5576,N_5252,N_5315);
and U5577 (N_5577,N_5331,N_5221);
and U5578 (N_5578,N_5240,N_5214);
nor U5579 (N_5579,N_5331,N_5338);
nor U5580 (N_5580,N_5327,N_5241);
or U5581 (N_5581,N_5315,N_5284);
or U5582 (N_5582,N_5282,N_5259);
or U5583 (N_5583,N_5226,N_5315);
and U5584 (N_5584,N_5291,N_5391);
nor U5585 (N_5585,N_5200,N_5350);
nor U5586 (N_5586,N_5229,N_5270);
nand U5587 (N_5587,N_5254,N_5209);
nor U5588 (N_5588,N_5226,N_5266);
nor U5589 (N_5589,N_5357,N_5240);
and U5590 (N_5590,N_5378,N_5340);
nand U5591 (N_5591,N_5239,N_5238);
or U5592 (N_5592,N_5331,N_5372);
or U5593 (N_5593,N_5282,N_5274);
nor U5594 (N_5594,N_5397,N_5398);
or U5595 (N_5595,N_5286,N_5201);
and U5596 (N_5596,N_5333,N_5282);
and U5597 (N_5597,N_5309,N_5393);
and U5598 (N_5598,N_5316,N_5297);
nor U5599 (N_5599,N_5296,N_5350);
and U5600 (N_5600,N_5432,N_5441);
or U5601 (N_5601,N_5470,N_5578);
nor U5602 (N_5602,N_5559,N_5537);
or U5603 (N_5603,N_5574,N_5501);
and U5604 (N_5604,N_5450,N_5454);
or U5605 (N_5605,N_5442,N_5464);
and U5606 (N_5606,N_5410,N_5407);
nor U5607 (N_5607,N_5451,N_5494);
and U5608 (N_5608,N_5506,N_5547);
and U5609 (N_5609,N_5504,N_5415);
nand U5610 (N_5610,N_5418,N_5516);
and U5611 (N_5611,N_5596,N_5431);
and U5612 (N_5612,N_5480,N_5587);
or U5613 (N_5613,N_5561,N_5565);
or U5614 (N_5614,N_5406,N_5509);
nor U5615 (N_5615,N_5488,N_5562);
and U5616 (N_5616,N_5496,N_5593);
or U5617 (N_5617,N_5419,N_5489);
nand U5618 (N_5618,N_5542,N_5524);
nand U5619 (N_5619,N_5446,N_5497);
nor U5620 (N_5620,N_5540,N_5523);
nor U5621 (N_5621,N_5533,N_5571);
nand U5622 (N_5622,N_5430,N_5412);
nor U5623 (N_5623,N_5428,N_5427);
nor U5624 (N_5624,N_5589,N_5474);
or U5625 (N_5625,N_5577,N_5538);
or U5626 (N_5626,N_5583,N_5536);
nor U5627 (N_5627,N_5564,N_5576);
and U5628 (N_5628,N_5586,N_5567);
nand U5629 (N_5629,N_5502,N_5569);
nand U5630 (N_5630,N_5411,N_5566);
and U5631 (N_5631,N_5429,N_5552);
or U5632 (N_5632,N_5452,N_5459);
and U5633 (N_5633,N_5493,N_5532);
and U5634 (N_5634,N_5585,N_5515);
nor U5635 (N_5635,N_5591,N_5437);
nor U5636 (N_5636,N_5468,N_5505);
or U5637 (N_5637,N_5558,N_5528);
nand U5638 (N_5638,N_5570,N_5522);
nor U5639 (N_5639,N_5405,N_5541);
nor U5640 (N_5640,N_5453,N_5449);
and U5641 (N_5641,N_5414,N_5420);
nor U5642 (N_5642,N_5485,N_5482);
or U5643 (N_5643,N_5503,N_5525);
or U5644 (N_5644,N_5499,N_5460);
or U5645 (N_5645,N_5425,N_5582);
nand U5646 (N_5646,N_5416,N_5467);
nor U5647 (N_5647,N_5556,N_5413);
nand U5648 (N_5648,N_5487,N_5495);
nand U5649 (N_5649,N_5498,N_5531);
nor U5650 (N_5650,N_5465,N_5534);
nor U5651 (N_5651,N_5421,N_5557);
nand U5652 (N_5652,N_5403,N_5584);
nand U5653 (N_5653,N_5550,N_5546);
nor U5654 (N_5654,N_5491,N_5599);
and U5655 (N_5655,N_5549,N_5520);
nor U5656 (N_5656,N_5477,N_5422);
nand U5657 (N_5657,N_5445,N_5457);
xnor U5658 (N_5658,N_5580,N_5481);
nand U5659 (N_5659,N_5483,N_5492);
nand U5660 (N_5660,N_5568,N_5544);
and U5661 (N_5661,N_5440,N_5526);
nand U5662 (N_5662,N_5517,N_5554);
nor U5663 (N_5663,N_5519,N_5458);
or U5664 (N_5664,N_5535,N_5443);
nor U5665 (N_5665,N_5448,N_5592);
or U5666 (N_5666,N_5597,N_5484);
or U5667 (N_5667,N_5475,N_5435);
or U5668 (N_5668,N_5466,N_5560);
and U5669 (N_5669,N_5426,N_5438);
xor U5670 (N_5670,N_5408,N_5490);
nor U5671 (N_5671,N_5472,N_5476);
nor U5672 (N_5672,N_5402,N_5513);
or U5673 (N_5673,N_5409,N_5434);
nand U5674 (N_5674,N_5548,N_5588);
nand U5675 (N_5675,N_5563,N_5527);
nand U5676 (N_5676,N_5461,N_5581);
nand U5677 (N_5677,N_5572,N_5404);
and U5678 (N_5678,N_5551,N_5595);
nor U5679 (N_5679,N_5469,N_5479);
and U5680 (N_5680,N_5555,N_5553);
nor U5681 (N_5681,N_5401,N_5439);
or U5682 (N_5682,N_5436,N_5598);
nor U5683 (N_5683,N_5508,N_5514);
nor U5684 (N_5684,N_5590,N_5463);
and U5685 (N_5685,N_5573,N_5521);
or U5686 (N_5686,N_5471,N_5486);
nor U5687 (N_5687,N_5500,N_5507);
nor U5688 (N_5688,N_5529,N_5433);
nor U5689 (N_5689,N_5423,N_5400);
nor U5690 (N_5690,N_5473,N_5424);
or U5691 (N_5691,N_5575,N_5417);
or U5692 (N_5692,N_5478,N_5511);
nor U5693 (N_5693,N_5539,N_5594);
and U5694 (N_5694,N_5518,N_5447);
nor U5695 (N_5695,N_5510,N_5462);
or U5696 (N_5696,N_5455,N_5512);
and U5697 (N_5697,N_5545,N_5579);
or U5698 (N_5698,N_5543,N_5530);
and U5699 (N_5699,N_5456,N_5444);
or U5700 (N_5700,N_5408,N_5494);
or U5701 (N_5701,N_5426,N_5541);
and U5702 (N_5702,N_5556,N_5571);
nor U5703 (N_5703,N_5543,N_5506);
and U5704 (N_5704,N_5518,N_5466);
nor U5705 (N_5705,N_5524,N_5557);
nand U5706 (N_5706,N_5567,N_5491);
and U5707 (N_5707,N_5509,N_5540);
nor U5708 (N_5708,N_5564,N_5533);
nand U5709 (N_5709,N_5528,N_5428);
nand U5710 (N_5710,N_5462,N_5540);
or U5711 (N_5711,N_5462,N_5539);
and U5712 (N_5712,N_5416,N_5471);
xnor U5713 (N_5713,N_5510,N_5537);
and U5714 (N_5714,N_5549,N_5514);
or U5715 (N_5715,N_5472,N_5421);
and U5716 (N_5716,N_5425,N_5512);
nor U5717 (N_5717,N_5478,N_5572);
or U5718 (N_5718,N_5587,N_5426);
nor U5719 (N_5719,N_5480,N_5415);
nand U5720 (N_5720,N_5578,N_5593);
or U5721 (N_5721,N_5425,N_5530);
or U5722 (N_5722,N_5486,N_5488);
nor U5723 (N_5723,N_5593,N_5547);
nor U5724 (N_5724,N_5485,N_5467);
nand U5725 (N_5725,N_5488,N_5502);
nor U5726 (N_5726,N_5419,N_5589);
and U5727 (N_5727,N_5555,N_5548);
nand U5728 (N_5728,N_5535,N_5458);
and U5729 (N_5729,N_5585,N_5520);
or U5730 (N_5730,N_5418,N_5407);
nand U5731 (N_5731,N_5569,N_5563);
and U5732 (N_5732,N_5463,N_5415);
or U5733 (N_5733,N_5558,N_5547);
nor U5734 (N_5734,N_5542,N_5470);
xnor U5735 (N_5735,N_5443,N_5453);
nor U5736 (N_5736,N_5455,N_5441);
nand U5737 (N_5737,N_5430,N_5496);
and U5738 (N_5738,N_5552,N_5465);
and U5739 (N_5739,N_5413,N_5408);
or U5740 (N_5740,N_5465,N_5546);
and U5741 (N_5741,N_5450,N_5587);
nor U5742 (N_5742,N_5472,N_5595);
and U5743 (N_5743,N_5553,N_5566);
or U5744 (N_5744,N_5418,N_5467);
and U5745 (N_5745,N_5442,N_5403);
or U5746 (N_5746,N_5508,N_5419);
nor U5747 (N_5747,N_5515,N_5402);
nor U5748 (N_5748,N_5457,N_5494);
or U5749 (N_5749,N_5484,N_5401);
nor U5750 (N_5750,N_5435,N_5563);
xnor U5751 (N_5751,N_5429,N_5532);
or U5752 (N_5752,N_5408,N_5407);
nor U5753 (N_5753,N_5414,N_5574);
nand U5754 (N_5754,N_5493,N_5526);
and U5755 (N_5755,N_5426,N_5511);
or U5756 (N_5756,N_5471,N_5453);
or U5757 (N_5757,N_5465,N_5431);
and U5758 (N_5758,N_5410,N_5512);
nand U5759 (N_5759,N_5575,N_5519);
or U5760 (N_5760,N_5514,N_5478);
nand U5761 (N_5761,N_5451,N_5436);
and U5762 (N_5762,N_5402,N_5528);
or U5763 (N_5763,N_5504,N_5414);
and U5764 (N_5764,N_5510,N_5574);
nand U5765 (N_5765,N_5586,N_5482);
nor U5766 (N_5766,N_5523,N_5552);
nand U5767 (N_5767,N_5465,N_5556);
nor U5768 (N_5768,N_5484,N_5534);
nor U5769 (N_5769,N_5426,N_5545);
or U5770 (N_5770,N_5512,N_5524);
nor U5771 (N_5771,N_5561,N_5529);
nor U5772 (N_5772,N_5491,N_5470);
or U5773 (N_5773,N_5492,N_5478);
or U5774 (N_5774,N_5447,N_5474);
nand U5775 (N_5775,N_5401,N_5482);
or U5776 (N_5776,N_5410,N_5421);
and U5777 (N_5777,N_5517,N_5531);
nor U5778 (N_5778,N_5436,N_5575);
or U5779 (N_5779,N_5567,N_5568);
nor U5780 (N_5780,N_5538,N_5502);
or U5781 (N_5781,N_5534,N_5444);
and U5782 (N_5782,N_5515,N_5431);
nor U5783 (N_5783,N_5514,N_5453);
nand U5784 (N_5784,N_5404,N_5548);
or U5785 (N_5785,N_5413,N_5577);
or U5786 (N_5786,N_5412,N_5418);
nand U5787 (N_5787,N_5424,N_5456);
and U5788 (N_5788,N_5594,N_5509);
or U5789 (N_5789,N_5569,N_5495);
nor U5790 (N_5790,N_5574,N_5537);
nor U5791 (N_5791,N_5584,N_5577);
nor U5792 (N_5792,N_5559,N_5507);
or U5793 (N_5793,N_5515,N_5418);
nor U5794 (N_5794,N_5487,N_5578);
or U5795 (N_5795,N_5410,N_5531);
nand U5796 (N_5796,N_5488,N_5446);
and U5797 (N_5797,N_5497,N_5531);
xnor U5798 (N_5798,N_5529,N_5555);
or U5799 (N_5799,N_5550,N_5585);
or U5800 (N_5800,N_5770,N_5706);
and U5801 (N_5801,N_5724,N_5785);
nor U5802 (N_5802,N_5687,N_5666);
and U5803 (N_5803,N_5690,N_5793);
nor U5804 (N_5804,N_5644,N_5692);
nand U5805 (N_5805,N_5714,N_5619);
nor U5806 (N_5806,N_5601,N_5676);
or U5807 (N_5807,N_5621,N_5671);
nand U5808 (N_5808,N_5708,N_5775);
or U5809 (N_5809,N_5614,N_5615);
nand U5810 (N_5810,N_5688,N_5656);
and U5811 (N_5811,N_5766,N_5751);
and U5812 (N_5812,N_5716,N_5630);
and U5813 (N_5813,N_5790,N_5602);
and U5814 (N_5814,N_5788,N_5629);
or U5815 (N_5815,N_5632,N_5761);
nand U5816 (N_5816,N_5682,N_5709);
or U5817 (N_5817,N_5611,N_5739);
or U5818 (N_5818,N_5633,N_5718);
nor U5819 (N_5819,N_5720,N_5675);
nor U5820 (N_5820,N_5684,N_5731);
nor U5821 (N_5821,N_5789,N_5725);
or U5822 (N_5822,N_5685,N_5722);
or U5823 (N_5823,N_5740,N_5796);
or U5824 (N_5824,N_5700,N_5647);
and U5825 (N_5825,N_5744,N_5733);
or U5826 (N_5826,N_5752,N_5641);
nand U5827 (N_5827,N_5681,N_5723);
or U5828 (N_5828,N_5750,N_5730);
and U5829 (N_5829,N_5627,N_5701);
nor U5830 (N_5830,N_5653,N_5639);
nand U5831 (N_5831,N_5604,N_5669);
and U5832 (N_5832,N_5735,N_5677);
or U5833 (N_5833,N_5697,N_5661);
nand U5834 (N_5834,N_5623,N_5712);
or U5835 (N_5835,N_5655,N_5736);
nand U5836 (N_5836,N_5662,N_5749);
and U5837 (N_5837,N_5649,N_5717);
nand U5838 (N_5838,N_5603,N_5711);
nand U5839 (N_5839,N_5791,N_5672);
xnor U5840 (N_5840,N_5783,N_5693);
nand U5841 (N_5841,N_5651,N_5646);
and U5842 (N_5842,N_5797,N_5747);
and U5843 (N_5843,N_5691,N_5636);
nor U5844 (N_5844,N_5650,N_5705);
nor U5845 (N_5845,N_5732,N_5786);
and U5846 (N_5846,N_5781,N_5794);
nor U5847 (N_5847,N_5607,N_5780);
nand U5848 (N_5848,N_5704,N_5771);
nand U5849 (N_5849,N_5713,N_5745);
nor U5850 (N_5850,N_5686,N_5624);
and U5851 (N_5851,N_5738,N_5742);
nor U5852 (N_5852,N_5753,N_5799);
nand U5853 (N_5853,N_5652,N_5776);
nor U5854 (N_5854,N_5618,N_5683);
and U5855 (N_5855,N_5698,N_5715);
nor U5856 (N_5856,N_5674,N_5635);
or U5857 (N_5857,N_5778,N_5643);
or U5858 (N_5858,N_5757,N_5665);
and U5859 (N_5859,N_5729,N_5625);
and U5860 (N_5860,N_5631,N_5710);
or U5861 (N_5861,N_5702,N_5734);
nor U5862 (N_5862,N_5748,N_5784);
or U5863 (N_5863,N_5727,N_5654);
nand U5864 (N_5864,N_5737,N_5759);
or U5865 (N_5865,N_5764,N_5657);
and U5866 (N_5866,N_5772,N_5660);
or U5867 (N_5867,N_5689,N_5695);
nand U5868 (N_5868,N_5755,N_5741);
and U5869 (N_5869,N_5626,N_5699);
or U5870 (N_5870,N_5798,N_5608);
nor U5871 (N_5871,N_5617,N_5645);
and U5872 (N_5872,N_5721,N_5616);
nor U5873 (N_5873,N_5609,N_5606);
nor U5874 (N_5874,N_5795,N_5726);
or U5875 (N_5875,N_5613,N_5622);
nor U5876 (N_5876,N_5758,N_5782);
and U5877 (N_5877,N_5679,N_5670);
or U5878 (N_5878,N_5640,N_5762);
nor U5879 (N_5879,N_5746,N_5768);
nand U5880 (N_5880,N_5678,N_5694);
and U5881 (N_5881,N_5667,N_5696);
nand U5882 (N_5882,N_5792,N_5648);
and U5883 (N_5883,N_5773,N_5600);
and U5884 (N_5884,N_5663,N_5658);
or U5885 (N_5885,N_5634,N_5668);
nor U5886 (N_5886,N_5787,N_5763);
or U5887 (N_5887,N_5754,N_5777);
nand U5888 (N_5888,N_5659,N_5610);
nor U5889 (N_5889,N_5743,N_5680);
nor U5890 (N_5890,N_5760,N_5620);
and U5891 (N_5891,N_5605,N_5664);
or U5892 (N_5892,N_5756,N_5769);
nor U5893 (N_5893,N_5638,N_5719);
nand U5894 (N_5894,N_5765,N_5728);
nand U5895 (N_5895,N_5637,N_5612);
nor U5896 (N_5896,N_5779,N_5673);
or U5897 (N_5897,N_5774,N_5628);
or U5898 (N_5898,N_5642,N_5767);
or U5899 (N_5899,N_5707,N_5703);
and U5900 (N_5900,N_5726,N_5634);
and U5901 (N_5901,N_5669,N_5633);
nor U5902 (N_5902,N_5796,N_5625);
nand U5903 (N_5903,N_5707,N_5643);
nor U5904 (N_5904,N_5628,N_5797);
nor U5905 (N_5905,N_5773,N_5655);
or U5906 (N_5906,N_5644,N_5625);
or U5907 (N_5907,N_5638,N_5681);
or U5908 (N_5908,N_5723,N_5606);
nand U5909 (N_5909,N_5698,N_5758);
nand U5910 (N_5910,N_5687,N_5741);
and U5911 (N_5911,N_5637,N_5705);
or U5912 (N_5912,N_5772,N_5606);
and U5913 (N_5913,N_5680,N_5661);
nand U5914 (N_5914,N_5796,N_5654);
and U5915 (N_5915,N_5707,N_5768);
and U5916 (N_5916,N_5764,N_5707);
nand U5917 (N_5917,N_5673,N_5664);
nand U5918 (N_5918,N_5613,N_5742);
nand U5919 (N_5919,N_5681,N_5641);
and U5920 (N_5920,N_5715,N_5794);
and U5921 (N_5921,N_5769,N_5676);
nand U5922 (N_5922,N_5729,N_5754);
or U5923 (N_5923,N_5641,N_5753);
nor U5924 (N_5924,N_5793,N_5640);
nand U5925 (N_5925,N_5788,N_5796);
and U5926 (N_5926,N_5780,N_5738);
nor U5927 (N_5927,N_5650,N_5794);
and U5928 (N_5928,N_5675,N_5685);
or U5929 (N_5929,N_5705,N_5717);
and U5930 (N_5930,N_5796,N_5680);
nand U5931 (N_5931,N_5735,N_5733);
and U5932 (N_5932,N_5639,N_5702);
nor U5933 (N_5933,N_5679,N_5731);
or U5934 (N_5934,N_5760,N_5720);
or U5935 (N_5935,N_5630,N_5610);
or U5936 (N_5936,N_5682,N_5730);
and U5937 (N_5937,N_5632,N_5754);
nor U5938 (N_5938,N_5786,N_5789);
nand U5939 (N_5939,N_5774,N_5606);
and U5940 (N_5940,N_5670,N_5688);
nand U5941 (N_5941,N_5707,N_5778);
and U5942 (N_5942,N_5633,N_5757);
nor U5943 (N_5943,N_5707,N_5786);
nand U5944 (N_5944,N_5711,N_5781);
nor U5945 (N_5945,N_5653,N_5645);
or U5946 (N_5946,N_5686,N_5662);
and U5947 (N_5947,N_5624,N_5696);
or U5948 (N_5948,N_5771,N_5718);
and U5949 (N_5949,N_5764,N_5794);
or U5950 (N_5950,N_5719,N_5717);
or U5951 (N_5951,N_5661,N_5628);
and U5952 (N_5952,N_5775,N_5740);
nor U5953 (N_5953,N_5777,N_5763);
nand U5954 (N_5954,N_5794,N_5604);
nand U5955 (N_5955,N_5629,N_5659);
nand U5956 (N_5956,N_5679,N_5706);
nor U5957 (N_5957,N_5748,N_5678);
nand U5958 (N_5958,N_5783,N_5785);
xnor U5959 (N_5959,N_5659,N_5732);
nand U5960 (N_5960,N_5719,N_5641);
and U5961 (N_5961,N_5725,N_5704);
or U5962 (N_5962,N_5675,N_5628);
nand U5963 (N_5963,N_5707,N_5623);
and U5964 (N_5964,N_5646,N_5767);
nor U5965 (N_5965,N_5784,N_5749);
nor U5966 (N_5966,N_5719,N_5699);
and U5967 (N_5967,N_5685,N_5786);
nor U5968 (N_5968,N_5687,N_5682);
nand U5969 (N_5969,N_5638,N_5623);
nor U5970 (N_5970,N_5746,N_5721);
xor U5971 (N_5971,N_5637,N_5653);
nand U5972 (N_5972,N_5710,N_5675);
or U5973 (N_5973,N_5629,N_5631);
and U5974 (N_5974,N_5761,N_5777);
nor U5975 (N_5975,N_5603,N_5796);
or U5976 (N_5976,N_5725,N_5778);
or U5977 (N_5977,N_5616,N_5725);
and U5978 (N_5978,N_5611,N_5653);
or U5979 (N_5979,N_5725,N_5669);
or U5980 (N_5980,N_5603,N_5742);
or U5981 (N_5981,N_5798,N_5604);
nand U5982 (N_5982,N_5764,N_5634);
nand U5983 (N_5983,N_5729,N_5665);
or U5984 (N_5984,N_5704,N_5618);
or U5985 (N_5985,N_5621,N_5662);
nor U5986 (N_5986,N_5769,N_5718);
or U5987 (N_5987,N_5607,N_5669);
nor U5988 (N_5988,N_5710,N_5680);
and U5989 (N_5989,N_5652,N_5737);
or U5990 (N_5990,N_5663,N_5608);
xnor U5991 (N_5991,N_5778,N_5685);
nand U5992 (N_5992,N_5688,N_5605);
or U5993 (N_5993,N_5769,N_5695);
nand U5994 (N_5994,N_5669,N_5671);
nor U5995 (N_5995,N_5794,N_5790);
nor U5996 (N_5996,N_5714,N_5642);
xnor U5997 (N_5997,N_5709,N_5699);
nor U5998 (N_5998,N_5790,N_5762);
and U5999 (N_5999,N_5776,N_5644);
nor U6000 (N_6000,N_5926,N_5912);
or U6001 (N_6001,N_5931,N_5910);
and U6002 (N_6002,N_5981,N_5904);
nand U6003 (N_6003,N_5844,N_5923);
nand U6004 (N_6004,N_5979,N_5906);
nor U6005 (N_6005,N_5824,N_5955);
and U6006 (N_6006,N_5930,N_5922);
or U6007 (N_6007,N_5925,N_5803);
and U6008 (N_6008,N_5882,N_5816);
and U6009 (N_6009,N_5935,N_5916);
and U6010 (N_6010,N_5850,N_5986);
nand U6011 (N_6011,N_5948,N_5908);
nand U6012 (N_6012,N_5895,N_5875);
and U6013 (N_6013,N_5915,N_5947);
or U6014 (N_6014,N_5961,N_5903);
nor U6015 (N_6015,N_5939,N_5886);
or U6016 (N_6016,N_5911,N_5848);
nor U6017 (N_6017,N_5980,N_5888);
nor U6018 (N_6018,N_5813,N_5829);
and U6019 (N_6019,N_5814,N_5846);
nand U6020 (N_6020,N_5837,N_5817);
nor U6021 (N_6021,N_5952,N_5800);
or U6022 (N_6022,N_5989,N_5826);
nor U6023 (N_6023,N_5874,N_5967);
nand U6024 (N_6024,N_5857,N_5806);
and U6025 (N_6025,N_5996,N_5985);
and U6026 (N_6026,N_5841,N_5864);
nand U6027 (N_6027,N_5958,N_5894);
nand U6028 (N_6028,N_5984,N_5914);
or U6029 (N_6029,N_5987,N_5859);
nor U6030 (N_6030,N_5851,N_5838);
nand U6031 (N_6031,N_5810,N_5990);
nor U6032 (N_6032,N_5869,N_5972);
and U6033 (N_6033,N_5960,N_5913);
nand U6034 (N_6034,N_5811,N_5956);
nand U6035 (N_6035,N_5878,N_5891);
and U6036 (N_6036,N_5883,N_5924);
or U6037 (N_6037,N_5860,N_5971);
nor U6038 (N_6038,N_5821,N_5887);
nand U6039 (N_6039,N_5862,N_5885);
nor U6040 (N_6040,N_5893,N_5968);
nand U6041 (N_6041,N_5872,N_5983);
nor U6042 (N_6042,N_5991,N_5998);
nand U6043 (N_6043,N_5808,N_5941);
and U6044 (N_6044,N_5871,N_5856);
and U6045 (N_6045,N_5946,N_5907);
or U6046 (N_6046,N_5853,N_5852);
nor U6047 (N_6047,N_5819,N_5954);
nor U6048 (N_6048,N_5896,N_5937);
nand U6049 (N_6049,N_5865,N_5950);
nand U6050 (N_6050,N_5839,N_5970);
nor U6051 (N_6051,N_5957,N_5963);
or U6052 (N_6052,N_5976,N_5953);
nor U6053 (N_6053,N_5802,N_5828);
or U6054 (N_6054,N_5951,N_5959);
or U6055 (N_6055,N_5977,N_5909);
nand U6056 (N_6056,N_5933,N_5934);
and U6057 (N_6057,N_5866,N_5901);
nand U6058 (N_6058,N_5928,N_5884);
xor U6059 (N_6059,N_5900,N_5944);
nor U6060 (N_6060,N_5988,N_5807);
and U6061 (N_6061,N_5831,N_5876);
nand U6062 (N_6062,N_5858,N_5902);
nor U6063 (N_6063,N_5849,N_5809);
nor U6064 (N_6064,N_5804,N_5833);
or U6065 (N_6065,N_5973,N_5992);
nand U6066 (N_6066,N_5995,N_5982);
and U6067 (N_6067,N_5975,N_5917);
nor U6068 (N_6068,N_5881,N_5805);
nor U6069 (N_6069,N_5815,N_5993);
nand U6070 (N_6070,N_5836,N_5845);
and U6071 (N_6071,N_5892,N_5994);
nor U6072 (N_6072,N_5898,N_5870);
nor U6073 (N_6073,N_5855,N_5827);
nor U6074 (N_6074,N_5854,N_5920);
and U6075 (N_6075,N_5822,N_5940);
nor U6076 (N_6076,N_5823,N_5818);
and U6077 (N_6077,N_5966,N_5832);
nand U6078 (N_6078,N_5861,N_5835);
or U6079 (N_6079,N_5942,N_5879);
or U6080 (N_6080,N_5880,N_5927);
or U6081 (N_6081,N_5899,N_5868);
or U6082 (N_6082,N_5919,N_5936);
nor U6083 (N_6083,N_5938,N_5867);
and U6084 (N_6084,N_5801,N_5820);
nor U6085 (N_6085,N_5962,N_5949);
nor U6086 (N_6086,N_5999,N_5834);
or U6087 (N_6087,N_5877,N_5929);
and U6088 (N_6088,N_5873,N_5897);
nor U6089 (N_6089,N_5890,N_5812);
and U6090 (N_6090,N_5997,N_5830);
nand U6091 (N_6091,N_5932,N_5964);
or U6092 (N_6092,N_5918,N_5965);
or U6093 (N_6093,N_5889,N_5978);
nor U6094 (N_6094,N_5905,N_5842);
nand U6095 (N_6095,N_5847,N_5974);
or U6096 (N_6096,N_5863,N_5945);
or U6097 (N_6097,N_5969,N_5843);
nand U6098 (N_6098,N_5943,N_5921);
and U6099 (N_6099,N_5825,N_5840);
nand U6100 (N_6100,N_5981,N_5859);
or U6101 (N_6101,N_5879,N_5805);
nand U6102 (N_6102,N_5932,N_5904);
and U6103 (N_6103,N_5886,N_5931);
nand U6104 (N_6104,N_5817,N_5852);
xnor U6105 (N_6105,N_5947,N_5858);
or U6106 (N_6106,N_5830,N_5841);
and U6107 (N_6107,N_5940,N_5854);
and U6108 (N_6108,N_5858,N_5976);
and U6109 (N_6109,N_5959,N_5979);
nand U6110 (N_6110,N_5985,N_5907);
nor U6111 (N_6111,N_5885,N_5877);
nor U6112 (N_6112,N_5891,N_5818);
and U6113 (N_6113,N_5917,N_5949);
or U6114 (N_6114,N_5999,N_5846);
or U6115 (N_6115,N_5924,N_5918);
and U6116 (N_6116,N_5954,N_5826);
nor U6117 (N_6117,N_5927,N_5950);
or U6118 (N_6118,N_5882,N_5912);
or U6119 (N_6119,N_5929,N_5853);
or U6120 (N_6120,N_5965,N_5944);
and U6121 (N_6121,N_5936,N_5931);
and U6122 (N_6122,N_5912,N_5998);
or U6123 (N_6123,N_5959,N_5974);
and U6124 (N_6124,N_5888,N_5837);
nor U6125 (N_6125,N_5867,N_5970);
or U6126 (N_6126,N_5825,N_5991);
nor U6127 (N_6127,N_5901,N_5885);
nand U6128 (N_6128,N_5986,N_5815);
and U6129 (N_6129,N_5801,N_5802);
and U6130 (N_6130,N_5966,N_5928);
nand U6131 (N_6131,N_5852,N_5975);
nor U6132 (N_6132,N_5901,N_5876);
and U6133 (N_6133,N_5915,N_5931);
or U6134 (N_6134,N_5864,N_5916);
and U6135 (N_6135,N_5911,N_5830);
nand U6136 (N_6136,N_5823,N_5829);
nand U6137 (N_6137,N_5859,N_5871);
and U6138 (N_6138,N_5953,N_5966);
and U6139 (N_6139,N_5995,N_5885);
nand U6140 (N_6140,N_5990,N_5985);
nor U6141 (N_6141,N_5914,N_5994);
or U6142 (N_6142,N_5935,N_5973);
nand U6143 (N_6143,N_5803,N_5959);
nand U6144 (N_6144,N_5819,N_5940);
or U6145 (N_6145,N_5938,N_5926);
and U6146 (N_6146,N_5831,N_5870);
nor U6147 (N_6147,N_5982,N_5933);
and U6148 (N_6148,N_5968,N_5984);
xor U6149 (N_6149,N_5987,N_5825);
nand U6150 (N_6150,N_5819,N_5907);
nor U6151 (N_6151,N_5904,N_5919);
or U6152 (N_6152,N_5844,N_5912);
nor U6153 (N_6153,N_5944,N_5866);
or U6154 (N_6154,N_5861,N_5849);
nor U6155 (N_6155,N_5900,N_5954);
nand U6156 (N_6156,N_5965,N_5931);
nand U6157 (N_6157,N_5937,N_5998);
and U6158 (N_6158,N_5870,N_5856);
nor U6159 (N_6159,N_5900,N_5863);
nor U6160 (N_6160,N_5854,N_5909);
nand U6161 (N_6161,N_5945,N_5926);
nand U6162 (N_6162,N_5958,N_5930);
nor U6163 (N_6163,N_5986,N_5993);
or U6164 (N_6164,N_5805,N_5937);
or U6165 (N_6165,N_5860,N_5954);
nor U6166 (N_6166,N_5982,N_5969);
and U6167 (N_6167,N_5929,N_5919);
or U6168 (N_6168,N_5976,N_5812);
nor U6169 (N_6169,N_5947,N_5989);
or U6170 (N_6170,N_5825,N_5896);
nor U6171 (N_6171,N_5869,N_5837);
or U6172 (N_6172,N_5932,N_5855);
nand U6173 (N_6173,N_5918,N_5956);
nor U6174 (N_6174,N_5896,N_5949);
nand U6175 (N_6175,N_5982,N_5958);
nand U6176 (N_6176,N_5936,N_5820);
or U6177 (N_6177,N_5925,N_5961);
nand U6178 (N_6178,N_5857,N_5888);
or U6179 (N_6179,N_5992,N_5836);
or U6180 (N_6180,N_5874,N_5837);
or U6181 (N_6181,N_5951,N_5816);
nand U6182 (N_6182,N_5851,N_5813);
and U6183 (N_6183,N_5860,N_5839);
or U6184 (N_6184,N_5850,N_5949);
or U6185 (N_6185,N_5807,N_5819);
and U6186 (N_6186,N_5960,N_5833);
nor U6187 (N_6187,N_5923,N_5997);
and U6188 (N_6188,N_5863,N_5855);
nand U6189 (N_6189,N_5833,N_5863);
or U6190 (N_6190,N_5966,N_5977);
and U6191 (N_6191,N_5858,N_5837);
or U6192 (N_6192,N_5899,N_5856);
and U6193 (N_6193,N_5843,N_5850);
nor U6194 (N_6194,N_5908,N_5824);
nor U6195 (N_6195,N_5910,N_5882);
and U6196 (N_6196,N_5842,N_5889);
nor U6197 (N_6197,N_5807,N_5926);
or U6198 (N_6198,N_5968,N_5985);
nand U6199 (N_6199,N_5903,N_5997);
nor U6200 (N_6200,N_6142,N_6006);
nand U6201 (N_6201,N_6121,N_6149);
nor U6202 (N_6202,N_6032,N_6172);
nand U6203 (N_6203,N_6182,N_6129);
or U6204 (N_6204,N_6199,N_6165);
or U6205 (N_6205,N_6005,N_6166);
nand U6206 (N_6206,N_6088,N_6020);
nand U6207 (N_6207,N_6095,N_6078);
or U6208 (N_6208,N_6062,N_6146);
and U6209 (N_6209,N_6080,N_6039);
and U6210 (N_6210,N_6027,N_6023);
or U6211 (N_6211,N_6184,N_6136);
nand U6212 (N_6212,N_6175,N_6069);
nand U6213 (N_6213,N_6124,N_6128);
or U6214 (N_6214,N_6178,N_6097);
and U6215 (N_6215,N_6125,N_6192);
or U6216 (N_6216,N_6042,N_6179);
nand U6217 (N_6217,N_6108,N_6091);
or U6218 (N_6218,N_6057,N_6197);
or U6219 (N_6219,N_6180,N_6044);
xor U6220 (N_6220,N_6103,N_6058);
nor U6221 (N_6221,N_6153,N_6074);
and U6222 (N_6222,N_6026,N_6111);
and U6223 (N_6223,N_6002,N_6018);
or U6224 (N_6224,N_6119,N_6191);
nor U6225 (N_6225,N_6076,N_6082);
nor U6226 (N_6226,N_6061,N_6019);
nor U6227 (N_6227,N_6056,N_6167);
or U6228 (N_6228,N_6170,N_6070);
or U6229 (N_6229,N_6152,N_6003);
nand U6230 (N_6230,N_6089,N_6000);
nor U6231 (N_6231,N_6059,N_6038);
nand U6232 (N_6232,N_6017,N_6140);
nor U6233 (N_6233,N_6060,N_6157);
nor U6234 (N_6234,N_6106,N_6035);
nand U6235 (N_6235,N_6141,N_6110);
nand U6236 (N_6236,N_6160,N_6054);
nor U6237 (N_6237,N_6137,N_6164);
nand U6238 (N_6238,N_6147,N_6099);
and U6239 (N_6239,N_6093,N_6105);
or U6240 (N_6240,N_6040,N_6181);
nand U6241 (N_6241,N_6196,N_6168);
nand U6242 (N_6242,N_6010,N_6025);
or U6243 (N_6243,N_6092,N_6077);
or U6244 (N_6244,N_6009,N_6037);
and U6245 (N_6245,N_6118,N_6133);
or U6246 (N_6246,N_6013,N_6198);
or U6247 (N_6247,N_6190,N_6143);
nand U6248 (N_6248,N_6139,N_6194);
nand U6249 (N_6249,N_6043,N_6159);
nand U6250 (N_6250,N_6134,N_6015);
and U6251 (N_6251,N_6156,N_6073);
nand U6252 (N_6252,N_6081,N_6011);
or U6253 (N_6253,N_6008,N_6031);
and U6254 (N_6254,N_6130,N_6055);
nor U6255 (N_6255,N_6132,N_6041);
nor U6256 (N_6256,N_6183,N_6187);
and U6257 (N_6257,N_6100,N_6066);
nor U6258 (N_6258,N_6096,N_6001);
nand U6259 (N_6259,N_6126,N_6085);
nand U6260 (N_6260,N_6155,N_6195);
and U6261 (N_6261,N_6030,N_6045);
nor U6262 (N_6262,N_6113,N_6075);
nand U6263 (N_6263,N_6016,N_6104);
nand U6264 (N_6264,N_6163,N_6115);
nand U6265 (N_6265,N_6186,N_6083);
xnor U6266 (N_6266,N_6049,N_6135);
nor U6267 (N_6267,N_6185,N_6050);
or U6268 (N_6268,N_6176,N_6193);
or U6269 (N_6269,N_6148,N_6084);
and U6270 (N_6270,N_6065,N_6053);
nor U6271 (N_6271,N_6067,N_6189);
or U6272 (N_6272,N_6004,N_6034);
and U6273 (N_6273,N_6029,N_6021);
nor U6274 (N_6274,N_6022,N_6007);
and U6275 (N_6275,N_6071,N_6123);
nor U6276 (N_6276,N_6068,N_6114);
and U6277 (N_6277,N_6047,N_6174);
nor U6278 (N_6278,N_6033,N_6151);
nand U6279 (N_6279,N_6014,N_6046);
nand U6280 (N_6280,N_6086,N_6090);
and U6281 (N_6281,N_6158,N_6079);
and U6282 (N_6282,N_6109,N_6138);
and U6283 (N_6283,N_6036,N_6064);
nor U6284 (N_6284,N_6122,N_6012);
and U6285 (N_6285,N_6177,N_6131);
nand U6286 (N_6286,N_6150,N_6116);
and U6287 (N_6287,N_6161,N_6154);
nand U6288 (N_6288,N_6098,N_6162);
nor U6289 (N_6289,N_6087,N_6173);
and U6290 (N_6290,N_6072,N_6063);
nor U6291 (N_6291,N_6051,N_6024);
or U6292 (N_6292,N_6048,N_6188);
nor U6293 (N_6293,N_6028,N_6102);
or U6294 (N_6294,N_6144,N_6117);
nand U6295 (N_6295,N_6101,N_6052);
and U6296 (N_6296,N_6094,N_6145);
nor U6297 (N_6297,N_6112,N_6171);
and U6298 (N_6298,N_6107,N_6127);
or U6299 (N_6299,N_6169,N_6120);
nor U6300 (N_6300,N_6084,N_6040);
or U6301 (N_6301,N_6020,N_6193);
nor U6302 (N_6302,N_6133,N_6062);
and U6303 (N_6303,N_6171,N_6139);
nor U6304 (N_6304,N_6115,N_6087);
and U6305 (N_6305,N_6030,N_6075);
nand U6306 (N_6306,N_6162,N_6076);
nor U6307 (N_6307,N_6158,N_6024);
or U6308 (N_6308,N_6155,N_6151);
or U6309 (N_6309,N_6033,N_6008);
nand U6310 (N_6310,N_6114,N_6080);
or U6311 (N_6311,N_6003,N_6069);
or U6312 (N_6312,N_6198,N_6122);
nor U6313 (N_6313,N_6165,N_6185);
and U6314 (N_6314,N_6183,N_6100);
nor U6315 (N_6315,N_6114,N_6082);
or U6316 (N_6316,N_6022,N_6103);
nand U6317 (N_6317,N_6104,N_6050);
nand U6318 (N_6318,N_6117,N_6126);
nand U6319 (N_6319,N_6097,N_6106);
or U6320 (N_6320,N_6079,N_6099);
nand U6321 (N_6321,N_6152,N_6018);
or U6322 (N_6322,N_6081,N_6189);
nor U6323 (N_6323,N_6179,N_6076);
nor U6324 (N_6324,N_6039,N_6142);
and U6325 (N_6325,N_6042,N_6110);
nand U6326 (N_6326,N_6167,N_6104);
nor U6327 (N_6327,N_6134,N_6078);
and U6328 (N_6328,N_6110,N_6092);
or U6329 (N_6329,N_6092,N_6082);
or U6330 (N_6330,N_6051,N_6050);
or U6331 (N_6331,N_6175,N_6185);
nand U6332 (N_6332,N_6053,N_6051);
or U6333 (N_6333,N_6166,N_6034);
nand U6334 (N_6334,N_6138,N_6119);
nor U6335 (N_6335,N_6063,N_6056);
nand U6336 (N_6336,N_6116,N_6070);
or U6337 (N_6337,N_6181,N_6047);
nand U6338 (N_6338,N_6094,N_6002);
nor U6339 (N_6339,N_6046,N_6110);
nand U6340 (N_6340,N_6107,N_6194);
nor U6341 (N_6341,N_6112,N_6131);
and U6342 (N_6342,N_6084,N_6118);
or U6343 (N_6343,N_6087,N_6133);
nor U6344 (N_6344,N_6179,N_6136);
or U6345 (N_6345,N_6096,N_6120);
nor U6346 (N_6346,N_6188,N_6020);
or U6347 (N_6347,N_6184,N_6103);
and U6348 (N_6348,N_6127,N_6036);
or U6349 (N_6349,N_6098,N_6048);
nor U6350 (N_6350,N_6182,N_6149);
nand U6351 (N_6351,N_6191,N_6075);
and U6352 (N_6352,N_6049,N_6057);
or U6353 (N_6353,N_6107,N_6044);
and U6354 (N_6354,N_6106,N_6008);
and U6355 (N_6355,N_6078,N_6035);
and U6356 (N_6356,N_6136,N_6047);
nand U6357 (N_6357,N_6013,N_6082);
nand U6358 (N_6358,N_6151,N_6132);
nand U6359 (N_6359,N_6065,N_6058);
nor U6360 (N_6360,N_6069,N_6187);
nor U6361 (N_6361,N_6088,N_6072);
nor U6362 (N_6362,N_6072,N_6086);
nor U6363 (N_6363,N_6086,N_6186);
or U6364 (N_6364,N_6176,N_6088);
or U6365 (N_6365,N_6011,N_6004);
or U6366 (N_6366,N_6152,N_6027);
or U6367 (N_6367,N_6119,N_6160);
nor U6368 (N_6368,N_6035,N_6164);
nand U6369 (N_6369,N_6120,N_6160);
nor U6370 (N_6370,N_6124,N_6063);
or U6371 (N_6371,N_6083,N_6169);
nand U6372 (N_6372,N_6054,N_6038);
nor U6373 (N_6373,N_6113,N_6069);
nand U6374 (N_6374,N_6113,N_6050);
or U6375 (N_6375,N_6053,N_6075);
nand U6376 (N_6376,N_6198,N_6082);
nor U6377 (N_6377,N_6111,N_6180);
nand U6378 (N_6378,N_6187,N_6079);
or U6379 (N_6379,N_6155,N_6187);
or U6380 (N_6380,N_6145,N_6177);
nand U6381 (N_6381,N_6031,N_6194);
and U6382 (N_6382,N_6058,N_6126);
and U6383 (N_6383,N_6064,N_6024);
nand U6384 (N_6384,N_6003,N_6153);
and U6385 (N_6385,N_6177,N_6157);
nor U6386 (N_6386,N_6098,N_6161);
or U6387 (N_6387,N_6152,N_6101);
or U6388 (N_6388,N_6164,N_6160);
nor U6389 (N_6389,N_6147,N_6140);
and U6390 (N_6390,N_6112,N_6047);
and U6391 (N_6391,N_6120,N_6070);
or U6392 (N_6392,N_6132,N_6123);
nand U6393 (N_6393,N_6010,N_6060);
or U6394 (N_6394,N_6194,N_6154);
nor U6395 (N_6395,N_6152,N_6047);
and U6396 (N_6396,N_6168,N_6125);
nor U6397 (N_6397,N_6035,N_6046);
or U6398 (N_6398,N_6040,N_6178);
nor U6399 (N_6399,N_6158,N_6075);
nand U6400 (N_6400,N_6399,N_6206);
nand U6401 (N_6401,N_6299,N_6228);
nand U6402 (N_6402,N_6305,N_6216);
or U6403 (N_6403,N_6300,N_6252);
nand U6404 (N_6404,N_6363,N_6222);
nand U6405 (N_6405,N_6295,N_6294);
nand U6406 (N_6406,N_6397,N_6273);
nand U6407 (N_6407,N_6351,N_6359);
nor U6408 (N_6408,N_6229,N_6379);
and U6409 (N_6409,N_6266,N_6296);
or U6410 (N_6410,N_6377,N_6395);
and U6411 (N_6411,N_6327,N_6245);
or U6412 (N_6412,N_6366,N_6388);
and U6413 (N_6413,N_6224,N_6272);
nor U6414 (N_6414,N_6251,N_6345);
nor U6415 (N_6415,N_6315,N_6372);
nand U6416 (N_6416,N_6217,N_6280);
nand U6417 (N_6417,N_6339,N_6244);
and U6418 (N_6418,N_6317,N_6328);
or U6419 (N_6419,N_6380,N_6355);
nor U6420 (N_6420,N_6258,N_6331);
or U6421 (N_6421,N_6354,N_6311);
or U6422 (N_6422,N_6264,N_6218);
and U6423 (N_6423,N_6236,N_6239);
and U6424 (N_6424,N_6277,N_6226);
or U6425 (N_6425,N_6319,N_6338);
nor U6426 (N_6426,N_6233,N_6282);
nand U6427 (N_6427,N_6361,N_6304);
and U6428 (N_6428,N_6204,N_6227);
or U6429 (N_6429,N_6394,N_6326);
nand U6430 (N_6430,N_6374,N_6215);
nor U6431 (N_6431,N_6383,N_6312);
nand U6432 (N_6432,N_6238,N_6265);
nand U6433 (N_6433,N_6353,N_6389);
nor U6434 (N_6434,N_6385,N_6332);
nor U6435 (N_6435,N_6203,N_6335);
and U6436 (N_6436,N_6302,N_6391);
nor U6437 (N_6437,N_6292,N_6316);
nor U6438 (N_6438,N_6211,N_6220);
or U6439 (N_6439,N_6314,N_6392);
or U6440 (N_6440,N_6358,N_6253);
nor U6441 (N_6441,N_6381,N_6221);
nor U6442 (N_6442,N_6369,N_6320);
nand U6443 (N_6443,N_6365,N_6364);
nand U6444 (N_6444,N_6207,N_6213);
nor U6445 (N_6445,N_6368,N_6370);
nand U6446 (N_6446,N_6376,N_6308);
nor U6447 (N_6447,N_6241,N_6254);
and U6448 (N_6448,N_6202,N_6200);
or U6449 (N_6449,N_6344,N_6293);
nand U6450 (N_6450,N_6356,N_6340);
nand U6451 (N_6451,N_6349,N_6271);
or U6452 (N_6452,N_6318,N_6255);
and U6453 (N_6453,N_6362,N_6303);
and U6454 (N_6454,N_6278,N_6274);
or U6455 (N_6455,N_6384,N_6260);
xor U6456 (N_6456,N_6256,N_6393);
nand U6457 (N_6457,N_6270,N_6343);
or U6458 (N_6458,N_6259,N_6350);
or U6459 (N_6459,N_6231,N_6262);
and U6460 (N_6460,N_6298,N_6247);
or U6461 (N_6461,N_6232,N_6219);
and U6462 (N_6462,N_6321,N_6285);
nor U6463 (N_6463,N_6284,N_6261);
or U6464 (N_6464,N_6223,N_6225);
nand U6465 (N_6465,N_6212,N_6240);
nand U6466 (N_6466,N_6230,N_6378);
or U6467 (N_6467,N_6382,N_6214);
or U6468 (N_6468,N_6337,N_6275);
or U6469 (N_6469,N_6333,N_6286);
or U6470 (N_6470,N_6267,N_6289);
and U6471 (N_6471,N_6210,N_6387);
or U6472 (N_6472,N_6242,N_6396);
nor U6473 (N_6473,N_6341,N_6234);
nor U6474 (N_6474,N_6324,N_6386);
nand U6475 (N_6475,N_6297,N_6243);
nand U6476 (N_6476,N_6309,N_6246);
nor U6477 (N_6477,N_6257,N_6360);
nor U6478 (N_6478,N_6334,N_6357);
and U6479 (N_6479,N_6310,N_6371);
nand U6480 (N_6480,N_6276,N_6279);
nor U6481 (N_6481,N_6250,N_6235);
nor U6482 (N_6482,N_6346,N_6249);
nor U6483 (N_6483,N_6352,N_6288);
nor U6484 (N_6484,N_6283,N_6237);
or U6485 (N_6485,N_6330,N_6201);
or U6486 (N_6486,N_6390,N_6268);
or U6487 (N_6487,N_6323,N_6208);
and U6488 (N_6488,N_6248,N_6306);
or U6489 (N_6489,N_6269,N_6301);
and U6490 (N_6490,N_6329,N_6281);
nor U6491 (N_6491,N_6209,N_6342);
nor U6492 (N_6492,N_6375,N_6348);
or U6493 (N_6493,N_6205,N_6336);
nor U6494 (N_6494,N_6263,N_6347);
nor U6495 (N_6495,N_6367,N_6373);
nor U6496 (N_6496,N_6325,N_6291);
nor U6497 (N_6497,N_6322,N_6307);
or U6498 (N_6498,N_6313,N_6290);
nand U6499 (N_6499,N_6287,N_6398);
nand U6500 (N_6500,N_6274,N_6351);
nand U6501 (N_6501,N_6263,N_6338);
or U6502 (N_6502,N_6263,N_6356);
or U6503 (N_6503,N_6275,N_6394);
nand U6504 (N_6504,N_6384,N_6211);
nand U6505 (N_6505,N_6295,N_6246);
nand U6506 (N_6506,N_6273,N_6373);
nand U6507 (N_6507,N_6281,N_6332);
or U6508 (N_6508,N_6279,N_6217);
or U6509 (N_6509,N_6301,N_6332);
or U6510 (N_6510,N_6203,N_6385);
nor U6511 (N_6511,N_6282,N_6361);
nand U6512 (N_6512,N_6381,N_6228);
or U6513 (N_6513,N_6328,N_6283);
and U6514 (N_6514,N_6369,N_6258);
nor U6515 (N_6515,N_6310,N_6202);
or U6516 (N_6516,N_6235,N_6324);
or U6517 (N_6517,N_6298,N_6231);
or U6518 (N_6518,N_6358,N_6207);
and U6519 (N_6519,N_6291,N_6370);
or U6520 (N_6520,N_6326,N_6390);
nand U6521 (N_6521,N_6397,N_6300);
and U6522 (N_6522,N_6207,N_6287);
or U6523 (N_6523,N_6343,N_6264);
nand U6524 (N_6524,N_6382,N_6259);
and U6525 (N_6525,N_6279,N_6271);
or U6526 (N_6526,N_6308,N_6209);
nand U6527 (N_6527,N_6319,N_6391);
nor U6528 (N_6528,N_6295,N_6285);
or U6529 (N_6529,N_6287,N_6386);
nand U6530 (N_6530,N_6265,N_6346);
nand U6531 (N_6531,N_6203,N_6276);
nor U6532 (N_6532,N_6369,N_6245);
or U6533 (N_6533,N_6356,N_6377);
nand U6534 (N_6534,N_6382,N_6309);
nor U6535 (N_6535,N_6389,N_6359);
nor U6536 (N_6536,N_6248,N_6264);
and U6537 (N_6537,N_6287,N_6229);
nor U6538 (N_6538,N_6201,N_6393);
and U6539 (N_6539,N_6341,N_6201);
and U6540 (N_6540,N_6287,N_6355);
xnor U6541 (N_6541,N_6340,N_6367);
or U6542 (N_6542,N_6269,N_6261);
or U6543 (N_6543,N_6330,N_6239);
nor U6544 (N_6544,N_6284,N_6388);
and U6545 (N_6545,N_6240,N_6306);
and U6546 (N_6546,N_6323,N_6343);
and U6547 (N_6547,N_6364,N_6246);
and U6548 (N_6548,N_6271,N_6362);
or U6549 (N_6549,N_6385,N_6390);
nor U6550 (N_6550,N_6304,N_6384);
nand U6551 (N_6551,N_6367,N_6310);
and U6552 (N_6552,N_6219,N_6223);
nor U6553 (N_6553,N_6343,N_6283);
and U6554 (N_6554,N_6211,N_6274);
nor U6555 (N_6555,N_6294,N_6371);
nand U6556 (N_6556,N_6284,N_6276);
nor U6557 (N_6557,N_6250,N_6242);
and U6558 (N_6558,N_6296,N_6290);
or U6559 (N_6559,N_6253,N_6368);
nor U6560 (N_6560,N_6363,N_6231);
and U6561 (N_6561,N_6235,N_6328);
or U6562 (N_6562,N_6386,N_6231);
nand U6563 (N_6563,N_6204,N_6282);
or U6564 (N_6564,N_6218,N_6246);
nor U6565 (N_6565,N_6208,N_6373);
and U6566 (N_6566,N_6223,N_6363);
xor U6567 (N_6567,N_6280,N_6335);
or U6568 (N_6568,N_6283,N_6314);
nor U6569 (N_6569,N_6302,N_6266);
nor U6570 (N_6570,N_6322,N_6273);
nor U6571 (N_6571,N_6258,N_6387);
nand U6572 (N_6572,N_6210,N_6300);
or U6573 (N_6573,N_6340,N_6216);
nor U6574 (N_6574,N_6366,N_6226);
nand U6575 (N_6575,N_6216,N_6296);
or U6576 (N_6576,N_6334,N_6276);
and U6577 (N_6577,N_6220,N_6389);
nor U6578 (N_6578,N_6380,N_6210);
nand U6579 (N_6579,N_6232,N_6379);
or U6580 (N_6580,N_6304,N_6339);
nor U6581 (N_6581,N_6374,N_6360);
or U6582 (N_6582,N_6297,N_6366);
and U6583 (N_6583,N_6279,N_6282);
or U6584 (N_6584,N_6298,N_6215);
and U6585 (N_6585,N_6258,N_6224);
and U6586 (N_6586,N_6390,N_6245);
nand U6587 (N_6587,N_6341,N_6259);
nand U6588 (N_6588,N_6203,N_6345);
nor U6589 (N_6589,N_6248,N_6298);
nand U6590 (N_6590,N_6250,N_6380);
nor U6591 (N_6591,N_6211,N_6279);
nand U6592 (N_6592,N_6229,N_6216);
nor U6593 (N_6593,N_6384,N_6246);
nand U6594 (N_6594,N_6371,N_6213);
and U6595 (N_6595,N_6285,N_6256);
and U6596 (N_6596,N_6355,N_6366);
nor U6597 (N_6597,N_6219,N_6371);
and U6598 (N_6598,N_6358,N_6229);
and U6599 (N_6599,N_6283,N_6361);
and U6600 (N_6600,N_6468,N_6479);
or U6601 (N_6601,N_6503,N_6437);
nand U6602 (N_6602,N_6554,N_6444);
nand U6603 (N_6603,N_6412,N_6555);
or U6604 (N_6604,N_6516,N_6509);
nor U6605 (N_6605,N_6404,N_6462);
nand U6606 (N_6606,N_6517,N_6576);
nand U6607 (N_6607,N_6442,N_6507);
xor U6608 (N_6608,N_6400,N_6458);
and U6609 (N_6609,N_6460,N_6480);
or U6610 (N_6610,N_6512,N_6569);
and U6611 (N_6611,N_6505,N_6408);
or U6612 (N_6612,N_6545,N_6514);
or U6613 (N_6613,N_6560,N_6574);
nand U6614 (N_6614,N_6584,N_6449);
or U6615 (N_6615,N_6448,N_6552);
and U6616 (N_6616,N_6414,N_6447);
and U6617 (N_6617,N_6575,N_6527);
nand U6618 (N_6618,N_6522,N_6543);
or U6619 (N_6619,N_6577,N_6453);
or U6620 (N_6620,N_6536,N_6487);
nand U6621 (N_6621,N_6562,N_6493);
nor U6622 (N_6622,N_6579,N_6494);
or U6623 (N_6623,N_6464,N_6565);
or U6624 (N_6624,N_6415,N_6586);
or U6625 (N_6625,N_6438,N_6525);
or U6626 (N_6626,N_6434,N_6417);
nor U6627 (N_6627,N_6418,N_6590);
nand U6628 (N_6628,N_6403,N_6549);
nor U6629 (N_6629,N_6583,N_6495);
and U6630 (N_6630,N_6591,N_6523);
and U6631 (N_6631,N_6445,N_6524);
nor U6632 (N_6632,N_6451,N_6465);
nor U6633 (N_6633,N_6508,N_6501);
or U6634 (N_6634,N_6567,N_6588);
nor U6635 (N_6635,N_6564,N_6500);
or U6636 (N_6636,N_6520,N_6497);
nor U6637 (N_6637,N_6419,N_6450);
nand U6638 (N_6638,N_6553,N_6413);
and U6639 (N_6639,N_6530,N_6506);
nor U6640 (N_6640,N_6484,N_6428);
and U6641 (N_6641,N_6513,N_6592);
or U6642 (N_6642,N_6573,N_6459);
nand U6643 (N_6643,N_6491,N_6425);
nand U6644 (N_6644,N_6597,N_6589);
and U6645 (N_6645,N_6538,N_6475);
nand U6646 (N_6646,N_6488,N_6572);
nor U6647 (N_6647,N_6593,N_6424);
nor U6648 (N_6648,N_6529,N_6594);
nor U6649 (N_6649,N_6490,N_6581);
nand U6650 (N_6650,N_6566,N_6481);
nand U6651 (N_6651,N_6433,N_6528);
nor U6652 (N_6652,N_6492,N_6410);
nand U6653 (N_6653,N_6446,N_6471);
or U6654 (N_6654,N_6580,N_6570);
nand U6655 (N_6655,N_6482,N_6466);
nand U6656 (N_6656,N_6532,N_6441);
or U6657 (N_6657,N_6443,N_6405);
or U6658 (N_6658,N_6456,N_6402);
or U6659 (N_6659,N_6539,N_6485);
or U6660 (N_6660,N_6546,N_6511);
nand U6661 (N_6661,N_6587,N_6498);
nor U6662 (N_6662,N_6502,N_6541);
nor U6663 (N_6663,N_6537,N_6401);
nor U6664 (N_6664,N_6432,N_6521);
and U6665 (N_6665,N_6440,N_6469);
nor U6666 (N_6666,N_6429,N_6473);
nor U6667 (N_6667,N_6457,N_6426);
nor U6668 (N_6668,N_6476,N_6470);
nand U6669 (N_6669,N_6435,N_6474);
nor U6670 (N_6670,N_6409,N_6406);
nor U6671 (N_6671,N_6550,N_6407);
and U6672 (N_6672,N_6531,N_6571);
or U6673 (N_6673,N_6430,N_6431);
nor U6674 (N_6674,N_6499,N_6518);
and U6675 (N_6675,N_6504,N_6422);
nand U6676 (N_6676,N_6472,N_6547);
and U6677 (N_6677,N_6535,N_6439);
and U6678 (N_6678,N_6578,N_6540);
or U6679 (N_6679,N_6533,N_6582);
or U6680 (N_6680,N_6452,N_6542);
nand U6681 (N_6681,N_6548,N_6568);
and U6682 (N_6682,N_6486,N_6599);
nand U6683 (N_6683,N_6436,N_6427);
or U6684 (N_6684,N_6461,N_6598);
and U6685 (N_6685,N_6519,N_6558);
nand U6686 (N_6686,N_6421,N_6455);
nand U6687 (N_6687,N_6551,N_6416);
nand U6688 (N_6688,N_6596,N_6477);
or U6689 (N_6689,N_6423,N_6585);
xor U6690 (N_6690,N_6557,N_6534);
or U6691 (N_6691,N_6496,N_6467);
nand U6692 (N_6692,N_6595,N_6411);
or U6693 (N_6693,N_6526,N_6561);
or U6694 (N_6694,N_6420,N_6556);
or U6695 (N_6695,N_6483,N_6454);
or U6696 (N_6696,N_6515,N_6463);
or U6697 (N_6697,N_6489,N_6563);
or U6698 (N_6698,N_6510,N_6478);
nor U6699 (N_6699,N_6544,N_6559);
nand U6700 (N_6700,N_6579,N_6516);
and U6701 (N_6701,N_6447,N_6479);
and U6702 (N_6702,N_6594,N_6571);
or U6703 (N_6703,N_6596,N_6552);
nor U6704 (N_6704,N_6401,N_6515);
nand U6705 (N_6705,N_6424,N_6449);
and U6706 (N_6706,N_6459,N_6471);
nor U6707 (N_6707,N_6551,N_6489);
nor U6708 (N_6708,N_6596,N_6509);
nand U6709 (N_6709,N_6543,N_6511);
nand U6710 (N_6710,N_6436,N_6556);
or U6711 (N_6711,N_6489,N_6529);
nand U6712 (N_6712,N_6573,N_6570);
nand U6713 (N_6713,N_6405,N_6529);
nand U6714 (N_6714,N_6550,N_6420);
and U6715 (N_6715,N_6444,N_6429);
or U6716 (N_6716,N_6516,N_6581);
nor U6717 (N_6717,N_6414,N_6527);
nand U6718 (N_6718,N_6455,N_6463);
and U6719 (N_6719,N_6497,N_6470);
and U6720 (N_6720,N_6575,N_6483);
or U6721 (N_6721,N_6439,N_6522);
nor U6722 (N_6722,N_6442,N_6476);
nor U6723 (N_6723,N_6417,N_6470);
nor U6724 (N_6724,N_6575,N_6458);
nand U6725 (N_6725,N_6474,N_6550);
or U6726 (N_6726,N_6561,N_6435);
nand U6727 (N_6727,N_6589,N_6440);
nand U6728 (N_6728,N_6559,N_6560);
nor U6729 (N_6729,N_6487,N_6542);
nor U6730 (N_6730,N_6458,N_6535);
nand U6731 (N_6731,N_6598,N_6550);
or U6732 (N_6732,N_6448,N_6589);
nor U6733 (N_6733,N_6514,N_6590);
or U6734 (N_6734,N_6498,N_6444);
or U6735 (N_6735,N_6558,N_6504);
or U6736 (N_6736,N_6528,N_6594);
nor U6737 (N_6737,N_6527,N_6402);
or U6738 (N_6738,N_6530,N_6477);
and U6739 (N_6739,N_6580,N_6503);
or U6740 (N_6740,N_6587,N_6491);
nor U6741 (N_6741,N_6549,N_6534);
nor U6742 (N_6742,N_6457,N_6531);
nand U6743 (N_6743,N_6554,N_6416);
nand U6744 (N_6744,N_6552,N_6518);
nand U6745 (N_6745,N_6590,N_6598);
nor U6746 (N_6746,N_6433,N_6447);
and U6747 (N_6747,N_6522,N_6571);
nand U6748 (N_6748,N_6426,N_6568);
nor U6749 (N_6749,N_6497,N_6458);
and U6750 (N_6750,N_6506,N_6434);
and U6751 (N_6751,N_6552,N_6425);
and U6752 (N_6752,N_6480,N_6566);
nor U6753 (N_6753,N_6421,N_6466);
nor U6754 (N_6754,N_6564,N_6532);
nor U6755 (N_6755,N_6580,N_6553);
nand U6756 (N_6756,N_6598,N_6576);
or U6757 (N_6757,N_6594,N_6527);
nor U6758 (N_6758,N_6566,N_6520);
and U6759 (N_6759,N_6409,N_6483);
nand U6760 (N_6760,N_6448,N_6462);
or U6761 (N_6761,N_6528,N_6579);
nand U6762 (N_6762,N_6554,N_6479);
nor U6763 (N_6763,N_6589,N_6483);
and U6764 (N_6764,N_6492,N_6506);
and U6765 (N_6765,N_6530,N_6523);
or U6766 (N_6766,N_6517,N_6442);
or U6767 (N_6767,N_6524,N_6575);
and U6768 (N_6768,N_6416,N_6586);
or U6769 (N_6769,N_6418,N_6450);
nand U6770 (N_6770,N_6586,N_6585);
or U6771 (N_6771,N_6437,N_6523);
nand U6772 (N_6772,N_6475,N_6485);
nor U6773 (N_6773,N_6474,N_6458);
nor U6774 (N_6774,N_6574,N_6436);
or U6775 (N_6775,N_6569,N_6555);
and U6776 (N_6776,N_6531,N_6408);
and U6777 (N_6777,N_6433,N_6450);
nand U6778 (N_6778,N_6451,N_6540);
nand U6779 (N_6779,N_6454,N_6591);
or U6780 (N_6780,N_6517,N_6539);
nor U6781 (N_6781,N_6462,N_6504);
nand U6782 (N_6782,N_6593,N_6452);
nand U6783 (N_6783,N_6491,N_6585);
nor U6784 (N_6784,N_6567,N_6560);
nand U6785 (N_6785,N_6536,N_6439);
or U6786 (N_6786,N_6580,N_6525);
nor U6787 (N_6787,N_6568,N_6419);
or U6788 (N_6788,N_6591,N_6416);
or U6789 (N_6789,N_6598,N_6463);
or U6790 (N_6790,N_6551,N_6568);
and U6791 (N_6791,N_6533,N_6558);
and U6792 (N_6792,N_6437,N_6422);
nor U6793 (N_6793,N_6475,N_6527);
or U6794 (N_6794,N_6519,N_6512);
and U6795 (N_6795,N_6536,N_6486);
nor U6796 (N_6796,N_6514,N_6589);
or U6797 (N_6797,N_6471,N_6434);
or U6798 (N_6798,N_6456,N_6440);
nand U6799 (N_6799,N_6430,N_6488);
nand U6800 (N_6800,N_6716,N_6782);
and U6801 (N_6801,N_6713,N_6650);
nor U6802 (N_6802,N_6726,N_6763);
nor U6803 (N_6803,N_6785,N_6731);
nand U6804 (N_6804,N_6610,N_6638);
and U6805 (N_6805,N_6669,N_6769);
and U6806 (N_6806,N_6693,N_6625);
and U6807 (N_6807,N_6639,N_6705);
and U6808 (N_6808,N_6766,N_6758);
nor U6809 (N_6809,N_6697,N_6706);
and U6810 (N_6810,N_6665,N_6779);
or U6811 (N_6811,N_6725,N_6608);
and U6812 (N_6812,N_6735,N_6702);
nor U6813 (N_6813,N_6688,N_6730);
and U6814 (N_6814,N_6627,N_6717);
or U6815 (N_6815,N_6745,N_6795);
nand U6816 (N_6816,N_6759,N_6695);
and U6817 (N_6817,N_6663,N_6617);
or U6818 (N_6818,N_6724,N_6704);
nor U6819 (N_6819,N_6799,N_6710);
nand U6820 (N_6820,N_6684,N_6618);
nand U6821 (N_6821,N_6788,N_6649);
nand U6822 (N_6822,N_6728,N_6753);
or U6823 (N_6823,N_6796,N_6708);
nand U6824 (N_6824,N_6683,N_6620);
or U6825 (N_6825,N_6700,N_6671);
nor U6826 (N_6826,N_6630,N_6622);
nand U6827 (N_6827,N_6668,N_6611);
or U6828 (N_6828,N_6723,N_6784);
nor U6829 (N_6829,N_6609,N_6616);
or U6830 (N_6830,N_6699,N_6628);
nor U6831 (N_6831,N_6774,N_6701);
nand U6832 (N_6832,N_6648,N_6748);
nor U6833 (N_6833,N_6743,N_6685);
nand U6834 (N_6834,N_6679,N_6652);
or U6835 (N_6835,N_6798,N_6780);
or U6836 (N_6836,N_6734,N_6692);
and U6837 (N_6837,N_6778,N_6757);
or U6838 (N_6838,N_6719,N_6689);
nand U6839 (N_6839,N_6667,N_6786);
nand U6840 (N_6840,N_6661,N_6658);
or U6841 (N_6841,N_6767,N_6793);
and U6842 (N_6842,N_6614,N_6764);
nor U6843 (N_6843,N_6605,N_6729);
nor U6844 (N_6844,N_6623,N_6682);
nor U6845 (N_6845,N_6612,N_6755);
or U6846 (N_6846,N_6613,N_6791);
or U6847 (N_6847,N_6727,N_6773);
or U6848 (N_6848,N_6742,N_6690);
or U6849 (N_6849,N_6637,N_6670);
and U6850 (N_6850,N_6740,N_6651);
nand U6851 (N_6851,N_6681,N_6624);
nor U6852 (N_6852,N_6747,N_6754);
xor U6853 (N_6853,N_6662,N_6744);
nand U6854 (N_6854,N_6765,N_6632);
or U6855 (N_6855,N_6736,N_6703);
and U6856 (N_6856,N_6711,N_6659);
nand U6857 (N_6857,N_6721,N_6790);
or U6858 (N_6858,N_6657,N_6646);
nor U6859 (N_6859,N_6672,N_6750);
nor U6860 (N_6860,N_6709,N_6633);
and U6861 (N_6861,N_6707,N_6676);
nor U6862 (N_6862,N_6615,N_6756);
nor U6863 (N_6863,N_6792,N_6698);
or U6864 (N_6864,N_6664,N_6635);
nor U6865 (N_6865,N_6660,N_6720);
nor U6866 (N_6866,N_6644,N_6601);
and U6867 (N_6867,N_6645,N_6797);
or U6868 (N_6868,N_6737,N_6762);
and U6869 (N_6869,N_6732,N_6783);
nor U6870 (N_6870,N_6600,N_6642);
or U6871 (N_6871,N_6654,N_6772);
and U6872 (N_6872,N_6718,N_6634);
nand U6873 (N_6873,N_6738,N_6640);
or U6874 (N_6874,N_6687,N_6673);
nand U6875 (N_6875,N_6770,N_6722);
nand U6876 (N_6876,N_6678,N_6636);
and U6877 (N_6877,N_6733,N_6787);
nor U6878 (N_6878,N_6775,N_6771);
or U6879 (N_6879,N_6604,N_6607);
nor U6880 (N_6880,N_6641,N_6696);
nor U6881 (N_6881,N_6666,N_6626);
and U6882 (N_6882,N_6746,N_6686);
nor U6883 (N_6883,N_6749,N_6619);
and U6884 (N_6884,N_6694,N_6655);
nor U6885 (N_6885,N_6629,N_6631);
or U6886 (N_6886,N_6606,N_6680);
or U6887 (N_6887,N_6777,N_6603);
nor U6888 (N_6888,N_6789,N_6647);
nand U6889 (N_6889,N_6643,N_6794);
or U6890 (N_6890,N_6761,N_6653);
and U6891 (N_6891,N_6781,N_6602);
nor U6892 (N_6892,N_6741,N_6712);
nor U6893 (N_6893,N_6751,N_6691);
and U6894 (N_6894,N_6677,N_6760);
nand U6895 (N_6895,N_6739,N_6675);
and U6896 (N_6896,N_6752,N_6621);
nor U6897 (N_6897,N_6715,N_6674);
and U6898 (N_6898,N_6768,N_6656);
or U6899 (N_6899,N_6714,N_6776);
and U6900 (N_6900,N_6716,N_6659);
nand U6901 (N_6901,N_6763,N_6689);
and U6902 (N_6902,N_6650,N_6719);
nand U6903 (N_6903,N_6609,N_6620);
or U6904 (N_6904,N_6704,N_6766);
and U6905 (N_6905,N_6650,N_6746);
nand U6906 (N_6906,N_6621,N_6639);
or U6907 (N_6907,N_6642,N_6771);
or U6908 (N_6908,N_6633,N_6625);
nand U6909 (N_6909,N_6739,N_6666);
nor U6910 (N_6910,N_6790,N_6745);
and U6911 (N_6911,N_6642,N_6666);
nand U6912 (N_6912,N_6648,N_6722);
or U6913 (N_6913,N_6647,N_6777);
nor U6914 (N_6914,N_6684,N_6794);
nand U6915 (N_6915,N_6763,N_6664);
nand U6916 (N_6916,N_6700,N_6789);
and U6917 (N_6917,N_6746,N_6784);
or U6918 (N_6918,N_6741,N_6732);
or U6919 (N_6919,N_6728,N_6762);
and U6920 (N_6920,N_6699,N_6601);
and U6921 (N_6921,N_6621,N_6660);
and U6922 (N_6922,N_6677,N_6651);
or U6923 (N_6923,N_6666,N_6629);
and U6924 (N_6924,N_6695,N_6628);
nand U6925 (N_6925,N_6639,N_6726);
and U6926 (N_6926,N_6788,N_6677);
nor U6927 (N_6927,N_6651,N_6769);
and U6928 (N_6928,N_6650,N_6720);
and U6929 (N_6929,N_6736,N_6727);
nand U6930 (N_6930,N_6694,N_6692);
nand U6931 (N_6931,N_6657,N_6716);
and U6932 (N_6932,N_6658,N_6734);
nand U6933 (N_6933,N_6792,N_6793);
and U6934 (N_6934,N_6679,N_6647);
and U6935 (N_6935,N_6707,N_6770);
nor U6936 (N_6936,N_6786,N_6675);
nor U6937 (N_6937,N_6763,N_6673);
nand U6938 (N_6938,N_6756,N_6745);
or U6939 (N_6939,N_6649,N_6729);
or U6940 (N_6940,N_6672,N_6787);
and U6941 (N_6941,N_6780,N_6734);
and U6942 (N_6942,N_6759,N_6746);
or U6943 (N_6943,N_6636,N_6624);
nand U6944 (N_6944,N_6625,N_6742);
and U6945 (N_6945,N_6657,N_6625);
nor U6946 (N_6946,N_6760,N_6636);
nor U6947 (N_6947,N_6769,N_6788);
nand U6948 (N_6948,N_6648,N_6730);
and U6949 (N_6949,N_6720,N_6768);
nand U6950 (N_6950,N_6750,N_6659);
or U6951 (N_6951,N_6773,N_6685);
or U6952 (N_6952,N_6638,N_6692);
nor U6953 (N_6953,N_6728,N_6616);
or U6954 (N_6954,N_6672,N_6658);
or U6955 (N_6955,N_6698,N_6714);
or U6956 (N_6956,N_6615,N_6667);
and U6957 (N_6957,N_6730,N_6764);
nand U6958 (N_6958,N_6706,N_6772);
nand U6959 (N_6959,N_6753,N_6657);
nand U6960 (N_6960,N_6695,N_6729);
or U6961 (N_6961,N_6746,N_6728);
and U6962 (N_6962,N_6731,N_6720);
or U6963 (N_6963,N_6612,N_6618);
or U6964 (N_6964,N_6783,N_6757);
and U6965 (N_6965,N_6769,N_6712);
or U6966 (N_6966,N_6610,N_6722);
and U6967 (N_6967,N_6668,N_6799);
and U6968 (N_6968,N_6716,N_6610);
nand U6969 (N_6969,N_6730,N_6659);
nor U6970 (N_6970,N_6735,N_6742);
or U6971 (N_6971,N_6726,N_6646);
and U6972 (N_6972,N_6675,N_6777);
nand U6973 (N_6973,N_6640,N_6716);
and U6974 (N_6974,N_6733,N_6732);
nor U6975 (N_6975,N_6765,N_6709);
and U6976 (N_6976,N_6699,N_6657);
and U6977 (N_6977,N_6629,N_6657);
nor U6978 (N_6978,N_6780,N_6773);
nand U6979 (N_6979,N_6626,N_6749);
and U6980 (N_6980,N_6790,N_6648);
or U6981 (N_6981,N_6776,N_6618);
nand U6982 (N_6982,N_6666,N_6699);
and U6983 (N_6983,N_6625,N_6678);
nand U6984 (N_6984,N_6747,N_6622);
nand U6985 (N_6985,N_6604,N_6643);
and U6986 (N_6986,N_6759,N_6658);
nand U6987 (N_6987,N_6652,N_6646);
and U6988 (N_6988,N_6695,N_6743);
and U6989 (N_6989,N_6721,N_6702);
and U6990 (N_6990,N_6711,N_6639);
and U6991 (N_6991,N_6642,N_6658);
and U6992 (N_6992,N_6656,N_6774);
nor U6993 (N_6993,N_6723,N_6682);
nand U6994 (N_6994,N_6761,N_6773);
nand U6995 (N_6995,N_6607,N_6774);
nand U6996 (N_6996,N_6776,N_6791);
and U6997 (N_6997,N_6656,N_6626);
nand U6998 (N_6998,N_6693,N_6708);
nor U6999 (N_6999,N_6793,N_6787);
nor U7000 (N_7000,N_6823,N_6997);
or U7001 (N_7001,N_6954,N_6821);
or U7002 (N_7002,N_6816,N_6933);
or U7003 (N_7003,N_6846,N_6886);
nand U7004 (N_7004,N_6803,N_6829);
and U7005 (N_7005,N_6976,N_6959);
and U7006 (N_7006,N_6894,N_6979);
nand U7007 (N_7007,N_6945,N_6918);
or U7008 (N_7008,N_6830,N_6801);
nor U7009 (N_7009,N_6833,N_6917);
nand U7010 (N_7010,N_6863,N_6855);
or U7011 (N_7011,N_6842,N_6991);
nand U7012 (N_7012,N_6968,N_6864);
nand U7013 (N_7013,N_6982,N_6893);
nor U7014 (N_7014,N_6929,N_6880);
or U7015 (N_7015,N_6818,N_6868);
or U7016 (N_7016,N_6998,N_6873);
or U7017 (N_7017,N_6857,N_6972);
nor U7018 (N_7018,N_6812,N_6879);
nor U7019 (N_7019,N_6937,N_6810);
or U7020 (N_7020,N_6966,N_6882);
nor U7021 (N_7021,N_6862,N_6804);
nand U7022 (N_7022,N_6844,N_6969);
and U7023 (N_7023,N_6885,N_6811);
nor U7024 (N_7024,N_6974,N_6944);
and U7025 (N_7025,N_6908,N_6853);
and U7026 (N_7026,N_6922,N_6876);
and U7027 (N_7027,N_6946,N_6978);
and U7028 (N_7028,N_6934,N_6836);
nor U7029 (N_7029,N_6874,N_6825);
nor U7030 (N_7030,N_6985,N_6884);
nand U7031 (N_7031,N_6955,N_6820);
nand U7032 (N_7032,N_6947,N_6904);
nor U7033 (N_7033,N_6926,N_6807);
nand U7034 (N_7034,N_6952,N_6980);
nand U7035 (N_7035,N_6819,N_6808);
nand U7036 (N_7036,N_6851,N_6900);
nor U7037 (N_7037,N_6941,N_6925);
and U7038 (N_7038,N_6861,N_6957);
and U7039 (N_7039,N_6964,N_6914);
nor U7040 (N_7040,N_6981,N_6865);
and U7041 (N_7041,N_6814,N_6907);
nand U7042 (N_7042,N_6815,N_6951);
nand U7043 (N_7043,N_6867,N_6877);
and U7044 (N_7044,N_6827,N_6860);
nand U7045 (N_7045,N_6870,N_6943);
nor U7046 (N_7046,N_6909,N_6965);
nor U7047 (N_7047,N_6809,N_6931);
nor U7048 (N_7048,N_6826,N_6845);
nand U7049 (N_7049,N_6813,N_6849);
nand U7050 (N_7050,N_6817,N_6989);
or U7051 (N_7051,N_6971,N_6986);
and U7052 (N_7052,N_6923,N_6948);
or U7053 (N_7053,N_6856,N_6839);
nand U7054 (N_7054,N_6924,N_6854);
and U7055 (N_7055,N_6837,N_6970);
nor U7056 (N_7056,N_6905,N_6866);
or U7057 (N_7057,N_6912,N_6953);
and U7058 (N_7058,N_6872,N_6805);
nand U7059 (N_7059,N_6987,N_6848);
and U7060 (N_7060,N_6967,N_6939);
nand U7061 (N_7061,N_6895,N_6901);
or U7062 (N_7062,N_6919,N_6938);
nor U7063 (N_7063,N_6962,N_6871);
nand U7064 (N_7064,N_6940,N_6834);
nor U7065 (N_7065,N_6913,N_6890);
and U7066 (N_7066,N_6960,N_6949);
nand U7067 (N_7067,N_6899,N_6992);
or U7068 (N_7068,N_6988,N_6878);
and U7069 (N_7069,N_6984,N_6994);
or U7070 (N_7070,N_6983,N_6843);
or U7071 (N_7071,N_6828,N_6806);
nor U7072 (N_7072,N_6892,N_6858);
and U7073 (N_7073,N_6869,N_6824);
nand U7074 (N_7074,N_6832,N_6936);
or U7075 (N_7075,N_6975,N_6915);
or U7076 (N_7076,N_6916,N_6928);
or U7077 (N_7077,N_6956,N_6896);
nand U7078 (N_7078,N_6996,N_6887);
nand U7079 (N_7079,N_6903,N_6950);
nand U7080 (N_7080,N_6831,N_6911);
or U7081 (N_7081,N_6888,N_6897);
or U7082 (N_7082,N_6881,N_6995);
nand U7083 (N_7083,N_6891,N_6822);
or U7084 (N_7084,N_6852,N_6920);
or U7085 (N_7085,N_6883,N_6906);
nand U7086 (N_7086,N_6841,N_6898);
nand U7087 (N_7087,N_6990,N_6921);
and U7088 (N_7088,N_6875,N_6930);
nand U7089 (N_7089,N_6977,N_6942);
nand U7090 (N_7090,N_6999,N_6859);
xor U7091 (N_7091,N_6850,N_6927);
nand U7092 (N_7092,N_6835,N_6840);
or U7093 (N_7093,N_6802,N_6993);
or U7094 (N_7094,N_6932,N_6800);
nor U7095 (N_7095,N_6902,N_6958);
nor U7096 (N_7096,N_6973,N_6889);
nand U7097 (N_7097,N_6935,N_6847);
and U7098 (N_7098,N_6838,N_6961);
and U7099 (N_7099,N_6910,N_6963);
nand U7100 (N_7100,N_6918,N_6890);
and U7101 (N_7101,N_6984,N_6906);
nor U7102 (N_7102,N_6881,N_6924);
or U7103 (N_7103,N_6830,N_6820);
and U7104 (N_7104,N_6881,N_6838);
or U7105 (N_7105,N_6993,N_6848);
nor U7106 (N_7106,N_6835,N_6816);
nor U7107 (N_7107,N_6941,N_6920);
or U7108 (N_7108,N_6961,N_6881);
nor U7109 (N_7109,N_6964,N_6942);
or U7110 (N_7110,N_6896,N_6873);
nand U7111 (N_7111,N_6966,N_6954);
or U7112 (N_7112,N_6921,N_6869);
nand U7113 (N_7113,N_6861,N_6813);
nor U7114 (N_7114,N_6841,N_6974);
nor U7115 (N_7115,N_6858,N_6817);
and U7116 (N_7116,N_6986,N_6954);
nor U7117 (N_7117,N_6971,N_6904);
or U7118 (N_7118,N_6864,N_6895);
and U7119 (N_7119,N_6943,N_6964);
nor U7120 (N_7120,N_6954,N_6806);
and U7121 (N_7121,N_6809,N_6968);
or U7122 (N_7122,N_6899,N_6862);
or U7123 (N_7123,N_6958,N_6878);
nand U7124 (N_7124,N_6895,N_6998);
nor U7125 (N_7125,N_6852,N_6952);
xnor U7126 (N_7126,N_6975,N_6866);
nand U7127 (N_7127,N_6816,N_6960);
and U7128 (N_7128,N_6889,N_6801);
nor U7129 (N_7129,N_6831,N_6877);
or U7130 (N_7130,N_6937,N_6973);
nand U7131 (N_7131,N_6923,N_6963);
nor U7132 (N_7132,N_6952,N_6863);
or U7133 (N_7133,N_6906,N_6988);
nor U7134 (N_7134,N_6885,N_6873);
or U7135 (N_7135,N_6892,N_6955);
nand U7136 (N_7136,N_6867,N_6955);
nand U7137 (N_7137,N_6997,N_6905);
and U7138 (N_7138,N_6879,N_6852);
or U7139 (N_7139,N_6960,N_6819);
nand U7140 (N_7140,N_6841,N_6928);
and U7141 (N_7141,N_6827,N_6932);
nand U7142 (N_7142,N_6945,N_6841);
nand U7143 (N_7143,N_6908,N_6848);
nor U7144 (N_7144,N_6926,N_6861);
xor U7145 (N_7145,N_6829,N_6990);
and U7146 (N_7146,N_6828,N_6947);
nor U7147 (N_7147,N_6849,N_6963);
nor U7148 (N_7148,N_6836,N_6964);
nand U7149 (N_7149,N_6924,N_6886);
nor U7150 (N_7150,N_6956,N_6899);
nor U7151 (N_7151,N_6877,N_6894);
and U7152 (N_7152,N_6847,N_6863);
nor U7153 (N_7153,N_6976,N_6905);
and U7154 (N_7154,N_6889,N_6966);
and U7155 (N_7155,N_6839,N_6878);
nor U7156 (N_7156,N_6939,N_6894);
and U7157 (N_7157,N_6805,N_6944);
or U7158 (N_7158,N_6904,N_6887);
or U7159 (N_7159,N_6816,N_6829);
nand U7160 (N_7160,N_6946,N_6917);
or U7161 (N_7161,N_6879,N_6923);
and U7162 (N_7162,N_6918,N_6849);
nand U7163 (N_7163,N_6804,N_6998);
nand U7164 (N_7164,N_6981,N_6861);
nand U7165 (N_7165,N_6855,N_6866);
nor U7166 (N_7166,N_6950,N_6863);
nor U7167 (N_7167,N_6820,N_6976);
nand U7168 (N_7168,N_6994,N_6995);
and U7169 (N_7169,N_6883,N_6988);
or U7170 (N_7170,N_6940,N_6854);
nand U7171 (N_7171,N_6904,N_6917);
and U7172 (N_7172,N_6898,N_6993);
and U7173 (N_7173,N_6968,N_6990);
or U7174 (N_7174,N_6932,N_6970);
nor U7175 (N_7175,N_6817,N_6856);
and U7176 (N_7176,N_6961,N_6832);
or U7177 (N_7177,N_6987,N_6981);
nor U7178 (N_7178,N_6830,N_6937);
nand U7179 (N_7179,N_6963,N_6941);
or U7180 (N_7180,N_6832,N_6835);
or U7181 (N_7181,N_6872,N_6917);
and U7182 (N_7182,N_6963,N_6888);
nor U7183 (N_7183,N_6891,N_6872);
xnor U7184 (N_7184,N_6929,N_6975);
or U7185 (N_7185,N_6920,N_6989);
and U7186 (N_7186,N_6841,N_6825);
or U7187 (N_7187,N_6923,N_6999);
and U7188 (N_7188,N_6857,N_6922);
nor U7189 (N_7189,N_6812,N_6899);
or U7190 (N_7190,N_6944,N_6893);
and U7191 (N_7191,N_6819,N_6854);
nor U7192 (N_7192,N_6954,N_6815);
nand U7193 (N_7193,N_6939,N_6840);
and U7194 (N_7194,N_6846,N_6801);
nand U7195 (N_7195,N_6803,N_6821);
nor U7196 (N_7196,N_6866,N_6999);
nor U7197 (N_7197,N_6858,N_6901);
and U7198 (N_7198,N_6872,N_6943);
nor U7199 (N_7199,N_6977,N_6959);
or U7200 (N_7200,N_7023,N_7131);
nor U7201 (N_7201,N_7024,N_7152);
or U7202 (N_7202,N_7027,N_7003);
and U7203 (N_7203,N_7187,N_7021);
or U7204 (N_7204,N_7054,N_7134);
nand U7205 (N_7205,N_7039,N_7140);
or U7206 (N_7206,N_7090,N_7053);
or U7207 (N_7207,N_7129,N_7035);
nor U7208 (N_7208,N_7103,N_7100);
nor U7209 (N_7209,N_7046,N_7083);
nand U7210 (N_7210,N_7040,N_7136);
nor U7211 (N_7211,N_7116,N_7061);
xor U7212 (N_7212,N_7169,N_7104);
or U7213 (N_7213,N_7171,N_7092);
and U7214 (N_7214,N_7042,N_7182);
and U7215 (N_7215,N_7001,N_7191);
or U7216 (N_7216,N_7009,N_7075);
and U7217 (N_7217,N_7007,N_7195);
nand U7218 (N_7218,N_7082,N_7148);
or U7219 (N_7219,N_7072,N_7161);
nand U7220 (N_7220,N_7055,N_7167);
or U7221 (N_7221,N_7133,N_7172);
and U7222 (N_7222,N_7034,N_7066);
and U7223 (N_7223,N_7177,N_7045);
nor U7224 (N_7224,N_7085,N_7000);
nand U7225 (N_7225,N_7178,N_7183);
nor U7226 (N_7226,N_7164,N_7163);
and U7227 (N_7227,N_7106,N_7097);
nor U7228 (N_7228,N_7196,N_7158);
or U7229 (N_7229,N_7173,N_7002);
nor U7230 (N_7230,N_7022,N_7105);
and U7231 (N_7231,N_7143,N_7049);
and U7232 (N_7232,N_7151,N_7154);
nand U7233 (N_7233,N_7036,N_7080);
or U7234 (N_7234,N_7010,N_7118);
nand U7235 (N_7235,N_7068,N_7110);
and U7236 (N_7236,N_7111,N_7101);
nand U7237 (N_7237,N_7168,N_7137);
nand U7238 (N_7238,N_7114,N_7056);
nand U7239 (N_7239,N_7032,N_7069);
nand U7240 (N_7240,N_7028,N_7044);
or U7241 (N_7241,N_7081,N_7165);
and U7242 (N_7242,N_7071,N_7155);
nand U7243 (N_7243,N_7125,N_7079);
and U7244 (N_7244,N_7124,N_7159);
nand U7245 (N_7245,N_7060,N_7199);
nor U7246 (N_7246,N_7098,N_7175);
nand U7247 (N_7247,N_7094,N_7025);
or U7248 (N_7248,N_7157,N_7166);
or U7249 (N_7249,N_7119,N_7073);
or U7250 (N_7250,N_7018,N_7139);
and U7251 (N_7251,N_7033,N_7058);
nand U7252 (N_7252,N_7070,N_7087);
or U7253 (N_7253,N_7038,N_7099);
nor U7254 (N_7254,N_7005,N_7051);
or U7255 (N_7255,N_7150,N_7128);
nor U7256 (N_7256,N_7186,N_7095);
and U7257 (N_7257,N_7108,N_7180);
nand U7258 (N_7258,N_7029,N_7126);
nor U7259 (N_7259,N_7144,N_7138);
nor U7260 (N_7260,N_7076,N_7188);
nand U7261 (N_7261,N_7016,N_7189);
nor U7262 (N_7262,N_7050,N_7153);
nor U7263 (N_7263,N_7123,N_7011);
nor U7264 (N_7264,N_7062,N_7047);
nor U7265 (N_7265,N_7113,N_7193);
nand U7266 (N_7266,N_7088,N_7091);
nand U7267 (N_7267,N_7181,N_7135);
or U7268 (N_7268,N_7160,N_7077);
and U7269 (N_7269,N_7145,N_7015);
nand U7270 (N_7270,N_7086,N_7043);
nor U7271 (N_7271,N_7176,N_7030);
nand U7272 (N_7272,N_7074,N_7026);
and U7273 (N_7273,N_7109,N_7115);
or U7274 (N_7274,N_7146,N_7141);
and U7275 (N_7275,N_7078,N_7102);
nor U7276 (N_7276,N_7052,N_7020);
and U7277 (N_7277,N_7194,N_7048);
nand U7278 (N_7278,N_7093,N_7008);
and U7279 (N_7279,N_7065,N_7122);
nor U7280 (N_7280,N_7184,N_7179);
nor U7281 (N_7281,N_7012,N_7156);
nor U7282 (N_7282,N_7147,N_7006);
nor U7283 (N_7283,N_7132,N_7198);
nand U7284 (N_7284,N_7031,N_7014);
nor U7285 (N_7285,N_7057,N_7013);
nand U7286 (N_7286,N_7121,N_7084);
or U7287 (N_7287,N_7089,N_7174);
or U7288 (N_7288,N_7037,N_7107);
nand U7289 (N_7289,N_7117,N_7130);
nor U7290 (N_7290,N_7192,N_7017);
and U7291 (N_7291,N_7120,N_7096);
nor U7292 (N_7292,N_7127,N_7197);
nor U7293 (N_7293,N_7190,N_7162);
nor U7294 (N_7294,N_7142,N_7041);
nor U7295 (N_7295,N_7059,N_7063);
and U7296 (N_7296,N_7112,N_7004);
nor U7297 (N_7297,N_7185,N_7019);
nand U7298 (N_7298,N_7064,N_7149);
nor U7299 (N_7299,N_7170,N_7067);
and U7300 (N_7300,N_7183,N_7194);
and U7301 (N_7301,N_7107,N_7138);
nand U7302 (N_7302,N_7094,N_7033);
or U7303 (N_7303,N_7176,N_7186);
and U7304 (N_7304,N_7135,N_7121);
and U7305 (N_7305,N_7092,N_7087);
nand U7306 (N_7306,N_7046,N_7106);
or U7307 (N_7307,N_7143,N_7034);
or U7308 (N_7308,N_7132,N_7056);
nand U7309 (N_7309,N_7081,N_7036);
or U7310 (N_7310,N_7184,N_7059);
nor U7311 (N_7311,N_7155,N_7070);
and U7312 (N_7312,N_7020,N_7028);
nand U7313 (N_7313,N_7129,N_7037);
or U7314 (N_7314,N_7100,N_7166);
nand U7315 (N_7315,N_7068,N_7132);
or U7316 (N_7316,N_7078,N_7179);
or U7317 (N_7317,N_7051,N_7179);
and U7318 (N_7318,N_7157,N_7149);
nor U7319 (N_7319,N_7018,N_7036);
or U7320 (N_7320,N_7089,N_7048);
nand U7321 (N_7321,N_7056,N_7010);
or U7322 (N_7322,N_7017,N_7001);
nor U7323 (N_7323,N_7139,N_7090);
or U7324 (N_7324,N_7175,N_7047);
or U7325 (N_7325,N_7022,N_7120);
nand U7326 (N_7326,N_7055,N_7146);
nor U7327 (N_7327,N_7182,N_7129);
nor U7328 (N_7328,N_7005,N_7032);
or U7329 (N_7329,N_7173,N_7028);
and U7330 (N_7330,N_7116,N_7146);
nor U7331 (N_7331,N_7128,N_7007);
and U7332 (N_7332,N_7142,N_7003);
and U7333 (N_7333,N_7012,N_7031);
nand U7334 (N_7334,N_7081,N_7005);
and U7335 (N_7335,N_7022,N_7198);
and U7336 (N_7336,N_7139,N_7030);
and U7337 (N_7337,N_7077,N_7122);
nor U7338 (N_7338,N_7112,N_7045);
nand U7339 (N_7339,N_7088,N_7052);
nand U7340 (N_7340,N_7099,N_7137);
nand U7341 (N_7341,N_7015,N_7053);
nand U7342 (N_7342,N_7090,N_7199);
nor U7343 (N_7343,N_7177,N_7187);
or U7344 (N_7344,N_7020,N_7129);
or U7345 (N_7345,N_7087,N_7160);
and U7346 (N_7346,N_7082,N_7109);
nor U7347 (N_7347,N_7109,N_7005);
nand U7348 (N_7348,N_7088,N_7032);
or U7349 (N_7349,N_7170,N_7053);
or U7350 (N_7350,N_7167,N_7114);
nor U7351 (N_7351,N_7149,N_7084);
and U7352 (N_7352,N_7090,N_7192);
and U7353 (N_7353,N_7097,N_7073);
or U7354 (N_7354,N_7111,N_7029);
nor U7355 (N_7355,N_7182,N_7141);
nor U7356 (N_7356,N_7049,N_7196);
nand U7357 (N_7357,N_7143,N_7094);
nor U7358 (N_7358,N_7166,N_7168);
and U7359 (N_7359,N_7064,N_7105);
or U7360 (N_7360,N_7154,N_7085);
and U7361 (N_7361,N_7148,N_7150);
nand U7362 (N_7362,N_7135,N_7093);
and U7363 (N_7363,N_7123,N_7078);
or U7364 (N_7364,N_7040,N_7052);
or U7365 (N_7365,N_7098,N_7150);
nor U7366 (N_7366,N_7063,N_7049);
nand U7367 (N_7367,N_7048,N_7138);
or U7368 (N_7368,N_7052,N_7050);
nand U7369 (N_7369,N_7156,N_7086);
or U7370 (N_7370,N_7084,N_7193);
and U7371 (N_7371,N_7023,N_7085);
and U7372 (N_7372,N_7097,N_7153);
and U7373 (N_7373,N_7119,N_7105);
or U7374 (N_7374,N_7123,N_7182);
nor U7375 (N_7375,N_7159,N_7025);
and U7376 (N_7376,N_7194,N_7147);
nand U7377 (N_7377,N_7020,N_7035);
or U7378 (N_7378,N_7168,N_7053);
nor U7379 (N_7379,N_7154,N_7136);
or U7380 (N_7380,N_7143,N_7142);
nor U7381 (N_7381,N_7069,N_7063);
nand U7382 (N_7382,N_7027,N_7092);
nand U7383 (N_7383,N_7129,N_7030);
nor U7384 (N_7384,N_7152,N_7022);
nand U7385 (N_7385,N_7120,N_7054);
and U7386 (N_7386,N_7008,N_7014);
nor U7387 (N_7387,N_7195,N_7171);
nand U7388 (N_7388,N_7135,N_7038);
or U7389 (N_7389,N_7067,N_7016);
nor U7390 (N_7390,N_7017,N_7129);
and U7391 (N_7391,N_7065,N_7184);
and U7392 (N_7392,N_7018,N_7035);
nand U7393 (N_7393,N_7001,N_7030);
nor U7394 (N_7394,N_7029,N_7086);
and U7395 (N_7395,N_7105,N_7140);
nand U7396 (N_7396,N_7172,N_7135);
nand U7397 (N_7397,N_7090,N_7029);
and U7398 (N_7398,N_7103,N_7089);
nor U7399 (N_7399,N_7089,N_7043);
nor U7400 (N_7400,N_7326,N_7394);
or U7401 (N_7401,N_7387,N_7242);
nand U7402 (N_7402,N_7249,N_7232);
or U7403 (N_7403,N_7360,N_7369);
nor U7404 (N_7404,N_7372,N_7377);
nand U7405 (N_7405,N_7207,N_7314);
and U7406 (N_7406,N_7382,N_7215);
nor U7407 (N_7407,N_7296,N_7307);
or U7408 (N_7408,N_7254,N_7252);
nor U7409 (N_7409,N_7333,N_7264);
and U7410 (N_7410,N_7325,N_7288);
or U7411 (N_7411,N_7376,N_7388);
nand U7412 (N_7412,N_7223,N_7362);
and U7413 (N_7413,N_7346,N_7344);
nor U7414 (N_7414,N_7374,N_7313);
and U7415 (N_7415,N_7238,N_7361);
nor U7416 (N_7416,N_7319,N_7318);
and U7417 (N_7417,N_7340,N_7265);
nor U7418 (N_7418,N_7277,N_7371);
nand U7419 (N_7419,N_7272,N_7304);
or U7420 (N_7420,N_7251,N_7363);
nor U7421 (N_7421,N_7225,N_7329);
and U7422 (N_7422,N_7308,N_7285);
nor U7423 (N_7423,N_7389,N_7212);
and U7424 (N_7424,N_7200,N_7391);
nor U7425 (N_7425,N_7298,N_7347);
nand U7426 (N_7426,N_7204,N_7399);
and U7427 (N_7427,N_7324,N_7213);
nor U7428 (N_7428,N_7332,N_7381);
and U7429 (N_7429,N_7370,N_7306);
and U7430 (N_7430,N_7257,N_7209);
nor U7431 (N_7431,N_7261,N_7241);
or U7432 (N_7432,N_7276,N_7226);
and U7433 (N_7433,N_7393,N_7357);
and U7434 (N_7434,N_7323,N_7219);
nand U7435 (N_7435,N_7202,N_7275);
and U7436 (N_7436,N_7355,N_7274);
or U7437 (N_7437,N_7284,N_7309);
and U7438 (N_7438,N_7224,N_7293);
nand U7439 (N_7439,N_7300,N_7231);
nor U7440 (N_7440,N_7336,N_7310);
nor U7441 (N_7441,N_7216,N_7237);
and U7442 (N_7442,N_7305,N_7273);
or U7443 (N_7443,N_7262,N_7246);
or U7444 (N_7444,N_7235,N_7348);
or U7445 (N_7445,N_7217,N_7255);
and U7446 (N_7446,N_7337,N_7349);
nand U7447 (N_7447,N_7342,N_7328);
xor U7448 (N_7448,N_7270,N_7205);
xor U7449 (N_7449,N_7398,N_7201);
nand U7450 (N_7450,N_7343,N_7208);
nand U7451 (N_7451,N_7334,N_7367);
nand U7452 (N_7452,N_7203,N_7320);
nand U7453 (N_7453,N_7383,N_7373);
or U7454 (N_7454,N_7244,N_7230);
and U7455 (N_7455,N_7206,N_7247);
nor U7456 (N_7456,N_7335,N_7386);
or U7457 (N_7457,N_7365,N_7339);
or U7458 (N_7458,N_7259,N_7236);
and U7459 (N_7459,N_7256,N_7283);
nor U7460 (N_7460,N_7303,N_7248);
xor U7461 (N_7461,N_7282,N_7280);
nand U7462 (N_7462,N_7295,N_7227);
nand U7463 (N_7463,N_7375,N_7287);
or U7464 (N_7464,N_7358,N_7297);
and U7465 (N_7465,N_7354,N_7253);
nor U7466 (N_7466,N_7292,N_7239);
nor U7467 (N_7467,N_7240,N_7350);
and U7468 (N_7468,N_7327,N_7353);
or U7469 (N_7469,N_7301,N_7245);
nor U7470 (N_7470,N_7384,N_7214);
or U7471 (N_7471,N_7281,N_7299);
nor U7472 (N_7472,N_7243,N_7211);
nand U7473 (N_7473,N_7315,N_7289);
nor U7474 (N_7474,N_7218,N_7278);
or U7475 (N_7475,N_7392,N_7379);
or U7476 (N_7476,N_7390,N_7351);
nor U7477 (N_7477,N_7368,N_7222);
or U7478 (N_7478,N_7229,N_7356);
and U7479 (N_7479,N_7258,N_7341);
nand U7480 (N_7480,N_7359,N_7271);
or U7481 (N_7481,N_7220,N_7263);
or U7482 (N_7482,N_7250,N_7378);
nand U7483 (N_7483,N_7228,N_7279);
nand U7484 (N_7484,N_7345,N_7366);
and U7485 (N_7485,N_7396,N_7302);
nor U7486 (N_7486,N_7269,N_7268);
and U7487 (N_7487,N_7352,N_7294);
nor U7488 (N_7488,N_7291,N_7322);
nor U7489 (N_7489,N_7317,N_7260);
or U7490 (N_7490,N_7395,N_7210);
nand U7491 (N_7491,N_7221,N_7266);
nand U7492 (N_7492,N_7330,N_7331);
or U7493 (N_7493,N_7380,N_7338);
or U7494 (N_7494,N_7286,N_7234);
nor U7495 (N_7495,N_7385,N_7290);
and U7496 (N_7496,N_7311,N_7312);
nand U7497 (N_7497,N_7321,N_7316);
or U7498 (N_7498,N_7233,N_7267);
nand U7499 (N_7499,N_7397,N_7364);
and U7500 (N_7500,N_7278,N_7213);
nand U7501 (N_7501,N_7276,N_7295);
nand U7502 (N_7502,N_7325,N_7207);
nand U7503 (N_7503,N_7250,N_7266);
or U7504 (N_7504,N_7214,N_7341);
nor U7505 (N_7505,N_7221,N_7359);
nor U7506 (N_7506,N_7235,N_7265);
and U7507 (N_7507,N_7352,N_7358);
or U7508 (N_7508,N_7292,N_7373);
and U7509 (N_7509,N_7367,N_7264);
nor U7510 (N_7510,N_7298,N_7207);
or U7511 (N_7511,N_7365,N_7286);
or U7512 (N_7512,N_7377,N_7242);
nand U7513 (N_7513,N_7333,N_7316);
or U7514 (N_7514,N_7278,N_7237);
or U7515 (N_7515,N_7294,N_7206);
nor U7516 (N_7516,N_7269,N_7267);
nand U7517 (N_7517,N_7252,N_7234);
nand U7518 (N_7518,N_7343,N_7217);
nor U7519 (N_7519,N_7262,N_7237);
or U7520 (N_7520,N_7360,N_7294);
and U7521 (N_7521,N_7286,N_7227);
nand U7522 (N_7522,N_7280,N_7247);
nor U7523 (N_7523,N_7279,N_7277);
nor U7524 (N_7524,N_7268,N_7211);
or U7525 (N_7525,N_7341,N_7324);
nor U7526 (N_7526,N_7376,N_7259);
nand U7527 (N_7527,N_7260,N_7237);
or U7528 (N_7528,N_7279,N_7338);
or U7529 (N_7529,N_7372,N_7295);
and U7530 (N_7530,N_7397,N_7242);
or U7531 (N_7531,N_7353,N_7269);
or U7532 (N_7532,N_7326,N_7279);
and U7533 (N_7533,N_7319,N_7362);
and U7534 (N_7534,N_7244,N_7387);
and U7535 (N_7535,N_7397,N_7391);
nand U7536 (N_7536,N_7318,N_7367);
or U7537 (N_7537,N_7268,N_7201);
or U7538 (N_7538,N_7298,N_7357);
or U7539 (N_7539,N_7390,N_7363);
nand U7540 (N_7540,N_7364,N_7353);
and U7541 (N_7541,N_7336,N_7239);
nand U7542 (N_7542,N_7265,N_7207);
or U7543 (N_7543,N_7387,N_7382);
nor U7544 (N_7544,N_7218,N_7299);
and U7545 (N_7545,N_7372,N_7299);
or U7546 (N_7546,N_7387,N_7202);
nand U7547 (N_7547,N_7311,N_7204);
or U7548 (N_7548,N_7315,N_7243);
nor U7549 (N_7549,N_7376,N_7370);
nand U7550 (N_7550,N_7315,N_7390);
and U7551 (N_7551,N_7330,N_7367);
or U7552 (N_7552,N_7254,N_7242);
nand U7553 (N_7553,N_7237,N_7316);
nor U7554 (N_7554,N_7348,N_7332);
or U7555 (N_7555,N_7220,N_7361);
and U7556 (N_7556,N_7256,N_7270);
nor U7557 (N_7557,N_7330,N_7372);
nand U7558 (N_7558,N_7326,N_7253);
nand U7559 (N_7559,N_7278,N_7238);
and U7560 (N_7560,N_7241,N_7284);
or U7561 (N_7561,N_7370,N_7372);
xor U7562 (N_7562,N_7341,N_7270);
and U7563 (N_7563,N_7323,N_7383);
and U7564 (N_7564,N_7226,N_7385);
nand U7565 (N_7565,N_7248,N_7395);
nor U7566 (N_7566,N_7362,N_7316);
or U7567 (N_7567,N_7375,N_7278);
nor U7568 (N_7568,N_7340,N_7363);
or U7569 (N_7569,N_7364,N_7235);
nor U7570 (N_7570,N_7379,N_7294);
nor U7571 (N_7571,N_7281,N_7218);
and U7572 (N_7572,N_7398,N_7246);
and U7573 (N_7573,N_7338,N_7225);
and U7574 (N_7574,N_7378,N_7320);
or U7575 (N_7575,N_7300,N_7245);
and U7576 (N_7576,N_7355,N_7290);
nor U7577 (N_7577,N_7321,N_7314);
or U7578 (N_7578,N_7271,N_7376);
nand U7579 (N_7579,N_7352,N_7374);
and U7580 (N_7580,N_7338,N_7200);
or U7581 (N_7581,N_7218,N_7340);
nor U7582 (N_7582,N_7263,N_7323);
or U7583 (N_7583,N_7311,N_7258);
nand U7584 (N_7584,N_7368,N_7201);
xor U7585 (N_7585,N_7317,N_7393);
nor U7586 (N_7586,N_7266,N_7214);
nand U7587 (N_7587,N_7300,N_7368);
and U7588 (N_7588,N_7222,N_7330);
nand U7589 (N_7589,N_7294,N_7295);
nand U7590 (N_7590,N_7396,N_7376);
or U7591 (N_7591,N_7294,N_7345);
and U7592 (N_7592,N_7310,N_7219);
nand U7593 (N_7593,N_7234,N_7290);
and U7594 (N_7594,N_7259,N_7226);
nand U7595 (N_7595,N_7250,N_7206);
nor U7596 (N_7596,N_7237,N_7259);
nor U7597 (N_7597,N_7354,N_7297);
nor U7598 (N_7598,N_7369,N_7215);
or U7599 (N_7599,N_7397,N_7367);
and U7600 (N_7600,N_7486,N_7577);
or U7601 (N_7601,N_7497,N_7401);
nand U7602 (N_7602,N_7570,N_7458);
or U7603 (N_7603,N_7503,N_7528);
nor U7604 (N_7604,N_7452,N_7477);
or U7605 (N_7605,N_7546,N_7468);
nand U7606 (N_7606,N_7408,N_7413);
or U7607 (N_7607,N_7469,N_7502);
nor U7608 (N_7608,N_7586,N_7563);
or U7609 (N_7609,N_7549,N_7485);
or U7610 (N_7610,N_7424,N_7463);
nor U7611 (N_7611,N_7566,N_7567);
nor U7612 (N_7612,N_7512,N_7533);
and U7613 (N_7613,N_7431,N_7561);
and U7614 (N_7614,N_7499,N_7482);
nor U7615 (N_7615,N_7474,N_7456);
nor U7616 (N_7616,N_7545,N_7592);
nand U7617 (N_7617,N_7415,N_7419);
nor U7618 (N_7618,N_7564,N_7483);
and U7619 (N_7619,N_7501,N_7529);
nand U7620 (N_7620,N_7426,N_7535);
and U7621 (N_7621,N_7557,N_7476);
or U7622 (N_7622,N_7583,N_7581);
nand U7623 (N_7623,N_7520,N_7542);
nand U7624 (N_7624,N_7446,N_7444);
nand U7625 (N_7625,N_7425,N_7489);
or U7626 (N_7626,N_7422,N_7579);
or U7627 (N_7627,N_7505,N_7437);
and U7628 (N_7628,N_7587,N_7578);
nand U7629 (N_7629,N_7438,N_7596);
nor U7630 (N_7630,N_7466,N_7461);
and U7631 (N_7631,N_7550,N_7400);
nand U7632 (N_7632,N_7462,N_7460);
and U7633 (N_7633,N_7555,N_7434);
and U7634 (N_7634,N_7481,N_7598);
and U7635 (N_7635,N_7548,N_7538);
nor U7636 (N_7636,N_7500,N_7417);
and U7637 (N_7637,N_7451,N_7521);
nand U7638 (N_7638,N_7543,N_7591);
or U7639 (N_7639,N_7589,N_7580);
nand U7640 (N_7640,N_7436,N_7506);
nor U7641 (N_7641,N_7547,N_7588);
or U7642 (N_7642,N_7585,N_7552);
nor U7643 (N_7643,N_7433,N_7554);
nand U7644 (N_7644,N_7492,N_7490);
nor U7645 (N_7645,N_7559,N_7459);
or U7646 (N_7646,N_7590,N_7568);
nor U7647 (N_7647,N_7488,N_7423);
or U7648 (N_7648,N_7487,N_7510);
or U7649 (N_7649,N_7407,N_7455);
nor U7650 (N_7650,N_7525,N_7551);
or U7651 (N_7651,N_7507,N_7475);
nor U7652 (N_7652,N_7553,N_7498);
nand U7653 (N_7653,N_7522,N_7516);
and U7654 (N_7654,N_7448,N_7519);
or U7655 (N_7655,N_7427,N_7571);
nand U7656 (N_7656,N_7471,N_7560);
nor U7657 (N_7657,N_7439,N_7402);
or U7658 (N_7658,N_7403,N_7409);
and U7659 (N_7659,N_7479,N_7411);
or U7660 (N_7660,N_7514,N_7518);
and U7661 (N_7661,N_7504,N_7532);
and U7662 (N_7662,N_7428,N_7541);
nand U7663 (N_7663,N_7450,N_7530);
nor U7664 (N_7664,N_7430,N_7496);
nor U7665 (N_7665,N_7406,N_7562);
nand U7666 (N_7666,N_7465,N_7416);
and U7667 (N_7667,N_7405,N_7464);
nand U7668 (N_7668,N_7457,N_7443);
or U7669 (N_7669,N_7597,N_7447);
nor U7670 (N_7670,N_7491,N_7593);
and U7671 (N_7671,N_7582,N_7495);
and U7672 (N_7672,N_7435,N_7404);
or U7673 (N_7673,N_7454,N_7537);
nor U7674 (N_7674,N_7429,N_7515);
nor U7675 (N_7675,N_7412,N_7418);
nor U7676 (N_7676,N_7575,N_7565);
nand U7677 (N_7677,N_7572,N_7467);
and U7678 (N_7678,N_7540,N_7576);
or U7679 (N_7679,N_7494,N_7453);
nand U7680 (N_7680,N_7484,N_7445);
and U7681 (N_7681,N_7573,N_7524);
or U7682 (N_7682,N_7508,N_7556);
nand U7683 (N_7683,N_7594,N_7513);
nor U7684 (N_7684,N_7569,N_7478);
and U7685 (N_7685,N_7511,N_7472);
nor U7686 (N_7686,N_7526,N_7574);
nand U7687 (N_7687,N_7531,N_7440);
or U7688 (N_7688,N_7473,N_7595);
or U7689 (N_7689,N_7527,N_7432);
or U7690 (N_7690,N_7517,N_7449);
and U7691 (N_7691,N_7480,N_7539);
nor U7692 (N_7692,N_7509,N_7414);
nor U7693 (N_7693,N_7470,N_7599);
and U7694 (N_7694,N_7536,N_7544);
nor U7695 (N_7695,N_7442,N_7410);
and U7696 (N_7696,N_7420,N_7584);
nand U7697 (N_7697,N_7534,N_7493);
and U7698 (N_7698,N_7421,N_7523);
or U7699 (N_7699,N_7558,N_7441);
or U7700 (N_7700,N_7592,N_7591);
or U7701 (N_7701,N_7446,N_7418);
or U7702 (N_7702,N_7481,N_7483);
nor U7703 (N_7703,N_7565,N_7496);
or U7704 (N_7704,N_7504,N_7476);
and U7705 (N_7705,N_7425,N_7411);
nor U7706 (N_7706,N_7417,N_7482);
or U7707 (N_7707,N_7437,N_7522);
and U7708 (N_7708,N_7454,N_7522);
nor U7709 (N_7709,N_7579,N_7429);
nand U7710 (N_7710,N_7462,N_7530);
nor U7711 (N_7711,N_7541,N_7513);
and U7712 (N_7712,N_7473,N_7578);
or U7713 (N_7713,N_7436,N_7431);
or U7714 (N_7714,N_7429,N_7566);
or U7715 (N_7715,N_7453,N_7407);
nand U7716 (N_7716,N_7453,N_7479);
and U7717 (N_7717,N_7408,N_7541);
or U7718 (N_7718,N_7425,N_7541);
and U7719 (N_7719,N_7401,N_7588);
nand U7720 (N_7720,N_7505,N_7576);
and U7721 (N_7721,N_7588,N_7437);
or U7722 (N_7722,N_7501,N_7425);
nor U7723 (N_7723,N_7519,N_7442);
or U7724 (N_7724,N_7483,N_7494);
nand U7725 (N_7725,N_7578,N_7478);
nand U7726 (N_7726,N_7424,N_7416);
and U7727 (N_7727,N_7528,N_7404);
or U7728 (N_7728,N_7478,N_7448);
nor U7729 (N_7729,N_7506,N_7431);
nand U7730 (N_7730,N_7520,N_7468);
nor U7731 (N_7731,N_7537,N_7402);
nor U7732 (N_7732,N_7418,N_7421);
and U7733 (N_7733,N_7416,N_7420);
nor U7734 (N_7734,N_7598,N_7574);
or U7735 (N_7735,N_7532,N_7401);
nor U7736 (N_7736,N_7410,N_7583);
and U7737 (N_7737,N_7523,N_7534);
and U7738 (N_7738,N_7481,N_7452);
and U7739 (N_7739,N_7511,N_7477);
or U7740 (N_7740,N_7405,N_7411);
and U7741 (N_7741,N_7545,N_7495);
nand U7742 (N_7742,N_7424,N_7467);
or U7743 (N_7743,N_7573,N_7527);
nor U7744 (N_7744,N_7548,N_7488);
nand U7745 (N_7745,N_7553,N_7468);
nor U7746 (N_7746,N_7469,N_7404);
nor U7747 (N_7747,N_7549,N_7518);
nor U7748 (N_7748,N_7508,N_7518);
nand U7749 (N_7749,N_7527,N_7468);
and U7750 (N_7750,N_7402,N_7425);
nor U7751 (N_7751,N_7447,N_7598);
and U7752 (N_7752,N_7485,N_7502);
nand U7753 (N_7753,N_7504,N_7419);
xnor U7754 (N_7754,N_7425,N_7518);
nor U7755 (N_7755,N_7475,N_7468);
or U7756 (N_7756,N_7564,N_7496);
nand U7757 (N_7757,N_7437,N_7465);
nor U7758 (N_7758,N_7524,N_7579);
nand U7759 (N_7759,N_7535,N_7446);
nor U7760 (N_7760,N_7512,N_7401);
and U7761 (N_7761,N_7442,N_7421);
or U7762 (N_7762,N_7503,N_7499);
nor U7763 (N_7763,N_7466,N_7584);
nor U7764 (N_7764,N_7435,N_7462);
or U7765 (N_7765,N_7534,N_7526);
and U7766 (N_7766,N_7498,N_7583);
nand U7767 (N_7767,N_7405,N_7467);
or U7768 (N_7768,N_7414,N_7561);
and U7769 (N_7769,N_7404,N_7448);
and U7770 (N_7770,N_7568,N_7548);
or U7771 (N_7771,N_7554,N_7461);
and U7772 (N_7772,N_7596,N_7490);
and U7773 (N_7773,N_7437,N_7547);
or U7774 (N_7774,N_7449,N_7558);
or U7775 (N_7775,N_7492,N_7450);
and U7776 (N_7776,N_7574,N_7502);
and U7777 (N_7777,N_7516,N_7509);
nor U7778 (N_7778,N_7572,N_7531);
nand U7779 (N_7779,N_7469,N_7506);
and U7780 (N_7780,N_7511,N_7543);
nor U7781 (N_7781,N_7551,N_7587);
nand U7782 (N_7782,N_7536,N_7579);
nor U7783 (N_7783,N_7422,N_7566);
nor U7784 (N_7784,N_7484,N_7426);
nor U7785 (N_7785,N_7417,N_7509);
nor U7786 (N_7786,N_7423,N_7464);
nand U7787 (N_7787,N_7524,N_7590);
and U7788 (N_7788,N_7412,N_7441);
nor U7789 (N_7789,N_7435,N_7436);
and U7790 (N_7790,N_7450,N_7582);
nor U7791 (N_7791,N_7556,N_7474);
or U7792 (N_7792,N_7453,N_7518);
nor U7793 (N_7793,N_7498,N_7588);
and U7794 (N_7794,N_7565,N_7459);
and U7795 (N_7795,N_7445,N_7572);
or U7796 (N_7796,N_7569,N_7517);
and U7797 (N_7797,N_7563,N_7465);
nor U7798 (N_7798,N_7594,N_7527);
and U7799 (N_7799,N_7574,N_7463);
or U7800 (N_7800,N_7700,N_7631);
and U7801 (N_7801,N_7722,N_7784);
nor U7802 (N_7802,N_7701,N_7602);
or U7803 (N_7803,N_7698,N_7629);
nor U7804 (N_7804,N_7619,N_7720);
or U7805 (N_7805,N_7751,N_7643);
nand U7806 (N_7806,N_7793,N_7735);
or U7807 (N_7807,N_7750,N_7748);
and U7808 (N_7808,N_7713,N_7708);
nand U7809 (N_7809,N_7678,N_7755);
nand U7810 (N_7810,N_7795,N_7799);
nand U7811 (N_7811,N_7703,N_7622);
nor U7812 (N_7812,N_7661,N_7646);
nand U7813 (N_7813,N_7625,N_7611);
nand U7814 (N_7814,N_7760,N_7671);
or U7815 (N_7815,N_7762,N_7758);
nand U7816 (N_7816,N_7695,N_7742);
nor U7817 (N_7817,N_7604,N_7741);
or U7818 (N_7818,N_7680,N_7617);
nand U7819 (N_7819,N_7718,N_7716);
nor U7820 (N_7820,N_7667,N_7739);
or U7821 (N_7821,N_7753,N_7668);
nor U7822 (N_7822,N_7651,N_7712);
and U7823 (N_7823,N_7771,N_7664);
nor U7824 (N_7824,N_7687,N_7707);
and U7825 (N_7825,N_7609,N_7724);
nand U7826 (N_7826,N_7696,N_7785);
nand U7827 (N_7827,N_7675,N_7764);
nor U7828 (N_7828,N_7647,N_7615);
nand U7829 (N_7829,N_7699,N_7770);
and U7830 (N_7830,N_7613,N_7705);
nor U7831 (N_7831,N_7607,N_7662);
nor U7832 (N_7832,N_7706,N_7633);
nand U7833 (N_7833,N_7688,N_7736);
nor U7834 (N_7834,N_7682,N_7768);
nand U7835 (N_7835,N_7640,N_7723);
nand U7836 (N_7836,N_7610,N_7637);
nand U7837 (N_7837,N_7690,N_7686);
or U7838 (N_7838,N_7636,N_7632);
or U7839 (N_7839,N_7623,N_7654);
or U7840 (N_7840,N_7618,N_7694);
or U7841 (N_7841,N_7757,N_7674);
nand U7842 (N_7842,N_7670,N_7666);
nor U7843 (N_7843,N_7780,N_7660);
nand U7844 (N_7844,N_7756,N_7676);
and U7845 (N_7845,N_7797,N_7638);
nor U7846 (N_7846,N_7767,N_7601);
or U7847 (N_7847,N_7774,N_7710);
nor U7848 (N_7848,N_7624,N_7659);
or U7849 (N_7849,N_7728,N_7792);
and U7850 (N_7850,N_7752,N_7776);
nand U7851 (N_7851,N_7684,N_7681);
nor U7852 (N_7852,N_7616,N_7693);
and U7853 (N_7853,N_7778,N_7691);
and U7854 (N_7854,N_7653,N_7747);
or U7855 (N_7855,N_7635,N_7772);
nand U7856 (N_7856,N_7605,N_7765);
or U7857 (N_7857,N_7683,N_7650);
or U7858 (N_7858,N_7642,N_7692);
nor U7859 (N_7859,N_7763,N_7652);
and U7860 (N_7860,N_7773,N_7743);
or U7861 (N_7861,N_7759,N_7738);
nor U7862 (N_7862,N_7733,N_7769);
or U7863 (N_7863,N_7714,N_7794);
nor U7864 (N_7864,N_7641,N_7737);
xor U7865 (N_7865,N_7783,N_7775);
nand U7866 (N_7866,N_7761,N_7719);
nand U7867 (N_7867,N_7614,N_7726);
nand U7868 (N_7868,N_7709,N_7704);
nor U7869 (N_7869,N_7730,N_7777);
nor U7870 (N_7870,N_7685,N_7679);
nor U7871 (N_7871,N_7620,N_7717);
nand U7872 (N_7872,N_7630,N_7621);
nor U7873 (N_7873,N_7702,N_7665);
nand U7874 (N_7874,N_7645,N_7786);
nor U7875 (N_7875,N_7790,N_7721);
and U7876 (N_7876,N_7608,N_7612);
nor U7877 (N_7877,N_7663,N_7689);
nand U7878 (N_7878,N_7725,N_7600);
or U7879 (N_7879,N_7796,N_7649);
and U7880 (N_7880,N_7672,N_7627);
nand U7881 (N_7881,N_7673,N_7791);
nand U7882 (N_7882,N_7658,N_7788);
and U7883 (N_7883,N_7669,N_7731);
nor U7884 (N_7884,N_7603,N_7729);
or U7885 (N_7885,N_7639,N_7744);
or U7886 (N_7886,N_7740,N_7734);
and U7887 (N_7887,N_7657,N_7732);
and U7888 (N_7888,N_7606,N_7781);
nor U7889 (N_7889,N_7754,N_7779);
or U7890 (N_7890,N_7766,N_7749);
and U7891 (N_7891,N_7626,N_7746);
nand U7892 (N_7892,N_7711,N_7745);
or U7893 (N_7893,N_7787,N_7782);
nand U7894 (N_7894,N_7634,N_7628);
nor U7895 (N_7895,N_7798,N_7648);
or U7896 (N_7896,N_7715,N_7656);
or U7897 (N_7897,N_7677,N_7655);
and U7898 (N_7898,N_7644,N_7789);
or U7899 (N_7899,N_7697,N_7727);
nand U7900 (N_7900,N_7711,N_7798);
or U7901 (N_7901,N_7664,N_7761);
nor U7902 (N_7902,N_7779,N_7766);
or U7903 (N_7903,N_7734,N_7790);
and U7904 (N_7904,N_7781,N_7696);
nand U7905 (N_7905,N_7651,N_7726);
xor U7906 (N_7906,N_7714,N_7730);
or U7907 (N_7907,N_7628,N_7603);
nor U7908 (N_7908,N_7765,N_7674);
nand U7909 (N_7909,N_7756,N_7648);
or U7910 (N_7910,N_7741,N_7763);
nand U7911 (N_7911,N_7615,N_7750);
or U7912 (N_7912,N_7707,N_7787);
nand U7913 (N_7913,N_7606,N_7682);
nand U7914 (N_7914,N_7710,N_7694);
or U7915 (N_7915,N_7771,N_7704);
nand U7916 (N_7916,N_7642,N_7633);
or U7917 (N_7917,N_7793,N_7750);
and U7918 (N_7918,N_7796,N_7638);
and U7919 (N_7919,N_7682,N_7787);
nor U7920 (N_7920,N_7642,N_7632);
nand U7921 (N_7921,N_7729,N_7616);
nor U7922 (N_7922,N_7769,N_7632);
nor U7923 (N_7923,N_7642,N_7766);
nand U7924 (N_7924,N_7703,N_7623);
nor U7925 (N_7925,N_7765,N_7708);
nand U7926 (N_7926,N_7729,N_7618);
nand U7927 (N_7927,N_7622,N_7656);
nand U7928 (N_7928,N_7645,N_7704);
nor U7929 (N_7929,N_7773,N_7690);
nand U7930 (N_7930,N_7722,N_7675);
nand U7931 (N_7931,N_7607,N_7720);
nand U7932 (N_7932,N_7738,N_7723);
and U7933 (N_7933,N_7634,N_7697);
or U7934 (N_7934,N_7760,N_7704);
nand U7935 (N_7935,N_7705,N_7694);
or U7936 (N_7936,N_7747,N_7770);
nand U7937 (N_7937,N_7689,N_7679);
nor U7938 (N_7938,N_7792,N_7651);
nor U7939 (N_7939,N_7758,N_7702);
nand U7940 (N_7940,N_7708,N_7679);
nor U7941 (N_7941,N_7673,N_7720);
and U7942 (N_7942,N_7660,N_7622);
nand U7943 (N_7943,N_7718,N_7784);
nor U7944 (N_7944,N_7754,N_7665);
nand U7945 (N_7945,N_7745,N_7615);
nor U7946 (N_7946,N_7749,N_7619);
nor U7947 (N_7947,N_7799,N_7723);
and U7948 (N_7948,N_7667,N_7671);
xnor U7949 (N_7949,N_7652,N_7663);
and U7950 (N_7950,N_7631,N_7721);
or U7951 (N_7951,N_7791,N_7764);
and U7952 (N_7952,N_7606,N_7721);
nand U7953 (N_7953,N_7665,N_7793);
nand U7954 (N_7954,N_7627,N_7685);
and U7955 (N_7955,N_7787,N_7798);
nand U7956 (N_7956,N_7666,N_7614);
nand U7957 (N_7957,N_7748,N_7740);
or U7958 (N_7958,N_7778,N_7649);
nand U7959 (N_7959,N_7773,N_7784);
nand U7960 (N_7960,N_7714,N_7662);
or U7961 (N_7961,N_7674,N_7626);
nor U7962 (N_7962,N_7623,N_7698);
nor U7963 (N_7963,N_7623,N_7678);
nand U7964 (N_7964,N_7642,N_7608);
and U7965 (N_7965,N_7651,N_7795);
nor U7966 (N_7966,N_7738,N_7686);
nand U7967 (N_7967,N_7604,N_7764);
or U7968 (N_7968,N_7752,N_7795);
and U7969 (N_7969,N_7693,N_7671);
nor U7970 (N_7970,N_7777,N_7671);
or U7971 (N_7971,N_7770,N_7782);
and U7972 (N_7972,N_7672,N_7721);
and U7973 (N_7973,N_7666,N_7657);
nand U7974 (N_7974,N_7623,N_7761);
and U7975 (N_7975,N_7739,N_7722);
or U7976 (N_7976,N_7778,N_7707);
or U7977 (N_7977,N_7637,N_7699);
nor U7978 (N_7978,N_7684,N_7665);
nand U7979 (N_7979,N_7780,N_7676);
or U7980 (N_7980,N_7621,N_7646);
and U7981 (N_7981,N_7610,N_7634);
or U7982 (N_7982,N_7733,N_7639);
or U7983 (N_7983,N_7613,N_7714);
and U7984 (N_7984,N_7778,N_7752);
nor U7985 (N_7985,N_7675,N_7641);
and U7986 (N_7986,N_7653,N_7788);
nor U7987 (N_7987,N_7692,N_7660);
and U7988 (N_7988,N_7781,N_7681);
and U7989 (N_7989,N_7680,N_7798);
or U7990 (N_7990,N_7735,N_7712);
and U7991 (N_7991,N_7763,N_7627);
nor U7992 (N_7992,N_7786,N_7766);
and U7993 (N_7993,N_7657,N_7774);
nand U7994 (N_7994,N_7690,N_7717);
nor U7995 (N_7995,N_7722,N_7626);
and U7996 (N_7996,N_7781,N_7704);
nor U7997 (N_7997,N_7655,N_7600);
nor U7998 (N_7998,N_7624,N_7705);
or U7999 (N_7999,N_7644,N_7769);
and U8000 (N_8000,N_7830,N_7898);
or U8001 (N_8001,N_7999,N_7823);
nor U8002 (N_8002,N_7983,N_7821);
and U8003 (N_8003,N_7961,N_7874);
and U8004 (N_8004,N_7833,N_7906);
and U8005 (N_8005,N_7811,N_7912);
and U8006 (N_8006,N_7952,N_7875);
nor U8007 (N_8007,N_7981,N_7896);
and U8008 (N_8008,N_7818,N_7815);
or U8009 (N_8009,N_7956,N_7938);
nor U8010 (N_8010,N_7856,N_7847);
or U8011 (N_8011,N_7939,N_7948);
nor U8012 (N_8012,N_7953,N_7834);
nand U8013 (N_8013,N_7998,N_7970);
nand U8014 (N_8014,N_7935,N_7976);
and U8015 (N_8015,N_7967,N_7929);
or U8016 (N_8016,N_7978,N_7972);
nand U8017 (N_8017,N_7853,N_7916);
nand U8018 (N_8018,N_7969,N_7840);
or U8019 (N_8019,N_7984,N_7934);
and U8020 (N_8020,N_7860,N_7841);
nor U8021 (N_8021,N_7927,N_7987);
nand U8022 (N_8022,N_7977,N_7985);
or U8023 (N_8023,N_7835,N_7836);
or U8024 (N_8024,N_7873,N_7975);
nand U8025 (N_8025,N_7880,N_7807);
or U8026 (N_8026,N_7950,N_7884);
nor U8027 (N_8027,N_7911,N_7892);
nor U8028 (N_8028,N_7918,N_7997);
or U8029 (N_8029,N_7806,N_7816);
nor U8030 (N_8030,N_7995,N_7982);
nor U8031 (N_8031,N_7960,N_7914);
nor U8032 (N_8032,N_7920,N_7812);
nor U8033 (N_8033,N_7851,N_7826);
nor U8034 (N_8034,N_7883,N_7996);
nor U8035 (N_8035,N_7825,N_7974);
or U8036 (N_8036,N_7846,N_7980);
nand U8037 (N_8037,N_7979,N_7936);
or U8038 (N_8038,N_7882,N_7890);
and U8039 (N_8039,N_7819,N_7990);
nand U8040 (N_8040,N_7885,N_7932);
nor U8041 (N_8041,N_7828,N_7813);
or U8042 (N_8042,N_7899,N_7910);
nand U8043 (N_8043,N_7859,N_7957);
and U8044 (N_8044,N_7829,N_7909);
or U8045 (N_8045,N_7824,N_7891);
and U8046 (N_8046,N_7852,N_7958);
nand U8047 (N_8047,N_7889,N_7964);
and U8048 (N_8048,N_7876,N_7837);
nand U8049 (N_8049,N_7888,N_7870);
and U8050 (N_8050,N_7921,N_7868);
or U8051 (N_8051,N_7871,N_7809);
nor U8052 (N_8052,N_7803,N_7965);
or U8053 (N_8053,N_7900,N_7915);
and U8054 (N_8054,N_7931,N_7872);
nand U8055 (N_8055,N_7902,N_7901);
and U8056 (N_8056,N_7937,N_7986);
nor U8057 (N_8057,N_7993,N_7801);
nand U8058 (N_8058,N_7861,N_7814);
nor U8059 (N_8059,N_7831,N_7849);
or U8060 (N_8060,N_7913,N_7854);
nor U8061 (N_8061,N_7949,N_7925);
nand U8062 (N_8062,N_7946,N_7855);
and U8063 (N_8063,N_7844,N_7994);
nand U8064 (N_8064,N_7930,N_7881);
or U8065 (N_8065,N_7842,N_7893);
or U8066 (N_8066,N_7804,N_7917);
nor U8067 (N_8067,N_7928,N_7827);
nor U8068 (N_8068,N_7887,N_7959);
nor U8069 (N_8069,N_7963,N_7800);
nor U8070 (N_8070,N_7905,N_7989);
nand U8071 (N_8071,N_7863,N_7848);
nand U8072 (N_8072,N_7805,N_7886);
and U8073 (N_8073,N_7877,N_7897);
and U8074 (N_8074,N_7857,N_7907);
nand U8075 (N_8075,N_7832,N_7904);
nor U8076 (N_8076,N_7947,N_7895);
or U8077 (N_8077,N_7924,N_7951);
or U8078 (N_8078,N_7988,N_7850);
and U8079 (N_8079,N_7941,N_7843);
nor U8080 (N_8080,N_7866,N_7968);
nand U8081 (N_8081,N_7864,N_7808);
nor U8082 (N_8082,N_7940,N_7820);
nor U8083 (N_8083,N_7839,N_7923);
nor U8084 (N_8084,N_7878,N_7992);
nor U8085 (N_8085,N_7973,N_7817);
nand U8086 (N_8086,N_7869,N_7867);
nor U8087 (N_8087,N_7944,N_7894);
or U8088 (N_8088,N_7908,N_7962);
or U8089 (N_8089,N_7919,N_7903);
nor U8090 (N_8090,N_7926,N_7879);
or U8091 (N_8091,N_7943,N_7838);
or U8092 (N_8092,N_7862,N_7865);
nand U8093 (N_8093,N_7955,N_7971);
nor U8094 (N_8094,N_7822,N_7810);
nor U8095 (N_8095,N_7945,N_7922);
nor U8096 (N_8096,N_7845,N_7858);
nor U8097 (N_8097,N_7942,N_7966);
or U8098 (N_8098,N_7991,N_7954);
nand U8099 (N_8099,N_7802,N_7933);
or U8100 (N_8100,N_7992,N_7942);
nor U8101 (N_8101,N_7878,N_7832);
or U8102 (N_8102,N_7891,N_7940);
nor U8103 (N_8103,N_7838,N_7821);
nor U8104 (N_8104,N_7847,N_7829);
xor U8105 (N_8105,N_7927,N_7848);
and U8106 (N_8106,N_7881,N_7839);
and U8107 (N_8107,N_7858,N_7904);
nand U8108 (N_8108,N_7968,N_7978);
nand U8109 (N_8109,N_7904,N_7863);
nand U8110 (N_8110,N_7888,N_7916);
nor U8111 (N_8111,N_7971,N_7873);
or U8112 (N_8112,N_7838,N_7997);
and U8113 (N_8113,N_7835,N_7867);
and U8114 (N_8114,N_7923,N_7895);
or U8115 (N_8115,N_7995,N_7844);
and U8116 (N_8116,N_7880,N_7960);
nand U8117 (N_8117,N_7987,N_7961);
and U8118 (N_8118,N_7962,N_7803);
nand U8119 (N_8119,N_7847,N_7914);
nand U8120 (N_8120,N_7896,N_7969);
nor U8121 (N_8121,N_7880,N_7949);
or U8122 (N_8122,N_7928,N_7821);
nand U8123 (N_8123,N_7986,N_7872);
nor U8124 (N_8124,N_7964,N_7879);
or U8125 (N_8125,N_7827,N_7921);
nand U8126 (N_8126,N_7949,N_7889);
nand U8127 (N_8127,N_7898,N_7923);
nor U8128 (N_8128,N_7982,N_7839);
or U8129 (N_8129,N_7942,N_7803);
nor U8130 (N_8130,N_7981,N_7803);
or U8131 (N_8131,N_7976,N_7881);
and U8132 (N_8132,N_7818,N_7958);
or U8133 (N_8133,N_7893,N_7847);
or U8134 (N_8134,N_7999,N_7828);
or U8135 (N_8135,N_7849,N_7852);
and U8136 (N_8136,N_7983,N_7975);
or U8137 (N_8137,N_7819,N_7837);
and U8138 (N_8138,N_7909,N_7818);
and U8139 (N_8139,N_7849,N_7830);
or U8140 (N_8140,N_7813,N_7966);
nand U8141 (N_8141,N_7846,N_7898);
nor U8142 (N_8142,N_7950,N_7843);
or U8143 (N_8143,N_7808,N_7846);
and U8144 (N_8144,N_7806,N_7948);
or U8145 (N_8145,N_7970,N_7869);
or U8146 (N_8146,N_7909,N_7924);
nand U8147 (N_8147,N_7889,N_7853);
nor U8148 (N_8148,N_7851,N_7887);
nor U8149 (N_8149,N_7827,N_7937);
and U8150 (N_8150,N_7953,N_7939);
nand U8151 (N_8151,N_7983,N_7943);
nor U8152 (N_8152,N_7979,N_7814);
and U8153 (N_8153,N_7940,N_7922);
and U8154 (N_8154,N_7820,N_7959);
and U8155 (N_8155,N_7932,N_7831);
and U8156 (N_8156,N_7911,N_7818);
nand U8157 (N_8157,N_7922,N_7931);
or U8158 (N_8158,N_7835,N_7977);
nor U8159 (N_8159,N_7831,N_7908);
or U8160 (N_8160,N_7999,N_7945);
nor U8161 (N_8161,N_7960,N_7843);
or U8162 (N_8162,N_7810,N_7911);
and U8163 (N_8163,N_7967,N_7908);
and U8164 (N_8164,N_7881,N_7890);
and U8165 (N_8165,N_7816,N_7809);
or U8166 (N_8166,N_7855,N_7914);
nand U8167 (N_8167,N_7921,N_7883);
nand U8168 (N_8168,N_7968,N_7907);
nor U8169 (N_8169,N_7803,N_7971);
or U8170 (N_8170,N_7906,N_7837);
and U8171 (N_8171,N_7935,N_7833);
or U8172 (N_8172,N_7825,N_7835);
and U8173 (N_8173,N_7858,N_7902);
and U8174 (N_8174,N_7857,N_7801);
nand U8175 (N_8175,N_7834,N_7991);
nor U8176 (N_8176,N_7877,N_7912);
nand U8177 (N_8177,N_7976,N_7925);
or U8178 (N_8178,N_7865,N_7836);
or U8179 (N_8179,N_7800,N_7817);
or U8180 (N_8180,N_7903,N_7867);
and U8181 (N_8181,N_7980,N_7928);
and U8182 (N_8182,N_7903,N_7856);
or U8183 (N_8183,N_7913,N_7983);
or U8184 (N_8184,N_7978,N_7871);
nor U8185 (N_8185,N_7923,N_7971);
and U8186 (N_8186,N_7821,N_7804);
nor U8187 (N_8187,N_7969,N_7947);
and U8188 (N_8188,N_7908,N_7993);
and U8189 (N_8189,N_7999,N_7982);
nand U8190 (N_8190,N_7935,N_7830);
or U8191 (N_8191,N_7908,N_7802);
and U8192 (N_8192,N_7834,N_7984);
and U8193 (N_8193,N_7907,N_7948);
or U8194 (N_8194,N_7801,N_7944);
or U8195 (N_8195,N_7882,N_7941);
nand U8196 (N_8196,N_7915,N_7815);
and U8197 (N_8197,N_7935,N_7802);
or U8198 (N_8198,N_7853,N_7845);
and U8199 (N_8199,N_7885,N_7890);
nor U8200 (N_8200,N_8008,N_8077);
nor U8201 (N_8201,N_8050,N_8063);
nor U8202 (N_8202,N_8188,N_8073);
or U8203 (N_8203,N_8173,N_8125);
or U8204 (N_8204,N_8115,N_8038);
nand U8205 (N_8205,N_8094,N_8084);
or U8206 (N_8206,N_8002,N_8139);
or U8207 (N_8207,N_8170,N_8099);
nand U8208 (N_8208,N_8070,N_8149);
nand U8209 (N_8209,N_8015,N_8141);
nor U8210 (N_8210,N_8054,N_8111);
nand U8211 (N_8211,N_8171,N_8059);
nor U8212 (N_8212,N_8080,N_8103);
nand U8213 (N_8213,N_8102,N_8184);
nand U8214 (N_8214,N_8035,N_8093);
and U8215 (N_8215,N_8065,N_8087);
or U8216 (N_8216,N_8071,N_8104);
or U8217 (N_8217,N_8058,N_8114);
and U8218 (N_8218,N_8025,N_8009);
or U8219 (N_8219,N_8082,N_8183);
nand U8220 (N_8220,N_8092,N_8194);
nor U8221 (N_8221,N_8024,N_8152);
nor U8222 (N_8222,N_8085,N_8081);
and U8223 (N_8223,N_8021,N_8055);
nor U8224 (N_8224,N_8068,N_8051);
nand U8225 (N_8225,N_8116,N_8143);
nand U8226 (N_8226,N_8067,N_8064);
nand U8227 (N_8227,N_8040,N_8052);
or U8228 (N_8228,N_8174,N_8083);
nor U8229 (N_8229,N_8126,N_8195);
and U8230 (N_8230,N_8120,N_8189);
nor U8231 (N_8231,N_8136,N_8107);
and U8232 (N_8232,N_8164,N_8098);
nand U8233 (N_8233,N_8047,N_8145);
nor U8234 (N_8234,N_8095,N_8033);
or U8235 (N_8235,N_8130,N_8165);
and U8236 (N_8236,N_8148,N_8016);
nor U8237 (N_8237,N_8131,N_8181);
nand U8238 (N_8238,N_8142,N_8182);
or U8239 (N_8239,N_8133,N_8113);
or U8240 (N_8240,N_8041,N_8122);
nand U8241 (N_8241,N_8167,N_8076);
nand U8242 (N_8242,N_8127,N_8062);
nand U8243 (N_8243,N_8043,N_8129);
or U8244 (N_8244,N_8155,N_8191);
and U8245 (N_8245,N_8049,N_8089);
nand U8246 (N_8246,N_8088,N_8180);
and U8247 (N_8247,N_8156,N_8109);
nand U8248 (N_8248,N_8079,N_8176);
nor U8249 (N_8249,N_8169,N_8010);
nor U8250 (N_8250,N_8190,N_8044);
and U8251 (N_8251,N_8100,N_8154);
or U8252 (N_8252,N_8056,N_8006);
nor U8253 (N_8253,N_8185,N_8177);
nand U8254 (N_8254,N_8161,N_8036);
and U8255 (N_8255,N_8000,N_8144);
nand U8256 (N_8256,N_8037,N_8066);
nor U8257 (N_8257,N_8121,N_8022);
nand U8258 (N_8258,N_8012,N_8005);
nor U8259 (N_8259,N_8192,N_8007);
or U8260 (N_8260,N_8001,N_8128);
or U8261 (N_8261,N_8186,N_8137);
nand U8262 (N_8262,N_8003,N_8159);
nand U8263 (N_8263,N_8060,N_8175);
or U8264 (N_8264,N_8091,N_8123);
nor U8265 (N_8265,N_8096,N_8075);
nand U8266 (N_8266,N_8197,N_8112);
nand U8267 (N_8267,N_8032,N_8042);
nor U8268 (N_8268,N_8030,N_8158);
or U8269 (N_8269,N_8105,N_8046);
nand U8270 (N_8270,N_8074,N_8019);
nor U8271 (N_8271,N_8048,N_8199);
or U8272 (N_8272,N_8187,N_8028);
nand U8273 (N_8273,N_8069,N_8086);
and U8274 (N_8274,N_8110,N_8108);
nand U8275 (N_8275,N_8078,N_8140);
or U8276 (N_8276,N_8146,N_8027);
and U8277 (N_8277,N_8134,N_8198);
nand U8278 (N_8278,N_8011,N_8196);
and U8279 (N_8279,N_8029,N_8097);
nand U8280 (N_8280,N_8132,N_8053);
nor U8281 (N_8281,N_8138,N_8135);
nor U8282 (N_8282,N_8014,N_8168);
nand U8283 (N_8283,N_8124,N_8178);
or U8284 (N_8284,N_8020,N_8106);
nor U8285 (N_8285,N_8117,N_8045);
nor U8286 (N_8286,N_8172,N_8031);
nand U8287 (N_8287,N_8160,N_8057);
and U8288 (N_8288,N_8017,N_8101);
xor U8289 (N_8289,N_8162,N_8151);
nand U8290 (N_8290,N_8004,N_8018);
nand U8291 (N_8291,N_8166,N_8193);
nand U8292 (N_8292,N_8147,N_8072);
nor U8293 (N_8293,N_8026,N_8179);
nand U8294 (N_8294,N_8118,N_8153);
nor U8295 (N_8295,N_8150,N_8013);
and U8296 (N_8296,N_8157,N_8163);
and U8297 (N_8297,N_8039,N_8090);
nor U8298 (N_8298,N_8119,N_8034);
or U8299 (N_8299,N_8061,N_8023);
nor U8300 (N_8300,N_8014,N_8151);
and U8301 (N_8301,N_8177,N_8195);
nand U8302 (N_8302,N_8050,N_8075);
nand U8303 (N_8303,N_8113,N_8101);
or U8304 (N_8304,N_8029,N_8107);
xor U8305 (N_8305,N_8104,N_8121);
and U8306 (N_8306,N_8088,N_8126);
or U8307 (N_8307,N_8068,N_8013);
nor U8308 (N_8308,N_8023,N_8108);
nor U8309 (N_8309,N_8135,N_8049);
or U8310 (N_8310,N_8136,N_8060);
nand U8311 (N_8311,N_8002,N_8137);
nand U8312 (N_8312,N_8150,N_8102);
or U8313 (N_8313,N_8001,N_8125);
nor U8314 (N_8314,N_8122,N_8057);
nand U8315 (N_8315,N_8022,N_8195);
nand U8316 (N_8316,N_8030,N_8046);
and U8317 (N_8317,N_8048,N_8188);
nand U8318 (N_8318,N_8009,N_8086);
and U8319 (N_8319,N_8022,N_8199);
nand U8320 (N_8320,N_8101,N_8024);
or U8321 (N_8321,N_8023,N_8065);
nor U8322 (N_8322,N_8066,N_8108);
nor U8323 (N_8323,N_8143,N_8174);
nor U8324 (N_8324,N_8034,N_8130);
and U8325 (N_8325,N_8084,N_8140);
or U8326 (N_8326,N_8111,N_8175);
nand U8327 (N_8327,N_8051,N_8114);
nand U8328 (N_8328,N_8128,N_8189);
and U8329 (N_8329,N_8117,N_8034);
nand U8330 (N_8330,N_8171,N_8022);
nand U8331 (N_8331,N_8028,N_8193);
nor U8332 (N_8332,N_8005,N_8196);
and U8333 (N_8333,N_8064,N_8065);
and U8334 (N_8334,N_8087,N_8179);
nand U8335 (N_8335,N_8198,N_8010);
nand U8336 (N_8336,N_8035,N_8017);
nand U8337 (N_8337,N_8114,N_8062);
and U8338 (N_8338,N_8198,N_8050);
nand U8339 (N_8339,N_8137,N_8106);
or U8340 (N_8340,N_8104,N_8108);
nand U8341 (N_8341,N_8167,N_8079);
and U8342 (N_8342,N_8059,N_8039);
and U8343 (N_8343,N_8068,N_8096);
and U8344 (N_8344,N_8069,N_8006);
nand U8345 (N_8345,N_8017,N_8177);
nand U8346 (N_8346,N_8086,N_8152);
nor U8347 (N_8347,N_8163,N_8019);
or U8348 (N_8348,N_8027,N_8167);
nand U8349 (N_8349,N_8073,N_8028);
nand U8350 (N_8350,N_8009,N_8088);
nand U8351 (N_8351,N_8087,N_8055);
and U8352 (N_8352,N_8040,N_8042);
and U8353 (N_8353,N_8026,N_8157);
nand U8354 (N_8354,N_8081,N_8155);
and U8355 (N_8355,N_8112,N_8021);
nor U8356 (N_8356,N_8142,N_8055);
or U8357 (N_8357,N_8165,N_8155);
or U8358 (N_8358,N_8050,N_8049);
or U8359 (N_8359,N_8106,N_8120);
and U8360 (N_8360,N_8171,N_8155);
and U8361 (N_8361,N_8086,N_8102);
and U8362 (N_8362,N_8005,N_8188);
and U8363 (N_8363,N_8079,N_8021);
nor U8364 (N_8364,N_8011,N_8192);
nor U8365 (N_8365,N_8134,N_8098);
and U8366 (N_8366,N_8018,N_8179);
and U8367 (N_8367,N_8060,N_8103);
or U8368 (N_8368,N_8006,N_8035);
or U8369 (N_8369,N_8179,N_8042);
and U8370 (N_8370,N_8138,N_8148);
or U8371 (N_8371,N_8129,N_8116);
and U8372 (N_8372,N_8088,N_8172);
and U8373 (N_8373,N_8129,N_8080);
and U8374 (N_8374,N_8056,N_8189);
or U8375 (N_8375,N_8011,N_8073);
and U8376 (N_8376,N_8163,N_8194);
nand U8377 (N_8377,N_8014,N_8035);
and U8378 (N_8378,N_8108,N_8116);
nor U8379 (N_8379,N_8170,N_8103);
or U8380 (N_8380,N_8186,N_8096);
nor U8381 (N_8381,N_8097,N_8030);
and U8382 (N_8382,N_8128,N_8100);
and U8383 (N_8383,N_8150,N_8040);
xor U8384 (N_8384,N_8150,N_8075);
nor U8385 (N_8385,N_8138,N_8188);
and U8386 (N_8386,N_8084,N_8023);
nor U8387 (N_8387,N_8038,N_8060);
and U8388 (N_8388,N_8194,N_8180);
nand U8389 (N_8389,N_8106,N_8018);
nor U8390 (N_8390,N_8054,N_8117);
nor U8391 (N_8391,N_8138,N_8167);
nand U8392 (N_8392,N_8049,N_8155);
and U8393 (N_8393,N_8053,N_8150);
nor U8394 (N_8394,N_8191,N_8040);
nand U8395 (N_8395,N_8175,N_8172);
and U8396 (N_8396,N_8110,N_8055);
or U8397 (N_8397,N_8029,N_8056);
nand U8398 (N_8398,N_8187,N_8061);
nand U8399 (N_8399,N_8099,N_8022);
nand U8400 (N_8400,N_8352,N_8227);
nor U8401 (N_8401,N_8296,N_8368);
nor U8402 (N_8402,N_8334,N_8340);
nor U8403 (N_8403,N_8283,N_8217);
or U8404 (N_8404,N_8268,N_8286);
or U8405 (N_8405,N_8232,N_8299);
nor U8406 (N_8406,N_8225,N_8273);
nor U8407 (N_8407,N_8295,N_8235);
and U8408 (N_8408,N_8318,N_8231);
and U8409 (N_8409,N_8350,N_8335);
nand U8410 (N_8410,N_8275,N_8282);
nand U8411 (N_8411,N_8255,N_8220);
nor U8412 (N_8412,N_8320,N_8381);
nor U8413 (N_8413,N_8358,N_8263);
nor U8414 (N_8414,N_8298,N_8397);
or U8415 (N_8415,N_8308,N_8214);
nor U8416 (N_8416,N_8256,N_8386);
nand U8417 (N_8417,N_8229,N_8343);
and U8418 (N_8418,N_8319,N_8223);
and U8419 (N_8419,N_8250,N_8267);
and U8420 (N_8420,N_8379,N_8242);
and U8421 (N_8421,N_8288,N_8251);
nor U8422 (N_8422,N_8233,N_8388);
or U8423 (N_8423,N_8376,N_8276);
and U8424 (N_8424,N_8355,N_8226);
xor U8425 (N_8425,N_8345,N_8322);
and U8426 (N_8426,N_8364,N_8359);
and U8427 (N_8427,N_8375,N_8324);
nor U8428 (N_8428,N_8351,N_8269);
nand U8429 (N_8429,N_8313,N_8248);
or U8430 (N_8430,N_8219,N_8237);
or U8431 (N_8431,N_8290,N_8395);
nand U8432 (N_8432,N_8245,N_8236);
nand U8433 (N_8433,N_8289,N_8385);
nor U8434 (N_8434,N_8384,N_8363);
nand U8435 (N_8435,N_8323,N_8253);
nand U8436 (N_8436,N_8371,N_8338);
nand U8437 (N_8437,N_8393,N_8241);
and U8438 (N_8438,N_8291,N_8314);
or U8439 (N_8439,N_8317,N_8218);
and U8440 (N_8440,N_8398,N_8292);
nor U8441 (N_8441,N_8344,N_8311);
and U8442 (N_8442,N_8331,N_8370);
nand U8443 (N_8443,N_8304,N_8302);
nor U8444 (N_8444,N_8391,N_8383);
and U8445 (N_8445,N_8202,N_8216);
and U8446 (N_8446,N_8339,N_8394);
nand U8447 (N_8447,N_8261,N_8309);
or U8448 (N_8448,N_8305,N_8208);
nand U8449 (N_8449,N_8215,N_8316);
nand U8450 (N_8450,N_8310,N_8347);
nand U8451 (N_8451,N_8209,N_8228);
or U8452 (N_8452,N_8265,N_8259);
or U8453 (N_8453,N_8260,N_8264);
nand U8454 (N_8454,N_8252,N_8207);
nor U8455 (N_8455,N_8287,N_8201);
and U8456 (N_8456,N_8306,N_8200);
or U8457 (N_8457,N_8377,N_8204);
nand U8458 (N_8458,N_8206,N_8378);
or U8459 (N_8459,N_8382,N_8281);
or U8460 (N_8460,N_8353,N_8303);
nand U8461 (N_8461,N_8238,N_8373);
or U8462 (N_8462,N_8239,N_8360);
nand U8463 (N_8463,N_8329,N_8222);
nor U8464 (N_8464,N_8224,N_8221);
nand U8465 (N_8465,N_8257,N_8234);
nand U8466 (N_8466,N_8399,N_8266);
and U8467 (N_8467,N_8346,N_8369);
nor U8468 (N_8468,N_8396,N_8300);
and U8469 (N_8469,N_8357,N_8367);
or U8470 (N_8470,N_8203,N_8244);
nor U8471 (N_8471,N_8328,N_8272);
xor U8472 (N_8472,N_8389,N_8332);
or U8473 (N_8473,N_8294,N_8284);
nor U8474 (N_8474,N_8213,N_8333);
or U8475 (N_8475,N_8243,N_8321);
or U8476 (N_8476,N_8274,N_8211);
or U8477 (N_8477,N_8348,N_8387);
or U8478 (N_8478,N_8212,N_8307);
nor U8479 (N_8479,N_8349,N_8277);
nor U8480 (N_8480,N_8278,N_8341);
nand U8481 (N_8481,N_8374,N_8254);
xnor U8482 (N_8482,N_8279,N_8293);
and U8483 (N_8483,N_8246,N_8325);
nand U8484 (N_8484,N_8326,N_8297);
nor U8485 (N_8485,N_8247,N_8271);
nor U8486 (N_8486,N_8301,N_8249);
or U8487 (N_8487,N_8280,N_8312);
nand U8488 (N_8488,N_8210,N_8356);
and U8489 (N_8489,N_8205,N_8327);
nand U8490 (N_8490,N_8342,N_8365);
and U8491 (N_8491,N_8366,N_8258);
nor U8492 (N_8492,N_8230,N_8270);
nor U8493 (N_8493,N_8315,N_8380);
or U8494 (N_8494,N_8337,N_8354);
or U8495 (N_8495,N_8390,N_8372);
or U8496 (N_8496,N_8285,N_8336);
and U8497 (N_8497,N_8262,N_8392);
nor U8498 (N_8498,N_8240,N_8361);
and U8499 (N_8499,N_8330,N_8362);
and U8500 (N_8500,N_8354,N_8227);
and U8501 (N_8501,N_8258,N_8232);
nand U8502 (N_8502,N_8286,N_8300);
or U8503 (N_8503,N_8330,N_8342);
nand U8504 (N_8504,N_8209,N_8317);
nor U8505 (N_8505,N_8393,N_8329);
nor U8506 (N_8506,N_8241,N_8267);
nor U8507 (N_8507,N_8231,N_8358);
and U8508 (N_8508,N_8344,N_8219);
and U8509 (N_8509,N_8352,N_8343);
and U8510 (N_8510,N_8276,N_8265);
nand U8511 (N_8511,N_8309,N_8394);
and U8512 (N_8512,N_8202,N_8300);
nor U8513 (N_8513,N_8243,N_8252);
and U8514 (N_8514,N_8313,N_8291);
nor U8515 (N_8515,N_8326,N_8222);
nor U8516 (N_8516,N_8344,N_8338);
or U8517 (N_8517,N_8373,N_8222);
or U8518 (N_8518,N_8315,N_8291);
nor U8519 (N_8519,N_8322,N_8315);
or U8520 (N_8520,N_8339,N_8319);
nor U8521 (N_8521,N_8327,N_8299);
or U8522 (N_8522,N_8358,N_8229);
nand U8523 (N_8523,N_8353,N_8377);
nand U8524 (N_8524,N_8350,N_8365);
or U8525 (N_8525,N_8328,N_8323);
and U8526 (N_8526,N_8268,N_8365);
and U8527 (N_8527,N_8283,N_8306);
nor U8528 (N_8528,N_8216,N_8322);
or U8529 (N_8529,N_8302,N_8373);
or U8530 (N_8530,N_8339,N_8284);
xnor U8531 (N_8531,N_8225,N_8243);
and U8532 (N_8532,N_8372,N_8373);
nand U8533 (N_8533,N_8205,N_8204);
nand U8534 (N_8534,N_8330,N_8351);
and U8535 (N_8535,N_8224,N_8344);
and U8536 (N_8536,N_8207,N_8343);
or U8537 (N_8537,N_8354,N_8363);
or U8538 (N_8538,N_8262,N_8327);
and U8539 (N_8539,N_8372,N_8339);
and U8540 (N_8540,N_8370,N_8380);
and U8541 (N_8541,N_8200,N_8363);
nand U8542 (N_8542,N_8258,N_8263);
or U8543 (N_8543,N_8221,N_8299);
or U8544 (N_8544,N_8285,N_8385);
and U8545 (N_8545,N_8301,N_8289);
and U8546 (N_8546,N_8369,N_8221);
or U8547 (N_8547,N_8203,N_8384);
or U8548 (N_8548,N_8232,N_8238);
nor U8549 (N_8549,N_8326,N_8369);
xor U8550 (N_8550,N_8247,N_8356);
or U8551 (N_8551,N_8347,N_8326);
or U8552 (N_8552,N_8212,N_8254);
nand U8553 (N_8553,N_8379,N_8345);
or U8554 (N_8554,N_8320,N_8245);
and U8555 (N_8555,N_8220,N_8223);
or U8556 (N_8556,N_8362,N_8279);
and U8557 (N_8557,N_8283,N_8385);
nand U8558 (N_8558,N_8352,N_8250);
or U8559 (N_8559,N_8295,N_8377);
and U8560 (N_8560,N_8343,N_8311);
nor U8561 (N_8561,N_8375,N_8333);
or U8562 (N_8562,N_8358,N_8350);
nand U8563 (N_8563,N_8382,N_8242);
and U8564 (N_8564,N_8384,N_8389);
and U8565 (N_8565,N_8288,N_8283);
nor U8566 (N_8566,N_8377,N_8328);
or U8567 (N_8567,N_8249,N_8361);
and U8568 (N_8568,N_8303,N_8227);
and U8569 (N_8569,N_8386,N_8384);
nand U8570 (N_8570,N_8352,N_8385);
nor U8571 (N_8571,N_8342,N_8359);
nand U8572 (N_8572,N_8274,N_8292);
and U8573 (N_8573,N_8257,N_8263);
nor U8574 (N_8574,N_8354,N_8298);
nand U8575 (N_8575,N_8397,N_8379);
nor U8576 (N_8576,N_8267,N_8397);
or U8577 (N_8577,N_8315,N_8339);
nand U8578 (N_8578,N_8298,N_8322);
and U8579 (N_8579,N_8269,N_8361);
xnor U8580 (N_8580,N_8376,N_8269);
and U8581 (N_8581,N_8367,N_8203);
and U8582 (N_8582,N_8297,N_8210);
and U8583 (N_8583,N_8291,N_8246);
nand U8584 (N_8584,N_8379,N_8388);
nor U8585 (N_8585,N_8259,N_8283);
nand U8586 (N_8586,N_8349,N_8326);
and U8587 (N_8587,N_8264,N_8237);
nand U8588 (N_8588,N_8386,N_8211);
or U8589 (N_8589,N_8219,N_8235);
nor U8590 (N_8590,N_8377,N_8227);
nor U8591 (N_8591,N_8342,N_8231);
or U8592 (N_8592,N_8375,N_8250);
xor U8593 (N_8593,N_8226,N_8345);
nor U8594 (N_8594,N_8354,N_8305);
nand U8595 (N_8595,N_8379,N_8253);
or U8596 (N_8596,N_8338,N_8397);
nand U8597 (N_8597,N_8280,N_8351);
or U8598 (N_8598,N_8356,N_8355);
or U8599 (N_8599,N_8256,N_8365);
or U8600 (N_8600,N_8492,N_8534);
and U8601 (N_8601,N_8566,N_8481);
nand U8602 (N_8602,N_8491,N_8418);
or U8603 (N_8603,N_8427,N_8458);
nor U8604 (N_8604,N_8408,N_8519);
and U8605 (N_8605,N_8426,N_8567);
nand U8606 (N_8606,N_8589,N_8553);
or U8607 (N_8607,N_8493,N_8510);
nand U8608 (N_8608,N_8490,N_8503);
and U8609 (N_8609,N_8524,N_8449);
nand U8610 (N_8610,N_8480,N_8414);
or U8611 (N_8611,N_8420,N_8558);
nand U8612 (N_8612,N_8516,N_8422);
and U8613 (N_8613,N_8591,N_8438);
and U8614 (N_8614,N_8451,N_8525);
and U8615 (N_8615,N_8499,N_8587);
and U8616 (N_8616,N_8563,N_8515);
and U8617 (N_8617,N_8544,N_8448);
nand U8618 (N_8618,N_8541,N_8407);
and U8619 (N_8619,N_8550,N_8527);
nand U8620 (N_8620,N_8454,N_8470);
or U8621 (N_8621,N_8538,N_8574);
nor U8622 (N_8622,N_8536,N_8500);
or U8623 (N_8623,N_8494,N_8496);
nand U8624 (N_8624,N_8512,N_8593);
or U8625 (N_8625,N_8529,N_8580);
nand U8626 (N_8626,N_8595,N_8495);
nor U8627 (N_8627,N_8437,N_8476);
or U8628 (N_8628,N_8513,N_8453);
or U8629 (N_8629,N_8522,N_8477);
and U8630 (N_8630,N_8533,N_8577);
and U8631 (N_8631,N_8526,N_8487);
nor U8632 (N_8632,N_8445,N_8401);
or U8633 (N_8633,N_8409,N_8552);
nand U8634 (N_8634,N_8464,N_8447);
and U8635 (N_8635,N_8471,N_8583);
nand U8636 (N_8636,N_8585,N_8540);
nor U8637 (N_8637,N_8537,N_8465);
nand U8638 (N_8638,N_8594,N_8561);
or U8639 (N_8639,N_8425,N_8456);
and U8640 (N_8640,N_8475,N_8459);
or U8641 (N_8641,N_8586,N_8545);
and U8642 (N_8642,N_8466,N_8483);
or U8643 (N_8643,N_8578,N_8472);
or U8644 (N_8644,N_8421,N_8575);
xnor U8645 (N_8645,N_8479,N_8506);
xnor U8646 (N_8646,N_8489,N_8528);
and U8647 (N_8647,N_8505,N_8497);
nand U8648 (N_8648,N_8597,N_8457);
and U8649 (N_8649,N_8570,N_8444);
and U8650 (N_8650,N_8554,N_8424);
and U8651 (N_8651,N_8435,N_8509);
nand U8652 (N_8652,N_8579,N_8441);
or U8653 (N_8653,N_8549,N_8571);
nor U8654 (N_8654,N_8588,N_8542);
and U8655 (N_8655,N_8598,N_8400);
nand U8656 (N_8656,N_8402,N_8461);
or U8657 (N_8657,N_8599,N_8547);
nor U8658 (N_8658,N_8485,N_8412);
and U8659 (N_8659,N_8562,N_8504);
or U8660 (N_8660,N_8436,N_8463);
or U8661 (N_8661,N_8439,N_8415);
nor U8662 (N_8662,N_8416,N_8428);
or U8663 (N_8663,N_8423,N_8507);
and U8664 (N_8664,N_8584,N_8548);
and U8665 (N_8665,N_8565,N_8560);
and U8666 (N_8666,N_8413,N_8521);
and U8667 (N_8667,N_8430,N_8468);
or U8668 (N_8668,N_8484,N_8531);
and U8669 (N_8669,N_8535,N_8462);
and U8670 (N_8670,N_8406,N_8569);
nand U8671 (N_8671,N_8469,N_8532);
nand U8672 (N_8672,N_8455,N_8517);
and U8673 (N_8673,N_8543,N_8411);
and U8674 (N_8674,N_8432,N_8482);
nand U8675 (N_8675,N_8508,N_8404);
nor U8676 (N_8676,N_8530,N_8478);
and U8677 (N_8677,N_8440,N_8596);
nand U8678 (N_8678,N_8473,N_8518);
or U8679 (N_8679,N_8498,N_8442);
and U8680 (N_8680,N_8564,N_8419);
nor U8681 (N_8681,N_8501,N_8581);
nor U8682 (N_8682,N_8502,N_8557);
nor U8683 (N_8683,N_8486,N_8582);
nand U8684 (N_8684,N_8410,N_8590);
nor U8685 (N_8685,N_8443,N_8434);
and U8686 (N_8686,N_8555,N_8546);
nor U8687 (N_8687,N_8514,N_8403);
nand U8688 (N_8688,N_8433,N_8450);
nand U8689 (N_8689,N_8405,N_8523);
or U8690 (N_8690,N_8488,N_8556);
nor U8691 (N_8691,N_8551,N_8592);
and U8692 (N_8692,N_8576,N_8511);
or U8693 (N_8693,N_8452,N_8417);
or U8694 (N_8694,N_8431,N_8559);
or U8695 (N_8695,N_8568,N_8446);
or U8696 (N_8696,N_8460,N_8474);
and U8697 (N_8697,N_8539,N_8573);
and U8698 (N_8698,N_8572,N_8520);
or U8699 (N_8699,N_8467,N_8429);
or U8700 (N_8700,N_8438,N_8419);
or U8701 (N_8701,N_8421,N_8490);
nand U8702 (N_8702,N_8432,N_8458);
or U8703 (N_8703,N_8514,N_8527);
nand U8704 (N_8704,N_8551,N_8520);
or U8705 (N_8705,N_8471,N_8595);
nor U8706 (N_8706,N_8470,N_8495);
xnor U8707 (N_8707,N_8591,N_8539);
nor U8708 (N_8708,N_8555,N_8442);
and U8709 (N_8709,N_8533,N_8479);
and U8710 (N_8710,N_8499,N_8470);
nor U8711 (N_8711,N_8423,N_8435);
nor U8712 (N_8712,N_8505,N_8589);
or U8713 (N_8713,N_8467,N_8434);
nand U8714 (N_8714,N_8414,N_8546);
nor U8715 (N_8715,N_8491,N_8425);
or U8716 (N_8716,N_8494,N_8554);
or U8717 (N_8717,N_8475,N_8402);
nand U8718 (N_8718,N_8409,N_8446);
nor U8719 (N_8719,N_8446,N_8463);
and U8720 (N_8720,N_8450,N_8570);
or U8721 (N_8721,N_8585,N_8454);
nor U8722 (N_8722,N_8502,N_8400);
nor U8723 (N_8723,N_8462,N_8534);
and U8724 (N_8724,N_8559,N_8564);
or U8725 (N_8725,N_8472,N_8425);
nand U8726 (N_8726,N_8560,N_8555);
nor U8727 (N_8727,N_8548,N_8409);
or U8728 (N_8728,N_8402,N_8476);
and U8729 (N_8729,N_8514,N_8568);
nor U8730 (N_8730,N_8487,N_8470);
nor U8731 (N_8731,N_8569,N_8413);
nor U8732 (N_8732,N_8481,N_8558);
nor U8733 (N_8733,N_8522,N_8455);
and U8734 (N_8734,N_8489,N_8425);
nand U8735 (N_8735,N_8598,N_8516);
and U8736 (N_8736,N_8465,N_8461);
nor U8737 (N_8737,N_8510,N_8590);
nor U8738 (N_8738,N_8501,N_8427);
nand U8739 (N_8739,N_8521,N_8538);
nand U8740 (N_8740,N_8441,N_8594);
nor U8741 (N_8741,N_8501,N_8585);
or U8742 (N_8742,N_8439,N_8504);
nor U8743 (N_8743,N_8418,N_8569);
nor U8744 (N_8744,N_8463,N_8447);
nand U8745 (N_8745,N_8512,N_8426);
and U8746 (N_8746,N_8504,N_8437);
nand U8747 (N_8747,N_8456,N_8501);
nor U8748 (N_8748,N_8451,N_8574);
and U8749 (N_8749,N_8463,N_8421);
nor U8750 (N_8750,N_8515,N_8494);
nand U8751 (N_8751,N_8503,N_8494);
nor U8752 (N_8752,N_8518,N_8588);
or U8753 (N_8753,N_8437,N_8539);
nand U8754 (N_8754,N_8423,N_8470);
and U8755 (N_8755,N_8542,N_8527);
nor U8756 (N_8756,N_8540,N_8497);
and U8757 (N_8757,N_8486,N_8464);
nand U8758 (N_8758,N_8457,N_8405);
nand U8759 (N_8759,N_8496,N_8597);
or U8760 (N_8760,N_8429,N_8534);
nand U8761 (N_8761,N_8443,N_8493);
and U8762 (N_8762,N_8542,N_8445);
nor U8763 (N_8763,N_8511,N_8446);
nand U8764 (N_8764,N_8552,N_8406);
nand U8765 (N_8765,N_8488,N_8436);
nor U8766 (N_8766,N_8478,N_8590);
or U8767 (N_8767,N_8409,N_8457);
and U8768 (N_8768,N_8491,N_8408);
or U8769 (N_8769,N_8547,N_8530);
or U8770 (N_8770,N_8445,N_8500);
or U8771 (N_8771,N_8415,N_8516);
nor U8772 (N_8772,N_8593,N_8526);
nor U8773 (N_8773,N_8493,N_8523);
nor U8774 (N_8774,N_8526,N_8589);
and U8775 (N_8775,N_8517,N_8521);
nor U8776 (N_8776,N_8441,N_8540);
nand U8777 (N_8777,N_8470,N_8531);
or U8778 (N_8778,N_8455,N_8499);
nor U8779 (N_8779,N_8521,N_8477);
nor U8780 (N_8780,N_8407,N_8431);
and U8781 (N_8781,N_8535,N_8579);
and U8782 (N_8782,N_8403,N_8447);
nor U8783 (N_8783,N_8420,N_8536);
or U8784 (N_8784,N_8421,N_8436);
or U8785 (N_8785,N_8426,N_8405);
and U8786 (N_8786,N_8595,N_8547);
nand U8787 (N_8787,N_8510,N_8550);
and U8788 (N_8788,N_8579,N_8439);
nand U8789 (N_8789,N_8402,N_8464);
and U8790 (N_8790,N_8479,N_8434);
or U8791 (N_8791,N_8431,N_8599);
or U8792 (N_8792,N_8441,N_8553);
nor U8793 (N_8793,N_8501,N_8550);
nand U8794 (N_8794,N_8427,N_8403);
nand U8795 (N_8795,N_8585,N_8410);
nand U8796 (N_8796,N_8441,N_8422);
nor U8797 (N_8797,N_8419,N_8529);
nor U8798 (N_8798,N_8477,N_8496);
and U8799 (N_8799,N_8498,N_8555);
nand U8800 (N_8800,N_8672,N_8674);
and U8801 (N_8801,N_8624,N_8701);
or U8802 (N_8802,N_8766,N_8751);
or U8803 (N_8803,N_8703,N_8603);
and U8804 (N_8804,N_8753,N_8640);
and U8805 (N_8805,N_8785,N_8699);
or U8806 (N_8806,N_8634,N_8739);
or U8807 (N_8807,N_8694,N_8736);
nand U8808 (N_8808,N_8649,N_8782);
and U8809 (N_8809,N_8648,N_8748);
or U8810 (N_8810,N_8673,N_8670);
or U8811 (N_8811,N_8617,N_8720);
nand U8812 (N_8812,N_8675,N_8615);
nand U8813 (N_8813,N_8793,N_8667);
and U8814 (N_8814,N_8600,N_8781);
nand U8815 (N_8815,N_8740,N_8714);
nor U8816 (N_8816,N_8795,N_8685);
nand U8817 (N_8817,N_8622,N_8663);
and U8818 (N_8818,N_8619,N_8724);
or U8819 (N_8819,N_8779,N_8770);
nand U8820 (N_8820,N_8635,N_8711);
nor U8821 (N_8821,N_8680,N_8655);
nand U8822 (N_8822,N_8741,N_8657);
and U8823 (N_8823,N_8723,N_8602);
and U8824 (N_8824,N_8641,N_8767);
or U8825 (N_8825,N_8721,N_8716);
nor U8826 (N_8826,N_8722,N_8726);
or U8827 (N_8827,N_8768,N_8661);
and U8828 (N_8828,N_8651,N_8778);
nor U8829 (N_8829,N_8611,N_8758);
and U8830 (N_8830,N_8623,N_8616);
or U8831 (N_8831,N_8700,N_8637);
nand U8832 (N_8832,N_8764,N_8790);
nor U8833 (N_8833,N_8752,N_8717);
and U8834 (N_8834,N_8710,N_8730);
nand U8835 (N_8835,N_8610,N_8747);
and U8836 (N_8836,N_8787,N_8712);
or U8837 (N_8837,N_8774,N_8702);
nor U8838 (N_8838,N_8731,N_8783);
and U8839 (N_8839,N_8705,N_8742);
nor U8840 (N_8840,N_8601,N_8695);
or U8841 (N_8841,N_8660,N_8765);
and U8842 (N_8842,N_8656,N_8628);
and U8843 (N_8843,N_8683,N_8643);
nor U8844 (N_8844,N_8646,N_8665);
nand U8845 (N_8845,N_8792,N_8604);
nor U8846 (N_8846,N_8664,N_8620);
or U8847 (N_8847,N_8608,N_8784);
or U8848 (N_8848,N_8677,N_8737);
nor U8849 (N_8849,N_8749,N_8627);
or U8850 (N_8850,N_8735,N_8773);
nand U8851 (N_8851,N_8750,N_8756);
and U8852 (N_8852,N_8757,N_8644);
or U8853 (N_8853,N_8798,N_8607);
nor U8854 (N_8854,N_8653,N_8780);
nor U8855 (N_8855,N_8679,N_8625);
nand U8856 (N_8856,N_8630,N_8733);
or U8857 (N_8857,N_8746,N_8686);
and U8858 (N_8858,N_8709,N_8659);
nor U8859 (N_8859,N_8638,N_8727);
nor U8860 (N_8860,N_8609,N_8734);
or U8861 (N_8861,N_8605,N_8642);
or U8862 (N_8862,N_8732,N_8718);
nand U8863 (N_8863,N_8763,N_8687);
nand U8864 (N_8864,N_8652,N_8698);
and U8865 (N_8865,N_8715,N_8691);
nor U8866 (N_8866,N_8725,N_8708);
and U8867 (N_8867,N_8632,N_8697);
or U8868 (N_8868,N_8743,N_8797);
and U8869 (N_8869,N_8707,N_8626);
and U8870 (N_8870,N_8706,N_8676);
xor U8871 (N_8871,N_8678,N_8755);
nand U8872 (N_8872,N_8738,N_8786);
or U8873 (N_8873,N_8729,N_8688);
nand U8874 (N_8874,N_8788,N_8704);
nor U8875 (N_8875,N_8639,N_8633);
and U8876 (N_8876,N_8794,N_8671);
or U8877 (N_8877,N_8719,N_8776);
nor U8878 (N_8878,N_8696,N_8692);
nand U8879 (N_8879,N_8669,N_8666);
or U8880 (N_8880,N_8769,N_8612);
nand U8881 (N_8881,N_8799,N_8760);
nor U8882 (N_8882,N_8668,N_8789);
and U8883 (N_8883,N_8654,N_8650);
nor U8884 (N_8884,N_8682,N_8761);
nand U8885 (N_8885,N_8631,N_8728);
nor U8886 (N_8886,N_8636,N_8658);
nor U8887 (N_8887,N_8744,N_8613);
nand U8888 (N_8888,N_8754,N_8681);
nor U8889 (N_8889,N_8693,N_8662);
nand U8890 (N_8890,N_8629,N_8689);
and U8891 (N_8891,N_8618,N_8690);
nand U8892 (N_8892,N_8759,N_8762);
nor U8893 (N_8893,N_8791,N_8684);
nand U8894 (N_8894,N_8645,N_8771);
nor U8895 (N_8895,N_8647,N_8621);
or U8896 (N_8896,N_8777,N_8772);
or U8897 (N_8897,N_8745,N_8775);
nor U8898 (N_8898,N_8614,N_8796);
nand U8899 (N_8899,N_8713,N_8606);
nor U8900 (N_8900,N_8758,N_8763);
or U8901 (N_8901,N_8678,N_8694);
or U8902 (N_8902,N_8701,N_8669);
or U8903 (N_8903,N_8762,N_8602);
and U8904 (N_8904,N_8642,N_8636);
nand U8905 (N_8905,N_8764,N_8748);
or U8906 (N_8906,N_8683,N_8788);
and U8907 (N_8907,N_8677,N_8694);
nand U8908 (N_8908,N_8643,N_8645);
nor U8909 (N_8909,N_8704,N_8772);
nand U8910 (N_8910,N_8785,N_8772);
nor U8911 (N_8911,N_8625,N_8683);
nand U8912 (N_8912,N_8709,N_8626);
or U8913 (N_8913,N_8757,N_8669);
or U8914 (N_8914,N_8679,N_8713);
nand U8915 (N_8915,N_8779,N_8636);
nor U8916 (N_8916,N_8738,N_8696);
nand U8917 (N_8917,N_8748,N_8752);
or U8918 (N_8918,N_8799,N_8637);
nand U8919 (N_8919,N_8745,N_8722);
and U8920 (N_8920,N_8768,N_8764);
nand U8921 (N_8921,N_8659,N_8702);
or U8922 (N_8922,N_8760,N_8785);
and U8923 (N_8923,N_8645,N_8706);
nand U8924 (N_8924,N_8748,N_8673);
and U8925 (N_8925,N_8600,N_8669);
and U8926 (N_8926,N_8772,N_8718);
nor U8927 (N_8927,N_8770,N_8709);
and U8928 (N_8928,N_8658,N_8793);
nand U8929 (N_8929,N_8784,N_8773);
nand U8930 (N_8930,N_8766,N_8742);
nor U8931 (N_8931,N_8794,N_8773);
or U8932 (N_8932,N_8695,N_8732);
nand U8933 (N_8933,N_8635,N_8640);
nor U8934 (N_8934,N_8684,N_8718);
nand U8935 (N_8935,N_8787,N_8662);
nand U8936 (N_8936,N_8753,N_8696);
or U8937 (N_8937,N_8780,N_8684);
and U8938 (N_8938,N_8643,N_8762);
and U8939 (N_8939,N_8762,N_8654);
nor U8940 (N_8940,N_8698,N_8678);
nor U8941 (N_8941,N_8743,N_8638);
and U8942 (N_8942,N_8755,N_8714);
nor U8943 (N_8943,N_8711,N_8648);
or U8944 (N_8944,N_8793,N_8741);
or U8945 (N_8945,N_8612,N_8688);
and U8946 (N_8946,N_8618,N_8613);
and U8947 (N_8947,N_8692,N_8798);
nand U8948 (N_8948,N_8752,N_8695);
or U8949 (N_8949,N_8713,N_8698);
or U8950 (N_8950,N_8742,N_8723);
and U8951 (N_8951,N_8651,N_8699);
nor U8952 (N_8952,N_8655,N_8701);
and U8953 (N_8953,N_8754,N_8785);
and U8954 (N_8954,N_8670,N_8718);
and U8955 (N_8955,N_8605,N_8797);
nand U8956 (N_8956,N_8612,N_8703);
or U8957 (N_8957,N_8746,N_8770);
nand U8958 (N_8958,N_8664,N_8713);
nor U8959 (N_8959,N_8737,N_8750);
and U8960 (N_8960,N_8701,N_8705);
or U8961 (N_8961,N_8635,N_8685);
xor U8962 (N_8962,N_8656,N_8725);
and U8963 (N_8963,N_8643,N_8786);
and U8964 (N_8964,N_8647,N_8730);
or U8965 (N_8965,N_8685,N_8727);
nand U8966 (N_8966,N_8785,N_8681);
or U8967 (N_8967,N_8772,N_8609);
and U8968 (N_8968,N_8706,N_8658);
nor U8969 (N_8969,N_8763,N_8680);
and U8970 (N_8970,N_8781,N_8701);
and U8971 (N_8971,N_8705,N_8713);
and U8972 (N_8972,N_8756,N_8609);
and U8973 (N_8973,N_8791,N_8754);
nor U8974 (N_8974,N_8781,N_8636);
and U8975 (N_8975,N_8769,N_8697);
nand U8976 (N_8976,N_8777,N_8634);
nor U8977 (N_8977,N_8638,N_8709);
nand U8978 (N_8978,N_8633,N_8671);
and U8979 (N_8979,N_8645,N_8750);
or U8980 (N_8980,N_8676,N_8688);
nand U8981 (N_8981,N_8748,N_8656);
or U8982 (N_8982,N_8742,N_8773);
nor U8983 (N_8983,N_8630,N_8731);
and U8984 (N_8984,N_8703,N_8798);
nor U8985 (N_8985,N_8724,N_8663);
and U8986 (N_8986,N_8642,N_8743);
or U8987 (N_8987,N_8648,N_8798);
nand U8988 (N_8988,N_8788,N_8656);
nor U8989 (N_8989,N_8632,N_8639);
nand U8990 (N_8990,N_8756,N_8697);
nand U8991 (N_8991,N_8668,N_8748);
and U8992 (N_8992,N_8741,N_8618);
nand U8993 (N_8993,N_8756,N_8676);
or U8994 (N_8994,N_8726,N_8601);
nand U8995 (N_8995,N_8652,N_8793);
or U8996 (N_8996,N_8745,N_8669);
nand U8997 (N_8997,N_8687,N_8675);
nor U8998 (N_8998,N_8665,N_8725);
and U8999 (N_8999,N_8731,N_8620);
or U9000 (N_9000,N_8874,N_8808);
nor U9001 (N_9001,N_8945,N_8957);
or U9002 (N_9002,N_8895,N_8818);
nand U9003 (N_9003,N_8908,N_8919);
nand U9004 (N_9004,N_8986,N_8865);
or U9005 (N_9005,N_8878,N_8998);
nand U9006 (N_9006,N_8907,N_8880);
nor U9007 (N_9007,N_8964,N_8873);
and U9008 (N_9008,N_8947,N_8830);
or U9009 (N_9009,N_8938,N_8820);
nor U9010 (N_9010,N_8970,N_8926);
nor U9011 (N_9011,N_8955,N_8840);
and U9012 (N_9012,N_8917,N_8891);
or U9013 (N_9013,N_8946,N_8900);
and U9014 (N_9014,N_8927,N_8995);
or U9015 (N_9015,N_8863,N_8897);
nor U9016 (N_9016,N_8975,N_8882);
nand U9017 (N_9017,N_8864,N_8956);
nor U9018 (N_9018,N_8931,N_8949);
and U9019 (N_9019,N_8823,N_8932);
nor U9020 (N_9020,N_8819,N_8839);
and U9021 (N_9021,N_8887,N_8915);
nor U9022 (N_9022,N_8816,N_8904);
and U9023 (N_9023,N_8966,N_8821);
and U9024 (N_9024,N_8834,N_8974);
nand U9025 (N_9025,N_8940,N_8971);
or U9026 (N_9026,N_8868,N_8948);
and U9027 (N_9027,N_8883,N_8866);
and U9028 (N_9028,N_8851,N_8936);
or U9029 (N_9029,N_8937,N_8829);
or U9030 (N_9030,N_8807,N_8871);
nand U9031 (N_9031,N_8824,N_8993);
and U9032 (N_9032,N_8958,N_8858);
nand U9033 (N_9033,N_8811,N_8852);
nor U9034 (N_9034,N_8848,N_8877);
and U9035 (N_9035,N_8916,N_8967);
nor U9036 (N_9036,N_8905,N_8982);
or U9037 (N_9037,N_8875,N_8922);
nor U9038 (N_9038,N_8896,N_8857);
or U9039 (N_9039,N_8827,N_8963);
and U9040 (N_9040,N_8906,N_8861);
and U9041 (N_9041,N_8989,N_8803);
or U9042 (N_9042,N_8968,N_8959);
nand U9043 (N_9043,N_8952,N_8994);
xor U9044 (N_9044,N_8969,N_8845);
or U9045 (N_9045,N_8849,N_8801);
nor U9046 (N_9046,N_8983,N_8941);
and U9047 (N_9047,N_8809,N_8844);
or U9048 (N_9048,N_8996,N_8929);
xnor U9049 (N_9049,N_8961,N_8912);
and U9050 (N_9050,N_8836,N_8889);
or U9051 (N_9051,N_8962,N_8832);
and U9052 (N_9052,N_8859,N_8979);
and U9053 (N_9053,N_8999,N_8997);
or U9054 (N_9054,N_8930,N_8881);
nor U9055 (N_9055,N_8911,N_8856);
or U9056 (N_9056,N_8853,N_8918);
nor U9057 (N_9057,N_8976,N_8893);
or U9058 (N_9058,N_8965,N_8843);
nor U9059 (N_9059,N_8978,N_8953);
nand U9060 (N_9060,N_8847,N_8842);
nand U9061 (N_9061,N_8828,N_8835);
nor U9062 (N_9062,N_8825,N_8909);
xnor U9063 (N_9063,N_8890,N_8888);
nand U9064 (N_9064,N_8972,N_8990);
and U9065 (N_9065,N_8867,N_8870);
and U9066 (N_9066,N_8804,N_8838);
nand U9067 (N_9067,N_8899,N_8901);
nand U9068 (N_9068,N_8923,N_8898);
nand U9069 (N_9069,N_8876,N_8992);
or U9070 (N_9070,N_8850,N_8805);
nor U9071 (N_9071,N_8987,N_8942);
nor U9072 (N_9072,N_8921,N_8988);
nand U9073 (N_9073,N_8831,N_8913);
nand U9074 (N_9074,N_8884,N_8934);
nor U9075 (N_9075,N_8817,N_8892);
or U9076 (N_9076,N_8810,N_8944);
nand U9077 (N_9077,N_8928,N_8939);
nand U9078 (N_9078,N_8862,N_8814);
or U9079 (N_9079,N_8826,N_8885);
and U9080 (N_9080,N_8854,N_8841);
nand U9081 (N_9081,N_8812,N_8935);
nand U9082 (N_9082,N_8879,N_8837);
nand U9083 (N_9083,N_8813,N_8855);
nor U9084 (N_9084,N_8950,N_8860);
nand U9085 (N_9085,N_8872,N_8920);
or U9086 (N_9086,N_8886,N_8985);
nand U9087 (N_9087,N_8802,N_8925);
nor U9088 (N_9088,N_8869,N_8806);
nor U9089 (N_9089,N_8800,N_8943);
nand U9090 (N_9090,N_8894,N_8914);
and U9091 (N_9091,N_8815,N_8910);
nor U9092 (N_9092,N_8980,N_8960);
nor U9093 (N_9093,N_8991,N_8984);
nor U9094 (N_9094,N_8846,N_8954);
or U9095 (N_9095,N_8902,N_8924);
and U9096 (N_9096,N_8822,N_8977);
nand U9097 (N_9097,N_8951,N_8981);
or U9098 (N_9098,N_8973,N_8903);
nand U9099 (N_9099,N_8833,N_8933);
nand U9100 (N_9100,N_8820,N_8956);
or U9101 (N_9101,N_8963,N_8856);
and U9102 (N_9102,N_8979,N_8842);
or U9103 (N_9103,N_8808,N_8920);
and U9104 (N_9104,N_8866,N_8848);
nor U9105 (N_9105,N_8859,N_8944);
nand U9106 (N_9106,N_8864,N_8863);
and U9107 (N_9107,N_8857,N_8893);
and U9108 (N_9108,N_8866,N_8980);
nor U9109 (N_9109,N_8888,N_8923);
nor U9110 (N_9110,N_8851,N_8815);
nor U9111 (N_9111,N_8920,N_8835);
or U9112 (N_9112,N_8904,N_8800);
nor U9113 (N_9113,N_8926,N_8981);
and U9114 (N_9114,N_8846,N_8951);
nor U9115 (N_9115,N_8833,N_8979);
nor U9116 (N_9116,N_8819,N_8856);
nand U9117 (N_9117,N_8805,N_8842);
nand U9118 (N_9118,N_8911,N_8931);
nor U9119 (N_9119,N_8956,N_8830);
or U9120 (N_9120,N_8990,N_8918);
nor U9121 (N_9121,N_8813,N_8990);
or U9122 (N_9122,N_8824,N_8953);
and U9123 (N_9123,N_8950,N_8981);
or U9124 (N_9124,N_8833,N_8950);
nor U9125 (N_9125,N_8888,N_8806);
and U9126 (N_9126,N_8945,N_8892);
or U9127 (N_9127,N_8815,N_8947);
nand U9128 (N_9128,N_8860,N_8920);
and U9129 (N_9129,N_8922,N_8988);
and U9130 (N_9130,N_8923,N_8842);
xnor U9131 (N_9131,N_8878,N_8896);
nand U9132 (N_9132,N_8860,N_8914);
nor U9133 (N_9133,N_8944,N_8849);
nor U9134 (N_9134,N_8899,N_8838);
and U9135 (N_9135,N_8968,N_8931);
nand U9136 (N_9136,N_8869,N_8873);
or U9137 (N_9137,N_8958,N_8942);
or U9138 (N_9138,N_8887,N_8940);
or U9139 (N_9139,N_8894,N_8954);
nand U9140 (N_9140,N_8818,N_8849);
or U9141 (N_9141,N_8850,N_8801);
or U9142 (N_9142,N_8825,N_8861);
and U9143 (N_9143,N_8906,N_8952);
or U9144 (N_9144,N_8847,N_8835);
and U9145 (N_9145,N_8802,N_8948);
nor U9146 (N_9146,N_8802,N_8899);
and U9147 (N_9147,N_8982,N_8808);
or U9148 (N_9148,N_8890,N_8872);
or U9149 (N_9149,N_8858,N_8999);
nand U9150 (N_9150,N_8852,N_8839);
nand U9151 (N_9151,N_8857,N_8842);
nor U9152 (N_9152,N_8973,N_8981);
and U9153 (N_9153,N_8952,N_8933);
and U9154 (N_9154,N_8939,N_8829);
or U9155 (N_9155,N_8925,N_8903);
or U9156 (N_9156,N_8947,N_8865);
or U9157 (N_9157,N_8917,N_8958);
nor U9158 (N_9158,N_8991,N_8923);
and U9159 (N_9159,N_8813,N_8882);
nand U9160 (N_9160,N_8906,N_8800);
or U9161 (N_9161,N_8859,N_8984);
or U9162 (N_9162,N_8969,N_8986);
nor U9163 (N_9163,N_8902,N_8987);
nand U9164 (N_9164,N_8864,N_8823);
and U9165 (N_9165,N_8809,N_8990);
nor U9166 (N_9166,N_8829,N_8992);
nand U9167 (N_9167,N_8990,N_8881);
or U9168 (N_9168,N_8875,N_8854);
and U9169 (N_9169,N_8819,N_8804);
or U9170 (N_9170,N_8876,N_8946);
nor U9171 (N_9171,N_8847,N_8944);
nor U9172 (N_9172,N_8869,N_8904);
and U9173 (N_9173,N_8982,N_8897);
and U9174 (N_9174,N_8890,N_8825);
or U9175 (N_9175,N_8912,N_8862);
nand U9176 (N_9176,N_8922,N_8884);
and U9177 (N_9177,N_8819,N_8906);
or U9178 (N_9178,N_8831,N_8829);
nand U9179 (N_9179,N_8865,N_8980);
or U9180 (N_9180,N_8874,N_8917);
or U9181 (N_9181,N_8905,N_8881);
or U9182 (N_9182,N_8986,N_8813);
nor U9183 (N_9183,N_8941,N_8886);
nor U9184 (N_9184,N_8954,N_8855);
or U9185 (N_9185,N_8816,N_8829);
nand U9186 (N_9186,N_8807,N_8980);
and U9187 (N_9187,N_8904,N_8880);
nand U9188 (N_9188,N_8879,N_8847);
nor U9189 (N_9189,N_8854,N_8962);
or U9190 (N_9190,N_8903,N_8842);
nor U9191 (N_9191,N_8979,N_8877);
and U9192 (N_9192,N_8804,N_8906);
nand U9193 (N_9193,N_8833,N_8909);
nor U9194 (N_9194,N_8997,N_8964);
nor U9195 (N_9195,N_8951,N_8870);
nor U9196 (N_9196,N_8989,N_8931);
nand U9197 (N_9197,N_8823,N_8922);
nor U9198 (N_9198,N_8829,N_8929);
or U9199 (N_9199,N_8863,N_8958);
nand U9200 (N_9200,N_9045,N_9062);
nand U9201 (N_9201,N_9057,N_9084);
nand U9202 (N_9202,N_9108,N_9058);
nand U9203 (N_9203,N_9111,N_9127);
xor U9204 (N_9204,N_9040,N_9077);
or U9205 (N_9205,N_9177,N_9125);
or U9206 (N_9206,N_9104,N_9129);
and U9207 (N_9207,N_9016,N_9001);
and U9208 (N_9208,N_9124,N_9056);
nand U9209 (N_9209,N_9152,N_9014);
nand U9210 (N_9210,N_9054,N_9188);
nor U9211 (N_9211,N_9048,N_9053);
nand U9212 (N_9212,N_9116,N_9128);
nor U9213 (N_9213,N_9191,N_9131);
or U9214 (N_9214,N_9034,N_9146);
and U9215 (N_9215,N_9052,N_9031);
nand U9216 (N_9216,N_9074,N_9066);
nand U9217 (N_9217,N_9165,N_9113);
or U9218 (N_9218,N_9013,N_9081);
nor U9219 (N_9219,N_9130,N_9067);
and U9220 (N_9220,N_9122,N_9163);
and U9221 (N_9221,N_9148,N_9068);
nor U9222 (N_9222,N_9193,N_9162);
nor U9223 (N_9223,N_9190,N_9006);
or U9224 (N_9224,N_9022,N_9147);
nand U9225 (N_9225,N_9123,N_9018);
nand U9226 (N_9226,N_9071,N_9186);
nor U9227 (N_9227,N_9042,N_9106);
nor U9228 (N_9228,N_9174,N_9026);
or U9229 (N_9229,N_9044,N_9118);
and U9230 (N_9230,N_9187,N_9033);
and U9231 (N_9231,N_9010,N_9183);
nor U9232 (N_9232,N_9030,N_9117);
and U9233 (N_9233,N_9095,N_9089);
nand U9234 (N_9234,N_9107,N_9137);
nand U9235 (N_9235,N_9171,N_9141);
nand U9236 (N_9236,N_9098,N_9167);
nand U9237 (N_9237,N_9105,N_9180);
nand U9238 (N_9238,N_9024,N_9020);
or U9239 (N_9239,N_9100,N_9017);
nand U9240 (N_9240,N_9019,N_9173);
or U9241 (N_9241,N_9115,N_9156);
nor U9242 (N_9242,N_9189,N_9132);
and U9243 (N_9243,N_9161,N_9170);
nand U9244 (N_9244,N_9175,N_9027);
or U9245 (N_9245,N_9126,N_9028);
nand U9246 (N_9246,N_9103,N_9009);
or U9247 (N_9247,N_9063,N_9011);
nor U9248 (N_9248,N_9094,N_9178);
and U9249 (N_9249,N_9079,N_9160);
nand U9250 (N_9250,N_9036,N_9060);
nand U9251 (N_9251,N_9075,N_9080);
nor U9252 (N_9252,N_9096,N_9157);
or U9253 (N_9253,N_9166,N_9004);
nand U9254 (N_9254,N_9083,N_9005);
nand U9255 (N_9255,N_9176,N_9000);
nand U9256 (N_9256,N_9002,N_9151);
or U9257 (N_9257,N_9133,N_9172);
nand U9258 (N_9258,N_9097,N_9192);
nand U9259 (N_9259,N_9070,N_9012);
and U9260 (N_9260,N_9155,N_9101);
nand U9261 (N_9261,N_9073,N_9158);
and U9262 (N_9262,N_9032,N_9090);
or U9263 (N_9263,N_9064,N_9196);
or U9264 (N_9264,N_9029,N_9088);
and U9265 (N_9265,N_9076,N_9007);
nor U9266 (N_9266,N_9085,N_9061);
nand U9267 (N_9267,N_9109,N_9069);
and U9268 (N_9268,N_9119,N_9199);
and U9269 (N_9269,N_9185,N_9134);
nand U9270 (N_9270,N_9135,N_9025);
nand U9271 (N_9271,N_9055,N_9149);
nand U9272 (N_9272,N_9037,N_9144);
nand U9273 (N_9273,N_9015,N_9082);
and U9274 (N_9274,N_9121,N_9159);
and U9275 (N_9275,N_9065,N_9091);
nand U9276 (N_9276,N_9182,N_9169);
nand U9277 (N_9277,N_9143,N_9051);
nand U9278 (N_9278,N_9043,N_9049);
and U9279 (N_9279,N_9008,N_9138);
or U9280 (N_9280,N_9145,N_9164);
nand U9281 (N_9281,N_9114,N_9047);
nor U9282 (N_9282,N_9092,N_9140);
and U9283 (N_9283,N_9072,N_9099);
and U9284 (N_9284,N_9154,N_9003);
nor U9285 (N_9285,N_9078,N_9021);
nor U9286 (N_9286,N_9153,N_9102);
and U9287 (N_9287,N_9110,N_9059);
and U9288 (N_9288,N_9038,N_9035);
nand U9289 (N_9289,N_9112,N_9136);
or U9290 (N_9290,N_9195,N_9046);
and U9291 (N_9291,N_9197,N_9086);
nor U9292 (N_9292,N_9093,N_9120);
nor U9293 (N_9293,N_9039,N_9142);
and U9294 (N_9294,N_9168,N_9181);
or U9295 (N_9295,N_9041,N_9198);
and U9296 (N_9296,N_9050,N_9139);
or U9297 (N_9297,N_9087,N_9194);
nand U9298 (N_9298,N_9184,N_9150);
and U9299 (N_9299,N_9023,N_9179);
or U9300 (N_9300,N_9145,N_9118);
or U9301 (N_9301,N_9047,N_9172);
or U9302 (N_9302,N_9115,N_9046);
nand U9303 (N_9303,N_9037,N_9019);
or U9304 (N_9304,N_9051,N_9123);
nand U9305 (N_9305,N_9002,N_9175);
and U9306 (N_9306,N_9123,N_9008);
nand U9307 (N_9307,N_9043,N_9173);
or U9308 (N_9308,N_9130,N_9136);
and U9309 (N_9309,N_9191,N_9068);
xnor U9310 (N_9310,N_9090,N_9049);
nor U9311 (N_9311,N_9071,N_9092);
nand U9312 (N_9312,N_9119,N_9035);
nor U9313 (N_9313,N_9018,N_9110);
or U9314 (N_9314,N_9016,N_9146);
nand U9315 (N_9315,N_9139,N_9092);
and U9316 (N_9316,N_9025,N_9169);
or U9317 (N_9317,N_9025,N_9172);
and U9318 (N_9318,N_9084,N_9179);
or U9319 (N_9319,N_9151,N_9195);
nor U9320 (N_9320,N_9082,N_9148);
nor U9321 (N_9321,N_9099,N_9046);
nand U9322 (N_9322,N_9151,N_9178);
nor U9323 (N_9323,N_9154,N_9098);
nand U9324 (N_9324,N_9116,N_9036);
nand U9325 (N_9325,N_9001,N_9193);
nand U9326 (N_9326,N_9114,N_9031);
and U9327 (N_9327,N_9149,N_9167);
nor U9328 (N_9328,N_9028,N_9161);
nand U9329 (N_9329,N_9031,N_9117);
nor U9330 (N_9330,N_9199,N_9087);
nor U9331 (N_9331,N_9021,N_9127);
and U9332 (N_9332,N_9015,N_9195);
nand U9333 (N_9333,N_9165,N_9138);
xnor U9334 (N_9334,N_9019,N_9001);
and U9335 (N_9335,N_9137,N_9169);
or U9336 (N_9336,N_9154,N_9136);
or U9337 (N_9337,N_9097,N_9115);
nor U9338 (N_9338,N_9102,N_9041);
or U9339 (N_9339,N_9104,N_9135);
and U9340 (N_9340,N_9154,N_9058);
nand U9341 (N_9341,N_9161,N_9097);
and U9342 (N_9342,N_9151,N_9072);
nand U9343 (N_9343,N_9196,N_9032);
or U9344 (N_9344,N_9159,N_9149);
and U9345 (N_9345,N_9152,N_9125);
or U9346 (N_9346,N_9198,N_9025);
or U9347 (N_9347,N_9080,N_9171);
nand U9348 (N_9348,N_9095,N_9137);
or U9349 (N_9349,N_9066,N_9011);
and U9350 (N_9350,N_9158,N_9018);
or U9351 (N_9351,N_9131,N_9082);
and U9352 (N_9352,N_9156,N_9035);
nor U9353 (N_9353,N_9147,N_9049);
or U9354 (N_9354,N_9108,N_9116);
nand U9355 (N_9355,N_9017,N_9049);
or U9356 (N_9356,N_9014,N_9147);
nor U9357 (N_9357,N_9000,N_9033);
xor U9358 (N_9358,N_9024,N_9064);
nand U9359 (N_9359,N_9141,N_9174);
nor U9360 (N_9360,N_9133,N_9064);
and U9361 (N_9361,N_9163,N_9116);
and U9362 (N_9362,N_9095,N_9105);
nor U9363 (N_9363,N_9050,N_9167);
and U9364 (N_9364,N_9114,N_9021);
nor U9365 (N_9365,N_9127,N_9171);
or U9366 (N_9366,N_9145,N_9001);
or U9367 (N_9367,N_9112,N_9128);
or U9368 (N_9368,N_9015,N_9013);
and U9369 (N_9369,N_9138,N_9039);
and U9370 (N_9370,N_9189,N_9062);
nor U9371 (N_9371,N_9134,N_9001);
and U9372 (N_9372,N_9175,N_9006);
nand U9373 (N_9373,N_9199,N_9154);
and U9374 (N_9374,N_9030,N_9003);
nand U9375 (N_9375,N_9197,N_9153);
or U9376 (N_9376,N_9166,N_9052);
nand U9377 (N_9377,N_9101,N_9126);
or U9378 (N_9378,N_9074,N_9079);
nand U9379 (N_9379,N_9151,N_9053);
or U9380 (N_9380,N_9134,N_9152);
or U9381 (N_9381,N_9015,N_9054);
or U9382 (N_9382,N_9000,N_9157);
nand U9383 (N_9383,N_9151,N_9099);
nand U9384 (N_9384,N_9178,N_9040);
nand U9385 (N_9385,N_9023,N_9102);
nand U9386 (N_9386,N_9104,N_9150);
or U9387 (N_9387,N_9095,N_9080);
nand U9388 (N_9388,N_9071,N_9038);
nand U9389 (N_9389,N_9072,N_9131);
nand U9390 (N_9390,N_9081,N_9130);
and U9391 (N_9391,N_9122,N_9041);
and U9392 (N_9392,N_9156,N_9166);
nor U9393 (N_9393,N_9024,N_9120);
nand U9394 (N_9394,N_9075,N_9131);
and U9395 (N_9395,N_9126,N_9157);
nor U9396 (N_9396,N_9150,N_9007);
and U9397 (N_9397,N_9123,N_9094);
and U9398 (N_9398,N_9168,N_9130);
nor U9399 (N_9399,N_9142,N_9068);
nand U9400 (N_9400,N_9322,N_9328);
nor U9401 (N_9401,N_9393,N_9381);
and U9402 (N_9402,N_9334,N_9387);
or U9403 (N_9403,N_9301,N_9292);
nor U9404 (N_9404,N_9361,N_9203);
nor U9405 (N_9405,N_9316,N_9291);
and U9406 (N_9406,N_9308,N_9202);
nand U9407 (N_9407,N_9245,N_9290);
nor U9408 (N_9408,N_9373,N_9293);
nor U9409 (N_9409,N_9214,N_9321);
nor U9410 (N_9410,N_9332,N_9287);
nor U9411 (N_9411,N_9315,N_9377);
or U9412 (N_9412,N_9279,N_9359);
nand U9413 (N_9413,N_9365,N_9216);
xor U9414 (N_9414,N_9337,N_9297);
nor U9415 (N_9415,N_9347,N_9223);
nor U9416 (N_9416,N_9319,N_9336);
and U9417 (N_9417,N_9229,N_9358);
and U9418 (N_9418,N_9272,N_9210);
or U9419 (N_9419,N_9344,N_9305);
nor U9420 (N_9420,N_9271,N_9284);
nand U9421 (N_9421,N_9259,N_9253);
nor U9422 (N_9422,N_9349,N_9234);
nand U9423 (N_9423,N_9302,N_9376);
nor U9424 (N_9424,N_9375,N_9273);
nand U9425 (N_9425,N_9261,N_9274);
nand U9426 (N_9426,N_9383,N_9260);
and U9427 (N_9427,N_9325,N_9209);
or U9428 (N_9428,N_9262,N_9257);
or U9429 (N_9429,N_9395,N_9230);
or U9430 (N_9430,N_9335,N_9220);
or U9431 (N_9431,N_9298,N_9281);
or U9432 (N_9432,N_9314,N_9294);
nor U9433 (N_9433,N_9239,N_9227);
nand U9434 (N_9434,N_9345,N_9283);
and U9435 (N_9435,N_9236,N_9215);
or U9436 (N_9436,N_9277,N_9224);
nor U9437 (N_9437,N_9248,N_9213);
or U9438 (N_9438,N_9382,N_9396);
or U9439 (N_9439,N_9364,N_9226);
or U9440 (N_9440,N_9385,N_9391);
or U9441 (N_9441,N_9235,N_9232);
nand U9442 (N_9442,N_9390,N_9346);
and U9443 (N_9443,N_9266,N_9285);
and U9444 (N_9444,N_9288,N_9366);
nor U9445 (N_9445,N_9369,N_9278);
nand U9446 (N_9446,N_9222,N_9267);
nor U9447 (N_9447,N_9205,N_9249);
or U9448 (N_9448,N_9237,N_9252);
or U9449 (N_9449,N_9217,N_9362);
nand U9450 (N_9450,N_9374,N_9368);
and U9451 (N_9451,N_9331,N_9299);
nand U9452 (N_9452,N_9309,N_9219);
or U9453 (N_9453,N_9221,N_9354);
nor U9454 (N_9454,N_9313,N_9268);
and U9455 (N_9455,N_9351,N_9211);
or U9456 (N_9456,N_9200,N_9339);
nand U9457 (N_9457,N_9247,N_9384);
nor U9458 (N_9458,N_9218,N_9295);
nand U9459 (N_9459,N_9280,N_9356);
nand U9460 (N_9460,N_9386,N_9225);
and U9461 (N_9461,N_9269,N_9353);
nand U9462 (N_9462,N_9348,N_9352);
and U9463 (N_9463,N_9208,N_9324);
and U9464 (N_9464,N_9333,N_9327);
or U9465 (N_9465,N_9378,N_9206);
xnor U9466 (N_9466,N_9398,N_9255);
and U9467 (N_9467,N_9370,N_9242);
and U9468 (N_9468,N_9265,N_9311);
nor U9469 (N_9469,N_9392,N_9289);
and U9470 (N_9470,N_9201,N_9244);
nor U9471 (N_9471,N_9254,N_9355);
nand U9472 (N_9472,N_9300,N_9204);
or U9473 (N_9473,N_9367,N_9304);
or U9474 (N_9474,N_9275,N_9251);
and U9475 (N_9475,N_9212,N_9380);
nand U9476 (N_9476,N_9246,N_9270);
and U9477 (N_9477,N_9397,N_9372);
nor U9478 (N_9478,N_9340,N_9343);
nor U9479 (N_9479,N_9231,N_9310);
nand U9480 (N_9480,N_9329,N_9371);
and U9481 (N_9481,N_9399,N_9233);
or U9482 (N_9482,N_9238,N_9307);
or U9483 (N_9483,N_9389,N_9306);
nor U9484 (N_9484,N_9312,N_9341);
nor U9485 (N_9485,N_9282,N_9241);
and U9486 (N_9486,N_9330,N_9264);
or U9487 (N_9487,N_9388,N_9394);
or U9488 (N_9488,N_9258,N_9323);
or U9489 (N_9489,N_9303,N_9357);
and U9490 (N_9490,N_9250,N_9379);
nor U9491 (N_9491,N_9363,N_9317);
or U9492 (N_9492,N_9286,N_9360);
and U9493 (N_9493,N_9263,N_9320);
nand U9494 (N_9494,N_9276,N_9207);
nand U9495 (N_9495,N_9240,N_9256);
nand U9496 (N_9496,N_9326,N_9296);
nand U9497 (N_9497,N_9318,N_9228);
nand U9498 (N_9498,N_9350,N_9338);
nand U9499 (N_9499,N_9342,N_9243);
and U9500 (N_9500,N_9373,N_9383);
nand U9501 (N_9501,N_9393,N_9286);
nor U9502 (N_9502,N_9221,N_9241);
and U9503 (N_9503,N_9215,N_9268);
and U9504 (N_9504,N_9313,N_9367);
nor U9505 (N_9505,N_9377,N_9384);
nand U9506 (N_9506,N_9320,N_9344);
nor U9507 (N_9507,N_9241,N_9353);
nand U9508 (N_9508,N_9289,N_9352);
or U9509 (N_9509,N_9207,N_9242);
nor U9510 (N_9510,N_9260,N_9305);
and U9511 (N_9511,N_9209,N_9339);
or U9512 (N_9512,N_9354,N_9300);
or U9513 (N_9513,N_9311,N_9301);
and U9514 (N_9514,N_9389,N_9341);
nand U9515 (N_9515,N_9227,N_9389);
or U9516 (N_9516,N_9212,N_9330);
and U9517 (N_9517,N_9319,N_9298);
and U9518 (N_9518,N_9267,N_9231);
and U9519 (N_9519,N_9306,N_9221);
nor U9520 (N_9520,N_9396,N_9231);
and U9521 (N_9521,N_9207,N_9305);
and U9522 (N_9522,N_9339,N_9258);
and U9523 (N_9523,N_9298,N_9211);
nor U9524 (N_9524,N_9355,N_9289);
and U9525 (N_9525,N_9391,N_9316);
and U9526 (N_9526,N_9258,N_9309);
nand U9527 (N_9527,N_9282,N_9222);
and U9528 (N_9528,N_9255,N_9257);
xor U9529 (N_9529,N_9209,N_9235);
and U9530 (N_9530,N_9292,N_9208);
nand U9531 (N_9531,N_9334,N_9221);
nor U9532 (N_9532,N_9394,N_9376);
nand U9533 (N_9533,N_9377,N_9321);
or U9534 (N_9534,N_9270,N_9333);
nand U9535 (N_9535,N_9221,N_9211);
or U9536 (N_9536,N_9259,N_9267);
and U9537 (N_9537,N_9316,N_9285);
nand U9538 (N_9538,N_9218,N_9222);
nand U9539 (N_9539,N_9272,N_9307);
nor U9540 (N_9540,N_9231,N_9243);
or U9541 (N_9541,N_9240,N_9363);
nand U9542 (N_9542,N_9316,N_9237);
and U9543 (N_9543,N_9287,N_9312);
nand U9544 (N_9544,N_9355,N_9250);
nand U9545 (N_9545,N_9349,N_9222);
and U9546 (N_9546,N_9368,N_9340);
nor U9547 (N_9547,N_9348,N_9240);
or U9548 (N_9548,N_9247,N_9394);
nand U9549 (N_9549,N_9204,N_9375);
or U9550 (N_9550,N_9217,N_9343);
and U9551 (N_9551,N_9398,N_9316);
and U9552 (N_9552,N_9316,N_9214);
or U9553 (N_9553,N_9238,N_9351);
or U9554 (N_9554,N_9341,N_9397);
xor U9555 (N_9555,N_9392,N_9394);
and U9556 (N_9556,N_9341,N_9214);
nand U9557 (N_9557,N_9283,N_9294);
or U9558 (N_9558,N_9238,N_9389);
or U9559 (N_9559,N_9346,N_9382);
nand U9560 (N_9560,N_9325,N_9334);
or U9561 (N_9561,N_9396,N_9325);
nand U9562 (N_9562,N_9204,N_9347);
nor U9563 (N_9563,N_9308,N_9318);
and U9564 (N_9564,N_9291,N_9288);
nor U9565 (N_9565,N_9370,N_9289);
nor U9566 (N_9566,N_9369,N_9391);
nor U9567 (N_9567,N_9233,N_9283);
nor U9568 (N_9568,N_9204,N_9224);
nor U9569 (N_9569,N_9340,N_9264);
nand U9570 (N_9570,N_9297,N_9209);
nor U9571 (N_9571,N_9356,N_9378);
nand U9572 (N_9572,N_9373,N_9309);
nand U9573 (N_9573,N_9352,N_9379);
nor U9574 (N_9574,N_9396,N_9324);
or U9575 (N_9575,N_9295,N_9217);
and U9576 (N_9576,N_9321,N_9295);
nand U9577 (N_9577,N_9291,N_9246);
and U9578 (N_9578,N_9282,N_9391);
nand U9579 (N_9579,N_9244,N_9258);
and U9580 (N_9580,N_9296,N_9255);
xnor U9581 (N_9581,N_9284,N_9370);
nor U9582 (N_9582,N_9273,N_9323);
nor U9583 (N_9583,N_9398,N_9226);
or U9584 (N_9584,N_9227,N_9303);
and U9585 (N_9585,N_9253,N_9318);
nand U9586 (N_9586,N_9223,N_9285);
nor U9587 (N_9587,N_9200,N_9229);
or U9588 (N_9588,N_9337,N_9233);
or U9589 (N_9589,N_9371,N_9335);
and U9590 (N_9590,N_9308,N_9394);
and U9591 (N_9591,N_9282,N_9317);
or U9592 (N_9592,N_9289,N_9367);
nand U9593 (N_9593,N_9320,N_9387);
and U9594 (N_9594,N_9389,N_9373);
or U9595 (N_9595,N_9339,N_9309);
or U9596 (N_9596,N_9372,N_9371);
nor U9597 (N_9597,N_9397,N_9322);
nand U9598 (N_9598,N_9340,N_9318);
nand U9599 (N_9599,N_9252,N_9340);
nor U9600 (N_9600,N_9593,N_9556);
nand U9601 (N_9601,N_9517,N_9497);
nand U9602 (N_9602,N_9445,N_9545);
or U9603 (N_9603,N_9540,N_9583);
and U9604 (N_9604,N_9435,N_9594);
or U9605 (N_9605,N_9586,N_9451);
nor U9606 (N_9606,N_9564,N_9483);
and U9607 (N_9607,N_9562,N_9454);
or U9608 (N_9608,N_9405,N_9481);
nor U9609 (N_9609,N_9538,N_9588);
or U9610 (N_9610,N_9459,N_9546);
xnor U9611 (N_9611,N_9541,N_9506);
and U9612 (N_9612,N_9431,N_9470);
nand U9613 (N_9613,N_9407,N_9513);
nand U9614 (N_9614,N_9515,N_9484);
and U9615 (N_9615,N_9507,N_9465);
or U9616 (N_9616,N_9424,N_9569);
nor U9617 (N_9617,N_9462,N_9508);
nand U9618 (N_9618,N_9559,N_9566);
and U9619 (N_9619,N_9539,N_9543);
and U9620 (N_9620,N_9437,N_9574);
or U9621 (N_9621,N_9489,N_9430);
nand U9622 (N_9622,N_9463,N_9477);
nand U9623 (N_9623,N_9487,N_9519);
nor U9624 (N_9624,N_9448,N_9510);
and U9625 (N_9625,N_9478,N_9522);
nor U9626 (N_9626,N_9573,N_9473);
and U9627 (N_9627,N_9422,N_9542);
and U9628 (N_9628,N_9576,N_9469);
or U9629 (N_9629,N_9485,N_9496);
or U9630 (N_9630,N_9499,N_9423);
or U9631 (N_9631,N_9547,N_9450);
and U9632 (N_9632,N_9511,N_9596);
nor U9633 (N_9633,N_9531,N_9549);
nor U9634 (N_9634,N_9417,N_9458);
nor U9635 (N_9635,N_9476,N_9486);
nor U9636 (N_9636,N_9537,N_9408);
nor U9637 (N_9637,N_9429,N_9558);
and U9638 (N_9638,N_9466,N_9460);
or U9639 (N_9639,N_9582,N_9587);
nand U9640 (N_9640,N_9495,N_9548);
and U9641 (N_9641,N_9552,N_9503);
nor U9642 (N_9642,N_9464,N_9500);
or U9643 (N_9643,N_9580,N_9516);
and U9644 (N_9644,N_9472,N_9488);
or U9645 (N_9645,N_9532,N_9453);
nor U9646 (N_9646,N_9468,N_9557);
and U9647 (N_9647,N_9525,N_9493);
or U9648 (N_9648,N_9452,N_9413);
nand U9649 (N_9649,N_9444,N_9425);
and U9650 (N_9650,N_9572,N_9551);
nand U9651 (N_9651,N_9440,N_9482);
and U9652 (N_9652,N_9427,N_9520);
nor U9653 (N_9653,N_9416,N_9599);
and U9654 (N_9654,N_9457,N_9567);
and U9655 (N_9655,N_9560,N_9456);
and U9656 (N_9656,N_9401,N_9432);
or U9657 (N_9657,N_9536,N_9400);
nor U9658 (N_9658,N_9442,N_9404);
nand U9659 (N_9659,N_9480,N_9512);
nand U9660 (N_9660,N_9490,N_9402);
and U9661 (N_9661,N_9589,N_9505);
nor U9662 (N_9662,N_9433,N_9428);
nand U9663 (N_9663,N_9524,N_9535);
or U9664 (N_9664,N_9563,N_9534);
and U9665 (N_9665,N_9578,N_9514);
nor U9666 (N_9666,N_9565,N_9406);
nand U9667 (N_9667,N_9523,N_9509);
nor U9668 (N_9668,N_9530,N_9529);
nor U9669 (N_9669,N_9554,N_9403);
or U9670 (N_9670,N_9434,N_9439);
nand U9671 (N_9671,N_9491,N_9438);
and U9672 (N_9672,N_9555,N_9414);
nor U9673 (N_9673,N_9570,N_9475);
xnor U9674 (N_9674,N_9449,N_9577);
and U9675 (N_9675,N_9411,N_9467);
nor U9676 (N_9676,N_9420,N_9494);
nand U9677 (N_9677,N_9501,N_9591);
nand U9678 (N_9678,N_9441,N_9544);
and U9679 (N_9679,N_9533,N_9597);
nand U9680 (N_9680,N_9579,N_9581);
nand U9681 (N_9681,N_9409,N_9585);
and U9682 (N_9682,N_9592,N_9436);
nand U9683 (N_9683,N_9575,N_9568);
or U9684 (N_9684,N_9415,N_9419);
nor U9685 (N_9685,N_9550,N_9443);
and U9686 (N_9686,N_9561,N_9590);
and U9687 (N_9687,N_9471,N_9446);
nand U9688 (N_9688,N_9598,N_9527);
nand U9689 (N_9689,N_9595,N_9528);
or U9690 (N_9690,N_9455,N_9498);
or U9691 (N_9691,N_9553,N_9410);
and U9692 (N_9692,N_9504,N_9526);
and U9693 (N_9693,N_9418,N_9474);
nor U9694 (N_9694,N_9521,N_9447);
nand U9695 (N_9695,N_9571,N_9421);
or U9696 (N_9696,N_9479,N_9502);
or U9697 (N_9697,N_9426,N_9412);
nor U9698 (N_9698,N_9518,N_9492);
nand U9699 (N_9699,N_9584,N_9461);
nor U9700 (N_9700,N_9497,N_9408);
or U9701 (N_9701,N_9543,N_9500);
and U9702 (N_9702,N_9474,N_9492);
or U9703 (N_9703,N_9559,N_9467);
nor U9704 (N_9704,N_9560,N_9435);
nand U9705 (N_9705,N_9529,N_9426);
or U9706 (N_9706,N_9595,N_9544);
and U9707 (N_9707,N_9436,N_9488);
and U9708 (N_9708,N_9524,N_9515);
and U9709 (N_9709,N_9472,N_9410);
and U9710 (N_9710,N_9466,N_9484);
and U9711 (N_9711,N_9495,N_9468);
nor U9712 (N_9712,N_9439,N_9558);
or U9713 (N_9713,N_9450,N_9406);
or U9714 (N_9714,N_9543,N_9579);
nor U9715 (N_9715,N_9510,N_9570);
and U9716 (N_9716,N_9504,N_9462);
nand U9717 (N_9717,N_9496,N_9575);
nand U9718 (N_9718,N_9540,N_9508);
and U9719 (N_9719,N_9549,N_9596);
nand U9720 (N_9720,N_9469,N_9425);
nor U9721 (N_9721,N_9456,N_9400);
and U9722 (N_9722,N_9531,N_9561);
nand U9723 (N_9723,N_9516,N_9537);
nand U9724 (N_9724,N_9415,N_9405);
nor U9725 (N_9725,N_9553,N_9480);
and U9726 (N_9726,N_9561,N_9540);
nand U9727 (N_9727,N_9419,N_9437);
nand U9728 (N_9728,N_9437,N_9492);
nand U9729 (N_9729,N_9580,N_9573);
nand U9730 (N_9730,N_9481,N_9501);
nand U9731 (N_9731,N_9458,N_9575);
or U9732 (N_9732,N_9424,N_9544);
or U9733 (N_9733,N_9467,N_9475);
or U9734 (N_9734,N_9472,N_9404);
nand U9735 (N_9735,N_9532,N_9462);
nand U9736 (N_9736,N_9513,N_9477);
or U9737 (N_9737,N_9457,N_9498);
nand U9738 (N_9738,N_9483,N_9439);
nand U9739 (N_9739,N_9584,N_9408);
and U9740 (N_9740,N_9551,N_9474);
or U9741 (N_9741,N_9519,N_9401);
or U9742 (N_9742,N_9574,N_9573);
nor U9743 (N_9743,N_9544,N_9505);
nand U9744 (N_9744,N_9459,N_9556);
nor U9745 (N_9745,N_9408,N_9566);
or U9746 (N_9746,N_9417,N_9475);
nand U9747 (N_9747,N_9421,N_9429);
nor U9748 (N_9748,N_9412,N_9421);
and U9749 (N_9749,N_9467,N_9413);
nand U9750 (N_9750,N_9579,N_9422);
and U9751 (N_9751,N_9424,N_9520);
nor U9752 (N_9752,N_9429,N_9439);
nand U9753 (N_9753,N_9574,N_9406);
and U9754 (N_9754,N_9457,N_9465);
or U9755 (N_9755,N_9457,N_9401);
nor U9756 (N_9756,N_9438,N_9520);
nor U9757 (N_9757,N_9577,N_9551);
or U9758 (N_9758,N_9412,N_9460);
and U9759 (N_9759,N_9409,N_9417);
or U9760 (N_9760,N_9510,N_9558);
or U9761 (N_9761,N_9556,N_9515);
or U9762 (N_9762,N_9491,N_9552);
nand U9763 (N_9763,N_9529,N_9489);
and U9764 (N_9764,N_9454,N_9511);
or U9765 (N_9765,N_9592,N_9453);
nand U9766 (N_9766,N_9503,N_9521);
nor U9767 (N_9767,N_9580,N_9538);
nand U9768 (N_9768,N_9587,N_9408);
and U9769 (N_9769,N_9520,N_9590);
or U9770 (N_9770,N_9582,N_9538);
or U9771 (N_9771,N_9586,N_9403);
or U9772 (N_9772,N_9452,N_9465);
or U9773 (N_9773,N_9491,N_9430);
nor U9774 (N_9774,N_9583,N_9492);
nand U9775 (N_9775,N_9448,N_9566);
and U9776 (N_9776,N_9575,N_9418);
and U9777 (N_9777,N_9583,N_9500);
nand U9778 (N_9778,N_9486,N_9589);
or U9779 (N_9779,N_9414,N_9504);
nand U9780 (N_9780,N_9576,N_9539);
or U9781 (N_9781,N_9505,N_9437);
and U9782 (N_9782,N_9404,N_9487);
or U9783 (N_9783,N_9432,N_9581);
nand U9784 (N_9784,N_9510,N_9589);
and U9785 (N_9785,N_9541,N_9513);
nor U9786 (N_9786,N_9537,N_9449);
nand U9787 (N_9787,N_9522,N_9553);
nor U9788 (N_9788,N_9571,N_9436);
or U9789 (N_9789,N_9544,N_9466);
nand U9790 (N_9790,N_9564,N_9462);
nand U9791 (N_9791,N_9583,N_9494);
and U9792 (N_9792,N_9530,N_9444);
nor U9793 (N_9793,N_9548,N_9532);
nor U9794 (N_9794,N_9404,N_9497);
nand U9795 (N_9795,N_9526,N_9452);
nand U9796 (N_9796,N_9574,N_9565);
nor U9797 (N_9797,N_9447,N_9468);
or U9798 (N_9798,N_9568,N_9467);
nor U9799 (N_9799,N_9487,N_9593);
and U9800 (N_9800,N_9784,N_9615);
or U9801 (N_9801,N_9609,N_9690);
nor U9802 (N_9802,N_9691,N_9616);
or U9803 (N_9803,N_9730,N_9606);
xnor U9804 (N_9804,N_9640,N_9694);
nand U9805 (N_9805,N_9758,N_9729);
and U9806 (N_9806,N_9713,N_9761);
and U9807 (N_9807,N_9610,N_9659);
or U9808 (N_9808,N_9663,N_9727);
nand U9809 (N_9809,N_9670,N_9737);
and U9810 (N_9810,N_9642,N_9756);
or U9811 (N_9811,N_9662,N_9604);
nand U9812 (N_9812,N_9620,N_9719);
nor U9813 (N_9813,N_9793,N_9769);
and U9814 (N_9814,N_9652,N_9718);
nand U9815 (N_9815,N_9723,N_9768);
nor U9816 (N_9816,N_9601,N_9708);
and U9817 (N_9817,N_9607,N_9765);
nor U9818 (N_9818,N_9704,N_9676);
nor U9819 (N_9819,N_9752,N_9643);
nand U9820 (N_9820,N_9791,N_9654);
nor U9821 (N_9821,N_9683,N_9753);
nand U9822 (N_9822,N_9754,N_9779);
nand U9823 (N_9823,N_9777,N_9759);
nor U9824 (N_9824,N_9638,N_9760);
nor U9825 (N_9825,N_9655,N_9624);
and U9826 (N_9826,N_9795,N_9798);
or U9827 (N_9827,N_9792,N_9650);
nand U9828 (N_9828,N_9619,N_9693);
or U9829 (N_9829,N_9748,N_9623);
or U9830 (N_9830,N_9614,N_9785);
and U9831 (N_9831,N_9681,N_9608);
nor U9832 (N_9832,N_9660,N_9726);
nand U9833 (N_9833,N_9688,N_9786);
and U9834 (N_9834,N_9771,N_9780);
nand U9835 (N_9835,N_9684,N_9627);
nor U9836 (N_9836,N_9762,N_9665);
and U9837 (N_9837,N_9702,N_9621);
and U9838 (N_9838,N_9757,N_9731);
and U9839 (N_9839,N_9668,N_9772);
nand U9840 (N_9840,N_9618,N_9613);
or U9841 (N_9841,N_9787,N_9799);
or U9842 (N_9842,N_9685,N_9782);
and U9843 (N_9843,N_9695,N_9736);
nand U9844 (N_9844,N_9696,N_9672);
nor U9845 (N_9845,N_9679,N_9766);
and U9846 (N_9846,N_9794,N_9612);
and U9847 (N_9847,N_9639,N_9673);
and U9848 (N_9848,N_9666,N_9686);
nor U9849 (N_9849,N_9721,N_9739);
nor U9850 (N_9850,N_9774,N_9781);
and U9851 (N_9851,N_9667,N_9653);
and U9852 (N_9852,N_9626,N_9743);
or U9853 (N_9853,N_9714,N_9680);
nand U9854 (N_9854,N_9649,N_9617);
nand U9855 (N_9855,N_9622,N_9778);
nand U9856 (N_9856,N_9661,N_9776);
nand U9857 (N_9857,N_9641,N_9755);
and U9858 (N_9858,N_9706,N_9796);
nor U9859 (N_9859,N_9692,N_9633);
nand U9860 (N_9860,N_9751,N_9644);
and U9861 (N_9861,N_9703,N_9605);
or U9862 (N_9862,N_9724,N_9716);
and U9863 (N_9863,N_9750,N_9735);
nor U9864 (N_9864,N_9602,N_9775);
and U9865 (N_9865,N_9677,N_9631);
nor U9866 (N_9866,N_9687,N_9629);
or U9867 (N_9867,N_9797,N_9600);
nand U9868 (N_9868,N_9783,N_9678);
nand U9869 (N_9869,N_9744,N_9669);
or U9870 (N_9870,N_9682,N_9656);
nand U9871 (N_9871,N_9709,N_9749);
and U9872 (N_9872,N_9741,N_9767);
or U9873 (N_9873,N_9764,N_9710);
or U9874 (N_9874,N_9740,N_9658);
and U9875 (N_9875,N_9742,N_9707);
nand U9876 (N_9876,N_9648,N_9711);
and U9877 (N_9877,N_9763,N_9747);
and U9878 (N_9878,N_9717,N_9634);
or U9879 (N_9879,N_9746,N_9603);
nand U9880 (N_9880,N_9732,N_9657);
nor U9881 (N_9881,N_9611,N_9632);
nor U9882 (N_9882,N_9675,N_9705);
or U9883 (N_9883,N_9697,N_9689);
and U9884 (N_9884,N_9630,N_9628);
and U9885 (N_9885,N_9637,N_9664);
and U9886 (N_9886,N_9773,N_9712);
nor U9887 (N_9887,N_9671,N_9645);
or U9888 (N_9888,N_9789,N_9733);
and U9889 (N_9889,N_9700,N_9720);
and U9890 (N_9890,N_9770,N_9722);
and U9891 (N_9891,N_9699,N_9725);
nor U9892 (N_9892,N_9738,N_9636);
or U9893 (N_9893,N_9651,N_9745);
and U9894 (N_9894,N_9674,N_9790);
or U9895 (N_9895,N_9698,N_9701);
nand U9896 (N_9896,N_9625,N_9734);
nand U9897 (N_9897,N_9788,N_9728);
nor U9898 (N_9898,N_9635,N_9647);
nand U9899 (N_9899,N_9715,N_9646);
and U9900 (N_9900,N_9797,N_9792);
or U9901 (N_9901,N_9663,N_9670);
and U9902 (N_9902,N_9627,N_9614);
nand U9903 (N_9903,N_9774,N_9664);
or U9904 (N_9904,N_9742,N_9611);
or U9905 (N_9905,N_9630,N_9676);
nor U9906 (N_9906,N_9690,N_9776);
nand U9907 (N_9907,N_9641,N_9777);
and U9908 (N_9908,N_9763,N_9701);
or U9909 (N_9909,N_9730,N_9628);
or U9910 (N_9910,N_9614,N_9669);
or U9911 (N_9911,N_9607,N_9601);
nand U9912 (N_9912,N_9712,N_9617);
nor U9913 (N_9913,N_9704,N_9702);
nand U9914 (N_9914,N_9747,N_9622);
nand U9915 (N_9915,N_9789,N_9690);
nor U9916 (N_9916,N_9639,N_9670);
nor U9917 (N_9917,N_9774,N_9747);
or U9918 (N_9918,N_9651,N_9664);
nand U9919 (N_9919,N_9699,N_9625);
nand U9920 (N_9920,N_9710,N_9672);
nor U9921 (N_9921,N_9635,N_9724);
nand U9922 (N_9922,N_9636,N_9660);
nor U9923 (N_9923,N_9725,N_9648);
nor U9924 (N_9924,N_9798,N_9775);
nand U9925 (N_9925,N_9612,N_9708);
or U9926 (N_9926,N_9669,N_9676);
nand U9927 (N_9927,N_9792,N_9689);
and U9928 (N_9928,N_9648,N_9729);
or U9929 (N_9929,N_9747,N_9662);
nor U9930 (N_9930,N_9701,N_9640);
or U9931 (N_9931,N_9763,N_9636);
nor U9932 (N_9932,N_9723,N_9629);
and U9933 (N_9933,N_9714,N_9763);
nand U9934 (N_9934,N_9639,N_9782);
and U9935 (N_9935,N_9711,N_9728);
or U9936 (N_9936,N_9787,N_9652);
or U9937 (N_9937,N_9796,N_9720);
or U9938 (N_9938,N_9652,N_9732);
and U9939 (N_9939,N_9732,N_9618);
or U9940 (N_9940,N_9608,N_9719);
nor U9941 (N_9941,N_9725,N_9746);
nor U9942 (N_9942,N_9794,N_9798);
or U9943 (N_9943,N_9710,N_9690);
nand U9944 (N_9944,N_9673,N_9731);
nand U9945 (N_9945,N_9727,N_9697);
xor U9946 (N_9946,N_9684,N_9654);
nor U9947 (N_9947,N_9673,N_9792);
nand U9948 (N_9948,N_9602,N_9660);
or U9949 (N_9949,N_9621,N_9708);
nor U9950 (N_9950,N_9732,N_9603);
nor U9951 (N_9951,N_9606,N_9762);
nor U9952 (N_9952,N_9752,N_9709);
and U9953 (N_9953,N_9702,N_9639);
or U9954 (N_9954,N_9696,N_9764);
and U9955 (N_9955,N_9607,N_9619);
nand U9956 (N_9956,N_9698,N_9679);
nor U9957 (N_9957,N_9656,N_9610);
and U9958 (N_9958,N_9762,N_9648);
or U9959 (N_9959,N_9600,N_9658);
or U9960 (N_9960,N_9744,N_9707);
nand U9961 (N_9961,N_9794,N_9704);
nor U9962 (N_9962,N_9779,N_9765);
or U9963 (N_9963,N_9677,N_9640);
or U9964 (N_9964,N_9611,N_9604);
nand U9965 (N_9965,N_9781,N_9744);
and U9966 (N_9966,N_9635,N_9760);
and U9967 (N_9967,N_9775,N_9690);
nor U9968 (N_9968,N_9617,N_9690);
or U9969 (N_9969,N_9649,N_9731);
nor U9970 (N_9970,N_9790,N_9692);
nor U9971 (N_9971,N_9708,N_9611);
nor U9972 (N_9972,N_9695,N_9649);
or U9973 (N_9973,N_9604,N_9750);
nand U9974 (N_9974,N_9735,N_9747);
and U9975 (N_9975,N_9667,N_9649);
and U9976 (N_9976,N_9664,N_9778);
nor U9977 (N_9977,N_9607,N_9794);
nor U9978 (N_9978,N_9738,N_9606);
or U9979 (N_9979,N_9695,N_9703);
and U9980 (N_9980,N_9786,N_9633);
or U9981 (N_9981,N_9700,N_9748);
or U9982 (N_9982,N_9789,N_9787);
and U9983 (N_9983,N_9643,N_9765);
nand U9984 (N_9984,N_9621,N_9726);
and U9985 (N_9985,N_9713,N_9764);
and U9986 (N_9986,N_9767,N_9665);
or U9987 (N_9987,N_9612,N_9745);
nand U9988 (N_9988,N_9697,N_9752);
nor U9989 (N_9989,N_9655,N_9621);
nand U9990 (N_9990,N_9708,N_9664);
and U9991 (N_9991,N_9717,N_9738);
xnor U9992 (N_9992,N_9623,N_9745);
or U9993 (N_9993,N_9746,N_9722);
or U9994 (N_9994,N_9644,N_9746);
or U9995 (N_9995,N_9609,N_9627);
or U9996 (N_9996,N_9775,N_9720);
and U9997 (N_9997,N_9713,N_9655);
or U9998 (N_9998,N_9710,N_9614);
and U9999 (N_9999,N_9746,N_9606);
or U10000 (N_10000,N_9870,N_9953);
nand U10001 (N_10001,N_9854,N_9993);
nand U10002 (N_10002,N_9852,N_9909);
and U10003 (N_10003,N_9992,N_9869);
and U10004 (N_10004,N_9940,N_9844);
nor U10005 (N_10005,N_9882,N_9866);
nand U10006 (N_10006,N_9919,N_9819);
or U10007 (N_10007,N_9996,N_9979);
nand U10008 (N_10008,N_9937,N_9820);
nor U10009 (N_10009,N_9950,N_9952);
or U10010 (N_10010,N_9803,N_9843);
or U10011 (N_10011,N_9802,N_9850);
nand U10012 (N_10012,N_9838,N_9855);
nor U10013 (N_10013,N_9833,N_9887);
or U10014 (N_10014,N_9834,N_9806);
nor U10015 (N_10015,N_9917,N_9972);
and U10016 (N_10016,N_9967,N_9825);
or U10017 (N_10017,N_9867,N_9921);
and U10018 (N_10018,N_9836,N_9821);
and U10019 (N_10019,N_9824,N_9856);
nor U10020 (N_10020,N_9878,N_9851);
or U10021 (N_10021,N_9975,N_9835);
nor U10022 (N_10022,N_9871,N_9800);
and U10023 (N_10023,N_9899,N_9900);
nor U10024 (N_10024,N_9897,N_9827);
nand U10025 (N_10025,N_9935,N_9970);
nand U10026 (N_10026,N_9942,N_9906);
or U10027 (N_10027,N_9884,N_9894);
and U10028 (N_10028,N_9847,N_9976);
nor U10029 (N_10029,N_9826,N_9808);
nand U10030 (N_10030,N_9896,N_9931);
nand U10031 (N_10031,N_9845,N_9918);
or U10032 (N_10032,N_9971,N_9928);
nand U10033 (N_10033,N_9903,N_9831);
nand U10034 (N_10034,N_9995,N_9859);
or U10035 (N_10035,N_9983,N_9905);
nand U10036 (N_10036,N_9955,N_9927);
or U10037 (N_10037,N_9868,N_9991);
nand U10038 (N_10038,N_9811,N_9832);
nand U10039 (N_10039,N_9924,N_9948);
and U10040 (N_10040,N_9920,N_9912);
nand U10041 (N_10041,N_9916,N_9889);
and U10042 (N_10042,N_9849,N_9857);
or U10043 (N_10043,N_9915,N_9914);
and U10044 (N_10044,N_9997,N_9938);
nand U10045 (N_10045,N_9874,N_9858);
nor U10046 (N_10046,N_9981,N_9960);
or U10047 (N_10047,N_9989,N_9959);
nand U10048 (N_10048,N_9958,N_9977);
nand U10049 (N_10049,N_9933,N_9877);
and U10050 (N_10050,N_9939,N_9923);
nand U10051 (N_10051,N_9886,N_9964);
nand U10052 (N_10052,N_9842,N_9865);
and U10053 (N_10053,N_9898,N_9880);
and U10054 (N_10054,N_9885,N_9986);
nand U10055 (N_10055,N_9980,N_9888);
or U10056 (N_10056,N_9839,N_9812);
or U10057 (N_10057,N_9965,N_9932);
nand U10058 (N_10058,N_9999,N_9837);
nor U10059 (N_10059,N_9973,N_9968);
nor U10060 (N_10060,N_9974,N_9904);
and U10061 (N_10061,N_9985,N_9810);
nor U10062 (N_10062,N_9901,N_9963);
or U10063 (N_10063,N_9817,N_9907);
or U10064 (N_10064,N_9892,N_9881);
nor U10065 (N_10065,N_9998,N_9966);
or U10066 (N_10066,N_9804,N_9818);
and U10067 (N_10067,N_9872,N_9969);
nor U10068 (N_10068,N_9862,N_9864);
nand U10069 (N_10069,N_9944,N_9910);
nand U10070 (N_10070,N_9925,N_9848);
and U10071 (N_10071,N_9809,N_9936);
nand U10072 (N_10072,N_9814,N_9873);
nor U10073 (N_10073,N_9807,N_9891);
or U10074 (N_10074,N_9956,N_9801);
nor U10075 (N_10075,N_9957,N_9853);
and U10076 (N_10076,N_9816,N_9805);
nor U10077 (N_10077,N_9893,N_9941);
and U10078 (N_10078,N_9951,N_9946);
nor U10079 (N_10079,N_9823,N_9954);
and U10080 (N_10080,N_9883,N_9943);
or U10081 (N_10081,N_9913,N_9994);
or U10082 (N_10082,N_9908,N_9829);
and U10083 (N_10083,N_9813,N_9846);
nand U10084 (N_10084,N_9895,N_9902);
nor U10085 (N_10085,N_9990,N_9930);
nor U10086 (N_10086,N_9863,N_9922);
or U10087 (N_10087,N_9840,N_9988);
nand U10088 (N_10088,N_9822,N_9929);
nand U10089 (N_10089,N_9947,N_9945);
and U10090 (N_10090,N_9987,N_9841);
nor U10091 (N_10091,N_9875,N_9876);
nor U10092 (N_10092,N_9830,N_9962);
or U10093 (N_10093,N_9926,N_9984);
nand U10094 (N_10094,N_9879,N_9934);
and U10095 (N_10095,N_9978,N_9861);
nor U10096 (N_10096,N_9961,N_9982);
nand U10097 (N_10097,N_9860,N_9949);
or U10098 (N_10098,N_9815,N_9890);
and U10099 (N_10099,N_9911,N_9828);
or U10100 (N_10100,N_9990,N_9896);
and U10101 (N_10101,N_9916,N_9925);
nor U10102 (N_10102,N_9829,N_9999);
nor U10103 (N_10103,N_9967,N_9810);
or U10104 (N_10104,N_9858,N_9993);
nand U10105 (N_10105,N_9860,N_9925);
nand U10106 (N_10106,N_9838,N_9805);
xor U10107 (N_10107,N_9952,N_9859);
nor U10108 (N_10108,N_9812,N_9882);
nor U10109 (N_10109,N_9865,N_9889);
or U10110 (N_10110,N_9848,N_9880);
and U10111 (N_10111,N_9904,N_9878);
nor U10112 (N_10112,N_9900,N_9802);
and U10113 (N_10113,N_9816,N_9830);
or U10114 (N_10114,N_9898,N_9983);
nor U10115 (N_10115,N_9884,N_9857);
or U10116 (N_10116,N_9881,N_9959);
and U10117 (N_10117,N_9980,N_9905);
or U10118 (N_10118,N_9986,N_9861);
and U10119 (N_10119,N_9849,N_9904);
nor U10120 (N_10120,N_9915,N_9846);
nor U10121 (N_10121,N_9842,N_9838);
or U10122 (N_10122,N_9888,N_9889);
nor U10123 (N_10123,N_9975,N_9969);
or U10124 (N_10124,N_9890,N_9964);
or U10125 (N_10125,N_9879,N_9902);
and U10126 (N_10126,N_9979,N_9963);
nand U10127 (N_10127,N_9816,N_9817);
nand U10128 (N_10128,N_9859,N_9983);
xnor U10129 (N_10129,N_9863,N_9804);
nor U10130 (N_10130,N_9951,N_9992);
or U10131 (N_10131,N_9830,N_9990);
nand U10132 (N_10132,N_9872,N_9954);
nor U10133 (N_10133,N_9958,N_9887);
or U10134 (N_10134,N_9806,N_9821);
nand U10135 (N_10135,N_9912,N_9844);
nor U10136 (N_10136,N_9944,N_9812);
or U10137 (N_10137,N_9896,N_9914);
nand U10138 (N_10138,N_9916,N_9824);
nand U10139 (N_10139,N_9964,N_9871);
nor U10140 (N_10140,N_9994,N_9968);
or U10141 (N_10141,N_9900,N_9984);
and U10142 (N_10142,N_9870,N_9913);
nand U10143 (N_10143,N_9935,N_9836);
nor U10144 (N_10144,N_9866,N_9965);
nand U10145 (N_10145,N_9916,N_9806);
and U10146 (N_10146,N_9905,N_9924);
and U10147 (N_10147,N_9956,N_9989);
nor U10148 (N_10148,N_9902,N_9933);
nand U10149 (N_10149,N_9933,N_9949);
or U10150 (N_10150,N_9822,N_9802);
or U10151 (N_10151,N_9829,N_9978);
nand U10152 (N_10152,N_9949,N_9984);
nor U10153 (N_10153,N_9824,N_9897);
or U10154 (N_10154,N_9838,N_9835);
nand U10155 (N_10155,N_9819,N_9838);
and U10156 (N_10156,N_9953,N_9903);
or U10157 (N_10157,N_9954,N_9936);
or U10158 (N_10158,N_9995,N_9990);
and U10159 (N_10159,N_9839,N_9915);
and U10160 (N_10160,N_9879,N_9811);
or U10161 (N_10161,N_9966,N_9853);
or U10162 (N_10162,N_9902,N_9999);
nor U10163 (N_10163,N_9956,N_9848);
and U10164 (N_10164,N_9966,N_9977);
and U10165 (N_10165,N_9917,N_9994);
or U10166 (N_10166,N_9946,N_9873);
or U10167 (N_10167,N_9818,N_9866);
and U10168 (N_10168,N_9992,N_9828);
nand U10169 (N_10169,N_9912,N_9993);
nand U10170 (N_10170,N_9906,N_9871);
and U10171 (N_10171,N_9819,N_9986);
or U10172 (N_10172,N_9867,N_9969);
or U10173 (N_10173,N_9984,N_9846);
nor U10174 (N_10174,N_9850,N_9939);
nor U10175 (N_10175,N_9971,N_9885);
nand U10176 (N_10176,N_9830,N_9969);
nand U10177 (N_10177,N_9957,N_9921);
nand U10178 (N_10178,N_9928,N_9919);
or U10179 (N_10179,N_9819,N_9821);
nand U10180 (N_10180,N_9834,N_9868);
and U10181 (N_10181,N_9811,N_9911);
nor U10182 (N_10182,N_9807,N_9895);
nor U10183 (N_10183,N_9885,N_9877);
nor U10184 (N_10184,N_9826,N_9917);
or U10185 (N_10185,N_9985,N_9865);
and U10186 (N_10186,N_9951,N_9889);
nor U10187 (N_10187,N_9813,N_9841);
or U10188 (N_10188,N_9829,N_9956);
or U10189 (N_10189,N_9983,N_9952);
nor U10190 (N_10190,N_9814,N_9904);
and U10191 (N_10191,N_9809,N_9941);
nor U10192 (N_10192,N_9830,N_9866);
or U10193 (N_10193,N_9983,N_9881);
and U10194 (N_10194,N_9843,N_9809);
and U10195 (N_10195,N_9867,N_9999);
or U10196 (N_10196,N_9875,N_9874);
xnor U10197 (N_10197,N_9951,N_9846);
or U10198 (N_10198,N_9900,N_9955);
or U10199 (N_10199,N_9881,N_9852);
nand U10200 (N_10200,N_10092,N_10030);
and U10201 (N_10201,N_10158,N_10042);
and U10202 (N_10202,N_10178,N_10033);
and U10203 (N_10203,N_10082,N_10189);
and U10204 (N_10204,N_10125,N_10116);
and U10205 (N_10205,N_10059,N_10155);
xor U10206 (N_10206,N_10071,N_10034);
nor U10207 (N_10207,N_10175,N_10080);
nor U10208 (N_10208,N_10144,N_10131);
and U10209 (N_10209,N_10112,N_10104);
nor U10210 (N_10210,N_10045,N_10078);
nand U10211 (N_10211,N_10090,N_10085);
and U10212 (N_10212,N_10004,N_10013);
or U10213 (N_10213,N_10166,N_10049);
and U10214 (N_10214,N_10063,N_10057);
nor U10215 (N_10215,N_10105,N_10048);
nor U10216 (N_10216,N_10014,N_10086);
nand U10217 (N_10217,N_10024,N_10194);
nand U10218 (N_10218,N_10109,N_10124);
xnor U10219 (N_10219,N_10132,N_10176);
or U10220 (N_10220,N_10142,N_10138);
nand U10221 (N_10221,N_10011,N_10008);
or U10222 (N_10222,N_10182,N_10040);
nand U10223 (N_10223,N_10139,N_10118);
or U10224 (N_10224,N_10198,N_10190);
nand U10225 (N_10225,N_10076,N_10007);
and U10226 (N_10226,N_10153,N_10172);
or U10227 (N_10227,N_10196,N_10121);
and U10228 (N_10228,N_10108,N_10119);
or U10229 (N_10229,N_10136,N_10046);
nand U10230 (N_10230,N_10020,N_10081);
or U10231 (N_10231,N_10152,N_10187);
and U10232 (N_10232,N_10170,N_10157);
nor U10233 (N_10233,N_10101,N_10199);
or U10234 (N_10234,N_10103,N_10114);
and U10235 (N_10235,N_10148,N_10061);
and U10236 (N_10236,N_10140,N_10137);
nor U10237 (N_10237,N_10188,N_10126);
and U10238 (N_10238,N_10097,N_10111);
nor U10239 (N_10239,N_10077,N_10134);
xor U10240 (N_10240,N_10197,N_10066);
nand U10241 (N_10241,N_10089,N_10181);
nor U10242 (N_10242,N_10053,N_10075);
and U10243 (N_10243,N_10120,N_10037);
and U10244 (N_10244,N_10050,N_10123);
or U10245 (N_10245,N_10073,N_10146);
nor U10246 (N_10246,N_10168,N_10010);
and U10247 (N_10247,N_10156,N_10099);
or U10248 (N_10248,N_10151,N_10068);
and U10249 (N_10249,N_10162,N_10160);
and U10250 (N_10250,N_10041,N_10058);
nand U10251 (N_10251,N_10018,N_10193);
or U10252 (N_10252,N_10102,N_10083);
nand U10253 (N_10253,N_10065,N_10022);
and U10254 (N_10254,N_10012,N_10032);
nand U10255 (N_10255,N_10035,N_10016);
and U10256 (N_10256,N_10159,N_10052);
or U10257 (N_10257,N_10147,N_10031);
and U10258 (N_10258,N_10106,N_10130);
nor U10259 (N_10259,N_10186,N_10021);
nand U10260 (N_10260,N_10150,N_10036);
nor U10261 (N_10261,N_10005,N_10173);
or U10262 (N_10262,N_10141,N_10094);
or U10263 (N_10263,N_10143,N_10002);
nand U10264 (N_10264,N_10128,N_10161);
nand U10265 (N_10265,N_10044,N_10110);
and U10266 (N_10266,N_10167,N_10100);
or U10267 (N_10267,N_10184,N_10174);
and U10268 (N_10268,N_10087,N_10093);
and U10269 (N_10269,N_10043,N_10072);
nor U10270 (N_10270,N_10054,N_10169);
nand U10271 (N_10271,N_10095,N_10000);
xor U10272 (N_10272,N_10069,N_10015);
or U10273 (N_10273,N_10183,N_10180);
nor U10274 (N_10274,N_10154,N_10026);
and U10275 (N_10275,N_10165,N_10074);
or U10276 (N_10276,N_10055,N_10113);
nand U10277 (N_10277,N_10019,N_10163);
nor U10278 (N_10278,N_10027,N_10088);
or U10279 (N_10279,N_10122,N_10091);
and U10280 (N_10280,N_10039,N_10164);
nor U10281 (N_10281,N_10115,N_10001);
nor U10282 (N_10282,N_10029,N_10062);
nor U10283 (N_10283,N_10064,N_10133);
and U10284 (N_10284,N_10051,N_10127);
and U10285 (N_10285,N_10195,N_10079);
or U10286 (N_10286,N_10098,N_10006);
and U10287 (N_10287,N_10003,N_10009);
and U10288 (N_10288,N_10070,N_10192);
and U10289 (N_10289,N_10023,N_10117);
nand U10290 (N_10290,N_10107,N_10056);
and U10291 (N_10291,N_10135,N_10025);
and U10292 (N_10292,N_10179,N_10129);
or U10293 (N_10293,N_10177,N_10084);
nand U10294 (N_10294,N_10149,N_10028);
nor U10295 (N_10295,N_10191,N_10171);
nor U10296 (N_10296,N_10047,N_10145);
nor U10297 (N_10297,N_10185,N_10060);
and U10298 (N_10298,N_10067,N_10096);
nand U10299 (N_10299,N_10017,N_10038);
nand U10300 (N_10300,N_10176,N_10074);
nor U10301 (N_10301,N_10151,N_10052);
and U10302 (N_10302,N_10154,N_10092);
or U10303 (N_10303,N_10050,N_10103);
nand U10304 (N_10304,N_10172,N_10026);
nor U10305 (N_10305,N_10061,N_10154);
nand U10306 (N_10306,N_10078,N_10150);
or U10307 (N_10307,N_10196,N_10050);
and U10308 (N_10308,N_10080,N_10143);
nor U10309 (N_10309,N_10138,N_10017);
and U10310 (N_10310,N_10131,N_10160);
nor U10311 (N_10311,N_10008,N_10141);
or U10312 (N_10312,N_10065,N_10094);
nand U10313 (N_10313,N_10108,N_10085);
and U10314 (N_10314,N_10146,N_10182);
nor U10315 (N_10315,N_10033,N_10000);
nand U10316 (N_10316,N_10039,N_10054);
and U10317 (N_10317,N_10004,N_10050);
or U10318 (N_10318,N_10128,N_10060);
and U10319 (N_10319,N_10129,N_10070);
nor U10320 (N_10320,N_10184,N_10191);
or U10321 (N_10321,N_10169,N_10132);
nor U10322 (N_10322,N_10031,N_10065);
nand U10323 (N_10323,N_10134,N_10115);
nand U10324 (N_10324,N_10119,N_10037);
nand U10325 (N_10325,N_10146,N_10134);
nor U10326 (N_10326,N_10142,N_10033);
nor U10327 (N_10327,N_10044,N_10046);
or U10328 (N_10328,N_10049,N_10045);
or U10329 (N_10329,N_10174,N_10004);
nand U10330 (N_10330,N_10152,N_10037);
nor U10331 (N_10331,N_10160,N_10104);
nor U10332 (N_10332,N_10122,N_10130);
nand U10333 (N_10333,N_10194,N_10139);
nand U10334 (N_10334,N_10026,N_10086);
or U10335 (N_10335,N_10112,N_10043);
nor U10336 (N_10336,N_10114,N_10014);
or U10337 (N_10337,N_10146,N_10178);
or U10338 (N_10338,N_10100,N_10001);
nor U10339 (N_10339,N_10189,N_10183);
nand U10340 (N_10340,N_10108,N_10040);
and U10341 (N_10341,N_10112,N_10019);
and U10342 (N_10342,N_10106,N_10192);
or U10343 (N_10343,N_10179,N_10125);
or U10344 (N_10344,N_10047,N_10172);
nor U10345 (N_10345,N_10003,N_10136);
or U10346 (N_10346,N_10047,N_10150);
or U10347 (N_10347,N_10163,N_10122);
and U10348 (N_10348,N_10133,N_10156);
nand U10349 (N_10349,N_10199,N_10123);
nor U10350 (N_10350,N_10046,N_10160);
or U10351 (N_10351,N_10087,N_10094);
xnor U10352 (N_10352,N_10081,N_10034);
or U10353 (N_10353,N_10114,N_10155);
or U10354 (N_10354,N_10037,N_10157);
or U10355 (N_10355,N_10163,N_10080);
or U10356 (N_10356,N_10046,N_10130);
or U10357 (N_10357,N_10051,N_10110);
or U10358 (N_10358,N_10139,N_10135);
or U10359 (N_10359,N_10123,N_10195);
xor U10360 (N_10360,N_10091,N_10186);
nor U10361 (N_10361,N_10197,N_10139);
and U10362 (N_10362,N_10179,N_10043);
and U10363 (N_10363,N_10143,N_10077);
or U10364 (N_10364,N_10095,N_10181);
nor U10365 (N_10365,N_10105,N_10154);
nor U10366 (N_10366,N_10187,N_10029);
nor U10367 (N_10367,N_10104,N_10090);
xor U10368 (N_10368,N_10199,N_10194);
or U10369 (N_10369,N_10014,N_10051);
or U10370 (N_10370,N_10173,N_10011);
or U10371 (N_10371,N_10195,N_10144);
nand U10372 (N_10372,N_10161,N_10010);
nand U10373 (N_10373,N_10180,N_10072);
or U10374 (N_10374,N_10060,N_10015);
nand U10375 (N_10375,N_10176,N_10118);
or U10376 (N_10376,N_10135,N_10042);
nand U10377 (N_10377,N_10078,N_10048);
nor U10378 (N_10378,N_10145,N_10093);
nor U10379 (N_10379,N_10173,N_10169);
xor U10380 (N_10380,N_10146,N_10196);
nor U10381 (N_10381,N_10032,N_10066);
and U10382 (N_10382,N_10034,N_10049);
or U10383 (N_10383,N_10072,N_10151);
nand U10384 (N_10384,N_10036,N_10187);
or U10385 (N_10385,N_10125,N_10016);
nor U10386 (N_10386,N_10112,N_10053);
or U10387 (N_10387,N_10161,N_10048);
nor U10388 (N_10388,N_10084,N_10140);
or U10389 (N_10389,N_10017,N_10078);
nand U10390 (N_10390,N_10046,N_10167);
and U10391 (N_10391,N_10030,N_10122);
or U10392 (N_10392,N_10134,N_10108);
nand U10393 (N_10393,N_10057,N_10070);
or U10394 (N_10394,N_10122,N_10008);
and U10395 (N_10395,N_10113,N_10027);
or U10396 (N_10396,N_10111,N_10086);
nor U10397 (N_10397,N_10006,N_10100);
or U10398 (N_10398,N_10047,N_10085);
nand U10399 (N_10399,N_10169,N_10094);
or U10400 (N_10400,N_10261,N_10231);
or U10401 (N_10401,N_10252,N_10279);
nor U10402 (N_10402,N_10248,N_10313);
nand U10403 (N_10403,N_10256,N_10225);
or U10404 (N_10404,N_10380,N_10298);
or U10405 (N_10405,N_10376,N_10323);
and U10406 (N_10406,N_10227,N_10396);
or U10407 (N_10407,N_10355,N_10278);
nor U10408 (N_10408,N_10300,N_10327);
and U10409 (N_10409,N_10282,N_10251);
or U10410 (N_10410,N_10209,N_10285);
and U10411 (N_10411,N_10254,N_10333);
or U10412 (N_10412,N_10260,N_10301);
and U10413 (N_10413,N_10351,N_10340);
or U10414 (N_10414,N_10360,N_10320);
nor U10415 (N_10415,N_10302,N_10369);
nand U10416 (N_10416,N_10325,N_10318);
nor U10417 (N_10417,N_10284,N_10316);
and U10418 (N_10418,N_10258,N_10264);
or U10419 (N_10419,N_10387,N_10393);
and U10420 (N_10420,N_10224,N_10277);
or U10421 (N_10421,N_10394,N_10346);
or U10422 (N_10422,N_10215,N_10253);
or U10423 (N_10423,N_10353,N_10343);
nand U10424 (N_10424,N_10220,N_10273);
nand U10425 (N_10425,N_10336,N_10200);
and U10426 (N_10426,N_10363,N_10219);
nand U10427 (N_10427,N_10212,N_10237);
or U10428 (N_10428,N_10234,N_10290);
nor U10429 (N_10429,N_10206,N_10372);
or U10430 (N_10430,N_10378,N_10321);
nand U10431 (N_10431,N_10388,N_10330);
or U10432 (N_10432,N_10337,N_10235);
nand U10433 (N_10433,N_10349,N_10335);
nand U10434 (N_10434,N_10203,N_10281);
and U10435 (N_10435,N_10359,N_10356);
or U10436 (N_10436,N_10287,N_10211);
nand U10437 (N_10437,N_10244,N_10345);
nor U10438 (N_10438,N_10391,N_10314);
or U10439 (N_10439,N_10202,N_10247);
and U10440 (N_10440,N_10310,N_10286);
or U10441 (N_10441,N_10241,N_10230);
nor U10442 (N_10442,N_10311,N_10390);
nor U10443 (N_10443,N_10319,N_10271);
nand U10444 (N_10444,N_10332,N_10242);
nor U10445 (N_10445,N_10347,N_10293);
or U10446 (N_10446,N_10386,N_10397);
nand U10447 (N_10447,N_10204,N_10266);
nor U10448 (N_10448,N_10331,N_10341);
nor U10449 (N_10449,N_10317,N_10309);
nor U10450 (N_10450,N_10374,N_10236);
or U10451 (N_10451,N_10348,N_10339);
nor U10452 (N_10452,N_10379,N_10315);
nor U10453 (N_10453,N_10223,N_10299);
and U10454 (N_10454,N_10250,N_10257);
xnor U10455 (N_10455,N_10213,N_10392);
and U10456 (N_10456,N_10322,N_10276);
or U10457 (N_10457,N_10304,N_10226);
xnor U10458 (N_10458,N_10229,N_10305);
or U10459 (N_10459,N_10205,N_10324);
or U10460 (N_10460,N_10344,N_10289);
nand U10461 (N_10461,N_10268,N_10245);
nand U10462 (N_10462,N_10214,N_10246);
nand U10463 (N_10463,N_10269,N_10395);
nand U10464 (N_10464,N_10328,N_10350);
and U10465 (N_10465,N_10207,N_10272);
or U10466 (N_10466,N_10383,N_10361);
or U10467 (N_10467,N_10265,N_10232);
or U10468 (N_10468,N_10294,N_10259);
nand U10469 (N_10469,N_10329,N_10288);
nor U10470 (N_10470,N_10399,N_10297);
nand U10471 (N_10471,N_10275,N_10274);
xor U10472 (N_10472,N_10283,N_10295);
and U10473 (N_10473,N_10240,N_10362);
or U10474 (N_10474,N_10357,N_10389);
nor U10475 (N_10475,N_10267,N_10373);
nand U10476 (N_10476,N_10385,N_10201);
nand U10477 (N_10477,N_10262,N_10210);
nor U10478 (N_10478,N_10217,N_10291);
and U10479 (N_10479,N_10239,N_10370);
and U10480 (N_10480,N_10280,N_10218);
or U10481 (N_10481,N_10384,N_10334);
and U10482 (N_10482,N_10352,N_10382);
nor U10483 (N_10483,N_10255,N_10358);
nor U10484 (N_10484,N_10296,N_10208);
and U10485 (N_10485,N_10375,N_10233);
nor U10486 (N_10486,N_10263,N_10342);
or U10487 (N_10487,N_10308,N_10366);
or U10488 (N_10488,N_10398,N_10238);
or U10489 (N_10489,N_10249,N_10216);
and U10490 (N_10490,N_10222,N_10354);
or U10491 (N_10491,N_10364,N_10326);
or U10492 (N_10492,N_10312,N_10377);
nor U10493 (N_10493,N_10381,N_10306);
nor U10494 (N_10494,N_10270,N_10371);
or U10495 (N_10495,N_10365,N_10307);
nand U10496 (N_10496,N_10292,N_10368);
nand U10497 (N_10497,N_10303,N_10243);
nor U10498 (N_10498,N_10367,N_10221);
nor U10499 (N_10499,N_10338,N_10228);
and U10500 (N_10500,N_10380,N_10211);
nand U10501 (N_10501,N_10358,N_10393);
nand U10502 (N_10502,N_10234,N_10340);
or U10503 (N_10503,N_10233,N_10205);
and U10504 (N_10504,N_10365,N_10227);
nor U10505 (N_10505,N_10387,N_10373);
nand U10506 (N_10506,N_10321,N_10398);
nand U10507 (N_10507,N_10369,N_10330);
and U10508 (N_10508,N_10214,N_10360);
and U10509 (N_10509,N_10238,N_10387);
nand U10510 (N_10510,N_10252,N_10344);
and U10511 (N_10511,N_10329,N_10311);
or U10512 (N_10512,N_10279,N_10231);
or U10513 (N_10513,N_10397,N_10372);
nand U10514 (N_10514,N_10328,N_10352);
nand U10515 (N_10515,N_10328,N_10272);
nand U10516 (N_10516,N_10236,N_10378);
nand U10517 (N_10517,N_10365,N_10388);
or U10518 (N_10518,N_10292,N_10211);
and U10519 (N_10519,N_10207,N_10390);
or U10520 (N_10520,N_10306,N_10352);
and U10521 (N_10521,N_10219,N_10267);
or U10522 (N_10522,N_10300,N_10337);
and U10523 (N_10523,N_10345,N_10239);
nor U10524 (N_10524,N_10204,N_10281);
nand U10525 (N_10525,N_10315,N_10258);
nor U10526 (N_10526,N_10221,N_10349);
or U10527 (N_10527,N_10209,N_10277);
nand U10528 (N_10528,N_10366,N_10365);
nor U10529 (N_10529,N_10220,N_10212);
nand U10530 (N_10530,N_10309,N_10329);
nor U10531 (N_10531,N_10385,N_10248);
nand U10532 (N_10532,N_10359,N_10214);
or U10533 (N_10533,N_10297,N_10395);
nor U10534 (N_10534,N_10294,N_10360);
or U10535 (N_10535,N_10223,N_10281);
and U10536 (N_10536,N_10352,N_10360);
and U10537 (N_10537,N_10315,N_10329);
and U10538 (N_10538,N_10206,N_10283);
and U10539 (N_10539,N_10284,N_10329);
nor U10540 (N_10540,N_10277,N_10300);
or U10541 (N_10541,N_10203,N_10315);
nand U10542 (N_10542,N_10343,N_10328);
nand U10543 (N_10543,N_10238,N_10262);
nor U10544 (N_10544,N_10247,N_10251);
or U10545 (N_10545,N_10262,N_10221);
nor U10546 (N_10546,N_10228,N_10328);
and U10547 (N_10547,N_10334,N_10240);
nor U10548 (N_10548,N_10294,N_10214);
nand U10549 (N_10549,N_10395,N_10205);
and U10550 (N_10550,N_10376,N_10230);
or U10551 (N_10551,N_10262,N_10215);
and U10552 (N_10552,N_10263,N_10208);
nand U10553 (N_10553,N_10361,N_10261);
nor U10554 (N_10554,N_10314,N_10313);
nand U10555 (N_10555,N_10263,N_10382);
and U10556 (N_10556,N_10304,N_10389);
nand U10557 (N_10557,N_10328,N_10258);
nor U10558 (N_10558,N_10307,N_10263);
and U10559 (N_10559,N_10323,N_10251);
nand U10560 (N_10560,N_10285,N_10260);
or U10561 (N_10561,N_10347,N_10282);
xnor U10562 (N_10562,N_10276,N_10399);
and U10563 (N_10563,N_10321,N_10337);
nor U10564 (N_10564,N_10200,N_10203);
nand U10565 (N_10565,N_10237,N_10329);
and U10566 (N_10566,N_10299,N_10222);
nor U10567 (N_10567,N_10221,N_10232);
xor U10568 (N_10568,N_10392,N_10287);
and U10569 (N_10569,N_10286,N_10350);
and U10570 (N_10570,N_10390,N_10357);
and U10571 (N_10571,N_10210,N_10232);
nor U10572 (N_10572,N_10358,N_10215);
or U10573 (N_10573,N_10311,N_10278);
nand U10574 (N_10574,N_10392,N_10343);
and U10575 (N_10575,N_10384,N_10257);
nand U10576 (N_10576,N_10263,N_10361);
and U10577 (N_10577,N_10215,N_10310);
nor U10578 (N_10578,N_10271,N_10336);
and U10579 (N_10579,N_10301,N_10298);
and U10580 (N_10580,N_10397,N_10364);
or U10581 (N_10581,N_10309,N_10283);
nand U10582 (N_10582,N_10273,N_10335);
nor U10583 (N_10583,N_10207,N_10368);
nand U10584 (N_10584,N_10297,N_10206);
nand U10585 (N_10585,N_10332,N_10223);
and U10586 (N_10586,N_10394,N_10367);
or U10587 (N_10587,N_10230,N_10344);
or U10588 (N_10588,N_10257,N_10398);
or U10589 (N_10589,N_10308,N_10335);
and U10590 (N_10590,N_10237,N_10282);
nand U10591 (N_10591,N_10318,N_10348);
and U10592 (N_10592,N_10260,N_10286);
or U10593 (N_10593,N_10279,N_10277);
nor U10594 (N_10594,N_10357,N_10309);
nor U10595 (N_10595,N_10393,N_10272);
or U10596 (N_10596,N_10366,N_10300);
nor U10597 (N_10597,N_10307,N_10257);
or U10598 (N_10598,N_10253,N_10232);
or U10599 (N_10599,N_10397,N_10323);
nand U10600 (N_10600,N_10534,N_10526);
nor U10601 (N_10601,N_10537,N_10566);
nor U10602 (N_10602,N_10422,N_10527);
nor U10603 (N_10603,N_10521,N_10428);
nor U10604 (N_10604,N_10429,N_10555);
and U10605 (N_10605,N_10472,N_10490);
nand U10606 (N_10606,N_10424,N_10467);
and U10607 (N_10607,N_10421,N_10433);
nor U10608 (N_10608,N_10561,N_10582);
nor U10609 (N_10609,N_10468,N_10584);
and U10610 (N_10610,N_10580,N_10516);
or U10611 (N_10611,N_10574,N_10460);
and U10612 (N_10612,N_10571,N_10570);
nor U10613 (N_10613,N_10479,N_10572);
or U10614 (N_10614,N_10585,N_10562);
nand U10615 (N_10615,N_10564,N_10499);
nand U10616 (N_10616,N_10568,N_10418);
and U10617 (N_10617,N_10559,N_10529);
xor U10618 (N_10618,N_10589,N_10423);
nand U10619 (N_10619,N_10547,N_10443);
xor U10620 (N_10620,N_10446,N_10497);
and U10621 (N_10621,N_10553,N_10464);
nor U10622 (N_10622,N_10569,N_10461);
nand U10623 (N_10623,N_10469,N_10451);
or U10624 (N_10624,N_10557,N_10411);
or U10625 (N_10625,N_10520,N_10401);
or U10626 (N_10626,N_10503,N_10427);
nand U10627 (N_10627,N_10415,N_10438);
nand U10628 (N_10628,N_10508,N_10578);
nand U10629 (N_10629,N_10463,N_10481);
nor U10630 (N_10630,N_10533,N_10560);
or U10631 (N_10631,N_10554,N_10471);
nor U10632 (N_10632,N_10437,N_10558);
and U10633 (N_10633,N_10593,N_10539);
nand U10634 (N_10634,N_10549,N_10551);
and U10635 (N_10635,N_10431,N_10483);
nor U10636 (N_10636,N_10514,N_10494);
and U10637 (N_10637,N_10538,N_10500);
or U10638 (N_10638,N_10405,N_10450);
nor U10639 (N_10639,N_10513,N_10439);
or U10640 (N_10640,N_10403,N_10419);
or U10641 (N_10641,N_10583,N_10476);
nand U10642 (N_10642,N_10432,N_10563);
and U10643 (N_10643,N_10542,N_10495);
or U10644 (N_10644,N_10407,N_10496);
or U10645 (N_10645,N_10412,N_10493);
or U10646 (N_10646,N_10525,N_10545);
nor U10647 (N_10647,N_10530,N_10459);
nand U10648 (N_10648,N_10546,N_10440);
and U10649 (N_10649,N_10489,N_10491);
and U10650 (N_10650,N_10409,N_10550);
xnor U10651 (N_10651,N_10591,N_10541);
and U10652 (N_10652,N_10445,N_10596);
or U10653 (N_10653,N_10414,N_10447);
and U10654 (N_10654,N_10532,N_10400);
nor U10655 (N_10655,N_10576,N_10434);
or U10656 (N_10656,N_10404,N_10579);
nand U10657 (N_10657,N_10498,N_10552);
or U10658 (N_10658,N_10473,N_10510);
nor U10659 (N_10659,N_10436,N_10524);
nor U10660 (N_10660,N_10512,N_10456);
and U10661 (N_10661,N_10592,N_10598);
nor U10662 (N_10662,N_10515,N_10453);
or U10663 (N_10663,N_10426,N_10448);
or U10664 (N_10664,N_10502,N_10586);
nand U10665 (N_10665,N_10548,N_10567);
or U10666 (N_10666,N_10581,N_10417);
and U10667 (N_10667,N_10455,N_10402);
and U10668 (N_10668,N_10536,N_10444);
and U10669 (N_10669,N_10588,N_10466);
nand U10670 (N_10670,N_10420,N_10556);
nand U10671 (N_10671,N_10594,N_10597);
or U10672 (N_10672,N_10531,N_10540);
nor U10673 (N_10673,N_10505,N_10577);
nor U10674 (N_10674,N_10482,N_10478);
and U10675 (N_10675,N_10462,N_10458);
nand U10676 (N_10676,N_10406,N_10475);
nand U10677 (N_10677,N_10509,N_10517);
nor U10678 (N_10678,N_10501,N_10507);
and U10679 (N_10679,N_10528,N_10487);
nor U10680 (N_10680,N_10543,N_10523);
nand U10681 (N_10681,N_10484,N_10518);
and U10682 (N_10682,N_10522,N_10416);
nor U10683 (N_10683,N_10544,N_10587);
or U10684 (N_10684,N_10441,N_10590);
and U10685 (N_10685,N_10480,N_10465);
nor U10686 (N_10686,N_10573,N_10485);
or U10687 (N_10687,N_10425,N_10575);
nand U10688 (N_10688,N_10452,N_10506);
nand U10689 (N_10689,N_10457,N_10474);
nor U10690 (N_10690,N_10435,N_10519);
and U10691 (N_10691,N_10408,N_10477);
nand U10692 (N_10692,N_10486,N_10449);
nor U10693 (N_10693,N_10413,N_10599);
and U10694 (N_10694,N_10430,N_10535);
nand U10695 (N_10695,N_10504,N_10595);
and U10696 (N_10696,N_10565,N_10488);
nand U10697 (N_10697,N_10442,N_10454);
and U10698 (N_10698,N_10470,N_10511);
or U10699 (N_10699,N_10410,N_10492);
or U10700 (N_10700,N_10505,N_10506);
nor U10701 (N_10701,N_10512,N_10551);
and U10702 (N_10702,N_10428,N_10543);
nor U10703 (N_10703,N_10427,N_10450);
nor U10704 (N_10704,N_10413,N_10595);
and U10705 (N_10705,N_10466,N_10547);
nand U10706 (N_10706,N_10463,N_10421);
or U10707 (N_10707,N_10453,N_10465);
nor U10708 (N_10708,N_10516,N_10433);
nand U10709 (N_10709,N_10557,N_10527);
and U10710 (N_10710,N_10551,N_10490);
nor U10711 (N_10711,N_10450,N_10463);
and U10712 (N_10712,N_10547,N_10463);
nand U10713 (N_10713,N_10465,N_10473);
or U10714 (N_10714,N_10582,N_10422);
or U10715 (N_10715,N_10460,N_10504);
nand U10716 (N_10716,N_10410,N_10499);
nor U10717 (N_10717,N_10403,N_10526);
or U10718 (N_10718,N_10521,N_10598);
and U10719 (N_10719,N_10458,N_10560);
and U10720 (N_10720,N_10586,N_10576);
nor U10721 (N_10721,N_10528,N_10451);
nand U10722 (N_10722,N_10497,N_10552);
nand U10723 (N_10723,N_10565,N_10520);
nor U10724 (N_10724,N_10412,N_10550);
or U10725 (N_10725,N_10559,N_10579);
and U10726 (N_10726,N_10521,N_10495);
nand U10727 (N_10727,N_10440,N_10587);
and U10728 (N_10728,N_10490,N_10402);
and U10729 (N_10729,N_10599,N_10549);
nor U10730 (N_10730,N_10408,N_10424);
and U10731 (N_10731,N_10503,N_10577);
or U10732 (N_10732,N_10412,N_10467);
or U10733 (N_10733,N_10528,N_10545);
nor U10734 (N_10734,N_10530,N_10442);
nand U10735 (N_10735,N_10496,N_10400);
nand U10736 (N_10736,N_10430,N_10546);
nor U10737 (N_10737,N_10407,N_10522);
nand U10738 (N_10738,N_10570,N_10592);
nor U10739 (N_10739,N_10428,N_10465);
xor U10740 (N_10740,N_10423,N_10537);
nand U10741 (N_10741,N_10596,N_10425);
or U10742 (N_10742,N_10425,N_10584);
or U10743 (N_10743,N_10508,N_10519);
nor U10744 (N_10744,N_10511,N_10437);
nand U10745 (N_10745,N_10400,N_10504);
nor U10746 (N_10746,N_10434,N_10552);
and U10747 (N_10747,N_10550,N_10531);
nand U10748 (N_10748,N_10567,N_10436);
and U10749 (N_10749,N_10421,N_10425);
xor U10750 (N_10750,N_10533,N_10425);
and U10751 (N_10751,N_10599,N_10589);
nor U10752 (N_10752,N_10503,N_10490);
nor U10753 (N_10753,N_10421,N_10445);
nand U10754 (N_10754,N_10455,N_10526);
and U10755 (N_10755,N_10470,N_10456);
or U10756 (N_10756,N_10414,N_10552);
nand U10757 (N_10757,N_10541,N_10494);
and U10758 (N_10758,N_10402,N_10551);
nor U10759 (N_10759,N_10581,N_10516);
nand U10760 (N_10760,N_10523,N_10536);
or U10761 (N_10761,N_10416,N_10420);
or U10762 (N_10762,N_10435,N_10525);
or U10763 (N_10763,N_10449,N_10430);
nor U10764 (N_10764,N_10483,N_10463);
or U10765 (N_10765,N_10422,N_10508);
nor U10766 (N_10766,N_10541,N_10498);
nand U10767 (N_10767,N_10560,N_10546);
or U10768 (N_10768,N_10453,N_10484);
or U10769 (N_10769,N_10591,N_10426);
and U10770 (N_10770,N_10478,N_10538);
and U10771 (N_10771,N_10492,N_10590);
nor U10772 (N_10772,N_10414,N_10497);
and U10773 (N_10773,N_10556,N_10529);
or U10774 (N_10774,N_10527,N_10554);
nor U10775 (N_10775,N_10570,N_10566);
nand U10776 (N_10776,N_10476,N_10462);
nand U10777 (N_10777,N_10404,N_10456);
or U10778 (N_10778,N_10451,N_10464);
and U10779 (N_10779,N_10459,N_10506);
nand U10780 (N_10780,N_10511,N_10577);
xor U10781 (N_10781,N_10593,N_10416);
and U10782 (N_10782,N_10552,N_10429);
and U10783 (N_10783,N_10484,N_10500);
nand U10784 (N_10784,N_10433,N_10500);
nor U10785 (N_10785,N_10509,N_10463);
or U10786 (N_10786,N_10599,N_10488);
nand U10787 (N_10787,N_10429,N_10466);
nand U10788 (N_10788,N_10585,N_10511);
and U10789 (N_10789,N_10499,N_10511);
and U10790 (N_10790,N_10579,N_10505);
nand U10791 (N_10791,N_10518,N_10537);
nor U10792 (N_10792,N_10478,N_10532);
or U10793 (N_10793,N_10428,N_10486);
nand U10794 (N_10794,N_10446,N_10418);
and U10795 (N_10795,N_10585,N_10512);
and U10796 (N_10796,N_10535,N_10543);
nand U10797 (N_10797,N_10440,N_10589);
nand U10798 (N_10798,N_10500,N_10534);
or U10799 (N_10799,N_10531,N_10593);
or U10800 (N_10800,N_10710,N_10699);
nand U10801 (N_10801,N_10733,N_10694);
or U10802 (N_10802,N_10680,N_10655);
nand U10803 (N_10803,N_10610,N_10715);
nand U10804 (N_10804,N_10721,N_10649);
and U10805 (N_10805,N_10614,N_10682);
or U10806 (N_10806,N_10734,N_10609);
or U10807 (N_10807,N_10769,N_10640);
nor U10808 (N_10808,N_10784,N_10653);
and U10809 (N_10809,N_10758,N_10776);
or U10810 (N_10810,N_10661,N_10778);
nor U10811 (N_10811,N_10777,N_10686);
or U10812 (N_10812,N_10623,N_10627);
and U10813 (N_10813,N_10665,N_10743);
and U10814 (N_10814,N_10648,N_10732);
nand U10815 (N_10815,N_10683,N_10727);
nand U10816 (N_10816,N_10621,N_10750);
nand U10817 (N_10817,N_10791,N_10687);
and U10818 (N_10818,N_10774,N_10644);
nand U10819 (N_10819,N_10798,N_10793);
nor U10820 (N_10820,N_10679,N_10681);
and U10821 (N_10821,N_10637,N_10670);
and U10822 (N_10822,N_10735,N_10691);
nand U10823 (N_10823,N_10775,N_10651);
nor U10824 (N_10824,N_10647,N_10722);
nand U10825 (N_10825,N_10783,N_10781);
nor U10826 (N_10826,N_10600,N_10690);
nand U10827 (N_10827,N_10754,N_10708);
and U10828 (N_10828,N_10759,N_10657);
nor U10829 (N_10829,N_10744,N_10730);
or U10830 (N_10830,N_10662,N_10713);
nand U10831 (N_10831,N_10756,N_10605);
nor U10832 (N_10832,N_10671,N_10619);
nand U10833 (N_10833,N_10703,N_10674);
or U10834 (N_10834,N_10630,N_10765);
and U10835 (N_10835,N_10764,N_10705);
nor U10836 (N_10836,N_10712,N_10612);
nor U10837 (N_10837,N_10684,N_10795);
and U10838 (N_10838,N_10745,N_10678);
or U10839 (N_10839,N_10707,N_10771);
nand U10840 (N_10840,N_10689,N_10717);
or U10841 (N_10841,N_10633,N_10692);
or U10842 (N_10842,N_10601,N_10796);
nand U10843 (N_10843,N_10728,N_10632);
and U10844 (N_10844,N_10746,N_10606);
and U10845 (N_10845,N_10654,N_10794);
or U10846 (N_10846,N_10731,N_10740);
nand U10847 (N_10847,N_10659,N_10626);
nand U10848 (N_10848,N_10737,N_10761);
or U10849 (N_10849,N_10716,N_10685);
and U10850 (N_10850,N_10641,N_10663);
nand U10851 (N_10851,N_10669,N_10747);
xor U10852 (N_10852,N_10620,N_10770);
and U10853 (N_10853,N_10782,N_10709);
nor U10854 (N_10854,N_10677,N_10675);
or U10855 (N_10855,N_10676,N_10673);
nor U10856 (N_10856,N_10757,N_10726);
nand U10857 (N_10857,N_10617,N_10650);
and U10858 (N_10858,N_10755,N_10767);
nor U10859 (N_10859,N_10688,N_10636);
or U10860 (N_10860,N_10706,N_10711);
or U10861 (N_10861,N_10719,N_10760);
nand U10862 (N_10862,N_10768,N_10741);
and U10863 (N_10863,N_10656,N_10611);
nor U10864 (N_10864,N_10799,N_10696);
or U10865 (N_10865,N_10664,N_10666);
or U10866 (N_10866,N_10700,N_10652);
and U10867 (N_10867,N_10718,N_10797);
and U10868 (N_10868,N_10748,N_10697);
nand U10869 (N_10869,N_10723,N_10668);
and U10870 (N_10870,N_10660,N_10639);
nand U10871 (N_10871,N_10792,N_10635);
or U10872 (N_10872,N_10702,N_10698);
nand U10873 (N_10873,N_10622,N_10714);
nand U10874 (N_10874,N_10643,N_10729);
nor U10875 (N_10875,N_10602,N_10751);
nand U10876 (N_10876,N_10701,N_10613);
and U10877 (N_10877,N_10608,N_10788);
nor U10878 (N_10878,N_10704,N_10628);
or U10879 (N_10879,N_10780,N_10789);
xnor U10880 (N_10880,N_10629,N_10725);
or U10881 (N_10881,N_10603,N_10753);
and U10882 (N_10882,N_10604,N_10772);
nand U10883 (N_10883,N_10638,N_10739);
and U10884 (N_10884,N_10790,N_10634);
nor U10885 (N_10885,N_10624,N_10645);
or U10886 (N_10886,N_10749,N_10786);
nor U10887 (N_10887,N_10631,N_10724);
or U10888 (N_10888,N_10779,N_10752);
nor U10889 (N_10889,N_10773,N_10763);
or U10890 (N_10890,N_10607,N_10738);
nand U10891 (N_10891,N_10742,N_10787);
nand U10892 (N_10892,N_10618,N_10615);
nand U10893 (N_10893,N_10785,N_10693);
or U10894 (N_10894,N_10736,N_10766);
nand U10895 (N_10895,N_10658,N_10642);
nor U10896 (N_10896,N_10672,N_10616);
or U10897 (N_10897,N_10667,N_10646);
nor U10898 (N_10898,N_10762,N_10625);
nor U10899 (N_10899,N_10720,N_10695);
or U10900 (N_10900,N_10728,N_10667);
nor U10901 (N_10901,N_10713,N_10671);
nand U10902 (N_10902,N_10713,N_10618);
nand U10903 (N_10903,N_10654,N_10662);
nor U10904 (N_10904,N_10782,N_10750);
and U10905 (N_10905,N_10746,N_10786);
and U10906 (N_10906,N_10734,N_10647);
or U10907 (N_10907,N_10796,N_10658);
nand U10908 (N_10908,N_10754,N_10685);
nor U10909 (N_10909,N_10761,N_10699);
or U10910 (N_10910,N_10770,N_10775);
nand U10911 (N_10911,N_10601,N_10775);
nand U10912 (N_10912,N_10684,N_10605);
nand U10913 (N_10913,N_10755,N_10621);
and U10914 (N_10914,N_10602,N_10698);
and U10915 (N_10915,N_10658,N_10728);
or U10916 (N_10916,N_10774,N_10723);
or U10917 (N_10917,N_10765,N_10712);
nor U10918 (N_10918,N_10684,N_10797);
nor U10919 (N_10919,N_10769,N_10647);
nor U10920 (N_10920,N_10613,N_10787);
nand U10921 (N_10921,N_10747,N_10688);
and U10922 (N_10922,N_10690,N_10700);
nand U10923 (N_10923,N_10733,N_10789);
and U10924 (N_10924,N_10733,N_10602);
nor U10925 (N_10925,N_10657,N_10799);
nand U10926 (N_10926,N_10773,N_10718);
nand U10927 (N_10927,N_10624,N_10704);
nor U10928 (N_10928,N_10681,N_10732);
nor U10929 (N_10929,N_10723,N_10780);
nand U10930 (N_10930,N_10609,N_10798);
nand U10931 (N_10931,N_10673,N_10764);
nand U10932 (N_10932,N_10773,N_10791);
and U10933 (N_10933,N_10646,N_10757);
and U10934 (N_10934,N_10746,N_10676);
nand U10935 (N_10935,N_10799,N_10729);
nand U10936 (N_10936,N_10792,N_10747);
nor U10937 (N_10937,N_10618,N_10673);
and U10938 (N_10938,N_10642,N_10649);
or U10939 (N_10939,N_10738,N_10753);
nor U10940 (N_10940,N_10600,N_10676);
and U10941 (N_10941,N_10753,N_10631);
or U10942 (N_10942,N_10707,N_10731);
nand U10943 (N_10943,N_10646,N_10729);
nand U10944 (N_10944,N_10686,N_10610);
nor U10945 (N_10945,N_10662,N_10605);
nor U10946 (N_10946,N_10614,N_10651);
nor U10947 (N_10947,N_10611,N_10639);
or U10948 (N_10948,N_10650,N_10741);
nand U10949 (N_10949,N_10783,N_10718);
nand U10950 (N_10950,N_10783,N_10601);
nand U10951 (N_10951,N_10798,N_10606);
and U10952 (N_10952,N_10638,N_10748);
nand U10953 (N_10953,N_10670,N_10788);
and U10954 (N_10954,N_10674,N_10705);
and U10955 (N_10955,N_10669,N_10758);
nand U10956 (N_10956,N_10606,N_10731);
nor U10957 (N_10957,N_10733,N_10717);
nor U10958 (N_10958,N_10697,N_10703);
nand U10959 (N_10959,N_10718,N_10655);
nand U10960 (N_10960,N_10760,N_10687);
nor U10961 (N_10961,N_10669,N_10790);
or U10962 (N_10962,N_10741,N_10712);
nand U10963 (N_10963,N_10759,N_10605);
nand U10964 (N_10964,N_10724,N_10719);
and U10965 (N_10965,N_10681,N_10692);
and U10966 (N_10966,N_10772,N_10639);
or U10967 (N_10967,N_10621,N_10720);
nand U10968 (N_10968,N_10626,N_10681);
nor U10969 (N_10969,N_10745,N_10719);
or U10970 (N_10970,N_10717,N_10704);
and U10971 (N_10971,N_10661,N_10799);
and U10972 (N_10972,N_10621,N_10784);
or U10973 (N_10973,N_10739,N_10779);
nand U10974 (N_10974,N_10637,N_10678);
and U10975 (N_10975,N_10739,N_10793);
or U10976 (N_10976,N_10757,N_10620);
and U10977 (N_10977,N_10691,N_10767);
and U10978 (N_10978,N_10632,N_10719);
nor U10979 (N_10979,N_10794,N_10715);
nand U10980 (N_10980,N_10749,N_10632);
nand U10981 (N_10981,N_10736,N_10611);
or U10982 (N_10982,N_10744,N_10643);
nand U10983 (N_10983,N_10658,N_10646);
nand U10984 (N_10984,N_10678,N_10622);
or U10985 (N_10985,N_10716,N_10684);
nand U10986 (N_10986,N_10608,N_10615);
nor U10987 (N_10987,N_10783,N_10673);
or U10988 (N_10988,N_10778,N_10615);
and U10989 (N_10989,N_10726,N_10768);
nor U10990 (N_10990,N_10610,N_10709);
and U10991 (N_10991,N_10682,N_10608);
nor U10992 (N_10992,N_10634,N_10648);
nand U10993 (N_10993,N_10750,N_10626);
and U10994 (N_10994,N_10653,N_10788);
nor U10995 (N_10995,N_10680,N_10669);
and U10996 (N_10996,N_10737,N_10753);
nor U10997 (N_10997,N_10603,N_10629);
nand U10998 (N_10998,N_10759,N_10709);
nand U10999 (N_10999,N_10604,N_10780);
xnor U11000 (N_11000,N_10918,N_10961);
and U11001 (N_11001,N_10919,N_10836);
and U11002 (N_11002,N_10986,N_10820);
nor U11003 (N_11003,N_10832,N_10834);
or U11004 (N_11004,N_10937,N_10897);
nor U11005 (N_11005,N_10873,N_10973);
and U11006 (N_11006,N_10946,N_10901);
nand U11007 (N_11007,N_10931,N_10876);
and U11008 (N_11008,N_10940,N_10978);
and U11009 (N_11009,N_10960,N_10968);
and U11010 (N_11010,N_10987,N_10895);
nand U11011 (N_11011,N_10877,N_10809);
nor U11012 (N_11012,N_10813,N_10913);
and U11013 (N_11013,N_10963,N_10842);
and U11014 (N_11014,N_10911,N_10823);
nand U11015 (N_11015,N_10951,N_10972);
nor U11016 (N_11016,N_10852,N_10945);
nand U11017 (N_11017,N_10910,N_10875);
and U11018 (N_11018,N_10824,N_10989);
nor U11019 (N_11019,N_10994,N_10970);
or U11020 (N_11020,N_10983,N_10802);
nand U11021 (N_11021,N_10930,N_10828);
xor U11022 (N_11022,N_10977,N_10953);
nand U11023 (N_11023,N_10835,N_10902);
or U11024 (N_11024,N_10866,N_10925);
and U11025 (N_11025,N_10858,N_10859);
or U11026 (N_11026,N_10964,N_10844);
or U11027 (N_11027,N_10915,N_10906);
nor U11028 (N_11028,N_10984,N_10878);
nand U11029 (N_11029,N_10860,N_10871);
or U11030 (N_11030,N_10991,N_10857);
nand U11031 (N_11031,N_10829,N_10950);
nor U11032 (N_11032,N_10988,N_10889);
nor U11033 (N_11033,N_10868,N_10936);
and U11034 (N_11034,N_10993,N_10803);
and U11035 (N_11035,N_10839,N_10998);
nor U11036 (N_11036,N_10801,N_10800);
nor U11037 (N_11037,N_10971,N_10948);
nand U11038 (N_11038,N_10874,N_10920);
nor U11039 (N_11039,N_10870,N_10849);
or U11040 (N_11040,N_10822,N_10811);
nor U11041 (N_11041,N_10841,N_10976);
nand U11042 (N_11042,N_10872,N_10893);
and U11043 (N_11043,N_10804,N_10947);
nor U11044 (N_11044,N_10838,N_10845);
nand U11045 (N_11045,N_10883,N_10997);
nand U11046 (N_11046,N_10921,N_10982);
or U11047 (N_11047,N_10818,N_10974);
or U11048 (N_11048,N_10958,N_10805);
nand U11049 (N_11049,N_10846,N_10995);
or U11050 (N_11050,N_10938,N_10856);
or U11051 (N_11051,N_10812,N_10851);
nand U11052 (N_11052,N_10882,N_10975);
nand U11053 (N_11053,N_10934,N_10815);
and U11054 (N_11054,N_10904,N_10905);
or U11055 (N_11055,N_10924,N_10810);
nand U11056 (N_11056,N_10955,N_10928);
or U11057 (N_11057,N_10996,N_10854);
and U11058 (N_11058,N_10843,N_10939);
nand U11059 (N_11059,N_10914,N_10985);
or U11060 (N_11060,N_10900,N_10833);
nand U11061 (N_11061,N_10933,N_10855);
nor U11062 (N_11062,N_10819,N_10869);
and U11063 (N_11063,N_10817,N_10808);
nor U11064 (N_11064,N_10980,N_10888);
nand U11065 (N_11065,N_10885,N_10935);
nor U11066 (N_11066,N_10892,N_10965);
nor U11067 (N_11067,N_10912,N_10990);
and U11068 (N_11068,N_10898,N_10816);
and U11069 (N_11069,N_10890,N_10853);
and U11070 (N_11070,N_10848,N_10929);
or U11071 (N_11071,N_10907,N_10899);
or U11072 (N_11072,N_10908,N_10999);
nand U11073 (N_11073,N_10814,N_10957);
xnor U11074 (N_11074,N_10887,N_10992);
xor U11075 (N_11075,N_10837,N_10861);
or U11076 (N_11076,N_10865,N_10850);
nor U11077 (N_11077,N_10922,N_10942);
and U11078 (N_11078,N_10956,N_10969);
or U11079 (N_11079,N_10943,N_10962);
nor U11080 (N_11080,N_10981,N_10831);
and U11081 (N_11081,N_10881,N_10867);
nor U11082 (N_11082,N_10840,N_10880);
or U11083 (N_11083,N_10806,N_10959);
and U11084 (N_11084,N_10894,N_10821);
and U11085 (N_11085,N_10891,N_10909);
or U11086 (N_11086,N_10941,N_10979);
nand U11087 (N_11087,N_10926,N_10917);
nor U11088 (N_11088,N_10923,N_10825);
nand U11089 (N_11089,N_10903,N_10967);
nor U11090 (N_11090,N_10862,N_10884);
nand U11091 (N_11091,N_10927,N_10826);
nand U11092 (N_11092,N_10896,N_10830);
nor U11093 (N_11093,N_10863,N_10944);
nand U11094 (N_11094,N_10966,N_10952);
nand U11095 (N_11095,N_10879,N_10847);
and U11096 (N_11096,N_10932,N_10864);
or U11097 (N_11097,N_10827,N_10807);
nand U11098 (N_11098,N_10954,N_10949);
or U11099 (N_11099,N_10886,N_10916);
nor U11100 (N_11100,N_10987,N_10992);
and U11101 (N_11101,N_10869,N_10914);
nand U11102 (N_11102,N_10959,N_10838);
nor U11103 (N_11103,N_10840,N_10860);
nand U11104 (N_11104,N_10886,N_10973);
nor U11105 (N_11105,N_10925,N_10938);
or U11106 (N_11106,N_10940,N_10814);
nor U11107 (N_11107,N_10964,N_10930);
or U11108 (N_11108,N_10838,N_10938);
or U11109 (N_11109,N_10947,N_10852);
and U11110 (N_11110,N_10920,N_10948);
nor U11111 (N_11111,N_10828,N_10950);
nand U11112 (N_11112,N_10986,N_10844);
and U11113 (N_11113,N_10902,N_10865);
and U11114 (N_11114,N_10869,N_10968);
and U11115 (N_11115,N_10839,N_10951);
or U11116 (N_11116,N_10904,N_10826);
nor U11117 (N_11117,N_10841,N_10844);
and U11118 (N_11118,N_10976,N_10855);
nor U11119 (N_11119,N_10946,N_10855);
xnor U11120 (N_11120,N_10929,N_10905);
nor U11121 (N_11121,N_10832,N_10938);
or U11122 (N_11122,N_10899,N_10933);
nand U11123 (N_11123,N_10951,N_10970);
and U11124 (N_11124,N_10864,N_10927);
and U11125 (N_11125,N_10888,N_10952);
or U11126 (N_11126,N_10988,N_10838);
and U11127 (N_11127,N_10831,N_10921);
or U11128 (N_11128,N_10823,N_10836);
and U11129 (N_11129,N_10915,N_10891);
nor U11130 (N_11130,N_10976,N_10843);
and U11131 (N_11131,N_10889,N_10979);
nand U11132 (N_11132,N_10885,N_10831);
or U11133 (N_11133,N_10832,N_10847);
or U11134 (N_11134,N_10940,N_10822);
nor U11135 (N_11135,N_10810,N_10877);
nand U11136 (N_11136,N_10892,N_10898);
and U11137 (N_11137,N_10850,N_10961);
and U11138 (N_11138,N_10824,N_10972);
and U11139 (N_11139,N_10849,N_10833);
nand U11140 (N_11140,N_10897,N_10869);
nor U11141 (N_11141,N_10868,N_10839);
or U11142 (N_11142,N_10987,N_10971);
and U11143 (N_11143,N_10862,N_10936);
nor U11144 (N_11144,N_10908,N_10846);
nor U11145 (N_11145,N_10910,N_10956);
nand U11146 (N_11146,N_10876,N_10935);
or U11147 (N_11147,N_10932,N_10941);
or U11148 (N_11148,N_10982,N_10899);
or U11149 (N_11149,N_10952,N_10844);
nor U11150 (N_11150,N_10834,N_10930);
nand U11151 (N_11151,N_10954,N_10930);
and U11152 (N_11152,N_10957,N_10993);
nand U11153 (N_11153,N_10852,N_10848);
xnor U11154 (N_11154,N_10819,N_10955);
and U11155 (N_11155,N_10947,N_10967);
nand U11156 (N_11156,N_10981,N_10846);
and U11157 (N_11157,N_10880,N_10827);
and U11158 (N_11158,N_10838,N_10867);
or U11159 (N_11159,N_10805,N_10976);
or U11160 (N_11160,N_10873,N_10969);
nor U11161 (N_11161,N_10998,N_10952);
nor U11162 (N_11162,N_10922,N_10988);
nand U11163 (N_11163,N_10908,N_10879);
nor U11164 (N_11164,N_10839,N_10911);
nor U11165 (N_11165,N_10932,N_10952);
or U11166 (N_11166,N_10878,N_10838);
nand U11167 (N_11167,N_10908,N_10896);
or U11168 (N_11168,N_10841,N_10982);
nor U11169 (N_11169,N_10907,N_10982);
nand U11170 (N_11170,N_10850,N_10915);
or U11171 (N_11171,N_10839,N_10806);
or U11172 (N_11172,N_10959,N_10908);
nand U11173 (N_11173,N_10897,N_10847);
or U11174 (N_11174,N_10810,N_10864);
nor U11175 (N_11175,N_10823,N_10894);
and U11176 (N_11176,N_10801,N_10814);
and U11177 (N_11177,N_10973,N_10802);
and U11178 (N_11178,N_10985,N_10958);
and U11179 (N_11179,N_10942,N_10959);
nand U11180 (N_11180,N_10846,N_10923);
nor U11181 (N_11181,N_10826,N_10852);
or U11182 (N_11182,N_10841,N_10833);
or U11183 (N_11183,N_10956,N_10850);
nand U11184 (N_11184,N_10828,N_10964);
nand U11185 (N_11185,N_10898,N_10842);
nand U11186 (N_11186,N_10945,N_10966);
nor U11187 (N_11187,N_10829,N_10914);
or U11188 (N_11188,N_10918,N_10854);
nor U11189 (N_11189,N_10885,N_10963);
nor U11190 (N_11190,N_10865,N_10818);
nor U11191 (N_11191,N_10875,N_10969);
nand U11192 (N_11192,N_10874,N_10852);
and U11193 (N_11193,N_10907,N_10960);
nor U11194 (N_11194,N_10825,N_10800);
nor U11195 (N_11195,N_10821,N_10850);
or U11196 (N_11196,N_10839,N_10959);
nor U11197 (N_11197,N_10981,N_10960);
or U11198 (N_11198,N_10800,N_10844);
or U11199 (N_11199,N_10963,N_10973);
or U11200 (N_11200,N_11154,N_11019);
nand U11201 (N_11201,N_11073,N_11021);
and U11202 (N_11202,N_11088,N_11065);
and U11203 (N_11203,N_11131,N_11002);
or U11204 (N_11204,N_11053,N_11118);
or U11205 (N_11205,N_11106,N_11020);
or U11206 (N_11206,N_11011,N_11098);
or U11207 (N_11207,N_11103,N_11046);
nand U11208 (N_11208,N_11096,N_11057);
nand U11209 (N_11209,N_11147,N_11105);
nor U11210 (N_11210,N_11100,N_11160);
nand U11211 (N_11211,N_11128,N_11030);
nand U11212 (N_11212,N_11083,N_11061);
nand U11213 (N_11213,N_11171,N_11164);
or U11214 (N_11214,N_11094,N_11024);
nand U11215 (N_11215,N_11185,N_11141);
nor U11216 (N_11216,N_11123,N_11155);
nor U11217 (N_11217,N_11191,N_11133);
and U11218 (N_11218,N_11135,N_11108);
nor U11219 (N_11219,N_11142,N_11091);
nor U11220 (N_11220,N_11013,N_11140);
and U11221 (N_11221,N_11014,N_11104);
nor U11222 (N_11222,N_11107,N_11113);
nand U11223 (N_11223,N_11080,N_11145);
and U11224 (N_11224,N_11033,N_11121);
and U11225 (N_11225,N_11012,N_11006);
or U11226 (N_11226,N_11023,N_11054);
or U11227 (N_11227,N_11127,N_11099);
or U11228 (N_11228,N_11195,N_11028);
nor U11229 (N_11229,N_11178,N_11040);
nand U11230 (N_11230,N_11163,N_11038);
nor U11231 (N_11231,N_11139,N_11007);
and U11232 (N_11232,N_11084,N_11157);
and U11233 (N_11233,N_11044,N_11165);
and U11234 (N_11234,N_11114,N_11159);
or U11235 (N_11235,N_11087,N_11109);
nand U11236 (N_11236,N_11036,N_11072);
and U11237 (N_11237,N_11015,N_11137);
nor U11238 (N_11238,N_11125,N_11052);
nor U11239 (N_11239,N_11049,N_11172);
nand U11240 (N_11240,N_11058,N_11097);
nor U11241 (N_11241,N_11051,N_11003);
nand U11242 (N_11242,N_11018,N_11126);
nand U11243 (N_11243,N_11010,N_11162);
nor U11244 (N_11244,N_11001,N_11188);
nand U11245 (N_11245,N_11166,N_11193);
or U11246 (N_11246,N_11068,N_11170);
and U11247 (N_11247,N_11184,N_11075);
nor U11248 (N_11248,N_11189,N_11136);
and U11249 (N_11249,N_11093,N_11143);
or U11250 (N_11250,N_11000,N_11062);
and U11251 (N_11251,N_11047,N_11064);
nand U11252 (N_11252,N_11196,N_11187);
nand U11253 (N_11253,N_11092,N_11130);
nand U11254 (N_11254,N_11186,N_11041);
nand U11255 (N_11255,N_11070,N_11037);
and U11256 (N_11256,N_11048,N_11176);
and U11257 (N_11257,N_11152,N_11081);
and U11258 (N_11258,N_11161,N_11150);
and U11259 (N_11259,N_11129,N_11056);
nor U11260 (N_11260,N_11032,N_11122);
nor U11261 (N_11261,N_11132,N_11004);
nor U11262 (N_11262,N_11190,N_11034);
or U11263 (N_11263,N_11146,N_11071);
or U11264 (N_11264,N_11095,N_11079);
nor U11265 (N_11265,N_11198,N_11063);
nand U11266 (N_11266,N_11138,N_11144);
or U11267 (N_11267,N_11025,N_11134);
and U11268 (N_11268,N_11115,N_11174);
or U11269 (N_11269,N_11017,N_11008);
and U11270 (N_11270,N_11060,N_11101);
and U11271 (N_11271,N_11177,N_11055);
nor U11272 (N_11272,N_11005,N_11117);
or U11273 (N_11273,N_11066,N_11149);
and U11274 (N_11274,N_11085,N_11182);
nand U11275 (N_11275,N_11175,N_11027);
nor U11276 (N_11276,N_11077,N_11169);
and U11277 (N_11277,N_11045,N_11090);
or U11278 (N_11278,N_11120,N_11086);
xnor U11279 (N_11279,N_11031,N_11111);
nor U11280 (N_11280,N_11059,N_11043);
nand U11281 (N_11281,N_11042,N_11116);
nand U11282 (N_11282,N_11158,N_11148);
nor U11283 (N_11283,N_11089,N_11074);
or U11284 (N_11284,N_11076,N_11039);
or U11285 (N_11285,N_11151,N_11173);
nor U11286 (N_11286,N_11156,N_11112);
and U11287 (N_11287,N_11029,N_11102);
and U11288 (N_11288,N_11197,N_11022);
nand U11289 (N_11289,N_11181,N_11016);
nor U11290 (N_11290,N_11035,N_11180);
and U11291 (N_11291,N_11168,N_11069);
nand U11292 (N_11292,N_11194,N_11119);
nand U11293 (N_11293,N_11153,N_11179);
and U11294 (N_11294,N_11082,N_11124);
nand U11295 (N_11295,N_11050,N_11110);
nand U11296 (N_11296,N_11078,N_11192);
or U11297 (N_11297,N_11067,N_11183);
and U11298 (N_11298,N_11026,N_11009);
nand U11299 (N_11299,N_11167,N_11199);
nor U11300 (N_11300,N_11059,N_11086);
or U11301 (N_11301,N_11191,N_11090);
or U11302 (N_11302,N_11144,N_11019);
or U11303 (N_11303,N_11029,N_11003);
or U11304 (N_11304,N_11181,N_11073);
nand U11305 (N_11305,N_11129,N_11088);
or U11306 (N_11306,N_11070,N_11014);
nand U11307 (N_11307,N_11081,N_11190);
nand U11308 (N_11308,N_11016,N_11023);
nand U11309 (N_11309,N_11173,N_11056);
nand U11310 (N_11310,N_11125,N_11104);
or U11311 (N_11311,N_11147,N_11139);
or U11312 (N_11312,N_11002,N_11160);
and U11313 (N_11313,N_11126,N_11077);
nand U11314 (N_11314,N_11177,N_11008);
nand U11315 (N_11315,N_11134,N_11015);
nand U11316 (N_11316,N_11160,N_11120);
and U11317 (N_11317,N_11108,N_11050);
and U11318 (N_11318,N_11129,N_11004);
and U11319 (N_11319,N_11013,N_11147);
or U11320 (N_11320,N_11095,N_11121);
and U11321 (N_11321,N_11006,N_11192);
or U11322 (N_11322,N_11029,N_11135);
or U11323 (N_11323,N_11105,N_11050);
and U11324 (N_11324,N_11030,N_11165);
and U11325 (N_11325,N_11120,N_11094);
or U11326 (N_11326,N_11001,N_11185);
nand U11327 (N_11327,N_11113,N_11194);
and U11328 (N_11328,N_11066,N_11003);
and U11329 (N_11329,N_11072,N_11066);
and U11330 (N_11330,N_11118,N_11068);
or U11331 (N_11331,N_11182,N_11134);
and U11332 (N_11332,N_11017,N_11072);
nand U11333 (N_11333,N_11107,N_11061);
nor U11334 (N_11334,N_11032,N_11082);
nand U11335 (N_11335,N_11028,N_11196);
nor U11336 (N_11336,N_11057,N_11134);
or U11337 (N_11337,N_11131,N_11033);
nand U11338 (N_11338,N_11162,N_11047);
nand U11339 (N_11339,N_11117,N_11180);
nor U11340 (N_11340,N_11191,N_11127);
or U11341 (N_11341,N_11008,N_11100);
or U11342 (N_11342,N_11197,N_11185);
nor U11343 (N_11343,N_11137,N_11154);
nor U11344 (N_11344,N_11137,N_11063);
nand U11345 (N_11345,N_11010,N_11161);
and U11346 (N_11346,N_11094,N_11096);
or U11347 (N_11347,N_11052,N_11005);
and U11348 (N_11348,N_11019,N_11032);
nor U11349 (N_11349,N_11141,N_11045);
and U11350 (N_11350,N_11001,N_11150);
and U11351 (N_11351,N_11028,N_11072);
or U11352 (N_11352,N_11194,N_11186);
nand U11353 (N_11353,N_11064,N_11058);
or U11354 (N_11354,N_11045,N_11162);
nor U11355 (N_11355,N_11125,N_11051);
or U11356 (N_11356,N_11060,N_11125);
and U11357 (N_11357,N_11184,N_11159);
nand U11358 (N_11358,N_11104,N_11042);
nor U11359 (N_11359,N_11133,N_11109);
or U11360 (N_11360,N_11068,N_11143);
and U11361 (N_11361,N_11075,N_11139);
nor U11362 (N_11362,N_11159,N_11004);
or U11363 (N_11363,N_11023,N_11065);
nand U11364 (N_11364,N_11176,N_11011);
nor U11365 (N_11365,N_11198,N_11141);
nor U11366 (N_11366,N_11004,N_11036);
nor U11367 (N_11367,N_11049,N_11018);
nor U11368 (N_11368,N_11187,N_11106);
xnor U11369 (N_11369,N_11082,N_11075);
nor U11370 (N_11370,N_11080,N_11002);
nor U11371 (N_11371,N_11090,N_11193);
or U11372 (N_11372,N_11060,N_11027);
nor U11373 (N_11373,N_11125,N_11094);
or U11374 (N_11374,N_11136,N_11124);
nand U11375 (N_11375,N_11149,N_11116);
nand U11376 (N_11376,N_11031,N_11054);
and U11377 (N_11377,N_11057,N_11018);
nand U11378 (N_11378,N_11180,N_11186);
nand U11379 (N_11379,N_11020,N_11152);
or U11380 (N_11380,N_11189,N_11115);
and U11381 (N_11381,N_11073,N_11198);
or U11382 (N_11382,N_11033,N_11082);
xnor U11383 (N_11383,N_11077,N_11007);
or U11384 (N_11384,N_11181,N_11011);
and U11385 (N_11385,N_11020,N_11030);
nor U11386 (N_11386,N_11035,N_11094);
nand U11387 (N_11387,N_11105,N_11144);
or U11388 (N_11388,N_11048,N_11001);
nand U11389 (N_11389,N_11078,N_11163);
or U11390 (N_11390,N_11115,N_11000);
and U11391 (N_11391,N_11095,N_11007);
or U11392 (N_11392,N_11058,N_11187);
or U11393 (N_11393,N_11195,N_11123);
nor U11394 (N_11394,N_11096,N_11051);
nor U11395 (N_11395,N_11158,N_11035);
nor U11396 (N_11396,N_11078,N_11184);
nor U11397 (N_11397,N_11089,N_11175);
nand U11398 (N_11398,N_11098,N_11014);
and U11399 (N_11399,N_11041,N_11076);
nand U11400 (N_11400,N_11311,N_11331);
or U11401 (N_11401,N_11249,N_11306);
nor U11402 (N_11402,N_11234,N_11358);
nand U11403 (N_11403,N_11394,N_11377);
and U11404 (N_11404,N_11239,N_11271);
nor U11405 (N_11405,N_11285,N_11359);
nor U11406 (N_11406,N_11215,N_11382);
nor U11407 (N_11407,N_11204,N_11373);
nor U11408 (N_11408,N_11381,N_11242);
nand U11409 (N_11409,N_11371,N_11384);
nand U11410 (N_11410,N_11240,N_11360);
nor U11411 (N_11411,N_11224,N_11289);
and U11412 (N_11412,N_11319,N_11262);
nand U11413 (N_11413,N_11243,N_11222);
or U11414 (N_11414,N_11304,N_11313);
and U11415 (N_11415,N_11203,N_11366);
or U11416 (N_11416,N_11380,N_11277);
nand U11417 (N_11417,N_11205,N_11374);
or U11418 (N_11418,N_11323,N_11322);
or U11419 (N_11419,N_11219,N_11300);
nor U11420 (N_11420,N_11303,N_11282);
or U11421 (N_11421,N_11307,N_11387);
nor U11422 (N_11422,N_11353,N_11356);
nand U11423 (N_11423,N_11274,N_11390);
or U11424 (N_11424,N_11372,N_11361);
and U11425 (N_11425,N_11352,N_11317);
nand U11426 (N_11426,N_11370,N_11218);
nor U11427 (N_11427,N_11325,N_11299);
nor U11428 (N_11428,N_11241,N_11276);
nand U11429 (N_11429,N_11367,N_11298);
nor U11430 (N_11430,N_11265,N_11320);
nand U11431 (N_11431,N_11208,N_11255);
or U11432 (N_11432,N_11201,N_11260);
or U11433 (N_11433,N_11258,N_11312);
and U11434 (N_11434,N_11268,N_11297);
nand U11435 (N_11435,N_11308,N_11330);
nor U11436 (N_11436,N_11273,N_11348);
nand U11437 (N_11437,N_11229,N_11388);
nand U11438 (N_11438,N_11280,N_11291);
nor U11439 (N_11439,N_11364,N_11264);
and U11440 (N_11440,N_11259,N_11252);
nor U11441 (N_11441,N_11345,N_11346);
xnor U11442 (N_11442,N_11376,N_11335);
xnor U11443 (N_11443,N_11396,N_11324);
nor U11444 (N_11444,N_11263,N_11232);
and U11445 (N_11445,N_11327,N_11290);
nor U11446 (N_11446,N_11309,N_11275);
or U11447 (N_11447,N_11278,N_11214);
and U11448 (N_11448,N_11340,N_11270);
or U11449 (N_11449,N_11216,N_11246);
and U11450 (N_11450,N_11294,N_11314);
nand U11451 (N_11451,N_11237,N_11329);
or U11452 (N_11452,N_11233,N_11302);
nand U11453 (N_11453,N_11293,N_11339);
nand U11454 (N_11454,N_11379,N_11343);
or U11455 (N_11455,N_11207,N_11230);
nand U11456 (N_11456,N_11391,N_11389);
nand U11457 (N_11457,N_11206,N_11213);
or U11458 (N_11458,N_11288,N_11200);
and U11459 (N_11459,N_11235,N_11223);
and U11460 (N_11460,N_11333,N_11338);
nand U11461 (N_11461,N_11281,N_11315);
and U11462 (N_11462,N_11256,N_11254);
nor U11463 (N_11463,N_11395,N_11245);
or U11464 (N_11464,N_11261,N_11383);
or U11465 (N_11465,N_11301,N_11226);
or U11466 (N_11466,N_11267,N_11357);
nand U11467 (N_11467,N_11272,N_11266);
nand U11468 (N_11468,N_11368,N_11250);
nor U11469 (N_11469,N_11210,N_11362);
nand U11470 (N_11470,N_11354,N_11296);
nor U11471 (N_11471,N_11209,N_11221);
nand U11472 (N_11472,N_11283,N_11347);
nand U11473 (N_11473,N_11295,N_11217);
and U11474 (N_11474,N_11326,N_11292);
nor U11475 (N_11475,N_11344,N_11341);
nor U11476 (N_11476,N_11231,N_11202);
nand U11477 (N_11477,N_11316,N_11211);
xnor U11478 (N_11478,N_11378,N_11385);
nor U11479 (N_11479,N_11251,N_11337);
or U11480 (N_11480,N_11392,N_11318);
and U11481 (N_11481,N_11397,N_11399);
or U11482 (N_11482,N_11247,N_11284);
nor U11483 (N_11483,N_11269,N_11393);
or U11484 (N_11484,N_11279,N_11365);
nor U11485 (N_11485,N_11342,N_11257);
and U11486 (N_11486,N_11349,N_11369);
nor U11487 (N_11487,N_11355,N_11212);
or U11488 (N_11488,N_11287,N_11386);
nand U11489 (N_11489,N_11363,N_11228);
nand U11490 (N_11490,N_11305,N_11238);
and U11491 (N_11491,N_11236,N_11336);
nand U11492 (N_11492,N_11248,N_11351);
nor U11493 (N_11493,N_11244,N_11328);
nand U11494 (N_11494,N_11398,N_11334);
nor U11495 (N_11495,N_11220,N_11253);
and U11496 (N_11496,N_11286,N_11227);
or U11497 (N_11497,N_11225,N_11310);
nand U11498 (N_11498,N_11321,N_11350);
nor U11499 (N_11499,N_11332,N_11375);
nand U11500 (N_11500,N_11363,N_11319);
nor U11501 (N_11501,N_11316,N_11356);
nand U11502 (N_11502,N_11229,N_11379);
or U11503 (N_11503,N_11297,N_11272);
nor U11504 (N_11504,N_11389,N_11301);
nand U11505 (N_11505,N_11390,N_11346);
and U11506 (N_11506,N_11276,N_11238);
nor U11507 (N_11507,N_11201,N_11204);
nor U11508 (N_11508,N_11259,N_11210);
nor U11509 (N_11509,N_11371,N_11312);
nor U11510 (N_11510,N_11330,N_11290);
nor U11511 (N_11511,N_11231,N_11267);
or U11512 (N_11512,N_11269,N_11253);
or U11513 (N_11513,N_11386,N_11282);
nand U11514 (N_11514,N_11264,N_11311);
or U11515 (N_11515,N_11251,N_11275);
nor U11516 (N_11516,N_11312,N_11216);
nor U11517 (N_11517,N_11323,N_11338);
and U11518 (N_11518,N_11223,N_11236);
or U11519 (N_11519,N_11299,N_11394);
nor U11520 (N_11520,N_11371,N_11256);
or U11521 (N_11521,N_11250,N_11201);
and U11522 (N_11522,N_11223,N_11233);
nand U11523 (N_11523,N_11343,N_11251);
and U11524 (N_11524,N_11339,N_11328);
nand U11525 (N_11525,N_11281,N_11267);
nor U11526 (N_11526,N_11228,N_11235);
or U11527 (N_11527,N_11318,N_11231);
or U11528 (N_11528,N_11227,N_11209);
nor U11529 (N_11529,N_11339,N_11291);
and U11530 (N_11530,N_11210,N_11367);
or U11531 (N_11531,N_11304,N_11327);
and U11532 (N_11532,N_11215,N_11238);
and U11533 (N_11533,N_11392,N_11336);
nor U11534 (N_11534,N_11258,N_11271);
or U11535 (N_11535,N_11242,N_11209);
or U11536 (N_11536,N_11206,N_11296);
nor U11537 (N_11537,N_11270,N_11336);
and U11538 (N_11538,N_11206,N_11328);
and U11539 (N_11539,N_11225,N_11354);
nor U11540 (N_11540,N_11309,N_11248);
and U11541 (N_11541,N_11232,N_11308);
or U11542 (N_11542,N_11265,N_11330);
nor U11543 (N_11543,N_11218,N_11397);
nor U11544 (N_11544,N_11390,N_11387);
or U11545 (N_11545,N_11370,N_11266);
nor U11546 (N_11546,N_11284,N_11316);
nor U11547 (N_11547,N_11327,N_11272);
nand U11548 (N_11548,N_11205,N_11364);
nor U11549 (N_11549,N_11253,N_11245);
or U11550 (N_11550,N_11318,N_11388);
xor U11551 (N_11551,N_11366,N_11228);
nor U11552 (N_11552,N_11293,N_11343);
and U11553 (N_11553,N_11203,N_11349);
and U11554 (N_11554,N_11369,N_11338);
nor U11555 (N_11555,N_11354,N_11333);
nand U11556 (N_11556,N_11374,N_11253);
or U11557 (N_11557,N_11387,N_11383);
nor U11558 (N_11558,N_11227,N_11201);
nand U11559 (N_11559,N_11253,N_11313);
nor U11560 (N_11560,N_11203,N_11301);
nor U11561 (N_11561,N_11358,N_11331);
and U11562 (N_11562,N_11313,N_11327);
or U11563 (N_11563,N_11325,N_11358);
nand U11564 (N_11564,N_11354,N_11373);
nor U11565 (N_11565,N_11220,N_11251);
and U11566 (N_11566,N_11319,N_11353);
nand U11567 (N_11567,N_11232,N_11399);
nor U11568 (N_11568,N_11322,N_11215);
and U11569 (N_11569,N_11327,N_11305);
nand U11570 (N_11570,N_11377,N_11320);
or U11571 (N_11571,N_11314,N_11322);
nor U11572 (N_11572,N_11398,N_11205);
and U11573 (N_11573,N_11351,N_11390);
or U11574 (N_11574,N_11267,N_11233);
nor U11575 (N_11575,N_11321,N_11304);
nand U11576 (N_11576,N_11286,N_11356);
or U11577 (N_11577,N_11326,N_11276);
nor U11578 (N_11578,N_11353,N_11301);
or U11579 (N_11579,N_11219,N_11200);
and U11580 (N_11580,N_11317,N_11307);
nand U11581 (N_11581,N_11305,N_11372);
or U11582 (N_11582,N_11359,N_11311);
nand U11583 (N_11583,N_11291,N_11299);
or U11584 (N_11584,N_11372,N_11311);
and U11585 (N_11585,N_11236,N_11370);
or U11586 (N_11586,N_11210,N_11297);
or U11587 (N_11587,N_11223,N_11230);
nand U11588 (N_11588,N_11327,N_11268);
nor U11589 (N_11589,N_11356,N_11207);
or U11590 (N_11590,N_11202,N_11235);
and U11591 (N_11591,N_11289,N_11383);
nor U11592 (N_11592,N_11260,N_11211);
and U11593 (N_11593,N_11353,N_11211);
nand U11594 (N_11594,N_11248,N_11348);
nand U11595 (N_11595,N_11206,N_11276);
or U11596 (N_11596,N_11336,N_11271);
nand U11597 (N_11597,N_11388,N_11378);
and U11598 (N_11598,N_11359,N_11318);
or U11599 (N_11599,N_11215,N_11266);
or U11600 (N_11600,N_11448,N_11406);
or U11601 (N_11601,N_11419,N_11559);
and U11602 (N_11602,N_11460,N_11586);
nand U11603 (N_11603,N_11437,N_11402);
and U11604 (N_11604,N_11536,N_11463);
nor U11605 (N_11605,N_11428,N_11582);
or U11606 (N_11606,N_11583,N_11566);
and U11607 (N_11607,N_11504,N_11507);
or U11608 (N_11608,N_11535,N_11537);
or U11609 (N_11609,N_11530,N_11579);
and U11610 (N_11610,N_11515,N_11540);
nand U11611 (N_11611,N_11409,N_11490);
nor U11612 (N_11612,N_11570,N_11455);
and U11613 (N_11613,N_11441,N_11426);
and U11614 (N_11614,N_11444,N_11564);
and U11615 (N_11615,N_11429,N_11459);
nand U11616 (N_11616,N_11424,N_11517);
nand U11617 (N_11617,N_11481,N_11442);
or U11618 (N_11618,N_11587,N_11422);
xnor U11619 (N_11619,N_11546,N_11458);
and U11620 (N_11620,N_11520,N_11525);
or U11621 (N_11621,N_11457,N_11433);
nand U11622 (N_11622,N_11413,N_11543);
and U11623 (N_11623,N_11462,N_11407);
and U11624 (N_11624,N_11423,N_11521);
nand U11625 (N_11625,N_11511,N_11508);
or U11626 (N_11626,N_11445,N_11486);
or U11627 (N_11627,N_11403,N_11558);
or U11628 (N_11628,N_11522,N_11539);
or U11629 (N_11629,N_11526,N_11461);
and U11630 (N_11630,N_11519,N_11534);
and U11631 (N_11631,N_11420,N_11538);
nor U11632 (N_11632,N_11593,N_11531);
or U11633 (N_11633,N_11557,N_11494);
and U11634 (N_11634,N_11509,N_11497);
nand U11635 (N_11635,N_11421,N_11430);
or U11636 (N_11636,N_11451,N_11405);
and U11637 (N_11637,N_11528,N_11597);
and U11638 (N_11638,N_11561,N_11483);
nor U11639 (N_11639,N_11529,N_11470);
nand U11640 (N_11640,N_11577,N_11434);
or U11641 (N_11641,N_11498,N_11552);
or U11642 (N_11642,N_11581,N_11542);
xor U11643 (N_11643,N_11450,N_11510);
or U11644 (N_11644,N_11449,N_11545);
nor U11645 (N_11645,N_11568,N_11411);
or U11646 (N_11646,N_11400,N_11469);
nand U11647 (N_11647,N_11495,N_11425);
and U11648 (N_11648,N_11474,N_11404);
or U11649 (N_11649,N_11479,N_11548);
and U11650 (N_11650,N_11456,N_11518);
and U11651 (N_11651,N_11482,N_11588);
nor U11652 (N_11652,N_11514,N_11550);
nor U11653 (N_11653,N_11574,N_11506);
or U11654 (N_11654,N_11447,N_11488);
or U11655 (N_11655,N_11527,N_11596);
nor U11656 (N_11656,N_11541,N_11547);
or U11657 (N_11657,N_11562,N_11473);
nand U11658 (N_11658,N_11565,N_11453);
nor U11659 (N_11659,N_11569,N_11468);
or U11660 (N_11660,N_11489,N_11464);
and U11661 (N_11661,N_11471,N_11553);
or U11662 (N_11662,N_11523,N_11502);
nor U11663 (N_11663,N_11415,N_11467);
nand U11664 (N_11664,N_11573,N_11478);
nor U11665 (N_11665,N_11524,N_11595);
nand U11666 (N_11666,N_11554,N_11414);
or U11667 (N_11667,N_11446,N_11499);
and U11668 (N_11668,N_11465,N_11598);
nand U11669 (N_11669,N_11452,N_11590);
nor U11670 (N_11670,N_11544,N_11578);
nand U11671 (N_11671,N_11503,N_11485);
nor U11672 (N_11672,N_11487,N_11513);
nor U11673 (N_11673,N_11501,N_11436);
or U11674 (N_11674,N_11532,N_11567);
or U11675 (N_11675,N_11443,N_11408);
nor U11676 (N_11676,N_11432,N_11599);
or U11677 (N_11677,N_11571,N_11454);
nand U11678 (N_11678,N_11492,N_11551);
nand U11679 (N_11679,N_11496,N_11491);
nor U11680 (N_11680,N_11431,N_11438);
or U11681 (N_11681,N_11439,N_11435);
or U11682 (N_11682,N_11476,N_11475);
nor U11683 (N_11683,N_11580,N_11500);
and U11684 (N_11684,N_11401,N_11484);
nor U11685 (N_11685,N_11585,N_11440);
or U11686 (N_11686,N_11416,N_11575);
or U11687 (N_11687,N_11516,N_11556);
nand U11688 (N_11688,N_11563,N_11576);
nand U11689 (N_11689,N_11591,N_11572);
nand U11690 (N_11690,N_11477,N_11560);
and U11691 (N_11691,N_11533,N_11412);
nor U11692 (N_11692,N_11472,N_11584);
or U11693 (N_11693,N_11589,N_11505);
nand U11694 (N_11694,N_11493,N_11418);
or U11695 (N_11695,N_11410,N_11592);
nor U11696 (N_11696,N_11466,N_11427);
nor U11697 (N_11697,N_11480,N_11417);
nand U11698 (N_11698,N_11555,N_11594);
nor U11699 (N_11699,N_11512,N_11549);
nor U11700 (N_11700,N_11402,N_11425);
or U11701 (N_11701,N_11499,N_11544);
or U11702 (N_11702,N_11481,N_11572);
and U11703 (N_11703,N_11511,N_11478);
and U11704 (N_11704,N_11585,N_11528);
nand U11705 (N_11705,N_11585,N_11460);
nor U11706 (N_11706,N_11493,N_11485);
and U11707 (N_11707,N_11543,N_11539);
nand U11708 (N_11708,N_11495,N_11400);
or U11709 (N_11709,N_11460,N_11542);
nor U11710 (N_11710,N_11513,N_11450);
nand U11711 (N_11711,N_11599,N_11572);
nor U11712 (N_11712,N_11418,N_11560);
or U11713 (N_11713,N_11599,N_11452);
nor U11714 (N_11714,N_11465,N_11558);
nand U11715 (N_11715,N_11481,N_11468);
nand U11716 (N_11716,N_11441,N_11492);
nand U11717 (N_11717,N_11480,N_11476);
xor U11718 (N_11718,N_11591,N_11448);
and U11719 (N_11719,N_11520,N_11589);
and U11720 (N_11720,N_11402,N_11576);
nor U11721 (N_11721,N_11505,N_11416);
and U11722 (N_11722,N_11409,N_11596);
nand U11723 (N_11723,N_11557,N_11424);
nand U11724 (N_11724,N_11544,N_11408);
and U11725 (N_11725,N_11412,N_11578);
and U11726 (N_11726,N_11498,N_11511);
and U11727 (N_11727,N_11561,N_11545);
or U11728 (N_11728,N_11524,N_11589);
nor U11729 (N_11729,N_11540,N_11524);
and U11730 (N_11730,N_11475,N_11421);
nor U11731 (N_11731,N_11463,N_11586);
and U11732 (N_11732,N_11540,N_11435);
or U11733 (N_11733,N_11495,N_11453);
and U11734 (N_11734,N_11473,N_11451);
nor U11735 (N_11735,N_11516,N_11542);
and U11736 (N_11736,N_11532,N_11541);
nor U11737 (N_11737,N_11598,N_11454);
nor U11738 (N_11738,N_11481,N_11576);
and U11739 (N_11739,N_11560,N_11444);
or U11740 (N_11740,N_11560,N_11534);
nand U11741 (N_11741,N_11571,N_11567);
or U11742 (N_11742,N_11588,N_11508);
nor U11743 (N_11743,N_11544,N_11472);
nand U11744 (N_11744,N_11564,N_11478);
nor U11745 (N_11745,N_11522,N_11531);
and U11746 (N_11746,N_11469,N_11552);
and U11747 (N_11747,N_11526,N_11566);
nand U11748 (N_11748,N_11599,N_11459);
or U11749 (N_11749,N_11526,N_11599);
nor U11750 (N_11750,N_11417,N_11597);
and U11751 (N_11751,N_11555,N_11403);
nand U11752 (N_11752,N_11529,N_11485);
and U11753 (N_11753,N_11480,N_11511);
or U11754 (N_11754,N_11414,N_11465);
and U11755 (N_11755,N_11562,N_11422);
or U11756 (N_11756,N_11576,N_11400);
nand U11757 (N_11757,N_11428,N_11430);
and U11758 (N_11758,N_11508,N_11514);
and U11759 (N_11759,N_11475,N_11405);
and U11760 (N_11760,N_11439,N_11453);
and U11761 (N_11761,N_11574,N_11534);
and U11762 (N_11762,N_11432,N_11577);
nand U11763 (N_11763,N_11561,N_11592);
nor U11764 (N_11764,N_11535,N_11444);
nor U11765 (N_11765,N_11597,N_11513);
and U11766 (N_11766,N_11400,N_11420);
or U11767 (N_11767,N_11541,N_11467);
nor U11768 (N_11768,N_11594,N_11499);
or U11769 (N_11769,N_11537,N_11424);
and U11770 (N_11770,N_11487,N_11427);
and U11771 (N_11771,N_11568,N_11420);
nor U11772 (N_11772,N_11429,N_11553);
nor U11773 (N_11773,N_11562,N_11409);
nand U11774 (N_11774,N_11571,N_11469);
or U11775 (N_11775,N_11426,N_11514);
xnor U11776 (N_11776,N_11517,N_11498);
nand U11777 (N_11777,N_11511,N_11400);
and U11778 (N_11778,N_11478,N_11438);
or U11779 (N_11779,N_11497,N_11538);
nand U11780 (N_11780,N_11429,N_11400);
or U11781 (N_11781,N_11404,N_11557);
nand U11782 (N_11782,N_11543,N_11457);
and U11783 (N_11783,N_11574,N_11561);
nand U11784 (N_11784,N_11443,N_11404);
or U11785 (N_11785,N_11508,N_11572);
and U11786 (N_11786,N_11543,N_11504);
nand U11787 (N_11787,N_11412,N_11409);
and U11788 (N_11788,N_11554,N_11461);
or U11789 (N_11789,N_11403,N_11511);
nor U11790 (N_11790,N_11535,N_11567);
or U11791 (N_11791,N_11414,N_11583);
or U11792 (N_11792,N_11583,N_11447);
or U11793 (N_11793,N_11455,N_11499);
and U11794 (N_11794,N_11467,N_11436);
and U11795 (N_11795,N_11559,N_11507);
or U11796 (N_11796,N_11539,N_11401);
nand U11797 (N_11797,N_11518,N_11460);
nor U11798 (N_11798,N_11581,N_11579);
nand U11799 (N_11799,N_11418,N_11523);
or U11800 (N_11800,N_11615,N_11673);
or U11801 (N_11801,N_11776,N_11654);
or U11802 (N_11802,N_11703,N_11702);
nor U11803 (N_11803,N_11726,N_11766);
nand U11804 (N_11804,N_11651,N_11609);
nor U11805 (N_11805,N_11704,N_11665);
nand U11806 (N_11806,N_11787,N_11670);
and U11807 (N_11807,N_11696,N_11718);
or U11808 (N_11808,N_11697,N_11752);
and U11809 (N_11809,N_11633,N_11616);
or U11810 (N_11810,N_11602,N_11764);
and U11811 (N_11811,N_11669,N_11680);
nand U11812 (N_11812,N_11793,N_11784);
or U11813 (N_11813,N_11610,N_11688);
or U11814 (N_11814,N_11652,N_11632);
or U11815 (N_11815,N_11711,N_11664);
and U11816 (N_11816,N_11644,N_11760);
and U11817 (N_11817,N_11732,N_11724);
and U11818 (N_11818,N_11601,N_11716);
and U11819 (N_11819,N_11740,N_11646);
nand U11820 (N_11820,N_11618,N_11627);
or U11821 (N_11821,N_11657,N_11775);
nor U11822 (N_11822,N_11628,N_11617);
or U11823 (N_11823,N_11743,N_11681);
or U11824 (N_11824,N_11727,N_11759);
or U11825 (N_11825,N_11631,N_11768);
xnor U11826 (N_11826,N_11663,N_11756);
or U11827 (N_11827,N_11771,N_11672);
or U11828 (N_11828,N_11734,N_11790);
nand U11829 (N_11829,N_11687,N_11643);
and U11830 (N_11830,N_11648,N_11721);
nor U11831 (N_11831,N_11736,N_11783);
or U11832 (N_11832,N_11640,N_11674);
nand U11833 (N_11833,N_11778,N_11638);
nor U11834 (N_11834,N_11773,N_11634);
nand U11835 (N_11835,N_11611,N_11765);
or U11836 (N_11836,N_11753,N_11695);
or U11837 (N_11837,N_11772,N_11662);
or U11838 (N_11838,N_11693,N_11751);
or U11839 (N_11839,N_11608,N_11710);
xnor U11840 (N_11840,N_11745,N_11733);
nand U11841 (N_11841,N_11746,N_11769);
or U11842 (N_11842,N_11698,N_11686);
and U11843 (N_11843,N_11699,N_11789);
or U11844 (N_11844,N_11679,N_11763);
and U11845 (N_11845,N_11641,N_11739);
nor U11846 (N_11846,N_11794,N_11781);
nor U11847 (N_11847,N_11712,N_11625);
and U11848 (N_11848,N_11770,N_11635);
or U11849 (N_11849,N_11639,N_11708);
nand U11850 (N_11850,N_11722,N_11676);
nor U11851 (N_11851,N_11700,N_11719);
and U11852 (N_11852,N_11767,N_11629);
and U11853 (N_11853,N_11797,N_11689);
nor U11854 (N_11854,N_11757,N_11701);
nor U11855 (N_11855,N_11796,N_11613);
or U11856 (N_11856,N_11649,N_11791);
nand U11857 (N_11857,N_11645,N_11655);
nor U11858 (N_11858,N_11777,N_11795);
nand U11859 (N_11859,N_11754,N_11709);
nand U11860 (N_11860,N_11706,N_11782);
nand U11861 (N_11861,N_11656,N_11675);
or U11862 (N_11862,N_11630,N_11637);
nand U11863 (N_11863,N_11642,N_11623);
xnor U11864 (N_11864,N_11605,N_11748);
or U11865 (N_11865,N_11624,N_11626);
nand U11866 (N_11866,N_11729,N_11620);
nand U11867 (N_11867,N_11666,N_11690);
and U11868 (N_11868,N_11730,N_11659);
or U11869 (N_11869,N_11668,N_11774);
and U11870 (N_11870,N_11622,N_11600);
nand U11871 (N_11871,N_11744,N_11762);
and U11872 (N_11872,N_11660,N_11661);
or U11873 (N_11873,N_11780,N_11742);
nor U11874 (N_11874,N_11677,N_11694);
nor U11875 (N_11875,N_11682,N_11720);
nand U11876 (N_11876,N_11705,N_11658);
nor U11877 (N_11877,N_11671,N_11685);
nor U11878 (N_11878,N_11755,N_11717);
nor U11879 (N_11879,N_11683,N_11738);
nand U11880 (N_11880,N_11741,N_11604);
nor U11881 (N_11881,N_11758,N_11750);
nor U11882 (N_11882,N_11786,N_11692);
nor U11883 (N_11883,N_11678,N_11650);
nor U11884 (N_11884,N_11707,N_11619);
or U11885 (N_11885,N_11647,N_11691);
nor U11886 (N_11886,N_11684,N_11636);
or U11887 (N_11887,N_11785,N_11792);
and U11888 (N_11888,N_11737,N_11723);
or U11889 (N_11889,N_11653,N_11607);
or U11890 (N_11890,N_11779,N_11731);
and U11891 (N_11891,N_11621,N_11614);
nand U11892 (N_11892,N_11612,N_11725);
or U11893 (N_11893,N_11799,N_11761);
and U11894 (N_11894,N_11728,N_11606);
nor U11895 (N_11895,N_11714,N_11603);
nand U11896 (N_11896,N_11735,N_11749);
and U11897 (N_11897,N_11747,N_11788);
nand U11898 (N_11898,N_11713,N_11667);
or U11899 (N_11899,N_11715,N_11798);
nor U11900 (N_11900,N_11697,N_11701);
nor U11901 (N_11901,N_11724,N_11730);
xor U11902 (N_11902,N_11791,N_11792);
nor U11903 (N_11903,N_11709,N_11758);
or U11904 (N_11904,N_11744,N_11734);
xor U11905 (N_11905,N_11798,N_11672);
nand U11906 (N_11906,N_11648,N_11676);
and U11907 (N_11907,N_11693,N_11659);
nor U11908 (N_11908,N_11601,N_11743);
or U11909 (N_11909,N_11769,N_11622);
and U11910 (N_11910,N_11648,N_11662);
nand U11911 (N_11911,N_11794,N_11751);
and U11912 (N_11912,N_11779,N_11637);
nor U11913 (N_11913,N_11799,N_11793);
and U11914 (N_11914,N_11628,N_11611);
and U11915 (N_11915,N_11620,N_11678);
nand U11916 (N_11916,N_11770,N_11622);
nor U11917 (N_11917,N_11734,N_11794);
nand U11918 (N_11918,N_11768,N_11748);
nand U11919 (N_11919,N_11778,N_11631);
nor U11920 (N_11920,N_11692,N_11722);
nor U11921 (N_11921,N_11693,N_11623);
nor U11922 (N_11922,N_11712,N_11795);
nand U11923 (N_11923,N_11610,N_11798);
nor U11924 (N_11924,N_11760,N_11675);
nand U11925 (N_11925,N_11706,N_11755);
and U11926 (N_11926,N_11653,N_11711);
nand U11927 (N_11927,N_11789,N_11755);
nor U11928 (N_11928,N_11755,N_11628);
nor U11929 (N_11929,N_11691,N_11706);
or U11930 (N_11930,N_11612,N_11741);
nand U11931 (N_11931,N_11663,N_11667);
nand U11932 (N_11932,N_11669,N_11711);
and U11933 (N_11933,N_11700,N_11756);
or U11934 (N_11934,N_11793,N_11656);
xnor U11935 (N_11935,N_11782,N_11682);
nor U11936 (N_11936,N_11639,N_11652);
nor U11937 (N_11937,N_11695,N_11650);
or U11938 (N_11938,N_11773,N_11704);
and U11939 (N_11939,N_11661,N_11751);
nor U11940 (N_11940,N_11687,N_11669);
and U11941 (N_11941,N_11791,N_11645);
or U11942 (N_11942,N_11656,N_11622);
nand U11943 (N_11943,N_11612,N_11779);
and U11944 (N_11944,N_11769,N_11723);
nand U11945 (N_11945,N_11717,N_11751);
and U11946 (N_11946,N_11689,N_11662);
and U11947 (N_11947,N_11633,N_11651);
or U11948 (N_11948,N_11778,N_11784);
nor U11949 (N_11949,N_11714,N_11730);
nand U11950 (N_11950,N_11692,N_11758);
and U11951 (N_11951,N_11680,N_11678);
and U11952 (N_11952,N_11655,N_11677);
or U11953 (N_11953,N_11768,N_11739);
nor U11954 (N_11954,N_11602,N_11637);
xor U11955 (N_11955,N_11728,N_11712);
and U11956 (N_11956,N_11626,N_11665);
or U11957 (N_11957,N_11713,N_11739);
nor U11958 (N_11958,N_11649,N_11672);
nand U11959 (N_11959,N_11755,N_11791);
or U11960 (N_11960,N_11684,N_11699);
and U11961 (N_11961,N_11678,N_11675);
and U11962 (N_11962,N_11605,N_11610);
or U11963 (N_11963,N_11779,N_11714);
or U11964 (N_11964,N_11633,N_11670);
nand U11965 (N_11965,N_11778,N_11642);
nor U11966 (N_11966,N_11666,N_11609);
or U11967 (N_11967,N_11757,N_11779);
and U11968 (N_11968,N_11652,N_11755);
nor U11969 (N_11969,N_11717,N_11725);
and U11970 (N_11970,N_11749,N_11696);
nor U11971 (N_11971,N_11654,N_11713);
or U11972 (N_11972,N_11767,N_11746);
or U11973 (N_11973,N_11621,N_11683);
or U11974 (N_11974,N_11738,N_11630);
xnor U11975 (N_11975,N_11712,N_11603);
nor U11976 (N_11976,N_11730,N_11765);
and U11977 (N_11977,N_11768,N_11673);
nor U11978 (N_11978,N_11767,N_11626);
nand U11979 (N_11979,N_11672,N_11739);
nand U11980 (N_11980,N_11665,N_11722);
or U11981 (N_11981,N_11616,N_11641);
nor U11982 (N_11982,N_11701,N_11656);
nand U11983 (N_11983,N_11733,N_11639);
nand U11984 (N_11984,N_11769,N_11664);
or U11985 (N_11985,N_11726,N_11774);
nor U11986 (N_11986,N_11768,N_11742);
and U11987 (N_11987,N_11722,N_11632);
xor U11988 (N_11988,N_11697,N_11729);
and U11989 (N_11989,N_11751,N_11799);
nor U11990 (N_11990,N_11686,N_11619);
nand U11991 (N_11991,N_11622,N_11695);
nand U11992 (N_11992,N_11755,N_11740);
xnor U11993 (N_11993,N_11613,N_11710);
nor U11994 (N_11994,N_11667,N_11736);
and U11995 (N_11995,N_11694,N_11758);
nand U11996 (N_11996,N_11729,N_11761);
or U11997 (N_11997,N_11666,N_11613);
nor U11998 (N_11998,N_11725,N_11705);
and U11999 (N_11999,N_11607,N_11675);
or U12000 (N_12000,N_11926,N_11875);
nor U12001 (N_12001,N_11826,N_11862);
nor U12002 (N_12002,N_11812,N_11852);
and U12003 (N_12003,N_11847,N_11915);
nand U12004 (N_12004,N_11971,N_11853);
or U12005 (N_12005,N_11833,N_11913);
nor U12006 (N_12006,N_11856,N_11949);
and U12007 (N_12007,N_11980,N_11948);
nor U12008 (N_12008,N_11902,N_11963);
nand U12009 (N_12009,N_11882,N_11842);
or U12010 (N_12010,N_11845,N_11953);
xnor U12011 (N_12011,N_11837,N_11828);
nor U12012 (N_12012,N_11806,N_11844);
nand U12013 (N_12013,N_11807,N_11923);
or U12014 (N_12014,N_11835,N_11878);
and U12015 (N_12015,N_11801,N_11995);
and U12016 (N_12016,N_11821,N_11904);
nand U12017 (N_12017,N_11909,N_11979);
or U12018 (N_12018,N_11900,N_11846);
nor U12019 (N_12019,N_11834,N_11892);
or U12020 (N_12020,N_11823,N_11973);
or U12021 (N_12021,N_11897,N_11962);
nor U12022 (N_12022,N_11860,N_11898);
or U12023 (N_12023,N_11800,N_11870);
and U12024 (N_12024,N_11903,N_11805);
or U12025 (N_12025,N_11886,N_11951);
nand U12026 (N_12026,N_11832,N_11854);
nand U12027 (N_12027,N_11955,N_11858);
nor U12028 (N_12028,N_11803,N_11864);
or U12029 (N_12029,N_11838,N_11901);
nand U12030 (N_12030,N_11929,N_11867);
and U12031 (N_12031,N_11932,N_11942);
nor U12032 (N_12032,N_11908,N_11937);
nand U12033 (N_12033,N_11907,N_11910);
nor U12034 (N_12034,N_11944,N_11936);
or U12035 (N_12035,N_11946,N_11820);
and U12036 (N_12036,N_11810,N_11885);
and U12037 (N_12037,N_11912,N_11859);
nor U12038 (N_12038,N_11802,N_11935);
nor U12039 (N_12039,N_11976,N_11814);
or U12040 (N_12040,N_11848,N_11871);
and U12041 (N_12041,N_11977,N_11829);
or U12042 (N_12042,N_11836,N_11952);
nand U12043 (N_12043,N_11968,N_11881);
and U12044 (N_12044,N_11997,N_11876);
nor U12045 (N_12045,N_11831,N_11991);
nand U12046 (N_12046,N_11855,N_11975);
nand U12047 (N_12047,N_11939,N_11960);
or U12048 (N_12048,N_11985,N_11933);
or U12049 (N_12049,N_11972,N_11906);
nand U12050 (N_12050,N_11865,N_11927);
and U12051 (N_12051,N_11917,N_11922);
or U12052 (N_12052,N_11815,N_11984);
or U12053 (N_12053,N_11850,N_11888);
or U12054 (N_12054,N_11887,N_11830);
and U12055 (N_12055,N_11827,N_11947);
nor U12056 (N_12056,N_11896,N_11839);
or U12057 (N_12057,N_11938,N_11964);
and U12058 (N_12058,N_11990,N_11811);
or U12059 (N_12059,N_11924,N_11925);
nor U12060 (N_12060,N_11994,N_11911);
or U12061 (N_12061,N_11861,N_11816);
nand U12062 (N_12062,N_11965,N_11956);
or U12063 (N_12063,N_11954,N_11974);
nor U12064 (N_12064,N_11824,N_11890);
nand U12065 (N_12065,N_11992,N_11804);
nor U12066 (N_12066,N_11921,N_11993);
nand U12067 (N_12067,N_11983,N_11808);
nor U12068 (N_12068,N_11872,N_11866);
nor U12069 (N_12069,N_11879,N_11884);
nor U12070 (N_12070,N_11899,N_11941);
nand U12071 (N_12071,N_11996,N_11840);
or U12072 (N_12072,N_11928,N_11957);
nor U12073 (N_12073,N_11843,N_11873);
nor U12074 (N_12074,N_11959,N_11869);
nand U12075 (N_12075,N_11874,N_11989);
and U12076 (N_12076,N_11982,N_11943);
nand U12077 (N_12077,N_11940,N_11905);
nand U12078 (N_12078,N_11891,N_11819);
or U12079 (N_12079,N_11851,N_11931);
or U12080 (N_12080,N_11916,N_11969);
and U12081 (N_12081,N_11822,N_11945);
and U12082 (N_12082,N_11841,N_11958);
or U12083 (N_12083,N_11895,N_11988);
nor U12084 (N_12084,N_11999,N_11809);
nor U12085 (N_12085,N_11857,N_11877);
and U12086 (N_12086,N_11868,N_11930);
and U12087 (N_12087,N_11998,N_11880);
and U12088 (N_12088,N_11919,N_11950);
nand U12089 (N_12089,N_11825,N_11920);
nor U12090 (N_12090,N_11970,N_11863);
or U12091 (N_12091,N_11889,N_11978);
nor U12092 (N_12092,N_11894,N_11961);
nor U12093 (N_12093,N_11818,N_11981);
nor U12094 (N_12094,N_11934,N_11918);
nand U12095 (N_12095,N_11893,N_11986);
nand U12096 (N_12096,N_11813,N_11914);
or U12097 (N_12097,N_11849,N_11966);
nand U12098 (N_12098,N_11883,N_11967);
and U12099 (N_12099,N_11987,N_11817);
nand U12100 (N_12100,N_11867,N_11817);
or U12101 (N_12101,N_11815,N_11949);
nor U12102 (N_12102,N_11805,N_11948);
nand U12103 (N_12103,N_11891,N_11809);
nand U12104 (N_12104,N_11915,N_11941);
nor U12105 (N_12105,N_11803,N_11907);
nor U12106 (N_12106,N_11924,N_11908);
and U12107 (N_12107,N_11930,N_11984);
or U12108 (N_12108,N_11903,N_11904);
and U12109 (N_12109,N_11948,N_11962);
and U12110 (N_12110,N_11940,N_11820);
or U12111 (N_12111,N_11813,N_11992);
or U12112 (N_12112,N_11820,N_11975);
or U12113 (N_12113,N_11959,N_11986);
and U12114 (N_12114,N_11998,N_11954);
nand U12115 (N_12115,N_11954,N_11914);
and U12116 (N_12116,N_11935,N_11962);
nor U12117 (N_12117,N_11921,N_11873);
nand U12118 (N_12118,N_11921,N_11802);
nand U12119 (N_12119,N_11936,N_11818);
or U12120 (N_12120,N_11967,N_11981);
nor U12121 (N_12121,N_11853,N_11897);
and U12122 (N_12122,N_11939,N_11934);
nor U12123 (N_12123,N_11853,N_11885);
nand U12124 (N_12124,N_11881,N_11814);
and U12125 (N_12125,N_11861,N_11932);
nor U12126 (N_12126,N_11967,N_11991);
and U12127 (N_12127,N_11816,N_11998);
nand U12128 (N_12128,N_11957,N_11946);
and U12129 (N_12129,N_11988,N_11949);
nand U12130 (N_12130,N_11801,N_11826);
nor U12131 (N_12131,N_11900,N_11802);
nor U12132 (N_12132,N_11941,N_11919);
nand U12133 (N_12133,N_11975,N_11949);
xnor U12134 (N_12134,N_11876,N_11843);
or U12135 (N_12135,N_11876,N_11980);
nor U12136 (N_12136,N_11841,N_11981);
and U12137 (N_12137,N_11866,N_11954);
nor U12138 (N_12138,N_11974,N_11890);
or U12139 (N_12139,N_11932,N_11926);
nand U12140 (N_12140,N_11872,N_11983);
nand U12141 (N_12141,N_11925,N_11821);
and U12142 (N_12142,N_11865,N_11916);
or U12143 (N_12143,N_11973,N_11856);
or U12144 (N_12144,N_11917,N_11900);
or U12145 (N_12145,N_11982,N_11826);
nor U12146 (N_12146,N_11925,N_11888);
nor U12147 (N_12147,N_11844,N_11855);
nand U12148 (N_12148,N_11855,N_11826);
and U12149 (N_12149,N_11814,N_11832);
nor U12150 (N_12150,N_11957,N_11948);
or U12151 (N_12151,N_11999,N_11831);
nand U12152 (N_12152,N_11968,N_11883);
nand U12153 (N_12153,N_11986,N_11883);
nand U12154 (N_12154,N_11981,N_11968);
or U12155 (N_12155,N_11863,N_11825);
or U12156 (N_12156,N_11941,N_11994);
nor U12157 (N_12157,N_11809,N_11863);
nand U12158 (N_12158,N_11800,N_11971);
nand U12159 (N_12159,N_11921,N_11813);
and U12160 (N_12160,N_11810,N_11888);
and U12161 (N_12161,N_11943,N_11860);
or U12162 (N_12162,N_11953,N_11803);
nor U12163 (N_12163,N_11879,N_11927);
nand U12164 (N_12164,N_11961,N_11901);
and U12165 (N_12165,N_11838,N_11892);
nor U12166 (N_12166,N_11911,N_11802);
or U12167 (N_12167,N_11952,N_11993);
nand U12168 (N_12168,N_11863,N_11940);
or U12169 (N_12169,N_11824,N_11928);
or U12170 (N_12170,N_11923,N_11990);
or U12171 (N_12171,N_11836,N_11828);
and U12172 (N_12172,N_11896,N_11854);
nand U12173 (N_12173,N_11828,N_11924);
nor U12174 (N_12174,N_11852,N_11959);
or U12175 (N_12175,N_11853,N_11964);
and U12176 (N_12176,N_11835,N_11919);
or U12177 (N_12177,N_11995,N_11880);
or U12178 (N_12178,N_11887,N_11869);
or U12179 (N_12179,N_11984,N_11884);
or U12180 (N_12180,N_11854,N_11987);
and U12181 (N_12181,N_11951,N_11852);
nor U12182 (N_12182,N_11849,N_11948);
nor U12183 (N_12183,N_11873,N_11922);
and U12184 (N_12184,N_11803,N_11875);
nor U12185 (N_12185,N_11814,N_11915);
nand U12186 (N_12186,N_11940,N_11960);
nand U12187 (N_12187,N_11895,N_11950);
or U12188 (N_12188,N_11905,N_11977);
xor U12189 (N_12189,N_11872,N_11925);
or U12190 (N_12190,N_11986,N_11877);
and U12191 (N_12191,N_11849,N_11840);
nand U12192 (N_12192,N_11856,N_11896);
and U12193 (N_12193,N_11881,N_11853);
nor U12194 (N_12194,N_11975,N_11967);
nand U12195 (N_12195,N_11836,N_11878);
or U12196 (N_12196,N_11908,N_11832);
or U12197 (N_12197,N_11937,N_11861);
nand U12198 (N_12198,N_11908,N_11985);
nor U12199 (N_12199,N_11935,N_11919);
and U12200 (N_12200,N_12058,N_12039);
nor U12201 (N_12201,N_12029,N_12157);
and U12202 (N_12202,N_12053,N_12104);
or U12203 (N_12203,N_12134,N_12151);
nand U12204 (N_12204,N_12191,N_12102);
or U12205 (N_12205,N_12019,N_12022);
and U12206 (N_12206,N_12085,N_12008);
nand U12207 (N_12207,N_12069,N_12090);
and U12208 (N_12208,N_12173,N_12142);
or U12209 (N_12209,N_12052,N_12178);
nor U12210 (N_12210,N_12198,N_12036);
and U12211 (N_12211,N_12097,N_12025);
or U12212 (N_12212,N_12035,N_12038);
and U12213 (N_12213,N_12083,N_12009);
nand U12214 (N_12214,N_12032,N_12141);
and U12215 (N_12215,N_12153,N_12093);
and U12216 (N_12216,N_12072,N_12079);
or U12217 (N_12217,N_12131,N_12189);
nor U12218 (N_12218,N_12040,N_12171);
nand U12219 (N_12219,N_12165,N_12100);
and U12220 (N_12220,N_12065,N_12066);
or U12221 (N_12221,N_12042,N_12106);
or U12222 (N_12222,N_12007,N_12091);
nand U12223 (N_12223,N_12051,N_12027);
or U12224 (N_12224,N_12168,N_12143);
and U12225 (N_12225,N_12084,N_12109);
nor U12226 (N_12226,N_12136,N_12192);
nand U12227 (N_12227,N_12043,N_12081);
nor U12228 (N_12228,N_12161,N_12125);
nand U12229 (N_12229,N_12119,N_12129);
nand U12230 (N_12230,N_12166,N_12121);
nor U12231 (N_12231,N_12179,N_12152);
nor U12232 (N_12232,N_12057,N_12064);
nand U12233 (N_12233,N_12094,N_12098);
and U12234 (N_12234,N_12010,N_12089);
and U12235 (N_12235,N_12174,N_12110);
nor U12236 (N_12236,N_12195,N_12167);
nor U12237 (N_12237,N_12183,N_12190);
nor U12238 (N_12238,N_12150,N_12082);
nand U12239 (N_12239,N_12138,N_12075);
nand U12240 (N_12240,N_12108,N_12193);
nand U12241 (N_12241,N_12194,N_12088);
nand U12242 (N_12242,N_12095,N_12067);
nand U12243 (N_12243,N_12068,N_12148);
nand U12244 (N_12244,N_12123,N_12062);
nand U12245 (N_12245,N_12101,N_12133);
nor U12246 (N_12246,N_12113,N_12001);
nand U12247 (N_12247,N_12112,N_12144);
nor U12248 (N_12248,N_12156,N_12199);
nor U12249 (N_12249,N_12004,N_12162);
and U12250 (N_12250,N_12078,N_12074);
and U12251 (N_12251,N_12023,N_12086);
or U12252 (N_12252,N_12158,N_12103);
and U12253 (N_12253,N_12177,N_12126);
and U12254 (N_12254,N_12117,N_12130);
and U12255 (N_12255,N_12163,N_12107);
nand U12256 (N_12256,N_12160,N_12122);
nand U12257 (N_12257,N_12147,N_12146);
or U12258 (N_12258,N_12030,N_12056);
nand U12259 (N_12259,N_12105,N_12132);
nand U12260 (N_12260,N_12018,N_12135);
and U12261 (N_12261,N_12092,N_12155);
and U12262 (N_12262,N_12055,N_12099);
nand U12263 (N_12263,N_12076,N_12197);
and U12264 (N_12264,N_12015,N_12028);
nor U12265 (N_12265,N_12061,N_12002);
nand U12266 (N_12266,N_12060,N_12041);
nand U12267 (N_12267,N_12059,N_12127);
or U12268 (N_12268,N_12115,N_12026);
nand U12269 (N_12269,N_12017,N_12031);
nor U12270 (N_12270,N_12050,N_12176);
or U12271 (N_12271,N_12188,N_12111);
nand U12272 (N_12272,N_12024,N_12003);
nand U12273 (N_12273,N_12021,N_12020);
nand U12274 (N_12274,N_12080,N_12005);
and U12275 (N_12275,N_12047,N_12114);
and U12276 (N_12276,N_12063,N_12012);
nor U12277 (N_12277,N_12187,N_12037);
nor U12278 (N_12278,N_12175,N_12054);
nand U12279 (N_12279,N_12045,N_12044);
and U12280 (N_12280,N_12124,N_12034);
and U12281 (N_12281,N_12186,N_12087);
nor U12282 (N_12282,N_12140,N_12006);
or U12283 (N_12283,N_12145,N_12184);
nand U12284 (N_12284,N_12011,N_12073);
or U12285 (N_12285,N_12164,N_12182);
or U12286 (N_12286,N_12154,N_12181);
nand U12287 (N_12287,N_12128,N_12077);
xnor U12288 (N_12288,N_12149,N_12196);
nor U12289 (N_12289,N_12116,N_12014);
and U12290 (N_12290,N_12120,N_12049);
or U12291 (N_12291,N_12070,N_12048);
nand U12292 (N_12292,N_12137,N_12118);
nand U12293 (N_12293,N_12013,N_12033);
nor U12294 (N_12294,N_12071,N_12159);
and U12295 (N_12295,N_12000,N_12096);
and U12296 (N_12296,N_12139,N_12046);
xor U12297 (N_12297,N_12172,N_12169);
and U12298 (N_12298,N_12185,N_12016);
and U12299 (N_12299,N_12180,N_12170);
nor U12300 (N_12300,N_12144,N_12089);
and U12301 (N_12301,N_12064,N_12167);
nand U12302 (N_12302,N_12129,N_12078);
or U12303 (N_12303,N_12137,N_12075);
nor U12304 (N_12304,N_12184,N_12063);
or U12305 (N_12305,N_12092,N_12037);
or U12306 (N_12306,N_12031,N_12148);
or U12307 (N_12307,N_12167,N_12041);
nor U12308 (N_12308,N_12181,N_12006);
and U12309 (N_12309,N_12158,N_12015);
and U12310 (N_12310,N_12119,N_12146);
xnor U12311 (N_12311,N_12052,N_12101);
and U12312 (N_12312,N_12099,N_12116);
nand U12313 (N_12313,N_12102,N_12182);
or U12314 (N_12314,N_12102,N_12170);
or U12315 (N_12315,N_12090,N_12073);
or U12316 (N_12316,N_12057,N_12029);
nor U12317 (N_12317,N_12065,N_12197);
nand U12318 (N_12318,N_12168,N_12192);
or U12319 (N_12319,N_12118,N_12129);
and U12320 (N_12320,N_12120,N_12117);
or U12321 (N_12321,N_12072,N_12057);
nor U12322 (N_12322,N_12188,N_12134);
or U12323 (N_12323,N_12093,N_12059);
and U12324 (N_12324,N_12102,N_12115);
nand U12325 (N_12325,N_12192,N_12019);
or U12326 (N_12326,N_12168,N_12001);
and U12327 (N_12327,N_12138,N_12100);
and U12328 (N_12328,N_12166,N_12164);
nor U12329 (N_12329,N_12078,N_12059);
or U12330 (N_12330,N_12188,N_12107);
nand U12331 (N_12331,N_12190,N_12011);
or U12332 (N_12332,N_12037,N_12184);
and U12333 (N_12333,N_12036,N_12014);
nor U12334 (N_12334,N_12062,N_12060);
nand U12335 (N_12335,N_12139,N_12176);
nor U12336 (N_12336,N_12100,N_12107);
nor U12337 (N_12337,N_12095,N_12001);
or U12338 (N_12338,N_12183,N_12119);
nand U12339 (N_12339,N_12109,N_12118);
or U12340 (N_12340,N_12094,N_12179);
nand U12341 (N_12341,N_12002,N_12130);
nor U12342 (N_12342,N_12095,N_12164);
and U12343 (N_12343,N_12085,N_12043);
or U12344 (N_12344,N_12173,N_12102);
nand U12345 (N_12345,N_12077,N_12098);
or U12346 (N_12346,N_12181,N_12090);
nor U12347 (N_12347,N_12050,N_12038);
nand U12348 (N_12348,N_12054,N_12141);
nor U12349 (N_12349,N_12033,N_12003);
nor U12350 (N_12350,N_12020,N_12170);
nor U12351 (N_12351,N_12011,N_12057);
nand U12352 (N_12352,N_12107,N_12005);
nor U12353 (N_12353,N_12000,N_12014);
or U12354 (N_12354,N_12169,N_12121);
nand U12355 (N_12355,N_12010,N_12126);
or U12356 (N_12356,N_12029,N_12017);
nor U12357 (N_12357,N_12019,N_12076);
and U12358 (N_12358,N_12061,N_12099);
or U12359 (N_12359,N_12103,N_12055);
or U12360 (N_12360,N_12125,N_12158);
and U12361 (N_12361,N_12163,N_12121);
nor U12362 (N_12362,N_12181,N_12118);
and U12363 (N_12363,N_12158,N_12129);
or U12364 (N_12364,N_12116,N_12142);
or U12365 (N_12365,N_12004,N_12005);
nor U12366 (N_12366,N_12175,N_12057);
or U12367 (N_12367,N_12125,N_12055);
nor U12368 (N_12368,N_12023,N_12036);
nand U12369 (N_12369,N_12049,N_12037);
and U12370 (N_12370,N_12171,N_12012);
nor U12371 (N_12371,N_12107,N_12047);
or U12372 (N_12372,N_12092,N_12081);
nor U12373 (N_12373,N_12116,N_12192);
and U12374 (N_12374,N_12121,N_12181);
nor U12375 (N_12375,N_12169,N_12043);
and U12376 (N_12376,N_12196,N_12190);
nor U12377 (N_12377,N_12071,N_12140);
nor U12378 (N_12378,N_12124,N_12164);
nor U12379 (N_12379,N_12083,N_12084);
or U12380 (N_12380,N_12079,N_12126);
nor U12381 (N_12381,N_12031,N_12047);
nor U12382 (N_12382,N_12095,N_12173);
or U12383 (N_12383,N_12122,N_12137);
and U12384 (N_12384,N_12168,N_12170);
or U12385 (N_12385,N_12107,N_12105);
nand U12386 (N_12386,N_12057,N_12147);
nor U12387 (N_12387,N_12048,N_12093);
nand U12388 (N_12388,N_12112,N_12109);
and U12389 (N_12389,N_12019,N_12077);
nand U12390 (N_12390,N_12152,N_12030);
nor U12391 (N_12391,N_12171,N_12198);
or U12392 (N_12392,N_12097,N_12005);
and U12393 (N_12393,N_12040,N_12162);
or U12394 (N_12394,N_12102,N_12198);
and U12395 (N_12395,N_12109,N_12081);
or U12396 (N_12396,N_12019,N_12146);
nand U12397 (N_12397,N_12178,N_12115);
and U12398 (N_12398,N_12033,N_12018);
nand U12399 (N_12399,N_12063,N_12005);
or U12400 (N_12400,N_12283,N_12305);
and U12401 (N_12401,N_12244,N_12300);
nor U12402 (N_12402,N_12375,N_12349);
nor U12403 (N_12403,N_12311,N_12367);
or U12404 (N_12404,N_12332,N_12277);
nand U12405 (N_12405,N_12260,N_12392);
or U12406 (N_12406,N_12322,N_12363);
and U12407 (N_12407,N_12396,N_12222);
nor U12408 (N_12408,N_12383,N_12347);
or U12409 (N_12409,N_12270,N_12236);
nor U12410 (N_12410,N_12211,N_12266);
and U12411 (N_12411,N_12296,N_12204);
or U12412 (N_12412,N_12224,N_12246);
nor U12413 (N_12413,N_12262,N_12342);
nand U12414 (N_12414,N_12388,N_12362);
and U12415 (N_12415,N_12216,N_12251);
nor U12416 (N_12416,N_12214,N_12237);
or U12417 (N_12417,N_12213,N_12239);
nor U12418 (N_12418,N_12365,N_12309);
or U12419 (N_12419,N_12379,N_12361);
or U12420 (N_12420,N_12380,N_12329);
nor U12421 (N_12421,N_12376,N_12324);
or U12422 (N_12422,N_12235,N_12327);
or U12423 (N_12423,N_12233,N_12387);
and U12424 (N_12424,N_12294,N_12368);
and U12425 (N_12425,N_12360,N_12301);
nand U12426 (N_12426,N_12346,N_12314);
nand U12427 (N_12427,N_12255,N_12345);
nor U12428 (N_12428,N_12374,N_12292);
and U12429 (N_12429,N_12297,N_12350);
nor U12430 (N_12430,N_12372,N_12293);
or U12431 (N_12431,N_12307,N_12355);
nor U12432 (N_12432,N_12354,N_12335);
and U12433 (N_12433,N_12366,N_12282);
or U12434 (N_12434,N_12364,N_12319);
nand U12435 (N_12435,N_12227,N_12303);
and U12436 (N_12436,N_12264,N_12280);
nor U12437 (N_12437,N_12261,N_12247);
or U12438 (N_12438,N_12358,N_12348);
and U12439 (N_12439,N_12208,N_12217);
or U12440 (N_12440,N_12397,N_12268);
nand U12441 (N_12441,N_12340,N_12321);
and U12442 (N_12442,N_12212,N_12339);
xor U12443 (N_12443,N_12353,N_12338);
nor U12444 (N_12444,N_12328,N_12206);
nand U12445 (N_12445,N_12291,N_12394);
and U12446 (N_12446,N_12250,N_12234);
nand U12447 (N_12447,N_12285,N_12267);
nor U12448 (N_12448,N_12389,N_12308);
and U12449 (N_12449,N_12325,N_12359);
nor U12450 (N_12450,N_12232,N_12316);
or U12451 (N_12451,N_12278,N_12238);
and U12452 (N_12452,N_12299,N_12371);
or U12453 (N_12453,N_12265,N_12295);
nor U12454 (N_12454,N_12352,N_12326);
nor U12455 (N_12455,N_12333,N_12302);
nor U12456 (N_12456,N_12310,N_12386);
nor U12457 (N_12457,N_12241,N_12223);
nand U12458 (N_12458,N_12248,N_12229);
and U12459 (N_12459,N_12289,N_12351);
and U12460 (N_12460,N_12207,N_12334);
and U12461 (N_12461,N_12385,N_12210);
nor U12462 (N_12462,N_12259,N_12344);
nor U12463 (N_12463,N_12317,N_12271);
and U12464 (N_12464,N_12377,N_12343);
nand U12465 (N_12465,N_12382,N_12218);
nand U12466 (N_12466,N_12315,N_12275);
or U12467 (N_12467,N_12231,N_12220);
and U12468 (N_12468,N_12395,N_12272);
nand U12469 (N_12469,N_12398,N_12378);
and U12470 (N_12470,N_12202,N_12356);
nor U12471 (N_12471,N_12240,N_12269);
or U12472 (N_12472,N_12252,N_12290);
nand U12473 (N_12473,N_12298,N_12287);
or U12474 (N_12474,N_12256,N_12253);
nand U12475 (N_12475,N_12323,N_12225);
and U12476 (N_12476,N_12219,N_12228);
nor U12477 (N_12477,N_12381,N_12370);
nor U12478 (N_12478,N_12391,N_12330);
nor U12479 (N_12479,N_12226,N_12304);
nand U12480 (N_12480,N_12254,N_12205);
and U12481 (N_12481,N_12320,N_12399);
nand U12482 (N_12482,N_12373,N_12393);
or U12483 (N_12483,N_12288,N_12337);
nand U12484 (N_12484,N_12341,N_12221);
and U12485 (N_12485,N_12331,N_12284);
or U12486 (N_12486,N_12313,N_12273);
nand U12487 (N_12487,N_12384,N_12201);
and U12488 (N_12488,N_12390,N_12369);
nand U12489 (N_12489,N_12230,N_12312);
or U12490 (N_12490,N_12276,N_12215);
or U12491 (N_12491,N_12243,N_12274);
nand U12492 (N_12492,N_12242,N_12286);
nand U12493 (N_12493,N_12279,N_12336);
or U12494 (N_12494,N_12200,N_12263);
nor U12495 (N_12495,N_12258,N_12318);
and U12496 (N_12496,N_12281,N_12209);
and U12497 (N_12497,N_12245,N_12203);
nand U12498 (N_12498,N_12249,N_12257);
or U12499 (N_12499,N_12357,N_12306);
nor U12500 (N_12500,N_12378,N_12225);
nor U12501 (N_12501,N_12354,N_12386);
nand U12502 (N_12502,N_12399,N_12375);
nand U12503 (N_12503,N_12288,N_12271);
nand U12504 (N_12504,N_12381,N_12397);
nand U12505 (N_12505,N_12308,N_12339);
nor U12506 (N_12506,N_12306,N_12261);
and U12507 (N_12507,N_12342,N_12224);
nor U12508 (N_12508,N_12268,N_12334);
or U12509 (N_12509,N_12331,N_12207);
and U12510 (N_12510,N_12264,N_12364);
nor U12511 (N_12511,N_12330,N_12293);
and U12512 (N_12512,N_12271,N_12346);
nand U12513 (N_12513,N_12318,N_12362);
or U12514 (N_12514,N_12238,N_12296);
nand U12515 (N_12515,N_12312,N_12297);
nor U12516 (N_12516,N_12270,N_12283);
nor U12517 (N_12517,N_12270,N_12305);
and U12518 (N_12518,N_12253,N_12226);
or U12519 (N_12519,N_12282,N_12287);
nand U12520 (N_12520,N_12310,N_12384);
and U12521 (N_12521,N_12372,N_12393);
and U12522 (N_12522,N_12374,N_12318);
nor U12523 (N_12523,N_12384,N_12287);
nand U12524 (N_12524,N_12241,N_12262);
nand U12525 (N_12525,N_12375,N_12200);
or U12526 (N_12526,N_12284,N_12260);
and U12527 (N_12527,N_12387,N_12248);
or U12528 (N_12528,N_12214,N_12372);
nor U12529 (N_12529,N_12326,N_12334);
xor U12530 (N_12530,N_12321,N_12210);
nor U12531 (N_12531,N_12250,N_12219);
nor U12532 (N_12532,N_12374,N_12329);
nor U12533 (N_12533,N_12297,N_12269);
and U12534 (N_12534,N_12252,N_12255);
nand U12535 (N_12535,N_12345,N_12393);
nor U12536 (N_12536,N_12241,N_12338);
and U12537 (N_12537,N_12351,N_12291);
or U12538 (N_12538,N_12330,N_12384);
nand U12539 (N_12539,N_12271,N_12331);
nor U12540 (N_12540,N_12340,N_12358);
nor U12541 (N_12541,N_12354,N_12356);
and U12542 (N_12542,N_12370,N_12326);
xnor U12543 (N_12543,N_12331,N_12385);
and U12544 (N_12544,N_12350,N_12341);
and U12545 (N_12545,N_12226,N_12354);
xnor U12546 (N_12546,N_12212,N_12232);
nor U12547 (N_12547,N_12348,N_12367);
nand U12548 (N_12548,N_12393,N_12292);
nand U12549 (N_12549,N_12216,N_12395);
and U12550 (N_12550,N_12338,N_12335);
or U12551 (N_12551,N_12228,N_12317);
or U12552 (N_12552,N_12371,N_12290);
nand U12553 (N_12553,N_12259,N_12382);
nor U12554 (N_12554,N_12259,N_12363);
nor U12555 (N_12555,N_12305,N_12375);
nand U12556 (N_12556,N_12260,N_12356);
nand U12557 (N_12557,N_12361,N_12213);
nand U12558 (N_12558,N_12238,N_12385);
nor U12559 (N_12559,N_12238,N_12288);
nand U12560 (N_12560,N_12251,N_12351);
and U12561 (N_12561,N_12201,N_12307);
and U12562 (N_12562,N_12308,N_12248);
or U12563 (N_12563,N_12223,N_12323);
or U12564 (N_12564,N_12300,N_12285);
or U12565 (N_12565,N_12381,N_12301);
nor U12566 (N_12566,N_12270,N_12391);
and U12567 (N_12567,N_12223,N_12296);
or U12568 (N_12568,N_12383,N_12362);
or U12569 (N_12569,N_12353,N_12347);
and U12570 (N_12570,N_12379,N_12333);
and U12571 (N_12571,N_12264,N_12209);
and U12572 (N_12572,N_12325,N_12367);
or U12573 (N_12573,N_12383,N_12371);
nand U12574 (N_12574,N_12308,N_12241);
and U12575 (N_12575,N_12311,N_12378);
or U12576 (N_12576,N_12392,N_12313);
nor U12577 (N_12577,N_12357,N_12286);
and U12578 (N_12578,N_12203,N_12335);
nor U12579 (N_12579,N_12296,N_12373);
or U12580 (N_12580,N_12358,N_12209);
and U12581 (N_12581,N_12239,N_12253);
and U12582 (N_12582,N_12313,N_12353);
nand U12583 (N_12583,N_12276,N_12380);
nand U12584 (N_12584,N_12374,N_12358);
and U12585 (N_12585,N_12321,N_12258);
nor U12586 (N_12586,N_12275,N_12396);
or U12587 (N_12587,N_12221,N_12294);
or U12588 (N_12588,N_12372,N_12263);
nor U12589 (N_12589,N_12334,N_12361);
and U12590 (N_12590,N_12332,N_12231);
nand U12591 (N_12591,N_12379,N_12364);
and U12592 (N_12592,N_12281,N_12299);
nor U12593 (N_12593,N_12235,N_12309);
nor U12594 (N_12594,N_12316,N_12238);
and U12595 (N_12595,N_12306,N_12374);
nand U12596 (N_12596,N_12328,N_12393);
or U12597 (N_12597,N_12341,N_12366);
nor U12598 (N_12598,N_12239,N_12250);
or U12599 (N_12599,N_12328,N_12285);
nand U12600 (N_12600,N_12460,N_12429);
nor U12601 (N_12601,N_12418,N_12453);
and U12602 (N_12602,N_12438,N_12446);
or U12603 (N_12603,N_12514,N_12535);
and U12604 (N_12604,N_12409,N_12492);
nor U12605 (N_12605,N_12543,N_12553);
or U12606 (N_12606,N_12545,N_12528);
or U12607 (N_12607,N_12539,N_12560);
nor U12608 (N_12608,N_12458,N_12402);
or U12609 (N_12609,N_12502,N_12530);
or U12610 (N_12610,N_12421,N_12470);
nor U12611 (N_12611,N_12435,N_12534);
or U12612 (N_12612,N_12574,N_12546);
and U12613 (N_12613,N_12519,N_12437);
nor U12614 (N_12614,N_12516,N_12433);
or U12615 (N_12615,N_12489,N_12548);
and U12616 (N_12616,N_12414,N_12477);
nand U12617 (N_12617,N_12593,N_12562);
and U12618 (N_12618,N_12499,N_12478);
and U12619 (N_12619,N_12581,N_12420);
and U12620 (N_12620,N_12599,N_12517);
nand U12621 (N_12621,N_12518,N_12454);
nand U12622 (N_12622,N_12552,N_12428);
or U12623 (N_12623,N_12413,N_12587);
nor U12624 (N_12624,N_12510,N_12467);
xor U12625 (N_12625,N_12583,N_12590);
and U12626 (N_12626,N_12584,N_12491);
nor U12627 (N_12627,N_12401,N_12423);
nor U12628 (N_12628,N_12588,N_12496);
and U12629 (N_12629,N_12494,N_12577);
or U12630 (N_12630,N_12415,N_12404);
nand U12631 (N_12631,N_12500,N_12472);
nor U12632 (N_12632,N_12531,N_12424);
or U12633 (N_12633,N_12445,N_12511);
or U12634 (N_12634,N_12484,N_12416);
nor U12635 (N_12635,N_12443,N_12427);
nor U12636 (N_12636,N_12469,N_12564);
nor U12637 (N_12637,N_12582,N_12439);
or U12638 (N_12638,N_12576,N_12448);
or U12639 (N_12639,N_12471,N_12464);
and U12640 (N_12640,N_12444,N_12512);
and U12641 (N_12641,N_12586,N_12480);
nand U12642 (N_12642,N_12533,N_12490);
or U12643 (N_12643,N_12468,N_12465);
or U12644 (N_12644,N_12547,N_12412);
nand U12645 (N_12645,N_12525,N_12567);
nand U12646 (N_12646,N_12425,N_12572);
nor U12647 (N_12647,N_12442,N_12506);
nor U12648 (N_12648,N_12456,N_12507);
nor U12649 (N_12649,N_12452,N_12495);
or U12650 (N_12650,N_12479,N_12488);
nand U12651 (N_12651,N_12554,N_12447);
nor U12652 (N_12652,N_12557,N_12434);
nand U12653 (N_12653,N_12509,N_12430);
or U12654 (N_12654,N_12573,N_12537);
nor U12655 (N_12655,N_12529,N_12570);
and U12656 (N_12656,N_12493,N_12596);
nand U12657 (N_12657,N_12410,N_12474);
and U12658 (N_12658,N_12522,N_12594);
nor U12659 (N_12659,N_12565,N_12563);
nor U12660 (N_12660,N_12550,N_12462);
nand U12661 (N_12661,N_12580,N_12486);
nand U12662 (N_12662,N_12417,N_12523);
and U12663 (N_12663,N_12501,N_12497);
nor U12664 (N_12664,N_12411,N_12589);
nand U12665 (N_12665,N_12451,N_12461);
or U12666 (N_12666,N_12559,N_12450);
xor U12667 (N_12667,N_12441,N_12455);
nand U12668 (N_12668,N_12575,N_12569);
nand U12669 (N_12669,N_12504,N_12431);
nor U12670 (N_12670,N_12463,N_12457);
nand U12671 (N_12671,N_12403,N_12526);
nor U12672 (N_12672,N_12481,N_12521);
and U12673 (N_12673,N_12422,N_12561);
and U12674 (N_12674,N_12542,N_12538);
xor U12675 (N_12675,N_12498,N_12515);
nor U12676 (N_12676,N_12520,N_12513);
nor U12677 (N_12677,N_12482,N_12524);
nor U12678 (N_12678,N_12558,N_12449);
and U12679 (N_12679,N_12549,N_12426);
nor U12680 (N_12680,N_12503,N_12406);
nand U12681 (N_12681,N_12568,N_12571);
or U12682 (N_12682,N_12540,N_12505);
and U12683 (N_12683,N_12466,N_12407);
nor U12684 (N_12684,N_12487,N_12527);
nor U12685 (N_12685,N_12544,N_12556);
nor U12686 (N_12686,N_12591,N_12532);
or U12687 (N_12687,N_12597,N_12551);
and U12688 (N_12688,N_12440,N_12555);
and U12689 (N_12689,N_12485,N_12483);
nor U12690 (N_12690,N_12508,N_12595);
and U12691 (N_12691,N_12566,N_12579);
nor U12692 (N_12692,N_12408,N_12419);
or U12693 (N_12693,N_12592,N_12400);
or U12694 (N_12694,N_12405,N_12585);
nor U12695 (N_12695,N_12536,N_12475);
nand U12696 (N_12696,N_12476,N_12541);
nand U12697 (N_12697,N_12432,N_12598);
nand U12698 (N_12698,N_12436,N_12459);
nand U12699 (N_12699,N_12473,N_12578);
or U12700 (N_12700,N_12530,N_12567);
and U12701 (N_12701,N_12479,N_12485);
nor U12702 (N_12702,N_12464,N_12577);
nand U12703 (N_12703,N_12412,N_12436);
nand U12704 (N_12704,N_12571,N_12442);
nor U12705 (N_12705,N_12558,N_12478);
nand U12706 (N_12706,N_12515,N_12536);
nor U12707 (N_12707,N_12420,N_12542);
or U12708 (N_12708,N_12509,N_12598);
or U12709 (N_12709,N_12477,N_12538);
and U12710 (N_12710,N_12589,N_12553);
and U12711 (N_12711,N_12539,N_12528);
and U12712 (N_12712,N_12469,N_12572);
and U12713 (N_12713,N_12531,N_12557);
nand U12714 (N_12714,N_12402,N_12443);
nand U12715 (N_12715,N_12535,N_12547);
and U12716 (N_12716,N_12417,N_12546);
nor U12717 (N_12717,N_12477,N_12411);
nor U12718 (N_12718,N_12541,N_12434);
and U12719 (N_12719,N_12517,N_12416);
nand U12720 (N_12720,N_12558,N_12505);
nor U12721 (N_12721,N_12547,N_12467);
nand U12722 (N_12722,N_12511,N_12578);
or U12723 (N_12723,N_12580,N_12465);
and U12724 (N_12724,N_12463,N_12578);
nor U12725 (N_12725,N_12472,N_12423);
and U12726 (N_12726,N_12555,N_12485);
nor U12727 (N_12727,N_12419,N_12502);
nand U12728 (N_12728,N_12457,N_12572);
or U12729 (N_12729,N_12487,N_12504);
nor U12730 (N_12730,N_12520,N_12477);
nor U12731 (N_12731,N_12516,N_12475);
nand U12732 (N_12732,N_12515,N_12458);
and U12733 (N_12733,N_12587,N_12555);
nand U12734 (N_12734,N_12578,N_12501);
nand U12735 (N_12735,N_12523,N_12447);
and U12736 (N_12736,N_12460,N_12417);
or U12737 (N_12737,N_12407,N_12574);
nor U12738 (N_12738,N_12415,N_12476);
and U12739 (N_12739,N_12428,N_12578);
nand U12740 (N_12740,N_12460,N_12406);
or U12741 (N_12741,N_12464,N_12547);
or U12742 (N_12742,N_12583,N_12480);
nand U12743 (N_12743,N_12574,N_12592);
or U12744 (N_12744,N_12545,N_12462);
nor U12745 (N_12745,N_12558,N_12576);
and U12746 (N_12746,N_12440,N_12594);
and U12747 (N_12747,N_12536,N_12491);
nor U12748 (N_12748,N_12428,N_12564);
nor U12749 (N_12749,N_12543,N_12594);
or U12750 (N_12750,N_12598,N_12531);
nand U12751 (N_12751,N_12458,N_12459);
nand U12752 (N_12752,N_12436,N_12414);
nor U12753 (N_12753,N_12432,N_12463);
or U12754 (N_12754,N_12544,N_12488);
and U12755 (N_12755,N_12421,N_12567);
and U12756 (N_12756,N_12443,N_12489);
nor U12757 (N_12757,N_12498,N_12585);
nor U12758 (N_12758,N_12529,N_12476);
and U12759 (N_12759,N_12584,N_12569);
or U12760 (N_12760,N_12562,N_12484);
and U12761 (N_12761,N_12497,N_12538);
or U12762 (N_12762,N_12483,N_12552);
nor U12763 (N_12763,N_12588,N_12482);
nor U12764 (N_12764,N_12528,N_12527);
and U12765 (N_12765,N_12412,N_12449);
and U12766 (N_12766,N_12564,N_12565);
nor U12767 (N_12767,N_12539,N_12412);
nand U12768 (N_12768,N_12489,N_12552);
nand U12769 (N_12769,N_12547,N_12482);
or U12770 (N_12770,N_12542,N_12474);
nand U12771 (N_12771,N_12585,N_12597);
nand U12772 (N_12772,N_12569,N_12465);
or U12773 (N_12773,N_12554,N_12486);
and U12774 (N_12774,N_12487,N_12534);
nand U12775 (N_12775,N_12459,N_12443);
or U12776 (N_12776,N_12584,N_12473);
or U12777 (N_12777,N_12552,N_12410);
nand U12778 (N_12778,N_12480,N_12448);
nand U12779 (N_12779,N_12442,N_12551);
nand U12780 (N_12780,N_12571,N_12512);
and U12781 (N_12781,N_12465,N_12492);
nor U12782 (N_12782,N_12592,N_12467);
or U12783 (N_12783,N_12410,N_12419);
or U12784 (N_12784,N_12453,N_12544);
nand U12785 (N_12785,N_12555,N_12483);
or U12786 (N_12786,N_12507,N_12434);
nor U12787 (N_12787,N_12466,N_12435);
and U12788 (N_12788,N_12481,N_12492);
nor U12789 (N_12789,N_12452,N_12459);
nor U12790 (N_12790,N_12530,N_12514);
or U12791 (N_12791,N_12590,N_12420);
nor U12792 (N_12792,N_12585,N_12512);
nand U12793 (N_12793,N_12556,N_12486);
nor U12794 (N_12794,N_12430,N_12558);
or U12795 (N_12795,N_12534,N_12449);
nor U12796 (N_12796,N_12529,N_12462);
nand U12797 (N_12797,N_12409,N_12478);
nor U12798 (N_12798,N_12542,N_12497);
or U12799 (N_12799,N_12464,N_12415);
and U12800 (N_12800,N_12605,N_12742);
and U12801 (N_12801,N_12648,N_12751);
xnor U12802 (N_12802,N_12694,N_12700);
nor U12803 (N_12803,N_12602,N_12707);
or U12804 (N_12804,N_12761,N_12792);
nand U12805 (N_12805,N_12716,N_12632);
and U12806 (N_12806,N_12623,N_12755);
and U12807 (N_12807,N_12651,N_12631);
and U12808 (N_12808,N_12685,N_12671);
or U12809 (N_12809,N_12799,N_12609);
and U12810 (N_12810,N_12713,N_12699);
nor U12811 (N_12811,N_12692,N_12744);
or U12812 (N_12812,N_12783,N_12669);
nand U12813 (N_12813,N_12712,N_12679);
nand U12814 (N_12814,N_12601,N_12624);
or U12815 (N_12815,N_12794,N_12657);
nand U12816 (N_12816,N_12750,N_12677);
or U12817 (N_12817,N_12723,N_12776);
or U12818 (N_12818,N_12698,N_12680);
or U12819 (N_12819,N_12633,N_12606);
and U12820 (N_12820,N_12666,N_12620);
or U12821 (N_12821,N_12619,N_12722);
and U12822 (N_12822,N_12736,N_12687);
nand U12823 (N_12823,N_12718,N_12791);
nor U12824 (N_12824,N_12613,N_12787);
nand U12825 (N_12825,N_12610,N_12778);
nor U12826 (N_12826,N_12705,N_12661);
nor U12827 (N_12827,N_12749,N_12681);
xor U12828 (N_12828,N_12603,N_12703);
and U12829 (N_12829,N_12745,N_12793);
nand U12830 (N_12830,N_12764,N_12754);
or U12831 (N_12831,N_12762,N_12630);
or U12832 (N_12832,N_12690,N_12636);
nand U12833 (N_12833,N_12717,N_12688);
nand U12834 (N_12834,N_12654,N_12765);
or U12835 (N_12835,N_12789,N_12627);
or U12836 (N_12836,N_12719,N_12650);
and U12837 (N_12837,N_12752,N_12786);
nor U12838 (N_12838,N_12614,N_12638);
and U12839 (N_12839,N_12686,N_12766);
or U12840 (N_12840,N_12612,N_12797);
nand U12841 (N_12841,N_12714,N_12656);
or U12842 (N_12842,N_12740,N_12796);
and U12843 (N_12843,N_12760,N_12780);
nand U12844 (N_12844,N_12781,N_12709);
nand U12845 (N_12845,N_12611,N_12637);
nand U12846 (N_12846,N_12746,N_12658);
nor U12847 (N_12847,N_12726,N_12634);
nand U12848 (N_12848,N_12735,N_12670);
nor U12849 (N_12849,N_12642,N_12668);
or U12850 (N_12850,N_12663,N_12691);
or U12851 (N_12851,N_12774,N_12711);
or U12852 (N_12852,N_12617,N_12772);
and U12853 (N_12853,N_12758,N_12779);
or U12854 (N_12854,N_12770,N_12662);
nand U12855 (N_12855,N_12682,N_12706);
nand U12856 (N_12856,N_12635,N_12738);
nand U12857 (N_12857,N_12753,N_12622);
and U12858 (N_12858,N_12626,N_12728);
nand U12859 (N_12859,N_12710,N_12673);
and U12860 (N_12860,N_12616,N_12600);
or U12861 (N_12861,N_12678,N_12795);
nand U12862 (N_12862,N_12621,N_12756);
nand U12863 (N_12863,N_12704,N_12775);
and U12864 (N_12864,N_12696,N_12743);
nor U12865 (N_12865,N_12618,N_12628);
nor U12866 (N_12866,N_12615,N_12737);
nand U12867 (N_12867,N_12784,N_12767);
and U12868 (N_12868,N_12676,N_12683);
or U12869 (N_12869,N_12608,N_12646);
and U12870 (N_12870,N_12720,N_12689);
nor U12871 (N_12871,N_12724,N_12715);
and U12872 (N_12872,N_12732,N_12741);
xor U12873 (N_12873,N_12675,N_12645);
nand U12874 (N_12874,N_12708,N_12644);
nor U12875 (N_12875,N_12771,N_12729);
nand U12876 (N_12876,N_12643,N_12730);
and U12877 (N_12877,N_12748,N_12727);
nor U12878 (N_12878,N_12667,N_12647);
nand U12879 (N_12879,N_12672,N_12625);
nand U12880 (N_12880,N_12785,N_12664);
nor U12881 (N_12881,N_12721,N_12763);
nand U12882 (N_12882,N_12629,N_12701);
nor U12883 (N_12883,N_12759,N_12702);
nand U12884 (N_12884,N_12693,N_12695);
nor U12885 (N_12885,N_12604,N_12697);
nand U12886 (N_12886,N_12773,N_12769);
nor U12887 (N_12887,N_12684,N_12768);
nor U12888 (N_12888,N_12649,N_12660);
and U12889 (N_12889,N_12798,N_12607);
nor U12890 (N_12890,N_12640,N_12739);
and U12891 (N_12891,N_12659,N_12665);
nor U12892 (N_12892,N_12639,N_12788);
xor U12893 (N_12893,N_12734,N_12652);
nor U12894 (N_12894,N_12653,N_12782);
or U12895 (N_12895,N_12757,N_12725);
and U12896 (N_12896,N_12733,N_12674);
nand U12897 (N_12897,N_12777,N_12731);
nor U12898 (N_12898,N_12747,N_12655);
and U12899 (N_12899,N_12790,N_12641);
nand U12900 (N_12900,N_12692,N_12776);
or U12901 (N_12901,N_12748,N_12704);
nor U12902 (N_12902,N_12679,N_12767);
nand U12903 (N_12903,N_12662,N_12715);
nand U12904 (N_12904,N_12689,N_12646);
or U12905 (N_12905,N_12704,N_12764);
or U12906 (N_12906,N_12731,N_12757);
nand U12907 (N_12907,N_12625,N_12782);
nand U12908 (N_12908,N_12790,N_12665);
nand U12909 (N_12909,N_12613,N_12605);
or U12910 (N_12910,N_12655,N_12716);
or U12911 (N_12911,N_12675,N_12777);
or U12912 (N_12912,N_12771,N_12631);
nand U12913 (N_12913,N_12791,N_12638);
and U12914 (N_12914,N_12677,N_12659);
or U12915 (N_12915,N_12683,N_12736);
or U12916 (N_12916,N_12708,N_12619);
and U12917 (N_12917,N_12672,N_12651);
nand U12918 (N_12918,N_12796,N_12602);
nand U12919 (N_12919,N_12760,N_12710);
and U12920 (N_12920,N_12699,N_12661);
and U12921 (N_12921,N_12668,N_12788);
nor U12922 (N_12922,N_12658,N_12692);
and U12923 (N_12923,N_12645,N_12796);
nand U12924 (N_12924,N_12753,N_12722);
nor U12925 (N_12925,N_12673,N_12760);
nor U12926 (N_12926,N_12790,N_12706);
xor U12927 (N_12927,N_12626,N_12664);
and U12928 (N_12928,N_12790,N_12780);
nand U12929 (N_12929,N_12733,N_12698);
nand U12930 (N_12930,N_12638,N_12636);
or U12931 (N_12931,N_12719,N_12798);
or U12932 (N_12932,N_12674,N_12714);
or U12933 (N_12933,N_12717,N_12663);
and U12934 (N_12934,N_12680,N_12780);
xor U12935 (N_12935,N_12635,N_12664);
nor U12936 (N_12936,N_12653,N_12798);
nor U12937 (N_12937,N_12773,N_12671);
and U12938 (N_12938,N_12724,N_12758);
nand U12939 (N_12939,N_12611,N_12774);
nor U12940 (N_12940,N_12638,N_12767);
or U12941 (N_12941,N_12690,N_12791);
or U12942 (N_12942,N_12779,N_12605);
or U12943 (N_12943,N_12629,N_12617);
nor U12944 (N_12944,N_12790,N_12759);
and U12945 (N_12945,N_12637,N_12780);
nand U12946 (N_12946,N_12703,N_12624);
nand U12947 (N_12947,N_12634,N_12659);
nand U12948 (N_12948,N_12648,N_12676);
nor U12949 (N_12949,N_12745,N_12740);
and U12950 (N_12950,N_12651,N_12794);
nand U12951 (N_12951,N_12784,N_12636);
and U12952 (N_12952,N_12635,N_12714);
nor U12953 (N_12953,N_12789,N_12658);
nor U12954 (N_12954,N_12630,N_12777);
or U12955 (N_12955,N_12745,N_12744);
xor U12956 (N_12956,N_12746,N_12646);
nand U12957 (N_12957,N_12727,N_12718);
nor U12958 (N_12958,N_12784,N_12608);
nor U12959 (N_12959,N_12737,N_12678);
and U12960 (N_12960,N_12680,N_12736);
or U12961 (N_12961,N_12795,N_12642);
and U12962 (N_12962,N_12768,N_12637);
or U12963 (N_12963,N_12641,N_12743);
nor U12964 (N_12964,N_12798,N_12698);
nor U12965 (N_12965,N_12731,N_12729);
nor U12966 (N_12966,N_12742,N_12793);
nand U12967 (N_12967,N_12734,N_12761);
and U12968 (N_12968,N_12674,N_12775);
or U12969 (N_12969,N_12644,N_12658);
nor U12970 (N_12970,N_12628,N_12656);
nor U12971 (N_12971,N_12725,N_12782);
or U12972 (N_12972,N_12609,N_12759);
nand U12973 (N_12973,N_12714,N_12682);
or U12974 (N_12974,N_12775,N_12785);
or U12975 (N_12975,N_12766,N_12724);
nand U12976 (N_12976,N_12635,N_12666);
nor U12977 (N_12977,N_12623,N_12719);
nand U12978 (N_12978,N_12634,N_12799);
nor U12979 (N_12979,N_12671,N_12738);
nand U12980 (N_12980,N_12629,N_12778);
nand U12981 (N_12981,N_12688,N_12774);
or U12982 (N_12982,N_12743,N_12738);
nor U12983 (N_12983,N_12798,N_12759);
nor U12984 (N_12984,N_12645,N_12673);
or U12985 (N_12985,N_12795,N_12754);
and U12986 (N_12986,N_12659,N_12638);
nor U12987 (N_12987,N_12685,N_12718);
nand U12988 (N_12988,N_12764,N_12791);
nand U12989 (N_12989,N_12724,N_12753);
or U12990 (N_12990,N_12692,N_12625);
nand U12991 (N_12991,N_12664,N_12769);
nand U12992 (N_12992,N_12763,N_12779);
or U12993 (N_12993,N_12791,N_12729);
nor U12994 (N_12994,N_12697,N_12701);
nand U12995 (N_12995,N_12612,N_12673);
nor U12996 (N_12996,N_12796,N_12750);
nor U12997 (N_12997,N_12636,N_12613);
or U12998 (N_12998,N_12790,N_12738);
and U12999 (N_12999,N_12729,N_12694);
or U13000 (N_13000,N_12955,N_12801);
nor U13001 (N_13001,N_12823,N_12919);
nand U13002 (N_13002,N_12877,N_12904);
xor U13003 (N_13003,N_12918,N_12997);
and U13004 (N_13004,N_12963,N_12950);
nor U13005 (N_13005,N_12864,N_12933);
nor U13006 (N_13006,N_12800,N_12935);
nand U13007 (N_13007,N_12913,N_12893);
and U13008 (N_13008,N_12829,N_12859);
and U13009 (N_13009,N_12890,N_12951);
or U13010 (N_13010,N_12966,N_12813);
nor U13011 (N_13011,N_12876,N_12880);
nand U13012 (N_13012,N_12807,N_12860);
nand U13013 (N_13013,N_12803,N_12920);
or U13014 (N_13014,N_12934,N_12802);
nand U13015 (N_13015,N_12806,N_12892);
nor U13016 (N_13016,N_12960,N_12992);
and U13017 (N_13017,N_12852,N_12957);
nand U13018 (N_13018,N_12910,N_12842);
and U13019 (N_13019,N_12894,N_12830);
and U13020 (N_13020,N_12871,N_12971);
or U13021 (N_13021,N_12975,N_12867);
nor U13022 (N_13022,N_12968,N_12887);
nand U13023 (N_13023,N_12926,N_12909);
nand U13024 (N_13024,N_12828,N_12949);
and U13025 (N_13025,N_12902,N_12814);
and U13026 (N_13026,N_12879,N_12982);
and U13027 (N_13027,N_12977,N_12845);
and U13028 (N_13028,N_12943,N_12849);
xor U13029 (N_13029,N_12939,N_12923);
and U13030 (N_13030,N_12886,N_12855);
nor U13031 (N_13031,N_12999,N_12872);
nand U13032 (N_13032,N_12907,N_12898);
and U13033 (N_13033,N_12932,N_12917);
nand U13034 (N_13034,N_12965,N_12834);
nand U13035 (N_13035,N_12967,N_12969);
nand U13036 (N_13036,N_12873,N_12838);
nor U13037 (N_13037,N_12888,N_12847);
or U13038 (N_13038,N_12991,N_12836);
and U13039 (N_13039,N_12862,N_12973);
and U13040 (N_13040,N_12974,N_12869);
nor U13041 (N_13041,N_12941,N_12812);
or U13042 (N_13042,N_12953,N_12911);
and U13043 (N_13043,N_12856,N_12927);
nor U13044 (N_13044,N_12840,N_12865);
nand U13045 (N_13045,N_12897,N_12881);
and U13046 (N_13046,N_12866,N_12874);
or U13047 (N_13047,N_12915,N_12922);
or U13048 (N_13048,N_12956,N_12818);
nand U13049 (N_13049,N_12850,N_12998);
nand U13050 (N_13050,N_12868,N_12895);
and U13051 (N_13051,N_12846,N_12905);
nand U13052 (N_13052,N_12958,N_12924);
nand U13053 (N_13053,N_12938,N_12844);
xnor U13054 (N_13054,N_12854,N_12899);
xnor U13055 (N_13055,N_12815,N_12821);
nand U13056 (N_13056,N_12947,N_12891);
nand U13057 (N_13057,N_12970,N_12816);
and U13058 (N_13058,N_12901,N_12983);
nand U13059 (N_13059,N_12896,N_12908);
or U13060 (N_13060,N_12839,N_12944);
or U13061 (N_13061,N_12995,N_12930);
and U13062 (N_13062,N_12835,N_12978);
nor U13063 (N_13063,N_12805,N_12870);
nand U13064 (N_13064,N_12851,N_12831);
nor U13065 (N_13065,N_12962,N_12996);
and U13066 (N_13066,N_12979,N_12980);
nor U13067 (N_13067,N_12952,N_12981);
and U13068 (N_13068,N_12972,N_12961);
or U13069 (N_13069,N_12804,N_12921);
or U13070 (N_13070,N_12937,N_12837);
or U13071 (N_13071,N_12843,N_12817);
nand U13072 (N_13072,N_12861,N_12841);
nor U13073 (N_13073,N_12878,N_12900);
or U13074 (N_13074,N_12990,N_12925);
or U13075 (N_13075,N_12857,N_12882);
nand U13076 (N_13076,N_12848,N_12875);
and U13077 (N_13077,N_12914,N_12994);
nor U13078 (N_13078,N_12825,N_12819);
nand U13079 (N_13079,N_12827,N_12858);
nand U13080 (N_13080,N_12928,N_12986);
nor U13081 (N_13081,N_12929,N_12889);
or U13082 (N_13082,N_12954,N_12826);
or U13083 (N_13083,N_12987,N_12820);
nand U13084 (N_13084,N_12912,N_12984);
and U13085 (N_13085,N_12811,N_12863);
and U13086 (N_13086,N_12985,N_12988);
and U13087 (N_13087,N_12959,N_12808);
nand U13088 (N_13088,N_12810,N_12906);
nor U13089 (N_13089,N_12940,N_12822);
nand U13090 (N_13090,N_12903,N_12989);
nand U13091 (N_13091,N_12824,N_12931);
and U13092 (N_13092,N_12993,N_12942);
and U13093 (N_13093,N_12976,N_12884);
xor U13094 (N_13094,N_12936,N_12964);
nand U13095 (N_13095,N_12885,N_12883);
and U13096 (N_13096,N_12809,N_12916);
and U13097 (N_13097,N_12833,N_12948);
nand U13098 (N_13098,N_12832,N_12946);
and U13099 (N_13099,N_12853,N_12945);
nor U13100 (N_13100,N_12865,N_12800);
or U13101 (N_13101,N_12857,N_12982);
nor U13102 (N_13102,N_12896,N_12921);
nand U13103 (N_13103,N_12845,N_12973);
nor U13104 (N_13104,N_12872,N_12996);
and U13105 (N_13105,N_12825,N_12820);
and U13106 (N_13106,N_12856,N_12809);
or U13107 (N_13107,N_12924,N_12928);
nand U13108 (N_13108,N_12993,N_12804);
nand U13109 (N_13109,N_12899,N_12900);
nor U13110 (N_13110,N_12826,N_12840);
or U13111 (N_13111,N_12892,N_12815);
nand U13112 (N_13112,N_12975,N_12913);
or U13113 (N_13113,N_12916,N_12842);
or U13114 (N_13114,N_12993,N_12938);
and U13115 (N_13115,N_12827,N_12856);
nand U13116 (N_13116,N_12958,N_12995);
or U13117 (N_13117,N_12853,N_12911);
or U13118 (N_13118,N_12929,N_12854);
nand U13119 (N_13119,N_12982,N_12873);
or U13120 (N_13120,N_12830,N_12941);
and U13121 (N_13121,N_12940,N_12949);
or U13122 (N_13122,N_12937,N_12984);
nand U13123 (N_13123,N_12893,N_12898);
or U13124 (N_13124,N_12851,N_12942);
or U13125 (N_13125,N_12867,N_12947);
or U13126 (N_13126,N_12821,N_12991);
and U13127 (N_13127,N_12893,N_12895);
nor U13128 (N_13128,N_12885,N_12803);
and U13129 (N_13129,N_12963,N_12937);
and U13130 (N_13130,N_12978,N_12812);
nand U13131 (N_13131,N_12917,N_12910);
nor U13132 (N_13132,N_12945,N_12893);
nand U13133 (N_13133,N_12884,N_12935);
nand U13134 (N_13134,N_12893,N_12849);
and U13135 (N_13135,N_12899,N_12851);
and U13136 (N_13136,N_12816,N_12858);
and U13137 (N_13137,N_12985,N_12904);
nor U13138 (N_13138,N_12963,N_12925);
nand U13139 (N_13139,N_12857,N_12807);
nand U13140 (N_13140,N_12855,N_12873);
and U13141 (N_13141,N_12879,N_12977);
or U13142 (N_13142,N_12924,N_12836);
and U13143 (N_13143,N_12896,N_12855);
nand U13144 (N_13144,N_12829,N_12944);
or U13145 (N_13145,N_12836,N_12813);
or U13146 (N_13146,N_12894,N_12998);
or U13147 (N_13147,N_12831,N_12975);
or U13148 (N_13148,N_12840,N_12944);
nor U13149 (N_13149,N_12832,N_12806);
nand U13150 (N_13150,N_12886,N_12927);
or U13151 (N_13151,N_12975,N_12969);
nor U13152 (N_13152,N_12886,N_12918);
nand U13153 (N_13153,N_12881,N_12904);
nand U13154 (N_13154,N_12831,N_12943);
and U13155 (N_13155,N_12879,N_12899);
or U13156 (N_13156,N_12990,N_12819);
or U13157 (N_13157,N_12884,N_12941);
nand U13158 (N_13158,N_12818,N_12847);
and U13159 (N_13159,N_12800,N_12828);
and U13160 (N_13160,N_12924,N_12919);
nand U13161 (N_13161,N_12949,N_12977);
or U13162 (N_13162,N_12993,N_12855);
and U13163 (N_13163,N_12945,N_12946);
and U13164 (N_13164,N_12893,N_12878);
xor U13165 (N_13165,N_12841,N_12851);
or U13166 (N_13166,N_12983,N_12973);
or U13167 (N_13167,N_12821,N_12877);
or U13168 (N_13168,N_12838,N_12977);
and U13169 (N_13169,N_12985,N_12971);
nand U13170 (N_13170,N_12814,N_12875);
or U13171 (N_13171,N_12916,N_12822);
nand U13172 (N_13172,N_12970,N_12942);
nor U13173 (N_13173,N_12857,N_12908);
xnor U13174 (N_13174,N_12947,N_12806);
and U13175 (N_13175,N_12840,N_12821);
or U13176 (N_13176,N_12812,N_12922);
nand U13177 (N_13177,N_12963,N_12991);
and U13178 (N_13178,N_12826,N_12820);
nor U13179 (N_13179,N_12908,N_12859);
xor U13180 (N_13180,N_12923,N_12947);
and U13181 (N_13181,N_12921,N_12840);
nand U13182 (N_13182,N_12915,N_12944);
or U13183 (N_13183,N_12820,N_12942);
or U13184 (N_13184,N_12801,N_12800);
and U13185 (N_13185,N_12830,N_12949);
nor U13186 (N_13186,N_12892,N_12989);
and U13187 (N_13187,N_12988,N_12936);
nor U13188 (N_13188,N_12801,N_12959);
nor U13189 (N_13189,N_12885,N_12927);
nand U13190 (N_13190,N_12885,N_12876);
and U13191 (N_13191,N_12893,N_12835);
nor U13192 (N_13192,N_12956,N_12922);
xor U13193 (N_13193,N_12931,N_12920);
nor U13194 (N_13194,N_12820,N_12874);
nor U13195 (N_13195,N_12903,N_12981);
nor U13196 (N_13196,N_12971,N_12856);
and U13197 (N_13197,N_12982,N_12823);
nand U13198 (N_13198,N_12865,N_12892);
and U13199 (N_13199,N_12847,N_12803);
and U13200 (N_13200,N_13119,N_13142);
nor U13201 (N_13201,N_13056,N_13013);
and U13202 (N_13202,N_13109,N_13102);
nor U13203 (N_13203,N_13091,N_13055);
and U13204 (N_13204,N_13086,N_13011);
or U13205 (N_13205,N_13042,N_13189);
nand U13206 (N_13206,N_13149,N_13083);
and U13207 (N_13207,N_13124,N_13146);
nor U13208 (N_13208,N_13043,N_13152);
nor U13209 (N_13209,N_13089,N_13178);
or U13210 (N_13210,N_13001,N_13133);
and U13211 (N_13211,N_13075,N_13058);
or U13212 (N_13212,N_13132,N_13123);
nand U13213 (N_13213,N_13150,N_13161);
nand U13214 (N_13214,N_13034,N_13054);
nand U13215 (N_13215,N_13108,N_13144);
or U13216 (N_13216,N_13100,N_13047);
nor U13217 (N_13217,N_13045,N_13076);
and U13218 (N_13218,N_13014,N_13136);
nor U13219 (N_13219,N_13179,N_13046);
and U13220 (N_13220,N_13065,N_13067);
nand U13221 (N_13221,N_13092,N_13016);
nand U13222 (N_13222,N_13022,N_13195);
and U13223 (N_13223,N_13027,N_13156);
or U13224 (N_13224,N_13103,N_13191);
nor U13225 (N_13225,N_13105,N_13098);
or U13226 (N_13226,N_13033,N_13052);
or U13227 (N_13227,N_13019,N_13114);
nor U13228 (N_13228,N_13173,N_13188);
nand U13229 (N_13229,N_13162,N_13194);
or U13230 (N_13230,N_13115,N_13186);
nand U13231 (N_13231,N_13177,N_13127);
nor U13232 (N_13232,N_13020,N_13085);
and U13233 (N_13233,N_13131,N_13041);
nand U13234 (N_13234,N_13095,N_13106);
or U13235 (N_13235,N_13035,N_13082);
nor U13236 (N_13236,N_13097,N_13073);
nand U13237 (N_13237,N_13155,N_13079);
nor U13238 (N_13238,N_13074,N_13005);
nand U13239 (N_13239,N_13008,N_13064);
nand U13240 (N_13240,N_13117,N_13000);
and U13241 (N_13241,N_13198,N_13190);
nor U13242 (N_13242,N_13071,N_13057);
and U13243 (N_13243,N_13025,N_13163);
nand U13244 (N_13244,N_13002,N_13110);
and U13245 (N_13245,N_13113,N_13143);
and U13246 (N_13246,N_13184,N_13187);
nor U13247 (N_13247,N_13037,N_13125);
and U13248 (N_13248,N_13126,N_13135);
and U13249 (N_13249,N_13015,N_13088);
and U13250 (N_13250,N_13066,N_13154);
nor U13251 (N_13251,N_13171,N_13138);
nand U13252 (N_13252,N_13199,N_13151);
nor U13253 (N_13253,N_13036,N_13157);
nand U13254 (N_13254,N_13006,N_13069);
or U13255 (N_13255,N_13050,N_13094);
nand U13256 (N_13256,N_13084,N_13175);
or U13257 (N_13257,N_13059,N_13120);
nand U13258 (N_13258,N_13077,N_13004);
nand U13259 (N_13259,N_13118,N_13101);
and U13260 (N_13260,N_13104,N_13018);
and U13261 (N_13261,N_13130,N_13026);
and U13262 (N_13262,N_13003,N_13140);
nand U13263 (N_13263,N_13061,N_13049);
or U13264 (N_13264,N_13172,N_13012);
nor U13265 (N_13265,N_13121,N_13159);
and U13266 (N_13266,N_13147,N_13145);
nor U13267 (N_13267,N_13166,N_13080);
or U13268 (N_13268,N_13023,N_13028);
or U13269 (N_13269,N_13134,N_13116);
or U13270 (N_13270,N_13167,N_13063);
or U13271 (N_13271,N_13111,N_13048);
nand U13272 (N_13272,N_13137,N_13182);
and U13273 (N_13273,N_13197,N_13176);
nor U13274 (N_13274,N_13090,N_13031);
nor U13275 (N_13275,N_13081,N_13129);
nor U13276 (N_13276,N_13044,N_13196);
nor U13277 (N_13277,N_13029,N_13053);
nor U13278 (N_13278,N_13141,N_13112);
and U13279 (N_13279,N_13107,N_13093);
and U13280 (N_13280,N_13038,N_13078);
nand U13281 (N_13281,N_13180,N_13039);
nand U13282 (N_13282,N_13040,N_13030);
nand U13283 (N_13283,N_13193,N_13072);
and U13284 (N_13284,N_13181,N_13051);
nand U13285 (N_13285,N_13021,N_13070);
xor U13286 (N_13286,N_13128,N_13174);
nand U13287 (N_13287,N_13096,N_13099);
and U13288 (N_13288,N_13160,N_13170);
nand U13289 (N_13289,N_13148,N_13007);
or U13290 (N_13290,N_13164,N_13192);
and U13291 (N_13291,N_13165,N_13158);
nor U13292 (N_13292,N_13024,N_13169);
nor U13293 (N_13293,N_13017,N_13183);
nand U13294 (N_13294,N_13168,N_13185);
or U13295 (N_13295,N_13032,N_13139);
and U13296 (N_13296,N_13010,N_13060);
nand U13297 (N_13297,N_13009,N_13153);
nand U13298 (N_13298,N_13068,N_13062);
and U13299 (N_13299,N_13087,N_13122);
and U13300 (N_13300,N_13032,N_13038);
xnor U13301 (N_13301,N_13099,N_13087);
nor U13302 (N_13302,N_13123,N_13190);
nor U13303 (N_13303,N_13104,N_13061);
or U13304 (N_13304,N_13180,N_13198);
nor U13305 (N_13305,N_13008,N_13132);
nand U13306 (N_13306,N_13064,N_13095);
nand U13307 (N_13307,N_13024,N_13083);
nand U13308 (N_13308,N_13098,N_13005);
nand U13309 (N_13309,N_13056,N_13034);
or U13310 (N_13310,N_13044,N_13182);
nor U13311 (N_13311,N_13188,N_13112);
nor U13312 (N_13312,N_13116,N_13179);
nor U13313 (N_13313,N_13035,N_13093);
or U13314 (N_13314,N_13116,N_13177);
or U13315 (N_13315,N_13081,N_13062);
nor U13316 (N_13316,N_13042,N_13187);
nor U13317 (N_13317,N_13153,N_13056);
and U13318 (N_13318,N_13189,N_13077);
and U13319 (N_13319,N_13160,N_13009);
and U13320 (N_13320,N_13192,N_13182);
and U13321 (N_13321,N_13198,N_13142);
nor U13322 (N_13322,N_13120,N_13085);
nand U13323 (N_13323,N_13008,N_13096);
or U13324 (N_13324,N_13166,N_13114);
and U13325 (N_13325,N_13099,N_13085);
nor U13326 (N_13326,N_13092,N_13024);
nor U13327 (N_13327,N_13143,N_13042);
nand U13328 (N_13328,N_13012,N_13097);
or U13329 (N_13329,N_13171,N_13128);
nor U13330 (N_13330,N_13103,N_13124);
or U13331 (N_13331,N_13169,N_13053);
nand U13332 (N_13332,N_13157,N_13055);
nor U13333 (N_13333,N_13007,N_13005);
and U13334 (N_13334,N_13091,N_13188);
nor U13335 (N_13335,N_13129,N_13072);
or U13336 (N_13336,N_13193,N_13082);
nor U13337 (N_13337,N_13021,N_13081);
nor U13338 (N_13338,N_13125,N_13036);
nand U13339 (N_13339,N_13186,N_13033);
nand U13340 (N_13340,N_13072,N_13059);
and U13341 (N_13341,N_13139,N_13116);
or U13342 (N_13342,N_13086,N_13095);
and U13343 (N_13343,N_13180,N_13042);
nand U13344 (N_13344,N_13186,N_13144);
and U13345 (N_13345,N_13173,N_13111);
nor U13346 (N_13346,N_13025,N_13079);
nor U13347 (N_13347,N_13104,N_13109);
or U13348 (N_13348,N_13040,N_13134);
nor U13349 (N_13349,N_13102,N_13067);
and U13350 (N_13350,N_13114,N_13006);
or U13351 (N_13351,N_13193,N_13128);
or U13352 (N_13352,N_13188,N_13013);
and U13353 (N_13353,N_13034,N_13154);
nor U13354 (N_13354,N_13013,N_13027);
nand U13355 (N_13355,N_13046,N_13015);
nor U13356 (N_13356,N_13116,N_13054);
and U13357 (N_13357,N_13067,N_13070);
or U13358 (N_13358,N_13068,N_13170);
nor U13359 (N_13359,N_13051,N_13066);
nor U13360 (N_13360,N_13126,N_13097);
or U13361 (N_13361,N_13048,N_13036);
and U13362 (N_13362,N_13046,N_13160);
nor U13363 (N_13363,N_13047,N_13187);
or U13364 (N_13364,N_13077,N_13142);
nand U13365 (N_13365,N_13103,N_13080);
nor U13366 (N_13366,N_13097,N_13136);
and U13367 (N_13367,N_13046,N_13170);
and U13368 (N_13368,N_13062,N_13182);
or U13369 (N_13369,N_13108,N_13121);
nor U13370 (N_13370,N_13033,N_13083);
nor U13371 (N_13371,N_13164,N_13095);
nand U13372 (N_13372,N_13034,N_13149);
or U13373 (N_13373,N_13125,N_13153);
or U13374 (N_13374,N_13076,N_13054);
or U13375 (N_13375,N_13021,N_13118);
nor U13376 (N_13376,N_13003,N_13024);
or U13377 (N_13377,N_13102,N_13020);
or U13378 (N_13378,N_13064,N_13048);
and U13379 (N_13379,N_13162,N_13190);
and U13380 (N_13380,N_13011,N_13162);
or U13381 (N_13381,N_13186,N_13027);
nor U13382 (N_13382,N_13085,N_13017);
or U13383 (N_13383,N_13131,N_13124);
nor U13384 (N_13384,N_13147,N_13105);
or U13385 (N_13385,N_13150,N_13140);
and U13386 (N_13386,N_13141,N_13145);
nand U13387 (N_13387,N_13041,N_13036);
and U13388 (N_13388,N_13058,N_13194);
nor U13389 (N_13389,N_13043,N_13073);
nand U13390 (N_13390,N_13197,N_13078);
or U13391 (N_13391,N_13162,N_13023);
nand U13392 (N_13392,N_13077,N_13165);
nor U13393 (N_13393,N_13178,N_13100);
nand U13394 (N_13394,N_13125,N_13064);
nor U13395 (N_13395,N_13054,N_13105);
nor U13396 (N_13396,N_13060,N_13145);
and U13397 (N_13397,N_13153,N_13104);
nand U13398 (N_13398,N_13167,N_13104);
nor U13399 (N_13399,N_13178,N_13197);
nand U13400 (N_13400,N_13206,N_13349);
nor U13401 (N_13401,N_13253,N_13259);
nor U13402 (N_13402,N_13254,N_13267);
nand U13403 (N_13403,N_13221,N_13227);
nor U13404 (N_13404,N_13292,N_13357);
and U13405 (N_13405,N_13204,N_13309);
and U13406 (N_13406,N_13249,N_13340);
nand U13407 (N_13407,N_13212,N_13304);
and U13408 (N_13408,N_13232,N_13243);
nand U13409 (N_13409,N_13203,N_13286);
nor U13410 (N_13410,N_13321,N_13308);
nand U13411 (N_13411,N_13345,N_13250);
nand U13412 (N_13412,N_13248,N_13266);
or U13413 (N_13413,N_13397,N_13343);
or U13414 (N_13414,N_13277,N_13202);
and U13415 (N_13415,N_13335,N_13242);
and U13416 (N_13416,N_13237,N_13394);
nand U13417 (N_13417,N_13228,N_13235);
nand U13418 (N_13418,N_13337,N_13294);
nor U13419 (N_13419,N_13222,N_13236);
and U13420 (N_13420,N_13284,N_13246);
and U13421 (N_13421,N_13334,N_13208);
nor U13422 (N_13422,N_13366,N_13320);
or U13423 (N_13423,N_13219,N_13326);
nor U13424 (N_13424,N_13365,N_13239);
nand U13425 (N_13425,N_13281,N_13378);
or U13426 (N_13426,N_13262,N_13234);
or U13427 (N_13427,N_13319,N_13325);
and U13428 (N_13428,N_13307,N_13328);
nor U13429 (N_13429,N_13216,N_13261);
nor U13430 (N_13430,N_13391,N_13229);
nand U13431 (N_13431,N_13329,N_13360);
nand U13432 (N_13432,N_13348,N_13382);
and U13433 (N_13433,N_13347,N_13257);
or U13434 (N_13434,N_13293,N_13217);
nand U13435 (N_13435,N_13385,N_13392);
nor U13436 (N_13436,N_13218,N_13388);
or U13437 (N_13437,N_13355,N_13240);
nor U13438 (N_13438,N_13341,N_13226);
and U13439 (N_13439,N_13295,N_13361);
and U13440 (N_13440,N_13374,N_13386);
and U13441 (N_13441,N_13332,N_13214);
and U13442 (N_13442,N_13356,N_13273);
nand U13443 (N_13443,N_13280,N_13323);
or U13444 (N_13444,N_13396,N_13313);
and U13445 (N_13445,N_13245,N_13367);
and U13446 (N_13446,N_13285,N_13258);
and U13447 (N_13447,N_13354,N_13271);
nor U13448 (N_13448,N_13230,N_13370);
nor U13449 (N_13449,N_13324,N_13389);
and U13450 (N_13450,N_13223,N_13279);
or U13451 (N_13451,N_13220,N_13398);
nand U13452 (N_13452,N_13299,N_13359);
or U13453 (N_13453,N_13376,N_13336);
nor U13454 (N_13454,N_13312,N_13282);
nor U13455 (N_13455,N_13290,N_13200);
nand U13456 (N_13456,N_13352,N_13265);
nor U13457 (N_13457,N_13231,N_13283);
nand U13458 (N_13458,N_13210,N_13314);
or U13459 (N_13459,N_13333,N_13233);
nor U13460 (N_13460,N_13207,N_13375);
and U13461 (N_13461,N_13368,N_13272);
or U13462 (N_13462,N_13316,N_13384);
and U13463 (N_13463,N_13330,N_13275);
nor U13464 (N_13464,N_13264,N_13393);
and U13465 (N_13465,N_13225,N_13296);
nand U13466 (N_13466,N_13276,N_13351);
or U13467 (N_13467,N_13346,N_13291);
nor U13468 (N_13468,N_13274,N_13209);
nand U13469 (N_13469,N_13390,N_13377);
nor U13470 (N_13470,N_13288,N_13251);
nand U13471 (N_13471,N_13301,N_13270);
nand U13472 (N_13472,N_13302,N_13269);
and U13473 (N_13473,N_13303,N_13252);
nand U13474 (N_13474,N_13278,N_13289);
or U13475 (N_13475,N_13298,N_13371);
and U13476 (N_13476,N_13383,N_13362);
nand U13477 (N_13477,N_13379,N_13317);
or U13478 (N_13478,N_13350,N_13255);
nand U13479 (N_13479,N_13287,N_13315);
nand U13480 (N_13480,N_13247,N_13305);
nand U13481 (N_13481,N_13311,N_13256);
and U13482 (N_13482,N_13358,N_13263);
and U13483 (N_13483,N_13310,N_13205);
or U13484 (N_13484,N_13268,N_13306);
or U13485 (N_13485,N_13381,N_13201);
and U13486 (N_13486,N_13297,N_13260);
and U13487 (N_13487,N_13372,N_13353);
nor U13488 (N_13488,N_13327,N_13238);
or U13489 (N_13489,N_13395,N_13363);
nand U13490 (N_13490,N_13344,N_13244);
nand U13491 (N_13491,N_13331,N_13399);
and U13492 (N_13492,N_13224,N_13380);
nor U13493 (N_13493,N_13339,N_13364);
and U13494 (N_13494,N_13373,N_13322);
or U13495 (N_13495,N_13300,N_13213);
and U13496 (N_13496,N_13387,N_13369);
and U13497 (N_13497,N_13338,N_13241);
nor U13498 (N_13498,N_13318,N_13215);
or U13499 (N_13499,N_13342,N_13211);
nand U13500 (N_13500,N_13254,N_13231);
or U13501 (N_13501,N_13371,N_13254);
nand U13502 (N_13502,N_13370,N_13217);
or U13503 (N_13503,N_13351,N_13326);
nand U13504 (N_13504,N_13392,N_13307);
and U13505 (N_13505,N_13354,N_13254);
nand U13506 (N_13506,N_13358,N_13261);
nor U13507 (N_13507,N_13213,N_13295);
nor U13508 (N_13508,N_13206,N_13262);
or U13509 (N_13509,N_13397,N_13216);
or U13510 (N_13510,N_13285,N_13326);
nand U13511 (N_13511,N_13328,N_13292);
and U13512 (N_13512,N_13300,N_13336);
and U13513 (N_13513,N_13261,N_13389);
and U13514 (N_13514,N_13341,N_13369);
and U13515 (N_13515,N_13261,N_13322);
nor U13516 (N_13516,N_13385,N_13253);
nor U13517 (N_13517,N_13234,N_13383);
or U13518 (N_13518,N_13395,N_13322);
nand U13519 (N_13519,N_13342,N_13276);
or U13520 (N_13520,N_13288,N_13339);
nand U13521 (N_13521,N_13335,N_13226);
nor U13522 (N_13522,N_13207,N_13333);
or U13523 (N_13523,N_13342,N_13248);
and U13524 (N_13524,N_13253,N_13210);
nor U13525 (N_13525,N_13256,N_13242);
and U13526 (N_13526,N_13240,N_13239);
nor U13527 (N_13527,N_13336,N_13294);
nand U13528 (N_13528,N_13273,N_13269);
nor U13529 (N_13529,N_13295,N_13328);
nand U13530 (N_13530,N_13382,N_13300);
or U13531 (N_13531,N_13360,N_13287);
and U13532 (N_13532,N_13272,N_13334);
nor U13533 (N_13533,N_13396,N_13364);
nor U13534 (N_13534,N_13384,N_13244);
nand U13535 (N_13535,N_13327,N_13323);
or U13536 (N_13536,N_13225,N_13299);
or U13537 (N_13537,N_13259,N_13256);
nand U13538 (N_13538,N_13321,N_13226);
and U13539 (N_13539,N_13239,N_13224);
nand U13540 (N_13540,N_13363,N_13337);
nor U13541 (N_13541,N_13230,N_13315);
or U13542 (N_13542,N_13227,N_13282);
nor U13543 (N_13543,N_13201,N_13397);
nand U13544 (N_13544,N_13280,N_13251);
nor U13545 (N_13545,N_13293,N_13223);
and U13546 (N_13546,N_13233,N_13337);
and U13547 (N_13547,N_13251,N_13342);
and U13548 (N_13548,N_13236,N_13293);
nand U13549 (N_13549,N_13329,N_13290);
nand U13550 (N_13550,N_13370,N_13391);
nand U13551 (N_13551,N_13382,N_13373);
and U13552 (N_13552,N_13300,N_13374);
or U13553 (N_13553,N_13396,N_13229);
nor U13554 (N_13554,N_13248,N_13281);
nand U13555 (N_13555,N_13356,N_13283);
nor U13556 (N_13556,N_13380,N_13393);
or U13557 (N_13557,N_13315,N_13320);
and U13558 (N_13558,N_13354,N_13326);
or U13559 (N_13559,N_13321,N_13251);
and U13560 (N_13560,N_13315,N_13265);
nand U13561 (N_13561,N_13238,N_13320);
nand U13562 (N_13562,N_13216,N_13289);
nor U13563 (N_13563,N_13227,N_13349);
and U13564 (N_13564,N_13230,N_13374);
and U13565 (N_13565,N_13249,N_13269);
and U13566 (N_13566,N_13224,N_13347);
or U13567 (N_13567,N_13304,N_13331);
or U13568 (N_13568,N_13233,N_13269);
and U13569 (N_13569,N_13225,N_13387);
nand U13570 (N_13570,N_13303,N_13351);
nor U13571 (N_13571,N_13282,N_13228);
or U13572 (N_13572,N_13380,N_13351);
nor U13573 (N_13573,N_13240,N_13255);
or U13574 (N_13574,N_13218,N_13210);
nand U13575 (N_13575,N_13287,N_13345);
nor U13576 (N_13576,N_13353,N_13289);
nor U13577 (N_13577,N_13382,N_13313);
and U13578 (N_13578,N_13277,N_13355);
and U13579 (N_13579,N_13268,N_13262);
or U13580 (N_13580,N_13343,N_13248);
and U13581 (N_13581,N_13228,N_13250);
or U13582 (N_13582,N_13259,N_13322);
nand U13583 (N_13583,N_13229,N_13326);
or U13584 (N_13584,N_13245,N_13286);
nand U13585 (N_13585,N_13326,N_13366);
nand U13586 (N_13586,N_13245,N_13269);
and U13587 (N_13587,N_13288,N_13303);
nand U13588 (N_13588,N_13388,N_13221);
or U13589 (N_13589,N_13313,N_13278);
or U13590 (N_13590,N_13231,N_13271);
nor U13591 (N_13591,N_13265,N_13234);
and U13592 (N_13592,N_13380,N_13299);
and U13593 (N_13593,N_13204,N_13364);
nor U13594 (N_13594,N_13335,N_13316);
and U13595 (N_13595,N_13292,N_13225);
nand U13596 (N_13596,N_13286,N_13262);
nand U13597 (N_13597,N_13377,N_13209);
nor U13598 (N_13598,N_13306,N_13305);
nor U13599 (N_13599,N_13398,N_13320);
or U13600 (N_13600,N_13484,N_13566);
nor U13601 (N_13601,N_13456,N_13490);
nand U13602 (N_13602,N_13538,N_13513);
or U13603 (N_13603,N_13545,N_13477);
and U13604 (N_13604,N_13596,N_13533);
nand U13605 (N_13605,N_13542,N_13475);
xor U13606 (N_13606,N_13585,N_13564);
and U13607 (N_13607,N_13402,N_13563);
nand U13608 (N_13608,N_13537,N_13559);
or U13609 (N_13609,N_13400,N_13519);
or U13610 (N_13610,N_13410,N_13429);
nor U13611 (N_13611,N_13425,N_13444);
nor U13612 (N_13612,N_13549,N_13448);
and U13613 (N_13613,N_13575,N_13462);
and U13614 (N_13614,N_13577,N_13547);
or U13615 (N_13615,N_13413,N_13569);
and U13616 (N_13616,N_13578,N_13481);
nand U13617 (N_13617,N_13594,N_13511);
nor U13618 (N_13618,N_13528,N_13408);
or U13619 (N_13619,N_13498,N_13555);
or U13620 (N_13620,N_13517,N_13487);
nor U13621 (N_13621,N_13554,N_13516);
or U13622 (N_13622,N_13436,N_13531);
or U13623 (N_13623,N_13534,N_13504);
and U13624 (N_13624,N_13532,N_13499);
or U13625 (N_13625,N_13454,N_13571);
nand U13626 (N_13626,N_13502,N_13421);
nor U13627 (N_13627,N_13597,N_13440);
nor U13628 (N_13628,N_13553,N_13485);
or U13629 (N_13629,N_13401,N_13595);
and U13630 (N_13630,N_13582,N_13535);
nor U13631 (N_13631,N_13403,N_13540);
nor U13632 (N_13632,N_13552,N_13407);
or U13633 (N_13633,N_13419,N_13438);
nor U13634 (N_13634,N_13491,N_13573);
and U13635 (N_13635,N_13591,N_13474);
and U13636 (N_13636,N_13526,N_13497);
nor U13637 (N_13637,N_13480,N_13509);
and U13638 (N_13638,N_13420,N_13417);
nor U13639 (N_13639,N_13459,N_13479);
nor U13640 (N_13640,N_13568,N_13579);
or U13641 (N_13641,N_13461,N_13524);
nor U13642 (N_13642,N_13576,N_13451);
and U13643 (N_13643,N_13476,N_13443);
nand U13644 (N_13644,N_13561,N_13494);
and U13645 (N_13645,N_13505,N_13503);
and U13646 (N_13646,N_13593,N_13469);
or U13647 (N_13647,N_13558,N_13515);
nor U13648 (N_13648,N_13464,N_13539);
nand U13649 (N_13649,N_13587,N_13529);
nor U13650 (N_13650,N_13508,N_13500);
nor U13651 (N_13651,N_13427,N_13586);
and U13652 (N_13652,N_13583,N_13589);
and U13653 (N_13653,N_13482,N_13424);
nand U13654 (N_13654,N_13458,N_13590);
nor U13655 (N_13655,N_13431,N_13453);
or U13656 (N_13656,N_13486,N_13409);
and U13657 (N_13657,N_13457,N_13536);
or U13658 (N_13658,N_13439,N_13478);
nand U13659 (N_13659,N_13557,N_13437);
nor U13660 (N_13660,N_13567,N_13510);
nand U13661 (N_13661,N_13404,N_13565);
nand U13662 (N_13662,N_13418,N_13460);
nor U13663 (N_13663,N_13506,N_13544);
or U13664 (N_13664,N_13541,N_13518);
nand U13665 (N_13665,N_13598,N_13446);
xor U13666 (N_13666,N_13525,N_13543);
nor U13667 (N_13667,N_13430,N_13496);
nand U13668 (N_13668,N_13562,N_13445);
or U13669 (N_13669,N_13570,N_13489);
or U13670 (N_13670,N_13514,N_13470);
nand U13671 (N_13671,N_13414,N_13455);
or U13672 (N_13672,N_13574,N_13467);
or U13673 (N_13673,N_13521,N_13452);
nor U13674 (N_13674,N_13501,N_13405);
or U13675 (N_13675,N_13522,N_13466);
or U13676 (N_13676,N_13551,N_13492);
and U13677 (N_13677,N_13422,N_13493);
nor U13678 (N_13678,N_13550,N_13411);
or U13679 (N_13679,N_13584,N_13435);
and U13680 (N_13680,N_13520,N_13432);
and U13681 (N_13681,N_13426,N_13495);
or U13682 (N_13682,N_13548,N_13415);
nand U13683 (N_13683,N_13488,N_13412);
and U13684 (N_13684,N_13588,N_13449);
nor U13685 (N_13685,N_13463,N_13473);
and U13686 (N_13686,N_13556,N_13472);
or U13687 (N_13687,N_13468,N_13580);
or U13688 (N_13688,N_13428,N_13572);
and U13689 (N_13689,N_13592,N_13447);
nor U13690 (N_13690,N_13546,N_13512);
or U13691 (N_13691,N_13450,N_13581);
or U13692 (N_13692,N_13406,N_13465);
or U13693 (N_13693,N_13527,N_13483);
nor U13694 (N_13694,N_13507,N_13530);
nand U13695 (N_13695,N_13423,N_13434);
and U13696 (N_13696,N_13471,N_13442);
xor U13697 (N_13697,N_13523,N_13599);
and U13698 (N_13698,N_13416,N_13433);
nand U13699 (N_13699,N_13441,N_13560);
and U13700 (N_13700,N_13552,N_13465);
and U13701 (N_13701,N_13450,N_13599);
nor U13702 (N_13702,N_13521,N_13535);
nand U13703 (N_13703,N_13582,N_13579);
and U13704 (N_13704,N_13463,N_13477);
and U13705 (N_13705,N_13429,N_13590);
and U13706 (N_13706,N_13511,N_13513);
nand U13707 (N_13707,N_13439,N_13584);
and U13708 (N_13708,N_13462,N_13487);
nor U13709 (N_13709,N_13440,N_13567);
and U13710 (N_13710,N_13435,N_13562);
or U13711 (N_13711,N_13505,N_13597);
and U13712 (N_13712,N_13555,N_13514);
or U13713 (N_13713,N_13402,N_13458);
nor U13714 (N_13714,N_13472,N_13541);
or U13715 (N_13715,N_13543,N_13403);
nand U13716 (N_13716,N_13444,N_13408);
and U13717 (N_13717,N_13447,N_13426);
nor U13718 (N_13718,N_13527,N_13584);
nand U13719 (N_13719,N_13444,N_13433);
or U13720 (N_13720,N_13558,N_13442);
or U13721 (N_13721,N_13415,N_13587);
and U13722 (N_13722,N_13502,N_13410);
and U13723 (N_13723,N_13589,N_13403);
or U13724 (N_13724,N_13527,N_13522);
nand U13725 (N_13725,N_13470,N_13537);
nand U13726 (N_13726,N_13510,N_13581);
nand U13727 (N_13727,N_13518,N_13470);
nor U13728 (N_13728,N_13508,N_13520);
nand U13729 (N_13729,N_13512,N_13460);
and U13730 (N_13730,N_13554,N_13567);
and U13731 (N_13731,N_13575,N_13593);
nand U13732 (N_13732,N_13575,N_13557);
nor U13733 (N_13733,N_13577,N_13420);
or U13734 (N_13734,N_13404,N_13508);
nand U13735 (N_13735,N_13582,N_13539);
nor U13736 (N_13736,N_13537,N_13569);
xnor U13737 (N_13737,N_13411,N_13534);
nand U13738 (N_13738,N_13581,N_13453);
nor U13739 (N_13739,N_13430,N_13529);
or U13740 (N_13740,N_13463,N_13456);
or U13741 (N_13741,N_13576,N_13559);
and U13742 (N_13742,N_13492,N_13547);
nor U13743 (N_13743,N_13509,N_13478);
or U13744 (N_13744,N_13496,N_13593);
xnor U13745 (N_13745,N_13585,N_13529);
nand U13746 (N_13746,N_13533,N_13514);
or U13747 (N_13747,N_13578,N_13477);
nor U13748 (N_13748,N_13400,N_13450);
or U13749 (N_13749,N_13586,N_13571);
nand U13750 (N_13750,N_13576,N_13484);
or U13751 (N_13751,N_13517,N_13595);
and U13752 (N_13752,N_13573,N_13500);
or U13753 (N_13753,N_13545,N_13462);
nor U13754 (N_13754,N_13564,N_13555);
nor U13755 (N_13755,N_13564,N_13546);
or U13756 (N_13756,N_13540,N_13464);
nand U13757 (N_13757,N_13551,N_13421);
nor U13758 (N_13758,N_13482,N_13522);
or U13759 (N_13759,N_13579,N_13424);
nand U13760 (N_13760,N_13534,N_13443);
nand U13761 (N_13761,N_13525,N_13417);
or U13762 (N_13762,N_13417,N_13512);
nor U13763 (N_13763,N_13591,N_13566);
and U13764 (N_13764,N_13526,N_13522);
nor U13765 (N_13765,N_13577,N_13513);
nand U13766 (N_13766,N_13474,N_13433);
nand U13767 (N_13767,N_13593,N_13598);
nor U13768 (N_13768,N_13486,N_13517);
nand U13769 (N_13769,N_13456,N_13419);
or U13770 (N_13770,N_13434,N_13460);
nor U13771 (N_13771,N_13588,N_13539);
nor U13772 (N_13772,N_13593,N_13408);
nor U13773 (N_13773,N_13438,N_13599);
nand U13774 (N_13774,N_13501,N_13591);
nor U13775 (N_13775,N_13461,N_13454);
nor U13776 (N_13776,N_13450,N_13493);
and U13777 (N_13777,N_13547,N_13474);
and U13778 (N_13778,N_13476,N_13521);
or U13779 (N_13779,N_13512,N_13449);
or U13780 (N_13780,N_13565,N_13442);
nand U13781 (N_13781,N_13599,N_13449);
and U13782 (N_13782,N_13534,N_13597);
and U13783 (N_13783,N_13556,N_13514);
nor U13784 (N_13784,N_13507,N_13570);
and U13785 (N_13785,N_13586,N_13558);
nand U13786 (N_13786,N_13500,N_13582);
and U13787 (N_13787,N_13472,N_13469);
nand U13788 (N_13788,N_13515,N_13533);
or U13789 (N_13789,N_13566,N_13454);
nand U13790 (N_13790,N_13514,N_13560);
or U13791 (N_13791,N_13413,N_13439);
or U13792 (N_13792,N_13593,N_13577);
nor U13793 (N_13793,N_13410,N_13426);
or U13794 (N_13794,N_13432,N_13449);
and U13795 (N_13795,N_13466,N_13441);
or U13796 (N_13796,N_13434,N_13534);
and U13797 (N_13797,N_13527,N_13438);
and U13798 (N_13798,N_13551,N_13554);
nor U13799 (N_13799,N_13403,N_13529);
and U13800 (N_13800,N_13630,N_13754);
and U13801 (N_13801,N_13794,N_13720);
and U13802 (N_13802,N_13738,N_13689);
and U13803 (N_13803,N_13706,N_13744);
or U13804 (N_13804,N_13679,N_13658);
nor U13805 (N_13805,N_13724,N_13626);
nor U13806 (N_13806,N_13713,N_13648);
and U13807 (N_13807,N_13790,N_13764);
or U13808 (N_13808,N_13780,N_13684);
and U13809 (N_13809,N_13692,N_13675);
nor U13810 (N_13810,N_13646,N_13717);
and U13811 (N_13811,N_13698,N_13791);
nor U13812 (N_13812,N_13796,N_13606);
or U13813 (N_13813,N_13633,N_13721);
nor U13814 (N_13814,N_13603,N_13678);
nand U13815 (N_13815,N_13743,N_13733);
and U13816 (N_13816,N_13642,N_13631);
nand U13817 (N_13817,N_13708,N_13704);
nand U13818 (N_13818,N_13641,N_13627);
nand U13819 (N_13819,N_13745,N_13690);
nand U13820 (N_13820,N_13783,N_13660);
nand U13821 (N_13821,N_13649,N_13644);
nand U13822 (N_13822,N_13673,N_13669);
nor U13823 (N_13823,N_13798,N_13670);
or U13824 (N_13824,N_13771,N_13760);
xnor U13825 (N_13825,N_13782,N_13766);
and U13826 (N_13826,N_13629,N_13664);
nand U13827 (N_13827,N_13740,N_13653);
nor U13828 (N_13828,N_13770,N_13750);
and U13829 (N_13829,N_13739,N_13773);
or U13830 (N_13830,N_13610,N_13614);
nor U13831 (N_13831,N_13752,N_13737);
or U13832 (N_13832,N_13608,N_13635);
and U13833 (N_13833,N_13699,N_13668);
and U13834 (N_13834,N_13657,N_13710);
nor U13835 (N_13835,N_13736,N_13615);
or U13836 (N_13836,N_13774,N_13718);
nor U13837 (N_13837,N_13655,N_13728);
or U13838 (N_13838,N_13703,N_13705);
and U13839 (N_13839,N_13767,N_13772);
nor U13840 (N_13840,N_13654,N_13793);
and U13841 (N_13841,N_13628,N_13676);
nor U13842 (N_13842,N_13776,N_13731);
or U13843 (N_13843,N_13778,N_13693);
nand U13844 (N_13844,N_13671,N_13709);
nand U13845 (N_13845,N_13691,N_13621);
and U13846 (N_13846,N_13726,N_13686);
and U13847 (N_13847,N_13645,N_13757);
or U13848 (N_13848,N_13638,N_13622);
nor U13849 (N_13849,N_13759,N_13623);
and U13850 (N_13850,N_13735,N_13702);
nor U13851 (N_13851,N_13751,N_13775);
or U13852 (N_13852,N_13650,N_13719);
nand U13853 (N_13853,N_13663,N_13761);
or U13854 (N_13854,N_13632,N_13612);
or U13855 (N_13855,N_13781,N_13749);
nor U13856 (N_13856,N_13707,N_13777);
nand U13857 (N_13857,N_13715,N_13651);
or U13858 (N_13858,N_13695,N_13662);
nor U13859 (N_13859,N_13787,N_13730);
and U13860 (N_13860,N_13665,N_13677);
and U13861 (N_13861,N_13674,N_13758);
or U13862 (N_13862,N_13661,N_13613);
and U13863 (N_13863,N_13755,N_13616);
and U13864 (N_13864,N_13711,N_13634);
nor U13865 (N_13865,N_13753,N_13799);
nor U13866 (N_13866,N_13748,N_13643);
and U13867 (N_13867,N_13768,N_13742);
nand U13868 (N_13868,N_13788,N_13732);
and U13869 (N_13869,N_13697,N_13672);
nand U13870 (N_13870,N_13694,N_13734);
nor U13871 (N_13871,N_13619,N_13639);
or U13872 (N_13872,N_13779,N_13602);
nand U13873 (N_13873,N_13700,N_13747);
nor U13874 (N_13874,N_13604,N_13652);
nor U13875 (N_13875,N_13636,N_13601);
nor U13876 (N_13876,N_13683,N_13656);
xor U13877 (N_13877,N_13605,N_13785);
and U13878 (N_13878,N_13792,N_13722);
nand U13879 (N_13879,N_13769,N_13620);
and U13880 (N_13880,N_13729,N_13609);
nand U13881 (N_13881,N_13666,N_13765);
nand U13882 (N_13882,N_13723,N_13687);
or U13883 (N_13883,N_13607,N_13637);
nand U13884 (N_13884,N_13725,N_13667);
and U13885 (N_13885,N_13688,N_13789);
nand U13886 (N_13886,N_13640,N_13659);
nor U13887 (N_13887,N_13600,N_13680);
and U13888 (N_13888,N_13625,N_13756);
nor U13889 (N_13889,N_13795,N_13746);
nor U13890 (N_13890,N_13624,N_13762);
and U13891 (N_13891,N_13617,N_13618);
and U13892 (N_13892,N_13727,N_13647);
or U13893 (N_13893,N_13712,N_13797);
or U13894 (N_13894,N_13714,N_13611);
nand U13895 (N_13895,N_13696,N_13682);
nand U13896 (N_13896,N_13741,N_13784);
nor U13897 (N_13897,N_13786,N_13685);
and U13898 (N_13898,N_13716,N_13701);
xnor U13899 (N_13899,N_13763,N_13681);
xnor U13900 (N_13900,N_13761,N_13628);
nand U13901 (N_13901,N_13740,N_13731);
or U13902 (N_13902,N_13664,N_13796);
and U13903 (N_13903,N_13797,N_13688);
xor U13904 (N_13904,N_13648,N_13673);
nand U13905 (N_13905,N_13713,N_13680);
nor U13906 (N_13906,N_13775,N_13720);
nand U13907 (N_13907,N_13688,N_13676);
and U13908 (N_13908,N_13602,N_13718);
nand U13909 (N_13909,N_13610,N_13645);
or U13910 (N_13910,N_13672,N_13742);
nor U13911 (N_13911,N_13731,N_13739);
and U13912 (N_13912,N_13794,N_13702);
nor U13913 (N_13913,N_13684,N_13781);
nor U13914 (N_13914,N_13638,N_13708);
and U13915 (N_13915,N_13605,N_13733);
nor U13916 (N_13916,N_13763,N_13632);
nand U13917 (N_13917,N_13688,N_13744);
and U13918 (N_13918,N_13665,N_13616);
nor U13919 (N_13919,N_13673,N_13742);
nor U13920 (N_13920,N_13632,N_13775);
nor U13921 (N_13921,N_13672,N_13765);
and U13922 (N_13922,N_13726,N_13775);
or U13923 (N_13923,N_13659,N_13672);
nand U13924 (N_13924,N_13742,N_13654);
nor U13925 (N_13925,N_13617,N_13766);
or U13926 (N_13926,N_13789,N_13797);
or U13927 (N_13927,N_13785,N_13625);
nor U13928 (N_13928,N_13772,N_13618);
nor U13929 (N_13929,N_13600,N_13764);
nor U13930 (N_13930,N_13694,N_13692);
or U13931 (N_13931,N_13607,N_13765);
nor U13932 (N_13932,N_13600,N_13687);
and U13933 (N_13933,N_13617,N_13624);
and U13934 (N_13934,N_13746,N_13634);
nand U13935 (N_13935,N_13795,N_13741);
nand U13936 (N_13936,N_13745,N_13643);
and U13937 (N_13937,N_13640,N_13682);
or U13938 (N_13938,N_13786,N_13684);
and U13939 (N_13939,N_13612,N_13718);
nor U13940 (N_13940,N_13632,N_13625);
or U13941 (N_13941,N_13714,N_13647);
and U13942 (N_13942,N_13637,N_13653);
and U13943 (N_13943,N_13766,N_13729);
or U13944 (N_13944,N_13758,N_13618);
or U13945 (N_13945,N_13792,N_13601);
or U13946 (N_13946,N_13626,N_13600);
nor U13947 (N_13947,N_13706,N_13747);
nand U13948 (N_13948,N_13637,N_13707);
or U13949 (N_13949,N_13637,N_13617);
nor U13950 (N_13950,N_13736,N_13710);
nand U13951 (N_13951,N_13783,N_13646);
nand U13952 (N_13952,N_13656,N_13746);
nor U13953 (N_13953,N_13776,N_13618);
nand U13954 (N_13954,N_13662,N_13760);
and U13955 (N_13955,N_13642,N_13750);
and U13956 (N_13956,N_13782,N_13601);
nor U13957 (N_13957,N_13754,N_13710);
or U13958 (N_13958,N_13652,N_13733);
nor U13959 (N_13959,N_13701,N_13785);
nor U13960 (N_13960,N_13765,N_13606);
and U13961 (N_13961,N_13783,N_13643);
nor U13962 (N_13962,N_13762,N_13654);
and U13963 (N_13963,N_13732,N_13626);
or U13964 (N_13964,N_13724,N_13762);
and U13965 (N_13965,N_13671,N_13768);
nand U13966 (N_13966,N_13706,N_13738);
and U13967 (N_13967,N_13756,N_13745);
and U13968 (N_13968,N_13671,N_13677);
or U13969 (N_13969,N_13749,N_13716);
nand U13970 (N_13970,N_13738,N_13758);
nand U13971 (N_13971,N_13675,N_13750);
nor U13972 (N_13972,N_13623,N_13765);
or U13973 (N_13973,N_13631,N_13637);
or U13974 (N_13974,N_13631,N_13665);
nand U13975 (N_13975,N_13721,N_13689);
nand U13976 (N_13976,N_13691,N_13755);
nor U13977 (N_13977,N_13723,N_13728);
or U13978 (N_13978,N_13619,N_13673);
or U13979 (N_13979,N_13770,N_13607);
nand U13980 (N_13980,N_13634,N_13704);
or U13981 (N_13981,N_13721,N_13716);
and U13982 (N_13982,N_13634,N_13778);
nor U13983 (N_13983,N_13662,N_13755);
and U13984 (N_13984,N_13659,N_13752);
or U13985 (N_13985,N_13677,N_13651);
and U13986 (N_13986,N_13692,N_13616);
nand U13987 (N_13987,N_13719,N_13611);
nand U13988 (N_13988,N_13676,N_13755);
nand U13989 (N_13989,N_13756,N_13707);
and U13990 (N_13990,N_13705,N_13666);
nor U13991 (N_13991,N_13701,N_13768);
nand U13992 (N_13992,N_13714,N_13636);
or U13993 (N_13993,N_13685,N_13625);
nor U13994 (N_13994,N_13699,N_13771);
nor U13995 (N_13995,N_13614,N_13696);
and U13996 (N_13996,N_13673,N_13765);
nor U13997 (N_13997,N_13766,N_13770);
and U13998 (N_13998,N_13658,N_13677);
nor U13999 (N_13999,N_13708,N_13794);
nor U14000 (N_14000,N_13973,N_13908);
and U14001 (N_14001,N_13896,N_13910);
or U14002 (N_14002,N_13866,N_13808);
and U14003 (N_14003,N_13846,N_13828);
nor U14004 (N_14004,N_13841,N_13969);
and U14005 (N_14005,N_13890,N_13899);
and U14006 (N_14006,N_13817,N_13833);
or U14007 (N_14007,N_13945,N_13867);
nand U14008 (N_14008,N_13949,N_13814);
and U14009 (N_14009,N_13864,N_13898);
nor U14010 (N_14010,N_13951,N_13960);
nand U14011 (N_14011,N_13830,N_13819);
nor U14012 (N_14012,N_13874,N_13940);
or U14013 (N_14013,N_13850,N_13991);
nand U14014 (N_14014,N_13880,N_13829);
nand U14015 (N_14015,N_13897,N_13947);
and U14016 (N_14016,N_13931,N_13835);
and U14017 (N_14017,N_13832,N_13886);
nand U14018 (N_14018,N_13987,N_13994);
or U14019 (N_14019,N_13831,N_13943);
and U14020 (N_14020,N_13974,N_13803);
nand U14021 (N_14021,N_13923,N_13844);
nand U14022 (N_14022,N_13920,N_13919);
or U14023 (N_14023,N_13975,N_13815);
and U14024 (N_14024,N_13964,N_13888);
nand U14025 (N_14025,N_13818,N_13934);
nor U14026 (N_14026,N_13900,N_13954);
nand U14027 (N_14027,N_13925,N_13996);
and U14028 (N_14028,N_13861,N_13858);
nor U14029 (N_14029,N_13849,N_13993);
nand U14030 (N_14030,N_13873,N_13988);
or U14031 (N_14031,N_13860,N_13807);
nor U14032 (N_14032,N_13990,N_13872);
or U14033 (N_14033,N_13962,N_13812);
nand U14034 (N_14034,N_13979,N_13946);
nand U14035 (N_14035,N_13827,N_13976);
and U14036 (N_14036,N_13909,N_13932);
or U14037 (N_14037,N_13985,N_13826);
nand U14038 (N_14038,N_13865,N_13917);
and U14039 (N_14039,N_13902,N_13970);
xnor U14040 (N_14040,N_13914,N_13971);
nor U14041 (N_14041,N_13884,N_13859);
and U14042 (N_14042,N_13984,N_13998);
nand U14043 (N_14043,N_13903,N_13845);
and U14044 (N_14044,N_13839,N_13941);
and U14045 (N_14045,N_13836,N_13922);
nor U14046 (N_14046,N_13825,N_13916);
nor U14047 (N_14047,N_13809,N_13882);
or U14048 (N_14048,N_13904,N_13977);
and U14049 (N_14049,N_13915,N_13823);
and U14050 (N_14050,N_13901,N_13857);
and U14051 (N_14051,N_13838,N_13967);
and U14052 (N_14052,N_13959,N_13927);
nand U14053 (N_14053,N_13997,N_13950);
or U14054 (N_14054,N_13869,N_13847);
or U14055 (N_14055,N_13989,N_13982);
nor U14056 (N_14056,N_13834,N_13905);
or U14057 (N_14057,N_13895,N_13871);
and U14058 (N_14058,N_13937,N_13820);
and U14059 (N_14059,N_13889,N_13840);
nand U14060 (N_14060,N_13942,N_13918);
nor U14061 (N_14061,N_13986,N_13939);
nor U14062 (N_14062,N_13891,N_13966);
or U14063 (N_14063,N_13856,N_13936);
nand U14064 (N_14064,N_13805,N_13876);
nand U14065 (N_14065,N_13938,N_13930);
and U14066 (N_14066,N_13928,N_13952);
or U14067 (N_14067,N_13883,N_13854);
or U14068 (N_14068,N_13862,N_13924);
and U14069 (N_14069,N_13953,N_13981);
nand U14070 (N_14070,N_13955,N_13911);
or U14071 (N_14071,N_13806,N_13821);
nand U14072 (N_14072,N_13853,N_13885);
xor U14073 (N_14073,N_13913,N_13811);
and U14074 (N_14074,N_13824,N_13965);
or U14075 (N_14075,N_13929,N_13968);
or U14076 (N_14076,N_13848,N_13837);
nand U14077 (N_14077,N_13992,N_13978);
or U14078 (N_14078,N_13802,N_13958);
nor U14079 (N_14079,N_13810,N_13906);
or U14080 (N_14080,N_13843,N_13842);
nand U14081 (N_14081,N_13881,N_13868);
and U14082 (N_14082,N_13963,N_13921);
nand U14083 (N_14083,N_13870,N_13801);
and U14084 (N_14084,N_13813,N_13855);
nand U14085 (N_14085,N_13851,N_13875);
and U14086 (N_14086,N_13956,N_13863);
nand U14087 (N_14087,N_13877,N_13816);
nand U14088 (N_14088,N_13957,N_13852);
nand U14089 (N_14089,N_13961,N_13926);
and U14090 (N_14090,N_13894,N_13887);
nor U14091 (N_14091,N_13948,N_13804);
nand U14092 (N_14092,N_13944,N_13892);
or U14093 (N_14093,N_13935,N_13995);
nor U14094 (N_14094,N_13878,N_13933);
and U14095 (N_14095,N_13800,N_13893);
nor U14096 (N_14096,N_13912,N_13972);
or U14097 (N_14097,N_13999,N_13983);
and U14098 (N_14098,N_13980,N_13879);
and U14099 (N_14099,N_13907,N_13822);
nand U14100 (N_14100,N_13992,N_13944);
or U14101 (N_14101,N_13811,N_13982);
and U14102 (N_14102,N_13918,N_13838);
nand U14103 (N_14103,N_13836,N_13841);
nand U14104 (N_14104,N_13855,N_13996);
nand U14105 (N_14105,N_13934,N_13803);
nand U14106 (N_14106,N_13945,N_13863);
nand U14107 (N_14107,N_13933,N_13864);
or U14108 (N_14108,N_13853,N_13989);
nor U14109 (N_14109,N_13915,N_13930);
or U14110 (N_14110,N_13906,N_13995);
nand U14111 (N_14111,N_13901,N_13974);
or U14112 (N_14112,N_13940,N_13860);
nand U14113 (N_14113,N_13948,N_13906);
nor U14114 (N_14114,N_13855,N_13960);
nand U14115 (N_14115,N_13956,N_13996);
or U14116 (N_14116,N_13825,N_13864);
nand U14117 (N_14117,N_13979,N_13846);
or U14118 (N_14118,N_13926,N_13936);
and U14119 (N_14119,N_13923,N_13809);
or U14120 (N_14120,N_13869,N_13958);
or U14121 (N_14121,N_13980,N_13844);
and U14122 (N_14122,N_13936,N_13970);
or U14123 (N_14123,N_13937,N_13896);
and U14124 (N_14124,N_13871,N_13883);
nor U14125 (N_14125,N_13839,N_13831);
nor U14126 (N_14126,N_13900,N_13890);
nor U14127 (N_14127,N_13852,N_13869);
and U14128 (N_14128,N_13875,N_13970);
or U14129 (N_14129,N_13992,N_13821);
nor U14130 (N_14130,N_13977,N_13812);
nor U14131 (N_14131,N_13930,N_13977);
and U14132 (N_14132,N_13962,N_13836);
nand U14133 (N_14133,N_13817,N_13905);
or U14134 (N_14134,N_13920,N_13928);
nor U14135 (N_14135,N_13959,N_13965);
or U14136 (N_14136,N_13834,N_13908);
nand U14137 (N_14137,N_13810,N_13916);
nand U14138 (N_14138,N_13827,N_13811);
xnor U14139 (N_14139,N_13980,N_13908);
or U14140 (N_14140,N_13905,N_13856);
nand U14141 (N_14141,N_13869,N_13863);
nor U14142 (N_14142,N_13872,N_13912);
nor U14143 (N_14143,N_13914,N_13807);
and U14144 (N_14144,N_13836,N_13812);
nor U14145 (N_14145,N_13865,N_13962);
nand U14146 (N_14146,N_13867,N_13986);
and U14147 (N_14147,N_13883,N_13801);
and U14148 (N_14148,N_13885,N_13979);
nor U14149 (N_14149,N_13999,N_13874);
and U14150 (N_14150,N_13879,N_13834);
or U14151 (N_14151,N_13871,N_13878);
or U14152 (N_14152,N_13978,N_13829);
nand U14153 (N_14153,N_13969,N_13886);
nor U14154 (N_14154,N_13833,N_13941);
nand U14155 (N_14155,N_13896,N_13839);
and U14156 (N_14156,N_13980,N_13904);
nor U14157 (N_14157,N_13845,N_13990);
nor U14158 (N_14158,N_13934,N_13902);
nand U14159 (N_14159,N_13966,N_13945);
nand U14160 (N_14160,N_13893,N_13806);
nand U14161 (N_14161,N_13807,N_13851);
nor U14162 (N_14162,N_13990,N_13896);
and U14163 (N_14163,N_13939,N_13948);
nand U14164 (N_14164,N_13899,N_13828);
and U14165 (N_14165,N_13830,N_13958);
or U14166 (N_14166,N_13800,N_13910);
nand U14167 (N_14167,N_13911,N_13824);
and U14168 (N_14168,N_13831,N_13966);
or U14169 (N_14169,N_13957,N_13846);
and U14170 (N_14170,N_13985,N_13959);
nor U14171 (N_14171,N_13907,N_13801);
and U14172 (N_14172,N_13975,N_13936);
nor U14173 (N_14173,N_13862,N_13868);
and U14174 (N_14174,N_13925,N_13898);
nand U14175 (N_14175,N_13903,N_13818);
nand U14176 (N_14176,N_13958,N_13981);
and U14177 (N_14177,N_13966,N_13886);
nand U14178 (N_14178,N_13906,N_13808);
nor U14179 (N_14179,N_13904,N_13871);
nand U14180 (N_14180,N_13924,N_13919);
nand U14181 (N_14181,N_13870,N_13888);
or U14182 (N_14182,N_13832,N_13911);
nor U14183 (N_14183,N_13808,N_13975);
or U14184 (N_14184,N_13824,N_13957);
nand U14185 (N_14185,N_13858,N_13931);
or U14186 (N_14186,N_13937,N_13823);
or U14187 (N_14187,N_13903,N_13978);
nor U14188 (N_14188,N_13861,N_13945);
and U14189 (N_14189,N_13965,N_13932);
and U14190 (N_14190,N_13870,N_13926);
nand U14191 (N_14191,N_13934,N_13868);
and U14192 (N_14192,N_13838,N_13907);
and U14193 (N_14193,N_13870,N_13921);
nor U14194 (N_14194,N_13826,N_13825);
nand U14195 (N_14195,N_13845,N_13887);
xor U14196 (N_14196,N_13931,N_13897);
or U14197 (N_14197,N_13871,N_13942);
and U14198 (N_14198,N_13802,N_13881);
and U14199 (N_14199,N_13921,N_13950);
or U14200 (N_14200,N_14081,N_14132);
or U14201 (N_14201,N_14092,N_14172);
or U14202 (N_14202,N_14115,N_14018);
nor U14203 (N_14203,N_14168,N_14113);
nand U14204 (N_14204,N_14090,N_14089);
or U14205 (N_14205,N_14065,N_14151);
nor U14206 (N_14206,N_14122,N_14180);
or U14207 (N_14207,N_14183,N_14163);
nand U14208 (N_14208,N_14068,N_14042);
nor U14209 (N_14209,N_14140,N_14061);
nor U14210 (N_14210,N_14072,N_14054);
or U14211 (N_14211,N_14159,N_14035);
or U14212 (N_14212,N_14044,N_14195);
nor U14213 (N_14213,N_14171,N_14004);
nor U14214 (N_14214,N_14015,N_14155);
nand U14215 (N_14215,N_14062,N_14067);
nor U14216 (N_14216,N_14166,N_14129);
or U14217 (N_14217,N_14037,N_14100);
and U14218 (N_14218,N_14136,N_14007);
and U14219 (N_14219,N_14077,N_14199);
or U14220 (N_14220,N_14008,N_14094);
and U14221 (N_14221,N_14116,N_14064);
nand U14222 (N_14222,N_14108,N_14154);
or U14223 (N_14223,N_14075,N_14079);
and U14224 (N_14224,N_14181,N_14028);
nor U14225 (N_14225,N_14139,N_14016);
and U14226 (N_14226,N_14146,N_14142);
or U14227 (N_14227,N_14121,N_14013);
or U14228 (N_14228,N_14191,N_14022);
nand U14229 (N_14229,N_14179,N_14125);
nor U14230 (N_14230,N_14073,N_14170);
or U14231 (N_14231,N_14109,N_14058);
and U14232 (N_14232,N_14034,N_14148);
or U14233 (N_14233,N_14112,N_14097);
and U14234 (N_14234,N_14133,N_14071);
or U14235 (N_14235,N_14128,N_14192);
nand U14236 (N_14236,N_14196,N_14167);
nor U14237 (N_14237,N_14083,N_14193);
and U14238 (N_14238,N_14052,N_14164);
nor U14239 (N_14239,N_14162,N_14012);
and U14240 (N_14240,N_14020,N_14105);
nor U14241 (N_14241,N_14010,N_14006);
or U14242 (N_14242,N_14025,N_14106);
and U14243 (N_14243,N_14048,N_14176);
and U14244 (N_14244,N_14069,N_14045);
or U14245 (N_14245,N_14150,N_14049);
nor U14246 (N_14246,N_14003,N_14189);
nand U14247 (N_14247,N_14085,N_14047);
nor U14248 (N_14248,N_14041,N_14091);
nor U14249 (N_14249,N_14103,N_14111);
nor U14250 (N_14250,N_14110,N_14057);
and U14251 (N_14251,N_14190,N_14169);
nand U14252 (N_14252,N_14144,N_14023);
nor U14253 (N_14253,N_14117,N_14138);
nand U14254 (N_14254,N_14114,N_14063);
nand U14255 (N_14255,N_14024,N_14178);
nor U14256 (N_14256,N_14039,N_14102);
or U14257 (N_14257,N_14011,N_14000);
or U14258 (N_14258,N_14093,N_14060);
nand U14259 (N_14259,N_14107,N_14005);
nand U14260 (N_14260,N_14141,N_14076);
or U14261 (N_14261,N_14036,N_14157);
or U14262 (N_14262,N_14149,N_14126);
nand U14263 (N_14263,N_14017,N_14032);
and U14264 (N_14264,N_14059,N_14029);
or U14265 (N_14265,N_14118,N_14194);
or U14266 (N_14266,N_14143,N_14070);
nor U14267 (N_14267,N_14087,N_14074);
or U14268 (N_14268,N_14158,N_14177);
nand U14269 (N_14269,N_14147,N_14182);
and U14270 (N_14270,N_14009,N_14027);
nor U14271 (N_14271,N_14099,N_14127);
and U14272 (N_14272,N_14038,N_14124);
and U14273 (N_14273,N_14156,N_14197);
and U14274 (N_14274,N_14056,N_14186);
nand U14275 (N_14275,N_14165,N_14019);
nand U14276 (N_14276,N_14001,N_14184);
xor U14277 (N_14277,N_14066,N_14098);
nor U14278 (N_14278,N_14040,N_14123);
and U14279 (N_14279,N_14078,N_14104);
nor U14280 (N_14280,N_14021,N_14096);
or U14281 (N_14281,N_14030,N_14135);
or U14282 (N_14282,N_14033,N_14101);
nand U14283 (N_14283,N_14046,N_14145);
nor U14284 (N_14284,N_14137,N_14119);
nor U14285 (N_14285,N_14188,N_14051);
or U14286 (N_14286,N_14031,N_14088);
and U14287 (N_14287,N_14084,N_14086);
or U14288 (N_14288,N_14134,N_14161);
nor U14289 (N_14289,N_14174,N_14055);
nor U14290 (N_14290,N_14187,N_14131);
and U14291 (N_14291,N_14130,N_14152);
or U14292 (N_14292,N_14120,N_14026);
and U14293 (N_14293,N_14002,N_14175);
and U14294 (N_14294,N_14185,N_14095);
and U14295 (N_14295,N_14082,N_14014);
or U14296 (N_14296,N_14043,N_14160);
and U14297 (N_14297,N_14080,N_14053);
nand U14298 (N_14298,N_14050,N_14173);
xor U14299 (N_14299,N_14153,N_14198);
and U14300 (N_14300,N_14168,N_14094);
or U14301 (N_14301,N_14105,N_14046);
nor U14302 (N_14302,N_14075,N_14190);
or U14303 (N_14303,N_14160,N_14009);
and U14304 (N_14304,N_14135,N_14178);
or U14305 (N_14305,N_14068,N_14133);
nand U14306 (N_14306,N_14155,N_14020);
nand U14307 (N_14307,N_14150,N_14022);
and U14308 (N_14308,N_14192,N_14075);
and U14309 (N_14309,N_14034,N_14054);
nor U14310 (N_14310,N_14131,N_14184);
nand U14311 (N_14311,N_14146,N_14190);
or U14312 (N_14312,N_14053,N_14031);
and U14313 (N_14313,N_14128,N_14017);
and U14314 (N_14314,N_14186,N_14007);
nor U14315 (N_14315,N_14090,N_14037);
and U14316 (N_14316,N_14141,N_14027);
and U14317 (N_14317,N_14146,N_14033);
and U14318 (N_14318,N_14062,N_14019);
nand U14319 (N_14319,N_14124,N_14048);
and U14320 (N_14320,N_14035,N_14140);
nor U14321 (N_14321,N_14146,N_14005);
and U14322 (N_14322,N_14065,N_14035);
and U14323 (N_14323,N_14158,N_14155);
nor U14324 (N_14324,N_14117,N_14034);
and U14325 (N_14325,N_14055,N_14111);
nor U14326 (N_14326,N_14184,N_14141);
or U14327 (N_14327,N_14030,N_14060);
nor U14328 (N_14328,N_14071,N_14011);
or U14329 (N_14329,N_14061,N_14137);
and U14330 (N_14330,N_14083,N_14174);
or U14331 (N_14331,N_14184,N_14178);
and U14332 (N_14332,N_14168,N_14071);
nor U14333 (N_14333,N_14027,N_14104);
nand U14334 (N_14334,N_14014,N_14013);
and U14335 (N_14335,N_14178,N_14112);
nor U14336 (N_14336,N_14045,N_14004);
and U14337 (N_14337,N_14003,N_14009);
nor U14338 (N_14338,N_14095,N_14195);
or U14339 (N_14339,N_14051,N_14122);
or U14340 (N_14340,N_14053,N_14113);
nor U14341 (N_14341,N_14088,N_14125);
and U14342 (N_14342,N_14061,N_14003);
and U14343 (N_14343,N_14042,N_14082);
nand U14344 (N_14344,N_14154,N_14042);
or U14345 (N_14345,N_14128,N_14096);
xor U14346 (N_14346,N_14087,N_14137);
or U14347 (N_14347,N_14082,N_14064);
xor U14348 (N_14348,N_14165,N_14048);
nand U14349 (N_14349,N_14126,N_14145);
and U14350 (N_14350,N_14050,N_14057);
and U14351 (N_14351,N_14067,N_14103);
nand U14352 (N_14352,N_14071,N_14081);
and U14353 (N_14353,N_14073,N_14157);
and U14354 (N_14354,N_14086,N_14194);
or U14355 (N_14355,N_14069,N_14017);
nand U14356 (N_14356,N_14166,N_14133);
or U14357 (N_14357,N_14025,N_14153);
and U14358 (N_14358,N_14103,N_14037);
or U14359 (N_14359,N_14022,N_14024);
or U14360 (N_14360,N_14080,N_14019);
nand U14361 (N_14361,N_14087,N_14009);
and U14362 (N_14362,N_14084,N_14107);
nor U14363 (N_14363,N_14137,N_14100);
nand U14364 (N_14364,N_14129,N_14135);
nand U14365 (N_14365,N_14086,N_14081);
and U14366 (N_14366,N_14134,N_14063);
nor U14367 (N_14367,N_14036,N_14123);
or U14368 (N_14368,N_14171,N_14153);
and U14369 (N_14369,N_14097,N_14150);
nand U14370 (N_14370,N_14040,N_14073);
nand U14371 (N_14371,N_14044,N_14121);
nor U14372 (N_14372,N_14059,N_14122);
or U14373 (N_14373,N_14090,N_14028);
nor U14374 (N_14374,N_14078,N_14060);
nor U14375 (N_14375,N_14112,N_14040);
nand U14376 (N_14376,N_14049,N_14168);
and U14377 (N_14377,N_14160,N_14161);
or U14378 (N_14378,N_14037,N_14013);
or U14379 (N_14379,N_14019,N_14000);
or U14380 (N_14380,N_14073,N_14033);
nand U14381 (N_14381,N_14085,N_14199);
nand U14382 (N_14382,N_14021,N_14137);
nand U14383 (N_14383,N_14168,N_14010);
or U14384 (N_14384,N_14115,N_14019);
and U14385 (N_14385,N_14138,N_14067);
or U14386 (N_14386,N_14001,N_14150);
and U14387 (N_14387,N_14013,N_14106);
or U14388 (N_14388,N_14068,N_14071);
or U14389 (N_14389,N_14046,N_14120);
and U14390 (N_14390,N_14053,N_14129);
nor U14391 (N_14391,N_14175,N_14139);
nand U14392 (N_14392,N_14014,N_14027);
or U14393 (N_14393,N_14116,N_14045);
nor U14394 (N_14394,N_14110,N_14003);
nor U14395 (N_14395,N_14176,N_14159);
and U14396 (N_14396,N_14162,N_14091);
nor U14397 (N_14397,N_14015,N_14112);
xnor U14398 (N_14398,N_14181,N_14163);
or U14399 (N_14399,N_14128,N_14027);
and U14400 (N_14400,N_14250,N_14381);
and U14401 (N_14401,N_14341,N_14357);
or U14402 (N_14402,N_14294,N_14355);
nor U14403 (N_14403,N_14227,N_14249);
nor U14404 (N_14404,N_14210,N_14332);
nand U14405 (N_14405,N_14329,N_14350);
and U14406 (N_14406,N_14277,N_14390);
and U14407 (N_14407,N_14279,N_14239);
or U14408 (N_14408,N_14334,N_14262);
nand U14409 (N_14409,N_14289,N_14288);
and U14410 (N_14410,N_14206,N_14300);
and U14411 (N_14411,N_14205,N_14395);
and U14412 (N_14412,N_14291,N_14325);
and U14413 (N_14413,N_14282,N_14237);
nand U14414 (N_14414,N_14240,N_14385);
nor U14415 (N_14415,N_14342,N_14321);
and U14416 (N_14416,N_14323,N_14312);
nand U14417 (N_14417,N_14219,N_14292);
nor U14418 (N_14418,N_14322,N_14269);
and U14419 (N_14419,N_14304,N_14271);
nor U14420 (N_14420,N_14351,N_14225);
nor U14421 (N_14421,N_14293,N_14232);
or U14422 (N_14422,N_14251,N_14336);
and U14423 (N_14423,N_14318,N_14333);
nand U14424 (N_14424,N_14203,N_14297);
nand U14425 (N_14425,N_14340,N_14295);
and U14426 (N_14426,N_14364,N_14223);
or U14427 (N_14427,N_14316,N_14306);
nor U14428 (N_14428,N_14246,N_14383);
nand U14429 (N_14429,N_14260,N_14243);
and U14430 (N_14430,N_14362,N_14359);
nor U14431 (N_14431,N_14274,N_14299);
nand U14432 (N_14432,N_14238,N_14356);
nand U14433 (N_14433,N_14265,N_14367);
nand U14434 (N_14434,N_14214,N_14200);
and U14435 (N_14435,N_14266,N_14216);
nand U14436 (N_14436,N_14270,N_14392);
nor U14437 (N_14437,N_14320,N_14261);
nor U14438 (N_14438,N_14388,N_14202);
and U14439 (N_14439,N_14382,N_14389);
or U14440 (N_14440,N_14324,N_14377);
or U14441 (N_14441,N_14308,N_14222);
nand U14442 (N_14442,N_14399,N_14303);
nand U14443 (N_14443,N_14281,N_14328);
and U14444 (N_14444,N_14365,N_14346);
nor U14445 (N_14445,N_14343,N_14327);
nor U14446 (N_14446,N_14201,N_14230);
nor U14447 (N_14447,N_14345,N_14369);
or U14448 (N_14448,N_14309,N_14301);
and U14449 (N_14449,N_14317,N_14287);
nor U14450 (N_14450,N_14344,N_14307);
or U14451 (N_14451,N_14373,N_14302);
or U14452 (N_14452,N_14268,N_14386);
nor U14453 (N_14453,N_14387,N_14349);
or U14454 (N_14454,N_14339,N_14348);
and U14455 (N_14455,N_14236,N_14290);
or U14456 (N_14456,N_14263,N_14253);
nor U14457 (N_14457,N_14361,N_14378);
or U14458 (N_14458,N_14217,N_14244);
nand U14459 (N_14459,N_14296,N_14226);
nor U14460 (N_14460,N_14257,N_14352);
nand U14461 (N_14461,N_14229,N_14248);
nand U14462 (N_14462,N_14273,N_14314);
nor U14463 (N_14463,N_14371,N_14326);
and U14464 (N_14464,N_14212,N_14285);
nor U14465 (N_14465,N_14204,N_14234);
nand U14466 (N_14466,N_14313,N_14363);
nor U14467 (N_14467,N_14331,N_14376);
and U14468 (N_14468,N_14375,N_14242);
and U14469 (N_14469,N_14353,N_14264);
nand U14470 (N_14470,N_14209,N_14393);
or U14471 (N_14471,N_14319,N_14255);
nand U14472 (N_14472,N_14228,N_14384);
nor U14473 (N_14473,N_14280,N_14207);
nand U14474 (N_14474,N_14254,N_14391);
nand U14475 (N_14475,N_14380,N_14258);
or U14476 (N_14476,N_14221,N_14394);
or U14477 (N_14477,N_14337,N_14218);
nand U14478 (N_14478,N_14347,N_14211);
or U14479 (N_14479,N_14259,N_14220);
or U14480 (N_14480,N_14275,N_14284);
nor U14481 (N_14481,N_14366,N_14241);
nand U14482 (N_14482,N_14272,N_14311);
nand U14483 (N_14483,N_14245,N_14379);
nand U14484 (N_14484,N_14397,N_14330);
and U14485 (N_14485,N_14335,N_14286);
or U14486 (N_14486,N_14315,N_14215);
nor U14487 (N_14487,N_14338,N_14235);
nand U14488 (N_14488,N_14252,N_14267);
or U14489 (N_14489,N_14276,N_14256);
nand U14490 (N_14490,N_14368,N_14278);
nand U14491 (N_14491,N_14310,N_14354);
and U14492 (N_14492,N_14374,N_14398);
and U14493 (N_14493,N_14360,N_14305);
or U14494 (N_14494,N_14247,N_14358);
nand U14495 (N_14495,N_14233,N_14396);
nor U14496 (N_14496,N_14298,N_14370);
nor U14497 (N_14497,N_14208,N_14213);
nand U14498 (N_14498,N_14283,N_14231);
nand U14499 (N_14499,N_14224,N_14372);
and U14500 (N_14500,N_14355,N_14266);
and U14501 (N_14501,N_14250,N_14391);
nor U14502 (N_14502,N_14269,N_14303);
nand U14503 (N_14503,N_14229,N_14255);
and U14504 (N_14504,N_14396,N_14241);
nand U14505 (N_14505,N_14293,N_14309);
and U14506 (N_14506,N_14207,N_14319);
nand U14507 (N_14507,N_14306,N_14379);
or U14508 (N_14508,N_14362,N_14296);
or U14509 (N_14509,N_14368,N_14284);
and U14510 (N_14510,N_14210,N_14289);
nor U14511 (N_14511,N_14287,N_14369);
and U14512 (N_14512,N_14304,N_14248);
or U14513 (N_14513,N_14265,N_14321);
nand U14514 (N_14514,N_14321,N_14221);
or U14515 (N_14515,N_14374,N_14229);
or U14516 (N_14516,N_14330,N_14285);
nand U14517 (N_14517,N_14234,N_14311);
xor U14518 (N_14518,N_14232,N_14388);
xnor U14519 (N_14519,N_14303,N_14256);
and U14520 (N_14520,N_14226,N_14398);
and U14521 (N_14521,N_14216,N_14259);
nand U14522 (N_14522,N_14202,N_14394);
and U14523 (N_14523,N_14310,N_14341);
and U14524 (N_14524,N_14314,N_14303);
nor U14525 (N_14525,N_14379,N_14226);
nor U14526 (N_14526,N_14260,N_14270);
nand U14527 (N_14527,N_14247,N_14369);
and U14528 (N_14528,N_14302,N_14389);
nor U14529 (N_14529,N_14257,N_14346);
or U14530 (N_14530,N_14210,N_14278);
nor U14531 (N_14531,N_14323,N_14340);
or U14532 (N_14532,N_14333,N_14382);
or U14533 (N_14533,N_14384,N_14351);
or U14534 (N_14534,N_14389,N_14249);
nor U14535 (N_14535,N_14288,N_14319);
nor U14536 (N_14536,N_14301,N_14331);
nor U14537 (N_14537,N_14315,N_14304);
nor U14538 (N_14538,N_14246,N_14347);
and U14539 (N_14539,N_14228,N_14258);
nand U14540 (N_14540,N_14335,N_14278);
and U14541 (N_14541,N_14216,N_14269);
nand U14542 (N_14542,N_14336,N_14271);
nor U14543 (N_14543,N_14386,N_14324);
nor U14544 (N_14544,N_14213,N_14212);
or U14545 (N_14545,N_14375,N_14298);
and U14546 (N_14546,N_14248,N_14264);
nor U14547 (N_14547,N_14335,N_14288);
nor U14548 (N_14548,N_14226,N_14305);
and U14549 (N_14549,N_14327,N_14240);
and U14550 (N_14550,N_14340,N_14348);
and U14551 (N_14551,N_14337,N_14342);
nor U14552 (N_14552,N_14269,N_14234);
nand U14553 (N_14553,N_14319,N_14311);
nor U14554 (N_14554,N_14276,N_14231);
or U14555 (N_14555,N_14396,N_14361);
or U14556 (N_14556,N_14275,N_14216);
or U14557 (N_14557,N_14260,N_14294);
and U14558 (N_14558,N_14371,N_14270);
nand U14559 (N_14559,N_14353,N_14312);
nand U14560 (N_14560,N_14356,N_14296);
and U14561 (N_14561,N_14344,N_14212);
or U14562 (N_14562,N_14366,N_14310);
and U14563 (N_14563,N_14235,N_14348);
nor U14564 (N_14564,N_14336,N_14326);
nand U14565 (N_14565,N_14258,N_14383);
and U14566 (N_14566,N_14288,N_14396);
and U14567 (N_14567,N_14367,N_14232);
nand U14568 (N_14568,N_14202,N_14344);
or U14569 (N_14569,N_14207,N_14278);
or U14570 (N_14570,N_14379,N_14258);
and U14571 (N_14571,N_14217,N_14332);
and U14572 (N_14572,N_14211,N_14247);
nor U14573 (N_14573,N_14336,N_14247);
and U14574 (N_14574,N_14336,N_14234);
and U14575 (N_14575,N_14374,N_14242);
or U14576 (N_14576,N_14330,N_14384);
nand U14577 (N_14577,N_14299,N_14278);
nor U14578 (N_14578,N_14238,N_14246);
and U14579 (N_14579,N_14285,N_14228);
nor U14580 (N_14580,N_14298,N_14230);
and U14581 (N_14581,N_14254,N_14395);
or U14582 (N_14582,N_14305,N_14337);
nor U14583 (N_14583,N_14364,N_14382);
or U14584 (N_14584,N_14284,N_14388);
and U14585 (N_14585,N_14278,N_14211);
and U14586 (N_14586,N_14374,N_14307);
and U14587 (N_14587,N_14378,N_14337);
and U14588 (N_14588,N_14355,N_14305);
and U14589 (N_14589,N_14323,N_14383);
nor U14590 (N_14590,N_14270,N_14223);
or U14591 (N_14591,N_14274,N_14257);
and U14592 (N_14592,N_14273,N_14390);
or U14593 (N_14593,N_14246,N_14371);
nor U14594 (N_14594,N_14316,N_14276);
and U14595 (N_14595,N_14391,N_14320);
xor U14596 (N_14596,N_14270,N_14312);
or U14597 (N_14597,N_14378,N_14397);
nand U14598 (N_14598,N_14339,N_14227);
nor U14599 (N_14599,N_14365,N_14394);
nand U14600 (N_14600,N_14486,N_14479);
nor U14601 (N_14601,N_14477,N_14490);
nor U14602 (N_14602,N_14571,N_14514);
nand U14603 (N_14603,N_14582,N_14584);
and U14604 (N_14604,N_14488,N_14452);
or U14605 (N_14605,N_14407,N_14579);
or U14606 (N_14606,N_14447,N_14495);
and U14607 (N_14607,N_14481,N_14501);
nand U14608 (N_14608,N_14468,N_14599);
and U14609 (N_14609,N_14478,N_14431);
and U14610 (N_14610,N_14554,N_14547);
nand U14611 (N_14611,N_14456,N_14517);
or U14612 (N_14612,N_14544,N_14442);
nor U14613 (N_14613,N_14402,N_14574);
nor U14614 (N_14614,N_14567,N_14408);
and U14615 (N_14615,N_14438,N_14570);
and U14616 (N_14616,N_14545,N_14586);
nor U14617 (N_14617,N_14469,N_14557);
nand U14618 (N_14618,N_14423,N_14404);
nand U14619 (N_14619,N_14529,N_14581);
nor U14620 (N_14620,N_14493,N_14508);
nand U14621 (N_14621,N_14418,N_14558);
and U14622 (N_14622,N_14569,N_14537);
nand U14623 (N_14623,N_14421,N_14448);
or U14624 (N_14624,N_14539,N_14577);
nor U14625 (N_14625,N_14572,N_14583);
and U14626 (N_14626,N_14453,N_14596);
nor U14627 (N_14627,N_14566,N_14565);
nor U14628 (N_14628,N_14461,N_14430);
nor U14629 (N_14629,N_14512,N_14549);
nor U14630 (N_14630,N_14428,N_14457);
nor U14631 (N_14631,N_14498,N_14410);
and U14632 (N_14632,N_14564,N_14470);
or U14633 (N_14633,N_14562,N_14521);
and U14634 (N_14634,N_14443,N_14502);
nand U14635 (N_14635,N_14482,N_14425);
nor U14636 (N_14636,N_14401,N_14411);
or U14637 (N_14637,N_14505,N_14597);
or U14638 (N_14638,N_14483,N_14429);
and U14639 (N_14639,N_14446,N_14489);
or U14640 (N_14640,N_14465,N_14585);
and U14641 (N_14641,N_14500,N_14413);
nand U14642 (N_14642,N_14523,N_14538);
or U14643 (N_14643,N_14432,N_14530);
or U14644 (N_14644,N_14471,N_14587);
nand U14645 (N_14645,N_14496,N_14476);
nor U14646 (N_14646,N_14506,N_14400);
or U14647 (N_14647,N_14563,N_14420);
nand U14648 (N_14648,N_14513,N_14590);
xor U14649 (N_14649,N_14409,N_14576);
nor U14650 (N_14650,N_14515,N_14588);
or U14651 (N_14651,N_14532,N_14541);
nand U14652 (N_14652,N_14528,N_14427);
nand U14653 (N_14653,N_14436,N_14504);
and U14654 (N_14654,N_14439,N_14459);
nand U14655 (N_14655,N_14540,N_14454);
or U14656 (N_14656,N_14426,N_14592);
and U14657 (N_14657,N_14458,N_14451);
or U14658 (N_14658,N_14499,N_14492);
or U14659 (N_14659,N_14424,N_14542);
or U14660 (N_14660,N_14526,N_14533);
and U14661 (N_14661,N_14475,N_14593);
or U14662 (N_14662,N_14524,N_14546);
and U14663 (N_14663,N_14445,N_14527);
or U14664 (N_14664,N_14511,N_14503);
and U14665 (N_14665,N_14591,N_14598);
or U14666 (N_14666,N_14464,N_14441);
or U14667 (N_14667,N_14551,N_14519);
and U14668 (N_14668,N_14487,N_14518);
nor U14669 (N_14669,N_14462,N_14485);
nand U14670 (N_14670,N_14403,N_14580);
and U14671 (N_14671,N_14437,N_14415);
and U14672 (N_14672,N_14531,N_14553);
and U14673 (N_14673,N_14520,N_14491);
nor U14674 (N_14674,N_14434,N_14522);
or U14675 (N_14675,N_14543,N_14550);
or U14676 (N_14676,N_14435,N_14422);
nand U14677 (N_14677,N_14472,N_14552);
nor U14678 (N_14678,N_14414,N_14536);
or U14679 (N_14679,N_14507,N_14473);
and U14680 (N_14680,N_14573,N_14463);
and U14681 (N_14681,N_14589,N_14417);
xnor U14682 (N_14682,N_14535,N_14561);
nor U14683 (N_14683,N_14578,N_14480);
nor U14684 (N_14684,N_14449,N_14405);
nand U14685 (N_14685,N_14412,N_14568);
nand U14686 (N_14686,N_14575,N_14525);
nand U14687 (N_14687,N_14450,N_14559);
nor U14688 (N_14688,N_14510,N_14494);
nand U14689 (N_14689,N_14484,N_14419);
nor U14690 (N_14690,N_14466,N_14594);
and U14691 (N_14691,N_14497,N_14474);
nor U14692 (N_14692,N_14516,N_14595);
nand U14693 (N_14693,N_14433,N_14440);
nand U14694 (N_14694,N_14444,N_14560);
nand U14695 (N_14695,N_14416,N_14556);
and U14696 (N_14696,N_14509,N_14460);
and U14697 (N_14697,N_14534,N_14555);
and U14698 (N_14698,N_14406,N_14467);
or U14699 (N_14699,N_14548,N_14455);
nand U14700 (N_14700,N_14443,N_14558);
nand U14701 (N_14701,N_14445,N_14466);
or U14702 (N_14702,N_14578,N_14487);
and U14703 (N_14703,N_14542,N_14462);
or U14704 (N_14704,N_14461,N_14485);
and U14705 (N_14705,N_14471,N_14448);
or U14706 (N_14706,N_14574,N_14499);
or U14707 (N_14707,N_14476,N_14556);
and U14708 (N_14708,N_14413,N_14587);
and U14709 (N_14709,N_14443,N_14592);
nand U14710 (N_14710,N_14588,N_14571);
or U14711 (N_14711,N_14560,N_14527);
nand U14712 (N_14712,N_14523,N_14473);
nand U14713 (N_14713,N_14525,N_14497);
nor U14714 (N_14714,N_14508,N_14457);
nand U14715 (N_14715,N_14488,N_14484);
and U14716 (N_14716,N_14410,N_14457);
nor U14717 (N_14717,N_14556,N_14568);
or U14718 (N_14718,N_14516,N_14562);
or U14719 (N_14719,N_14541,N_14474);
xnor U14720 (N_14720,N_14449,N_14569);
or U14721 (N_14721,N_14422,N_14473);
or U14722 (N_14722,N_14583,N_14470);
nor U14723 (N_14723,N_14496,N_14505);
nand U14724 (N_14724,N_14497,N_14599);
nor U14725 (N_14725,N_14400,N_14409);
nand U14726 (N_14726,N_14569,N_14454);
and U14727 (N_14727,N_14547,N_14502);
nand U14728 (N_14728,N_14519,N_14439);
nor U14729 (N_14729,N_14589,N_14505);
nor U14730 (N_14730,N_14462,N_14458);
nor U14731 (N_14731,N_14560,N_14477);
and U14732 (N_14732,N_14464,N_14428);
or U14733 (N_14733,N_14529,N_14477);
and U14734 (N_14734,N_14488,N_14404);
nor U14735 (N_14735,N_14579,N_14453);
and U14736 (N_14736,N_14463,N_14598);
nand U14737 (N_14737,N_14484,N_14585);
and U14738 (N_14738,N_14595,N_14487);
and U14739 (N_14739,N_14573,N_14590);
nand U14740 (N_14740,N_14475,N_14494);
and U14741 (N_14741,N_14425,N_14555);
nand U14742 (N_14742,N_14560,N_14496);
and U14743 (N_14743,N_14558,N_14422);
or U14744 (N_14744,N_14431,N_14535);
nor U14745 (N_14745,N_14487,N_14474);
nor U14746 (N_14746,N_14432,N_14446);
nand U14747 (N_14747,N_14434,N_14505);
nand U14748 (N_14748,N_14585,N_14475);
nand U14749 (N_14749,N_14494,N_14430);
nor U14750 (N_14750,N_14402,N_14414);
nor U14751 (N_14751,N_14586,N_14467);
or U14752 (N_14752,N_14532,N_14519);
nand U14753 (N_14753,N_14548,N_14418);
and U14754 (N_14754,N_14493,N_14578);
or U14755 (N_14755,N_14525,N_14583);
or U14756 (N_14756,N_14409,N_14436);
nor U14757 (N_14757,N_14546,N_14523);
nand U14758 (N_14758,N_14504,N_14423);
nor U14759 (N_14759,N_14420,N_14414);
nor U14760 (N_14760,N_14490,N_14416);
nand U14761 (N_14761,N_14442,N_14497);
nand U14762 (N_14762,N_14410,N_14515);
nor U14763 (N_14763,N_14467,N_14559);
nand U14764 (N_14764,N_14457,N_14572);
and U14765 (N_14765,N_14573,N_14500);
and U14766 (N_14766,N_14488,N_14481);
and U14767 (N_14767,N_14498,N_14423);
and U14768 (N_14768,N_14494,N_14592);
and U14769 (N_14769,N_14486,N_14449);
and U14770 (N_14770,N_14419,N_14476);
xor U14771 (N_14771,N_14404,N_14556);
nor U14772 (N_14772,N_14533,N_14505);
nor U14773 (N_14773,N_14404,N_14434);
and U14774 (N_14774,N_14411,N_14510);
or U14775 (N_14775,N_14521,N_14456);
nor U14776 (N_14776,N_14578,N_14569);
nand U14777 (N_14777,N_14425,N_14568);
or U14778 (N_14778,N_14555,N_14421);
or U14779 (N_14779,N_14443,N_14414);
nor U14780 (N_14780,N_14467,N_14523);
or U14781 (N_14781,N_14528,N_14437);
nand U14782 (N_14782,N_14590,N_14538);
nor U14783 (N_14783,N_14426,N_14577);
or U14784 (N_14784,N_14449,N_14441);
and U14785 (N_14785,N_14595,N_14596);
and U14786 (N_14786,N_14425,N_14523);
nand U14787 (N_14787,N_14470,N_14597);
nand U14788 (N_14788,N_14403,N_14448);
or U14789 (N_14789,N_14414,N_14572);
nor U14790 (N_14790,N_14485,N_14458);
and U14791 (N_14791,N_14562,N_14553);
nor U14792 (N_14792,N_14417,N_14490);
or U14793 (N_14793,N_14531,N_14528);
nand U14794 (N_14794,N_14409,N_14419);
nor U14795 (N_14795,N_14423,N_14539);
nand U14796 (N_14796,N_14413,N_14537);
and U14797 (N_14797,N_14457,N_14570);
nand U14798 (N_14798,N_14491,N_14583);
nor U14799 (N_14799,N_14528,N_14464);
or U14800 (N_14800,N_14785,N_14765);
nand U14801 (N_14801,N_14731,N_14775);
nor U14802 (N_14802,N_14619,N_14709);
nand U14803 (N_14803,N_14725,N_14728);
and U14804 (N_14804,N_14751,N_14770);
nand U14805 (N_14805,N_14767,N_14786);
nor U14806 (N_14806,N_14720,N_14636);
and U14807 (N_14807,N_14658,N_14788);
and U14808 (N_14808,N_14721,N_14620);
nand U14809 (N_14809,N_14653,N_14707);
and U14810 (N_14810,N_14714,N_14698);
nand U14811 (N_14811,N_14790,N_14673);
and U14812 (N_14812,N_14700,N_14694);
nor U14813 (N_14813,N_14647,N_14799);
xor U14814 (N_14814,N_14662,N_14645);
xnor U14815 (N_14815,N_14795,N_14683);
nor U14816 (N_14816,N_14702,N_14665);
nor U14817 (N_14817,N_14697,N_14724);
and U14818 (N_14818,N_14742,N_14611);
nor U14819 (N_14819,N_14743,N_14678);
nor U14820 (N_14820,N_14753,N_14618);
or U14821 (N_14821,N_14607,N_14726);
and U14822 (N_14822,N_14652,N_14614);
and U14823 (N_14823,N_14613,N_14755);
nand U14824 (N_14824,N_14679,N_14686);
nor U14825 (N_14825,N_14628,N_14756);
and U14826 (N_14826,N_14666,N_14732);
nand U14827 (N_14827,N_14670,N_14741);
or U14828 (N_14828,N_14669,N_14643);
or U14829 (N_14829,N_14794,N_14701);
and U14830 (N_14830,N_14718,N_14609);
or U14831 (N_14831,N_14605,N_14735);
or U14832 (N_14832,N_14740,N_14602);
nand U14833 (N_14833,N_14739,N_14604);
or U14834 (N_14834,N_14608,N_14637);
nand U14835 (N_14835,N_14733,N_14648);
or U14836 (N_14836,N_14633,N_14668);
and U14837 (N_14837,N_14711,N_14677);
nor U14838 (N_14838,N_14603,N_14684);
nand U14839 (N_14839,N_14760,N_14695);
nand U14840 (N_14840,N_14624,N_14761);
nor U14841 (N_14841,N_14617,N_14764);
or U14842 (N_14842,N_14708,N_14716);
or U14843 (N_14843,N_14749,N_14699);
and U14844 (N_14844,N_14746,N_14793);
nand U14845 (N_14845,N_14623,N_14690);
nor U14846 (N_14846,N_14771,N_14693);
and U14847 (N_14847,N_14757,N_14789);
or U14848 (N_14848,N_14622,N_14736);
and U14849 (N_14849,N_14696,N_14675);
and U14850 (N_14850,N_14766,N_14631);
and U14851 (N_14851,N_14655,N_14730);
or U14852 (N_14852,N_14774,N_14745);
or U14853 (N_14853,N_14649,N_14776);
nand U14854 (N_14854,N_14710,N_14606);
or U14855 (N_14855,N_14763,N_14674);
nor U14856 (N_14856,N_14772,N_14657);
or U14857 (N_14857,N_14600,N_14682);
nor U14858 (N_14858,N_14722,N_14797);
nor U14859 (N_14859,N_14712,N_14621);
and U14860 (N_14860,N_14689,N_14681);
or U14861 (N_14861,N_14784,N_14717);
or U14862 (N_14862,N_14773,N_14676);
nor U14863 (N_14863,N_14651,N_14632);
and U14864 (N_14864,N_14642,N_14644);
nand U14865 (N_14865,N_14692,N_14646);
nor U14866 (N_14866,N_14758,N_14672);
and U14867 (N_14867,N_14792,N_14659);
or U14868 (N_14868,N_14738,N_14744);
or U14869 (N_14869,N_14664,N_14635);
nand U14870 (N_14870,N_14660,N_14791);
and U14871 (N_14871,N_14782,N_14705);
nor U14872 (N_14872,N_14727,N_14729);
nor U14873 (N_14873,N_14734,N_14612);
and U14874 (N_14874,N_14601,N_14796);
nand U14875 (N_14875,N_14610,N_14777);
nand U14876 (N_14876,N_14661,N_14750);
nor U14877 (N_14877,N_14687,N_14783);
nor U14878 (N_14878,N_14754,N_14667);
nand U14879 (N_14879,N_14768,N_14703);
and U14880 (N_14880,N_14639,N_14656);
and U14881 (N_14881,N_14630,N_14723);
and U14882 (N_14882,N_14778,N_14663);
or U14883 (N_14883,N_14634,N_14737);
nor U14884 (N_14884,N_14779,N_14638);
or U14885 (N_14885,N_14625,N_14706);
and U14886 (N_14886,N_14654,N_14715);
nand U14887 (N_14887,N_14616,N_14650);
or U14888 (N_14888,N_14615,N_14719);
nor U14889 (N_14889,N_14691,N_14629);
nor U14890 (N_14890,N_14780,N_14627);
nor U14891 (N_14891,N_14781,N_14762);
and U14892 (N_14892,N_14688,N_14626);
or U14893 (N_14893,N_14787,N_14769);
and U14894 (N_14894,N_14671,N_14747);
nor U14895 (N_14895,N_14713,N_14759);
nor U14896 (N_14896,N_14680,N_14748);
nor U14897 (N_14897,N_14752,N_14640);
nor U14898 (N_14898,N_14798,N_14685);
nand U14899 (N_14899,N_14641,N_14704);
nor U14900 (N_14900,N_14603,N_14774);
nor U14901 (N_14901,N_14787,N_14679);
nand U14902 (N_14902,N_14741,N_14631);
or U14903 (N_14903,N_14788,N_14784);
nand U14904 (N_14904,N_14606,N_14752);
or U14905 (N_14905,N_14688,N_14689);
or U14906 (N_14906,N_14721,N_14621);
nand U14907 (N_14907,N_14707,N_14756);
nor U14908 (N_14908,N_14792,N_14741);
and U14909 (N_14909,N_14640,N_14704);
and U14910 (N_14910,N_14791,N_14666);
xor U14911 (N_14911,N_14632,N_14795);
nand U14912 (N_14912,N_14663,N_14628);
and U14913 (N_14913,N_14715,N_14718);
or U14914 (N_14914,N_14688,N_14649);
and U14915 (N_14915,N_14776,N_14610);
nor U14916 (N_14916,N_14787,N_14695);
nor U14917 (N_14917,N_14780,N_14741);
and U14918 (N_14918,N_14794,N_14629);
nor U14919 (N_14919,N_14639,N_14600);
nand U14920 (N_14920,N_14731,N_14601);
or U14921 (N_14921,N_14752,N_14712);
nand U14922 (N_14922,N_14798,N_14645);
nand U14923 (N_14923,N_14600,N_14655);
nor U14924 (N_14924,N_14646,N_14716);
nor U14925 (N_14925,N_14631,N_14796);
nor U14926 (N_14926,N_14624,N_14640);
nand U14927 (N_14927,N_14773,N_14684);
or U14928 (N_14928,N_14796,N_14674);
nand U14929 (N_14929,N_14667,N_14680);
or U14930 (N_14930,N_14668,N_14657);
and U14931 (N_14931,N_14756,N_14787);
nand U14932 (N_14932,N_14641,N_14675);
or U14933 (N_14933,N_14648,N_14637);
and U14934 (N_14934,N_14782,N_14608);
nor U14935 (N_14935,N_14709,N_14647);
and U14936 (N_14936,N_14786,N_14743);
nor U14937 (N_14937,N_14616,N_14699);
nand U14938 (N_14938,N_14601,N_14798);
nand U14939 (N_14939,N_14636,N_14713);
nor U14940 (N_14940,N_14791,N_14686);
nor U14941 (N_14941,N_14690,N_14709);
or U14942 (N_14942,N_14666,N_14725);
and U14943 (N_14943,N_14687,N_14784);
or U14944 (N_14944,N_14753,N_14620);
nor U14945 (N_14945,N_14659,N_14653);
and U14946 (N_14946,N_14646,N_14673);
or U14947 (N_14947,N_14637,N_14711);
nor U14948 (N_14948,N_14717,N_14611);
nand U14949 (N_14949,N_14747,N_14692);
and U14950 (N_14950,N_14650,N_14770);
nor U14951 (N_14951,N_14708,N_14726);
nand U14952 (N_14952,N_14644,N_14732);
and U14953 (N_14953,N_14750,N_14601);
nand U14954 (N_14954,N_14744,N_14705);
nand U14955 (N_14955,N_14757,N_14663);
or U14956 (N_14956,N_14707,N_14602);
and U14957 (N_14957,N_14655,N_14608);
and U14958 (N_14958,N_14699,N_14697);
nor U14959 (N_14959,N_14717,N_14648);
or U14960 (N_14960,N_14762,N_14644);
nand U14961 (N_14961,N_14694,N_14630);
nand U14962 (N_14962,N_14701,N_14642);
and U14963 (N_14963,N_14764,N_14724);
and U14964 (N_14964,N_14617,N_14723);
nand U14965 (N_14965,N_14684,N_14659);
nor U14966 (N_14966,N_14693,N_14647);
nor U14967 (N_14967,N_14708,N_14631);
and U14968 (N_14968,N_14633,N_14667);
and U14969 (N_14969,N_14618,N_14624);
nor U14970 (N_14970,N_14737,N_14608);
nand U14971 (N_14971,N_14648,N_14724);
nand U14972 (N_14972,N_14631,N_14794);
nand U14973 (N_14973,N_14617,N_14644);
nor U14974 (N_14974,N_14772,N_14633);
or U14975 (N_14975,N_14622,N_14741);
or U14976 (N_14976,N_14778,N_14799);
nand U14977 (N_14977,N_14769,N_14701);
nand U14978 (N_14978,N_14620,N_14742);
or U14979 (N_14979,N_14745,N_14711);
nand U14980 (N_14980,N_14717,N_14632);
or U14981 (N_14981,N_14617,N_14799);
nand U14982 (N_14982,N_14636,N_14678);
and U14983 (N_14983,N_14728,N_14775);
nand U14984 (N_14984,N_14662,N_14648);
or U14985 (N_14985,N_14741,N_14607);
nand U14986 (N_14986,N_14638,N_14783);
and U14987 (N_14987,N_14777,N_14612);
or U14988 (N_14988,N_14683,N_14692);
nor U14989 (N_14989,N_14651,N_14709);
and U14990 (N_14990,N_14654,N_14734);
nor U14991 (N_14991,N_14739,N_14736);
or U14992 (N_14992,N_14660,N_14760);
and U14993 (N_14993,N_14708,N_14792);
nor U14994 (N_14994,N_14701,N_14653);
and U14995 (N_14995,N_14745,N_14616);
or U14996 (N_14996,N_14631,N_14729);
and U14997 (N_14997,N_14651,N_14615);
nor U14998 (N_14998,N_14683,N_14688);
and U14999 (N_14999,N_14767,N_14648);
or U15000 (N_15000,N_14981,N_14955);
nand U15001 (N_15001,N_14992,N_14947);
nand U15002 (N_15002,N_14970,N_14968);
nor U15003 (N_15003,N_14809,N_14959);
nor U15004 (N_15004,N_14816,N_14935);
or U15005 (N_15005,N_14908,N_14838);
nor U15006 (N_15006,N_14821,N_14817);
nor U15007 (N_15007,N_14983,N_14842);
or U15008 (N_15008,N_14899,N_14876);
nand U15009 (N_15009,N_14930,N_14934);
and U15010 (N_15010,N_14931,N_14898);
and U15011 (N_15011,N_14951,N_14907);
or U15012 (N_15012,N_14818,N_14873);
nor U15013 (N_15013,N_14895,N_14807);
nor U15014 (N_15014,N_14962,N_14990);
and U15015 (N_15015,N_14946,N_14917);
or U15016 (N_15016,N_14815,N_14841);
nor U15017 (N_15017,N_14830,N_14874);
nor U15018 (N_15018,N_14918,N_14997);
nand U15019 (N_15019,N_14912,N_14958);
or U15020 (N_15020,N_14971,N_14919);
nor U15021 (N_15021,N_14848,N_14902);
or U15022 (N_15022,N_14984,N_14871);
nand U15023 (N_15023,N_14857,N_14800);
nand U15024 (N_15024,N_14811,N_14808);
and U15025 (N_15025,N_14836,N_14826);
and U15026 (N_15026,N_14878,N_14843);
or U15027 (N_15027,N_14952,N_14945);
or U15028 (N_15028,N_14977,N_14846);
nor U15029 (N_15029,N_14812,N_14966);
nand U15030 (N_15030,N_14802,N_14923);
nand U15031 (N_15031,N_14890,N_14999);
nand U15032 (N_15032,N_14996,N_14879);
or U15033 (N_15033,N_14928,N_14906);
or U15034 (N_15034,N_14853,N_14834);
or U15035 (N_15035,N_14850,N_14900);
nor U15036 (N_15036,N_14921,N_14889);
nor U15037 (N_15037,N_14832,N_14909);
nand U15038 (N_15038,N_14941,N_14974);
nand U15039 (N_15039,N_14915,N_14922);
nor U15040 (N_15040,N_14861,N_14979);
nor U15041 (N_15041,N_14901,N_14872);
or U15042 (N_15042,N_14953,N_14829);
nand U15043 (N_15043,N_14804,N_14998);
nor U15044 (N_15044,N_14885,N_14939);
and U15045 (N_15045,N_14880,N_14932);
nor U15046 (N_15046,N_14867,N_14839);
nor U15047 (N_15047,N_14882,N_14913);
and U15048 (N_15048,N_14852,N_14929);
nand U15049 (N_15049,N_14863,N_14933);
nand U15050 (N_15050,N_14956,N_14875);
nor U15051 (N_15051,N_14858,N_14859);
and U15052 (N_15052,N_14987,N_14887);
and U15053 (N_15053,N_14914,N_14856);
and U15054 (N_15054,N_14940,N_14963);
and U15055 (N_15055,N_14891,N_14969);
or U15056 (N_15056,N_14851,N_14820);
nand U15057 (N_15057,N_14944,N_14903);
and U15058 (N_15058,N_14866,N_14868);
and U15059 (N_15059,N_14877,N_14828);
nor U15060 (N_15060,N_14835,N_14831);
and U15061 (N_15061,N_14936,N_14973);
nand U15062 (N_15062,N_14991,N_14823);
nand U15063 (N_15063,N_14819,N_14814);
nand U15064 (N_15064,N_14911,N_14943);
or U15065 (N_15065,N_14884,N_14972);
or U15066 (N_15066,N_14822,N_14916);
or U15067 (N_15067,N_14950,N_14849);
nor U15068 (N_15068,N_14942,N_14869);
nand U15069 (N_15069,N_14905,N_14982);
nor U15070 (N_15070,N_14833,N_14840);
nand U15071 (N_15071,N_14847,N_14825);
and U15072 (N_15072,N_14813,N_14926);
and U15073 (N_15073,N_14976,N_14855);
nand U15074 (N_15074,N_14961,N_14938);
and U15075 (N_15075,N_14967,N_14949);
or U15076 (N_15076,N_14827,N_14965);
and U15077 (N_15077,N_14986,N_14978);
or U15078 (N_15078,N_14960,N_14892);
and U15079 (N_15079,N_14844,N_14881);
nor U15080 (N_15080,N_14925,N_14870);
or U15081 (N_15081,N_14888,N_14837);
nor U15082 (N_15082,N_14862,N_14805);
nand U15083 (N_15083,N_14824,N_14893);
nor U15084 (N_15084,N_14806,N_14860);
and U15085 (N_15085,N_14896,N_14994);
nor U15086 (N_15086,N_14988,N_14985);
or U15087 (N_15087,N_14937,N_14995);
nand U15088 (N_15088,N_14904,N_14886);
nor U15089 (N_15089,N_14883,N_14865);
nor U15090 (N_15090,N_14989,N_14927);
nand U15091 (N_15091,N_14845,N_14801);
and U15092 (N_15092,N_14957,N_14803);
and U15093 (N_15093,N_14810,N_14894);
or U15094 (N_15094,N_14910,N_14897);
nor U15095 (N_15095,N_14948,N_14993);
nand U15096 (N_15096,N_14954,N_14920);
and U15097 (N_15097,N_14924,N_14980);
and U15098 (N_15098,N_14975,N_14864);
or U15099 (N_15099,N_14854,N_14964);
and U15100 (N_15100,N_14885,N_14808);
nand U15101 (N_15101,N_14979,N_14961);
nor U15102 (N_15102,N_14828,N_14819);
or U15103 (N_15103,N_14941,N_14897);
and U15104 (N_15104,N_14995,N_14846);
nor U15105 (N_15105,N_14989,N_14858);
or U15106 (N_15106,N_14954,N_14870);
nand U15107 (N_15107,N_14939,N_14849);
or U15108 (N_15108,N_14903,N_14825);
nor U15109 (N_15109,N_14939,N_14949);
nand U15110 (N_15110,N_14817,N_14998);
nand U15111 (N_15111,N_14840,N_14874);
nand U15112 (N_15112,N_14827,N_14921);
and U15113 (N_15113,N_14820,N_14871);
or U15114 (N_15114,N_14915,N_14808);
or U15115 (N_15115,N_14900,N_14849);
nor U15116 (N_15116,N_14967,N_14894);
xnor U15117 (N_15117,N_14859,N_14944);
nand U15118 (N_15118,N_14863,N_14804);
or U15119 (N_15119,N_14990,N_14868);
or U15120 (N_15120,N_14894,N_14977);
nor U15121 (N_15121,N_14828,N_14917);
or U15122 (N_15122,N_14892,N_14947);
and U15123 (N_15123,N_14820,N_14965);
or U15124 (N_15124,N_14855,N_14939);
and U15125 (N_15125,N_14958,N_14979);
and U15126 (N_15126,N_14883,N_14866);
and U15127 (N_15127,N_14820,N_14824);
and U15128 (N_15128,N_14879,N_14831);
or U15129 (N_15129,N_14957,N_14925);
or U15130 (N_15130,N_14889,N_14837);
nand U15131 (N_15131,N_14806,N_14978);
and U15132 (N_15132,N_14895,N_14901);
nand U15133 (N_15133,N_14843,N_14886);
nand U15134 (N_15134,N_14942,N_14991);
or U15135 (N_15135,N_14987,N_14810);
and U15136 (N_15136,N_14962,N_14852);
nand U15137 (N_15137,N_14805,N_14956);
and U15138 (N_15138,N_14991,N_14870);
nor U15139 (N_15139,N_14859,N_14845);
and U15140 (N_15140,N_14908,N_14933);
xnor U15141 (N_15141,N_14945,N_14950);
nand U15142 (N_15142,N_14817,N_14865);
or U15143 (N_15143,N_14942,N_14911);
nand U15144 (N_15144,N_14974,N_14888);
and U15145 (N_15145,N_14984,N_14854);
nand U15146 (N_15146,N_14955,N_14835);
and U15147 (N_15147,N_14986,N_14865);
or U15148 (N_15148,N_14871,N_14962);
nand U15149 (N_15149,N_14944,N_14892);
and U15150 (N_15150,N_14829,N_14986);
and U15151 (N_15151,N_14809,N_14921);
or U15152 (N_15152,N_14996,N_14979);
nor U15153 (N_15153,N_14986,N_14875);
or U15154 (N_15154,N_14898,N_14905);
or U15155 (N_15155,N_14903,N_14898);
and U15156 (N_15156,N_14878,N_14865);
or U15157 (N_15157,N_14915,N_14863);
or U15158 (N_15158,N_14965,N_14805);
nor U15159 (N_15159,N_14856,N_14885);
or U15160 (N_15160,N_14863,N_14883);
nor U15161 (N_15161,N_14836,N_14974);
nand U15162 (N_15162,N_14824,N_14938);
nand U15163 (N_15163,N_14819,N_14897);
nor U15164 (N_15164,N_14833,N_14888);
nand U15165 (N_15165,N_14898,N_14996);
nor U15166 (N_15166,N_14924,N_14973);
nor U15167 (N_15167,N_14910,N_14913);
and U15168 (N_15168,N_14804,N_14824);
and U15169 (N_15169,N_14875,N_14914);
and U15170 (N_15170,N_14840,N_14819);
and U15171 (N_15171,N_14878,N_14968);
and U15172 (N_15172,N_14948,N_14990);
nand U15173 (N_15173,N_14926,N_14943);
and U15174 (N_15174,N_14985,N_14995);
nand U15175 (N_15175,N_14985,N_14908);
and U15176 (N_15176,N_14805,N_14917);
nor U15177 (N_15177,N_14846,N_14864);
or U15178 (N_15178,N_14873,N_14864);
nor U15179 (N_15179,N_14959,N_14820);
nor U15180 (N_15180,N_14981,N_14991);
or U15181 (N_15181,N_14997,N_14840);
nand U15182 (N_15182,N_14964,N_14853);
or U15183 (N_15183,N_14855,N_14892);
nor U15184 (N_15184,N_14808,N_14889);
or U15185 (N_15185,N_14870,N_14823);
and U15186 (N_15186,N_14978,N_14913);
or U15187 (N_15187,N_14846,N_14842);
or U15188 (N_15188,N_14877,N_14848);
and U15189 (N_15189,N_14963,N_14907);
or U15190 (N_15190,N_14922,N_14887);
nor U15191 (N_15191,N_14822,N_14863);
nor U15192 (N_15192,N_14918,N_14945);
and U15193 (N_15193,N_14868,N_14896);
or U15194 (N_15194,N_14869,N_14967);
and U15195 (N_15195,N_14828,N_14919);
and U15196 (N_15196,N_14886,N_14954);
and U15197 (N_15197,N_14858,N_14807);
nand U15198 (N_15198,N_14836,N_14817);
or U15199 (N_15199,N_14801,N_14885);
or U15200 (N_15200,N_15196,N_15165);
nand U15201 (N_15201,N_15081,N_15099);
nor U15202 (N_15202,N_15025,N_15054);
or U15203 (N_15203,N_15132,N_15193);
nand U15204 (N_15204,N_15169,N_15119);
nor U15205 (N_15205,N_15114,N_15166);
nor U15206 (N_15206,N_15194,N_15195);
or U15207 (N_15207,N_15177,N_15189);
nor U15208 (N_15208,N_15153,N_15098);
nand U15209 (N_15209,N_15125,N_15120);
nor U15210 (N_15210,N_15086,N_15064);
and U15211 (N_15211,N_15101,N_15142);
or U15212 (N_15212,N_15073,N_15012);
nand U15213 (N_15213,N_15009,N_15109);
or U15214 (N_15214,N_15106,N_15036);
nand U15215 (N_15215,N_15097,N_15160);
and U15216 (N_15216,N_15066,N_15171);
or U15217 (N_15217,N_15157,N_15181);
and U15218 (N_15218,N_15108,N_15198);
or U15219 (N_15219,N_15063,N_15031);
nor U15220 (N_15220,N_15071,N_15137);
and U15221 (N_15221,N_15183,N_15180);
and U15222 (N_15222,N_15000,N_15083);
nand U15223 (N_15223,N_15069,N_15013);
nand U15224 (N_15224,N_15028,N_15006);
nor U15225 (N_15225,N_15050,N_15035);
and U15226 (N_15226,N_15123,N_15082);
and U15227 (N_15227,N_15131,N_15170);
nor U15228 (N_15228,N_15162,N_15041);
and U15229 (N_15229,N_15161,N_15156);
nand U15230 (N_15230,N_15053,N_15058);
nand U15231 (N_15231,N_15047,N_15048);
or U15232 (N_15232,N_15004,N_15010);
nand U15233 (N_15233,N_15062,N_15118);
nor U15234 (N_15234,N_15045,N_15024);
nor U15235 (N_15235,N_15061,N_15184);
nand U15236 (N_15236,N_15027,N_15002);
and U15237 (N_15237,N_15107,N_15017);
and U15238 (N_15238,N_15136,N_15147);
nand U15239 (N_15239,N_15032,N_15164);
nor U15240 (N_15240,N_15130,N_15117);
nand U15241 (N_15241,N_15080,N_15011);
and U15242 (N_15242,N_15085,N_15178);
xor U15243 (N_15243,N_15043,N_15057);
xor U15244 (N_15244,N_15140,N_15089);
nand U15245 (N_15245,N_15187,N_15105);
nand U15246 (N_15246,N_15172,N_15020);
nand U15247 (N_15247,N_15015,N_15021);
and U15248 (N_15248,N_15019,N_15126);
nor U15249 (N_15249,N_15093,N_15176);
nand U15250 (N_15250,N_15168,N_15092);
or U15251 (N_15251,N_15110,N_15113);
nor U15252 (N_15252,N_15135,N_15016);
or U15253 (N_15253,N_15128,N_15046);
nor U15254 (N_15254,N_15077,N_15145);
nor U15255 (N_15255,N_15173,N_15072);
nor U15256 (N_15256,N_15040,N_15138);
and U15257 (N_15257,N_15174,N_15076);
and U15258 (N_15258,N_15056,N_15129);
or U15259 (N_15259,N_15005,N_15094);
nor U15260 (N_15260,N_15008,N_15122);
nor U15261 (N_15261,N_15014,N_15095);
and U15262 (N_15262,N_15112,N_15087);
nor U15263 (N_15263,N_15154,N_15018);
nand U15264 (N_15264,N_15111,N_15022);
or U15265 (N_15265,N_15052,N_15148);
nand U15266 (N_15266,N_15182,N_15023);
nor U15267 (N_15267,N_15175,N_15103);
nor U15268 (N_15268,N_15116,N_15084);
or U15269 (N_15269,N_15030,N_15078);
nor U15270 (N_15270,N_15060,N_15075);
or U15271 (N_15271,N_15143,N_15074);
nor U15272 (N_15272,N_15096,N_15124);
or U15273 (N_15273,N_15034,N_15144);
and U15274 (N_15274,N_15197,N_15067);
or U15275 (N_15275,N_15146,N_15091);
nor U15276 (N_15276,N_15199,N_15029);
and U15277 (N_15277,N_15100,N_15121);
and U15278 (N_15278,N_15186,N_15167);
and U15279 (N_15279,N_15051,N_15104);
and U15280 (N_15280,N_15163,N_15150);
nor U15281 (N_15281,N_15151,N_15133);
or U15282 (N_15282,N_15155,N_15134);
and U15283 (N_15283,N_15068,N_15044);
nor U15284 (N_15284,N_15039,N_15159);
and U15285 (N_15285,N_15042,N_15033);
or U15286 (N_15286,N_15001,N_15127);
or U15287 (N_15287,N_15079,N_15038);
or U15288 (N_15288,N_15115,N_15049);
nand U15289 (N_15289,N_15188,N_15055);
or U15290 (N_15290,N_15192,N_15152);
and U15291 (N_15291,N_15090,N_15088);
nor U15292 (N_15292,N_15190,N_15026);
or U15293 (N_15293,N_15102,N_15007);
nor U15294 (N_15294,N_15065,N_15059);
nor U15295 (N_15295,N_15158,N_15191);
or U15296 (N_15296,N_15037,N_15149);
nand U15297 (N_15297,N_15141,N_15003);
and U15298 (N_15298,N_15185,N_15179);
nand U15299 (N_15299,N_15139,N_15070);
and U15300 (N_15300,N_15059,N_15001);
or U15301 (N_15301,N_15178,N_15009);
or U15302 (N_15302,N_15108,N_15035);
nand U15303 (N_15303,N_15045,N_15030);
nand U15304 (N_15304,N_15155,N_15104);
nor U15305 (N_15305,N_15075,N_15036);
nand U15306 (N_15306,N_15044,N_15082);
nand U15307 (N_15307,N_15190,N_15057);
or U15308 (N_15308,N_15136,N_15126);
or U15309 (N_15309,N_15020,N_15189);
or U15310 (N_15310,N_15034,N_15134);
or U15311 (N_15311,N_15017,N_15023);
and U15312 (N_15312,N_15025,N_15171);
nor U15313 (N_15313,N_15090,N_15040);
or U15314 (N_15314,N_15093,N_15019);
nand U15315 (N_15315,N_15038,N_15195);
nor U15316 (N_15316,N_15142,N_15182);
nor U15317 (N_15317,N_15060,N_15177);
or U15318 (N_15318,N_15195,N_15080);
xor U15319 (N_15319,N_15184,N_15091);
nand U15320 (N_15320,N_15025,N_15030);
nand U15321 (N_15321,N_15128,N_15148);
nor U15322 (N_15322,N_15170,N_15169);
nand U15323 (N_15323,N_15002,N_15192);
nand U15324 (N_15324,N_15073,N_15128);
nand U15325 (N_15325,N_15079,N_15054);
nand U15326 (N_15326,N_15163,N_15118);
nor U15327 (N_15327,N_15080,N_15082);
xnor U15328 (N_15328,N_15196,N_15077);
nor U15329 (N_15329,N_15198,N_15045);
nor U15330 (N_15330,N_15194,N_15079);
and U15331 (N_15331,N_15023,N_15016);
nand U15332 (N_15332,N_15056,N_15024);
nand U15333 (N_15333,N_15013,N_15121);
nand U15334 (N_15334,N_15150,N_15114);
nor U15335 (N_15335,N_15136,N_15007);
nand U15336 (N_15336,N_15125,N_15072);
nand U15337 (N_15337,N_15027,N_15163);
and U15338 (N_15338,N_15077,N_15146);
nor U15339 (N_15339,N_15039,N_15049);
nand U15340 (N_15340,N_15085,N_15056);
nand U15341 (N_15341,N_15120,N_15034);
and U15342 (N_15342,N_15067,N_15051);
nor U15343 (N_15343,N_15089,N_15079);
nand U15344 (N_15344,N_15061,N_15082);
nand U15345 (N_15345,N_15159,N_15176);
nand U15346 (N_15346,N_15085,N_15184);
nand U15347 (N_15347,N_15032,N_15119);
and U15348 (N_15348,N_15125,N_15028);
nor U15349 (N_15349,N_15180,N_15081);
nand U15350 (N_15350,N_15130,N_15047);
or U15351 (N_15351,N_15083,N_15088);
or U15352 (N_15352,N_15016,N_15121);
and U15353 (N_15353,N_15195,N_15104);
or U15354 (N_15354,N_15054,N_15037);
or U15355 (N_15355,N_15035,N_15069);
and U15356 (N_15356,N_15135,N_15024);
nor U15357 (N_15357,N_15045,N_15085);
or U15358 (N_15358,N_15085,N_15042);
nor U15359 (N_15359,N_15057,N_15051);
and U15360 (N_15360,N_15042,N_15157);
or U15361 (N_15361,N_15042,N_15126);
or U15362 (N_15362,N_15001,N_15159);
or U15363 (N_15363,N_15134,N_15115);
nor U15364 (N_15364,N_15083,N_15181);
and U15365 (N_15365,N_15045,N_15104);
and U15366 (N_15366,N_15199,N_15066);
or U15367 (N_15367,N_15049,N_15141);
or U15368 (N_15368,N_15035,N_15196);
nor U15369 (N_15369,N_15076,N_15059);
nor U15370 (N_15370,N_15102,N_15079);
nor U15371 (N_15371,N_15058,N_15087);
nand U15372 (N_15372,N_15085,N_15180);
nand U15373 (N_15373,N_15159,N_15065);
or U15374 (N_15374,N_15136,N_15030);
or U15375 (N_15375,N_15118,N_15179);
nand U15376 (N_15376,N_15008,N_15117);
nand U15377 (N_15377,N_15028,N_15190);
nor U15378 (N_15378,N_15042,N_15060);
nand U15379 (N_15379,N_15167,N_15178);
xor U15380 (N_15380,N_15144,N_15127);
and U15381 (N_15381,N_15142,N_15151);
and U15382 (N_15382,N_15012,N_15185);
nor U15383 (N_15383,N_15019,N_15117);
nand U15384 (N_15384,N_15163,N_15178);
and U15385 (N_15385,N_15006,N_15112);
or U15386 (N_15386,N_15037,N_15116);
and U15387 (N_15387,N_15166,N_15038);
nand U15388 (N_15388,N_15056,N_15014);
nor U15389 (N_15389,N_15189,N_15182);
nor U15390 (N_15390,N_15199,N_15044);
nand U15391 (N_15391,N_15100,N_15041);
nor U15392 (N_15392,N_15101,N_15049);
and U15393 (N_15393,N_15113,N_15026);
and U15394 (N_15394,N_15087,N_15079);
nand U15395 (N_15395,N_15093,N_15161);
and U15396 (N_15396,N_15197,N_15129);
and U15397 (N_15397,N_15008,N_15162);
nand U15398 (N_15398,N_15117,N_15054);
and U15399 (N_15399,N_15140,N_15110);
nor U15400 (N_15400,N_15265,N_15325);
and U15401 (N_15401,N_15260,N_15218);
or U15402 (N_15402,N_15298,N_15305);
nor U15403 (N_15403,N_15248,N_15376);
and U15404 (N_15404,N_15324,N_15285);
and U15405 (N_15405,N_15261,N_15322);
or U15406 (N_15406,N_15219,N_15399);
or U15407 (N_15407,N_15317,N_15269);
and U15408 (N_15408,N_15366,N_15396);
or U15409 (N_15409,N_15283,N_15313);
or U15410 (N_15410,N_15337,N_15223);
or U15411 (N_15411,N_15369,N_15217);
and U15412 (N_15412,N_15276,N_15206);
nand U15413 (N_15413,N_15247,N_15339);
nand U15414 (N_15414,N_15213,N_15304);
nand U15415 (N_15415,N_15352,N_15258);
nand U15416 (N_15416,N_15377,N_15364);
nand U15417 (N_15417,N_15245,N_15240);
nand U15418 (N_15418,N_15365,N_15264);
or U15419 (N_15419,N_15312,N_15379);
nor U15420 (N_15420,N_15381,N_15386);
nand U15421 (N_15421,N_15235,N_15303);
and U15422 (N_15422,N_15343,N_15233);
nand U15423 (N_15423,N_15315,N_15387);
and U15424 (N_15424,N_15268,N_15336);
and U15425 (N_15425,N_15210,N_15200);
nor U15426 (N_15426,N_15277,N_15393);
nand U15427 (N_15427,N_15249,N_15342);
or U15428 (N_15428,N_15215,N_15358);
nor U15429 (N_15429,N_15267,N_15321);
nor U15430 (N_15430,N_15284,N_15212);
nand U15431 (N_15431,N_15203,N_15356);
nor U15432 (N_15432,N_15344,N_15397);
and U15433 (N_15433,N_15238,N_15237);
nand U15434 (N_15434,N_15357,N_15348);
nor U15435 (N_15435,N_15263,N_15306);
nand U15436 (N_15436,N_15380,N_15333);
or U15437 (N_15437,N_15273,N_15241);
nand U15438 (N_15438,N_15394,N_15355);
nor U15439 (N_15439,N_15271,N_15205);
and U15440 (N_15440,N_15359,N_15328);
or U15441 (N_15441,N_15391,N_15289);
nor U15442 (N_15442,N_15367,N_15294);
and U15443 (N_15443,N_15278,N_15214);
nand U15444 (N_15444,N_15299,N_15346);
nor U15445 (N_15445,N_15291,N_15384);
or U15446 (N_15446,N_15310,N_15383);
nand U15447 (N_15447,N_15287,N_15202);
nor U15448 (N_15448,N_15349,N_15388);
and U15449 (N_15449,N_15266,N_15209);
nand U15450 (N_15450,N_15272,N_15234);
nand U15451 (N_15451,N_15253,N_15300);
nor U15452 (N_15452,N_15373,N_15318);
nand U15453 (N_15453,N_15230,N_15224);
nand U15454 (N_15454,N_15243,N_15208);
or U15455 (N_15455,N_15309,N_15329);
nand U15456 (N_15456,N_15244,N_15251);
or U15457 (N_15457,N_15341,N_15362);
and U15458 (N_15458,N_15374,N_15211);
and U15459 (N_15459,N_15331,N_15389);
nor U15460 (N_15460,N_15281,N_15257);
nor U15461 (N_15461,N_15347,N_15262);
nand U15462 (N_15462,N_15232,N_15368);
nor U15463 (N_15463,N_15293,N_15330);
and U15464 (N_15464,N_15351,N_15274);
nand U15465 (N_15465,N_15398,N_15220);
nand U15466 (N_15466,N_15207,N_15334);
nand U15467 (N_15467,N_15361,N_15259);
nor U15468 (N_15468,N_15239,N_15255);
nand U15469 (N_15469,N_15226,N_15320);
nor U15470 (N_15470,N_15382,N_15372);
or U15471 (N_15471,N_15360,N_15326);
or U15472 (N_15472,N_15280,N_15201);
nand U15473 (N_15473,N_15363,N_15275);
nand U15474 (N_15474,N_15345,N_15254);
nor U15475 (N_15475,N_15395,N_15270);
xnor U15476 (N_15476,N_15282,N_15332);
nor U15477 (N_15477,N_15250,N_15290);
nand U15478 (N_15478,N_15296,N_15375);
and U15479 (N_15479,N_15301,N_15231);
nand U15480 (N_15480,N_15246,N_15390);
nor U15481 (N_15481,N_15204,N_15221);
nor U15482 (N_15482,N_15319,N_15385);
and U15483 (N_15483,N_15314,N_15316);
and U15484 (N_15484,N_15236,N_15295);
and U15485 (N_15485,N_15279,N_15256);
nor U15486 (N_15486,N_15392,N_15340);
or U15487 (N_15487,N_15371,N_15353);
or U15488 (N_15488,N_15216,N_15242);
or U15489 (N_15489,N_15335,N_15228);
nand U15490 (N_15490,N_15292,N_15350);
or U15491 (N_15491,N_15327,N_15302);
or U15492 (N_15492,N_15370,N_15222);
nor U15493 (N_15493,N_15307,N_15227);
and U15494 (N_15494,N_15229,N_15311);
or U15495 (N_15495,N_15378,N_15308);
nor U15496 (N_15496,N_15286,N_15354);
or U15497 (N_15497,N_15323,N_15338);
or U15498 (N_15498,N_15252,N_15288);
nand U15499 (N_15499,N_15297,N_15225);
nand U15500 (N_15500,N_15397,N_15212);
xnor U15501 (N_15501,N_15374,N_15323);
nand U15502 (N_15502,N_15215,N_15364);
nor U15503 (N_15503,N_15204,N_15383);
nand U15504 (N_15504,N_15390,N_15232);
and U15505 (N_15505,N_15201,N_15229);
and U15506 (N_15506,N_15256,N_15330);
or U15507 (N_15507,N_15295,N_15376);
or U15508 (N_15508,N_15200,N_15362);
nand U15509 (N_15509,N_15301,N_15310);
or U15510 (N_15510,N_15232,N_15358);
or U15511 (N_15511,N_15357,N_15224);
or U15512 (N_15512,N_15364,N_15356);
nand U15513 (N_15513,N_15200,N_15345);
and U15514 (N_15514,N_15270,N_15293);
nor U15515 (N_15515,N_15283,N_15296);
nand U15516 (N_15516,N_15268,N_15355);
or U15517 (N_15517,N_15225,N_15279);
and U15518 (N_15518,N_15232,N_15270);
nand U15519 (N_15519,N_15272,N_15216);
or U15520 (N_15520,N_15230,N_15283);
nor U15521 (N_15521,N_15230,N_15213);
or U15522 (N_15522,N_15306,N_15283);
or U15523 (N_15523,N_15268,N_15231);
nand U15524 (N_15524,N_15395,N_15248);
nand U15525 (N_15525,N_15362,N_15277);
nand U15526 (N_15526,N_15309,N_15242);
nor U15527 (N_15527,N_15258,N_15338);
or U15528 (N_15528,N_15336,N_15338);
or U15529 (N_15529,N_15299,N_15219);
nand U15530 (N_15530,N_15310,N_15289);
or U15531 (N_15531,N_15347,N_15284);
nand U15532 (N_15532,N_15328,N_15286);
xnor U15533 (N_15533,N_15296,N_15217);
xnor U15534 (N_15534,N_15372,N_15350);
nand U15535 (N_15535,N_15397,N_15366);
nand U15536 (N_15536,N_15317,N_15265);
nand U15537 (N_15537,N_15304,N_15317);
or U15538 (N_15538,N_15216,N_15377);
nand U15539 (N_15539,N_15398,N_15360);
nor U15540 (N_15540,N_15367,N_15244);
nor U15541 (N_15541,N_15351,N_15305);
or U15542 (N_15542,N_15212,N_15319);
or U15543 (N_15543,N_15299,N_15246);
or U15544 (N_15544,N_15317,N_15372);
or U15545 (N_15545,N_15242,N_15363);
and U15546 (N_15546,N_15270,N_15256);
nor U15547 (N_15547,N_15337,N_15354);
or U15548 (N_15548,N_15363,N_15345);
xor U15549 (N_15549,N_15296,N_15383);
and U15550 (N_15550,N_15242,N_15376);
and U15551 (N_15551,N_15395,N_15259);
nand U15552 (N_15552,N_15246,N_15315);
and U15553 (N_15553,N_15235,N_15289);
nor U15554 (N_15554,N_15254,N_15309);
nor U15555 (N_15555,N_15330,N_15221);
nor U15556 (N_15556,N_15324,N_15371);
or U15557 (N_15557,N_15200,N_15316);
nand U15558 (N_15558,N_15287,N_15249);
or U15559 (N_15559,N_15356,N_15378);
or U15560 (N_15560,N_15367,N_15356);
nand U15561 (N_15561,N_15234,N_15371);
nor U15562 (N_15562,N_15386,N_15345);
nor U15563 (N_15563,N_15320,N_15275);
or U15564 (N_15564,N_15233,N_15284);
nor U15565 (N_15565,N_15257,N_15363);
and U15566 (N_15566,N_15347,N_15293);
nand U15567 (N_15567,N_15375,N_15392);
or U15568 (N_15568,N_15355,N_15380);
nand U15569 (N_15569,N_15324,N_15346);
nor U15570 (N_15570,N_15370,N_15300);
and U15571 (N_15571,N_15236,N_15350);
or U15572 (N_15572,N_15290,N_15316);
nand U15573 (N_15573,N_15230,N_15212);
nor U15574 (N_15574,N_15398,N_15349);
and U15575 (N_15575,N_15362,N_15350);
and U15576 (N_15576,N_15387,N_15304);
nand U15577 (N_15577,N_15244,N_15299);
nor U15578 (N_15578,N_15339,N_15203);
nor U15579 (N_15579,N_15288,N_15311);
nor U15580 (N_15580,N_15232,N_15384);
and U15581 (N_15581,N_15301,N_15233);
nand U15582 (N_15582,N_15323,N_15383);
nand U15583 (N_15583,N_15379,N_15257);
or U15584 (N_15584,N_15349,N_15246);
nand U15585 (N_15585,N_15230,N_15288);
nand U15586 (N_15586,N_15204,N_15276);
and U15587 (N_15587,N_15220,N_15384);
and U15588 (N_15588,N_15314,N_15287);
nand U15589 (N_15589,N_15373,N_15242);
and U15590 (N_15590,N_15247,N_15350);
nor U15591 (N_15591,N_15381,N_15232);
and U15592 (N_15592,N_15207,N_15299);
nand U15593 (N_15593,N_15266,N_15202);
nor U15594 (N_15594,N_15319,N_15234);
nor U15595 (N_15595,N_15383,N_15382);
and U15596 (N_15596,N_15276,N_15273);
or U15597 (N_15597,N_15258,N_15313);
nor U15598 (N_15598,N_15234,N_15280);
nor U15599 (N_15599,N_15365,N_15223);
nand U15600 (N_15600,N_15508,N_15518);
nor U15601 (N_15601,N_15534,N_15567);
nand U15602 (N_15602,N_15452,N_15459);
nor U15603 (N_15603,N_15410,N_15494);
nand U15604 (N_15604,N_15476,N_15573);
and U15605 (N_15605,N_15524,N_15414);
and U15606 (N_15606,N_15598,N_15539);
and U15607 (N_15607,N_15544,N_15487);
or U15608 (N_15608,N_15563,N_15477);
and U15609 (N_15609,N_15596,N_15435);
and U15610 (N_15610,N_15504,N_15427);
or U15611 (N_15611,N_15403,N_15515);
or U15612 (N_15612,N_15446,N_15506);
nand U15613 (N_15613,N_15569,N_15555);
and U15614 (N_15614,N_15480,N_15583);
or U15615 (N_15615,N_15439,N_15431);
and U15616 (N_15616,N_15428,N_15526);
and U15617 (N_15617,N_15478,N_15517);
or U15618 (N_15618,N_15562,N_15547);
xnor U15619 (N_15619,N_15599,N_15455);
and U15620 (N_15620,N_15527,N_15406);
nand U15621 (N_15621,N_15484,N_15570);
or U15622 (N_15622,N_15579,N_15499);
or U15623 (N_15623,N_15482,N_15591);
nand U15624 (N_15624,N_15580,N_15442);
or U15625 (N_15625,N_15528,N_15516);
nor U15626 (N_15626,N_15525,N_15537);
and U15627 (N_15627,N_15419,N_15460);
and U15628 (N_15628,N_15404,N_15535);
nand U15629 (N_15629,N_15514,N_15566);
nor U15630 (N_15630,N_15469,N_15492);
or U15631 (N_15631,N_15443,N_15522);
nor U15632 (N_15632,N_15401,N_15481);
nor U15633 (N_15633,N_15429,N_15521);
or U15634 (N_15634,N_15557,N_15572);
nor U15635 (N_15635,N_15584,N_15491);
or U15636 (N_15636,N_15493,N_15432);
and U15637 (N_15637,N_15543,N_15479);
nor U15638 (N_15638,N_15447,N_15502);
nor U15639 (N_15639,N_15457,N_15507);
or U15640 (N_15640,N_15418,N_15445);
nand U15641 (N_15641,N_15430,N_15560);
or U15642 (N_15642,N_15454,N_15588);
or U15643 (N_15643,N_15467,N_15451);
nor U15644 (N_15644,N_15510,N_15400);
nand U15645 (N_15645,N_15495,N_15587);
nor U15646 (N_15646,N_15595,N_15470);
nand U15647 (N_15647,N_15564,N_15578);
nand U15648 (N_15648,N_15464,N_15474);
or U15649 (N_15649,N_15412,N_15423);
and U15650 (N_15650,N_15444,N_15574);
and U15651 (N_15651,N_15590,N_15512);
or U15652 (N_15652,N_15458,N_15505);
and U15653 (N_15653,N_15550,N_15558);
nor U15654 (N_15654,N_15441,N_15576);
nor U15655 (N_15655,N_15413,N_15422);
nand U15656 (N_15656,N_15548,N_15575);
and U15657 (N_15657,N_15501,N_15577);
nand U15658 (N_15658,N_15471,N_15436);
nor U15659 (N_15659,N_15483,N_15540);
and U15660 (N_15660,N_15497,N_15533);
nor U15661 (N_15661,N_15503,N_15453);
or U15662 (N_15662,N_15490,N_15589);
or U15663 (N_15663,N_15408,N_15592);
nand U15664 (N_15664,N_15415,N_15417);
nand U15665 (N_15665,N_15586,N_15498);
nand U15666 (N_15666,N_15568,N_15475);
nand U15667 (N_15667,N_15559,N_15473);
and U15668 (N_15668,N_15461,N_15538);
and U15669 (N_15669,N_15437,N_15565);
and U15670 (N_15670,N_15407,N_15489);
nor U15671 (N_15671,N_15530,N_15511);
and U15672 (N_15672,N_15440,N_15509);
or U15673 (N_15673,N_15409,N_15472);
and U15674 (N_15674,N_15425,N_15531);
nand U15675 (N_15675,N_15546,N_15554);
nand U15676 (N_15676,N_15552,N_15593);
nor U15677 (N_15677,N_15496,N_15434);
nand U15678 (N_15678,N_15532,N_15465);
and U15679 (N_15679,N_15597,N_15416);
or U15680 (N_15680,N_15405,N_15536);
nor U15681 (N_15681,N_15545,N_15488);
nand U15682 (N_15682,N_15449,N_15411);
nor U15683 (N_15683,N_15561,N_15520);
nor U15684 (N_15684,N_15585,N_15581);
nand U15685 (N_15685,N_15513,N_15463);
nor U15686 (N_15686,N_15549,N_15450);
nand U15687 (N_15687,N_15402,N_15556);
or U15688 (N_15688,N_15594,N_15542);
and U15689 (N_15689,N_15529,N_15553);
and U15690 (N_15690,N_15468,N_15485);
or U15691 (N_15691,N_15519,N_15438);
nand U15692 (N_15692,N_15541,N_15448);
or U15693 (N_15693,N_15456,N_15500);
and U15694 (N_15694,N_15523,N_15582);
nor U15695 (N_15695,N_15426,N_15571);
and U15696 (N_15696,N_15486,N_15466);
or U15697 (N_15697,N_15462,N_15433);
nand U15698 (N_15698,N_15424,N_15421);
nand U15699 (N_15699,N_15551,N_15420);
nand U15700 (N_15700,N_15560,N_15482);
nor U15701 (N_15701,N_15545,N_15421);
nand U15702 (N_15702,N_15510,N_15539);
nand U15703 (N_15703,N_15520,N_15518);
or U15704 (N_15704,N_15470,N_15465);
nand U15705 (N_15705,N_15566,N_15462);
nor U15706 (N_15706,N_15534,N_15578);
and U15707 (N_15707,N_15584,N_15540);
and U15708 (N_15708,N_15460,N_15546);
and U15709 (N_15709,N_15403,N_15449);
and U15710 (N_15710,N_15447,N_15409);
and U15711 (N_15711,N_15436,N_15567);
nand U15712 (N_15712,N_15426,N_15596);
or U15713 (N_15713,N_15475,N_15518);
or U15714 (N_15714,N_15428,N_15521);
and U15715 (N_15715,N_15408,N_15427);
nand U15716 (N_15716,N_15516,N_15400);
nor U15717 (N_15717,N_15596,N_15424);
and U15718 (N_15718,N_15478,N_15560);
nand U15719 (N_15719,N_15427,N_15462);
and U15720 (N_15720,N_15459,N_15589);
and U15721 (N_15721,N_15596,N_15403);
or U15722 (N_15722,N_15516,N_15584);
nor U15723 (N_15723,N_15573,N_15449);
and U15724 (N_15724,N_15550,N_15504);
and U15725 (N_15725,N_15526,N_15573);
or U15726 (N_15726,N_15469,N_15535);
nand U15727 (N_15727,N_15508,N_15436);
or U15728 (N_15728,N_15545,N_15406);
and U15729 (N_15729,N_15564,N_15537);
and U15730 (N_15730,N_15426,N_15545);
nand U15731 (N_15731,N_15520,N_15440);
xor U15732 (N_15732,N_15449,N_15559);
or U15733 (N_15733,N_15441,N_15426);
nor U15734 (N_15734,N_15403,N_15538);
nor U15735 (N_15735,N_15563,N_15462);
or U15736 (N_15736,N_15454,N_15532);
nand U15737 (N_15737,N_15455,N_15401);
nor U15738 (N_15738,N_15529,N_15416);
or U15739 (N_15739,N_15427,N_15489);
and U15740 (N_15740,N_15435,N_15511);
nor U15741 (N_15741,N_15421,N_15416);
nor U15742 (N_15742,N_15449,N_15514);
nor U15743 (N_15743,N_15480,N_15516);
and U15744 (N_15744,N_15492,N_15480);
and U15745 (N_15745,N_15418,N_15464);
nor U15746 (N_15746,N_15443,N_15428);
or U15747 (N_15747,N_15402,N_15541);
or U15748 (N_15748,N_15510,N_15556);
or U15749 (N_15749,N_15470,N_15582);
and U15750 (N_15750,N_15483,N_15440);
nand U15751 (N_15751,N_15477,N_15590);
nor U15752 (N_15752,N_15415,N_15577);
nand U15753 (N_15753,N_15513,N_15450);
nor U15754 (N_15754,N_15578,N_15565);
nand U15755 (N_15755,N_15526,N_15543);
nor U15756 (N_15756,N_15441,N_15532);
nor U15757 (N_15757,N_15450,N_15453);
and U15758 (N_15758,N_15494,N_15527);
nand U15759 (N_15759,N_15470,N_15539);
or U15760 (N_15760,N_15504,N_15566);
or U15761 (N_15761,N_15566,N_15487);
nand U15762 (N_15762,N_15471,N_15561);
or U15763 (N_15763,N_15507,N_15500);
or U15764 (N_15764,N_15557,N_15504);
and U15765 (N_15765,N_15477,N_15408);
nand U15766 (N_15766,N_15447,N_15497);
nand U15767 (N_15767,N_15491,N_15481);
nand U15768 (N_15768,N_15405,N_15533);
and U15769 (N_15769,N_15431,N_15421);
or U15770 (N_15770,N_15473,N_15505);
nor U15771 (N_15771,N_15460,N_15542);
or U15772 (N_15772,N_15492,N_15500);
nor U15773 (N_15773,N_15467,N_15537);
and U15774 (N_15774,N_15508,N_15468);
nand U15775 (N_15775,N_15495,N_15514);
nor U15776 (N_15776,N_15505,N_15578);
nor U15777 (N_15777,N_15410,N_15567);
or U15778 (N_15778,N_15438,N_15479);
nand U15779 (N_15779,N_15489,N_15498);
and U15780 (N_15780,N_15447,N_15462);
and U15781 (N_15781,N_15414,N_15519);
nor U15782 (N_15782,N_15533,N_15429);
and U15783 (N_15783,N_15546,N_15444);
and U15784 (N_15784,N_15527,N_15462);
nand U15785 (N_15785,N_15427,N_15573);
nand U15786 (N_15786,N_15468,N_15578);
nand U15787 (N_15787,N_15485,N_15508);
and U15788 (N_15788,N_15550,N_15411);
or U15789 (N_15789,N_15528,N_15465);
and U15790 (N_15790,N_15442,N_15490);
or U15791 (N_15791,N_15438,N_15458);
nor U15792 (N_15792,N_15459,N_15569);
nand U15793 (N_15793,N_15512,N_15511);
nor U15794 (N_15794,N_15424,N_15442);
nand U15795 (N_15795,N_15552,N_15586);
and U15796 (N_15796,N_15408,N_15548);
nand U15797 (N_15797,N_15490,N_15569);
nand U15798 (N_15798,N_15500,N_15490);
and U15799 (N_15799,N_15415,N_15544);
nand U15800 (N_15800,N_15653,N_15756);
or U15801 (N_15801,N_15650,N_15665);
nor U15802 (N_15802,N_15615,N_15656);
or U15803 (N_15803,N_15683,N_15686);
nand U15804 (N_15804,N_15667,N_15761);
nor U15805 (N_15805,N_15716,N_15658);
or U15806 (N_15806,N_15773,N_15793);
nand U15807 (N_15807,N_15721,N_15700);
nand U15808 (N_15808,N_15742,N_15642);
nor U15809 (N_15809,N_15647,N_15673);
or U15810 (N_15810,N_15774,N_15736);
or U15811 (N_15811,N_15798,N_15677);
nor U15812 (N_15812,N_15726,N_15762);
and U15813 (N_15813,N_15661,N_15747);
nand U15814 (N_15814,N_15685,N_15625);
and U15815 (N_15815,N_15708,N_15606);
nand U15816 (N_15816,N_15733,N_15776);
or U15817 (N_15817,N_15679,N_15754);
nand U15818 (N_15818,N_15792,N_15639);
nor U15819 (N_15819,N_15724,N_15796);
nor U15820 (N_15820,N_15640,N_15714);
or U15821 (N_15821,N_15669,N_15668);
nor U15822 (N_15822,N_15770,N_15623);
and U15823 (N_15823,N_15725,N_15713);
and U15824 (N_15824,N_15689,N_15600);
nand U15825 (N_15825,N_15672,N_15707);
nand U15826 (N_15826,N_15791,N_15630);
nand U15827 (N_15827,N_15655,N_15618);
nor U15828 (N_15828,N_15750,N_15624);
nor U15829 (N_15829,N_15780,N_15727);
nand U15830 (N_15830,N_15779,N_15757);
or U15831 (N_15831,N_15735,N_15734);
nor U15832 (N_15832,N_15751,N_15701);
and U15833 (N_15833,N_15691,N_15633);
or U15834 (N_15834,N_15752,N_15641);
nor U15835 (N_15835,N_15765,N_15654);
nand U15836 (N_15836,N_15741,N_15755);
and U15837 (N_15837,N_15728,N_15787);
nor U15838 (N_15838,N_15737,N_15645);
or U15839 (N_15839,N_15788,N_15766);
and U15840 (N_15840,N_15695,N_15619);
nand U15841 (N_15841,N_15722,N_15769);
or U15842 (N_15842,N_15730,N_15610);
nor U15843 (N_15843,N_15767,N_15732);
nand U15844 (N_15844,N_15664,N_15768);
nor U15845 (N_15845,N_15602,N_15682);
or U15846 (N_15846,N_15617,N_15785);
and U15847 (N_15847,N_15745,N_15703);
nor U15848 (N_15848,N_15782,N_15616);
nor U15849 (N_15849,N_15760,N_15651);
nand U15850 (N_15850,N_15620,N_15764);
nand U15851 (N_15851,N_15704,N_15636);
and U15852 (N_15852,N_15797,N_15626);
and U15853 (N_15853,N_15676,N_15772);
nand U15854 (N_15854,N_15646,N_15711);
nor U15855 (N_15855,N_15740,N_15698);
nand U15856 (N_15856,N_15697,N_15675);
and U15857 (N_15857,N_15758,N_15778);
nand U15858 (N_15858,N_15709,N_15671);
nand U15859 (N_15859,N_15660,N_15688);
and U15860 (N_15860,N_15608,N_15729);
and U15861 (N_15861,N_15603,N_15693);
nand U15862 (N_15862,N_15723,N_15643);
and U15863 (N_15863,N_15621,N_15712);
nand U15864 (N_15864,N_15702,N_15657);
and U15865 (N_15865,N_15648,N_15696);
and U15866 (N_15866,N_15666,N_15635);
and U15867 (N_15867,N_15759,N_15634);
xnor U15868 (N_15868,N_15720,N_15605);
or U15869 (N_15869,N_15629,N_15710);
nor U15870 (N_15870,N_15789,N_15637);
or U15871 (N_15871,N_15662,N_15799);
nand U15872 (N_15872,N_15631,N_15719);
nor U15873 (N_15873,N_15748,N_15622);
or U15874 (N_15874,N_15699,N_15738);
nor U15875 (N_15875,N_15684,N_15649);
and U15876 (N_15876,N_15690,N_15790);
or U15877 (N_15877,N_15692,N_15680);
nor U15878 (N_15878,N_15784,N_15628);
nand U15879 (N_15879,N_15638,N_15674);
nand U15880 (N_15880,N_15609,N_15687);
nand U15881 (N_15881,N_15775,N_15607);
nand U15882 (N_15882,N_15795,N_15771);
nand U15883 (N_15883,N_15627,N_15794);
and U15884 (N_15884,N_15753,N_15763);
or U15885 (N_15885,N_15611,N_15749);
nand U15886 (N_15886,N_15718,N_15670);
nor U15887 (N_15887,N_15681,N_15744);
nor U15888 (N_15888,N_15652,N_15632);
nand U15889 (N_15889,N_15659,N_15613);
and U15890 (N_15890,N_15601,N_15783);
nor U15891 (N_15891,N_15746,N_15663);
and U15892 (N_15892,N_15786,N_15781);
nand U15893 (N_15893,N_15612,N_15604);
and U15894 (N_15894,N_15706,N_15705);
and U15895 (N_15895,N_15777,N_15678);
nand U15896 (N_15896,N_15614,N_15694);
or U15897 (N_15897,N_15739,N_15717);
nand U15898 (N_15898,N_15743,N_15644);
or U15899 (N_15899,N_15731,N_15715);
nor U15900 (N_15900,N_15773,N_15637);
or U15901 (N_15901,N_15737,N_15665);
nand U15902 (N_15902,N_15723,N_15759);
or U15903 (N_15903,N_15724,N_15653);
or U15904 (N_15904,N_15701,N_15617);
and U15905 (N_15905,N_15779,N_15638);
nand U15906 (N_15906,N_15677,N_15639);
nand U15907 (N_15907,N_15774,N_15685);
nor U15908 (N_15908,N_15763,N_15696);
and U15909 (N_15909,N_15707,N_15769);
or U15910 (N_15910,N_15787,N_15674);
nand U15911 (N_15911,N_15709,N_15724);
nor U15912 (N_15912,N_15782,N_15632);
nor U15913 (N_15913,N_15692,N_15670);
and U15914 (N_15914,N_15652,N_15646);
nand U15915 (N_15915,N_15694,N_15663);
nor U15916 (N_15916,N_15639,N_15775);
or U15917 (N_15917,N_15703,N_15676);
and U15918 (N_15918,N_15745,N_15642);
nor U15919 (N_15919,N_15738,N_15697);
nand U15920 (N_15920,N_15612,N_15716);
and U15921 (N_15921,N_15699,N_15677);
nand U15922 (N_15922,N_15602,N_15612);
nand U15923 (N_15923,N_15781,N_15761);
nand U15924 (N_15924,N_15718,N_15773);
nor U15925 (N_15925,N_15703,N_15750);
and U15926 (N_15926,N_15730,N_15655);
nand U15927 (N_15927,N_15759,N_15649);
nand U15928 (N_15928,N_15752,N_15757);
nor U15929 (N_15929,N_15611,N_15772);
or U15930 (N_15930,N_15766,N_15769);
and U15931 (N_15931,N_15794,N_15616);
nand U15932 (N_15932,N_15601,N_15662);
nand U15933 (N_15933,N_15648,N_15612);
nand U15934 (N_15934,N_15720,N_15647);
and U15935 (N_15935,N_15672,N_15741);
or U15936 (N_15936,N_15666,N_15619);
nand U15937 (N_15937,N_15753,N_15671);
nor U15938 (N_15938,N_15751,N_15666);
nand U15939 (N_15939,N_15617,N_15682);
or U15940 (N_15940,N_15738,N_15677);
nand U15941 (N_15941,N_15602,N_15712);
nor U15942 (N_15942,N_15695,N_15757);
nand U15943 (N_15943,N_15640,N_15604);
nor U15944 (N_15944,N_15625,N_15724);
and U15945 (N_15945,N_15762,N_15722);
nor U15946 (N_15946,N_15619,N_15686);
and U15947 (N_15947,N_15680,N_15785);
and U15948 (N_15948,N_15748,N_15743);
and U15949 (N_15949,N_15603,N_15742);
nor U15950 (N_15950,N_15600,N_15756);
or U15951 (N_15951,N_15735,N_15635);
and U15952 (N_15952,N_15615,N_15691);
nand U15953 (N_15953,N_15773,N_15762);
nand U15954 (N_15954,N_15699,N_15602);
nand U15955 (N_15955,N_15726,N_15670);
xor U15956 (N_15956,N_15763,N_15679);
nor U15957 (N_15957,N_15718,N_15680);
nor U15958 (N_15958,N_15680,N_15621);
nor U15959 (N_15959,N_15678,N_15701);
or U15960 (N_15960,N_15674,N_15605);
nor U15961 (N_15961,N_15733,N_15706);
and U15962 (N_15962,N_15674,N_15640);
and U15963 (N_15963,N_15797,N_15716);
and U15964 (N_15964,N_15743,N_15668);
nor U15965 (N_15965,N_15731,N_15712);
nor U15966 (N_15966,N_15733,N_15688);
or U15967 (N_15967,N_15768,N_15609);
nor U15968 (N_15968,N_15685,N_15730);
or U15969 (N_15969,N_15604,N_15677);
or U15970 (N_15970,N_15605,N_15682);
or U15971 (N_15971,N_15773,N_15698);
nand U15972 (N_15972,N_15687,N_15742);
nor U15973 (N_15973,N_15651,N_15675);
nor U15974 (N_15974,N_15685,N_15670);
nand U15975 (N_15975,N_15659,N_15610);
and U15976 (N_15976,N_15740,N_15665);
and U15977 (N_15977,N_15609,N_15645);
or U15978 (N_15978,N_15795,N_15601);
and U15979 (N_15979,N_15795,N_15633);
and U15980 (N_15980,N_15654,N_15667);
or U15981 (N_15981,N_15711,N_15621);
or U15982 (N_15982,N_15673,N_15619);
nor U15983 (N_15983,N_15791,N_15793);
nor U15984 (N_15984,N_15756,N_15649);
nand U15985 (N_15985,N_15794,N_15786);
or U15986 (N_15986,N_15702,N_15644);
and U15987 (N_15987,N_15656,N_15710);
nand U15988 (N_15988,N_15684,N_15791);
and U15989 (N_15989,N_15614,N_15729);
nand U15990 (N_15990,N_15677,N_15731);
nand U15991 (N_15991,N_15722,N_15691);
nand U15992 (N_15992,N_15647,N_15773);
or U15993 (N_15993,N_15645,N_15736);
or U15994 (N_15994,N_15648,N_15695);
or U15995 (N_15995,N_15649,N_15656);
or U15996 (N_15996,N_15793,N_15639);
and U15997 (N_15997,N_15794,N_15651);
nor U15998 (N_15998,N_15646,N_15797);
or U15999 (N_15999,N_15675,N_15737);
and U16000 (N_16000,N_15931,N_15806);
or U16001 (N_16001,N_15983,N_15938);
nand U16002 (N_16002,N_15945,N_15903);
or U16003 (N_16003,N_15844,N_15875);
and U16004 (N_16004,N_15829,N_15987);
nand U16005 (N_16005,N_15973,N_15962);
nand U16006 (N_16006,N_15879,N_15892);
nand U16007 (N_16007,N_15848,N_15957);
nor U16008 (N_16008,N_15940,N_15923);
nand U16009 (N_16009,N_15807,N_15873);
and U16010 (N_16010,N_15910,N_15905);
and U16011 (N_16011,N_15835,N_15937);
nor U16012 (N_16012,N_15907,N_15929);
nand U16013 (N_16013,N_15820,N_15958);
nor U16014 (N_16014,N_15954,N_15979);
nor U16015 (N_16015,N_15819,N_15846);
nor U16016 (N_16016,N_15856,N_15857);
or U16017 (N_16017,N_15864,N_15843);
nor U16018 (N_16018,N_15964,N_15992);
or U16019 (N_16019,N_15827,N_15939);
or U16020 (N_16020,N_15975,N_15996);
nor U16021 (N_16021,N_15961,N_15935);
and U16022 (N_16022,N_15988,N_15909);
or U16023 (N_16023,N_15853,N_15831);
nor U16024 (N_16024,N_15825,N_15915);
nor U16025 (N_16025,N_15816,N_15981);
nand U16026 (N_16026,N_15860,N_15952);
nand U16027 (N_16027,N_15978,N_15883);
or U16028 (N_16028,N_15881,N_15956);
or U16029 (N_16029,N_15814,N_15951);
xnor U16030 (N_16030,N_15895,N_15890);
nor U16031 (N_16031,N_15885,N_15876);
nand U16032 (N_16032,N_15891,N_15801);
or U16033 (N_16033,N_15994,N_15934);
or U16034 (N_16034,N_15805,N_15901);
nand U16035 (N_16035,N_15986,N_15972);
or U16036 (N_16036,N_15974,N_15838);
or U16037 (N_16037,N_15911,N_15989);
xnor U16038 (N_16038,N_15818,N_15899);
and U16039 (N_16039,N_15809,N_15865);
nand U16040 (N_16040,N_15916,N_15925);
nand U16041 (N_16041,N_15904,N_15894);
nand U16042 (N_16042,N_15977,N_15993);
and U16043 (N_16043,N_15963,N_15863);
and U16044 (N_16044,N_15948,N_15833);
or U16045 (N_16045,N_15810,N_15870);
and U16046 (N_16046,N_15811,N_15800);
and U16047 (N_16047,N_15824,N_15847);
nand U16048 (N_16048,N_15884,N_15817);
nor U16049 (N_16049,N_15917,N_15998);
nor U16050 (N_16050,N_15913,N_15893);
or U16051 (N_16051,N_15867,N_15868);
or U16052 (N_16052,N_15880,N_15947);
nand U16053 (N_16053,N_15997,N_15866);
nor U16054 (N_16054,N_15837,N_15918);
or U16055 (N_16055,N_15821,N_15849);
nand U16056 (N_16056,N_15926,N_15971);
or U16057 (N_16057,N_15841,N_15840);
nor U16058 (N_16058,N_15855,N_15830);
nand U16059 (N_16059,N_15812,N_15960);
or U16060 (N_16060,N_15914,N_15928);
nand U16061 (N_16061,N_15808,N_15887);
and U16062 (N_16062,N_15984,N_15967);
nand U16063 (N_16063,N_15955,N_15976);
and U16064 (N_16064,N_15861,N_15927);
or U16065 (N_16065,N_15919,N_15858);
or U16066 (N_16066,N_15980,N_15999);
nand U16067 (N_16067,N_15839,N_15902);
xor U16068 (N_16068,N_15932,N_15906);
nor U16069 (N_16069,N_15965,N_15850);
nor U16070 (N_16070,N_15985,N_15822);
or U16071 (N_16071,N_15990,N_15968);
nor U16072 (N_16072,N_15804,N_15908);
nand U16073 (N_16073,N_15836,N_15953);
xor U16074 (N_16074,N_15828,N_15871);
nor U16075 (N_16075,N_15852,N_15920);
or U16076 (N_16076,N_15941,N_15851);
nand U16077 (N_16077,N_15886,N_15949);
or U16078 (N_16078,N_15930,N_15942);
nand U16079 (N_16079,N_15882,N_15813);
nand U16080 (N_16080,N_15802,N_15888);
and U16081 (N_16081,N_15991,N_15936);
or U16082 (N_16082,N_15877,N_15922);
and U16083 (N_16083,N_15900,N_15872);
nand U16084 (N_16084,N_15950,N_15874);
and U16085 (N_16085,N_15921,N_15842);
nor U16086 (N_16086,N_15859,N_15878);
and U16087 (N_16087,N_15982,N_15823);
nor U16088 (N_16088,N_15912,N_15943);
nand U16089 (N_16089,N_15970,N_15889);
or U16090 (N_16090,N_15869,N_15832);
nor U16091 (N_16091,N_15946,N_15966);
and U16092 (N_16092,N_15898,N_15896);
and U16093 (N_16093,N_15897,N_15924);
nor U16094 (N_16094,N_15959,N_15803);
and U16095 (N_16095,N_15969,N_15815);
or U16096 (N_16096,N_15995,N_15834);
nor U16097 (N_16097,N_15845,N_15862);
nor U16098 (N_16098,N_15933,N_15944);
or U16099 (N_16099,N_15826,N_15854);
or U16100 (N_16100,N_15991,N_15885);
nand U16101 (N_16101,N_15934,N_15885);
and U16102 (N_16102,N_15976,N_15993);
and U16103 (N_16103,N_15924,N_15809);
and U16104 (N_16104,N_15991,N_15838);
and U16105 (N_16105,N_15929,N_15994);
nand U16106 (N_16106,N_15809,N_15914);
nor U16107 (N_16107,N_15970,N_15996);
or U16108 (N_16108,N_15808,N_15883);
or U16109 (N_16109,N_15928,N_15811);
or U16110 (N_16110,N_15992,N_15971);
nor U16111 (N_16111,N_15824,N_15881);
nand U16112 (N_16112,N_15966,N_15933);
nor U16113 (N_16113,N_15865,N_15813);
or U16114 (N_16114,N_15944,N_15998);
xnor U16115 (N_16115,N_15955,N_15866);
nor U16116 (N_16116,N_15872,N_15978);
and U16117 (N_16117,N_15993,N_15937);
nor U16118 (N_16118,N_15924,N_15907);
nor U16119 (N_16119,N_15952,N_15810);
nand U16120 (N_16120,N_15870,N_15886);
or U16121 (N_16121,N_15842,N_15998);
nor U16122 (N_16122,N_15873,N_15972);
and U16123 (N_16123,N_15892,N_15933);
nor U16124 (N_16124,N_15898,N_15992);
nand U16125 (N_16125,N_15887,N_15844);
and U16126 (N_16126,N_15957,N_15852);
nor U16127 (N_16127,N_15871,N_15847);
or U16128 (N_16128,N_15815,N_15807);
and U16129 (N_16129,N_15837,N_15946);
or U16130 (N_16130,N_15907,N_15886);
nand U16131 (N_16131,N_15822,N_15888);
and U16132 (N_16132,N_15946,N_15952);
and U16133 (N_16133,N_15822,N_15849);
or U16134 (N_16134,N_15978,N_15939);
or U16135 (N_16135,N_15866,N_15867);
and U16136 (N_16136,N_15823,N_15812);
nor U16137 (N_16137,N_15954,N_15816);
nor U16138 (N_16138,N_15893,N_15844);
or U16139 (N_16139,N_15814,N_15944);
nor U16140 (N_16140,N_15960,N_15928);
or U16141 (N_16141,N_15889,N_15929);
nand U16142 (N_16142,N_15963,N_15939);
or U16143 (N_16143,N_15842,N_15852);
and U16144 (N_16144,N_15840,N_15864);
and U16145 (N_16145,N_15822,N_15987);
nor U16146 (N_16146,N_15942,N_15818);
or U16147 (N_16147,N_15845,N_15959);
nor U16148 (N_16148,N_15963,N_15979);
or U16149 (N_16149,N_15918,N_15903);
nor U16150 (N_16150,N_15981,N_15997);
xor U16151 (N_16151,N_15906,N_15911);
nand U16152 (N_16152,N_15810,N_15964);
nor U16153 (N_16153,N_15849,N_15833);
nor U16154 (N_16154,N_15916,N_15893);
or U16155 (N_16155,N_15862,N_15898);
or U16156 (N_16156,N_15953,N_15958);
or U16157 (N_16157,N_15893,N_15928);
nand U16158 (N_16158,N_15929,N_15862);
and U16159 (N_16159,N_15910,N_15813);
nand U16160 (N_16160,N_15864,N_15807);
or U16161 (N_16161,N_15971,N_15804);
nor U16162 (N_16162,N_15940,N_15992);
or U16163 (N_16163,N_15923,N_15995);
nor U16164 (N_16164,N_15830,N_15951);
and U16165 (N_16165,N_15830,N_15967);
nand U16166 (N_16166,N_15970,N_15831);
and U16167 (N_16167,N_15871,N_15820);
and U16168 (N_16168,N_15871,N_15998);
or U16169 (N_16169,N_15815,N_15983);
and U16170 (N_16170,N_15952,N_15908);
nand U16171 (N_16171,N_15947,N_15969);
nand U16172 (N_16172,N_15965,N_15996);
nand U16173 (N_16173,N_15925,N_15819);
and U16174 (N_16174,N_15941,N_15943);
nor U16175 (N_16175,N_15805,N_15835);
and U16176 (N_16176,N_15823,N_15910);
nand U16177 (N_16177,N_15886,N_15871);
nand U16178 (N_16178,N_15967,N_15960);
and U16179 (N_16179,N_15940,N_15854);
nor U16180 (N_16180,N_15904,N_15901);
and U16181 (N_16181,N_15905,N_15975);
nand U16182 (N_16182,N_15941,N_15995);
nand U16183 (N_16183,N_15908,N_15849);
and U16184 (N_16184,N_15948,N_15839);
nand U16185 (N_16185,N_15822,N_15978);
and U16186 (N_16186,N_15883,N_15999);
nand U16187 (N_16187,N_15967,N_15895);
or U16188 (N_16188,N_15923,N_15820);
and U16189 (N_16189,N_15868,N_15908);
or U16190 (N_16190,N_15993,N_15830);
and U16191 (N_16191,N_15967,N_15808);
or U16192 (N_16192,N_15820,N_15858);
nor U16193 (N_16193,N_15903,N_15828);
nor U16194 (N_16194,N_15887,N_15954);
nor U16195 (N_16195,N_15908,N_15968);
nor U16196 (N_16196,N_15803,N_15987);
or U16197 (N_16197,N_15972,N_15831);
and U16198 (N_16198,N_15879,N_15861);
nor U16199 (N_16199,N_15866,N_15974);
nand U16200 (N_16200,N_16042,N_16136);
nor U16201 (N_16201,N_16160,N_16152);
and U16202 (N_16202,N_16101,N_16054);
nand U16203 (N_16203,N_16058,N_16045);
or U16204 (N_16204,N_16081,N_16142);
nor U16205 (N_16205,N_16121,N_16009);
nor U16206 (N_16206,N_16004,N_16082);
or U16207 (N_16207,N_16112,N_16105);
nand U16208 (N_16208,N_16055,N_16083);
or U16209 (N_16209,N_16175,N_16090);
nor U16210 (N_16210,N_16040,N_16176);
nor U16211 (N_16211,N_16046,N_16130);
and U16212 (N_16212,N_16149,N_16100);
nand U16213 (N_16213,N_16150,N_16030);
nand U16214 (N_16214,N_16056,N_16106);
nand U16215 (N_16215,N_16018,N_16148);
and U16216 (N_16216,N_16051,N_16166);
and U16217 (N_16217,N_16041,N_16174);
and U16218 (N_16218,N_16008,N_16049);
nor U16219 (N_16219,N_16027,N_16158);
or U16220 (N_16220,N_16162,N_16195);
nand U16221 (N_16221,N_16170,N_16111);
nand U16222 (N_16222,N_16062,N_16085);
and U16223 (N_16223,N_16086,N_16137);
and U16224 (N_16224,N_16124,N_16145);
and U16225 (N_16225,N_16188,N_16161);
nand U16226 (N_16226,N_16013,N_16193);
nor U16227 (N_16227,N_16017,N_16061);
and U16228 (N_16228,N_16139,N_16169);
or U16229 (N_16229,N_16173,N_16116);
or U16230 (N_16230,N_16095,N_16065);
and U16231 (N_16231,N_16118,N_16198);
or U16232 (N_16232,N_16001,N_16068);
and U16233 (N_16233,N_16037,N_16057);
nor U16234 (N_16234,N_16167,N_16135);
and U16235 (N_16235,N_16067,N_16184);
or U16236 (N_16236,N_16172,N_16075);
nand U16237 (N_16237,N_16134,N_16102);
and U16238 (N_16238,N_16031,N_16153);
or U16239 (N_16239,N_16122,N_16197);
and U16240 (N_16240,N_16036,N_16157);
or U16241 (N_16241,N_16039,N_16129);
nand U16242 (N_16242,N_16154,N_16127);
and U16243 (N_16243,N_16147,N_16094);
nor U16244 (N_16244,N_16138,N_16131);
or U16245 (N_16245,N_16074,N_16053);
and U16246 (N_16246,N_16171,N_16003);
nand U16247 (N_16247,N_16126,N_16113);
and U16248 (N_16248,N_16144,N_16132);
or U16249 (N_16249,N_16115,N_16016);
nor U16250 (N_16250,N_16010,N_16070);
nor U16251 (N_16251,N_16024,N_16038);
or U16252 (N_16252,N_16097,N_16151);
or U16253 (N_16253,N_16181,N_16014);
or U16254 (N_16254,N_16191,N_16063);
nand U16255 (N_16255,N_16103,N_16064);
nor U16256 (N_16256,N_16078,N_16059);
nand U16257 (N_16257,N_16091,N_16023);
nand U16258 (N_16258,N_16159,N_16060);
or U16259 (N_16259,N_16178,N_16156);
and U16260 (N_16260,N_16026,N_16096);
nor U16261 (N_16261,N_16079,N_16050);
nor U16262 (N_16262,N_16072,N_16012);
nor U16263 (N_16263,N_16199,N_16044);
and U16264 (N_16264,N_16114,N_16125);
and U16265 (N_16265,N_16019,N_16155);
or U16266 (N_16266,N_16011,N_16034);
nand U16267 (N_16267,N_16133,N_16183);
nand U16268 (N_16268,N_16092,N_16164);
nand U16269 (N_16269,N_16120,N_16189);
nand U16270 (N_16270,N_16005,N_16179);
and U16271 (N_16271,N_16032,N_16168);
nor U16272 (N_16272,N_16033,N_16071);
and U16273 (N_16273,N_16021,N_16002);
nor U16274 (N_16274,N_16022,N_16006);
and U16275 (N_16275,N_16007,N_16165);
nor U16276 (N_16276,N_16104,N_16029);
nor U16277 (N_16277,N_16087,N_16047);
and U16278 (N_16278,N_16107,N_16196);
nor U16279 (N_16279,N_16192,N_16093);
nand U16280 (N_16280,N_16089,N_16025);
nand U16281 (N_16281,N_16119,N_16110);
or U16282 (N_16282,N_16194,N_16146);
nand U16283 (N_16283,N_16088,N_16000);
nand U16284 (N_16284,N_16066,N_16084);
or U16285 (N_16285,N_16141,N_16069);
nand U16286 (N_16286,N_16052,N_16163);
and U16287 (N_16287,N_16140,N_16128);
or U16288 (N_16288,N_16015,N_16077);
nor U16289 (N_16289,N_16076,N_16190);
or U16290 (N_16290,N_16186,N_16028);
and U16291 (N_16291,N_16182,N_16187);
nor U16292 (N_16292,N_16185,N_16143);
nand U16293 (N_16293,N_16073,N_16035);
nand U16294 (N_16294,N_16108,N_16099);
or U16295 (N_16295,N_16123,N_16180);
nand U16296 (N_16296,N_16177,N_16043);
nor U16297 (N_16297,N_16109,N_16048);
nor U16298 (N_16298,N_16020,N_16080);
and U16299 (N_16299,N_16117,N_16098);
nor U16300 (N_16300,N_16162,N_16163);
nand U16301 (N_16301,N_16066,N_16105);
and U16302 (N_16302,N_16053,N_16037);
nand U16303 (N_16303,N_16108,N_16058);
or U16304 (N_16304,N_16119,N_16041);
and U16305 (N_16305,N_16152,N_16108);
nand U16306 (N_16306,N_16150,N_16018);
and U16307 (N_16307,N_16192,N_16146);
nor U16308 (N_16308,N_16095,N_16084);
and U16309 (N_16309,N_16147,N_16118);
or U16310 (N_16310,N_16028,N_16121);
nor U16311 (N_16311,N_16121,N_16010);
and U16312 (N_16312,N_16085,N_16107);
or U16313 (N_16313,N_16188,N_16197);
or U16314 (N_16314,N_16112,N_16140);
nor U16315 (N_16315,N_16195,N_16194);
or U16316 (N_16316,N_16113,N_16112);
or U16317 (N_16317,N_16186,N_16150);
and U16318 (N_16318,N_16071,N_16094);
and U16319 (N_16319,N_16181,N_16035);
or U16320 (N_16320,N_16035,N_16142);
and U16321 (N_16321,N_16083,N_16064);
nand U16322 (N_16322,N_16171,N_16032);
nor U16323 (N_16323,N_16071,N_16198);
nand U16324 (N_16324,N_16078,N_16126);
nand U16325 (N_16325,N_16151,N_16022);
nand U16326 (N_16326,N_16049,N_16160);
nand U16327 (N_16327,N_16148,N_16145);
and U16328 (N_16328,N_16056,N_16169);
nor U16329 (N_16329,N_16040,N_16036);
nor U16330 (N_16330,N_16081,N_16065);
nor U16331 (N_16331,N_16043,N_16026);
nor U16332 (N_16332,N_16088,N_16061);
or U16333 (N_16333,N_16029,N_16149);
nor U16334 (N_16334,N_16169,N_16147);
nand U16335 (N_16335,N_16143,N_16179);
or U16336 (N_16336,N_16180,N_16107);
or U16337 (N_16337,N_16075,N_16057);
nand U16338 (N_16338,N_16054,N_16114);
or U16339 (N_16339,N_16199,N_16174);
or U16340 (N_16340,N_16163,N_16141);
nor U16341 (N_16341,N_16043,N_16075);
nand U16342 (N_16342,N_16033,N_16041);
or U16343 (N_16343,N_16056,N_16142);
nor U16344 (N_16344,N_16004,N_16003);
or U16345 (N_16345,N_16040,N_16183);
nor U16346 (N_16346,N_16050,N_16075);
and U16347 (N_16347,N_16115,N_16093);
and U16348 (N_16348,N_16147,N_16194);
and U16349 (N_16349,N_16076,N_16019);
or U16350 (N_16350,N_16184,N_16043);
or U16351 (N_16351,N_16062,N_16009);
nor U16352 (N_16352,N_16031,N_16119);
nand U16353 (N_16353,N_16126,N_16171);
and U16354 (N_16354,N_16054,N_16088);
nand U16355 (N_16355,N_16100,N_16135);
nor U16356 (N_16356,N_16162,N_16107);
and U16357 (N_16357,N_16066,N_16167);
or U16358 (N_16358,N_16181,N_16007);
or U16359 (N_16359,N_16125,N_16193);
nand U16360 (N_16360,N_16187,N_16014);
or U16361 (N_16361,N_16196,N_16080);
or U16362 (N_16362,N_16136,N_16186);
and U16363 (N_16363,N_16182,N_16057);
nand U16364 (N_16364,N_16009,N_16013);
or U16365 (N_16365,N_16112,N_16147);
nand U16366 (N_16366,N_16102,N_16009);
nor U16367 (N_16367,N_16165,N_16107);
and U16368 (N_16368,N_16083,N_16060);
or U16369 (N_16369,N_16189,N_16165);
nand U16370 (N_16370,N_16032,N_16122);
and U16371 (N_16371,N_16044,N_16173);
nand U16372 (N_16372,N_16055,N_16030);
or U16373 (N_16373,N_16163,N_16041);
or U16374 (N_16374,N_16101,N_16195);
nor U16375 (N_16375,N_16174,N_16067);
nor U16376 (N_16376,N_16166,N_16145);
nor U16377 (N_16377,N_16104,N_16048);
or U16378 (N_16378,N_16031,N_16051);
nor U16379 (N_16379,N_16153,N_16017);
or U16380 (N_16380,N_16080,N_16031);
or U16381 (N_16381,N_16181,N_16045);
or U16382 (N_16382,N_16057,N_16022);
or U16383 (N_16383,N_16078,N_16088);
or U16384 (N_16384,N_16041,N_16012);
nor U16385 (N_16385,N_16075,N_16136);
nand U16386 (N_16386,N_16104,N_16062);
or U16387 (N_16387,N_16156,N_16177);
and U16388 (N_16388,N_16072,N_16078);
nor U16389 (N_16389,N_16187,N_16017);
nand U16390 (N_16390,N_16140,N_16081);
or U16391 (N_16391,N_16065,N_16018);
and U16392 (N_16392,N_16110,N_16109);
and U16393 (N_16393,N_16064,N_16144);
and U16394 (N_16394,N_16061,N_16009);
nand U16395 (N_16395,N_16035,N_16164);
nor U16396 (N_16396,N_16199,N_16080);
nand U16397 (N_16397,N_16139,N_16087);
and U16398 (N_16398,N_16128,N_16188);
nor U16399 (N_16399,N_16113,N_16143);
nand U16400 (N_16400,N_16307,N_16333);
nand U16401 (N_16401,N_16314,N_16399);
and U16402 (N_16402,N_16335,N_16386);
or U16403 (N_16403,N_16354,N_16304);
nand U16404 (N_16404,N_16311,N_16325);
nand U16405 (N_16405,N_16316,N_16371);
and U16406 (N_16406,N_16204,N_16249);
nor U16407 (N_16407,N_16360,N_16381);
nand U16408 (N_16408,N_16280,N_16298);
and U16409 (N_16409,N_16357,N_16268);
and U16410 (N_16410,N_16284,N_16374);
nor U16411 (N_16411,N_16341,N_16200);
or U16412 (N_16412,N_16344,N_16369);
or U16413 (N_16413,N_16237,N_16397);
nor U16414 (N_16414,N_16309,N_16342);
nor U16415 (N_16415,N_16212,N_16283);
nand U16416 (N_16416,N_16323,N_16225);
nor U16417 (N_16417,N_16390,N_16279);
nor U16418 (N_16418,N_16391,N_16294);
nand U16419 (N_16419,N_16208,N_16286);
nand U16420 (N_16420,N_16243,N_16329);
nand U16421 (N_16421,N_16278,N_16332);
nor U16422 (N_16422,N_16241,N_16218);
or U16423 (N_16423,N_16376,N_16264);
nand U16424 (N_16424,N_16231,N_16326);
or U16425 (N_16425,N_16258,N_16306);
and U16426 (N_16426,N_16217,N_16203);
or U16427 (N_16427,N_16205,N_16343);
nor U16428 (N_16428,N_16246,N_16312);
nand U16429 (N_16429,N_16269,N_16229);
and U16430 (N_16430,N_16260,N_16221);
or U16431 (N_16431,N_16387,N_16349);
or U16432 (N_16432,N_16257,N_16255);
nand U16433 (N_16433,N_16261,N_16202);
and U16434 (N_16434,N_16305,N_16353);
or U16435 (N_16435,N_16345,N_16364);
or U16436 (N_16436,N_16248,N_16293);
or U16437 (N_16437,N_16336,N_16396);
nand U16438 (N_16438,N_16380,N_16285);
nor U16439 (N_16439,N_16273,N_16289);
nand U16440 (N_16440,N_16313,N_16373);
and U16441 (N_16441,N_16334,N_16253);
or U16442 (N_16442,N_16230,N_16377);
nor U16443 (N_16443,N_16211,N_16247);
nand U16444 (N_16444,N_16275,N_16240);
or U16445 (N_16445,N_16219,N_16395);
and U16446 (N_16446,N_16352,N_16392);
or U16447 (N_16447,N_16365,N_16256);
or U16448 (N_16448,N_16213,N_16393);
and U16449 (N_16449,N_16251,N_16301);
nor U16450 (N_16450,N_16224,N_16287);
and U16451 (N_16451,N_16389,N_16348);
or U16452 (N_16452,N_16226,N_16362);
and U16453 (N_16453,N_16295,N_16347);
nand U16454 (N_16454,N_16252,N_16288);
and U16455 (N_16455,N_16321,N_16356);
nand U16456 (N_16456,N_16245,N_16337);
nor U16457 (N_16457,N_16207,N_16359);
or U16458 (N_16458,N_16398,N_16274);
nand U16459 (N_16459,N_16265,N_16378);
nor U16460 (N_16460,N_16201,N_16222);
nand U16461 (N_16461,N_16367,N_16216);
nor U16462 (N_16462,N_16228,N_16238);
nand U16463 (N_16463,N_16319,N_16262);
nand U16464 (N_16464,N_16234,N_16322);
or U16465 (N_16465,N_16340,N_16368);
and U16466 (N_16466,N_16384,N_16233);
or U16467 (N_16467,N_16351,N_16303);
and U16468 (N_16468,N_16382,N_16244);
or U16469 (N_16469,N_16206,N_16267);
and U16470 (N_16470,N_16297,N_16259);
and U16471 (N_16471,N_16254,N_16282);
nor U16472 (N_16472,N_16308,N_16232);
nor U16473 (N_16473,N_16361,N_16350);
and U16474 (N_16474,N_16339,N_16320);
nor U16475 (N_16475,N_16214,N_16263);
nor U16476 (N_16476,N_16366,N_16331);
nand U16477 (N_16477,N_16292,N_16394);
or U16478 (N_16478,N_16223,N_16266);
or U16479 (N_16479,N_16355,N_16235);
nand U16480 (N_16480,N_16310,N_16338);
and U16481 (N_16481,N_16272,N_16327);
or U16482 (N_16482,N_16358,N_16239);
nor U16483 (N_16483,N_16281,N_16302);
and U16484 (N_16484,N_16363,N_16271);
nand U16485 (N_16485,N_16215,N_16276);
and U16486 (N_16486,N_16270,N_16210);
nand U16487 (N_16487,N_16370,N_16388);
or U16488 (N_16488,N_16236,N_16346);
nand U16489 (N_16489,N_16330,N_16209);
and U16490 (N_16490,N_16300,N_16385);
and U16491 (N_16491,N_16324,N_16296);
nand U16492 (N_16492,N_16242,N_16379);
nor U16493 (N_16493,N_16317,N_16375);
and U16494 (N_16494,N_16291,N_16372);
nor U16495 (N_16495,N_16250,N_16227);
nand U16496 (N_16496,N_16318,N_16383);
nand U16497 (N_16497,N_16277,N_16328);
nor U16498 (N_16498,N_16220,N_16315);
nor U16499 (N_16499,N_16299,N_16290);
or U16500 (N_16500,N_16209,N_16267);
nor U16501 (N_16501,N_16234,N_16373);
and U16502 (N_16502,N_16375,N_16357);
nand U16503 (N_16503,N_16227,N_16390);
nand U16504 (N_16504,N_16240,N_16230);
nand U16505 (N_16505,N_16214,N_16348);
and U16506 (N_16506,N_16239,N_16342);
or U16507 (N_16507,N_16361,N_16349);
nand U16508 (N_16508,N_16330,N_16394);
nand U16509 (N_16509,N_16381,N_16227);
or U16510 (N_16510,N_16390,N_16253);
nor U16511 (N_16511,N_16340,N_16256);
nand U16512 (N_16512,N_16323,N_16240);
nand U16513 (N_16513,N_16341,N_16279);
and U16514 (N_16514,N_16350,N_16278);
nor U16515 (N_16515,N_16285,N_16375);
nor U16516 (N_16516,N_16335,N_16292);
or U16517 (N_16517,N_16390,N_16357);
nor U16518 (N_16518,N_16281,N_16278);
nand U16519 (N_16519,N_16314,N_16254);
and U16520 (N_16520,N_16243,N_16207);
nand U16521 (N_16521,N_16334,N_16306);
or U16522 (N_16522,N_16215,N_16399);
nor U16523 (N_16523,N_16306,N_16224);
nor U16524 (N_16524,N_16394,N_16273);
or U16525 (N_16525,N_16290,N_16259);
nor U16526 (N_16526,N_16323,N_16264);
nor U16527 (N_16527,N_16271,N_16305);
nor U16528 (N_16528,N_16349,N_16386);
nor U16529 (N_16529,N_16373,N_16222);
nand U16530 (N_16530,N_16393,N_16365);
or U16531 (N_16531,N_16362,N_16388);
or U16532 (N_16532,N_16348,N_16355);
or U16533 (N_16533,N_16276,N_16208);
or U16534 (N_16534,N_16368,N_16392);
and U16535 (N_16535,N_16235,N_16372);
and U16536 (N_16536,N_16309,N_16200);
nand U16537 (N_16537,N_16335,N_16341);
nand U16538 (N_16538,N_16296,N_16362);
nand U16539 (N_16539,N_16369,N_16340);
and U16540 (N_16540,N_16230,N_16396);
or U16541 (N_16541,N_16278,N_16306);
nor U16542 (N_16542,N_16323,N_16205);
nand U16543 (N_16543,N_16308,N_16305);
and U16544 (N_16544,N_16248,N_16391);
or U16545 (N_16545,N_16309,N_16219);
or U16546 (N_16546,N_16252,N_16228);
nand U16547 (N_16547,N_16326,N_16209);
and U16548 (N_16548,N_16261,N_16370);
nand U16549 (N_16549,N_16282,N_16242);
nor U16550 (N_16550,N_16209,N_16286);
and U16551 (N_16551,N_16337,N_16393);
and U16552 (N_16552,N_16251,N_16329);
nor U16553 (N_16553,N_16265,N_16272);
or U16554 (N_16554,N_16348,N_16263);
nor U16555 (N_16555,N_16335,N_16307);
and U16556 (N_16556,N_16348,N_16333);
and U16557 (N_16557,N_16203,N_16216);
or U16558 (N_16558,N_16268,N_16337);
or U16559 (N_16559,N_16239,N_16397);
or U16560 (N_16560,N_16362,N_16243);
xnor U16561 (N_16561,N_16273,N_16340);
or U16562 (N_16562,N_16219,N_16373);
or U16563 (N_16563,N_16306,N_16303);
or U16564 (N_16564,N_16375,N_16251);
and U16565 (N_16565,N_16394,N_16247);
and U16566 (N_16566,N_16292,N_16313);
nor U16567 (N_16567,N_16350,N_16374);
or U16568 (N_16568,N_16213,N_16214);
nand U16569 (N_16569,N_16377,N_16252);
or U16570 (N_16570,N_16396,N_16374);
and U16571 (N_16571,N_16265,N_16271);
nand U16572 (N_16572,N_16387,N_16383);
nor U16573 (N_16573,N_16316,N_16266);
nor U16574 (N_16574,N_16273,N_16333);
nor U16575 (N_16575,N_16216,N_16329);
nand U16576 (N_16576,N_16286,N_16389);
or U16577 (N_16577,N_16274,N_16339);
nand U16578 (N_16578,N_16301,N_16247);
nor U16579 (N_16579,N_16273,N_16297);
nor U16580 (N_16580,N_16284,N_16323);
nand U16581 (N_16581,N_16355,N_16309);
or U16582 (N_16582,N_16317,N_16209);
nor U16583 (N_16583,N_16319,N_16304);
and U16584 (N_16584,N_16389,N_16254);
nand U16585 (N_16585,N_16353,N_16359);
or U16586 (N_16586,N_16202,N_16200);
nor U16587 (N_16587,N_16318,N_16214);
or U16588 (N_16588,N_16307,N_16390);
nand U16589 (N_16589,N_16397,N_16316);
and U16590 (N_16590,N_16256,N_16381);
nor U16591 (N_16591,N_16209,N_16307);
and U16592 (N_16592,N_16277,N_16373);
and U16593 (N_16593,N_16360,N_16375);
nand U16594 (N_16594,N_16341,N_16390);
nor U16595 (N_16595,N_16374,N_16204);
or U16596 (N_16596,N_16263,N_16301);
nor U16597 (N_16597,N_16306,N_16383);
and U16598 (N_16598,N_16364,N_16396);
and U16599 (N_16599,N_16345,N_16397);
nor U16600 (N_16600,N_16577,N_16462);
or U16601 (N_16601,N_16435,N_16421);
nor U16602 (N_16602,N_16575,N_16452);
and U16603 (N_16603,N_16484,N_16445);
nor U16604 (N_16604,N_16409,N_16524);
nand U16605 (N_16605,N_16415,N_16589);
and U16606 (N_16606,N_16581,N_16533);
nand U16607 (N_16607,N_16429,N_16478);
nand U16608 (N_16608,N_16460,N_16471);
and U16609 (N_16609,N_16441,N_16586);
or U16610 (N_16610,N_16416,N_16528);
nand U16611 (N_16611,N_16578,N_16582);
nor U16612 (N_16612,N_16483,N_16593);
or U16613 (N_16613,N_16555,N_16564);
nor U16614 (N_16614,N_16514,N_16463);
and U16615 (N_16615,N_16442,N_16494);
nor U16616 (N_16616,N_16572,N_16591);
nor U16617 (N_16617,N_16438,N_16482);
nand U16618 (N_16618,N_16449,N_16481);
nor U16619 (N_16619,N_16426,N_16502);
or U16620 (N_16620,N_16579,N_16504);
nor U16621 (N_16621,N_16541,N_16527);
and U16622 (N_16622,N_16427,N_16477);
nor U16623 (N_16623,N_16574,N_16436);
and U16624 (N_16624,N_16414,N_16457);
nand U16625 (N_16625,N_16570,N_16490);
nor U16626 (N_16626,N_16497,N_16598);
or U16627 (N_16627,N_16443,N_16444);
nor U16628 (N_16628,N_16525,N_16402);
or U16629 (N_16629,N_16454,N_16515);
nor U16630 (N_16630,N_16534,N_16539);
or U16631 (N_16631,N_16401,N_16506);
or U16632 (N_16632,N_16508,N_16537);
nor U16633 (N_16633,N_16465,N_16556);
and U16634 (N_16634,N_16561,N_16447);
nand U16635 (N_16635,N_16542,N_16458);
and U16636 (N_16636,N_16407,N_16571);
nand U16637 (N_16637,N_16476,N_16473);
nand U16638 (N_16638,N_16585,N_16526);
or U16639 (N_16639,N_16400,N_16428);
or U16640 (N_16640,N_16479,N_16432);
and U16641 (N_16641,N_16594,N_16520);
or U16642 (N_16642,N_16470,N_16487);
nand U16643 (N_16643,N_16425,N_16544);
or U16644 (N_16644,N_16545,N_16511);
nor U16645 (N_16645,N_16560,N_16540);
or U16646 (N_16646,N_16472,N_16433);
or U16647 (N_16647,N_16538,N_16567);
or U16648 (N_16648,N_16559,N_16453);
or U16649 (N_16649,N_16410,N_16486);
and U16650 (N_16650,N_16553,N_16512);
and U16651 (N_16651,N_16569,N_16501);
or U16652 (N_16652,N_16547,N_16568);
and U16653 (N_16653,N_16562,N_16498);
and U16654 (N_16654,N_16576,N_16451);
or U16655 (N_16655,N_16565,N_16434);
or U16656 (N_16656,N_16408,N_16509);
nor U16657 (N_16657,N_16440,N_16584);
nand U16658 (N_16658,N_16522,N_16422);
nand U16659 (N_16659,N_16588,N_16491);
or U16660 (N_16660,N_16455,N_16456);
or U16661 (N_16661,N_16531,N_16423);
nor U16662 (N_16662,N_16595,N_16543);
nand U16663 (N_16663,N_16437,N_16554);
and U16664 (N_16664,N_16590,N_16505);
nand U16665 (N_16665,N_16495,N_16446);
nand U16666 (N_16666,N_16566,N_16475);
and U16667 (N_16667,N_16469,N_16510);
nand U16668 (N_16668,N_16563,N_16466);
nor U16669 (N_16669,N_16523,N_16496);
and U16670 (N_16670,N_16503,N_16485);
or U16671 (N_16671,N_16558,N_16499);
and U16672 (N_16672,N_16596,N_16599);
nor U16673 (N_16673,N_16489,N_16551);
and U16674 (N_16674,N_16439,N_16532);
and U16675 (N_16675,N_16430,N_16530);
and U16676 (N_16676,N_16403,N_16405);
or U16677 (N_16677,N_16557,N_16474);
nand U16678 (N_16678,N_16536,N_16420);
or U16679 (N_16679,N_16500,N_16431);
nand U16680 (N_16680,N_16406,N_16552);
nand U16681 (N_16681,N_16518,N_16464);
or U16682 (N_16682,N_16467,N_16424);
nand U16683 (N_16683,N_16448,N_16535);
nand U16684 (N_16684,N_16516,N_16492);
or U16685 (N_16685,N_16468,N_16597);
nand U16686 (N_16686,N_16419,N_16548);
and U16687 (N_16687,N_16413,N_16450);
or U16688 (N_16688,N_16546,N_16417);
and U16689 (N_16689,N_16513,N_16521);
or U16690 (N_16690,N_16587,N_16550);
and U16691 (N_16691,N_16412,N_16507);
or U16692 (N_16692,N_16461,N_16592);
nand U16693 (N_16693,N_16519,N_16549);
or U16694 (N_16694,N_16573,N_16480);
or U16695 (N_16695,N_16411,N_16418);
nor U16696 (N_16696,N_16529,N_16580);
and U16697 (N_16697,N_16583,N_16517);
nor U16698 (N_16698,N_16488,N_16404);
and U16699 (N_16699,N_16493,N_16459);
nand U16700 (N_16700,N_16525,N_16505);
or U16701 (N_16701,N_16585,N_16520);
or U16702 (N_16702,N_16458,N_16575);
nand U16703 (N_16703,N_16430,N_16462);
nand U16704 (N_16704,N_16418,N_16436);
nand U16705 (N_16705,N_16412,N_16561);
and U16706 (N_16706,N_16487,N_16446);
or U16707 (N_16707,N_16507,N_16409);
nand U16708 (N_16708,N_16563,N_16556);
nand U16709 (N_16709,N_16408,N_16581);
nor U16710 (N_16710,N_16561,N_16584);
nor U16711 (N_16711,N_16464,N_16447);
and U16712 (N_16712,N_16555,N_16488);
nand U16713 (N_16713,N_16437,N_16560);
and U16714 (N_16714,N_16479,N_16480);
and U16715 (N_16715,N_16559,N_16417);
and U16716 (N_16716,N_16499,N_16579);
nor U16717 (N_16717,N_16581,N_16551);
nand U16718 (N_16718,N_16482,N_16401);
nand U16719 (N_16719,N_16445,N_16548);
nor U16720 (N_16720,N_16458,N_16530);
nor U16721 (N_16721,N_16541,N_16560);
or U16722 (N_16722,N_16429,N_16565);
nand U16723 (N_16723,N_16563,N_16463);
nor U16724 (N_16724,N_16480,N_16587);
nor U16725 (N_16725,N_16492,N_16574);
nor U16726 (N_16726,N_16501,N_16446);
nor U16727 (N_16727,N_16538,N_16506);
and U16728 (N_16728,N_16582,N_16463);
nor U16729 (N_16729,N_16525,N_16457);
nor U16730 (N_16730,N_16420,N_16438);
or U16731 (N_16731,N_16539,N_16414);
or U16732 (N_16732,N_16510,N_16541);
nor U16733 (N_16733,N_16490,N_16522);
nand U16734 (N_16734,N_16414,N_16468);
and U16735 (N_16735,N_16503,N_16444);
or U16736 (N_16736,N_16491,N_16407);
nand U16737 (N_16737,N_16477,N_16452);
nand U16738 (N_16738,N_16435,N_16439);
nor U16739 (N_16739,N_16510,N_16489);
nor U16740 (N_16740,N_16536,N_16418);
or U16741 (N_16741,N_16452,N_16552);
or U16742 (N_16742,N_16541,N_16561);
and U16743 (N_16743,N_16434,N_16542);
or U16744 (N_16744,N_16434,N_16570);
or U16745 (N_16745,N_16450,N_16404);
nand U16746 (N_16746,N_16421,N_16491);
or U16747 (N_16747,N_16555,N_16585);
nand U16748 (N_16748,N_16416,N_16455);
or U16749 (N_16749,N_16593,N_16468);
nand U16750 (N_16750,N_16404,N_16451);
xor U16751 (N_16751,N_16467,N_16481);
nand U16752 (N_16752,N_16460,N_16574);
nor U16753 (N_16753,N_16575,N_16410);
nand U16754 (N_16754,N_16546,N_16563);
or U16755 (N_16755,N_16455,N_16433);
nand U16756 (N_16756,N_16475,N_16565);
or U16757 (N_16757,N_16472,N_16596);
and U16758 (N_16758,N_16434,N_16474);
and U16759 (N_16759,N_16577,N_16470);
or U16760 (N_16760,N_16488,N_16431);
nor U16761 (N_16761,N_16416,N_16579);
nand U16762 (N_16762,N_16439,N_16557);
and U16763 (N_16763,N_16589,N_16587);
nand U16764 (N_16764,N_16485,N_16452);
or U16765 (N_16765,N_16563,N_16441);
nor U16766 (N_16766,N_16599,N_16564);
and U16767 (N_16767,N_16518,N_16506);
xnor U16768 (N_16768,N_16402,N_16412);
and U16769 (N_16769,N_16410,N_16501);
nor U16770 (N_16770,N_16496,N_16511);
nor U16771 (N_16771,N_16404,N_16516);
nand U16772 (N_16772,N_16582,N_16516);
nand U16773 (N_16773,N_16596,N_16436);
nor U16774 (N_16774,N_16470,N_16483);
and U16775 (N_16775,N_16466,N_16458);
nor U16776 (N_16776,N_16559,N_16420);
or U16777 (N_16777,N_16573,N_16481);
nand U16778 (N_16778,N_16463,N_16478);
and U16779 (N_16779,N_16489,N_16473);
and U16780 (N_16780,N_16437,N_16579);
and U16781 (N_16781,N_16591,N_16586);
nand U16782 (N_16782,N_16572,N_16571);
nor U16783 (N_16783,N_16417,N_16420);
nor U16784 (N_16784,N_16537,N_16460);
and U16785 (N_16785,N_16465,N_16461);
nand U16786 (N_16786,N_16501,N_16469);
and U16787 (N_16787,N_16522,N_16478);
and U16788 (N_16788,N_16564,N_16561);
nand U16789 (N_16789,N_16572,N_16550);
nor U16790 (N_16790,N_16408,N_16587);
nand U16791 (N_16791,N_16514,N_16544);
and U16792 (N_16792,N_16505,N_16510);
nor U16793 (N_16793,N_16498,N_16470);
nand U16794 (N_16794,N_16507,N_16425);
nor U16795 (N_16795,N_16447,N_16493);
and U16796 (N_16796,N_16499,N_16555);
or U16797 (N_16797,N_16464,N_16511);
and U16798 (N_16798,N_16425,N_16599);
or U16799 (N_16799,N_16578,N_16420);
nor U16800 (N_16800,N_16643,N_16605);
nor U16801 (N_16801,N_16739,N_16762);
and U16802 (N_16802,N_16781,N_16716);
nand U16803 (N_16803,N_16797,N_16774);
and U16804 (N_16804,N_16743,N_16661);
and U16805 (N_16805,N_16744,N_16657);
nand U16806 (N_16806,N_16734,N_16690);
xnor U16807 (N_16807,N_16784,N_16705);
nand U16808 (N_16808,N_16709,N_16720);
nand U16809 (N_16809,N_16601,N_16652);
and U16810 (N_16810,N_16730,N_16752);
nand U16811 (N_16811,N_16741,N_16669);
xnor U16812 (N_16812,N_16722,N_16733);
nand U16813 (N_16813,N_16764,N_16653);
and U16814 (N_16814,N_16702,N_16768);
nor U16815 (N_16815,N_16607,N_16721);
and U16816 (N_16816,N_16685,N_16651);
nand U16817 (N_16817,N_16629,N_16732);
or U16818 (N_16818,N_16723,N_16632);
nor U16819 (N_16819,N_16694,N_16606);
nand U16820 (N_16820,N_16700,N_16623);
or U16821 (N_16821,N_16794,N_16790);
nand U16822 (N_16822,N_16742,N_16612);
and U16823 (N_16823,N_16628,N_16672);
or U16824 (N_16824,N_16780,N_16656);
nand U16825 (N_16825,N_16618,N_16688);
or U16826 (N_16826,N_16624,N_16736);
and U16827 (N_16827,N_16756,N_16675);
nand U16828 (N_16828,N_16738,N_16726);
or U16829 (N_16829,N_16799,N_16600);
or U16830 (N_16830,N_16769,N_16613);
nand U16831 (N_16831,N_16602,N_16636);
nand U16832 (N_16832,N_16758,N_16682);
nand U16833 (N_16833,N_16621,N_16697);
or U16834 (N_16834,N_16788,N_16637);
nor U16835 (N_16835,N_16753,N_16708);
nor U16836 (N_16836,N_16763,N_16670);
nand U16837 (N_16837,N_16660,N_16728);
and U16838 (N_16838,N_16667,N_16666);
nor U16839 (N_16839,N_16662,N_16619);
or U16840 (N_16840,N_16766,N_16631);
nand U16841 (N_16841,N_16692,N_16772);
nand U16842 (N_16842,N_16646,N_16689);
nand U16843 (N_16843,N_16683,N_16659);
or U16844 (N_16844,N_16668,N_16749);
nand U16845 (N_16845,N_16717,N_16777);
and U16846 (N_16846,N_16617,N_16699);
and U16847 (N_16847,N_16610,N_16796);
or U16848 (N_16848,N_16770,N_16746);
or U16849 (N_16849,N_16686,N_16663);
and U16850 (N_16850,N_16755,N_16696);
and U16851 (N_16851,N_16750,N_16775);
nand U16852 (N_16852,N_16782,N_16620);
or U16853 (N_16853,N_16776,N_16664);
nor U16854 (N_16854,N_16704,N_16603);
or U16855 (N_16855,N_16681,N_16707);
or U16856 (N_16856,N_16765,N_16614);
nor U16857 (N_16857,N_16634,N_16622);
nor U16858 (N_16858,N_16706,N_16633);
or U16859 (N_16859,N_16779,N_16648);
and U16860 (N_16860,N_16748,N_16626);
nand U16861 (N_16861,N_16655,N_16654);
nor U16862 (N_16862,N_16630,N_16644);
nand U16863 (N_16863,N_16674,N_16761);
or U16864 (N_16864,N_16650,N_16671);
and U16865 (N_16865,N_16785,N_16787);
and U16866 (N_16866,N_16731,N_16676);
and U16867 (N_16867,N_16791,N_16680);
and U16868 (N_16868,N_16604,N_16701);
nor U16869 (N_16869,N_16665,N_16798);
nand U16870 (N_16870,N_16608,N_16793);
and U16871 (N_16871,N_16737,N_16792);
nand U16872 (N_16872,N_16687,N_16754);
or U16873 (N_16873,N_16740,N_16645);
nor U16874 (N_16874,N_16635,N_16649);
nand U16875 (N_16875,N_16691,N_16751);
and U16876 (N_16876,N_16714,N_16638);
and U16877 (N_16877,N_16786,N_16625);
nor U16878 (N_16878,N_16759,N_16639);
or U16879 (N_16879,N_16725,N_16789);
nand U16880 (N_16880,N_16641,N_16693);
or U16881 (N_16881,N_16773,N_16647);
nand U16882 (N_16882,N_16609,N_16711);
nand U16883 (N_16883,N_16735,N_16713);
or U16884 (N_16884,N_16767,N_16684);
nand U16885 (N_16885,N_16710,N_16615);
nand U16886 (N_16886,N_16640,N_16783);
nand U16887 (N_16887,N_16715,N_16673);
or U16888 (N_16888,N_16771,N_16745);
nand U16889 (N_16889,N_16678,N_16795);
or U16890 (N_16890,N_16642,N_16727);
or U16891 (N_16891,N_16718,N_16747);
and U16892 (N_16892,N_16695,N_16616);
nand U16893 (N_16893,N_16757,N_16760);
nand U16894 (N_16894,N_16611,N_16729);
nand U16895 (N_16895,N_16627,N_16677);
and U16896 (N_16896,N_16719,N_16658);
nor U16897 (N_16897,N_16679,N_16724);
or U16898 (N_16898,N_16778,N_16698);
xor U16899 (N_16899,N_16703,N_16712);
nor U16900 (N_16900,N_16705,N_16688);
nand U16901 (N_16901,N_16621,N_16711);
and U16902 (N_16902,N_16716,N_16776);
or U16903 (N_16903,N_16618,N_16624);
or U16904 (N_16904,N_16612,N_16720);
and U16905 (N_16905,N_16623,N_16767);
and U16906 (N_16906,N_16694,N_16626);
and U16907 (N_16907,N_16649,N_16621);
nor U16908 (N_16908,N_16679,N_16763);
and U16909 (N_16909,N_16798,N_16651);
and U16910 (N_16910,N_16771,N_16712);
nor U16911 (N_16911,N_16669,N_16722);
and U16912 (N_16912,N_16775,N_16725);
and U16913 (N_16913,N_16780,N_16620);
or U16914 (N_16914,N_16662,N_16694);
nand U16915 (N_16915,N_16603,N_16751);
xor U16916 (N_16916,N_16686,N_16786);
or U16917 (N_16917,N_16677,N_16672);
or U16918 (N_16918,N_16685,N_16723);
nor U16919 (N_16919,N_16703,N_16791);
or U16920 (N_16920,N_16640,N_16799);
nand U16921 (N_16921,N_16730,N_16657);
and U16922 (N_16922,N_16772,N_16666);
nor U16923 (N_16923,N_16674,N_16738);
nor U16924 (N_16924,N_16786,N_16787);
and U16925 (N_16925,N_16716,N_16644);
and U16926 (N_16926,N_16788,N_16782);
nand U16927 (N_16927,N_16747,N_16720);
nand U16928 (N_16928,N_16708,N_16777);
nand U16929 (N_16929,N_16602,N_16695);
or U16930 (N_16930,N_16690,N_16674);
or U16931 (N_16931,N_16718,N_16720);
nor U16932 (N_16932,N_16693,N_16634);
or U16933 (N_16933,N_16685,N_16773);
and U16934 (N_16934,N_16693,N_16760);
and U16935 (N_16935,N_16643,N_16624);
and U16936 (N_16936,N_16629,N_16668);
nand U16937 (N_16937,N_16603,N_16765);
and U16938 (N_16938,N_16717,N_16687);
or U16939 (N_16939,N_16725,N_16652);
or U16940 (N_16940,N_16697,N_16639);
or U16941 (N_16941,N_16687,N_16758);
nor U16942 (N_16942,N_16746,N_16723);
nor U16943 (N_16943,N_16600,N_16689);
nor U16944 (N_16944,N_16741,N_16638);
nor U16945 (N_16945,N_16749,N_16793);
or U16946 (N_16946,N_16759,N_16761);
or U16947 (N_16947,N_16763,N_16650);
and U16948 (N_16948,N_16666,N_16682);
nor U16949 (N_16949,N_16758,N_16716);
or U16950 (N_16950,N_16661,N_16789);
nor U16951 (N_16951,N_16684,N_16646);
nand U16952 (N_16952,N_16742,N_16715);
nand U16953 (N_16953,N_16729,N_16608);
nor U16954 (N_16954,N_16775,N_16712);
nor U16955 (N_16955,N_16723,N_16652);
and U16956 (N_16956,N_16716,N_16735);
and U16957 (N_16957,N_16679,N_16615);
nor U16958 (N_16958,N_16731,N_16634);
or U16959 (N_16959,N_16725,N_16729);
nand U16960 (N_16960,N_16640,N_16681);
or U16961 (N_16961,N_16676,N_16695);
and U16962 (N_16962,N_16784,N_16726);
and U16963 (N_16963,N_16636,N_16764);
nand U16964 (N_16964,N_16603,N_16695);
nor U16965 (N_16965,N_16624,N_16666);
and U16966 (N_16966,N_16727,N_16627);
and U16967 (N_16967,N_16656,N_16689);
and U16968 (N_16968,N_16675,N_16717);
or U16969 (N_16969,N_16726,N_16670);
nand U16970 (N_16970,N_16669,N_16767);
nor U16971 (N_16971,N_16733,N_16720);
nand U16972 (N_16972,N_16739,N_16629);
nand U16973 (N_16973,N_16621,N_16743);
or U16974 (N_16974,N_16734,N_16663);
nor U16975 (N_16975,N_16633,N_16747);
nor U16976 (N_16976,N_16692,N_16664);
nor U16977 (N_16977,N_16631,N_16650);
and U16978 (N_16978,N_16617,N_16708);
or U16979 (N_16979,N_16738,N_16685);
and U16980 (N_16980,N_16730,N_16644);
nand U16981 (N_16981,N_16626,N_16633);
or U16982 (N_16982,N_16746,N_16797);
and U16983 (N_16983,N_16657,N_16679);
nor U16984 (N_16984,N_16796,N_16659);
nand U16985 (N_16985,N_16769,N_16733);
nor U16986 (N_16986,N_16782,N_16765);
nand U16987 (N_16987,N_16610,N_16625);
nand U16988 (N_16988,N_16786,N_16754);
or U16989 (N_16989,N_16745,N_16702);
nand U16990 (N_16990,N_16602,N_16672);
and U16991 (N_16991,N_16702,N_16708);
nor U16992 (N_16992,N_16618,N_16636);
nor U16993 (N_16993,N_16607,N_16673);
nand U16994 (N_16994,N_16630,N_16764);
or U16995 (N_16995,N_16793,N_16705);
nor U16996 (N_16996,N_16619,N_16648);
and U16997 (N_16997,N_16751,N_16724);
or U16998 (N_16998,N_16766,N_16739);
and U16999 (N_16999,N_16689,N_16714);
and U17000 (N_17000,N_16942,N_16855);
nor U17001 (N_17001,N_16843,N_16966);
or U17002 (N_17002,N_16852,N_16915);
nand U17003 (N_17003,N_16978,N_16943);
and U17004 (N_17004,N_16839,N_16933);
nor U17005 (N_17005,N_16880,N_16901);
or U17006 (N_17006,N_16895,N_16863);
nor U17007 (N_17007,N_16869,N_16914);
or U17008 (N_17008,N_16975,N_16964);
nor U17009 (N_17009,N_16916,N_16939);
and U17010 (N_17010,N_16889,N_16954);
and U17011 (N_17011,N_16849,N_16835);
xnor U17012 (N_17012,N_16924,N_16818);
and U17013 (N_17013,N_16807,N_16864);
or U17014 (N_17014,N_16833,N_16931);
and U17015 (N_17015,N_16859,N_16968);
or U17016 (N_17016,N_16947,N_16983);
nor U17017 (N_17017,N_16891,N_16845);
nand U17018 (N_17018,N_16999,N_16925);
and U17019 (N_17019,N_16866,N_16995);
nor U17020 (N_17020,N_16888,N_16912);
and U17021 (N_17021,N_16937,N_16971);
nand U17022 (N_17022,N_16827,N_16965);
nand U17023 (N_17023,N_16918,N_16879);
or U17024 (N_17024,N_16900,N_16950);
and U17025 (N_17025,N_16875,N_16962);
nor U17026 (N_17026,N_16809,N_16870);
nor U17027 (N_17027,N_16981,N_16885);
nor U17028 (N_17028,N_16936,N_16890);
nor U17029 (N_17029,N_16867,N_16928);
nand U17030 (N_17030,N_16957,N_16988);
nand U17031 (N_17031,N_16874,N_16823);
or U17032 (N_17032,N_16934,N_16961);
nor U17033 (N_17033,N_16882,N_16911);
nor U17034 (N_17034,N_16877,N_16932);
nor U17035 (N_17035,N_16920,N_16994);
nand U17036 (N_17036,N_16938,N_16850);
xor U17037 (N_17037,N_16853,N_16980);
nand U17038 (N_17038,N_16856,N_16930);
or U17039 (N_17039,N_16808,N_16829);
nor U17040 (N_17040,N_16814,N_16842);
nor U17041 (N_17041,N_16860,N_16910);
nand U17042 (N_17042,N_16972,N_16984);
or U17043 (N_17043,N_16926,N_16892);
nor U17044 (N_17044,N_16812,N_16871);
and U17045 (N_17045,N_16944,N_16830);
or U17046 (N_17046,N_16953,N_16949);
xnor U17047 (N_17047,N_16941,N_16876);
nand U17048 (N_17048,N_16990,N_16913);
nor U17049 (N_17049,N_16886,N_16973);
or U17050 (N_17050,N_16878,N_16997);
nor U17051 (N_17051,N_16907,N_16991);
nand U17052 (N_17052,N_16817,N_16834);
and U17053 (N_17053,N_16952,N_16987);
nor U17054 (N_17054,N_16861,N_16917);
and U17055 (N_17055,N_16946,N_16841);
nand U17056 (N_17056,N_16948,N_16893);
nand U17057 (N_17057,N_16803,N_16919);
nand U17058 (N_17058,N_16847,N_16846);
nand U17059 (N_17059,N_16896,N_16923);
nand U17060 (N_17060,N_16959,N_16970);
or U17061 (N_17061,N_16825,N_16862);
nor U17062 (N_17062,N_16935,N_16868);
and U17063 (N_17063,N_16824,N_16921);
or U17064 (N_17064,N_16821,N_16977);
nand U17065 (N_17065,N_16906,N_16940);
nor U17066 (N_17066,N_16887,N_16902);
and U17067 (N_17067,N_16967,N_16993);
nand U17068 (N_17068,N_16826,N_16884);
nand U17069 (N_17069,N_16806,N_16894);
or U17070 (N_17070,N_16989,N_16945);
and U17071 (N_17071,N_16810,N_16903);
nor U17072 (N_17072,N_16815,N_16831);
and U17073 (N_17073,N_16816,N_16801);
and U17074 (N_17074,N_16857,N_16828);
nor U17075 (N_17075,N_16905,N_16883);
nor U17076 (N_17076,N_16840,N_16813);
nand U17077 (N_17077,N_16820,N_16897);
and U17078 (N_17078,N_16960,N_16838);
and U17079 (N_17079,N_16844,N_16976);
nor U17080 (N_17080,N_16822,N_16929);
or U17081 (N_17081,N_16963,N_16805);
and U17082 (N_17082,N_16998,N_16985);
or U17083 (N_17083,N_16851,N_16819);
nand U17084 (N_17084,N_16872,N_16881);
or U17085 (N_17085,N_16837,N_16909);
nor U17086 (N_17086,N_16922,N_16865);
xnor U17087 (N_17087,N_16802,N_16858);
nand U17088 (N_17088,N_16986,N_16982);
and U17089 (N_17089,N_16804,N_16848);
or U17090 (N_17090,N_16873,N_16927);
nand U17091 (N_17091,N_16836,N_16992);
nand U17092 (N_17092,N_16904,N_16899);
or U17093 (N_17093,N_16979,N_16800);
or U17094 (N_17094,N_16951,N_16958);
or U17095 (N_17095,N_16956,N_16854);
and U17096 (N_17096,N_16969,N_16974);
nor U17097 (N_17097,N_16811,N_16908);
nand U17098 (N_17098,N_16898,N_16955);
and U17099 (N_17099,N_16996,N_16832);
or U17100 (N_17100,N_16804,N_16980);
or U17101 (N_17101,N_16957,N_16825);
nand U17102 (N_17102,N_16841,N_16979);
nand U17103 (N_17103,N_16886,N_16949);
nor U17104 (N_17104,N_16819,N_16907);
or U17105 (N_17105,N_16853,N_16934);
nor U17106 (N_17106,N_16877,N_16879);
and U17107 (N_17107,N_16913,N_16907);
and U17108 (N_17108,N_16999,N_16929);
and U17109 (N_17109,N_16961,N_16840);
nor U17110 (N_17110,N_16993,N_16998);
or U17111 (N_17111,N_16904,N_16934);
and U17112 (N_17112,N_16843,N_16972);
nand U17113 (N_17113,N_16992,N_16988);
and U17114 (N_17114,N_16928,N_16864);
or U17115 (N_17115,N_16899,N_16848);
or U17116 (N_17116,N_16905,N_16906);
or U17117 (N_17117,N_16979,N_16912);
or U17118 (N_17118,N_16903,N_16985);
or U17119 (N_17119,N_16872,N_16951);
nor U17120 (N_17120,N_16907,N_16800);
nand U17121 (N_17121,N_16955,N_16807);
nor U17122 (N_17122,N_16897,N_16921);
or U17123 (N_17123,N_16900,N_16850);
nor U17124 (N_17124,N_16897,N_16850);
nand U17125 (N_17125,N_16817,N_16973);
nand U17126 (N_17126,N_16966,N_16877);
and U17127 (N_17127,N_16841,N_16840);
nand U17128 (N_17128,N_16863,N_16801);
and U17129 (N_17129,N_16908,N_16844);
and U17130 (N_17130,N_16991,N_16950);
and U17131 (N_17131,N_16909,N_16934);
or U17132 (N_17132,N_16951,N_16824);
nor U17133 (N_17133,N_16986,N_16902);
nor U17134 (N_17134,N_16881,N_16938);
or U17135 (N_17135,N_16970,N_16890);
nor U17136 (N_17136,N_16893,N_16999);
xnor U17137 (N_17137,N_16909,N_16916);
nor U17138 (N_17138,N_16800,N_16881);
or U17139 (N_17139,N_16887,N_16848);
and U17140 (N_17140,N_16822,N_16828);
or U17141 (N_17141,N_16855,N_16847);
nor U17142 (N_17142,N_16805,N_16956);
or U17143 (N_17143,N_16865,N_16978);
nor U17144 (N_17144,N_16834,N_16894);
and U17145 (N_17145,N_16900,N_16824);
and U17146 (N_17146,N_16912,N_16841);
or U17147 (N_17147,N_16810,N_16809);
xnor U17148 (N_17148,N_16892,N_16976);
nor U17149 (N_17149,N_16967,N_16831);
or U17150 (N_17150,N_16950,N_16853);
and U17151 (N_17151,N_16819,N_16903);
nand U17152 (N_17152,N_16832,N_16856);
nand U17153 (N_17153,N_16970,N_16903);
nand U17154 (N_17154,N_16838,N_16986);
nand U17155 (N_17155,N_16947,N_16996);
or U17156 (N_17156,N_16865,N_16833);
nor U17157 (N_17157,N_16903,N_16920);
nor U17158 (N_17158,N_16928,N_16956);
nor U17159 (N_17159,N_16987,N_16849);
and U17160 (N_17160,N_16801,N_16805);
nand U17161 (N_17161,N_16829,N_16804);
nor U17162 (N_17162,N_16803,N_16863);
or U17163 (N_17163,N_16919,N_16926);
or U17164 (N_17164,N_16919,N_16833);
nor U17165 (N_17165,N_16894,N_16852);
or U17166 (N_17166,N_16945,N_16869);
and U17167 (N_17167,N_16828,N_16910);
or U17168 (N_17168,N_16995,N_16841);
or U17169 (N_17169,N_16987,N_16839);
nor U17170 (N_17170,N_16983,N_16831);
and U17171 (N_17171,N_16842,N_16877);
nor U17172 (N_17172,N_16844,N_16980);
and U17173 (N_17173,N_16993,N_16899);
nand U17174 (N_17174,N_16921,N_16945);
and U17175 (N_17175,N_16835,N_16979);
and U17176 (N_17176,N_16954,N_16809);
nand U17177 (N_17177,N_16904,N_16935);
nor U17178 (N_17178,N_16990,N_16842);
nor U17179 (N_17179,N_16834,N_16822);
or U17180 (N_17180,N_16873,N_16803);
nand U17181 (N_17181,N_16904,N_16898);
and U17182 (N_17182,N_16842,N_16932);
or U17183 (N_17183,N_16806,N_16828);
or U17184 (N_17184,N_16964,N_16859);
or U17185 (N_17185,N_16983,N_16835);
nand U17186 (N_17186,N_16921,N_16943);
and U17187 (N_17187,N_16804,N_16999);
nand U17188 (N_17188,N_16880,N_16923);
and U17189 (N_17189,N_16873,N_16959);
or U17190 (N_17190,N_16845,N_16967);
or U17191 (N_17191,N_16815,N_16889);
nand U17192 (N_17192,N_16806,N_16808);
nand U17193 (N_17193,N_16971,N_16892);
and U17194 (N_17194,N_16854,N_16867);
nor U17195 (N_17195,N_16914,N_16980);
or U17196 (N_17196,N_16965,N_16909);
or U17197 (N_17197,N_16859,N_16920);
and U17198 (N_17198,N_16887,N_16966);
nor U17199 (N_17199,N_16998,N_16877);
or U17200 (N_17200,N_17039,N_17089);
nor U17201 (N_17201,N_17077,N_17132);
and U17202 (N_17202,N_17022,N_17188);
nor U17203 (N_17203,N_17195,N_17027);
nor U17204 (N_17204,N_17145,N_17103);
xnor U17205 (N_17205,N_17137,N_17197);
nor U17206 (N_17206,N_17163,N_17014);
or U17207 (N_17207,N_17151,N_17166);
nand U17208 (N_17208,N_17120,N_17033);
nor U17209 (N_17209,N_17141,N_17059);
nand U17210 (N_17210,N_17152,N_17026);
or U17211 (N_17211,N_17093,N_17168);
and U17212 (N_17212,N_17175,N_17143);
and U17213 (N_17213,N_17034,N_17123);
nor U17214 (N_17214,N_17119,N_17165);
and U17215 (N_17215,N_17199,N_17196);
or U17216 (N_17216,N_17020,N_17184);
nor U17217 (N_17217,N_17111,N_17019);
and U17218 (N_17218,N_17098,N_17158);
and U17219 (N_17219,N_17063,N_17045);
nor U17220 (N_17220,N_17105,N_17065);
and U17221 (N_17221,N_17162,N_17174);
or U17222 (N_17222,N_17154,N_17189);
nor U17223 (N_17223,N_17032,N_17040);
nand U17224 (N_17224,N_17044,N_17046);
nor U17225 (N_17225,N_17138,N_17112);
nor U17226 (N_17226,N_17085,N_17128);
nand U17227 (N_17227,N_17161,N_17191);
or U17228 (N_17228,N_17125,N_17172);
or U17229 (N_17229,N_17001,N_17179);
nand U17230 (N_17230,N_17198,N_17150);
and U17231 (N_17231,N_17011,N_17048);
or U17232 (N_17232,N_17104,N_17185);
and U17233 (N_17233,N_17121,N_17091);
or U17234 (N_17234,N_17095,N_17181);
or U17235 (N_17235,N_17117,N_17017);
or U17236 (N_17236,N_17101,N_17008);
nand U17237 (N_17237,N_17167,N_17072);
nand U17238 (N_17238,N_17142,N_17130);
nand U17239 (N_17239,N_17133,N_17030);
xnor U17240 (N_17240,N_17157,N_17109);
and U17241 (N_17241,N_17180,N_17002);
or U17242 (N_17242,N_17097,N_17135);
nor U17243 (N_17243,N_17094,N_17164);
nor U17244 (N_17244,N_17038,N_17087);
or U17245 (N_17245,N_17066,N_17170);
nor U17246 (N_17246,N_17193,N_17074);
nand U17247 (N_17247,N_17054,N_17136);
or U17248 (N_17248,N_17069,N_17041);
or U17249 (N_17249,N_17155,N_17025);
nand U17250 (N_17250,N_17187,N_17062);
and U17251 (N_17251,N_17052,N_17090);
nor U17252 (N_17252,N_17192,N_17176);
xnor U17253 (N_17253,N_17183,N_17144);
or U17254 (N_17254,N_17140,N_17139);
or U17255 (N_17255,N_17043,N_17000);
or U17256 (N_17256,N_17073,N_17114);
nand U17257 (N_17257,N_17178,N_17083);
nor U17258 (N_17258,N_17115,N_17042);
and U17259 (N_17259,N_17028,N_17071);
and U17260 (N_17260,N_17035,N_17056);
nor U17261 (N_17261,N_17182,N_17118);
or U17262 (N_17262,N_17160,N_17129);
or U17263 (N_17263,N_17024,N_17096);
nor U17264 (N_17264,N_17009,N_17190);
nor U17265 (N_17265,N_17021,N_17092);
nand U17266 (N_17266,N_17081,N_17080);
nand U17267 (N_17267,N_17088,N_17116);
and U17268 (N_17268,N_17159,N_17029);
nand U17269 (N_17269,N_17061,N_17075);
and U17270 (N_17270,N_17004,N_17055);
and U17271 (N_17271,N_17005,N_17127);
nor U17272 (N_17272,N_17057,N_17194);
nor U17273 (N_17273,N_17050,N_17079);
and U17274 (N_17274,N_17070,N_17134);
or U17275 (N_17275,N_17113,N_17102);
and U17276 (N_17276,N_17012,N_17126);
nor U17277 (N_17277,N_17067,N_17013);
and U17278 (N_17278,N_17007,N_17147);
and U17279 (N_17279,N_17131,N_17099);
and U17280 (N_17280,N_17010,N_17047);
and U17281 (N_17281,N_17049,N_17110);
nor U17282 (N_17282,N_17146,N_17060);
nor U17283 (N_17283,N_17173,N_17086);
nor U17284 (N_17284,N_17058,N_17169);
nand U17285 (N_17285,N_17076,N_17068);
or U17286 (N_17286,N_17106,N_17149);
and U17287 (N_17287,N_17148,N_17186);
and U17288 (N_17288,N_17064,N_17023);
and U17289 (N_17289,N_17015,N_17051);
and U17290 (N_17290,N_17100,N_17082);
and U17291 (N_17291,N_17171,N_17177);
nand U17292 (N_17292,N_17122,N_17078);
and U17293 (N_17293,N_17108,N_17016);
nand U17294 (N_17294,N_17006,N_17037);
nand U17295 (N_17295,N_17084,N_17003);
nand U17296 (N_17296,N_17107,N_17156);
and U17297 (N_17297,N_17018,N_17053);
nor U17298 (N_17298,N_17036,N_17031);
nor U17299 (N_17299,N_17124,N_17153);
or U17300 (N_17300,N_17196,N_17141);
nand U17301 (N_17301,N_17188,N_17045);
or U17302 (N_17302,N_17121,N_17054);
nand U17303 (N_17303,N_17056,N_17023);
or U17304 (N_17304,N_17099,N_17031);
or U17305 (N_17305,N_17167,N_17173);
or U17306 (N_17306,N_17127,N_17126);
nand U17307 (N_17307,N_17107,N_17198);
and U17308 (N_17308,N_17077,N_17178);
or U17309 (N_17309,N_17127,N_17096);
and U17310 (N_17310,N_17002,N_17199);
nand U17311 (N_17311,N_17146,N_17054);
or U17312 (N_17312,N_17184,N_17191);
nor U17313 (N_17313,N_17045,N_17061);
or U17314 (N_17314,N_17044,N_17117);
or U17315 (N_17315,N_17126,N_17005);
nand U17316 (N_17316,N_17142,N_17012);
and U17317 (N_17317,N_17177,N_17119);
or U17318 (N_17318,N_17102,N_17011);
nand U17319 (N_17319,N_17018,N_17017);
and U17320 (N_17320,N_17018,N_17158);
or U17321 (N_17321,N_17072,N_17155);
nand U17322 (N_17322,N_17056,N_17160);
and U17323 (N_17323,N_17113,N_17179);
or U17324 (N_17324,N_17020,N_17135);
or U17325 (N_17325,N_17009,N_17124);
or U17326 (N_17326,N_17119,N_17088);
and U17327 (N_17327,N_17160,N_17060);
and U17328 (N_17328,N_17128,N_17133);
nand U17329 (N_17329,N_17053,N_17113);
and U17330 (N_17330,N_17183,N_17126);
and U17331 (N_17331,N_17060,N_17081);
or U17332 (N_17332,N_17072,N_17123);
or U17333 (N_17333,N_17069,N_17091);
or U17334 (N_17334,N_17099,N_17051);
nor U17335 (N_17335,N_17170,N_17175);
and U17336 (N_17336,N_17079,N_17118);
and U17337 (N_17337,N_17129,N_17016);
and U17338 (N_17338,N_17045,N_17172);
or U17339 (N_17339,N_17014,N_17006);
and U17340 (N_17340,N_17079,N_17072);
or U17341 (N_17341,N_17135,N_17090);
or U17342 (N_17342,N_17170,N_17108);
nor U17343 (N_17343,N_17050,N_17002);
nand U17344 (N_17344,N_17132,N_17131);
nor U17345 (N_17345,N_17036,N_17198);
nor U17346 (N_17346,N_17046,N_17048);
nor U17347 (N_17347,N_17185,N_17190);
nor U17348 (N_17348,N_17129,N_17138);
nor U17349 (N_17349,N_17017,N_17163);
or U17350 (N_17350,N_17196,N_17193);
and U17351 (N_17351,N_17198,N_17033);
or U17352 (N_17352,N_17065,N_17169);
and U17353 (N_17353,N_17169,N_17144);
nor U17354 (N_17354,N_17106,N_17185);
nand U17355 (N_17355,N_17061,N_17195);
and U17356 (N_17356,N_17067,N_17069);
nor U17357 (N_17357,N_17132,N_17051);
and U17358 (N_17358,N_17120,N_17056);
xor U17359 (N_17359,N_17109,N_17173);
and U17360 (N_17360,N_17019,N_17071);
nor U17361 (N_17361,N_17079,N_17067);
nand U17362 (N_17362,N_17037,N_17105);
or U17363 (N_17363,N_17073,N_17023);
nor U17364 (N_17364,N_17141,N_17009);
nand U17365 (N_17365,N_17057,N_17116);
or U17366 (N_17366,N_17093,N_17103);
nand U17367 (N_17367,N_17057,N_17125);
nor U17368 (N_17368,N_17132,N_17050);
nor U17369 (N_17369,N_17197,N_17083);
and U17370 (N_17370,N_17058,N_17135);
or U17371 (N_17371,N_17182,N_17100);
or U17372 (N_17372,N_17112,N_17044);
nand U17373 (N_17373,N_17116,N_17191);
nor U17374 (N_17374,N_17199,N_17180);
or U17375 (N_17375,N_17147,N_17104);
nand U17376 (N_17376,N_17028,N_17027);
nand U17377 (N_17377,N_17050,N_17189);
nor U17378 (N_17378,N_17037,N_17091);
nor U17379 (N_17379,N_17044,N_17174);
and U17380 (N_17380,N_17096,N_17045);
nor U17381 (N_17381,N_17038,N_17048);
nor U17382 (N_17382,N_17029,N_17177);
nand U17383 (N_17383,N_17019,N_17170);
and U17384 (N_17384,N_17060,N_17074);
or U17385 (N_17385,N_17004,N_17136);
nand U17386 (N_17386,N_17088,N_17046);
or U17387 (N_17387,N_17025,N_17096);
nand U17388 (N_17388,N_17089,N_17082);
or U17389 (N_17389,N_17007,N_17112);
nand U17390 (N_17390,N_17051,N_17043);
or U17391 (N_17391,N_17149,N_17039);
and U17392 (N_17392,N_17124,N_17116);
and U17393 (N_17393,N_17061,N_17165);
and U17394 (N_17394,N_17127,N_17029);
or U17395 (N_17395,N_17070,N_17157);
and U17396 (N_17396,N_17016,N_17191);
nor U17397 (N_17397,N_17161,N_17178);
nand U17398 (N_17398,N_17133,N_17060);
and U17399 (N_17399,N_17061,N_17035);
or U17400 (N_17400,N_17333,N_17270);
and U17401 (N_17401,N_17353,N_17382);
nand U17402 (N_17402,N_17218,N_17209);
nand U17403 (N_17403,N_17386,N_17280);
and U17404 (N_17404,N_17349,N_17297);
or U17405 (N_17405,N_17221,N_17294);
nor U17406 (N_17406,N_17291,N_17376);
or U17407 (N_17407,N_17346,N_17360);
nor U17408 (N_17408,N_17358,N_17251);
nor U17409 (N_17409,N_17398,N_17310);
nor U17410 (N_17410,N_17350,N_17230);
or U17411 (N_17411,N_17332,N_17240);
or U17412 (N_17412,N_17264,N_17306);
nor U17413 (N_17413,N_17385,N_17371);
and U17414 (N_17414,N_17277,N_17312);
or U17415 (N_17415,N_17212,N_17387);
nand U17416 (N_17416,N_17330,N_17394);
nand U17417 (N_17417,N_17399,N_17302);
nand U17418 (N_17418,N_17229,N_17228);
nand U17419 (N_17419,N_17362,N_17288);
or U17420 (N_17420,N_17274,N_17241);
nand U17421 (N_17421,N_17269,N_17282);
or U17422 (N_17422,N_17328,N_17260);
nand U17423 (N_17423,N_17359,N_17308);
and U17424 (N_17424,N_17276,N_17272);
or U17425 (N_17425,N_17369,N_17388);
and U17426 (N_17426,N_17314,N_17357);
nand U17427 (N_17427,N_17342,N_17204);
nor U17428 (N_17428,N_17313,N_17324);
or U17429 (N_17429,N_17256,N_17309);
nor U17430 (N_17430,N_17389,N_17210);
nand U17431 (N_17431,N_17372,N_17345);
or U17432 (N_17432,N_17374,N_17238);
and U17433 (N_17433,N_17242,N_17225);
or U17434 (N_17434,N_17370,N_17396);
and U17435 (N_17435,N_17379,N_17275);
nor U17436 (N_17436,N_17223,N_17364);
or U17437 (N_17437,N_17239,N_17261);
nand U17438 (N_17438,N_17319,N_17356);
or U17439 (N_17439,N_17395,N_17208);
and U17440 (N_17440,N_17232,N_17205);
nor U17441 (N_17441,N_17340,N_17284);
nand U17442 (N_17442,N_17258,N_17327);
nor U17443 (N_17443,N_17317,N_17321);
nand U17444 (N_17444,N_17281,N_17263);
nand U17445 (N_17445,N_17303,N_17219);
or U17446 (N_17446,N_17366,N_17207);
nor U17447 (N_17447,N_17202,N_17335);
or U17448 (N_17448,N_17391,N_17311);
or U17449 (N_17449,N_17273,N_17300);
or U17450 (N_17450,N_17380,N_17206);
or U17451 (N_17451,N_17293,N_17338);
or U17452 (N_17452,N_17355,N_17244);
nand U17453 (N_17453,N_17249,N_17341);
or U17454 (N_17454,N_17247,N_17334);
or U17455 (N_17455,N_17336,N_17320);
or U17456 (N_17456,N_17354,N_17290);
nand U17457 (N_17457,N_17268,N_17234);
or U17458 (N_17458,N_17254,N_17255);
nand U17459 (N_17459,N_17315,N_17326);
and U17460 (N_17460,N_17233,N_17292);
nor U17461 (N_17461,N_17286,N_17226);
nand U17462 (N_17462,N_17316,N_17213);
or U17463 (N_17463,N_17217,N_17262);
and U17464 (N_17464,N_17243,N_17211);
nor U17465 (N_17465,N_17250,N_17305);
and U17466 (N_17466,N_17237,N_17325);
and U17467 (N_17467,N_17289,N_17278);
nand U17468 (N_17468,N_17351,N_17304);
or U17469 (N_17469,N_17363,N_17331);
or U17470 (N_17470,N_17279,N_17267);
nand U17471 (N_17471,N_17236,N_17347);
and U17472 (N_17472,N_17339,N_17283);
nand U17473 (N_17473,N_17322,N_17298);
and U17474 (N_17474,N_17220,N_17253);
nor U17475 (N_17475,N_17295,N_17344);
nand U17476 (N_17476,N_17235,N_17231);
and U17477 (N_17477,N_17266,N_17390);
or U17478 (N_17478,N_17348,N_17271);
or U17479 (N_17479,N_17384,N_17299);
and U17480 (N_17480,N_17318,N_17381);
nand U17481 (N_17481,N_17287,N_17285);
and U17482 (N_17482,N_17365,N_17296);
nor U17483 (N_17483,N_17227,N_17329);
or U17484 (N_17484,N_17392,N_17377);
or U17485 (N_17485,N_17248,N_17383);
or U17486 (N_17486,N_17224,N_17307);
nand U17487 (N_17487,N_17343,N_17245);
and U17488 (N_17488,N_17397,N_17378);
nand U17489 (N_17489,N_17301,N_17246);
or U17490 (N_17490,N_17259,N_17203);
and U17491 (N_17491,N_17216,N_17214);
xor U17492 (N_17492,N_17373,N_17352);
or U17493 (N_17493,N_17252,N_17222);
nand U17494 (N_17494,N_17337,N_17367);
and U17495 (N_17495,N_17323,N_17265);
or U17496 (N_17496,N_17201,N_17361);
nand U17497 (N_17497,N_17393,N_17200);
nand U17498 (N_17498,N_17257,N_17375);
or U17499 (N_17499,N_17215,N_17368);
nor U17500 (N_17500,N_17361,N_17340);
nor U17501 (N_17501,N_17395,N_17244);
nor U17502 (N_17502,N_17329,N_17377);
nor U17503 (N_17503,N_17332,N_17366);
or U17504 (N_17504,N_17279,N_17238);
or U17505 (N_17505,N_17298,N_17358);
nand U17506 (N_17506,N_17280,N_17360);
or U17507 (N_17507,N_17338,N_17220);
and U17508 (N_17508,N_17315,N_17357);
nand U17509 (N_17509,N_17242,N_17356);
or U17510 (N_17510,N_17389,N_17249);
nor U17511 (N_17511,N_17202,N_17367);
nor U17512 (N_17512,N_17210,N_17353);
or U17513 (N_17513,N_17248,N_17258);
nor U17514 (N_17514,N_17344,N_17292);
nor U17515 (N_17515,N_17331,N_17275);
and U17516 (N_17516,N_17217,N_17263);
and U17517 (N_17517,N_17261,N_17225);
or U17518 (N_17518,N_17372,N_17214);
nand U17519 (N_17519,N_17232,N_17349);
or U17520 (N_17520,N_17371,N_17275);
or U17521 (N_17521,N_17327,N_17331);
nor U17522 (N_17522,N_17391,N_17216);
and U17523 (N_17523,N_17368,N_17224);
nand U17524 (N_17524,N_17375,N_17356);
or U17525 (N_17525,N_17388,N_17280);
nand U17526 (N_17526,N_17379,N_17351);
nand U17527 (N_17527,N_17374,N_17266);
and U17528 (N_17528,N_17251,N_17275);
nor U17529 (N_17529,N_17279,N_17292);
and U17530 (N_17530,N_17363,N_17254);
nor U17531 (N_17531,N_17228,N_17216);
or U17532 (N_17532,N_17256,N_17366);
and U17533 (N_17533,N_17227,N_17385);
and U17534 (N_17534,N_17312,N_17297);
nor U17535 (N_17535,N_17368,N_17218);
and U17536 (N_17536,N_17276,N_17315);
and U17537 (N_17537,N_17253,N_17338);
nand U17538 (N_17538,N_17267,N_17240);
nand U17539 (N_17539,N_17347,N_17336);
and U17540 (N_17540,N_17302,N_17230);
nor U17541 (N_17541,N_17266,N_17386);
nor U17542 (N_17542,N_17391,N_17346);
or U17543 (N_17543,N_17228,N_17203);
nand U17544 (N_17544,N_17379,N_17297);
or U17545 (N_17545,N_17339,N_17290);
nand U17546 (N_17546,N_17392,N_17370);
and U17547 (N_17547,N_17203,N_17300);
nor U17548 (N_17548,N_17205,N_17297);
and U17549 (N_17549,N_17200,N_17265);
or U17550 (N_17550,N_17376,N_17312);
or U17551 (N_17551,N_17293,N_17230);
nand U17552 (N_17552,N_17346,N_17397);
and U17553 (N_17553,N_17253,N_17347);
nand U17554 (N_17554,N_17246,N_17388);
and U17555 (N_17555,N_17359,N_17334);
or U17556 (N_17556,N_17265,N_17253);
nor U17557 (N_17557,N_17260,N_17350);
and U17558 (N_17558,N_17336,N_17229);
nand U17559 (N_17559,N_17391,N_17277);
and U17560 (N_17560,N_17367,N_17332);
and U17561 (N_17561,N_17274,N_17344);
and U17562 (N_17562,N_17375,N_17240);
nor U17563 (N_17563,N_17301,N_17240);
or U17564 (N_17564,N_17350,N_17204);
or U17565 (N_17565,N_17349,N_17224);
nand U17566 (N_17566,N_17232,N_17297);
xnor U17567 (N_17567,N_17357,N_17233);
nand U17568 (N_17568,N_17383,N_17322);
and U17569 (N_17569,N_17381,N_17283);
or U17570 (N_17570,N_17211,N_17297);
or U17571 (N_17571,N_17334,N_17386);
or U17572 (N_17572,N_17255,N_17272);
nor U17573 (N_17573,N_17332,N_17294);
nand U17574 (N_17574,N_17286,N_17374);
or U17575 (N_17575,N_17268,N_17277);
and U17576 (N_17576,N_17228,N_17261);
nor U17577 (N_17577,N_17225,N_17393);
nor U17578 (N_17578,N_17261,N_17283);
nor U17579 (N_17579,N_17251,N_17312);
and U17580 (N_17580,N_17299,N_17208);
nand U17581 (N_17581,N_17254,N_17333);
and U17582 (N_17582,N_17214,N_17290);
nand U17583 (N_17583,N_17323,N_17279);
nand U17584 (N_17584,N_17228,N_17327);
and U17585 (N_17585,N_17386,N_17377);
nor U17586 (N_17586,N_17307,N_17229);
and U17587 (N_17587,N_17275,N_17337);
and U17588 (N_17588,N_17214,N_17223);
or U17589 (N_17589,N_17383,N_17368);
and U17590 (N_17590,N_17206,N_17366);
nor U17591 (N_17591,N_17345,N_17278);
and U17592 (N_17592,N_17239,N_17312);
nand U17593 (N_17593,N_17203,N_17337);
and U17594 (N_17594,N_17222,N_17249);
nor U17595 (N_17595,N_17211,N_17227);
nor U17596 (N_17596,N_17356,N_17321);
or U17597 (N_17597,N_17297,N_17396);
or U17598 (N_17598,N_17228,N_17333);
or U17599 (N_17599,N_17235,N_17293);
or U17600 (N_17600,N_17559,N_17405);
nand U17601 (N_17601,N_17459,N_17419);
nor U17602 (N_17602,N_17521,N_17560);
nor U17603 (N_17603,N_17415,N_17501);
and U17604 (N_17604,N_17580,N_17575);
and U17605 (N_17605,N_17451,N_17408);
and U17606 (N_17606,N_17538,N_17541);
and U17607 (N_17607,N_17561,N_17482);
and U17608 (N_17608,N_17484,N_17534);
and U17609 (N_17609,N_17495,N_17444);
nor U17610 (N_17610,N_17587,N_17545);
and U17611 (N_17611,N_17514,N_17585);
nand U17612 (N_17612,N_17450,N_17567);
nor U17613 (N_17613,N_17491,N_17520);
nor U17614 (N_17614,N_17410,N_17557);
nor U17615 (N_17615,N_17518,N_17493);
and U17616 (N_17616,N_17463,N_17583);
or U17617 (N_17617,N_17490,N_17531);
nand U17618 (N_17618,N_17515,N_17417);
nor U17619 (N_17619,N_17533,N_17414);
nand U17620 (N_17620,N_17548,N_17547);
nor U17621 (N_17621,N_17599,N_17523);
nand U17622 (N_17622,N_17563,N_17421);
and U17623 (N_17623,N_17413,N_17588);
nor U17624 (N_17624,N_17467,N_17532);
or U17625 (N_17625,N_17566,N_17464);
or U17626 (N_17626,N_17589,N_17420);
nor U17627 (N_17627,N_17553,N_17497);
nor U17628 (N_17628,N_17437,N_17487);
or U17629 (N_17629,N_17546,N_17506);
nand U17630 (N_17630,N_17452,N_17536);
and U17631 (N_17631,N_17586,N_17594);
or U17632 (N_17632,N_17574,N_17539);
nor U17633 (N_17633,N_17425,N_17412);
nand U17634 (N_17634,N_17512,N_17552);
nand U17635 (N_17635,N_17436,N_17542);
and U17636 (N_17636,N_17554,N_17486);
or U17637 (N_17637,N_17446,N_17462);
or U17638 (N_17638,N_17424,N_17492);
nand U17639 (N_17639,N_17505,N_17562);
nand U17640 (N_17640,N_17481,N_17576);
nand U17641 (N_17641,N_17422,N_17433);
and U17642 (N_17642,N_17503,N_17418);
and U17643 (N_17643,N_17579,N_17440);
nor U17644 (N_17644,N_17590,N_17525);
nor U17645 (N_17645,N_17569,N_17456);
nor U17646 (N_17646,N_17428,N_17537);
or U17647 (N_17647,N_17592,N_17455);
nor U17648 (N_17648,N_17477,N_17475);
nand U17649 (N_17649,N_17488,N_17435);
nor U17650 (N_17650,N_17595,N_17401);
nand U17651 (N_17651,N_17441,N_17578);
and U17652 (N_17652,N_17544,N_17406);
nor U17653 (N_17653,N_17485,N_17517);
nand U17654 (N_17654,N_17598,N_17522);
and U17655 (N_17655,N_17502,N_17483);
and U17656 (N_17656,N_17411,N_17403);
nor U17657 (N_17657,N_17543,N_17478);
nor U17658 (N_17658,N_17442,N_17527);
xor U17659 (N_17659,N_17572,N_17516);
nor U17660 (N_17660,N_17584,N_17509);
xor U17661 (N_17661,N_17510,N_17458);
nor U17662 (N_17662,N_17429,N_17461);
or U17663 (N_17663,N_17489,N_17472);
nor U17664 (N_17664,N_17551,N_17581);
or U17665 (N_17665,N_17404,N_17558);
nand U17666 (N_17666,N_17573,N_17582);
nor U17667 (N_17667,N_17568,N_17471);
nand U17668 (N_17668,N_17508,N_17409);
and U17669 (N_17669,N_17480,N_17550);
or U17670 (N_17670,N_17479,N_17565);
or U17671 (N_17671,N_17528,N_17474);
or U17672 (N_17672,N_17524,N_17476);
or U17673 (N_17673,N_17457,N_17494);
or U17674 (N_17674,N_17473,N_17454);
nand U17675 (N_17675,N_17564,N_17469);
nand U17676 (N_17676,N_17439,N_17519);
or U17677 (N_17677,N_17468,N_17407);
nor U17678 (N_17678,N_17593,N_17453);
nand U17679 (N_17679,N_17465,N_17438);
and U17680 (N_17680,N_17499,N_17577);
nor U17681 (N_17681,N_17445,N_17498);
nor U17682 (N_17682,N_17535,N_17596);
nand U17683 (N_17683,N_17400,N_17426);
and U17684 (N_17684,N_17432,N_17434);
nand U17685 (N_17685,N_17402,N_17443);
and U17686 (N_17686,N_17427,N_17526);
or U17687 (N_17687,N_17556,N_17570);
nor U17688 (N_17688,N_17549,N_17449);
and U17689 (N_17689,N_17448,N_17513);
or U17690 (N_17690,N_17529,N_17530);
nand U17691 (N_17691,N_17496,N_17447);
and U17692 (N_17692,N_17416,N_17500);
or U17693 (N_17693,N_17504,N_17470);
and U17694 (N_17694,N_17431,N_17597);
and U17695 (N_17695,N_17466,N_17555);
or U17696 (N_17696,N_17591,N_17511);
nand U17697 (N_17697,N_17430,N_17460);
nand U17698 (N_17698,N_17423,N_17507);
nor U17699 (N_17699,N_17571,N_17540);
nor U17700 (N_17700,N_17533,N_17428);
or U17701 (N_17701,N_17424,N_17538);
nor U17702 (N_17702,N_17594,N_17481);
and U17703 (N_17703,N_17426,N_17549);
or U17704 (N_17704,N_17402,N_17446);
nand U17705 (N_17705,N_17577,N_17423);
nand U17706 (N_17706,N_17434,N_17421);
or U17707 (N_17707,N_17439,N_17596);
and U17708 (N_17708,N_17454,N_17442);
nor U17709 (N_17709,N_17416,N_17443);
or U17710 (N_17710,N_17434,N_17505);
and U17711 (N_17711,N_17577,N_17432);
nand U17712 (N_17712,N_17435,N_17464);
and U17713 (N_17713,N_17464,N_17549);
or U17714 (N_17714,N_17595,N_17448);
nand U17715 (N_17715,N_17546,N_17431);
or U17716 (N_17716,N_17508,N_17442);
nand U17717 (N_17717,N_17443,N_17533);
or U17718 (N_17718,N_17535,N_17594);
nor U17719 (N_17719,N_17535,N_17536);
nand U17720 (N_17720,N_17506,N_17552);
xor U17721 (N_17721,N_17521,N_17485);
nor U17722 (N_17722,N_17545,N_17425);
nor U17723 (N_17723,N_17495,N_17550);
nand U17724 (N_17724,N_17405,N_17538);
or U17725 (N_17725,N_17451,N_17447);
nor U17726 (N_17726,N_17571,N_17406);
or U17727 (N_17727,N_17460,N_17531);
and U17728 (N_17728,N_17446,N_17578);
and U17729 (N_17729,N_17400,N_17440);
nor U17730 (N_17730,N_17427,N_17423);
or U17731 (N_17731,N_17431,N_17435);
and U17732 (N_17732,N_17457,N_17447);
nand U17733 (N_17733,N_17569,N_17502);
nand U17734 (N_17734,N_17424,N_17597);
nor U17735 (N_17735,N_17454,N_17413);
nand U17736 (N_17736,N_17539,N_17564);
nor U17737 (N_17737,N_17413,N_17571);
or U17738 (N_17738,N_17411,N_17421);
and U17739 (N_17739,N_17475,N_17402);
nor U17740 (N_17740,N_17467,N_17482);
or U17741 (N_17741,N_17528,N_17452);
or U17742 (N_17742,N_17563,N_17497);
nand U17743 (N_17743,N_17438,N_17400);
or U17744 (N_17744,N_17576,N_17419);
nand U17745 (N_17745,N_17537,N_17476);
and U17746 (N_17746,N_17504,N_17536);
and U17747 (N_17747,N_17488,N_17442);
and U17748 (N_17748,N_17526,N_17474);
nand U17749 (N_17749,N_17433,N_17540);
nand U17750 (N_17750,N_17585,N_17460);
nand U17751 (N_17751,N_17408,N_17593);
nor U17752 (N_17752,N_17499,N_17578);
nor U17753 (N_17753,N_17486,N_17511);
and U17754 (N_17754,N_17560,N_17510);
nand U17755 (N_17755,N_17512,N_17594);
nor U17756 (N_17756,N_17538,N_17524);
nor U17757 (N_17757,N_17492,N_17449);
nor U17758 (N_17758,N_17453,N_17410);
or U17759 (N_17759,N_17508,N_17400);
or U17760 (N_17760,N_17400,N_17541);
and U17761 (N_17761,N_17473,N_17505);
nand U17762 (N_17762,N_17580,N_17447);
or U17763 (N_17763,N_17528,N_17587);
nor U17764 (N_17764,N_17443,N_17424);
nand U17765 (N_17765,N_17416,N_17402);
or U17766 (N_17766,N_17542,N_17501);
xnor U17767 (N_17767,N_17518,N_17454);
or U17768 (N_17768,N_17536,N_17462);
nand U17769 (N_17769,N_17403,N_17562);
nand U17770 (N_17770,N_17410,N_17503);
nand U17771 (N_17771,N_17452,N_17566);
and U17772 (N_17772,N_17537,N_17449);
or U17773 (N_17773,N_17593,N_17495);
nand U17774 (N_17774,N_17436,N_17480);
nand U17775 (N_17775,N_17477,N_17412);
and U17776 (N_17776,N_17584,N_17504);
nor U17777 (N_17777,N_17587,N_17560);
nor U17778 (N_17778,N_17494,N_17566);
nor U17779 (N_17779,N_17413,N_17482);
and U17780 (N_17780,N_17455,N_17419);
nor U17781 (N_17781,N_17589,N_17417);
nand U17782 (N_17782,N_17482,N_17570);
or U17783 (N_17783,N_17523,N_17559);
nor U17784 (N_17784,N_17512,N_17528);
or U17785 (N_17785,N_17412,N_17593);
and U17786 (N_17786,N_17531,N_17561);
or U17787 (N_17787,N_17506,N_17573);
or U17788 (N_17788,N_17568,N_17430);
nor U17789 (N_17789,N_17460,N_17492);
nor U17790 (N_17790,N_17412,N_17424);
or U17791 (N_17791,N_17445,N_17546);
and U17792 (N_17792,N_17444,N_17501);
or U17793 (N_17793,N_17491,N_17446);
nand U17794 (N_17794,N_17463,N_17425);
nor U17795 (N_17795,N_17596,N_17533);
nor U17796 (N_17796,N_17520,N_17528);
nand U17797 (N_17797,N_17505,N_17570);
nor U17798 (N_17798,N_17500,N_17512);
xor U17799 (N_17799,N_17436,N_17457);
or U17800 (N_17800,N_17733,N_17710);
or U17801 (N_17801,N_17704,N_17785);
or U17802 (N_17802,N_17631,N_17609);
and U17803 (N_17803,N_17762,N_17787);
nor U17804 (N_17804,N_17638,N_17669);
or U17805 (N_17805,N_17628,N_17684);
nand U17806 (N_17806,N_17707,N_17650);
or U17807 (N_17807,N_17616,N_17709);
and U17808 (N_17808,N_17685,N_17747);
nand U17809 (N_17809,N_17605,N_17770);
nand U17810 (N_17810,N_17720,N_17600);
nor U17811 (N_17811,N_17651,N_17672);
nor U17812 (N_17812,N_17696,N_17758);
nand U17813 (N_17813,N_17798,N_17659);
nand U17814 (N_17814,N_17732,N_17649);
and U17815 (N_17815,N_17752,N_17694);
and U17816 (N_17816,N_17686,N_17719);
nor U17817 (N_17817,N_17602,N_17708);
and U17818 (N_17818,N_17679,N_17794);
nor U17819 (N_17819,N_17706,N_17682);
nor U17820 (N_17820,N_17663,N_17639);
or U17821 (N_17821,N_17671,N_17613);
nor U17822 (N_17822,N_17763,N_17657);
and U17823 (N_17823,N_17665,N_17648);
nand U17824 (N_17824,N_17676,N_17797);
and U17825 (N_17825,N_17703,N_17624);
nand U17826 (N_17826,N_17683,N_17788);
nor U17827 (N_17827,N_17688,N_17637);
or U17828 (N_17828,N_17796,N_17627);
and U17829 (N_17829,N_17674,N_17635);
nand U17830 (N_17830,N_17606,N_17718);
and U17831 (N_17831,N_17656,N_17791);
nand U17832 (N_17832,N_17781,N_17601);
or U17833 (N_17833,N_17626,N_17615);
nor U17834 (N_17834,N_17701,N_17714);
nor U17835 (N_17835,N_17652,N_17730);
nor U17836 (N_17836,N_17632,N_17680);
nand U17837 (N_17837,N_17670,N_17799);
nor U17838 (N_17838,N_17617,N_17748);
and U17839 (N_17839,N_17729,N_17761);
nor U17840 (N_17840,N_17692,N_17724);
and U17841 (N_17841,N_17666,N_17677);
nor U17842 (N_17842,N_17608,N_17689);
xor U17843 (N_17843,N_17619,N_17612);
or U17844 (N_17844,N_17636,N_17646);
nand U17845 (N_17845,N_17695,N_17661);
and U17846 (N_17846,N_17765,N_17620);
or U17847 (N_17847,N_17630,N_17725);
nand U17848 (N_17848,N_17726,N_17634);
nor U17849 (N_17849,N_17717,N_17705);
nand U17850 (N_17850,N_17793,N_17690);
or U17851 (N_17851,N_17739,N_17660);
and U17852 (N_17852,N_17603,N_17764);
and U17853 (N_17853,N_17675,N_17751);
nor U17854 (N_17854,N_17643,N_17776);
and U17855 (N_17855,N_17711,N_17697);
nand U17856 (N_17856,N_17778,N_17712);
nand U17857 (N_17857,N_17702,N_17644);
nand U17858 (N_17858,N_17723,N_17795);
or U17859 (N_17859,N_17716,N_17755);
or U17860 (N_17860,N_17611,N_17750);
xnor U17861 (N_17861,N_17654,N_17662);
and U17862 (N_17862,N_17784,N_17618);
nor U17863 (N_17863,N_17771,N_17792);
nor U17864 (N_17864,N_17610,N_17741);
and U17865 (N_17865,N_17740,N_17721);
nand U17866 (N_17866,N_17667,N_17713);
or U17867 (N_17867,N_17773,N_17736);
nand U17868 (N_17868,N_17744,N_17746);
or U17869 (N_17869,N_17737,N_17715);
nand U17870 (N_17870,N_17743,N_17623);
nor U17871 (N_17871,N_17780,N_17699);
and U17872 (N_17872,N_17777,N_17673);
nand U17873 (N_17873,N_17607,N_17664);
or U17874 (N_17874,N_17772,N_17621);
nand U17875 (N_17875,N_17789,N_17653);
xor U17876 (N_17876,N_17678,N_17658);
nor U17877 (N_17877,N_17645,N_17691);
and U17878 (N_17878,N_17754,N_17735);
or U17879 (N_17879,N_17641,N_17745);
nand U17880 (N_17880,N_17687,N_17614);
and U17881 (N_17881,N_17738,N_17700);
nand U17882 (N_17882,N_17779,N_17642);
or U17883 (N_17883,N_17742,N_17749);
nand U17884 (N_17884,N_17633,N_17625);
xor U17885 (N_17885,N_17655,N_17731);
nand U17886 (N_17886,N_17722,N_17734);
and U17887 (N_17887,N_17604,N_17629);
nor U17888 (N_17888,N_17769,N_17768);
nand U17889 (N_17889,N_17756,N_17757);
and U17890 (N_17890,N_17681,N_17783);
nand U17891 (N_17891,N_17786,N_17782);
or U17892 (N_17892,N_17790,N_17693);
nand U17893 (N_17893,N_17698,N_17760);
nand U17894 (N_17894,N_17767,N_17766);
or U17895 (N_17895,N_17668,N_17640);
and U17896 (N_17896,N_17775,N_17727);
or U17897 (N_17897,N_17647,N_17759);
or U17898 (N_17898,N_17753,N_17728);
nand U17899 (N_17899,N_17774,N_17622);
nand U17900 (N_17900,N_17719,N_17762);
or U17901 (N_17901,N_17775,N_17761);
nand U17902 (N_17902,N_17607,N_17750);
nand U17903 (N_17903,N_17763,N_17692);
nor U17904 (N_17904,N_17653,N_17634);
or U17905 (N_17905,N_17609,N_17695);
nor U17906 (N_17906,N_17648,N_17725);
and U17907 (N_17907,N_17700,N_17602);
nor U17908 (N_17908,N_17785,N_17708);
and U17909 (N_17909,N_17684,N_17642);
nand U17910 (N_17910,N_17734,N_17788);
or U17911 (N_17911,N_17655,N_17725);
nor U17912 (N_17912,N_17794,N_17785);
or U17913 (N_17913,N_17646,N_17700);
or U17914 (N_17914,N_17773,N_17714);
xnor U17915 (N_17915,N_17698,N_17629);
nand U17916 (N_17916,N_17618,N_17777);
or U17917 (N_17917,N_17769,N_17688);
or U17918 (N_17918,N_17774,N_17677);
nand U17919 (N_17919,N_17689,N_17715);
and U17920 (N_17920,N_17774,N_17767);
or U17921 (N_17921,N_17725,N_17707);
or U17922 (N_17922,N_17782,N_17693);
or U17923 (N_17923,N_17753,N_17716);
nor U17924 (N_17924,N_17761,N_17769);
nor U17925 (N_17925,N_17684,N_17773);
and U17926 (N_17926,N_17754,N_17718);
or U17927 (N_17927,N_17695,N_17644);
nand U17928 (N_17928,N_17610,N_17608);
or U17929 (N_17929,N_17764,N_17602);
nand U17930 (N_17930,N_17776,N_17777);
nor U17931 (N_17931,N_17688,N_17677);
nor U17932 (N_17932,N_17613,N_17607);
and U17933 (N_17933,N_17606,N_17702);
or U17934 (N_17934,N_17787,N_17638);
nand U17935 (N_17935,N_17738,N_17602);
nor U17936 (N_17936,N_17619,N_17722);
and U17937 (N_17937,N_17656,N_17683);
and U17938 (N_17938,N_17709,N_17766);
nand U17939 (N_17939,N_17766,N_17790);
nor U17940 (N_17940,N_17637,N_17712);
or U17941 (N_17941,N_17640,N_17744);
or U17942 (N_17942,N_17765,N_17693);
nand U17943 (N_17943,N_17780,N_17741);
nor U17944 (N_17944,N_17680,N_17620);
nand U17945 (N_17945,N_17733,N_17796);
nand U17946 (N_17946,N_17768,N_17689);
or U17947 (N_17947,N_17768,N_17690);
and U17948 (N_17948,N_17712,N_17711);
nand U17949 (N_17949,N_17642,N_17655);
or U17950 (N_17950,N_17692,N_17658);
nor U17951 (N_17951,N_17741,N_17747);
or U17952 (N_17952,N_17770,N_17722);
and U17953 (N_17953,N_17631,N_17792);
nor U17954 (N_17954,N_17756,N_17788);
nor U17955 (N_17955,N_17615,N_17682);
and U17956 (N_17956,N_17627,N_17789);
nor U17957 (N_17957,N_17604,N_17614);
nand U17958 (N_17958,N_17776,N_17773);
and U17959 (N_17959,N_17640,N_17670);
and U17960 (N_17960,N_17770,N_17639);
nand U17961 (N_17961,N_17712,N_17718);
xnor U17962 (N_17962,N_17718,N_17725);
or U17963 (N_17963,N_17646,N_17623);
or U17964 (N_17964,N_17669,N_17763);
and U17965 (N_17965,N_17746,N_17605);
or U17966 (N_17966,N_17769,N_17700);
nand U17967 (N_17967,N_17797,N_17745);
and U17968 (N_17968,N_17685,N_17638);
nand U17969 (N_17969,N_17773,N_17713);
nand U17970 (N_17970,N_17796,N_17693);
nor U17971 (N_17971,N_17733,N_17781);
or U17972 (N_17972,N_17730,N_17638);
nor U17973 (N_17973,N_17783,N_17759);
nor U17974 (N_17974,N_17606,N_17625);
nor U17975 (N_17975,N_17734,N_17752);
nand U17976 (N_17976,N_17706,N_17635);
xnor U17977 (N_17977,N_17714,N_17696);
nand U17978 (N_17978,N_17633,N_17661);
nor U17979 (N_17979,N_17767,N_17687);
or U17980 (N_17980,N_17666,N_17685);
nand U17981 (N_17981,N_17737,N_17667);
nand U17982 (N_17982,N_17660,N_17723);
nor U17983 (N_17983,N_17625,N_17665);
or U17984 (N_17984,N_17679,N_17690);
nand U17985 (N_17985,N_17705,N_17653);
nor U17986 (N_17986,N_17685,N_17627);
or U17987 (N_17987,N_17694,N_17791);
nor U17988 (N_17988,N_17740,N_17768);
nand U17989 (N_17989,N_17755,N_17724);
or U17990 (N_17990,N_17760,N_17711);
or U17991 (N_17991,N_17780,N_17671);
and U17992 (N_17992,N_17613,N_17736);
or U17993 (N_17993,N_17688,N_17674);
nor U17994 (N_17994,N_17793,N_17753);
or U17995 (N_17995,N_17625,N_17760);
nor U17996 (N_17996,N_17607,N_17697);
or U17997 (N_17997,N_17602,N_17643);
and U17998 (N_17998,N_17734,N_17616);
nor U17999 (N_17999,N_17716,N_17674);
and U18000 (N_18000,N_17839,N_17807);
nor U18001 (N_18001,N_17994,N_17969);
or U18002 (N_18002,N_17973,N_17997);
or U18003 (N_18003,N_17992,N_17963);
or U18004 (N_18004,N_17935,N_17873);
nor U18005 (N_18005,N_17898,N_17888);
or U18006 (N_18006,N_17837,N_17900);
nor U18007 (N_18007,N_17890,N_17891);
nand U18008 (N_18008,N_17852,N_17803);
nor U18009 (N_18009,N_17908,N_17828);
nand U18010 (N_18010,N_17966,N_17948);
nand U18011 (N_18011,N_17910,N_17868);
or U18012 (N_18012,N_17814,N_17860);
and U18013 (N_18013,N_17938,N_17939);
and U18014 (N_18014,N_17915,N_17981);
or U18015 (N_18015,N_17818,N_17974);
nand U18016 (N_18016,N_17995,N_17960);
and U18017 (N_18017,N_17846,N_17902);
and U18018 (N_18018,N_17949,N_17866);
or U18019 (N_18019,N_17806,N_17876);
nor U18020 (N_18020,N_17858,N_17917);
or U18021 (N_18021,N_17820,N_17952);
nor U18022 (N_18022,N_17930,N_17827);
nand U18023 (N_18023,N_17894,N_17850);
and U18024 (N_18024,N_17861,N_17901);
nor U18025 (N_18025,N_17853,N_17926);
and U18026 (N_18026,N_17986,N_17905);
nor U18027 (N_18027,N_17847,N_17921);
nor U18028 (N_18028,N_17931,N_17836);
nand U18029 (N_18029,N_17881,N_17976);
or U18030 (N_18030,N_17811,N_17843);
and U18031 (N_18031,N_17849,N_17989);
nand U18032 (N_18032,N_17810,N_17991);
or U18033 (N_18033,N_17877,N_17867);
and U18034 (N_18034,N_17848,N_17903);
nor U18035 (N_18035,N_17914,N_17895);
nor U18036 (N_18036,N_17862,N_17904);
nand U18037 (N_18037,N_17922,N_17943);
or U18038 (N_18038,N_17808,N_17856);
or U18039 (N_18039,N_17805,N_17893);
and U18040 (N_18040,N_17851,N_17979);
nor U18041 (N_18041,N_17800,N_17944);
nor U18042 (N_18042,N_17959,N_17940);
nor U18043 (N_18043,N_17968,N_17831);
nor U18044 (N_18044,N_17967,N_17998);
nand U18045 (N_18045,N_17886,N_17878);
nor U18046 (N_18046,N_17855,N_17845);
nand U18047 (N_18047,N_17971,N_17899);
nand U18048 (N_18048,N_17871,N_17869);
nand U18049 (N_18049,N_17859,N_17834);
nor U18050 (N_18050,N_17897,N_17980);
and U18051 (N_18051,N_17934,N_17880);
and U18052 (N_18052,N_17913,N_17985);
nor U18053 (N_18053,N_17887,N_17854);
or U18054 (N_18054,N_17835,N_17978);
nor U18055 (N_18055,N_17954,N_17865);
and U18056 (N_18056,N_17870,N_17955);
nor U18057 (N_18057,N_17924,N_17912);
xnor U18058 (N_18058,N_17885,N_17830);
nand U18059 (N_18059,N_17990,N_17923);
and U18060 (N_18060,N_17906,N_17947);
nand U18061 (N_18061,N_17984,N_17929);
nor U18062 (N_18062,N_17920,N_17925);
and U18063 (N_18063,N_17951,N_17829);
nor U18064 (N_18064,N_17961,N_17802);
nor U18065 (N_18065,N_17884,N_17987);
or U18066 (N_18066,N_17819,N_17909);
nand U18067 (N_18067,N_17993,N_17937);
and U18068 (N_18068,N_17950,N_17953);
and U18069 (N_18069,N_17932,N_17857);
nor U18070 (N_18070,N_17815,N_17941);
or U18071 (N_18071,N_17918,N_17942);
nand U18072 (N_18072,N_17824,N_17962);
and U18073 (N_18073,N_17911,N_17817);
or U18074 (N_18074,N_17833,N_17822);
nand U18075 (N_18075,N_17874,N_17889);
nor U18076 (N_18076,N_17936,N_17999);
or U18077 (N_18077,N_17832,N_17840);
and U18078 (N_18078,N_17896,N_17982);
or U18079 (N_18079,N_17842,N_17804);
and U18080 (N_18080,N_17970,N_17945);
and U18081 (N_18081,N_17879,N_17975);
nor U18082 (N_18082,N_17823,N_17864);
and U18083 (N_18083,N_17872,N_17916);
and U18084 (N_18084,N_17996,N_17957);
or U18085 (N_18085,N_17965,N_17927);
and U18086 (N_18086,N_17813,N_17825);
and U18087 (N_18087,N_17946,N_17983);
and U18088 (N_18088,N_17838,N_17928);
nor U18089 (N_18089,N_17977,N_17801);
nor U18090 (N_18090,N_17863,N_17821);
or U18091 (N_18091,N_17841,N_17812);
and U18092 (N_18092,N_17882,N_17892);
nand U18093 (N_18093,N_17809,N_17907);
nor U18094 (N_18094,N_17919,N_17883);
or U18095 (N_18095,N_17933,N_17956);
and U18096 (N_18096,N_17972,N_17826);
nand U18097 (N_18097,N_17875,N_17844);
or U18098 (N_18098,N_17958,N_17988);
or U18099 (N_18099,N_17964,N_17816);
nand U18100 (N_18100,N_17984,N_17832);
and U18101 (N_18101,N_17854,N_17839);
nand U18102 (N_18102,N_17869,N_17944);
and U18103 (N_18103,N_17926,N_17826);
or U18104 (N_18104,N_17934,N_17902);
nor U18105 (N_18105,N_17990,N_17907);
and U18106 (N_18106,N_17974,N_17831);
or U18107 (N_18107,N_17871,N_17929);
nor U18108 (N_18108,N_17989,N_17833);
or U18109 (N_18109,N_17891,N_17970);
nor U18110 (N_18110,N_17940,N_17812);
and U18111 (N_18111,N_17854,N_17810);
nand U18112 (N_18112,N_17915,N_17957);
or U18113 (N_18113,N_17805,N_17831);
nand U18114 (N_18114,N_17828,N_17899);
or U18115 (N_18115,N_17815,N_17899);
and U18116 (N_18116,N_17954,N_17997);
nand U18117 (N_18117,N_17929,N_17983);
and U18118 (N_18118,N_17998,N_17993);
or U18119 (N_18119,N_17868,N_17818);
nor U18120 (N_18120,N_17936,N_17981);
and U18121 (N_18121,N_17928,N_17936);
nor U18122 (N_18122,N_17973,N_17914);
and U18123 (N_18123,N_17957,N_17912);
or U18124 (N_18124,N_17898,N_17816);
nor U18125 (N_18125,N_17911,N_17941);
nand U18126 (N_18126,N_17935,N_17805);
nand U18127 (N_18127,N_17893,N_17989);
and U18128 (N_18128,N_17953,N_17805);
or U18129 (N_18129,N_17945,N_17809);
and U18130 (N_18130,N_17891,N_17847);
or U18131 (N_18131,N_17856,N_17921);
or U18132 (N_18132,N_17959,N_17980);
or U18133 (N_18133,N_17942,N_17971);
and U18134 (N_18134,N_17809,N_17925);
nand U18135 (N_18135,N_17820,N_17909);
nor U18136 (N_18136,N_17896,N_17867);
nor U18137 (N_18137,N_17825,N_17941);
nor U18138 (N_18138,N_17837,N_17980);
or U18139 (N_18139,N_17889,N_17861);
nand U18140 (N_18140,N_17809,N_17903);
nand U18141 (N_18141,N_17989,N_17899);
nand U18142 (N_18142,N_17939,N_17822);
or U18143 (N_18143,N_17975,N_17867);
or U18144 (N_18144,N_17921,N_17898);
or U18145 (N_18145,N_17818,N_17977);
nor U18146 (N_18146,N_17980,N_17885);
and U18147 (N_18147,N_17970,N_17835);
or U18148 (N_18148,N_17961,N_17876);
or U18149 (N_18149,N_17924,N_17805);
nand U18150 (N_18150,N_17823,N_17901);
nand U18151 (N_18151,N_17867,N_17988);
and U18152 (N_18152,N_17983,N_17944);
or U18153 (N_18153,N_17812,N_17846);
and U18154 (N_18154,N_17851,N_17805);
or U18155 (N_18155,N_17983,N_17962);
or U18156 (N_18156,N_17940,N_17845);
or U18157 (N_18157,N_17949,N_17884);
or U18158 (N_18158,N_17969,N_17995);
or U18159 (N_18159,N_17940,N_17867);
nand U18160 (N_18160,N_17832,N_17988);
nand U18161 (N_18161,N_17989,N_17810);
nor U18162 (N_18162,N_17813,N_17846);
nor U18163 (N_18163,N_17808,N_17998);
and U18164 (N_18164,N_17951,N_17898);
nor U18165 (N_18165,N_17833,N_17898);
nand U18166 (N_18166,N_17810,N_17953);
or U18167 (N_18167,N_17851,N_17901);
nor U18168 (N_18168,N_17964,N_17808);
nand U18169 (N_18169,N_17934,N_17973);
and U18170 (N_18170,N_17857,N_17960);
and U18171 (N_18171,N_17830,N_17973);
xnor U18172 (N_18172,N_17812,N_17833);
and U18173 (N_18173,N_17850,N_17801);
nand U18174 (N_18174,N_17910,N_17929);
nor U18175 (N_18175,N_17921,N_17933);
nor U18176 (N_18176,N_17889,N_17867);
nand U18177 (N_18177,N_17916,N_17832);
nor U18178 (N_18178,N_17851,N_17914);
or U18179 (N_18179,N_17814,N_17868);
and U18180 (N_18180,N_17814,N_17936);
and U18181 (N_18181,N_17847,N_17875);
nor U18182 (N_18182,N_17849,N_17872);
nor U18183 (N_18183,N_17859,N_17833);
nand U18184 (N_18184,N_17898,N_17890);
or U18185 (N_18185,N_17840,N_17947);
and U18186 (N_18186,N_17813,N_17908);
or U18187 (N_18187,N_17973,N_17982);
or U18188 (N_18188,N_17977,N_17828);
nand U18189 (N_18189,N_17903,N_17955);
nand U18190 (N_18190,N_17965,N_17992);
or U18191 (N_18191,N_17894,N_17994);
or U18192 (N_18192,N_17925,N_17960);
and U18193 (N_18193,N_17900,N_17975);
or U18194 (N_18194,N_17867,N_17826);
nor U18195 (N_18195,N_17889,N_17811);
and U18196 (N_18196,N_17824,N_17872);
nor U18197 (N_18197,N_17944,N_17919);
and U18198 (N_18198,N_17891,N_17976);
nor U18199 (N_18199,N_17998,N_17942);
and U18200 (N_18200,N_18179,N_18192);
nand U18201 (N_18201,N_18000,N_18075);
nand U18202 (N_18202,N_18188,N_18143);
nand U18203 (N_18203,N_18012,N_18044);
nand U18204 (N_18204,N_18017,N_18103);
or U18205 (N_18205,N_18057,N_18193);
and U18206 (N_18206,N_18168,N_18014);
nor U18207 (N_18207,N_18087,N_18151);
and U18208 (N_18208,N_18049,N_18113);
or U18209 (N_18209,N_18086,N_18079);
or U18210 (N_18210,N_18045,N_18165);
nand U18211 (N_18211,N_18154,N_18155);
nor U18212 (N_18212,N_18003,N_18195);
nand U18213 (N_18213,N_18080,N_18139);
and U18214 (N_18214,N_18136,N_18174);
and U18215 (N_18215,N_18076,N_18125);
or U18216 (N_18216,N_18041,N_18119);
and U18217 (N_18217,N_18043,N_18120);
nand U18218 (N_18218,N_18035,N_18163);
xnor U18219 (N_18219,N_18077,N_18110);
and U18220 (N_18220,N_18101,N_18009);
or U18221 (N_18221,N_18062,N_18095);
or U18222 (N_18222,N_18021,N_18112);
nand U18223 (N_18223,N_18169,N_18107);
or U18224 (N_18224,N_18197,N_18050);
and U18225 (N_18225,N_18097,N_18167);
nor U18226 (N_18226,N_18114,N_18130);
nor U18227 (N_18227,N_18156,N_18022);
or U18228 (N_18228,N_18088,N_18063);
nor U18229 (N_18229,N_18115,N_18127);
and U18230 (N_18230,N_18137,N_18019);
nand U18231 (N_18231,N_18160,N_18187);
or U18232 (N_18232,N_18198,N_18132);
nor U18233 (N_18233,N_18142,N_18084);
and U18234 (N_18234,N_18031,N_18164);
nor U18235 (N_18235,N_18007,N_18048);
nand U18236 (N_18236,N_18147,N_18189);
nand U18237 (N_18237,N_18094,N_18038);
or U18238 (N_18238,N_18129,N_18028);
nor U18239 (N_18239,N_18024,N_18148);
nor U18240 (N_18240,N_18046,N_18146);
nand U18241 (N_18241,N_18039,N_18191);
nor U18242 (N_18242,N_18020,N_18068);
nor U18243 (N_18243,N_18073,N_18074);
or U18244 (N_18244,N_18059,N_18099);
or U18245 (N_18245,N_18016,N_18036);
and U18246 (N_18246,N_18121,N_18047);
nor U18247 (N_18247,N_18054,N_18015);
xnor U18248 (N_18248,N_18173,N_18052);
nand U18249 (N_18249,N_18170,N_18064);
nand U18250 (N_18250,N_18051,N_18183);
and U18251 (N_18251,N_18098,N_18096);
nor U18252 (N_18252,N_18067,N_18199);
or U18253 (N_18253,N_18070,N_18141);
nor U18254 (N_18254,N_18030,N_18140);
or U18255 (N_18255,N_18008,N_18161);
or U18256 (N_18256,N_18056,N_18172);
nand U18257 (N_18257,N_18181,N_18069);
nand U18258 (N_18258,N_18032,N_18105);
nor U18259 (N_18259,N_18158,N_18134);
nor U18260 (N_18260,N_18128,N_18196);
or U18261 (N_18261,N_18033,N_18010);
or U18262 (N_18262,N_18018,N_18109);
or U18263 (N_18263,N_18133,N_18034);
and U18264 (N_18264,N_18006,N_18194);
and U18265 (N_18265,N_18058,N_18023);
and U18266 (N_18266,N_18144,N_18066);
or U18267 (N_18267,N_18124,N_18180);
or U18268 (N_18268,N_18159,N_18090);
nand U18269 (N_18269,N_18182,N_18004);
and U18270 (N_18270,N_18111,N_18190);
or U18271 (N_18271,N_18138,N_18001);
and U18272 (N_18272,N_18089,N_18011);
nor U18273 (N_18273,N_18152,N_18117);
nand U18274 (N_18274,N_18166,N_18027);
nand U18275 (N_18275,N_18175,N_18037);
nor U18276 (N_18276,N_18157,N_18185);
nand U18277 (N_18277,N_18072,N_18145);
and U18278 (N_18278,N_18065,N_18184);
nand U18279 (N_18279,N_18162,N_18093);
nand U18280 (N_18280,N_18153,N_18078);
nor U18281 (N_18281,N_18106,N_18013);
and U18282 (N_18282,N_18091,N_18186);
or U18283 (N_18283,N_18126,N_18150);
or U18284 (N_18284,N_18131,N_18082);
and U18285 (N_18285,N_18104,N_18040);
or U18286 (N_18286,N_18102,N_18177);
nand U18287 (N_18287,N_18071,N_18122);
nand U18288 (N_18288,N_18116,N_18092);
and U18289 (N_18289,N_18171,N_18100);
nor U18290 (N_18290,N_18108,N_18029);
and U18291 (N_18291,N_18123,N_18149);
nor U18292 (N_18292,N_18026,N_18176);
nor U18293 (N_18293,N_18081,N_18061);
and U18294 (N_18294,N_18135,N_18118);
nor U18295 (N_18295,N_18060,N_18005);
nand U18296 (N_18296,N_18055,N_18053);
or U18297 (N_18297,N_18042,N_18083);
or U18298 (N_18298,N_18085,N_18025);
or U18299 (N_18299,N_18002,N_18178);
nand U18300 (N_18300,N_18064,N_18171);
nor U18301 (N_18301,N_18123,N_18092);
or U18302 (N_18302,N_18021,N_18105);
nor U18303 (N_18303,N_18104,N_18058);
nand U18304 (N_18304,N_18095,N_18192);
or U18305 (N_18305,N_18066,N_18009);
nand U18306 (N_18306,N_18141,N_18154);
or U18307 (N_18307,N_18117,N_18026);
nor U18308 (N_18308,N_18086,N_18016);
and U18309 (N_18309,N_18027,N_18111);
or U18310 (N_18310,N_18055,N_18066);
or U18311 (N_18311,N_18130,N_18124);
nand U18312 (N_18312,N_18172,N_18068);
or U18313 (N_18313,N_18029,N_18100);
or U18314 (N_18314,N_18061,N_18151);
and U18315 (N_18315,N_18141,N_18161);
nor U18316 (N_18316,N_18027,N_18155);
and U18317 (N_18317,N_18117,N_18124);
nor U18318 (N_18318,N_18021,N_18090);
or U18319 (N_18319,N_18037,N_18132);
or U18320 (N_18320,N_18121,N_18042);
nand U18321 (N_18321,N_18002,N_18135);
nand U18322 (N_18322,N_18022,N_18080);
and U18323 (N_18323,N_18019,N_18100);
or U18324 (N_18324,N_18121,N_18007);
nor U18325 (N_18325,N_18059,N_18012);
or U18326 (N_18326,N_18062,N_18154);
and U18327 (N_18327,N_18138,N_18116);
nand U18328 (N_18328,N_18105,N_18022);
nor U18329 (N_18329,N_18082,N_18101);
nand U18330 (N_18330,N_18041,N_18142);
nand U18331 (N_18331,N_18074,N_18142);
and U18332 (N_18332,N_18029,N_18121);
or U18333 (N_18333,N_18127,N_18174);
nand U18334 (N_18334,N_18156,N_18139);
or U18335 (N_18335,N_18025,N_18189);
nand U18336 (N_18336,N_18014,N_18117);
nor U18337 (N_18337,N_18041,N_18031);
nand U18338 (N_18338,N_18023,N_18180);
nand U18339 (N_18339,N_18133,N_18097);
or U18340 (N_18340,N_18134,N_18005);
or U18341 (N_18341,N_18007,N_18011);
and U18342 (N_18342,N_18045,N_18057);
nand U18343 (N_18343,N_18073,N_18098);
and U18344 (N_18344,N_18175,N_18070);
nand U18345 (N_18345,N_18182,N_18082);
or U18346 (N_18346,N_18163,N_18066);
or U18347 (N_18347,N_18039,N_18012);
or U18348 (N_18348,N_18092,N_18018);
nor U18349 (N_18349,N_18139,N_18000);
or U18350 (N_18350,N_18113,N_18082);
nor U18351 (N_18351,N_18070,N_18061);
or U18352 (N_18352,N_18065,N_18121);
nor U18353 (N_18353,N_18154,N_18189);
nand U18354 (N_18354,N_18028,N_18067);
nor U18355 (N_18355,N_18076,N_18135);
and U18356 (N_18356,N_18120,N_18046);
and U18357 (N_18357,N_18083,N_18073);
nand U18358 (N_18358,N_18094,N_18129);
and U18359 (N_18359,N_18125,N_18175);
and U18360 (N_18360,N_18056,N_18181);
nand U18361 (N_18361,N_18029,N_18061);
nor U18362 (N_18362,N_18151,N_18124);
or U18363 (N_18363,N_18176,N_18084);
or U18364 (N_18364,N_18104,N_18010);
nor U18365 (N_18365,N_18099,N_18046);
nand U18366 (N_18366,N_18130,N_18041);
nor U18367 (N_18367,N_18176,N_18044);
or U18368 (N_18368,N_18102,N_18077);
nand U18369 (N_18369,N_18191,N_18030);
or U18370 (N_18370,N_18035,N_18039);
nor U18371 (N_18371,N_18024,N_18091);
and U18372 (N_18372,N_18083,N_18167);
and U18373 (N_18373,N_18116,N_18022);
nand U18374 (N_18374,N_18189,N_18008);
nor U18375 (N_18375,N_18060,N_18105);
nand U18376 (N_18376,N_18144,N_18178);
nand U18377 (N_18377,N_18096,N_18040);
and U18378 (N_18378,N_18163,N_18175);
or U18379 (N_18379,N_18155,N_18011);
nor U18380 (N_18380,N_18182,N_18113);
and U18381 (N_18381,N_18056,N_18148);
or U18382 (N_18382,N_18078,N_18101);
and U18383 (N_18383,N_18160,N_18094);
nor U18384 (N_18384,N_18144,N_18198);
nor U18385 (N_18385,N_18059,N_18009);
or U18386 (N_18386,N_18190,N_18169);
or U18387 (N_18387,N_18050,N_18106);
or U18388 (N_18388,N_18048,N_18029);
nand U18389 (N_18389,N_18092,N_18181);
and U18390 (N_18390,N_18157,N_18005);
nand U18391 (N_18391,N_18107,N_18052);
and U18392 (N_18392,N_18140,N_18073);
and U18393 (N_18393,N_18056,N_18018);
nor U18394 (N_18394,N_18034,N_18171);
nand U18395 (N_18395,N_18015,N_18151);
or U18396 (N_18396,N_18122,N_18035);
and U18397 (N_18397,N_18113,N_18054);
and U18398 (N_18398,N_18088,N_18156);
and U18399 (N_18399,N_18129,N_18089);
nand U18400 (N_18400,N_18237,N_18269);
or U18401 (N_18401,N_18333,N_18305);
or U18402 (N_18402,N_18255,N_18208);
and U18403 (N_18403,N_18320,N_18213);
or U18404 (N_18404,N_18304,N_18284);
and U18405 (N_18405,N_18245,N_18279);
nand U18406 (N_18406,N_18234,N_18392);
or U18407 (N_18407,N_18293,N_18277);
and U18408 (N_18408,N_18314,N_18313);
nor U18409 (N_18409,N_18387,N_18311);
and U18410 (N_18410,N_18356,N_18306);
nand U18411 (N_18411,N_18334,N_18246);
or U18412 (N_18412,N_18384,N_18330);
or U18413 (N_18413,N_18324,N_18364);
and U18414 (N_18414,N_18357,N_18201);
and U18415 (N_18415,N_18270,N_18256);
and U18416 (N_18416,N_18217,N_18244);
or U18417 (N_18417,N_18276,N_18362);
nor U18418 (N_18418,N_18302,N_18210);
or U18419 (N_18419,N_18370,N_18315);
or U18420 (N_18420,N_18274,N_18229);
and U18421 (N_18421,N_18369,N_18321);
nand U18422 (N_18422,N_18331,N_18233);
or U18423 (N_18423,N_18204,N_18212);
nor U18424 (N_18424,N_18346,N_18242);
or U18425 (N_18425,N_18398,N_18254);
nor U18426 (N_18426,N_18281,N_18259);
or U18427 (N_18427,N_18375,N_18264);
or U18428 (N_18428,N_18211,N_18286);
nor U18429 (N_18429,N_18382,N_18273);
nor U18430 (N_18430,N_18235,N_18263);
or U18431 (N_18431,N_18253,N_18261);
and U18432 (N_18432,N_18338,N_18348);
or U18433 (N_18433,N_18266,N_18345);
nor U18434 (N_18434,N_18301,N_18395);
and U18435 (N_18435,N_18388,N_18258);
or U18436 (N_18436,N_18354,N_18223);
nand U18437 (N_18437,N_18206,N_18230);
nor U18438 (N_18438,N_18372,N_18294);
and U18439 (N_18439,N_18241,N_18252);
or U18440 (N_18440,N_18290,N_18226);
nand U18441 (N_18441,N_18296,N_18232);
nor U18442 (N_18442,N_18272,N_18355);
and U18443 (N_18443,N_18215,N_18365);
and U18444 (N_18444,N_18291,N_18216);
nand U18445 (N_18445,N_18358,N_18238);
nand U18446 (N_18446,N_18374,N_18275);
and U18447 (N_18447,N_18295,N_18225);
and U18448 (N_18448,N_18312,N_18366);
nor U18449 (N_18449,N_18396,N_18247);
and U18450 (N_18450,N_18318,N_18342);
or U18451 (N_18451,N_18373,N_18227);
nor U18452 (N_18452,N_18250,N_18379);
nor U18453 (N_18453,N_18383,N_18202);
nand U18454 (N_18454,N_18271,N_18260);
nor U18455 (N_18455,N_18323,N_18361);
or U18456 (N_18456,N_18205,N_18298);
nor U18457 (N_18457,N_18267,N_18359);
or U18458 (N_18458,N_18310,N_18278);
and U18459 (N_18459,N_18220,N_18282);
nand U18460 (N_18460,N_18343,N_18292);
nor U18461 (N_18461,N_18283,N_18380);
or U18462 (N_18462,N_18236,N_18265);
nor U18463 (N_18463,N_18397,N_18371);
or U18464 (N_18464,N_18329,N_18309);
and U18465 (N_18465,N_18337,N_18399);
or U18466 (N_18466,N_18390,N_18353);
and U18467 (N_18467,N_18207,N_18228);
or U18468 (N_18468,N_18288,N_18325);
or U18469 (N_18469,N_18221,N_18249);
and U18470 (N_18470,N_18341,N_18287);
or U18471 (N_18471,N_18209,N_18391);
or U18472 (N_18472,N_18386,N_18239);
nand U18473 (N_18473,N_18214,N_18332);
nor U18474 (N_18474,N_18376,N_18200);
or U18475 (N_18475,N_18367,N_18335);
or U18476 (N_18476,N_18300,N_18339);
nand U18477 (N_18477,N_18240,N_18381);
nand U18478 (N_18478,N_18297,N_18385);
nand U18479 (N_18479,N_18307,N_18319);
nand U18480 (N_18480,N_18243,N_18317);
and U18481 (N_18481,N_18350,N_18248);
or U18482 (N_18482,N_18360,N_18378);
nand U18483 (N_18483,N_18219,N_18336);
nand U18484 (N_18484,N_18280,N_18328);
nand U18485 (N_18485,N_18262,N_18347);
or U18486 (N_18486,N_18368,N_18285);
nand U18487 (N_18487,N_18231,N_18389);
and U18488 (N_18488,N_18257,N_18251);
nor U18489 (N_18489,N_18349,N_18393);
and U18490 (N_18490,N_18299,N_18222);
or U18491 (N_18491,N_18352,N_18322);
nand U18492 (N_18492,N_18327,N_18394);
or U18493 (N_18493,N_18351,N_18308);
nand U18494 (N_18494,N_18316,N_18340);
nor U18495 (N_18495,N_18224,N_18363);
and U18496 (N_18496,N_18289,N_18344);
nand U18497 (N_18497,N_18326,N_18203);
nor U18498 (N_18498,N_18303,N_18268);
nand U18499 (N_18499,N_18218,N_18377);
nor U18500 (N_18500,N_18399,N_18218);
nand U18501 (N_18501,N_18367,N_18219);
nor U18502 (N_18502,N_18249,N_18344);
nand U18503 (N_18503,N_18315,N_18275);
nor U18504 (N_18504,N_18381,N_18347);
nor U18505 (N_18505,N_18213,N_18307);
nor U18506 (N_18506,N_18290,N_18214);
and U18507 (N_18507,N_18397,N_18214);
or U18508 (N_18508,N_18310,N_18205);
nand U18509 (N_18509,N_18240,N_18397);
or U18510 (N_18510,N_18332,N_18204);
nand U18511 (N_18511,N_18214,N_18342);
or U18512 (N_18512,N_18370,N_18247);
xnor U18513 (N_18513,N_18226,N_18250);
and U18514 (N_18514,N_18286,N_18356);
nor U18515 (N_18515,N_18348,N_18367);
and U18516 (N_18516,N_18306,N_18376);
and U18517 (N_18517,N_18201,N_18352);
nor U18518 (N_18518,N_18323,N_18345);
and U18519 (N_18519,N_18327,N_18204);
or U18520 (N_18520,N_18208,N_18358);
nor U18521 (N_18521,N_18315,N_18287);
nand U18522 (N_18522,N_18271,N_18394);
and U18523 (N_18523,N_18359,N_18329);
or U18524 (N_18524,N_18232,N_18270);
or U18525 (N_18525,N_18319,N_18299);
nand U18526 (N_18526,N_18215,N_18256);
nor U18527 (N_18527,N_18297,N_18353);
nor U18528 (N_18528,N_18295,N_18229);
nand U18529 (N_18529,N_18381,N_18277);
or U18530 (N_18530,N_18329,N_18336);
xor U18531 (N_18531,N_18250,N_18213);
or U18532 (N_18532,N_18286,N_18284);
nand U18533 (N_18533,N_18244,N_18321);
nor U18534 (N_18534,N_18251,N_18333);
nor U18535 (N_18535,N_18268,N_18301);
nor U18536 (N_18536,N_18392,N_18240);
or U18537 (N_18537,N_18226,N_18291);
and U18538 (N_18538,N_18377,N_18212);
and U18539 (N_18539,N_18211,N_18229);
nor U18540 (N_18540,N_18332,N_18242);
nor U18541 (N_18541,N_18326,N_18332);
and U18542 (N_18542,N_18278,N_18301);
nand U18543 (N_18543,N_18398,N_18376);
and U18544 (N_18544,N_18328,N_18275);
and U18545 (N_18545,N_18392,N_18365);
or U18546 (N_18546,N_18271,N_18216);
and U18547 (N_18547,N_18289,N_18273);
or U18548 (N_18548,N_18394,N_18286);
nor U18549 (N_18549,N_18358,N_18218);
or U18550 (N_18550,N_18220,N_18358);
nor U18551 (N_18551,N_18203,N_18363);
and U18552 (N_18552,N_18224,N_18387);
nor U18553 (N_18553,N_18389,N_18296);
or U18554 (N_18554,N_18336,N_18364);
nand U18555 (N_18555,N_18345,N_18319);
and U18556 (N_18556,N_18284,N_18258);
nand U18557 (N_18557,N_18298,N_18268);
nand U18558 (N_18558,N_18388,N_18307);
or U18559 (N_18559,N_18304,N_18376);
and U18560 (N_18560,N_18242,N_18223);
nand U18561 (N_18561,N_18351,N_18220);
nand U18562 (N_18562,N_18277,N_18383);
nor U18563 (N_18563,N_18232,N_18234);
nor U18564 (N_18564,N_18282,N_18344);
or U18565 (N_18565,N_18240,N_18258);
or U18566 (N_18566,N_18279,N_18344);
nand U18567 (N_18567,N_18370,N_18331);
nor U18568 (N_18568,N_18334,N_18224);
nor U18569 (N_18569,N_18238,N_18295);
nor U18570 (N_18570,N_18301,N_18394);
and U18571 (N_18571,N_18247,N_18232);
and U18572 (N_18572,N_18327,N_18373);
or U18573 (N_18573,N_18260,N_18203);
nor U18574 (N_18574,N_18391,N_18229);
nor U18575 (N_18575,N_18223,N_18356);
and U18576 (N_18576,N_18327,N_18336);
and U18577 (N_18577,N_18250,N_18252);
nor U18578 (N_18578,N_18370,N_18364);
and U18579 (N_18579,N_18221,N_18370);
nor U18580 (N_18580,N_18321,N_18283);
or U18581 (N_18581,N_18311,N_18396);
nor U18582 (N_18582,N_18315,N_18269);
and U18583 (N_18583,N_18389,N_18289);
or U18584 (N_18584,N_18306,N_18355);
nor U18585 (N_18585,N_18387,N_18288);
or U18586 (N_18586,N_18295,N_18279);
or U18587 (N_18587,N_18303,N_18315);
or U18588 (N_18588,N_18200,N_18222);
nand U18589 (N_18589,N_18387,N_18270);
and U18590 (N_18590,N_18278,N_18230);
nand U18591 (N_18591,N_18251,N_18235);
nand U18592 (N_18592,N_18222,N_18313);
nor U18593 (N_18593,N_18339,N_18249);
or U18594 (N_18594,N_18359,N_18360);
nor U18595 (N_18595,N_18313,N_18348);
and U18596 (N_18596,N_18356,N_18314);
and U18597 (N_18597,N_18255,N_18342);
and U18598 (N_18598,N_18368,N_18206);
and U18599 (N_18599,N_18304,N_18267);
nor U18600 (N_18600,N_18421,N_18512);
nor U18601 (N_18601,N_18490,N_18558);
nor U18602 (N_18602,N_18483,N_18590);
nand U18603 (N_18603,N_18419,N_18426);
or U18604 (N_18604,N_18442,N_18538);
or U18605 (N_18605,N_18561,N_18433);
nand U18606 (N_18606,N_18533,N_18551);
or U18607 (N_18607,N_18539,N_18534);
nor U18608 (N_18608,N_18581,N_18436);
xor U18609 (N_18609,N_18573,N_18530);
or U18610 (N_18610,N_18544,N_18477);
and U18611 (N_18611,N_18423,N_18487);
nand U18612 (N_18612,N_18552,N_18464);
or U18613 (N_18613,N_18452,N_18574);
nor U18614 (N_18614,N_18577,N_18567);
and U18615 (N_18615,N_18536,N_18566);
and U18616 (N_18616,N_18444,N_18473);
nor U18617 (N_18617,N_18499,N_18402);
nor U18618 (N_18618,N_18410,N_18559);
or U18619 (N_18619,N_18470,N_18424);
nor U18620 (N_18620,N_18493,N_18523);
nor U18621 (N_18621,N_18441,N_18593);
or U18622 (N_18622,N_18443,N_18463);
xnor U18623 (N_18623,N_18511,N_18518);
and U18624 (N_18624,N_18492,N_18554);
nand U18625 (N_18625,N_18506,N_18411);
nor U18626 (N_18626,N_18589,N_18471);
xor U18627 (N_18627,N_18501,N_18446);
and U18628 (N_18628,N_18569,N_18570);
nor U18629 (N_18629,N_18595,N_18422);
or U18630 (N_18630,N_18549,N_18434);
nand U18631 (N_18631,N_18472,N_18562);
and U18632 (N_18632,N_18578,N_18481);
nor U18633 (N_18633,N_18435,N_18404);
or U18634 (N_18634,N_18458,N_18405);
or U18635 (N_18635,N_18479,N_18502);
or U18636 (N_18636,N_18427,N_18572);
nand U18637 (N_18637,N_18548,N_18579);
or U18638 (N_18638,N_18594,N_18571);
or U18639 (N_18639,N_18505,N_18556);
or U18640 (N_18640,N_18503,N_18488);
nor U18641 (N_18641,N_18519,N_18460);
or U18642 (N_18642,N_18508,N_18555);
nand U18643 (N_18643,N_18430,N_18517);
nor U18644 (N_18644,N_18486,N_18532);
nor U18645 (N_18645,N_18409,N_18510);
or U18646 (N_18646,N_18489,N_18575);
nand U18647 (N_18647,N_18412,N_18513);
and U18648 (N_18648,N_18531,N_18437);
or U18649 (N_18649,N_18408,N_18540);
and U18650 (N_18650,N_18432,N_18583);
and U18651 (N_18651,N_18485,N_18468);
nor U18652 (N_18652,N_18401,N_18557);
nor U18653 (N_18653,N_18529,N_18495);
nor U18654 (N_18654,N_18445,N_18484);
or U18655 (N_18655,N_18521,N_18456);
or U18656 (N_18656,N_18415,N_18465);
or U18657 (N_18657,N_18429,N_18466);
and U18658 (N_18658,N_18497,N_18550);
or U18659 (N_18659,N_18565,N_18448);
or U18660 (N_18660,N_18447,N_18407);
or U18661 (N_18661,N_18564,N_18537);
nor U18662 (N_18662,N_18449,N_18599);
and U18663 (N_18663,N_18450,N_18509);
nor U18664 (N_18664,N_18475,N_18563);
and U18665 (N_18665,N_18568,N_18597);
and U18666 (N_18666,N_18469,N_18526);
nand U18667 (N_18667,N_18461,N_18428);
nor U18668 (N_18668,N_18507,N_18462);
or U18669 (N_18669,N_18416,N_18520);
or U18670 (N_18670,N_18586,N_18431);
or U18671 (N_18671,N_18582,N_18482);
nor U18672 (N_18672,N_18584,N_18496);
nand U18673 (N_18673,N_18474,N_18498);
or U18674 (N_18674,N_18553,N_18494);
nand U18675 (N_18675,N_18400,N_18504);
and U18676 (N_18676,N_18535,N_18587);
nand U18677 (N_18677,N_18545,N_18453);
and U18678 (N_18678,N_18455,N_18560);
nand U18679 (N_18679,N_18591,N_18598);
or U18680 (N_18680,N_18547,N_18528);
nor U18681 (N_18681,N_18438,N_18525);
and U18682 (N_18682,N_18515,N_18585);
and U18683 (N_18683,N_18457,N_18440);
nand U18684 (N_18684,N_18418,N_18524);
nor U18685 (N_18685,N_18514,N_18454);
and U18686 (N_18686,N_18451,N_18500);
nand U18687 (N_18687,N_18527,N_18576);
or U18688 (N_18688,N_18596,N_18420);
or U18689 (N_18689,N_18480,N_18425);
nor U18690 (N_18690,N_18476,N_18459);
nand U18691 (N_18691,N_18522,N_18417);
or U18692 (N_18692,N_18414,N_18467);
nand U18693 (N_18693,N_18580,N_18413);
or U18694 (N_18694,N_18516,N_18541);
nor U18695 (N_18695,N_18588,N_18439);
or U18696 (N_18696,N_18546,N_18478);
or U18697 (N_18697,N_18403,N_18543);
and U18698 (N_18698,N_18542,N_18592);
nand U18699 (N_18699,N_18406,N_18491);
nand U18700 (N_18700,N_18444,N_18575);
xnor U18701 (N_18701,N_18545,N_18428);
nor U18702 (N_18702,N_18401,N_18476);
nor U18703 (N_18703,N_18551,N_18475);
nand U18704 (N_18704,N_18507,N_18556);
and U18705 (N_18705,N_18518,N_18559);
and U18706 (N_18706,N_18573,N_18457);
nor U18707 (N_18707,N_18476,N_18580);
or U18708 (N_18708,N_18402,N_18519);
nand U18709 (N_18709,N_18588,N_18448);
and U18710 (N_18710,N_18540,N_18497);
and U18711 (N_18711,N_18501,N_18477);
and U18712 (N_18712,N_18542,N_18554);
nand U18713 (N_18713,N_18430,N_18453);
nand U18714 (N_18714,N_18512,N_18409);
nand U18715 (N_18715,N_18525,N_18557);
nor U18716 (N_18716,N_18439,N_18488);
nor U18717 (N_18717,N_18521,N_18545);
and U18718 (N_18718,N_18572,N_18547);
and U18719 (N_18719,N_18447,N_18436);
or U18720 (N_18720,N_18404,N_18460);
nand U18721 (N_18721,N_18422,N_18437);
nor U18722 (N_18722,N_18515,N_18531);
or U18723 (N_18723,N_18496,N_18593);
nand U18724 (N_18724,N_18479,N_18547);
and U18725 (N_18725,N_18426,N_18502);
nor U18726 (N_18726,N_18404,N_18447);
or U18727 (N_18727,N_18541,N_18460);
and U18728 (N_18728,N_18449,N_18403);
and U18729 (N_18729,N_18441,N_18486);
or U18730 (N_18730,N_18470,N_18536);
and U18731 (N_18731,N_18530,N_18455);
and U18732 (N_18732,N_18518,N_18548);
or U18733 (N_18733,N_18557,N_18461);
nor U18734 (N_18734,N_18443,N_18552);
nand U18735 (N_18735,N_18482,N_18492);
and U18736 (N_18736,N_18520,N_18538);
and U18737 (N_18737,N_18493,N_18471);
or U18738 (N_18738,N_18548,N_18409);
and U18739 (N_18739,N_18526,N_18595);
or U18740 (N_18740,N_18427,N_18544);
nor U18741 (N_18741,N_18516,N_18511);
and U18742 (N_18742,N_18540,N_18441);
or U18743 (N_18743,N_18421,N_18540);
nand U18744 (N_18744,N_18537,N_18558);
xnor U18745 (N_18745,N_18518,N_18496);
nor U18746 (N_18746,N_18404,N_18551);
or U18747 (N_18747,N_18476,N_18565);
nand U18748 (N_18748,N_18487,N_18580);
nand U18749 (N_18749,N_18402,N_18494);
and U18750 (N_18750,N_18427,N_18431);
and U18751 (N_18751,N_18468,N_18438);
and U18752 (N_18752,N_18520,N_18573);
nor U18753 (N_18753,N_18475,N_18598);
and U18754 (N_18754,N_18555,N_18559);
nand U18755 (N_18755,N_18538,N_18569);
nor U18756 (N_18756,N_18467,N_18527);
nand U18757 (N_18757,N_18457,N_18460);
nor U18758 (N_18758,N_18422,N_18474);
or U18759 (N_18759,N_18415,N_18466);
and U18760 (N_18760,N_18554,N_18471);
or U18761 (N_18761,N_18560,N_18436);
xnor U18762 (N_18762,N_18509,N_18586);
nor U18763 (N_18763,N_18403,N_18445);
or U18764 (N_18764,N_18598,N_18463);
and U18765 (N_18765,N_18597,N_18435);
nor U18766 (N_18766,N_18448,N_18402);
nand U18767 (N_18767,N_18586,N_18467);
and U18768 (N_18768,N_18542,N_18585);
nand U18769 (N_18769,N_18474,N_18581);
and U18770 (N_18770,N_18553,N_18438);
and U18771 (N_18771,N_18416,N_18430);
nand U18772 (N_18772,N_18443,N_18405);
or U18773 (N_18773,N_18409,N_18418);
nand U18774 (N_18774,N_18585,N_18521);
and U18775 (N_18775,N_18528,N_18581);
nor U18776 (N_18776,N_18532,N_18475);
nand U18777 (N_18777,N_18515,N_18424);
or U18778 (N_18778,N_18578,N_18553);
nand U18779 (N_18779,N_18418,N_18460);
nor U18780 (N_18780,N_18466,N_18583);
nor U18781 (N_18781,N_18457,N_18491);
and U18782 (N_18782,N_18520,N_18553);
nor U18783 (N_18783,N_18428,N_18476);
nand U18784 (N_18784,N_18483,N_18542);
nand U18785 (N_18785,N_18537,N_18431);
or U18786 (N_18786,N_18581,N_18599);
or U18787 (N_18787,N_18559,N_18437);
nor U18788 (N_18788,N_18484,N_18595);
nor U18789 (N_18789,N_18499,N_18519);
and U18790 (N_18790,N_18516,N_18535);
and U18791 (N_18791,N_18464,N_18577);
and U18792 (N_18792,N_18461,N_18497);
nand U18793 (N_18793,N_18591,N_18489);
and U18794 (N_18794,N_18467,N_18564);
nor U18795 (N_18795,N_18452,N_18404);
and U18796 (N_18796,N_18555,N_18492);
and U18797 (N_18797,N_18402,N_18405);
or U18798 (N_18798,N_18519,N_18406);
or U18799 (N_18799,N_18465,N_18481);
and U18800 (N_18800,N_18735,N_18694);
or U18801 (N_18801,N_18744,N_18747);
or U18802 (N_18802,N_18678,N_18793);
nor U18803 (N_18803,N_18654,N_18635);
nand U18804 (N_18804,N_18755,N_18788);
nand U18805 (N_18805,N_18682,N_18787);
or U18806 (N_18806,N_18776,N_18783);
nor U18807 (N_18807,N_18731,N_18690);
and U18808 (N_18808,N_18688,N_18664);
or U18809 (N_18809,N_18626,N_18612);
nand U18810 (N_18810,N_18738,N_18695);
nand U18811 (N_18811,N_18679,N_18666);
nor U18812 (N_18812,N_18657,N_18624);
or U18813 (N_18813,N_18729,N_18725);
and U18814 (N_18814,N_18683,N_18702);
and U18815 (N_18815,N_18705,N_18633);
and U18816 (N_18816,N_18677,N_18641);
nor U18817 (N_18817,N_18645,N_18711);
or U18818 (N_18818,N_18704,N_18734);
nor U18819 (N_18819,N_18648,N_18797);
nor U18820 (N_18820,N_18775,N_18622);
nand U18821 (N_18821,N_18779,N_18650);
or U18822 (N_18822,N_18617,N_18600);
or U18823 (N_18823,N_18728,N_18651);
and U18824 (N_18824,N_18615,N_18699);
or U18825 (N_18825,N_18778,N_18609);
and U18826 (N_18826,N_18748,N_18760);
nor U18827 (N_18827,N_18685,N_18662);
and U18828 (N_18828,N_18659,N_18669);
and U18829 (N_18829,N_18630,N_18764);
nor U18830 (N_18830,N_18637,N_18723);
nor U18831 (N_18831,N_18716,N_18799);
nor U18832 (N_18832,N_18647,N_18753);
nor U18833 (N_18833,N_18717,N_18674);
nor U18834 (N_18834,N_18608,N_18741);
or U18835 (N_18835,N_18710,N_18649);
nand U18836 (N_18836,N_18634,N_18794);
nand U18837 (N_18837,N_18743,N_18684);
nor U18838 (N_18838,N_18767,N_18675);
nor U18839 (N_18839,N_18707,N_18642);
nand U18840 (N_18840,N_18605,N_18719);
nand U18841 (N_18841,N_18713,N_18696);
nor U18842 (N_18842,N_18698,N_18620);
and U18843 (N_18843,N_18602,N_18757);
nor U18844 (N_18844,N_18610,N_18692);
nor U18845 (N_18845,N_18661,N_18606);
nor U18846 (N_18846,N_18780,N_18715);
and U18847 (N_18847,N_18724,N_18680);
nand U18848 (N_18848,N_18795,N_18756);
or U18849 (N_18849,N_18751,N_18709);
and U18850 (N_18850,N_18623,N_18613);
nor U18851 (N_18851,N_18639,N_18737);
nand U18852 (N_18852,N_18646,N_18625);
nor U18853 (N_18853,N_18644,N_18718);
nor U18854 (N_18854,N_18628,N_18730);
nand U18855 (N_18855,N_18643,N_18672);
and U18856 (N_18856,N_18660,N_18722);
and U18857 (N_18857,N_18604,N_18771);
nor U18858 (N_18858,N_18784,N_18763);
or U18859 (N_18859,N_18786,N_18790);
or U18860 (N_18860,N_18614,N_18652);
and U18861 (N_18861,N_18703,N_18673);
nand U18862 (N_18862,N_18720,N_18670);
or U18863 (N_18863,N_18700,N_18706);
xor U18864 (N_18864,N_18754,N_18691);
and U18865 (N_18865,N_18712,N_18750);
nor U18866 (N_18866,N_18777,N_18689);
and U18867 (N_18867,N_18714,N_18655);
or U18868 (N_18868,N_18621,N_18785);
and U18869 (N_18869,N_18721,N_18619);
or U18870 (N_18870,N_18761,N_18727);
or U18871 (N_18871,N_18726,N_18640);
nor U18872 (N_18872,N_18789,N_18616);
nor U18873 (N_18873,N_18631,N_18758);
or U18874 (N_18874,N_18671,N_18638);
or U18875 (N_18875,N_18782,N_18796);
nor U18876 (N_18876,N_18676,N_18627);
nand U18877 (N_18877,N_18740,N_18601);
nand U18878 (N_18878,N_18749,N_18629);
and U18879 (N_18879,N_18769,N_18687);
nand U18880 (N_18880,N_18658,N_18762);
or U18881 (N_18881,N_18791,N_18632);
nand U18882 (N_18882,N_18752,N_18736);
or U18883 (N_18883,N_18697,N_18607);
nand U18884 (N_18884,N_18745,N_18611);
nand U18885 (N_18885,N_18781,N_18770);
nor U18886 (N_18886,N_18746,N_18618);
or U18887 (N_18887,N_18739,N_18668);
nand U18888 (N_18888,N_18774,N_18732);
and U18889 (N_18889,N_18693,N_18759);
nand U18890 (N_18890,N_18765,N_18773);
and U18891 (N_18891,N_18603,N_18667);
nor U18892 (N_18892,N_18742,N_18708);
nor U18893 (N_18893,N_18798,N_18681);
or U18894 (N_18894,N_18653,N_18656);
and U18895 (N_18895,N_18768,N_18665);
nand U18896 (N_18896,N_18686,N_18772);
nor U18897 (N_18897,N_18701,N_18792);
nand U18898 (N_18898,N_18766,N_18733);
nor U18899 (N_18899,N_18636,N_18663);
nor U18900 (N_18900,N_18791,N_18647);
and U18901 (N_18901,N_18683,N_18716);
and U18902 (N_18902,N_18736,N_18600);
and U18903 (N_18903,N_18752,N_18648);
or U18904 (N_18904,N_18627,N_18601);
and U18905 (N_18905,N_18614,N_18690);
and U18906 (N_18906,N_18629,N_18651);
nor U18907 (N_18907,N_18613,N_18669);
and U18908 (N_18908,N_18704,N_18788);
nor U18909 (N_18909,N_18639,N_18610);
nand U18910 (N_18910,N_18741,N_18691);
nor U18911 (N_18911,N_18795,N_18787);
nand U18912 (N_18912,N_18707,N_18725);
nand U18913 (N_18913,N_18689,N_18631);
nor U18914 (N_18914,N_18679,N_18691);
nor U18915 (N_18915,N_18654,N_18629);
or U18916 (N_18916,N_18740,N_18693);
or U18917 (N_18917,N_18726,N_18671);
and U18918 (N_18918,N_18681,N_18706);
nor U18919 (N_18919,N_18738,N_18645);
or U18920 (N_18920,N_18680,N_18761);
or U18921 (N_18921,N_18779,N_18720);
nand U18922 (N_18922,N_18772,N_18746);
nand U18923 (N_18923,N_18729,N_18684);
nand U18924 (N_18924,N_18752,N_18764);
nor U18925 (N_18925,N_18657,N_18656);
or U18926 (N_18926,N_18770,N_18752);
nand U18927 (N_18927,N_18659,N_18648);
or U18928 (N_18928,N_18744,N_18659);
or U18929 (N_18929,N_18609,N_18699);
nand U18930 (N_18930,N_18715,N_18632);
nor U18931 (N_18931,N_18701,N_18642);
and U18932 (N_18932,N_18716,N_18784);
nand U18933 (N_18933,N_18628,N_18624);
nor U18934 (N_18934,N_18783,N_18762);
nand U18935 (N_18935,N_18606,N_18752);
and U18936 (N_18936,N_18681,N_18657);
or U18937 (N_18937,N_18718,N_18716);
nor U18938 (N_18938,N_18680,N_18627);
nor U18939 (N_18939,N_18698,N_18794);
nor U18940 (N_18940,N_18643,N_18654);
or U18941 (N_18941,N_18653,N_18679);
nand U18942 (N_18942,N_18636,N_18775);
or U18943 (N_18943,N_18666,N_18756);
nor U18944 (N_18944,N_18748,N_18763);
nand U18945 (N_18945,N_18615,N_18679);
xnor U18946 (N_18946,N_18766,N_18719);
nand U18947 (N_18947,N_18635,N_18605);
nand U18948 (N_18948,N_18746,N_18792);
nand U18949 (N_18949,N_18790,N_18683);
nor U18950 (N_18950,N_18724,N_18760);
nor U18951 (N_18951,N_18699,N_18772);
nand U18952 (N_18952,N_18668,N_18606);
and U18953 (N_18953,N_18788,N_18715);
nor U18954 (N_18954,N_18784,N_18633);
or U18955 (N_18955,N_18758,N_18797);
nand U18956 (N_18956,N_18629,N_18763);
or U18957 (N_18957,N_18636,N_18667);
nor U18958 (N_18958,N_18700,N_18790);
and U18959 (N_18959,N_18723,N_18796);
nor U18960 (N_18960,N_18622,N_18668);
or U18961 (N_18961,N_18732,N_18656);
and U18962 (N_18962,N_18724,N_18727);
nand U18963 (N_18963,N_18754,N_18695);
or U18964 (N_18964,N_18615,N_18603);
or U18965 (N_18965,N_18609,N_18695);
nor U18966 (N_18966,N_18749,N_18706);
nand U18967 (N_18967,N_18792,N_18627);
nand U18968 (N_18968,N_18752,N_18688);
xor U18969 (N_18969,N_18647,N_18601);
and U18970 (N_18970,N_18784,N_18758);
or U18971 (N_18971,N_18659,N_18730);
nand U18972 (N_18972,N_18791,N_18792);
nand U18973 (N_18973,N_18774,N_18785);
or U18974 (N_18974,N_18628,N_18738);
or U18975 (N_18975,N_18613,N_18608);
and U18976 (N_18976,N_18718,N_18628);
nand U18977 (N_18977,N_18701,N_18743);
or U18978 (N_18978,N_18658,N_18654);
and U18979 (N_18979,N_18629,N_18637);
or U18980 (N_18980,N_18638,N_18643);
nor U18981 (N_18981,N_18781,N_18741);
and U18982 (N_18982,N_18691,N_18633);
nor U18983 (N_18983,N_18739,N_18655);
nand U18984 (N_18984,N_18661,N_18748);
nand U18985 (N_18985,N_18751,N_18734);
and U18986 (N_18986,N_18726,N_18601);
nand U18987 (N_18987,N_18754,N_18790);
or U18988 (N_18988,N_18606,N_18749);
nor U18989 (N_18989,N_18787,N_18656);
nand U18990 (N_18990,N_18620,N_18622);
nand U18991 (N_18991,N_18770,N_18662);
nor U18992 (N_18992,N_18635,N_18742);
nor U18993 (N_18993,N_18638,N_18647);
nor U18994 (N_18994,N_18676,N_18745);
nor U18995 (N_18995,N_18683,N_18739);
and U18996 (N_18996,N_18767,N_18612);
nand U18997 (N_18997,N_18782,N_18753);
nor U18998 (N_18998,N_18785,N_18782);
nor U18999 (N_18999,N_18663,N_18674);
nor U19000 (N_19000,N_18860,N_18838);
nor U19001 (N_19001,N_18847,N_18803);
nand U19002 (N_19002,N_18962,N_18912);
and U19003 (N_19003,N_18923,N_18997);
or U19004 (N_19004,N_18963,N_18864);
nand U19005 (N_19005,N_18842,N_18824);
nor U19006 (N_19006,N_18922,N_18807);
and U19007 (N_19007,N_18843,N_18900);
and U19008 (N_19008,N_18934,N_18894);
nor U19009 (N_19009,N_18820,N_18953);
or U19010 (N_19010,N_18806,N_18938);
and U19011 (N_19011,N_18883,N_18932);
and U19012 (N_19012,N_18835,N_18837);
nor U19013 (N_19013,N_18839,N_18970);
or U19014 (N_19014,N_18878,N_18898);
and U19015 (N_19015,N_18821,N_18901);
or U19016 (N_19016,N_18939,N_18859);
or U19017 (N_19017,N_18930,N_18831);
nand U19018 (N_19018,N_18915,N_18907);
and U19019 (N_19019,N_18999,N_18988);
nand U19020 (N_19020,N_18814,N_18980);
and U19021 (N_19021,N_18986,N_18949);
nand U19022 (N_19022,N_18950,N_18882);
nor U19023 (N_19023,N_18952,N_18909);
nor U19024 (N_19024,N_18879,N_18959);
or U19025 (N_19025,N_18816,N_18853);
nand U19026 (N_19026,N_18913,N_18892);
and U19027 (N_19027,N_18976,N_18931);
and U19028 (N_19028,N_18940,N_18925);
or U19029 (N_19029,N_18858,N_18867);
xor U19030 (N_19030,N_18848,N_18929);
or U19031 (N_19031,N_18895,N_18979);
nand U19032 (N_19032,N_18924,N_18902);
nor U19033 (N_19033,N_18891,N_18822);
nand U19034 (N_19034,N_18927,N_18872);
nand U19035 (N_19035,N_18948,N_18893);
or U19036 (N_19036,N_18996,N_18828);
or U19037 (N_19037,N_18857,N_18871);
nand U19038 (N_19038,N_18802,N_18886);
nand U19039 (N_19039,N_18942,N_18861);
and U19040 (N_19040,N_18875,N_18995);
or U19041 (N_19041,N_18955,N_18967);
nor U19042 (N_19042,N_18851,N_18916);
nand U19043 (N_19043,N_18812,N_18983);
nand U19044 (N_19044,N_18978,N_18868);
or U19045 (N_19045,N_18844,N_18887);
and U19046 (N_19046,N_18852,N_18947);
and U19047 (N_19047,N_18877,N_18840);
or U19048 (N_19048,N_18805,N_18823);
or U19049 (N_19049,N_18965,N_18817);
nor U19050 (N_19050,N_18982,N_18889);
nor U19051 (N_19051,N_18935,N_18825);
and U19052 (N_19052,N_18808,N_18973);
and U19053 (N_19053,N_18917,N_18841);
nor U19054 (N_19054,N_18914,N_18881);
and U19055 (N_19055,N_18869,N_18946);
nor U19056 (N_19056,N_18870,N_18921);
nor U19057 (N_19057,N_18818,N_18829);
or U19058 (N_19058,N_18928,N_18903);
or U19059 (N_19059,N_18890,N_18998);
nand U19060 (N_19060,N_18984,N_18800);
and U19061 (N_19061,N_18993,N_18957);
nand U19062 (N_19062,N_18854,N_18933);
or U19063 (N_19063,N_18911,N_18856);
nand U19064 (N_19064,N_18888,N_18813);
nor U19065 (N_19065,N_18846,N_18863);
or U19066 (N_19066,N_18885,N_18977);
nor U19067 (N_19067,N_18966,N_18919);
nand U19068 (N_19068,N_18876,N_18918);
nand U19069 (N_19069,N_18954,N_18849);
and U19070 (N_19070,N_18811,N_18956);
nand U19071 (N_19071,N_18809,N_18972);
nand U19072 (N_19072,N_18968,N_18832);
or U19073 (N_19073,N_18906,N_18985);
and U19074 (N_19074,N_18810,N_18941);
nor U19075 (N_19075,N_18884,N_18936);
nor U19076 (N_19076,N_18964,N_18834);
and U19077 (N_19077,N_18880,N_18944);
nand U19078 (N_19078,N_18873,N_18874);
or U19079 (N_19079,N_18926,N_18975);
or U19080 (N_19080,N_18981,N_18937);
or U19081 (N_19081,N_18855,N_18899);
or U19082 (N_19082,N_18910,N_18920);
nor U19083 (N_19083,N_18908,N_18905);
and U19084 (N_19084,N_18897,N_18866);
or U19085 (N_19085,N_18945,N_18974);
or U19086 (N_19086,N_18990,N_18951);
nor U19087 (N_19087,N_18801,N_18826);
and U19088 (N_19088,N_18971,N_18865);
or U19089 (N_19089,N_18850,N_18969);
and U19090 (N_19090,N_18819,N_18989);
nand U19091 (N_19091,N_18827,N_18833);
or U19092 (N_19092,N_18958,N_18943);
and U19093 (N_19093,N_18896,N_18987);
and U19094 (N_19094,N_18994,N_18904);
and U19095 (N_19095,N_18845,N_18830);
and U19096 (N_19096,N_18992,N_18804);
or U19097 (N_19097,N_18815,N_18991);
nor U19098 (N_19098,N_18836,N_18961);
nor U19099 (N_19099,N_18960,N_18862);
nor U19100 (N_19100,N_18996,N_18986);
and U19101 (N_19101,N_18873,N_18965);
or U19102 (N_19102,N_18854,N_18923);
and U19103 (N_19103,N_18820,N_18949);
and U19104 (N_19104,N_18894,N_18834);
nand U19105 (N_19105,N_18938,N_18856);
and U19106 (N_19106,N_18962,N_18968);
nor U19107 (N_19107,N_18806,N_18874);
and U19108 (N_19108,N_18897,N_18970);
and U19109 (N_19109,N_18803,N_18859);
or U19110 (N_19110,N_18947,N_18892);
nand U19111 (N_19111,N_18952,N_18997);
nor U19112 (N_19112,N_18934,N_18877);
xor U19113 (N_19113,N_18837,N_18946);
and U19114 (N_19114,N_18810,N_18910);
nand U19115 (N_19115,N_18988,N_18877);
nand U19116 (N_19116,N_18820,N_18973);
nand U19117 (N_19117,N_18924,N_18975);
and U19118 (N_19118,N_18833,N_18863);
nand U19119 (N_19119,N_18939,N_18917);
and U19120 (N_19120,N_18866,N_18994);
or U19121 (N_19121,N_18970,N_18999);
nor U19122 (N_19122,N_18846,N_18942);
nand U19123 (N_19123,N_18988,N_18836);
and U19124 (N_19124,N_18944,N_18890);
or U19125 (N_19125,N_18913,N_18824);
nand U19126 (N_19126,N_18861,N_18846);
and U19127 (N_19127,N_18934,N_18876);
nor U19128 (N_19128,N_18950,N_18840);
nand U19129 (N_19129,N_18868,N_18826);
and U19130 (N_19130,N_18894,N_18818);
and U19131 (N_19131,N_18894,N_18805);
nand U19132 (N_19132,N_18927,N_18934);
nor U19133 (N_19133,N_18944,N_18843);
or U19134 (N_19134,N_18852,N_18989);
nor U19135 (N_19135,N_18890,N_18967);
and U19136 (N_19136,N_18867,N_18919);
nand U19137 (N_19137,N_18994,N_18911);
nand U19138 (N_19138,N_18880,N_18856);
and U19139 (N_19139,N_18972,N_18885);
and U19140 (N_19140,N_18827,N_18898);
or U19141 (N_19141,N_18975,N_18880);
and U19142 (N_19142,N_18979,N_18998);
nor U19143 (N_19143,N_18878,N_18861);
nand U19144 (N_19144,N_18881,N_18877);
and U19145 (N_19145,N_18904,N_18927);
and U19146 (N_19146,N_18821,N_18902);
nand U19147 (N_19147,N_18969,N_18813);
nand U19148 (N_19148,N_18904,N_18931);
nor U19149 (N_19149,N_18905,N_18933);
nor U19150 (N_19150,N_18871,N_18840);
and U19151 (N_19151,N_18933,N_18956);
and U19152 (N_19152,N_18992,N_18815);
nor U19153 (N_19153,N_18855,N_18830);
and U19154 (N_19154,N_18847,N_18958);
nor U19155 (N_19155,N_18936,N_18808);
nand U19156 (N_19156,N_18990,N_18987);
or U19157 (N_19157,N_18936,N_18944);
and U19158 (N_19158,N_18855,N_18972);
nor U19159 (N_19159,N_18816,N_18965);
and U19160 (N_19160,N_18976,N_18899);
or U19161 (N_19161,N_18904,N_18894);
nor U19162 (N_19162,N_18843,N_18989);
nand U19163 (N_19163,N_18818,N_18858);
or U19164 (N_19164,N_18923,N_18934);
nor U19165 (N_19165,N_18877,N_18953);
or U19166 (N_19166,N_18998,N_18842);
nor U19167 (N_19167,N_18944,N_18851);
or U19168 (N_19168,N_18836,N_18816);
nor U19169 (N_19169,N_18940,N_18802);
nand U19170 (N_19170,N_18929,N_18898);
xnor U19171 (N_19171,N_18973,N_18889);
or U19172 (N_19172,N_18905,N_18831);
nor U19173 (N_19173,N_18968,N_18883);
nor U19174 (N_19174,N_18832,N_18985);
and U19175 (N_19175,N_18812,N_18968);
and U19176 (N_19176,N_18885,N_18816);
nand U19177 (N_19177,N_18891,N_18819);
nor U19178 (N_19178,N_18816,N_18849);
and U19179 (N_19179,N_18841,N_18832);
nand U19180 (N_19180,N_18886,N_18881);
or U19181 (N_19181,N_18927,N_18932);
xor U19182 (N_19182,N_18972,N_18913);
nor U19183 (N_19183,N_18818,N_18820);
and U19184 (N_19184,N_18864,N_18845);
nand U19185 (N_19185,N_18821,N_18812);
xnor U19186 (N_19186,N_18992,N_18933);
nand U19187 (N_19187,N_18876,N_18959);
nand U19188 (N_19188,N_18890,N_18901);
and U19189 (N_19189,N_18829,N_18950);
nand U19190 (N_19190,N_18837,N_18803);
nand U19191 (N_19191,N_18894,N_18893);
nand U19192 (N_19192,N_18886,N_18867);
nand U19193 (N_19193,N_18992,N_18900);
nand U19194 (N_19194,N_18819,N_18888);
nor U19195 (N_19195,N_18904,N_18861);
or U19196 (N_19196,N_18936,N_18912);
nand U19197 (N_19197,N_18802,N_18861);
nand U19198 (N_19198,N_18954,N_18969);
nor U19199 (N_19199,N_18901,N_18938);
and U19200 (N_19200,N_19145,N_19170);
nor U19201 (N_19201,N_19131,N_19122);
nand U19202 (N_19202,N_19016,N_19015);
or U19203 (N_19203,N_19076,N_19161);
nor U19204 (N_19204,N_19133,N_19088);
nor U19205 (N_19205,N_19130,N_19199);
nor U19206 (N_19206,N_19094,N_19022);
nand U19207 (N_19207,N_19101,N_19193);
nand U19208 (N_19208,N_19182,N_19143);
nor U19209 (N_19209,N_19045,N_19175);
nor U19210 (N_19210,N_19119,N_19001);
or U19211 (N_19211,N_19085,N_19194);
nand U19212 (N_19212,N_19025,N_19113);
or U19213 (N_19213,N_19116,N_19059);
or U19214 (N_19214,N_19018,N_19047);
or U19215 (N_19215,N_19051,N_19083);
nand U19216 (N_19216,N_19033,N_19035);
or U19217 (N_19217,N_19055,N_19006);
and U19218 (N_19218,N_19102,N_19177);
nand U19219 (N_19219,N_19013,N_19089);
or U19220 (N_19220,N_19106,N_19180);
and U19221 (N_19221,N_19136,N_19184);
and U19222 (N_19222,N_19112,N_19171);
and U19223 (N_19223,N_19117,N_19123);
nor U19224 (N_19224,N_19169,N_19030);
nand U19225 (N_19225,N_19172,N_19084);
nor U19226 (N_19226,N_19107,N_19026);
and U19227 (N_19227,N_19140,N_19056);
nor U19228 (N_19228,N_19192,N_19178);
nand U19229 (N_19229,N_19086,N_19103);
nand U19230 (N_19230,N_19114,N_19005);
and U19231 (N_19231,N_19142,N_19160);
nand U19232 (N_19232,N_19121,N_19141);
or U19233 (N_19233,N_19064,N_19146);
nor U19234 (N_19234,N_19167,N_19037);
nor U19235 (N_19235,N_19154,N_19111);
nand U19236 (N_19236,N_19007,N_19072);
and U19237 (N_19237,N_19100,N_19189);
and U19238 (N_19238,N_19050,N_19173);
or U19239 (N_19239,N_19129,N_19069);
nor U19240 (N_19240,N_19183,N_19097);
nand U19241 (N_19241,N_19004,N_19048);
or U19242 (N_19242,N_19075,N_19179);
and U19243 (N_19243,N_19165,N_19021);
or U19244 (N_19244,N_19078,N_19127);
nand U19245 (N_19245,N_19115,N_19009);
nand U19246 (N_19246,N_19042,N_19063);
nor U19247 (N_19247,N_19020,N_19155);
or U19248 (N_19248,N_19062,N_19126);
or U19249 (N_19249,N_19185,N_19068);
nand U19250 (N_19250,N_19176,N_19124);
nand U19251 (N_19251,N_19036,N_19073);
nand U19252 (N_19252,N_19144,N_19087);
or U19253 (N_19253,N_19156,N_19028);
nand U19254 (N_19254,N_19061,N_19091);
or U19255 (N_19255,N_19197,N_19044);
or U19256 (N_19256,N_19152,N_19137);
and U19257 (N_19257,N_19120,N_19057);
nand U19258 (N_19258,N_19108,N_19039);
nor U19259 (N_19259,N_19032,N_19034);
or U19260 (N_19260,N_19198,N_19077);
nor U19261 (N_19261,N_19168,N_19052);
nor U19262 (N_19262,N_19149,N_19027);
and U19263 (N_19263,N_19181,N_19002);
and U19264 (N_19264,N_19000,N_19067);
and U19265 (N_19265,N_19053,N_19138);
and U19266 (N_19266,N_19139,N_19024);
or U19267 (N_19267,N_19003,N_19110);
nand U19268 (N_19268,N_19095,N_19065);
nor U19269 (N_19269,N_19099,N_19186);
nand U19270 (N_19270,N_19014,N_19038);
nand U19271 (N_19271,N_19066,N_19040);
or U19272 (N_19272,N_19096,N_19188);
xor U19273 (N_19273,N_19118,N_19031);
nand U19274 (N_19274,N_19151,N_19054);
nand U19275 (N_19275,N_19148,N_19159);
and U19276 (N_19276,N_19109,N_19191);
nor U19277 (N_19277,N_19125,N_19019);
nand U19278 (N_19278,N_19104,N_19081);
or U19279 (N_19279,N_19058,N_19079);
and U19280 (N_19280,N_19012,N_19150);
nor U19281 (N_19281,N_19132,N_19092);
xor U19282 (N_19282,N_19105,N_19158);
nand U19283 (N_19283,N_19060,N_19147);
xor U19284 (N_19284,N_19196,N_19011);
nand U19285 (N_19285,N_19017,N_19164);
or U19286 (N_19286,N_19134,N_19082);
and U19287 (N_19287,N_19041,N_19174);
nand U19288 (N_19288,N_19190,N_19029);
nor U19289 (N_19289,N_19153,N_19163);
nor U19290 (N_19290,N_19135,N_19090);
xor U19291 (N_19291,N_19093,N_19043);
and U19292 (N_19292,N_19074,N_19010);
or U19293 (N_19293,N_19128,N_19098);
or U19294 (N_19294,N_19008,N_19049);
and U19295 (N_19295,N_19162,N_19080);
or U19296 (N_19296,N_19046,N_19195);
xnor U19297 (N_19297,N_19071,N_19023);
and U19298 (N_19298,N_19187,N_19070);
nor U19299 (N_19299,N_19157,N_19166);
nor U19300 (N_19300,N_19055,N_19136);
nor U19301 (N_19301,N_19039,N_19035);
or U19302 (N_19302,N_19141,N_19043);
or U19303 (N_19303,N_19131,N_19022);
nand U19304 (N_19304,N_19162,N_19081);
and U19305 (N_19305,N_19065,N_19018);
or U19306 (N_19306,N_19083,N_19066);
and U19307 (N_19307,N_19056,N_19052);
and U19308 (N_19308,N_19115,N_19199);
nand U19309 (N_19309,N_19179,N_19062);
and U19310 (N_19310,N_19042,N_19122);
or U19311 (N_19311,N_19029,N_19158);
nor U19312 (N_19312,N_19022,N_19104);
nand U19313 (N_19313,N_19019,N_19096);
and U19314 (N_19314,N_19105,N_19195);
nor U19315 (N_19315,N_19019,N_19016);
or U19316 (N_19316,N_19045,N_19055);
or U19317 (N_19317,N_19161,N_19105);
nor U19318 (N_19318,N_19046,N_19093);
and U19319 (N_19319,N_19155,N_19029);
and U19320 (N_19320,N_19069,N_19095);
nand U19321 (N_19321,N_19019,N_19115);
and U19322 (N_19322,N_19161,N_19007);
and U19323 (N_19323,N_19175,N_19078);
nand U19324 (N_19324,N_19095,N_19084);
nor U19325 (N_19325,N_19166,N_19062);
nor U19326 (N_19326,N_19065,N_19108);
and U19327 (N_19327,N_19051,N_19056);
nand U19328 (N_19328,N_19017,N_19068);
or U19329 (N_19329,N_19038,N_19198);
or U19330 (N_19330,N_19117,N_19113);
nor U19331 (N_19331,N_19084,N_19173);
and U19332 (N_19332,N_19129,N_19177);
nor U19333 (N_19333,N_19073,N_19168);
nor U19334 (N_19334,N_19119,N_19076);
or U19335 (N_19335,N_19006,N_19117);
nand U19336 (N_19336,N_19050,N_19081);
and U19337 (N_19337,N_19123,N_19157);
or U19338 (N_19338,N_19039,N_19045);
or U19339 (N_19339,N_19091,N_19132);
nand U19340 (N_19340,N_19041,N_19017);
nand U19341 (N_19341,N_19110,N_19163);
nor U19342 (N_19342,N_19127,N_19183);
or U19343 (N_19343,N_19192,N_19142);
nand U19344 (N_19344,N_19123,N_19106);
nand U19345 (N_19345,N_19001,N_19161);
and U19346 (N_19346,N_19107,N_19173);
and U19347 (N_19347,N_19159,N_19130);
nand U19348 (N_19348,N_19124,N_19083);
and U19349 (N_19349,N_19067,N_19009);
or U19350 (N_19350,N_19186,N_19009);
and U19351 (N_19351,N_19198,N_19024);
or U19352 (N_19352,N_19079,N_19115);
and U19353 (N_19353,N_19000,N_19137);
or U19354 (N_19354,N_19087,N_19118);
or U19355 (N_19355,N_19051,N_19129);
and U19356 (N_19356,N_19046,N_19033);
and U19357 (N_19357,N_19133,N_19074);
and U19358 (N_19358,N_19093,N_19085);
or U19359 (N_19359,N_19076,N_19094);
nor U19360 (N_19360,N_19057,N_19190);
nand U19361 (N_19361,N_19099,N_19060);
and U19362 (N_19362,N_19113,N_19067);
or U19363 (N_19363,N_19120,N_19079);
or U19364 (N_19364,N_19173,N_19092);
nand U19365 (N_19365,N_19006,N_19100);
or U19366 (N_19366,N_19030,N_19185);
and U19367 (N_19367,N_19061,N_19175);
or U19368 (N_19368,N_19015,N_19088);
nand U19369 (N_19369,N_19076,N_19096);
nand U19370 (N_19370,N_19102,N_19165);
nand U19371 (N_19371,N_19174,N_19086);
nand U19372 (N_19372,N_19097,N_19017);
and U19373 (N_19373,N_19192,N_19193);
nand U19374 (N_19374,N_19121,N_19021);
or U19375 (N_19375,N_19015,N_19046);
nand U19376 (N_19376,N_19020,N_19196);
and U19377 (N_19377,N_19099,N_19156);
nor U19378 (N_19378,N_19004,N_19179);
nor U19379 (N_19379,N_19182,N_19108);
nand U19380 (N_19380,N_19064,N_19135);
nand U19381 (N_19381,N_19193,N_19020);
nand U19382 (N_19382,N_19012,N_19102);
nor U19383 (N_19383,N_19192,N_19032);
nor U19384 (N_19384,N_19162,N_19026);
or U19385 (N_19385,N_19097,N_19181);
nand U19386 (N_19386,N_19033,N_19106);
or U19387 (N_19387,N_19151,N_19183);
or U19388 (N_19388,N_19155,N_19002);
or U19389 (N_19389,N_19031,N_19121);
and U19390 (N_19390,N_19096,N_19178);
and U19391 (N_19391,N_19153,N_19180);
nand U19392 (N_19392,N_19079,N_19105);
nand U19393 (N_19393,N_19057,N_19177);
nor U19394 (N_19394,N_19173,N_19067);
nor U19395 (N_19395,N_19048,N_19031);
nor U19396 (N_19396,N_19185,N_19071);
nand U19397 (N_19397,N_19179,N_19012);
and U19398 (N_19398,N_19051,N_19019);
or U19399 (N_19399,N_19118,N_19139);
nand U19400 (N_19400,N_19241,N_19271);
nor U19401 (N_19401,N_19243,N_19329);
nand U19402 (N_19402,N_19349,N_19317);
or U19403 (N_19403,N_19345,N_19307);
and U19404 (N_19404,N_19259,N_19244);
or U19405 (N_19405,N_19256,N_19223);
nor U19406 (N_19406,N_19293,N_19253);
nor U19407 (N_19407,N_19354,N_19363);
nor U19408 (N_19408,N_19252,N_19397);
or U19409 (N_19409,N_19234,N_19261);
nor U19410 (N_19410,N_19388,N_19267);
or U19411 (N_19411,N_19394,N_19284);
nor U19412 (N_19412,N_19327,N_19297);
nand U19413 (N_19413,N_19260,N_19213);
nor U19414 (N_19414,N_19298,N_19233);
and U19415 (N_19415,N_19254,N_19276);
nor U19416 (N_19416,N_19396,N_19302);
nor U19417 (N_19417,N_19375,N_19226);
nand U19418 (N_19418,N_19371,N_19391);
nor U19419 (N_19419,N_19376,N_19247);
nor U19420 (N_19420,N_19257,N_19323);
nor U19421 (N_19421,N_19255,N_19258);
or U19422 (N_19422,N_19335,N_19389);
nor U19423 (N_19423,N_19320,N_19315);
and U19424 (N_19424,N_19299,N_19357);
and U19425 (N_19425,N_19339,N_19246);
or U19426 (N_19426,N_19344,N_19285);
nor U19427 (N_19427,N_19273,N_19319);
and U19428 (N_19428,N_19203,N_19304);
and U19429 (N_19429,N_19381,N_19263);
or U19430 (N_19430,N_19309,N_19240);
nor U19431 (N_19431,N_19303,N_19379);
or U19432 (N_19432,N_19300,N_19272);
nor U19433 (N_19433,N_19236,N_19383);
nor U19434 (N_19434,N_19294,N_19331);
or U19435 (N_19435,N_19370,N_19237);
and U19436 (N_19436,N_19217,N_19204);
or U19437 (N_19437,N_19269,N_19205);
nor U19438 (N_19438,N_19248,N_19295);
nor U19439 (N_19439,N_19367,N_19313);
and U19440 (N_19440,N_19326,N_19333);
nor U19441 (N_19441,N_19242,N_19201);
nor U19442 (N_19442,N_19321,N_19372);
or U19443 (N_19443,N_19336,N_19245);
nor U19444 (N_19444,N_19206,N_19220);
nor U19445 (N_19445,N_19274,N_19310);
nor U19446 (N_19446,N_19291,N_19387);
or U19447 (N_19447,N_19270,N_19341);
nor U19448 (N_19448,N_19377,N_19399);
nor U19449 (N_19449,N_19359,N_19338);
nor U19450 (N_19450,N_19228,N_19250);
or U19451 (N_19451,N_19325,N_19222);
nand U19452 (N_19452,N_19292,N_19282);
or U19453 (N_19453,N_19356,N_19347);
and U19454 (N_19454,N_19361,N_19268);
nor U19455 (N_19455,N_19279,N_19211);
nor U19456 (N_19456,N_19229,N_19390);
nor U19457 (N_19457,N_19306,N_19221);
or U19458 (N_19458,N_19322,N_19382);
nor U19459 (N_19459,N_19227,N_19350);
or U19460 (N_19460,N_19262,N_19219);
nand U19461 (N_19461,N_19353,N_19374);
nand U19462 (N_19462,N_19348,N_19230);
nand U19463 (N_19463,N_19360,N_19373);
and U19464 (N_19464,N_19231,N_19385);
nor U19465 (N_19465,N_19316,N_19378);
or U19466 (N_19466,N_19318,N_19398);
and U19467 (N_19467,N_19288,N_19311);
nor U19468 (N_19468,N_19395,N_19314);
xnor U19469 (N_19469,N_19209,N_19355);
and U19470 (N_19470,N_19384,N_19278);
nor U19471 (N_19471,N_19366,N_19343);
or U19472 (N_19472,N_19296,N_19312);
nand U19473 (N_19473,N_19200,N_19281);
nand U19474 (N_19474,N_19251,N_19214);
nor U19475 (N_19475,N_19308,N_19328);
or U19476 (N_19476,N_19207,N_19238);
nor U19477 (N_19477,N_19264,N_19224);
or U19478 (N_19478,N_19351,N_19301);
or U19479 (N_19479,N_19340,N_19235);
and U19480 (N_19480,N_19208,N_19287);
nor U19481 (N_19481,N_19332,N_19386);
nor U19482 (N_19482,N_19289,N_19265);
nor U19483 (N_19483,N_19218,N_19368);
nor U19484 (N_19484,N_19330,N_19283);
nand U19485 (N_19485,N_19324,N_19393);
or U19486 (N_19486,N_19249,N_19342);
nor U19487 (N_19487,N_19275,N_19365);
nor U19488 (N_19488,N_19337,N_19352);
nor U19489 (N_19489,N_19280,N_19210);
or U19490 (N_19490,N_19369,N_19380);
nand U19491 (N_19491,N_19266,N_19216);
nand U19492 (N_19492,N_19202,N_19232);
nand U19493 (N_19493,N_19225,N_19239);
nor U19494 (N_19494,N_19212,N_19362);
and U19495 (N_19495,N_19277,N_19358);
nor U19496 (N_19496,N_19346,N_19286);
nor U19497 (N_19497,N_19215,N_19392);
or U19498 (N_19498,N_19364,N_19290);
and U19499 (N_19499,N_19334,N_19305);
nand U19500 (N_19500,N_19389,N_19291);
nor U19501 (N_19501,N_19350,N_19229);
nand U19502 (N_19502,N_19231,N_19359);
or U19503 (N_19503,N_19288,N_19259);
nand U19504 (N_19504,N_19397,N_19304);
or U19505 (N_19505,N_19211,N_19246);
or U19506 (N_19506,N_19383,N_19388);
nor U19507 (N_19507,N_19246,N_19256);
and U19508 (N_19508,N_19324,N_19388);
nand U19509 (N_19509,N_19382,N_19243);
and U19510 (N_19510,N_19284,N_19300);
nor U19511 (N_19511,N_19212,N_19232);
and U19512 (N_19512,N_19240,N_19210);
or U19513 (N_19513,N_19329,N_19355);
and U19514 (N_19514,N_19328,N_19237);
or U19515 (N_19515,N_19259,N_19219);
nand U19516 (N_19516,N_19391,N_19399);
nand U19517 (N_19517,N_19263,N_19311);
or U19518 (N_19518,N_19364,N_19232);
and U19519 (N_19519,N_19394,N_19313);
and U19520 (N_19520,N_19378,N_19365);
nor U19521 (N_19521,N_19363,N_19291);
nor U19522 (N_19522,N_19291,N_19344);
nor U19523 (N_19523,N_19298,N_19281);
and U19524 (N_19524,N_19396,N_19383);
and U19525 (N_19525,N_19303,N_19330);
nor U19526 (N_19526,N_19240,N_19347);
nor U19527 (N_19527,N_19372,N_19227);
or U19528 (N_19528,N_19385,N_19255);
and U19529 (N_19529,N_19249,N_19354);
or U19530 (N_19530,N_19391,N_19237);
nor U19531 (N_19531,N_19267,N_19254);
or U19532 (N_19532,N_19291,N_19218);
nand U19533 (N_19533,N_19308,N_19221);
nand U19534 (N_19534,N_19233,N_19302);
and U19535 (N_19535,N_19309,N_19230);
or U19536 (N_19536,N_19334,N_19261);
nor U19537 (N_19537,N_19348,N_19387);
or U19538 (N_19538,N_19274,N_19350);
and U19539 (N_19539,N_19345,N_19269);
nand U19540 (N_19540,N_19246,N_19218);
nand U19541 (N_19541,N_19231,N_19236);
or U19542 (N_19542,N_19246,N_19297);
and U19543 (N_19543,N_19355,N_19214);
or U19544 (N_19544,N_19226,N_19389);
nor U19545 (N_19545,N_19297,N_19360);
and U19546 (N_19546,N_19289,N_19308);
nand U19547 (N_19547,N_19382,N_19225);
or U19548 (N_19548,N_19234,N_19210);
and U19549 (N_19549,N_19384,N_19389);
nand U19550 (N_19550,N_19298,N_19216);
and U19551 (N_19551,N_19243,N_19336);
and U19552 (N_19552,N_19221,N_19251);
nor U19553 (N_19553,N_19331,N_19368);
or U19554 (N_19554,N_19309,N_19269);
or U19555 (N_19555,N_19311,N_19286);
and U19556 (N_19556,N_19296,N_19220);
nand U19557 (N_19557,N_19258,N_19236);
nor U19558 (N_19558,N_19240,N_19255);
nand U19559 (N_19559,N_19376,N_19289);
and U19560 (N_19560,N_19385,N_19306);
nand U19561 (N_19561,N_19231,N_19232);
nor U19562 (N_19562,N_19296,N_19321);
or U19563 (N_19563,N_19341,N_19351);
nand U19564 (N_19564,N_19295,N_19385);
nor U19565 (N_19565,N_19273,N_19330);
nand U19566 (N_19566,N_19271,N_19342);
nand U19567 (N_19567,N_19300,N_19276);
and U19568 (N_19568,N_19353,N_19260);
nand U19569 (N_19569,N_19286,N_19325);
xnor U19570 (N_19570,N_19357,N_19378);
and U19571 (N_19571,N_19303,N_19336);
nand U19572 (N_19572,N_19353,N_19270);
nand U19573 (N_19573,N_19227,N_19311);
nor U19574 (N_19574,N_19260,N_19357);
or U19575 (N_19575,N_19258,N_19342);
nor U19576 (N_19576,N_19228,N_19276);
and U19577 (N_19577,N_19305,N_19315);
or U19578 (N_19578,N_19334,N_19230);
nor U19579 (N_19579,N_19283,N_19219);
and U19580 (N_19580,N_19223,N_19233);
xor U19581 (N_19581,N_19305,N_19359);
nor U19582 (N_19582,N_19246,N_19326);
and U19583 (N_19583,N_19397,N_19390);
and U19584 (N_19584,N_19365,N_19235);
nand U19585 (N_19585,N_19259,N_19325);
nand U19586 (N_19586,N_19268,N_19320);
and U19587 (N_19587,N_19233,N_19202);
or U19588 (N_19588,N_19382,N_19252);
or U19589 (N_19589,N_19335,N_19221);
nand U19590 (N_19590,N_19274,N_19369);
and U19591 (N_19591,N_19204,N_19364);
and U19592 (N_19592,N_19229,N_19221);
nor U19593 (N_19593,N_19379,N_19305);
nand U19594 (N_19594,N_19350,N_19311);
nand U19595 (N_19595,N_19351,N_19230);
or U19596 (N_19596,N_19328,N_19391);
and U19597 (N_19597,N_19241,N_19397);
and U19598 (N_19598,N_19291,N_19293);
and U19599 (N_19599,N_19255,N_19201);
nand U19600 (N_19600,N_19565,N_19454);
or U19601 (N_19601,N_19418,N_19438);
and U19602 (N_19602,N_19548,N_19465);
or U19603 (N_19603,N_19592,N_19506);
and U19604 (N_19604,N_19415,N_19480);
or U19605 (N_19605,N_19582,N_19424);
and U19606 (N_19606,N_19487,N_19597);
nand U19607 (N_19607,N_19514,N_19492);
xor U19608 (N_19608,N_19484,N_19446);
nor U19609 (N_19609,N_19490,N_19491);
nor U19610 (N_19610,N_19502,N_19545);
and U19611 (N_19611,N_19432,N_19584);
and U19612 (N_19612,N_19586,N_19554);
nand U19613 (N_19613,N_19587,N_19580);
nand U19614 (N_19614,N_19429,N_19590);
nor U19615 (N_19615,N_19523,N_19441);
or U19616 (N_19616,N_19516,N_19403);
nand U19617 (N_19617,N_19569,N_19439);
or U19618 (N_19618,N_19483,N_19504);
nor U19619 (N_19619,N_19411,N_19528);
nand U19620 (N_19620,N_19486,N_19508);
or U19621 (N_19621,N_19416,N_19517);
nor U19622 (N_19622,N_19570,N_19522);
or U19623 (N_19623,N_19420,N_19477);
xor U19624 (N_19624,N_19470,N_19524);
nor U19625 (N_19625,N_19437,N_19573);
nor U19626 (N_19626,N_19534,N_19594);
or U19627 (N_19627,N_19460,N_19469);
nand U19628 (N_19628,N_19510,N_19550);
or U19629 (N_19629,N_19450,N_19464);
nor U19630 (N_19630,N_19479,N_19551);
nand U19631 (N_19631,N_19585,N_19478);
nor U19632 (N_19632,N_19596,N_19501);
nand U19633 (N_19633,N_19560,N_19567);
nor U19634 (N_19634,N_19414,N_19507);
nor U19635 (N_19635,N_19494,N_19476);
or U19636 (N_19636,N_19520,N_19406);
and U19637 (N_19637,N_19595,N_19557);
or U19638 (N_19638,N_19509,N_19530);
nand U19639 (N_19639,N_19515,N_19559);
and U19640 (N_19640,N_19453,N_19422);
nand U19641 (N_19641,N_19579,N_19417);
or U19642 (N_19642,N_19404,N_19410);
nor U19643 (N_19643,N_19500,N_19461);
or U19644 (N_19644,N_19433,N_19436);
nand U19645 (N_19645,N_19529,N_19525);
nand U19646 (N_19646,N_19430,N_19442);
nand U19647 (N_19647,N_19571,N_19544);
xnor U19648 (N_19648,N_19543,N_19549);
nor U19649 (N_19649,N_19527,N_19493);
nor U19650 (N_19650,N_19540,N_19497);
nand U19651 (N_19651,N_19466,N_19568);
and U19652 (N_19652,N_19405,N_19558);
nand U19653 (N_19653,N_19519,N_19496);
nor U19654 (N_19654,N_19577,N_19566);
and U19655 (N_19655,N_19532,N_19481);
or U19656 (N_19656,N_19408,N_19456);
or U19657 (N_19657,N_19407,N_19458);
xor U19658 (N_19658,N_19434,N_19448);
nor U19659 (N_19659,N_19537,N_19400);
nor U19660 (N_19660,N_19463,N_19447);
nor U19661 (N_19661,N_19511,N_19402);
and U19662 (N_19662,N_19563,N_19435);
nor U19663 (N_19663,N_19427,N_19588);
nor U19664 (N_19664,N_19547,N_19574);
and U19665 (N_19665,N_19518,N_19452);
nand U19666 (N_19666,N_19553,N_19451);
or U19667 (N_19667,N_19489,N_19462);
nand U19668 (N_19668,N_19555,N_19485);
nor U19669 (N_19669,N_19538,N_19419);
and U19670 (N_19670,N_19526,N_19505);
or U19671 (N_19671,N_19425,N_19457);
and U19672 (N_19672,N_19512,N_19473);
nand U19673 (N_19673,N_19591,N_19546);
nor U19674 (N_19674,N_19426,N_19536);
nor U19675 (N_19675,N_19589,N_19583);
and U19676 (N_19676,N_19572,N_19541);
nor U19677 (N_19677,N_19535,N_19421);
nor U19678 (N_19678,N_19413,N_19495);
or U19679 (N_19679,N_19423,N_19471);
nor U19680 (N_19680,N_19521,N_19468);
or U19681 (N_19681,N_19459,N_19564);
or U19682 (N_19682,N_19533,N_19576);
nor U19683 (N_19683,N_19575,N_19482);
nor U19684 (N_19684,N_19542,N_19499);
or U19685 (N_19685,N_19578,N_19475);
nor U19686 (N_19686,N_19472,N_19561);
or U19687 (N_19687,N_19401,N_19412);
nand U19688 (N_19688,N_19498,N_19467);
nor U19689 (N_19689,N_19593,N_19503);
and U19690 (N_19690,N_19581,N_19539);
or U19691 (N_19691,N_19552,N_19474);
and U19692 (N_19692,N_19440,N_19443);
or U19693 (N_19693,N_19556,N_19455);
nor U19694 (N_19694,N_19431,N_19444);
nor U19695 (N_19695,N_19445,N_19598);
nor U19696 (N_19696,N_19513,N_19599);
or U19697 (N_19697,N_19449,N_19562);
nor U19698 (N_19698,N_19531,N_19409);
or U19699 (N_19699,N_19488,N_19428);
and U19700 (N_19700,N_19528,N_19443);
and U19701 (N_19701,N_19443,N_19587);
nand U19702 (N_19702,N_19440,N_19521);
and U19703 (N_19703,N_19461,N_19453);
nor U19704 (N_19704,N_19523,N_19570);
nor U19705 (N_19705,N_19489,N_19459);
nand U19706 (N_19706,N_19574,N_19568);
and U19707 (N_19707,N_19411,N_19504);
nor U19708 (N_19708,N_19515,N_19420);
nand U19709 (N_19709,N_19496,N_19489);
nand U19710 (N_19710,N_19544,N_19589);
nand U19711 (N_19711,N_19430,N_19467);
nand U19712 (N_19712,N_19479,N_19584);
or U19713 (N_19713,N_19450,N_19572);
nor U19714 (N_19714,N_19452,N_19446);
or U19715 (N_19715,N_19511,N_19417);
and U19716 (N_19716,N_19432,N_19442);
xor U19717 (N_19717,N_19481,N_19527);
or U19718 (N_19718,N_19579,N_19488);
and U19719 (N_19719,N_19434,N_19464);
or U19720 (N_19720,N_19583,N_19547);
nand U19721 (N_19721,N_19431,N_19515);
or U19722 (N_19722,N_19539,N_19420);
nor U19723 (N_19723,N_19445,N_19576);
nand U19724 (N_19724,N_19485,N_19562);
nor U19725 (N_19725,N_19539,N_19459);
nor U19726 (N_19726,N_19467,N_19521);
or U19727 (N_19727,N_19427,N_19482);
nand U19728 (N_19728,N_19438,N_19598);
or U19729 (N_19729,N_19550,N_19443);
nand U19730 (N_19730,N_19508,N_19445);
nor U19731 (N_19731,N_19488,N_19467);
nand U19732 (N_19732,N_19433,N_19546);
and U19733 (N_19733,N_19560,N_19545);
nand U19734 (N_19734,N_19424,N_19423);
nor U19735 (N_19735,N_19406,N_19454);
nand U19736 (N_19736,N_19576,N_19413);
nand U19737 (N_19737,N_19470,N_19420);
and U19738 (N_19738,N_19439,N_19492);
nor U19739 (N_19739,N_19424,N_19535);
and U19740 (N_19740,N_19473,N_19422);
or U19741 (N_19741,N_19436,N_19401);
nor U19742 (N_19742,N_19510,N_19514);
and U19743 (N_19743,N_19419,N_19401);
nand U19744 (N_19744,N_19528,N_19555);
nor U19745 (N_19745,N_19426,N_19503);
and U19746 (N_19746,N_19474,N_19493);
or U19747 (N_19747,N_19570,N_19486);
nor U19748 (N_19748,N_19426,N_19499);
and U19749 (N_19749,N_19584,N_19522);
nor U19750 (N_19750,N_19584,N_19418);
and U19751 (N_19751,N_19507,N_19495);
and U19752 (N_19752,N_19505,N_19411);
nor U19753 (N_19753,N_19418,N_19567);
nor U19754 (N_19754,N_19568,N_19502);
or U19755 (N_19755,N_19520,N_19545);
nand U19756 (N_19756,N_19527,N_19591);
xor U19757 (N_19757,N_19454,N_19457);
nor U19758 (N_19758,N_19548,N_19546);
nand U19759 (N_19759,N_19411,N_19550);
nor U19760 (N_19760,N_19409,N_19525);
or U19761 (N_19761,N_19553,N_19599);
nand U19762 (N_19762,N_19560,N_19412);
or U19763 (N_19763,N_19486,N_19465);
and U19764 (N_19764,N_19526,N_19500);
and U19765 (N_19765,N_19598,N_19407);
nor U19766 (N_19766,N_19574,N_19412);
nand U19767 (N_19767,N_19499,N_19430);
or U19768 (N_19768,N_19400,N_19542);
or U19769 (N_19769,N_19491,N_19560);
nand U19770 (N_19770,N_19421,N_19508);
and U19771 (N_19771,N_19483,N_19581);
or U19772 (N_19772,N_19465,N_19435);
or U19773 (N_19773,N_19409,N_19424);
or U19774 (N_19774,N_19498,N_19506);
nor U19775 (N_19775,N_19592,N_19515);
or U19776 (N_19776,N_19599,N_19516);
or U19777 (N_19777,N_19561,N_19513);
nand U19778 (N_19778,N_19516,N_19430);
and U19779 (N_19779,N_19507,N_19561);
nor U19780 (N_19780,N_19422,N_19441);
nor U19781 (N_19781,N_19496,N_19483);
nor U19782 (N_19782,N_19518,N_19479);
nor U19783 (N_19783,N_19401,N_19536);
or U19784 (N_19784,N_19533,N_19545);
nor U19785 (N_19785,N_19542,N_19564);
and U19786 (N_19786,N_19468,N_19582);
and U19787 (N_19787,N_19497,N_19528);
or U19788 (N_19788,N_19521,N_19497);
nor U19789 (N_19789,N_19510,N_19405);
or U19790 (N_19790,N_19411,N_19571);
and U19791 (N_19791,N_19432,N_19463);
nor U19792 (N_19792,N_19461,N_19411);
nand U19793 (N_19793,N_19507,N_19484);
or U19794 (N_19794,N_19595,N_19412);
or U19795 (N_19795,N_19570,N_19589);
nand U19796 (N_19796,N_19571,N_19427);
nor U19797 (N_19797,N_19505,N_19563);
nor U19798 (N_19798,N_19436,N_19555);
and U19799 (N_19799,N_19448,N_19486);
nor U19800 (N_19800,N_19703,N_19693);
nor U19801 (N_19801,N_19765,N_19768);
and U19802 (N_19802,N_19780,N_19620);
nor U19803 (N_19803,N_19770,N_19760);
and U19804 (N_19804,N_19719,N_19792);
and U19805 (N_19805,N_19762,N_19680);
or U19806 (N_19806,N_19751,N_19746);
and U19807 (N_19807,N_19646,N_19720);
nand U19808 (N_19808,N_19637,N_19655);
xnor U19809 (N_19809,N_19615,N_19725);
nand U19810 (N_19810,N_19619,N_19748);
or U19811 (N_19811,N_19672,N_19614);
or U19812 (N_19812,N_19629,N_19624);
nor U19813 (N_19813,N_19721,N_19755);
and U19814 (N_19814,N_19658,N_19716);
nor U19815 (N_19815,N_19769,N_19652);
nand U19816 (N_19816,N_19709,N_19666);
nor U19817 (N_19817,N_19722,N_19673);
nand U19818 (N_19818,N_19700,N_19790);
or U19819 (N_19819,N_19698,N_19735);
nor U19820 (N_19820,N_19712,N_19657);
nor U19821 (N_19821,N_19633,N_19627);
nand U19822 (N_19822,N_19718,N_19695);
and U19823 (N_19823,N_19643,N_19608);
nor U19824 (N_19824,N_19617,N_19711);
or U19825 (N_19825,N_19616,N_19640);
and U19826 (N_19826,N_19767,N_19759);
nor U19827 (N_19827,N_19732,N_19649);
nor U19828 (N_19828,N_19723,N_19731);
and U19829 (N_19829,N_19789,N_19682);
nand U19830 (N_19830,N_19650,N_19785);
nand U19831 (N_19831,N_19788,N_19784);
or U19832 (N_19832,N_19795,N_19604);
or U19833 (N_19833,N_19609,N_19744);
nand U19834 (N_19834,N_19713,N_19737);
and U19835 (N_19835,N_19613,N_19674);
and U19836 (N_19836,N_19684,N_19738);
and U19837 (N_19837,N_19661,N_19726);
nor U19838 (N_19838,N_19699,N_19749);
and U19839 (N_19839,N_19696,N_19648);
nor U19840 (N_19840,N_19638,N_19610);
or U19841 (N_19841,N_19662,N_19659);
nor U19842 (N_19842,N_19605,N_19690);
or U19843 (N_19843,N_19777,N_19664);
nor U19844 (N_19844,N_19791,N_19628);
nand U19845 (N_19845,N_19799,N_19741);
nor U19846 (N_19846,N_19641,N_19702);
nand U19847 (N_19847,N_19715,N_19794);
or U19848 (N_19848,N_19773,N_19606);
or U19849 (N_19849,N_19647,N_19639);
and U19850 (N_19850,N_19634,N_19651);
nand U19851 (N_19851,N_19654,N_19714);
nor U19852 (N_19852,N_19603,N_19694);
nor U19853 (N_19853,N_19636,N_19665);
nand U19854 (N_19854,N_19747,N_19697);
and U19855 (N_19855,N_19670,N_19687);
nor U19856 (N_19856,N_19757,N_19685);
nand U19857 (N_19857,N_19623,N_19763);
or U19858 (N_19858,N_19667,N_19754);
or U19859 (N_19859,N_19602,N_19796);
nand U19860 (N_19860,N_19739,N_19752);
and U19861 (N_19861,N_19645,N_19728);
nand U19862 (N_19862,N_19787,N_19668);
and U19863 (N_19863,N_19742,N_19676);
and U19864 (N_19864,N_19675,N_19692);
or U19865 (N_19865,N_19734,N_19771);
nor U19866 (N_19866,N_19793,N_19622);
and U19867 (N_19867,N_19601,N_19660);
or U19868 (N_19868,N_19706,N_19612);
nor U19869 (N_19869,N_19635,N_19669);
nor U19870 (N_19870,N_19733,N_19772);
nand U19871 (N_19871,N_19631,N_19708);
or U19872 (N_19872,N_19764,N_19786);
or U19873 (N_19873,N_19701,N_19724);
nor U19874 (N_19874,N_19766,N_19681);
and U19875 (N_19875,N_19686,N_19797);
nand U19876 (N_19876,N_19678,N_19776);
and U19877 (N_19877,N_19782,N_19679);
or U19878 (N_19878,N_19600,N_19632);
nand U19879 (N_19879,N_19656,N_19621);
and U19880 (N_19880,N_19625,N_19677);
or U19881 (N_19881,N_19642,N_19683);
nand U19882 (N_19882,N_19671,N_19707);
nor U19883 (N_19883,N_19688,N_19781);
and U19884 (N_19884,N_19618,N_19729);
nand U19885 (N_19885,N_19743,N_19710);
and U19886 (N_19886,N_19689,N_19626);
nor U19887 (N_19887,N_19663,N_19630);
or U19888 (N_19888,N_19727,N_19753);
and U19889 (N_19889,N_19653,N_19745);
nand U19890 (N_19890,N_19736,N_19740);
nand U19891 (N_19891,N_19704,N_19644);
and U19892 (N_19892,N_19717,N_19611);
nand U19893 (N_19893,N_19783,N_19691);
or U19894 (N_19894,N_19705,N_19758);
or U19895 (N_19895,N_19778,N_19730);
nand U19896 (N_19896,N_19756,N_19775);
or U19897 (N_19897,N_19774,N_19761);
and U19898 (N_19898,N_19607,N_19750);
or U19899 (N_19899,N_19779,N_19798);
or U19900 (N_19900,N_19720,N_19616);
nor U19901 (N_19901,N_19783,N_19718);
nor U19902 (N_19902,N_19639,N_19677);
nor U19903 (N_19903,N_19727,N_19606);
and U19904 (N_19904,N_19702,N_19705);
nand U19905 (N_19905,N_19648,N_19765);
and U19906 (N_19906,N_19792,N_19715);
nor U19907 (N_19907,N_19679,N_19674);
nor U19908 (N_19908,N_19619,N_19642);
and U19909 (N_19909,N_19677,N_19688);
or U19910 (N_19910,N_19743,N_19665);
and U19911 (N_19911,N_19768,N_19648);
or U19912 (N_19912,N_19682,N_19672);
and U19913 (N_19913,N_19720,N_19680);
or U19914 (N_19914,N_19644,N_19617);
and U19915 (N_19915,N_19680,N_19633);
or U19916 (N_19916,N_19640,N_19774);
or U19917 (N_19917,N_19695,N_19639);
and U19918 (N_19918,N_19683,N_19749);
and U19919 (N_19919,N_19659,N_19656);
nor U19920 (N_19920,N_19697,N_19766);
nand U19921 (N_19921,N_19650,N_19610);
nor U19922 (N_19922,N_19792,N_19629);
and U19923 (N_19923,N_19769,N_19622);
nand U19924 (N_19924,N_19726,N_19698);
nand U19925 (N_19925,N_19690,N_19771);
nand U19926 (N_19926,N_19755,N_19713);
and U19927 (N_19927,N_19729,N_19771);
and U19928 (N_19928,N_19797,N_19722);
nand U19929 (N_19929,N_19654,N_19636);
nor U19930 (N_19930,N_19608,N_19675);
nor U19931 (N_19931,N_19728,N_19643);
and U19932 (N_19932,N_19686,N_19637);
or U19933 (N_19933,N_19757,N_19639);
or U19934 (N_19934,N_19731,N_19734);
and U19935 (N_19935,N_19656,N_19671);
or U19936 (N_19936,N_19631,N_19621);
nor U19937 (N_19937,N_19747,N_19672);
or U19938 (N_19938,N_19711,N_19754);
or U19939 (N_19939,N_19767,N_19782);
and U19940 (N_19940,N_19673,N_19717);
nand U19941 (N_19941,N_19670,N_19656);
nand U19942 (N_19942,N_19643,N_19659);
and U19943 (N_19943,N_19641,N_19695);
and U19944 (N_19944,N_19603,N_19740);
or U19945 (N_19945,N_19657,N_19680);
nand U19946 (N_19946,N_19716,N_19685);
and U19947 (N_19947,N_19672,N_19769);
and U19948 (N_19948,N_19738,N_19799);
nand U19949 (N_19949,N_19797,N_19756);
nor U19950 (N_19950,N_19659,N_19681);
nor U19951 (N_19951,N_19661,N_19759);
nor U19952 (N_19952,N_19756,N_19632);
nand U19953 (N_19953,N_19762,N_19614);
or U19954 (N_19954,N_19738,N_19640);
or U19955 (N_19955,N_19781,N_19760);
nor U19956 (N_19956,N_19783,N_19612);
and U19957 (N_19957,N_19713,N_19798);
nor U19958 (N_19958,N_19665,N_19718);
nor U19959 (N_19959,N_19744,N_19783);
or U19960 (N_19960,N_19696,N_19753);
and U19961 (N_19961,N_19685,N_19614);
and U19962 (N_19962,N_19687,N_19784);
and U19963 (N_19963,N_19781,N_19603);
and U19964 (N_19964,N_19639,N_19787);
or U19965 (N_19965,N_19687,N_19718);
nand U19966 (N_19966,N_19668,N_19786);
and U19967 (N_19967,N_19690,N_19630);
nand U19968 (N_19968,N_19655,N_19750);
or U19969 (N_19969,N_19797,N_19684);
nand U19970 (N_19970,N_19766,N_19789);
nor U19971 (N_19971,N_19670,N_19633);
or U19972 (N_19972,N_19661,N_19607);
nand U19973 (N_19973,N_19701,N_19668);
and U19974 (N_19974,N_19641,N_19749);
and U19975 (N_19975,N_19608,N_19741);
nand U19976 (N_19976,N_19772,N_19669);
and U19977 (N_19977,N_19751,N_19711);
and U19978 (N_19978,N_19737,N_19719);
or U19979 (N_19979,N_19766,N_19774);
nor U19980 (N_19980,N_19606,N_19631);
or U19981 (N_19981,N_19756,N_19680);
and U19982 (N_19982,N_19636,N_19653);
nor U19983 (N_19983,N_19690,N_19654);
nor U19984 (N_19984,N_19748,N_19734);
or U19985 (N_19985,N_19797,N_19663);
nand U19986 (N_19986,N_19693,N_19749);
and U19987 (N_19987,N_19638,N_19643);
nand U19988 (N_19988,N_19626,N_19630);
nand U19989 (N_19989,N_19675,N_19696);
and U19990 (N_19990,N_19628,N_19680);
or U19991 (N_19991,N_19759,N_19728);
and U19992 (N_19992,N_19601,N_19748);
nand U19993 (N_19993,N_19617,N_19741);
nor U19994 (N_19994,N_19748,N_19770);
and U19995 (N_19995,N_19667,N_19779);
nor U19996 (N_19996,N_19717,N_19693);
and U19997 (N_19997,N_19703,N_19694);
nand U19998 (N_19998,N_19607,N_19606);
nand U19999 (N_19999,N_19673,N_19788);
and UO_0 (O_0,N_19941,N_19872);
or UO_1 (O_1,N_19972,N_19958);
nor UO_2 (O_2,N_19846,N_19829);
or UO_3 (O_3,N_19983,N_19924);
nor UO_4 (O_4,N_19892,N_19848);
nand UO_5 (O_5,N_19805,N_19912);
and UO_6 (O_6,N_19841,N_19957);
nand UO_7 (O_7,N_19979,N_19899);
or UO_8 (O_8,N_19859,N_19951);
and UO_9 (O_9,N_19923,N_19948);
nor UO_10 (O_10,N_19894,N_19930);
and UO_11 (O_11,N_19882,N_19967);
and UO_12 (O_12,N_19952,N_19936);
nor UO_13 (O_13,N_19934,N_19993);
nand UO_14 (O_14,N_19835,N_19870);
or UO_15 (O_15,N_19836,N_19854);
and UO_16 (O_16,N_19898,N_19911);
and UO_17 (O_17,N_19864,N_19804);
and UO_18 (O_18,N_19878,N_19927);
or UO_19 (O_19,N_19820,N_19896);
or UO_20 (O_20,N_19996,N_19965);
and UO_21 (O_21,N_19974,N_19862);
and UO_22 (O_22,N_19840,N_19945);
and UO_23 (O_23,N_19918,N_19831);
nand UO_24 (O_24,N_19909,N_19869);
nor UO_25 (O_25,N_19984,N_19976);
nor UO_26 (O_26,N_19943,N_19937);
and UO_27 (O_27,N_19959,N_19853);
or UO_28 (O_28,N_19814,N_19906);
or UO_29 (O_29,N_19889,N_19931);
nand UO_30 (O_30,N_19816,N_19887);
and UO_31 (O_31,N_19802,N_19933);
or UO_32 (O_32,N_19962,N_19865);
nor UO_33 (O_33,N_19975,N_19947);
nor UO_34 (O_34,N_19886,N_19818);
or UO_35 (O_35,N_19877,N_19997);
and UO_36 (O_36,N_19832,N_19895);
nand UO_37 (O_37,N_19910,N_19830);
or UO_38 (O_38,N_19966,N_19833);
nand UO_39 (O_39,N_19985,N_19860);
nand UO_40 (O_40,N_19817,N_19914);
and UO_41 (O_41,N_19987,N_19970);
nor UO_42 (O_42,N_19956,N_19935);
or UO_43 (O_43,N_19903,N_19990);
nor UO_44 (O_44,N_19982,N_19824);
and UO_45 (O_45,N_19961,N_19954);
nand UO_46 (O_46,N_19857,N_19850);
nor UO_47 (O_47,N_19808,N_19999);
or UO_48 (O_48,N_19938,N_19916);
nor UO_49 (O_49,N_19867,N_19880);
or UO_50 (O_50,N_19893,N_19875);
and UO_51 (O_51,N_19838,N_19825);
nand UO_52 (O_52,N_19807,N_19849);
nand UO_53 (O_53,N_19828,N_19968);
and UO_54 (O_54,N_19939,N_19823);
or UO_55 (O_55,N_19991,N_19842);
nand UO_56 (O_56,N_19811,N_19843);
nand UO_57 (O_57,N_19855,N_19815);
and UO_58 (O_58,N_19921,N_19913);
or UO_59 (O_59,N_19977,N_19980);
and UO_60 (O_60,N_19922,N_19803);
or UO_61 (O_61,N_19800,N_19940);
nor UO_62 (O_62,N_19928,N_19866);
xnor UO_63 (O_63,N_19873,N_19981);
or UO_64 (O_64,N_19891,N_19876);
or UO_65 (O_65,N_19858,N_19801);
nor UO_66 (O_66,N_19821,N_19847);
nand UO_67 (O_67,N_19863,N_19953);
or UO_68 (O_68,N_19908,N_19890);
nor UO_69 (O_69,N_19874,N_19994);
nand UO_70 (O_70,N_19856,N_19950);
and UO_71 (O_71,N_19907,N_19915);
and UO_72 (O_72,N_19809,N_19920);
nand UO_73 (O_73,N_19988,N_19963);
nand UO_74 (O_74,N_19837,N_19926);
nor UO_75 (O_75,N_19885,N_19844);
nand UO_76 (O_76,N_19971,N_19810);
or UO_77 (O_77,N_19826,N_19955);
nor UO_78 (O_78,N_19812,N_19905);
nand UO_79 (O_79,N_19932,N_19861);
nand UO_80 (O_80,N_19897,N_19884);
nor UO_81 (O_81,N_19883,N_19998);
and UO_82 (O_82,N_19944,N_19827);
or UO_83 (O_83,N_19919,N_19960);
or UO_84 (O_84,N_19851,N_19946);
and UO_85 (O_85,N_19995,N_19879);
and UO_86 (O_86,N_19964,N_19868);
and UO_87 (O_87,N_19902,N_19917);
and UO_88 (O_88,N_19839,N_19806);
or UO_89 (O_89,N_19819,N_19949);
nor UO_90 (O_90,N_19901,N_19969);
nor UO_91 (O_91,N_19834,N_19925);
and UO_92 (O_92,N_19871,N_19904);
and UO_93 (O_93,N_19978,N_19881);
nand UO_94 (O_94,N_19852,N_19992);
nand UO_95 (O_95,N_19942,N_19900);
nand UO_96 (O_96,N_19929,N_19888);
nand UO_97 (O_97,N_19822,N_19986);
nor UO_98 (O_98,N_19845,N_19989);
nor UO_99 (O_99,N_19973,N_19813);
nor UO_100 (O_100,N_19856,N_19846);
nand UO_101 (O_101,N_19883,N_19865);
and UO_102 (O_102,N_19931,N_19920);
or UO_103 (O_103,N_19863,N_19985);
and UO_104 (O_104,N_19916,N_19977);
or UO_105 (O_105,N_19804,N_19830);
and UO_106 (O_106,N_19918,N_19855);
nand UO_107 (O_107,N_19996,N_19876);
nand UO_108 (O_108,N_19983,N_19963);
and UO_109 (O_109,N_19841,N_19892);
nor UO_110 (O_110,N_19843,N_19809);
or UO_111 (O_111,N_19862,N_19928);
nor UO_112 (O_112,N_19877,N_19810);
and UO_113 (O_113,N_19918,N_19888);
and UO_114 (O_114,N_19827,N_19931);
and UO_115 (O_115,N_19868,N_19883);
nand UO_116 (O_116,N_19828,N_19800);
or UO_117 (O_117,N_19928,N_19964);
or UO_118 (O_118,N_19997,N_19832);
and UO_119 (O_119,N_19969,N_19930);
and UO_120 (O_120,N_19821,N_19900);
or UO_121 (O_121,N_19898,N_19830);
and UO_122 (O_122,N_19945,N_19985);
nor UO_123 (O_123,N_19870,N_19944);
and UO_124 (O_124,N_19808,N_19981);
nor UO_125 (O_125,N_19940,N_19923);
nand UO_126 (O_126,N_19800,N_19879);
nor UO_127 (O_127,N_19867,N_19828);
and UO_128 (O_128,N_19811,N_19913);
nand UO_129 (O_129,N_19805,N_19946);
or UO_130 (O_130,N_19916,N_19861);
and UO_131 (O_131,N_19944,N_19850);
or UO_132 (O_132,N_19833,N_19873);
nand UO_133 (O_133,N_19808,N_19819);
or UO_134 (O_134,N_19941,N_19809);
nand UO_135 (O_135,N_19888,N_19825);
and UO_136 (O_136,N_19917,N_19957);
nor UO_137 (O_137,N_19957,N_19918);
or UO_138 (O_138,N_19915,N_19843);
or UO_139 (O_139,N_19808,N_19851);
nand UO_140 (O_140,N_19884,N_19802);
and UO_141 (O_141,N_19981,N_19819);
and UO_142 (O_142,N_19978,N_19865);
nor UO_143 (O_143,N_19959,N_19965);
or UO_144 (O_144,N_19885,N_19975);
or UO_145 (O_145,N_19886,N_19942);
or UO_146 (O_146,N_19988,N_19900);
nor UO_147 (O_147,N_19866,N_19850);
nand UO_148 (O_148,N_19847,N_19865);
or UO_149 (O_149,N_19996,N_19823);
or UO_150 (O_150,N_19900,N_19911);
nand UO_151 (O_151,N_19863,N_19977);
nor UO_152 (O_152,N_19945,N_19845);
or UO_153 (O_153,N_19914,N_19975);
or UO_154 (O_154,N_19930,N_19964);
or UO_155 (O_155,N_19932,N_19874);
or UO_156 (O_156,N_19956,N_19906);
nand UO_157 (O_157,N_19816,N_19978);
nor UO_158 (O_158,N_19943,N_19888);
nand UO_159 (O_159,N_19892,N_19832);
and UO_160 (O_160,N_19914,N_19957);
nor UO_161 (O_161,N_19909,N_19809);
xor UO_162 (O_162,N_19931,N_19982);
or UO_163 (O_163,N_19975,N_19971);
nand UO_164 (O_164,N_19857,N_19879);
nand UO_165 (O_165,N_19846,N_19881);
nand UO_166 (O_166,N_19930,N_19895);
nor UO_167 (O_167,N_19812,N_19931);
and UO_168 (O_168,N_19948,N_19989);
and UO_169 (O_169,N_19924,N_19914);
and UO_170 (O_170,N_19845,N_19949);
nor UO_171 (O_171,N_19855,N_19831);
nor UO_172 (O_172,N_19926,N_19898);
or UO_173 (O_173,N_19963,N_19989);
nand UO_174 (O_174,N_19817,N_19950);
or UO_175 (O_175,N_19813,N_19809);
nor UO_176 (O_176,N_19945,N_19871);
nor UO_177 (O_177,N_19907,N_19950);
nand UO_178 (O_178,N_19902,N_19806);
nor UO_179 (O_179,N_19989,N_19901);
nand UO_180 (O_180,N_19845,N_19865);
and UO_181 (O_181,N_19990,N_19892);
and UO_182 (O_182,N_19985,N_19824);
nor UO_183 (O_183,N_19923,N_19832);
and UO_184 (O_184,N_19915,N_19810);
and UO_185 (O_185,N_19840,N_19998);
nor UO_186 (O_186,N_19936,N_19988);
nand UO_187 (O_187,N_19894,N_19910);
and UO_188 (O_188,N_19947,N_19921);
nand UO_189 (O_189,N_19905,N_19889);
or UO_190 (O_190,N_19926,N_19960);
and UO_191 (O_191,N_19991,N_19959);
or UO_192 (O_192,N_19808,N_19894);
nand UO_193 (O_193,N_19884,N_19808);
nor UO_194 (O_194,N_19804,N_19993);
or UO_195 (O_195,N_19873,N_19835);
or UO_196 (O_196,N_19900,N_19938);
nand UO_197 (O_197,N_19866,N_19983);
nor UO_198 (O_198,N_19830,N_19837);
or UO_199 (O_199,N_19987,N_19855);
and UO_200 (O_200,N_19812,N_19858);
nor UO_201 (O_201,N_19950,N_19937);
nand UO_202 (O_202,N_19943,N_19805);
nand UO_203 (O_203,N_19890,N_19905);
nor UO_204 (O_204,N_19936,N_19995);
nor UO_205 (O_205,N_19867,N_19843);
nand UO_206 (O_206,N_19839,N_19866);
nand UO_207 (O_207,N_19982,N_19918);
nor UO_208 (O_208,N_19890,N_19999);
nand UO_209 (O_209,N_19913,N_19862);
nand UO_210 (O_210,N_19920,N_19970);
and UO_211 (O_211,N_19822,N_19896);
or UO_212 (O_212,N_19932,N_19807);
or UO_213 (O_213,N_19802,N_19854);
nand UO_214 (O_214,N_19986,N_19984);
nand UO_215 (O_215,N_19810,N_19972);
or UO_216 (O_216,N_19849,N_19962);
nand UO_217 (O_217,N_19831,N_19975);
and UO_218 (O_218,N_19843,N_19807);
and UO_219 (O_219,N_19833,N_19895);
nand UO_220 (O_220,N_19911,N_19830);
nand UO_221 (O_221,N_19843,N_19881);
and UO_222 (O_222,N_19822,N_19860);
nor UO_223 (O_223,N_19877,N_19949);
or UO_224 (O_224,N_19969,N_19851);
or UO_225 (O_225,N_19888,N_19873);
xnor UO_226 (O_226,N_19906,N_19809);
or UO_227 (O_227,N_19828,N_19817);
and UO_228 (O_228,N_19873,N_19942);
and UO_229 (O_229,N_19840,N_19979);
and UO_230 (O_230,N_19948,N_19971);
xnor UO_231 (O_231,N_19996,N_19966);
or UO_232 (O_232,N_19942,N_19829);
xor UO_233 (O_233,N_19896,N_19835);
and UO_234 (O_234,N_19897,N_19888);
nor UO_235 (O_235,N_19841,N_19829);
nand UO_236 (O_236,N_19988,N_19990);
and UO_237 (O_237,N_19908,N_19922);
nand UO_238 (O_238,N_19807,N_19841);
nand UO_239 (O_239,N_19801,N_19946);
nor UO_240 (O_240,N_19826,N_19883);
or UO_241 (O_241,N_19860,N_19853);
and UO_242 (O_242,N_19975,N_19861);
or UO_243 (O_243,N_19987,N_19800);
nor UO_244 (O_244,N_19868,N_19847);
or UO_245 (O_245,N_19889,N_19846);
nor UO_246 (O_246,N_19908,N_19983);
and UO_247 (O_247,N_19823,N_19997);
nand UO_248 (O_248,N_19867,N_19899);
xor UO_249 (O_249,N_19871,N_19837);
and UO_250 (O_250,N_19910,N_19945);
nor UO_251 (O_251,N_19885,N_19821);
and UO_252 (O_252,N_19882,N_19846);
and UO_253 (O_253,N_19937,N_19964);
nand UO_254 (O_254,N_19949,N_19879);
and UO_255 (O_255,N_19917,N_19980);
or UO_256 (O_256,N_19976,N_19912);
and UO_257 (O_257,N_19834,N_19910);
nor UO_258 (O_258,N_19997,N_19827);
and UO_259 (O_259,N_19909,N_19913);
or UO_260 (O_260,N_19836,N_19959);
nand UO_261 (O_261,N_19882,N_19930);
nand UO_262 (O_262,N_19874,N_19996);
nand UO_263 (O_263,N_19897,N_19995);
nand UO_264 (O_264,N_19824,N_19986);
nand UO_265 (O_265,N_19826,N_19939);
nand UO_266 (O_266,N_19931,N_19945);
or UO_267 (O_267,N_19867,N_19987);
or UO_268 (O_268,N_19932,N_19864);
xor UO_269 (O_269,N_19880,N_19892);
or UO_270 (O_270,N_19806,N_19985);
and UO_271 (O_271,N_19856,N_19911);
nand UO_272 (O_272,N_19926,N_19930);
nor UO_273 (O_273,N_19858,N_19906);
or UO_274 (O_274,N_19888,N_19854);
nor UO_275 (O_275,N_19813,N_19904);
nor UO_276 (O_276,N_19846,N_19869);
and UO_277 (O_277,N_19893,N_19865);
or UO_278 (O_278,N_19860,N_19895);
or UO_279 (O_279,N_19857,N_19889);
and UO_280 (O_280,N_19925,N_19963);
nor UO_281 (O_281,N_19937,N_19811);
nor UO_282 (O_282,N_19841,N_19913);
and UO_283 (O_283,N_19912,N_19921);
nor UO_284 (O_284,N_19870,N_19919);
nor UO_285 (O_285,N_19915,N_19875);
nor UO_286 (O_286,N_19817,N_19909);
nand UO_287 (O_287,N_19969,N_19955);
nor UO_288 (O_288,N_19825,N_19881);
and UO_289 (O_289,N_19886,N_19810);
xor UO_290 (O_290,N_19974,N_19880);
and UO_291 (O_291,N_19814,N_19853);
nor UO_292 (O_292,N_19914,N_19965);
nor UO_293 (O_293,N_19950,N_19967);
nand UO_294 (O_294,N_19882,N_19983);
nand UO_295 (O_295,N_19958,N_19898);
nand UO_296 (O_296,N_19959,N_19810);
nand UO_297 (O_297,N_19877,N_19986);
or UO_298 (O_298,N_19899,N_19855);
xnor UO_299 (O_299,N_19920,N_19952);
or UO_300 (O_300,N_19924,N_19838);
nand UO_301 (O_301,N_19867,N_19834);
and UO_302 (O_302,N_19806,N_19800);
and UO_303 (O_303,N_19890,N_19988);
and UO_304 (O_304,N_19926,N_19992);
nor UO_305 (O_305,N_19905,N_19990);
nand UO_306 (O_306,N_19943,N_19857);
nand UO_307 (O_307,N_19831,N_19908);
nand UO_308 (O_308,N_19833,N_19935);
and UO_309 (O_309,N_19840,N_19932);
nand UO_310 (O_310,N_19845,N_19834);
nor UO_311 (O_311,N_19877,N_19874);
and UO_312 (O_312,N_19812,N_19857);
nand UO_313 (O_313,N_19993,N_19972);
nand UO_314 (O_314,N_19859,N_19827);
nor UO_315 (O_315,N_19886,N_19831);
nor UO_316 (O_316,N_19893,N_19880);
nor UO_317 (O_317,N_19814,N_19818);
or UO_318 (O_318,N_19835,N_19906);
xnor UO_319 (O_319,N_19843,N_19888);
nand UO_320 (O_320,N_19811,N_19918);
nand UO_321 (O_321,N_19881,N_19926);
nor UO_322 (O_322,N_19858,N_19888);
nand UO_323 (O_323,N_19950,N_19989);
or UO_324 (O_324,N_19801,N_19942);
nand UO_325 (O_325,N_19872,N_19827);
or UO_326 (O_326,N_19887,N_19936);
and UO_327 (O_327,N_19863,N_19907);
or UO_328 (O_328,N_19807,N_19820);
and UO_329 (O_329,N_19841,N_19835);
or UO_330 (O_330,N_19862,N_19907);
nor UO_331 (O_331,N_19923,N_19833);
nand UO_332 (O_332,N_19969,N_19946);
or UO_333 (O_333,N_19901,N_19829);
nand UO_334 (O_334,N_19936,N_19858);
nand UO_335 (O_335,N_19919,N_19820);
nand UO_336 (O_336,N_19924,N_19884);
or UO_337 (O_337,N_19974,N_19832);
and UO_338 (O_338,N_19843,N_19891);
or UO_339 (O_339,N_19999,N_19933);
and UO_340 (O_340,N_19863,N_19855);
nand UO_341 (O_341,N_19878,N_19810);
nand UO_342 (O_342,N_19874,N_19835);
nand UO_343 (O_343,N_19857,N_19885);
and UO_344 (O_344,N_19912,N_19849);
nand UO_345 (O_345,N_19983,N_19967);
nand UO_346 (O_346,N_19959,N_19862);
nor UO_347 (O_347,N_19993,N_19854);
nor UO_348 (O_348,N_19895,N_19910);
and UO_349 (O_349,N_19993,N_19847);
and UO_350 (O_350,N_19884,N_19928);
nand UO_351 (O_351,N_19844,N_19851);
nand UO_352 (O_352,N_19974,N_19908);
and UO_353 (O_353,N_19998,N_19905);
and UO_354 (O_354,N_19852,N_19810);
or UO_355 (O_355,N_19991,N_19940);
nand UO_356 (O_356,N_19813,N_19876);
and UO_357 (O_357,N_19860,N_19949);
nor UO_358 (O_358,N_19836,N_19990);
nor UO_359 (O_359,N_19888,N_19848);
and UO_360 (O_360,N_19867,N_19824);
nor UO_361 (O_361,N_19844,N_19984);
and UO_362 (O_362,N_19849,N_19855);
nor UO_363 (O_363,N_19915,N_19923);
or UO_364 (O_364,N_19917,N_19863);
nand UO_365 (O_365,N_19964,N_19820);
nand UO_366 (O_366,N_19884,N_19989);
nand UO_367 (O_367,N_19951,N_19850);
nor UO_368 (O_368,N_19812,N_19970);
or UO_369 (O_369,N_19932,N_19934);
nand UO_370 (O_370,N_19850,N_19997);
nand UO_371 (O_371,N_19925,N_19919);
nand UO_372 (O_372,N_19914,N_19941);
and UO_373 (O_373,N_19981,N_19913);
nand UO_374 (O_374,N_19849,N_19913);
nand UO_375 (O_375,N_19814,N_19839);
and UO_376 (O_376,N_19816,N_19896);
nand UO_377 (O_377,N_19816,N_19811);
and UO_378 (O_378,N_19934,N_19911);
nor UO_379 (O_379,N_19926,N_19808);
nor UO_380 (O_380,N_19924,N_19919);
and UO_381 (O_381,N_19963,N_19911);
or UO_382 (O_382,N_19805,N_19861);
and UO_383 (O_383,N_19880,N_19825);
and UO_384 (O_384,N_19858,N_19919);
and UO_385 (O_385,N_19934,N_19844);
or UO_386 (O_386,N_19865,N_19984);
and UO_387 (O_387,N_19810,N_19887);
and UO_388 (O_388,N_19841,N_19891);
and UO_389 (O_389,N_19858,N_19931);
nand UO_390 (O_390,N_19982,N_19894);
and UO_391 (O_391,N_19882,N_19920);
nand UO_392 (O_392,N_19908,N_19907);
nor UO_393 (O_393,N_19813,N_19984);
or UO_394 (O_394,N_19838,N_19907);
nand UO_395 (O_395,N_19886,N_19927);
nand UO_396 (O_396,N_19877,N_19826);
or UO_397 (O_397,N_19821,N_19969);
and UO_398 (O_398,N_19894,N_19887);
nor UO_399 (O_399,N_19852,N_19998);
nand UO_400 (O_400,N_19883,N_19846);
or UO_401 (O_401,N_19906,N_19839);
nand UO_402 (O_402,N_19977,N_19800);
and UO_403 (O_403,N_19945,N_19802);
and UO_404 (O_404,N_19999,N_19810);
nor UO_405 (O_405,N_19878,N_19919);
and UO_406 (O_406,N_19885,N_19995);
or UO_407 (O_407,N_19836,N_19986);
or UO_408 (O_408,N_19842,N_19834);
nor UO_409 (O_409,N_19816,N_19947);
or UO_410 (O_410,N_19825,N_19855);
nand UO_411 (O_411,N_19895,N_19837);
nor UO_412 (O_412,N_19955,N_19984);
nor UO_413 (O_413,N_19854,N_19918);
or UO_414 (O_414,N_19894,N_19881);
and UO_415 (O_415,N_19947,N_19919);
and UO_416 (O_416,N_19899,N_19950);
nand UO_417 (O_417,N_19873,N_19866);
or UO_418 (O_418,N_19942,N_19825);
nand UO_419 (O_419,N_19826,N_19876);
nand UO_420 (O_420,N_19904,N_19852);
or UO_421 (O_421,N_19958,N_19838);
nand UO_422 (O_422,N_19864,N_19820);
nor UO_423 (O_423,N_19985,N_19894);
and UO_424 (O_424,N_19903,N_19834);
or UO_425 (O_425,N_19858,N_19904);
nor UO_426 (O_426,N_19840,N_19879);
or UO_427 (O_427,N_19952,N_19899);
nand UO_428 (O_428,N_19812,N_19979);
nor UO_429 (O_429,N_19996,N_19837);
nand UO_430 (O_430,N_19898,N_19906);
or UO_431 (O_431,N_19929,N_19931);
or UO_432 (O_432,N_19840,N_19833);
or UO_433 (O_433,N_19990,N_19854);
nor UO_434 (O_434,N_19851,N_19823);
or UO_435 (O_435,N_19891,N_19990);
and UO_436 (O_436,N_19923,N_19825);
nand UO_437 (O_437,N_19825,N_19863);
or UO_438 (O_438,N_19979,N_19876);
and UO_439 (O_439,N_19880,N_19866);
or UO_440 (O_440,N_19846,N_19929);
or UO_441 (O_441,N_19877,N_19929);
and UO_442 (O_442,N_19923,N_19891);
and UO_443 (O_443,N_19881,N_19955);
or UO_444 (O_444,N_19813,N_19915);
or UO_445 (O_445,N_19885,N_19917);
or UO_446 (O_446,N_19841,N_19908);
nand UO_447 (O_447,N_19962,N_19810);
nor UO_448 (O_448,N_19824,N_19951);
or UO_449 (O_449,N_19859,N_19867);
nand UO_450 (O_450,N_19991,N_19938);
nand UO_451 (O_451,N_19891,N_19877);
nand UO_452 (O_452,N_19977,N_19826);
nor UO_453 (O_453,N_19938,N_19891);
and UO_454 (O_454,N_19957,N_19978);
or UO_455 (O_455,N_19820,N_19986);
nand UO_456 (O_456,N_19842,N_19802);
nand UO_457 (O_457,N_19939,N_19806);
or UO_458 (O_458,N_19919,N_19818);
nor UO_459 (O_459,N_19845,N_19913);
and UO_460 (O_460,N_19996,N_19805);
or UO_461 (O_461,N_19855,N_19904);
or UO_462 (O_462,N_19917,N_19913);
and UO_463 (O_463,N_19815,N_19942);
or UO_464 (O_464,N_19960,N_19901);
or UO_465 (O_465,N_19944,N_19972);
nor UO_466 (O_466,N_19830,N_19870);
nor UO_467 (O_467,N_19943,N_19955);
or UO_468 (O_468,N_19947,N_19993);
nand UO_469 (O_469,N_19850,N_19846);
nor UO_470 (O_470,N_19865,N_19937);
and UO_471 (O_471,N_19810,N_19836);
and UO_472 (O_472,N_19818,N_19925);
nand UO_473 (O_473,N_19925,N_19904);
nand UO_474 (O_474,N_19951,N_19846);
nand UO_475 (O_475,N_19844,N_19834);
and UO_476 (O_476,N_19995,N_19872);
or UO_477 (O_477,N_19993,N_19878);
nand UO_478 (O_478,N_19849,N_19862);
nor UO_479 (O_479,N_19832,N_19950);
nand UO_480 (O_480,N_19969,N_19833);
and UO_481 (O_481,N_19854,N_19816);
and UO_482 (O_482,N_19960,N_19929);
nor UO_483 (O_483,N_19987,N_19962);
nand UO_484 (O_484,N_19800,N_19849);
nand UO_485 (O_485,N_19914,N_19936);
xor UO_486 (O_486,N_19981,N_19901);
or UO_487 (O_487,N_19962,N_19893);
nand UO_488 (O_488,N_19814,N_19874);
or UO_489 (O_489,N_19836,N_19878);
nor UO_490 (O_490,N_19974,N_19939);
nand UO_491 (O_491,N_19946,N_19925);
nand UO_492 (O_492,N_19900,N_19978);
nand UO_493 (O_493,N_19826,N_19889);
or UO_494 (O_494,N_19830,N_19871);
or UO_495 (O_495,N_19997,N_19963);
nor UO_496 (O_496,N_19855,N_19898);
and UO_497 (O_497,N_19874,N_19804);
and UO_498 (O_498,N_19967,N_19836);
nor UO_499 (O_499,N_19930,N_19965);
and UO_500 (O_500,N_19879,N_19832);
nand UO_501 (O_501,N_19874,N_19806);
nor UO_502 (O_502,N_19890,N_19934);
nand UO_503 (O_503,N_19981,N_19844);
nand UO_504 (O_504,N_19959,N_19930);
or UO_505 (O_505,N_19849,N_19863);
nand UO_506 (O_506,N_19999,N_19976);
nand UO_507 (O_507,N_19811,N_19980);
nand UO_508 (O_508,N_19945,N_19938);
nand UO_509 (O_509,N_19922,N_19919);
and UO_510 (O_510,N_19962,N_19982);
and UO_511 (O_511,N_19852,N_19818);
nand UO_512 (O_512,N_19818,N_19839);
or UO_513 (O_513,N_19858,N_19887);
xor UO_514 (O_514,N_19826,N_19923);
or UO_515 (O_515,N_19804,N_19817);
and UO_516 (O_516,N_19948,N_19831);
or UO_517 (O_517,N_19947,N_19958);
nor UO_518 (O_518,N_19991,N_19827);
nand UO_519 (O_519,N_19954,N_19892);
nor UO_520 (O_520,N_19913,N_19930);
or UO_521 (O_521,N_19912,N_19818);
and UO_522 (O_522,N_19863,N_19807);
nor UO_523 (O_523,N_19889,N_19993);
or UO_524 (O_524,N_19993,N_19841);
and UO_525 (O_525,N_19965,N_19972);
and UO_526 (O_526,N_19817,N_19902);
nand UO_527 (O_527,N_19992,N_19962);
or UO_528 (O_528,N_19862,N_19935);
or UO_529 (O_529,N_19882,N_19884);
and UO_530 (O_530,N_19881,N_19924);
or UO_531 (O_531,N_19880,N_19878);
or UO_532 (O_532,N_19947,N_19933);
and UO_533 (O_533,N_19966,N_19997);
and UO_534 (O_534,N_19962,N_19952);
nand UO_535 (O_535,N_19904,N_19910);
and UO_536 (O_536,N_19899,N_19997);
or UO_537 (O_537,N_19977,N_19892);
and UO_538 (O_538,N_19849,N_19846);
nor UO_539 (O_539,N_19995,N_19899);
nand UO_540 (O_540,N_19815,N_19837);
nand UO_541 (O_541,N_19903,N_19977);
nand UO_542 (O_542,N_19855,N_19913);
or UO_543 (O_543,N_19918,N_19876);
nor UO_544 (O_544,N_19881,N_19806);
nor UO_545 (O_545,N_19855,N_19912);
nand UO_546 (O_546,N_19964,N_19949);
and UO_547 (O_547,N_19998,N_19958);
and UO_548 (O_548,N_19867,N_19974);
or UO_549 (O_549,N_19980,N_19869);
or UO_550 (O_550,N_19803,N_19991);
and UO_551 (O_551,N_19828,N_19881);
nand UO_552 (O_552,N_19864,N_19973);
or UO_553 (O_553,N_19997,N_19803);
or UO_554 (O_554,N_19852,N_19937);
or UO_555 (O_555,N_19909,N_19981);
nand UO_556 (O_556,N_19963,N_19894);
or UO_557 (O_557,N_19883,N_19967);
nand UO_558 (O_558,N_19835,N_19920);
and UO_559 (O_559,N_19962,N_19889);
nand UO_560 (O_560,N_19923,N_19855);
nor UO_561 (O_561,N_19909,N_19942);
and UO_562 (O_562,N_19869,N_19867);
nor UO_563 (O_563,N_19941,N_19939);
nor UO_564 (O_564,N_19998,N_19899);
nor UO_565 (O_565,N_19900,N_19889);
and UO_566 (O_566,N_19807,N_19855);
and UO_567 (O_567,N_19930,N_19967);
and UO_568 (O_568,N_19938,N_19930);
nor UO_569 (O_569,N_19930,N_19966);
or UO_570 (O_570,N_19837,N_19861);
nand UO_571 (O_571,N_19914,N_19821);
nand UO_572 (O_572,N_19826,N_19987);
or UO_573 (O_573,N_19897,N_19868);
nand UO_574 (O_574,N_19872,N_19939);
nor UO_575 (O_575,N_19874,N_19896);
or UO_576 (O_576,N_19917,N_19858);
nor UO_577 (O_577,N_19931,N_19887);
and UO_578 (O_578,N_19926,N_19873);
or UO_579 (O_579,N_19936,N_19921);
or UO_580 (O_580,N_19910,N_19969);
nand UO_581 (O_581,N_19963,N_19979);
or UO_582 (O_582,N_19911,N_19839);
or UO_583 (O_583,N_19936,N_19870);
nor UO_584 (O_584,N_19926,N_19983);
nand UO_585 (O_585,N_19900,N_19865);
nand UO_586 (O_586,N_19833,N_19816);
nand UO_587 (O_587,N_19864,N_19831);
or UO_588 (O_588,N_19852,N_19975);
nor UO_589 (O_589,N_19867,N_19881);
nor UO_590 (O_590,N_19800,N_19982);
nor UO_591 (O_591,N_19889,N_19949);
nand UO_592 (O_592,N_19965,N_19874);
nor UO_593 (O_593,N_19815,N_19895);
xnor UO_594 (O_594,N_19870,N_19833);
nand UO_595 (O_595,N_19830,N_19907);
or UO_596 (O_596,N_19967,N_19964);
and UO_597 (O_597,N_19900,N_19879);
nor UO_598 (O_598,N_19900,N_19929);
or UO_599 (O_599,N_19955,N_19963);
nand UO_600 (O_600,N_19949,N_19829);
or UO_601 (O_601,N_19898,N_19961);
nand UO_602 (O_602,N_19825,N_19879);
and UO_603 (O_603,N_19956,N_19937);
nand UO_604 (O_604,N_19935,N_19838);
and UO_605 (O_605,N_19833,N_19802);
nand UO_606 (O_606,N_19974,N_19982);
or UO_607 (O_607,N_19881,N_19839);
nor UO_608 (O_608,N_19948,N_19835);
and UO_609 (O_609,N_19910,N_19998);
and UO_610 (O_610,N_19977,N_19944);
or UO_611 (O_611,N_19943,N_19946);
nor UO_612 (O_612,N_19834,N_19870);
nand UO_613 (O_613,N_19975,N_19998);
nand UO_614 (O_614,N_19938,N_19899);
nor UO_615 (O_615,N_19921,N_19862);
nor UO_616 (O_616,N_19870,N_19917);
nor UO_617 (O_617,N_19910,N_19977);
or UO_618 (O_618,N_19889,N_19882);
nand UO_619 (O_619,N_19959,N_19920);
nand UO_620 (O_620,N_19907,N_19923);
nand UO_621 (O_621,N_19891,N_19860);
or UO_622 (O_622,N_19884,N_19983);
nor UO_623 (O_623,N_19824,N_19973);
nand UO_624 (O_624,N_19851,N_19995);
nand UO_625 (O_625,N_19800,N_19853);
and UO_626 (O_626,N_19893,N_19852);
or UO_627 (O_627,N_19918,N_19895);
nor UO_628 (O_628,N_19970,N_19930);
or UO_629 (O_629,N_19910,N_19964);
nand UO_630 (O_630,N_19877,N_19824);
and UO_631 (O_631,N_19995,N_19930);
or UO_632 (O_632,N_19811,N_19827);
nor UO_633 (O_633,N_19818,N_19987);
and UO_634 (O_634,N_19818,N_19927);
nand UO_635 (O_635,N_19889,N_19804);
nor UO_636 (O_636,N_19928,N_19830);
nand UO_637 (O_637,N_19832,N_19882);
nand UO_638 (O_638,N_19946,N_19857);
nor UO_639 (O_639,N_19848,N_19815);
and UO_640 (O_640,N_19892,N_19857);
and UO_641 (O_641,N_19859,N_19837);
or UO_642 (O_642,N_19857,N_19818);
and UO_643 (O_643,N_19909,N_19908);
or UO_644 (O_644,N_19856,N_19802);
nor UO_645 (O_645,N_19919,N_19970);
nor UO_646 (O_646,N_19815,N_19987);
xor UO_647 (O_647,N_19967,N_19951);
and UO_648 (O_648,N_19815,N_19804);
and UO_649 (O_649,N_19938,N_19808);
and UO_650 (O_650,N_19938,N_19933);
xor UO_651 (O_651,N_19866,N_19902);
nor UO_652 (O_652,N_19954,N_19943);
nor UO_653 (O_653,N_19980,N_19967);
nor UO_654 (O_654,N_19828,N_19961);
nand UO_655 (O_655,N_19820,N_19895);
nor UO_656 (O_656,N_19910,N_19881);
nand UO_657 (O_657,N_19994,N_19802);
nand UO_658 (O_658,N_19912,N_19932);
or UO_659 (O_659,N_19862,N_19998);
or UO_660 (O_660,N_19864,N_19902);
nor UO_661 (O_661,N_19991,N_19862);
and UO_662 (O_662,N_19834,N_19838);
nor UO_663 (O_663,N_19899,N_19800);
or UO_664 (O_664,N_19988,N_19881);
nor UO_665 (O_665,N_19988,N_19961);
nand UO_666 (O_666,N_19801,N_19822);
nor UO_667 (O_667,N_19936,N_19855);
nor UO_668 (O_668,N_19905,N_19804);
xor UO_669 (O_669,N_19910,N_19898);
or UO_670 (O_670,N_19853,N_19953);
and UO_671 (O_671,N_19902,N_19878);
nor UO_672 (O_672,N_19857,N_19989);
nor UO_673 (O_673,N_19850,N_19962);
nand UO_674 (O_674,N_19877,N_19961);
xor UO_675 (O_675,N_19859,N_19901);
or UO_676 (O_676,N_19847,N_19890);
and UO_677 (O_677,N_19909,N_19857);
or UO_678 (O_678,N_19848,N_19857);
or UO_679 (O_679,N_19991,N_19870);
and UO_680 (O_680,N_19990,N_19979);
or UO_681 (O_681,N_19944,N_19967);
nand UO_682 (O_682,N_19925,N_19847);
nand UO_683 (O_683,N_19840,N_19938);
nand UO_684 (O_684,N_19999,N_19803);
nor UO_685 (O_685,N_19937,N_19872);
nand UO_686 (O_686,N_19923,N_19991);
nor UO_687 (O_687,N_19931,N_19906);
or UO_688 (O_688,N_19933,N_19912);
and UO_689 (O_689,N_19879,N_19911);
nand UO_690 (O_690,N_19909,N_19984);
xnor UO_691 (O_691,N_19977,N_19935);
or UO_692 (O_692,N_19869,N_19982);
or UO_693 (O_693,N_19889,N_19894);
and UO_694 (O_694,N_19990,N_19874);
nand UO_695 (O_695,N_19927,N_19896);
nor UO_696 (O_696,N_19904,N_19878);
nor UO_697 (O_697,N_19911,N_19986);
and UO_698 (O_698,N_19999,N_19824);
nor UO_699 (O_699,N_19904,N_19830);
or UO_700 (O_700,N_19855,N_19988);
nor UO_701 (O_701,N_19808,N_19888);
or UO_702 (O_702,N_19965,N_19841);
nand UO_703 (O_703,N_19810,N_19874);
and UO_704 (O_704,N_19907,N_19906);
and UO_705 (O_705,N_19915,N_19816);
nand UO_706 (O_706,N_19976,N_19833);
nor UO_707 (O_707,N_19934,N_19880);
or UO_708 (O_708,N_19842,N_19906);
nor UO_709 (O_709,N_19841,N_19867);
nand UO_710 (O_710,N_19905,N_19830);
and UO_711 (O_711,N_19876,N_19829);
nand UO_712 (O_712,N_19911,N_19971);
xnor UO_713 (O_713,N_19846,N_19895);
nand UO_714 (O_714,N_19820,N_19918);
nand UO_715 (O_715,N_19944,N_19813);
nand UO_716 (O_716,N_19924,N_19970);
and UO_717 (O_717,N_19809,N_19819);
or UO_718 (O_718,N_19962,N_19926);
or UO_719 (O_719,N_19830,N_19944);
nor UO_720 (O_720,N_19941,N_19928);
nand UO_721 (O_721,N_19862,N_19870);
nand UO_722 (O_722,N_19852,N_19872);
nor UO_723 (O_723,N_19981,N_19806);
or UO_724 (O_724,N_19810,N_19929);
nand UO_725 (O_725,N_19817,N_19988);
and UO_726 (O_726,N_19881,N_19949);
nor UO_727 (O_727,N_19987,N_19802);
nor UO_728 (O_728,N_19865,N_19913);
and UO_729 (O_729,N_19980,N_19826);
nand UO_730 (O_730,N_19822,N_19828);
nor UO_731 (O_731,N_19849,N_19872);
nand UO_732 (O_732,N_19842,N_19850);
and UO_733 (O_733,N_19849,N_19828);
or UO_734 (O_734,N_19832,N_19814);
and UO_735 (O_735,N_19879,N_19962);
nor UO_736 (O_736,N_19860,N_19989);
and UO_737 (O_737,N_19815,N_19986);
nor UO_738 (O_738,N_19949,N_19841);
nor UO_739 (O_739,N_19857,N_19918);
or UO_740 (O_740,N_19905,N_19946);
and UO_741 (O_741,N_19944,N_19822);
nor UO_742 (O_742,N_19904,N_19831);
nand UO_743 (O_743,N_19821,N_19916);
nand UO_744 (O_744,N_19851,N_19999);
or UO_745 (O_745,N_19935,N_19847);
nand UO_746 (O_746,N_19848,N_19992);
nor UO_747 (O_747,N_19813,N_19841);
and UO_748 (O_748,N_19965,N_19955);
or UO_749 (O_749,N_19992,N_19939);
nand UO_750 (O_750,N_19999,N_19939);
nor UO_751 (O_751,N_19999,N_19855);
nand UO_752 (O_752,N_19811,N_19984);
or UO_753 (O_753,N_19864,N_19949);
nand UO_754 (O_754,N_19972,N_19882);
nand UO_755 (O_755,N_19920,N_19984);
or UO_756 (O_756,N_19983,N_19903);
nand UO_757 (O_757,N_19839,N_19918);
and UO_758 (O_758,N_19926,N_19816);
and UO_759 (O_759,N_19957,N_19960);
or UO_760 (O_760,N_19914,N_19829);
nor UO_761 (O_761,N_19815,N_19866);
and UO_762 (O_762,N_19985,N_19915);
nor UO_763 (O_763,N_19986,N_19957);
and UO_764 (O_764,N_19949,N_19966);
or UO_765 (O_765,N_19872,N_19824);
or UO_766 (O_766,N_19921,N_19930);
nor UO_767 (O_767,N_19828,N_19971);
or UO_768 (O_768,N_19810,N_19947);
or UO_769 (O_769,N_19995,N_19826);
nor UO_770 (O_770,N_19870,N_19954);
nand UO_771 (O_771,N_19977,N_19876);
and UO_772 (O_772,N_19916,N_19935);
or UO_773 (O_773,N_19828,N_19943);
or UO_774 (O_774,N_19823,N_19960);
nor UO_775 (O_775,N_19801,N_19824);
nor UO_776 (O_776,N_19859,N_19909);
nor UO_777 (O_777,N_19948,N_19930);
nor UO_778 (O_778,N_19883,N_19984);
and UO_779 (O_779,N_19837,N_19863);
nor UO_780 (O_780,N_19916,N_19999);
nor UO_781 (O_781,N_19922,N_19836);
nand UO_782 (O_782,N_19979,N_19974);
and UO_783 (O_783,N_19906,N_19802);
nor UO_784 (O_784,N_19934,N_19887);
nor UO_785 (O_785,N_19961,N_19992);
nor UO_786 (O_786,N_19989,N_19843);
nor UO_787 (O_787,N_19957,N_19985);
nand UO_788 (O_788,N_19939,N_19878);
and UO_789 (O_789,N_19936,N_19832);
and UO_790 (O_790,N_19807,N_19952);
and UO_791 (O_791,N_19961,N_19991);
nand UO_792 (O_792,N_19827,N_19923);
nor UO_793 (O_793,N_19953,N_19970);
or UO_794 (O_794,N_19801,N_19955);
or UO_795 (O_795,N_19935,N_19839);
or UO_796 (O_796,N_19911,N_19806);
nor UO_797 (O_797,N_19853,N_19920);
and UO_798 (O_798,N_19837,N_19883);
and UO_799 (O_799,N_19965,N_19807);
or UO_800 (O_800,N_19855,N_19984);
and UO_801 (O_801,N_19816,N_19886);
or UO_802 (O_802,N_19970,N_19888);
or UO_803 (O_803,N_19932,N_19981);
nor UO_804 (O_804,N_19885,N_19957);
or UO_805 (O_805,N_19891,N_19998);
nand UO_806 (O_806,N_19841,N_19820);
and UO_807 (O_807,N_19991,N_19946);
nand UO_808 (O_808,N_19838,N_19836);
or UO_809 (O_809,N_19887,N_19967);
and UO_810 (O_810,N_19807,N_19941);
nand UO_811 (O_811,N_19898,N_19834);
and UO_812 (O_812,N_19800,N_19807);
or UO_813 (O_813,N_19936,N_19960);
and UO_814 (O_814,N_19905,N_19991);
nand UO_815 (O_815,N_19909,N_19923);
nor UO_816 (O_816,N_19989,N_19953);
and UO_817 (O_817,N_19993,N_19960);
nand UO_818 (O_818,N_19939,N_19957);
and UO_819 (O_819,N_19881,N_19947);
nand UO_820 (O_820,N_19959,N_19893);
or UO_821 (O_821,N_19883,N_19934);
and UO_822 (O_822,N_19964,N_19979);
or UO_823 (O_823,N_19811,N_19853);
nor UO_824 (O_824,N_19853,N_19823);
nand UO_825 (O_825,N_19993,N_19920);
or UO_826 (O_826,N_19929,N_19845);
and UO_827 (O_827,N_19842,N_19875);
nand UO_828 (O_828,N_19838,N_19960);
nor UO_829 (O_829,N_19988,N_19903);
xnor UO_830 (O_830,N_19994,N_19859);
and UO_831 (O_831,N_19875,N_19986);
nand UO_832 (O_832,N_19923,N_19945);
or UO_833 (O_833,N_19835,N_19875);
and UO_834 (O_834,N_19875,N_19947);
or UO_835 (O_835,N_19943,N_19942);
nand UO_836 (O_836,N_19973,N_19981);
nor UO_837 (O_837,N_19871,N_19824);
or UO_838 (O_838,N_19956,N_19926);
nand UO_839 (O_839,N_19802,N_19857);
nor UO_840 (O_840,N_19940,N_19924);
nor UO_841 (O_841,N_19992,N_19880);
and UO_842 (O_842,N_19858,N_19925);
or UO_843 (O_843,N_19869,N_19883);
nor UO_844 (O_844,N_19877,N_19848);
or UO_845 (O_845,N_19851,N_19833);
nand UO_846 (O_846,N_19954,N_19851);
nand UO_847 (O_847,N_19894,N_19952);
nor UO_848 (O_848,N_19869,N_19933);
nand UO_849 (O_849,N_19960,N_19912);
and UO_850 (O_850,N_19858,N_19984);
or UO_851 (O_851,N_19829,N_19975);
or UO_852 (O_852,N_19812,N_19942);
nor UO_853 (O_853,N_19988,N_19927);
or UO_854 (O_854,N_19897,N_19960);
nor UO_855 (O_855,N_19976,N_19844);
or UO_856 (O_856,N_19815,N_19813);
nand UO_857 (O_857,N_19933,N_19924);
nand UO_858 (O_858,N_19801,N_19810);
nor UO_859 (O_859,N_19848,N_19957);
or UO_860 (O_860,N_19849,N_19844);
xnor UO_861 (O_861,N_19901,N_19875);
nor UO_862 (O_862,N_19947,N_19883);
nor UO_863 (O_863,N_19912,N_19809);
and UO_864 (O_864,N_19806,N_19805);
or UO_865 (O_865,N_19850,N_19913);
nor UO_866 (O_866,N_19976,N_19869);
nand UO_867 (O_867,N_19854,N_19904);
nor UO_868 (O_868,N_19949,N_19811);
or UO_869 (O_869,N_19952,N_19905);
and UO_870 (O_870,N_19939,N_19871);
and UO_871 (O_871,N_19983,N_19927);
nand UO_872 (O_872,N_19968,N_19803);
nand UO_873 (O_873,N_19847,N_19952);
and UO_874 (O_874,N_19841,N_19854);
nand UO_875 (O_875,N_19993,N_19816);
and UO_876 (O_876,N_19834,N_19848);
or UO_877 (O_877,N_19809,N_19981);
nor UO_878 (O_878,N_19934,N_19858);
or UO_879 (O_879,N_19817,N_19982);
nor UO_880 (O_880,N_19843,N_19983);
and UO_881 (O_881,N_19899,N_19913);
nand UO_882 (O_882,N_19937,N_19905);
or UO_883 (O_883,N_19988,N_19841);
nand UO_884 (O_884,N_19887,N_19929);
or UO_885 (O_885,N_19896,N_19956);
or UO_886 (O_886,N_19989,N_19924);
nand UO_887 (O_887,N_19843,N_19821);
nand UO_888 (O_888,N_19934,N_19942);
and UO_889 (O_889,N_19815,N_19850);
and UO_890 (O_890,N_19947,N_19957);
or UO_891 (O_891,N_19891,N_19859);
nor UO_892 (O_892,N_19815,N_19803);
or UO_893 (O_893,N_19858,N_19824);
or UO_894 (O_894,N_19924,N_19957);
or UO_895 (O_895,N_19863,N_19844);
nor UO_896 (O_896,N_19858,N_19844);
or UO_897 (O_897,N_19928,N_19959);
and UO_898 (O_898,N_19904,N_19844);
nor UO_899 (O_899,N_19839,N_19913);
or UO_900 (O_900,N_19885,N_19973);
nand UO_901 (O_901,N_19871,N_19901);
nor UO_902 (O_902,N_19898,N_19901);
or UO_903 (O_903,N_19941,N_19811);
nand UO_904 (O_904,N_19847,N_19931);
nand UO_905 (O_905,N_19944,N_19942);
nor UO_906 (O_906,N_19957,N_19896);
and UO_907 (O_907,N_19992,N_19959);
nand UO_908 (O_908,N_19858,N_19979);
nor UO_909 (O_909,N_19895,N_19950);
nand UO_910 (O_910,N_19954,N_19988);
nor UO_911 (O_911,N_19853,N_19981);
nor UO_912 (O_912,N_19801,N_19923);
nand UO_913 (O_913,N_19920,N_19918);
nor UO_914 (O_914,N_19977,N_19943);
or UO_915 (O_915,N_19952,N_19904);
nand UO_916 (O_916,N_19908,N_19851);
and UO_917 (O_917,N_19929,N_19977);
and UO_918 (O_918,N_19855,N_19915);
nand UO_919 (O_919,N_19972,N_19943);
nor UO_920 (O_920,N_19950,N_19852);
nor UO_921 (O_921,N_19935,N_19813);
nand UO_922 (O_922,N_19870,N_19933);
nand UO_923 (O_923,N_19875,N_19958);
and UO_924 (O_924,N_19848,N_19854);
nand UO_925 (O_925,N_19965,N_19892);
nor UO_926 (O_926,N_19812,N_19809);
nand UO_927 (O_927,N_19993,N_19974);
or UO_928 (O_928,N_19976,N_19845);
and UO_929 (O_929,N_19965,N_19872);
nor UO_930 (O_930,N_19860,N_19934);
nand UO_931 (O_931,N_19895,N_19999);
nand UO_932 (O_932,N_19957,N_19932);
or UO_933 (O_933,N_19911,N_19958);
nand UO_934 (O_934,N_19892,N_19956);
nand UO_935 (O_935,N_19837,N_19999);
and UO_936 (O_936,N_19815,N_19921);
and UO_937 (O_937,N_19885,N_19811);
and UO_938 (O_938,N_19893,N_19817);
or UO_939 (O_939,N_19963,N_19897);
and UO_940 (O_940,N_19874,N_19865);
nor UO_941 (O_941,N_19814,N_19817);
and UO_942 (O_942,N_19919,N_19867);
nor UO_943 (O_943,N_19832,N_19934);
nand UO_944 (O_944,N_19826,N_19857);
or UO_945 (O_945,N_19935,N_19825);
and UO_946 (O_946,N_19843,N_19903);
nor UO_947 (O_947,N_19895,N_19881);
nand UO_948 (O_948,N_19869,N_19809);
nor UO_949 (O_949,N_19893,N_19997);
nor UO_950 (O_950,N_19943,N_19831);
nand UO_951 (O_951,N_19923,N_19985);
or UO_952 (O_952,N_19910,N_19996);
nand UO_953 (O_953,N_19883,N_19907);
nor UO_954 (O_954,N_19943,N_19823);
nand UO_955 (O_955,N_19939,N_19929);
nand UO_956 (O_956,N_19895,N_19801);
nand UO_957 (O_957,N_19906,N_19832);
or UO_958 (O_958,N_19918,N_19821);
nand UO_959 (O_959,N_19923,N_19927);
and UO_960 (O_960,N_19815,N_19925);
and UO_961 (O_961,N_19864,N_19988);
xnor UO_962 (O_962,N_19891,N_19832);
nor UO_963 (O_963,N_19989,N_19848);
nand UO_964 (O_964,N_19822,N_19903);
and UO_965 (O_965,N_19846,N_19832);
or UO_966 (O_966,N_19902,N_19823);
and UO_967 (O_967,N_19925,N_19972);
nand UO_968 (O_968,N_19832,N_19989);
or UO_969 (O_969,N_19927,N_19920);
or UO_970 (O_970,N_19895,N_19969);
and UO_971 (O_971,N_19864,N_19928);
nand UO_972 (O_972,N_19830,N_19819);
nor UO_973 (O_973,N_19815,N_19849);
nor UO_974 (O_974,N_19854,N_19837);
nand UO_975 (O_975,N_19803,N_19812);
nand UO_976 (O_976,N_19896,N_19934);
nor UO_977 (O_977,N_19904,N_19978);
nand UO_978 (O_978,N_19938,N_19855);
nor UO_979 (O_979,N_19940,N_19913);
nor UO_980 (O_980,N_19941,N_19885);
nor UO_981 (O_981,N_19886,N_19903);
and UO_982 (O_982,N_19823,N_19999);
or UO_983 (O_983,N_19878,N_19848);
or UO_984 (O_984,N_19917,N_19871);
or UO_985 (O_985,N_19809,N_19991);
nand UO_986 (O_986,N_19902,N_19840);
nor UO_987 (O_987,N_19863,N_19961);
or UO_988 (O_988,N_19907,N_19887);
and UO_989 (O_989,N_19891,N_19871);
and UO_990 (O_990,N_19900,N_19835);
nand UO_991 (O_991,N_19987,N_19998);
nand UO_992 (O_992,N_19934,N_19959);
xnor UO_993 (O_993,N_19936,N_19954);
nor UO_994 (O_994,N_19942,N_19908);
or UO_995 (O_995,N_19815,N_19805);
and UO_996 (O_996,N_19966,N_19944);
nor UO_997 (O_997,N_19950,N_19910);
or UO_998 (O_998,N_19929,N_19842);
nand UO_999 (O_999,N_19871,N_19861);
and UO_1000 (O_1000,N_19943,N_19810);
and UO_1001 (O_1001,N_19881,N_19999);
or UO_1002 (O_1002,N_19831,N_19819);
nor UO_1003 (O_1003,N_19813,N_19891);
nand UO_1004 (O_1004,N_19916,N_19862);
nand UO_1005 (O_1005,N_19910,N_19848);
or UO_1006 (O_1006,N_19836,N_19814);
or UO_1007 (O_1007,N_19837,N_19938);
nor UO_1008 (O_1008,N_19801,N_19957);
and UO_1009 (O_1009,N_19939,N_19838);
and UO_1010 (O_1010,N_19957,N_19899);
or UO_1011 (O_1011,N_19830,N_19846);
and UO_1012 (O_1012,N_19874,N_19858);
and UO_1013 (O_1013,N_19822,N_19902);
and UO_1014 (O_1014,N_19921,N_19852);
nor UO_1015 (O_1015,N_19807,N_19978);
or UO_1016 (O_1016,N_19933,N_19843);
nor UO_1017 (O_1017,N_19985,N_19812);
and UO_1018 (O_1018,N_19913,N_19977);
nor UO_1019 (O_1019,N_19826,N_19848);
or UO_1020 (O_1020,N_19957,N_19891);
or UO_1021 (O_1021,N_19939,N_19854);
nand UO_1022 (O_1022,N_19869,N_19963);
nor UO_1023 (O_1023,N_19962,N_19997);
nand UO_1024 (O_1024,N_19815,N_19835);
or UO_1025 (O_1025,N_19836,N_19865);
or UO_1026 (O_1026,N_19964,N_19883);
and UO_1027 (O_1027,N_19831,N_19836);
and UO_1028 (O_1028,N_19807,N_19918);
nor UO_1029 (O_1029,N_19842,N_19976);
nand UO_1030 (O_1030,N_19823,N_19922);
nor UO_1031 (O_1031,N_19930,N_19958);
and UO_1032 (O_1032,N_19876,N_19848);
or UO_1033 (O_1033,N_19887,N_19848);
and UO_1034 (O_1034,N_19990,N_19839);
or UO_1035 (O_1035,N_19833,N_19937);
and UO_1036 (O_1036,N_19804,N_19890);
or UO_1037 (O_1037,N_19899,N_19812);
nor UO_1038 (O_1038,N_19920,N_19943);
nor UO_1039 (O_1039,N_19902,N_19800);
nand UO_1040 (O_1040,N_19851,N_19885);
and UO_1041 (O_1041,N_19959,N_19860);
or UO_1042 (O_1042,N_19884,N_19906);
or UO_1043 (O_1043,N_19805,N_19892);
nand UO_1044 (O_1044,N_19880,N_19843);
nor UO_1045 (O_1045,N_19866,N_19930);
and UO_1046 (O_1046,N_19835,N_19996);
nand UO_1047 (O_1047,N_19978,N_19969);
or UO_1048 (O_1048,N_19949,N_19973);
or UO_1049 (O_1049,N_19998,N_19865);
and UO_1050 (O_1050,N_19949,N_19900);
nor UO_1051 (O_1051,N_19871,N_19965);
and UO_1052 (O_1052,N_19837,N_19898);
or UO_1053 (O_1053,N_19976,N_19898);
nand UO_1054 (O_1054,N_19819,N_19883);
nor UO_1055 (O_1055,N_19942,N_19866);
and UO_1056 (O_1056,N_19956,N_19984);
and UO_1057 (O_1057,N_19910,N_19988);
nor UO_1058 (O_1058,N_19873,N_19841);
nand UO_1059 (O_1059,N_19996,N_19988);
or UO_1060 (O_1060,N_19836,N_19941);
and UO_1061 (O_1061,N_19842,N_19823);
nand UO_1062 (O_1062,N_19922,N_19982);
nand UO_1063 (O_1063,N_19965,N_19883);
or UO_1064 (O_1064,N_19867,N_19878);
nor UO_1065 (O_1065,N_19931,N_19971);
or UO_1066 (O_1066,N_19906,N_19848);
nor UO_1067 (O_1067,N_19989,N_19898);
and UO_1068 (O_1068,N_19877,N_19873);
and UO_1069 (O_1069,N_19853,N_19990);
or UO_1070 (O_1070,N_19874,N_19945);
or UO_1071 (O_1071,N_19965,N_19925);
nor UO_1072 (O_1072,N_19820,N_19839);
and UO_1073 (O_1073,N_19847,N_19816);
or UO_1074 (O_1074,N_19991,N_19899);
nor UO_1075 (O_1075,N_19895,N_19935);
or UO_1076 (O_1076,N_19994,N_19896);
nand UO_1077 (O_1077,N_19908,N_19985);
xor UO_1078 (O_1078,N_19989,N_19804);
nand UO_1079 (O_1079,N_19801,N_19873);
or UO_1080 (O_1080,N_19811,N_19872);
or UO_1081 (O_1081,N_19949,N_19936);
nand UO_1082 (O_1082,N_19842,N_19923);
or UO_1083 (O_1083,N_19953,N_19959);
nor UO_1084 (O_1084,N_19889,N_19908);
and UO_1085 (O_1085,N_19875,N_19910);
nor UO_1086 (O_1086,N_19930,N_19838);
nand UO_1087 (O_1087,N_19832,N_19861);
or UO_1088 (O_1088,N_19835,N_19953);
or UO_1089 (O_1089,N_19853,N_19896);
and UO_1090 (O_1090,N_19841,N_19804);
nand UO_1091 (O_1091,N_19889,N_19955);
nand UO_1092 (O_1092,N_19996,N_19926);
and UO_1093 (O_1093,N_19835,N_19934);
or UO_1094 (O_1094,N_19805,N_19944);
or UO_1095 (O_1095,N_19859,N_19865);
nand UO_1096 (O_1096,N_19889,N_19849);
or UO_1097 (O_1097,N_19840,N_19807);
or UO_1098 (O_1098,N_19893,N_19924);
nor UO_1099 (O_1099,N_19915,N_19842);
or UO_1100 (O_1100,N_19891,N_19999);
or UO_1101 (O_1101,N_19865,N_19992);
nor UO_1102 (O_1102,N_19822,N_19931);
or UO_1103 (O_1103,N_19921,N_19844);
and UO_1104 (O_1104,N_19805,N_19850);
or UO_1105 (O_1105,N_19997,N_19815);
nor UO_1106 (O_1106,N_19930,N_19876);
or UO_1107 (O_1107,N_19917,N_19866);
nand UO_1108 (O_1108,N_19855,N_19942);
nor UO_1109 (O_1109,N_19868,N_19898);
nor UO_1110 (O_1110,N_19926,N_19814);
nor UO_1111 (O_1111,N_19910,N_19920);
or UO_1112 (O_1112,N_19960,N_19953);
or UO_1113 (O_1113,N_19964,N_19902);
nand UO_1114 (O_1114,N_19925,N_19981);
and UO_1115 (O_1115,N_19802,N_19824);
nor UO_1116 (O_1116,N_19929,N_19959);
or UO_1117 (O_1117,N_19998,N_19866);
and UO_1118 (O_1118,N_19985,N_19996);
nor UO_1119 (O_1119,N_19834,N_19865);
nand UO_1120 (O_1120,N_19940,N_19920);
nand UO_1121 (O_1121,N_19997,N_19842);
nor UO_1122 (O_1122,N_19904,N_19872);
or UO_1123 (O_1123,N_19916,N_19996);
nor UO_1124 (O_1124,N_19946,N_19995);
nand UO_1125 (O_1125,N_19985,N_19831);
or UO_1126 (O_1126,N_19976,N_19946);
nand UO_1127 (O_1127,N_19899,N_19929);
or UO_1128 (O_1128,N_19866,N_19919);
and UO_1129 (O_1129,N_19963,N_19959);
or UO_1130 (O_1130,N_19911,N_19842);
nor UO_1131 (O_1131,N_19992,N_19893);
nor UO_1132 (O_1132,N_19924,N_19819);
nand UO_1133 (O_1133,N_19807,N_19817);
nor UO_1134 (O_1134,N_19829,N_19960);
nor UO_1135 (O_1135,N_19991,N_19939);
nand UO_1136 (O_1136,N_19898,N_19931);
and UO_1137 (O_1137,N_19872,N_19845);
or UO_1138 (O_1138,N_19987,N_19888);
and UO_1139 (O_1139,N_19888,N_19805);
or UO_1140 (O_1140,N_19818,N_19992);
nor UO_1141 (O_1141,N_19987,N_19977);
or UO_1142 (O_1142,N_19996,N_19978);
and UO_1143 (O_1143,N_19923,N_19816);
nand UO_1144 (O_1144,N_19875,N_19866);
nor UO_1145 (O_1145,N_19940,N_19804);
nor UO_1146 (O_1146,N_19930,N_19826);
nor UO_1147 (O_1147,N_19934,N_19951);
nor UO_1148 (O_1148,N_19992,N_19966);
or UO_1149 (O_1149,N_19802,N_19800);
or UO_1150 (O_1150,N_19916,N_19958);
and UO_1151 (O_1151,N_19905,N_19993);
or UO_1152 (O_1152,N_19960,N_19854);
nor UO_1153 (O_1153,N_19938,N_19902);
and UO_1154 (O_1154,N_19978,N_19956);
nand UO_1155 (O_1155,N_19810,N_19808);
and UO_1156 (O_1156,N_19979,N_19834);
and UO_1157 (O_1157,N_19857,N_19862);
nor UO_1158 (O_1158,N_19976,N_19882);
or UO_1159 (O_1159,N_19906,N_19959);
and UO_1160 (O_1160,N_19853,N_19837);
nand UO_1161 (O_1161,N_19968,N_19973);
or UO_1162 (O_1162,N_19939,N_19975);
and UO_1163 (O_1163,N_19874,N_19918);
and UO_1164 (O_1164,N_19987,N_19841);
or UO_1165 (O_1165,N_19917,N_19933);
and UO_1166 (O_1166,N_19987,N_19811);
or UO_1167 (O_1167,N_19943,N_19908);
and UO_1168 (O_1168,N_19829,N_19920);
or UO_1169 (O_1169,N_19956,N_19945);
nand UO_1170 (O_1170,N_19890,N_19906);
or UO_1171 (O_1171,N_19996,N_19813);
nor UO_1172 (O_1172,N_19868,N_19984);
or UO_1173 (O_1173,N_19996,N_19984);
or UO_1174 (O_1174,N_19863,N_19809);
xnor UO_1175 (O_1175,N_19996,N_19856);
nor UO_1176 (O_1176,N_19878,N_19911);
or UO_1177 (O_1177,N_19996,N_19998);
nand UO_1178 (O_1178,N_19917,N_19930);
nor UO_1179 (O_1179,N_19876,N_19853);
nor UO_1180 (O_1180,N_19819,N_19987);
nand UO_1181 (O_1181,N_19868,N_19840);
nand UO_1182 (O_1182,N_19829,N_19954);
nor UO_1183 (O_1183,N_19984,N_19834);
and UO_1184 (O_1184,N_19978,N_19842);
nand UO_1185 (O_1185,N_19840,N_19800);
nand UO_1186 (O_1186,N_19953,N_19904);
nand UO_1187 (O_1187,N_19862,N_19894);
nor UO_1188 (O_1188,N_19826,N_19838);
and UO_1189 (O_1189,N_19978,N_19869);
nor UO_1190 (O_1190,N_19863,N_19988);
nand UO_1191 (O_1191,N_19847,N_19809);
nand UO_1192 (O_1192,N_19920,N_19949);
nor UO_1193 (O_1193,N_19806,N_19849);
nand UO_1194 (O_1194,N_19836,N_19848);
or UO_1195 (O_1195,N_19987,N_19919);
nor UO_1196 (O_1196,N_19816,N_19873);
or UO_1197 (O_1197,N_19838,N_19800);
or UO_1198 (O_1198,N_19896,N_19971);
nand UO_1199 (O_1199,N_19906,N_19881);
nand UO_1200 (O_1200,N_19806,N_19907);
or UO_1201 (O_1201,N_19954,N_19972);
and UO_1202 (O_1202,N_19856,N_19990);
nand UO_1203 (O_1203,N_19983,N_19982);
nor UO_1204 (O_1204,N_19877,N_19927);
nand UO_1205 (O_1205,N_19943,N_19803);
nor UO_1206 (O_1206,N_19995,N_19924);
nor UO_1207 (O_1207,N_19888,N_19819);
nand UO_1208 (O_1208,N_19814,N_19862);
or UO_1209 (O_1209,N_19946,N_19993);
or UO_1210 (O_1210,N_19805,N_19916);
and UO_1211 (O_1211,N_19951,N_19827);
and UO_1212 (O_1212,N_19975,N_19887);
and UO_1213 (O_1213,N_19966,N_19890);
and UO_1214 (O_1214,N_19804,N_19824);
nand UO_1215 (O_1215,N_19806,N_19926);
and UO_1216 (O_1216,N_19940,N_19864);
and UO_1217 (O_1217,N_19926,N_19899);
and UO_1218 (O_1218,N_19973,N_19945);
and UO_1219 (O_1219,N_19874,N_19930);
nor UO_1220 (O_1220,N_19936,N_19953);
nand UO_1221 (O_1221,N_19980,N_19944);
nand UO_1222 (O_1222,N_19911,N_19967);
or UO_1223 (O_1223,N_19846,N_19946);
or UO_1224 (O_1224,N_19894,N_19800);
nor UO_1225 (O_1225,N_19869,N_19956);
and UO_1226 (O_1226,N_19925,N_19978);
nand UO_1227 (O_1227,N_19936,N_19917);
and UO_1228 (O_1228,N_19982,N_19876);
and UO_1229 (O_1229,N_19964,N_19897);
nor UO_1230 (O_1230,N_19840,N_19806);
xor UO_1231 (O_1231,N_19940,N_19966);
nand UO_1232 (O_1232,N_19984,N_19927);
and UO_1233 (O_1233,N_19908,N_19927);
or UO_1234 (O_1234,N_19911,N_19929);
and UO_1235 (O_1235,N_19941,N_19981);
and UO_1236 (O_1236,N_19924,N_19817);
nor UO_1237 (O_1237,N_19980,N_19981);
or UO_1238 (O_1238,N_19956,N_19825);
or UO_1239 (O_1239,N_19854,N_19901);
nand UO_1240 (O_1240,N_19829,N_19880);
and UO_1241 (O_1241,N_19800,N_19949);
nor UO_1242 (O_1242,N_19907,N_19827);
nor UO_1243 (O_1243,N_19835,N_19851);
and UO_1244 (O_1244,N_19835,N_19805);
nand UO_1245 (O_1245,N_19841,N_19827);
and UO_1246 (O_1246,N_19846,N_19914);
nor UO_1247 (O_1247,N_19919,N_19923);
and UO_1248 (O_1248,N_19889,N_19880);
nor UO_1249 (O_1249,N_19905,N_19872);
or UO_1250 (O_1250,N_19959,N_19917);
or UO_1251 (O_1251,N_19911,N_19866);
nand UO_1252 (O_1252,N_19978,N_19859);
nand UO_1253 (O_1253,N_19847,N_19998);
nor UO_1254 (O_1254,N_19947,N_19902);
nand UO_1255 (O_1255,N_19976,N_19885);
and UO_1256 (O_1256,N_19833,N_19881);
nor UO_1257 (O_1257,N_19890,N_19989);
nor UO_1258 (O_1258,N_19898,N_19975);
nand UO_1259 (O_1259,N_19810,N_19901);
nor UO_1260 (O_1260,N_19809,N_19873);
or UO_1261 (O_1261,N_19915,N_19939);
or UO_1262 (O_1262,N_19829,N_19912);
or UO_1263 (O_1263,N_19863,N_19877);
nand UO_1264 (O_1264,N_19807,N_19878);
or UO_1265 (O_1265,N_19818,N_19890);
or UO_1266 (O_1266,N_19834,N_19861);
nand UO_1267 (O_1267,N_19866,N_19883);
nand UO_1268 (O_1268,N_19990,N_19816);
nor UO_1269 (O_1269,N_19863,N_19898);
and UO_1270 (O_1270,N_19813,N_19845);
nor UO_1271 (O_1271,N_19931,N_19914);
nor UO_1272 (O_1272,N_19929,N_19844);
or UO_1273 (O_1273,N_19876,N_19965);
and UO_1274 (O_1274,N_19848,N_19901);
or UO_1275 (O_1275,N_19863,N_19811);
or UO_1276 (O_1276,N_19916,N_19951);
and UO_1277 (O_1277,N_19831,N_19910);
nor UO_1278 (O_1278,N_19925,N_19870);
or UO_1279 (O_1279,N_19965,N_19830);
nand UO_1280 (O_1280,N_19886,N_19860);
nand UO_1281 (O_1281,N_19901,N_19974);
nand UO_1282 (O_1282,N_19972,N_19999);
nand UO_1283 (O_1283,N_19945,N_19909);
nand UO_1284 (O_1284,N_19879,N_19849);
nor UO_1285 (O_1285,N_19948,N_19872);
or UO_1286 (O_1286,N_19978,N_19823);
or UO_1287 (O_1287,N_19960,N_19990);
or UO_1288 (O_1288,N_19868,N_19995);
nand UO_1289 (O_1289,N_19837,N_19903);
or UO_1290 (O_1290,N_19965,N_19853);
or UO_1291 (O_1291,N_19873,N_19913);
nand UO_1292 (O_1292,N_19856,N_19961);
nor UO_1293 (O_1293,N_19999,N_19914);
or UO_1294 (O_1294,N_19881,N_19891);
nand UO_1295 (O_1295,N_19883,N_19962);
or UO_1296 (O_1296,N_19936,N_19881);
nor UO_1297 (O_1297,N_19876,N_19993);
or UO_1298 (O_1298,N_19962,N_19964);
nor UO_1299 (O_1299,N_19860,N_19893);
or UO_1300 (O_1300,N_19954,N_19990);
nand UO_1301 (O_1301,N_19864,N_19873);
nor UO_1302 (O_1302,N_19823,N_19917);
or UO_1303 (O_1303,N_19963,N_19891);
or UO_1304 (O_1304,N_19818,N_19918);
or UO_1305 (O_1305,N_19822,N_19824);
or UO_1306 (O_1306,N_19852,N_19827);
nand UO_1307 (O_1307,N_19950,N_19892);
nor UO_1308 (O_1308,N_19808,N_19932);
nor UO_1309 (O_1309,N_19892,N_19804);
nand UO_1310 (O_1310,N_19987,N_19821);
or UO_1311 (O_1311,N_19845,N_19903);
and UO_1312 (O_1312,N_19973,N_19818);
or UO_1313 (O_1313,N_19855,N_19889);
xnor UO_1314 (O_1314,N_19943,N_19986);
nand UO_1315 (O_1315,N_19867,N_19992);
nand UO_1316 (O_1316,N_19906,N_19815);
and UO_1317 (O_1317,N_19962,N_19885);
nand UO_1318 (O_1318,N_19972,N_19878);
and UO_1319 (O_1319,N_19930,N_19971);
nand UO_1320 (O_1320,N_19813,N_19857);
xnor UO_1321 (O_1321,N_19957,N_19887);
and UO_1322 (O_1322,N_19806,N_19991);
nor UO_1323 (O_1323,N_19819,N_19939);
xor UO_1324 (O_1324,N_19926,N_19980);
or UO_1325 (O_1325,N_19952,N_19977);
nand UO_1326 (O_1326,N_19874,N_19961);
or UO_1327 (O_1327,N_19856,N_19876);
nor UO_1328 (O_1328,N_19964,N_19974);
nor UO_1329 (O_1329,N_19919,N_19973);
and UO_1330 (O_1330,N_19813,N_19999);
and UO_1331 (O_1331,N_19829,N_19923);
or UO_1332 (O_1332,N_19952,N_19837);
or UO_1333 (O_1333,N_19941,N_19846);
or UO_1334 (O_1334,N_19800,N_19974);
nand UO_1335 (O_1335,N_19922,N_19913);
and UO_1336 (O_1336,N_19972,N_19902);
or UO_1337 (O_1337,N_19968,N_19933);
nor UO_1338 (O_1338,N_19943,N_19895);
nand UO_1339 (O_1339,N_19839,N_19867);
nand UO_1340 (O_1340,N_19876,N_19914);
or UO_1341 (O_1341,N_19884,N_19996);
and UO_1342 (O_1342,N_19915,N_19898);
nor UO_1343 (O_1343,N_19858,N_19878);
nor UO_1344 (O_1344,N_19961,N_19899);
and UO_1345 (O_1345,N_19824,N_19827);
nor UO_1346 (O_1346,N_19828,N_19820);
and UO_1347 (O_1347,N_19906,N_19859);
or UO_1348 (O_1348,N_19829,N_19959);
nand UO_1349 (O_1349,N_19893,N_19908);
nand UO_1350 (O_1350,N_19915,N_19952);
and UO_1351 (O_1351,N_19994,N_19914);
or UO_1352 (O_1352,N_19995,N_19820);
nand UO_1353 (O_1353,N_19832,N_19968);
and UO_1354 (O_1354,N_19816,N_19980);
or UO_1355 (O_1355,N_19924,N_19984);
or UO_1356 (O_1356,N_19850,N_19802);
and UO_1357 (O_1357,N_19885,N_19891);
nand UO_1358 (O_1358,N_19813,N_19972);
or UO_1359 (O_1359,N_19875,N_19941);
and UO_1360 (O_1360,N_19889,N_19810);
nand UO_1361 (O_1361,N_19943,N_19912);
nand UO_1362 (O_1362,N_19953,N_19875);
and UO_1363 (O_1363,N_19906,N_19882);
and UO_1364 (O_1364,N_19807,N_19994);
or UO_1365 (O_1365,N_19987,N_19850);
nand UO_1366 (O_1366,N_19981,N_19825);
and UO_1367 (O_1367,N_19943,N_19904);
nor UO_1368 (O_1368,N_19879,N_19872);
and UO_1369 (O_1369,N_19819,N_19813);
nor UO_1370 (O_1370,N_19898,N_19840);
and UO_1371 (O_1371,N_19960,N_19951);
and UO_1372 (O_1372,N_19955,N_19872);
or UO_1373 (O_1373,N_19864,N_19983);
nand UO_1374 (O_1374,N_19961,N_19945);
nand UO_1375 (O_1375,N_19900,N_19826);
and UO_1376 (O_1376,N_19975,N_19986);
or UO_1377 (O_1377,N_19898,N_19991);
nor UO_1378 (O_1378,N_19937,N_19928);
nand UO_1379 (O_1379,N_19904,N_19896);
nor UO_1380 (O_1380,N_19960,N_19882);
nor UO_1381 (O_1381,N_19978,N_19976);
and UO_1382 (O_1382,N_19820,N_19826);
and UO_1383 (O_1383,N_19920,N_19938);
nand UO_1384 (O_1384,N_19874,N_19940);
and UO_1385 (O_1385,N_19988,N_19875);
and UO_1386 (O_1386,N_19840,N_19944);
nor UO_1387 (O_1387,N_19910,N_19942);
or UO_1388 (O_1388,N_19807,N_19861);
nor UO_1389 (O_1389,N_19824,N_19820);
xor UO_1390 (O_1390,N_19874,N_19875);
and UO_1391 (O_1391,N_19871,N_19994);
nor UO_1392 (O_1392,N_19868,N_19972);
nand UO_1393 (O_1393,N_19900,N_19917);
nand UO_1394 (O_1394,N_19864,N_19946);
nand UO_1395 (O_1395,N_19958,N_19878);
and UO_1396 (O_1396,N_19838,N_19803);
or UO_1397 (O_1397,N_19802,N_19939);
and UO_1398 (O_1398,N_19833,N_19849);
or UO_1399 (O_1399,N_19823,N_19838);
or UO_1400 (O_1400,N_19927,N_19887);
or UO_1401 (O_1401,N_19864,N_19836);
nor UO_1402 (O_1402,N_19892,N_19812);
nor UO_1403 (O_1403,N_19992,N_19846);
nor UO_1404 (O_1404,N_19978,N_19831);
nand UO_1405 (O_1405,N_19856,N_19977);
or UO_1406 (O_1406,N_19904,N_19987);
nand UO_1407 (O_1407,N_19950,N_19903);
and UO_1408 (O_1408,N_19932,N_19966);
and UO_1409 (O_1409,N_19835,N_19846);
nor UO_1410 (O_1410,N_19880,N_19858);
or UO_1411 (O_1411,N_19880,N_19965);
and UO_1412 (O_1412,N_19831,N_19865);
and UO_1413 (O_1413,N_19834,N_19935);
nor UO_1414 (O_1414,N_19801,N_19893);
nand UO_1415 (O_1415,N_19996,N_19947);
nor UO_1416 (O_1416,N_19902,N_19894);
and UO_1417 (O_1417,N_19887,N_19928);
nand UO_1418 (O_1418,N_19897,N_19883);
and UO_1419 (O_1419,N_19952,N_19978);
and UO_1420 (O_1420,N_19814,N_19835);
nor UO_1421 (O_1421,N_19829,N_19958);
nor UO_1422 (O_1422,N_19817,N_19859);
and UO_1423 (O_1423,N_19863,N_19903);
and UO_1424 (O_1424,N_19956,N_19972);
and UO_1425 (O_1425,N_19981,N_19937);
nor UO_1426 (O_1426,N_19958,N_19880);
and UO_1427 (O_1427,N_19900,N_19943);
and UO_1428 (O_1428,N_19818,N_19938);
nand UO_1429 (O_1429,N_19997,N_19918);
and UO_1430 (O_1430,N_19825,N_19839);
and UO_1431 (O_1431,N_19957,N_19898);
and UO_1432 (O_1432,N_19871,N_19959);
nor UO_1433 (O_1433,N_19927,N_19914);
nand UO_1434 (O_1434,N_19819,N_19928);
and UO_1435 (O_1435,N_19948,N_19916);
nor UO_1436 (O_1436,N_19968,N_19843);
nand UO_1437 (O_1437,N_19850,N_19807);
and UO_1438 (O_1438,N_19801,N_19806);
nor UO_1439 (O_1439,N_19859,N_19933);
nand UO_1440 (O_1440,N_19966,N_19970);
and UO_1441 (O_1441,N_19989,N_19863);
and UO_1442 (O_1442,N_19835,N_19923);
nand UO_1443 (O_1443,N_19876,N_19945);
nor UO_1444 (O_1444,N_19847,N_19943);
or UO_1445 (O_1445,N_19996,N_19807);
and UO_1446 (O_1446,N_19860,N_19900);
and UO_1447 (O_1447,N_19830,N_19964);
nor UO_1448 (O_1448,N_19814,N_19915);
or UO_1449 (O_1449,N_19893,N_19907);
nor UO_1450 (O_1450,N_19976,N_19834);
and UO_1451 (O_1451,N_19849,N_19981);
nor UO_1452 (O_1452,N_19820,N_19904);
nand UO_1453 (O_1453,N_19831,N_19912);
and UO_1454 (O_1454,N_19870,N_19977);
nand UO_1455 (O_1455,N_19887,N_19913);
nand UO_1456 (O_1456,N_19844,N_19875);
nand UO_1457 (O_1457,N_19990,N_19864);
and UO_1458 (O_1458,N_19983,N_19934);
or UO_1459 (O_1459,N_19871,N_19958);
or UO_1460 (O_1460,N_19856,N_19814);
nand UO_1461 (O_1461,N_19838,N_19828);
nor UO_1462 (O_1462,N_19938,N_19958);
nand UO_1463 (O_1463,N_19913,N_19932);
or UO_1464 (O_1464,N_19939,N_19856);
or UO_1465 (O_1465,N_19810,N_19922);
nor UO_1466 (O_1466,N_19972,N_19941);
and UO_1467 (O_1467,N_19858,N_19907);
nor UO_1468 (O_1468,N_19860,N_19896);
nor UO_1469 (O_1469,N_19928,N_19853);
nor UO_1470 (O_1470,N_19853,N_19878);
nand UO_1471 (O_1471,N_19905,N_19850);
xnor UO_1472 (O_1472,N_19931,N_19921);
or UO_1473 (O_1473,N_19872,N_19988);
nand UO_1474 (O_1474,N_19858,N_19974);
nor UO_1475 (O_1475,N_19822,N_19865);
nand UO_1476 (O_1476,N_19920,N_19900);
nor UO_1477 (O_1477,N_19911,N_19922);
nand UO_1478 (O_1478,N_19979,N_19932);
or UO_1479 (O_1479,N_19845,N_19833);
nor UO_1480 (O_1480,N_19810,N_19840);
nand UO_1481 (O_1481,N_19856,N_19930);
or UO_1482 (O_1482,N_19838,N_19848);
and UO_1483 (O_1483,N_19991,N_19874);
or UO_1484 (O_1484,N_19842,N_19891);
nand UO_1485 (O_1485,N_19945,N_19966);
or UO_1486 (O_1486,N_19818,N_19935);
or UO_1487 (O_1487,N_19908,N_19950);
or UO_1488 (O_1488,N_19944,N_19869);
nand UO_1489 (O_1489,N_19909,N_19841);
and UO_1490 (O_1490,N_19934,N_19904);
nor UO_1491 (O_1491,N_19879,N_19932);
or UO_1492 (O_1492,N_19886,N_19806);
and UO_1493 (O_1493,N_19868,N_19926);
and UO_1494 (O_1494,N_19830,N_19998);
nand UO_1495 (O_1495,N_19863,N_19862);
nor UO_1496 (O_1496,N_19836,N_19929);
and UO_1497 (O_1497,N_19846,N_19841);
or UO_1498 (O_1498,N_19947,N_19897);
and UO_1499 (O_1499,N_19949,N_19836);
nand UO_1500 (O_1500,N_19921,N_19833);
and UO_1501 (O_1501,N_19928,N_19929);
and UO_1502 (O_1502,N_19908,N_19919);
nand UO_1503 (O_1503,N_19995,N_19800);
or UO_1504 (O_1504,N_19924,N_19903);
or UO_1505 (O_1505,N_19924,N_19977);
nand UO_1506 (O_1506,N_19921,N_19943);
and UO_1507 (O_1507,N_19970,N_19915);
nand UO_1508 (O_1508,N_19953,N_19938);
and UO_1509 (O_1509,N_19924,N_19922);
nand UO_1510 (O_1510,N_19834,N_19929);
and UO_1511 (O_1511,N_19811,N_19975);
nand UO_1512 (O_1512,N_19839,N_19853);
or UO_1513 (O_1513,N_19802,N_19852);
nor UO_1514 (O_1514,N_19930,N_19800);
nand UO_1515 (O_1515,N_19825,N_19874);
nor UO_1516 (O_1516,N_19855,N_19928);
and UO_1517 (O_1517,N_19881,N_19832);
nand UO_1518 (O_1518,N_19965,N_19809);
nor UO_1519 (O_1519,N_19961,N_19926);
or UO_1520 (O_1520,N_19907,N_19979);
or UO_1521 (O_1521,N_19837,N_19914);
nor UO_1522 (O_1522,N_19881,N_19990);
and UO_1523 (O_1523,N_19982,N_19904);
and UO_1524 (O_1524,N_19963,N_19899);
and UO_1525 (O_1525,N_19877,N_19969);
or UO_1526 (O_1526,N_19911,N_19886);
and UO_1527 (O_1527,N_19911,N_19805);
or UO_1528 (O_1528,N_19932,N_19982);
nor UO_1529 (O_1529,N_19863,N_19979);
and UO_1530 (O_1530,N_19967,N_19924);
nor UO_1531 (O_1531,N_19845,N_19862);
nor UO_1532 (O_1532,N_19880,N_19997);
nand UO_1533 (O_1533,N_19877,N_19800);
nand UO_1534 (O_1534,N_19896,N_19841);
nand UO_1535 (O_1535,N_19997,N_19986);
or UO_1536 (O_1536,N_19831,N_19987);
nand UO_1537 (O_1537,N_19969,N_19966);
or UO_1538 (O_1538,N_19816,N_19906);
and UO_1539 (O_1539,N_19952,N_19829);
or UO_1540 (O_1540,N_19972,N_19840);
nor UO_1541 (O_1541,N_19849,N_19944);
nand UO_1542 (O_1542,N_19938,N_19967);
nand UO_1543 (O_1543,N_19996,N_19938);
and UO_1544 (O_1544,N_19914,N_19851);
or UO_1545 (O_1545,N_19977,N_19938);
nand UO_1546 (O_1546,N_19975,N_19864);
nor UO_1547 (O_1547,N_19972,N_19811);
nor UO_1548 (O_1548,N_19868,N_19881);
nand UO_1549 (O_1549,N_19836,N_19829);
nor UO_1550 (O_1550,N_19955,N_19884);
nand UO_1551 (O_1551,N_19839,N_19815);
nor UO_1552 (O_1552,N_19959,N_19985);
and UO_1553 (O_1553,N_19827,N_19836);
nand UO_1554 (O_1554,N_19936,N_19869);
nor UO_1555 (O_1555,N_19951,N_19966);
and UO_1556 (O_1556,N_19944,N_19853);
or UO_1557 (O_1557,N_19807,N_19848);
and UO_1558 (O_1558,N_19837,N_19814);
and UO_1559 (O_1559,N_19944,N_19823);
and UO_1560 (O_1560,N_19905,N_19943);
or UO_1561 (O_1561,N_19835,N_19817);
or UO_1562 (O_1562,N_19916,N_19881);
and UO_1563 (O_1563,N_19945,N_19898);
nand UO_1564 (O_1564,N_19881,N_19842);
nand UO_1565 (O_1565,N_19813,N_19918);
nor UO_1566 (O_1566,N_19980,N_19988);
nand UO_1567 (O_1567,N_19842,N_19840);
nand UO_1568 (O_1568,N_19853,N_19906);
nor UO_1569 (O_1569,N_19827,N_19835);
nand UO_1570 (O_1570,N_19882,N_19988);
and UO_1571 (O_1571,N_19802,N_19955);
or UO_1572 (O_1572,N_19842,N_19894);
or UO_1573 (O_1573,N_19916,N_19840);
nand UO_1574 (O_1574,N_19969,N_19989);
nand UO_1575 (O_1575,N_19820,N_19960);
nand UO_1576 (O_1576,N_19950,N_19970);
or UO_1577 (O_1577,N_19898,N_19822);
nand UO_1578 (O_1578,N_19981,N_19831);
or UO_1579 (O_1579,N_19956,N_19999);
nand UO_1580 (O_1580,N_19859,N_19884);
nor UO_1581 (O_1581,N_19838,N_19931);
nor UO_1582 (O_1582,N_19851,N_19889);
or UO_1583 (O_1583,N_19996,N_19824);
nor UO_1584 (O_1584,N_19824,N_19934);
and UO_1585 (O_1585,N_19844,N_19967);
nor UO_1586 (O_1586,N_19935,N_19845);
nand UO_1587 (O_1587,N_19931,N_19909);
or UO_1588 (O_1588,N_19915,N_19817);
or UO_1589 (O_1589,N_19925,N_19843);
nand UO_1590 (O_1590,N_19974,N_19965);
or UO_1591 (O_1591,N_19961,N_19972);
or UO_1592 (O_1592,N_19926,N_19878);
nor UO_1593 (O_1593,N_19815,N_19972);
nor UO_1594 (O_1594,N_19991,N_19969);
xor UO_1595 (O_1595,N_19854,N_19840);
and UO_1596 (O_1596,N_19885,N_19922);
nor UO_1597 (O_1597,N_19932,N_19830);
or UO_1598 (O_1598,N_19814,N_19921);
or UO_1599 (O_1599,N_19819,N_19835);
nor UO_1600 (O_1600,N_19833,N_19803);
and UO_1601 (O_1601,N_19957,N_19822);
nand UO_1602 (O_1602,N_19972,N_19981);
and UO_1603 (O_1603,N_19886,N_19983);
nor UO_1604 (O_1604,N_19937,N_19862);
and UO_1605 (O_1605,N_19944,N_19985);
nor UO_1606 (O_1606,N_19822,N_19919);
and UO_1607 (O_1607,N_19993,N_19919);
nor UO_1608 (O_1608,N_19913,N_19944);
nand UO_1609 (O_1609,N_19803,N_19863);
and UO_1610 (O_1610,N_19832,N_19931);
nor UO_1611 (O_1611,N_19805,N_19894);
nand UO_1612 (O_1612,N_19881,N_19996);
nand UO_1613 (O_1613,N_19894,N_19938);
and UO_1614 (O_1614,N_19999,N_19817);
nor UO_1615 (O_1615,N_19932,N_19924);
or UO_1616 (O_1616,N_19855,N_19818);
and UO_1617 (O_1617,N_19906,N_19921);
nand UO_1618 (O_1618,N_19803,N_19892);
or UO_1619 (O_1619,N_19834,N_19897);
nor UO_1620 (O_1620,N_19996,N_19839);
or UO_1621 (O_1621,N_19872,N_19830);
or UO_1622 (O_1622,N_19832,N_19976);
or UO_1623 (O_1623,N_19928,N_19888);
or UO_1624 (O_1624,N_19999,N_19990);
and UO_1625 (O_1625,N_19976,N_19883);
nand UO_1626 (O_1626,N_19912,N_19872);
or UO_1627 (O_1627,N_19981,N_19854);
and UO_1628 (O_1628,N_19814,N_19809);
and UO_1629 (O_1629,N_19994,N_19912);
or UO_1630 (O_1630,N_19898,N_19902);
nand UO_1631 (O_1631,N_19974,N_19826);
or UO_1632 (O_1632,N_19994,N_19824);
or UO_1633 (O_1633,N_19940,N_19872);
or UO_1634 (O_1634,N_19853,N_19901);
or UO_1635 (O_1635,N_19860,N_19931);
nand UO_1636 (O_1636,N_19899,N_19914);
and UO_1637 (O_1637,N_19953,N_19894);
and UO_1638 (O_1638,N_19830,N_19937);
xnor UO_1639 (O_1639,N_19937,N_19940);
nand UO_1640 (O_1640,N_19800,N_19956);
nor UO_1641 (O_1641,N_19948,N_19810);
and UO_1642 (O_1642,N_19970,N_19904);
nor UO_1643 (O_1643,N_19859,N_19979);
nor UO_1644 (O_1644,N_19818,N_19894);
and UO_1645 (O_1645,N_19926,N_19989);
nand UO_1646 (O_1646,N_19932,N_19961);
and UO_1647 (O_1647,N_19866,N_19977);
and UO_1648 (O_1648,N_19846,N_19828);
nand UO_1649 (O_1649,N_19998,N_19922);
nor UO_1650 (O_1650,N_19958,N_19804);
or UO_1651 (O_1651,N_19964,N_19864);
or UO_1652 (O_1652,N_19980,N_19971);
or UO_1653 (O_1653,N_19929,N_19883);
and UO_1654 (O_1654,N_19854,N_19808);
nor UO_1655 (O_1655,N_19965,N_19884);
nor UO_1656 (O_1656,N_19966,N_19828);
and UO_1657 (O_1657,N_19898,N_19861);
and UO_1658 (O_1658,N_19839,N_19991);
nor UO_1659 (O_1659,N_19853,N_19864);
or UO_1660 (O_1660,N_19807,N_19842);
nor UO_1661 (O_1661,N_19800,N_19817);
and UO_1662 (O_1662,N_19874,N_19964);
nand UO_1663 (O_1663,N_19885,N_19870);
or UO_1664 (O_1664,N_19861,N_19940);
or UO_1665 (O_1665,N_19887,N_19815);
nor UO_1666 (O_1666,N_19968,N_19822);
and UO_1667 (O_1667,N_19972,N_19945);
nor UO_1668 (O_1668,N_19854,N_19876);
nor UO_1669 (O_1669,N_19826,N_19976);
nand UO_1670 (O_1670,N_19854,N_19919);
and UO_1671 (O_1671,N_19919,N_19971);
nand UO_1672 (O_1672,N_19882,N_19842);
nor UO_1673 (O_1673,N_19841,N_19874);
nor UO_1674 (O_1674,N_19894,N_19867);
xnor UO_1675 (O_1675,N_19982,N_19892);
nor UO_1676 (O_1676,N_19992,N_19815);
and UO_1677 (O_1677,N_19993,N_19914);
and UO_1678 (O_1678,N_19998,N_19854);
or UO_1679 (O_1679,N_19810,N_19829);
nor UO_1680 (O_1680,N_19887,N_19990);
nand UO_1681 (O_1681,N_19851,N_19867);
and UO_1682 (O_1682,N_19978,N_19931);
and UO_1683 (O_1683,N_19876,N_19960);
or UO_1684 (O_1684,N_19999,N_19863);
nand UO_1685 (O_1685,N_19987,N_19835);
nor UO_1686 (O_1686,N_19837,N_19825);
and UO_1687 (O_1687,N_19974,N_19995);
nand UO_1688 (O_1688,N_19903,N_19939);
and UO_1689 (O_1689,N_19909,N_19969);
nor UO_1690 (O_1690,N_19835,N_19980);
and UO_1691 (O_1691,N_19880,N_19970);
nand UO_1692 (O_1692,N_19848,N_19825);
and UO_1693 (O_1693,N_19967,N_19931);
nor UO_1694 (O_1694,N_19895,N_19852);
nor UO_1695 (O_1695,N_19865,N_19928);
nand UO_1696 (O_1696,N_19821,N_19982);
nor UO_1697 (O_1697,N_19914,N_19938);
nor UO_1698 (O_1698,N_19824,N_19905);
or UO_1699 (O_1699,N_19815,N_19820);
or UO_1700 (O_1700,N_19908,N_19804);
nor UO_1701 (O_1701,N_19904,N_19849);
nand UO_1702 (O_1702,N_19981,N_19951);
or UO_1703 (O_1703,N_19970,N_19913);
nor UO_1704 (O_1704,N_19906,N_19901);
nor UO_1705 (O_1705,N_19969,N_19800);
or UO_1706 (O_1706,N_19854,N_19902);
nor UO_1707 (O_1707,N_19936,N_19866);
xnor UO_1708 (O_1708,N_19979,N_19872);
or UO_1709 (O_1709,N_19935,N_19918);
or UO_1710 (O_1710,N_19927,N_19942);
or UO_1711 (O_1711,N_19905,N_19828);
or UO_1712 (O_1712,N_19818,N_19846);
and UO_1713 (O_1713,N_19990,N_19950);
nand UO_1714 (O_1714,N_19878,N_19914);
nor UO_1715 (O_1715,N_19854,N_19847);
nor UO_1716 (O_1716,N_19848,N_19839);
or UO_1717 (O_1717,N_19973,N_19810);
nor UO_1718 (O_1718,N_19993,N_19990);
nand UO_1719 (O_1719,N_19876,N_19846);
or UO_1720 (O_1720,N_19850,N_19926);
nand UO_1721 (O_1721,N_19914,N_19961);
or UO_1722 (O_1722,N_19973,N_19892);
nand UO_1723 (O_1723,N_19967,N_19854);
or UO_1724 (O_1724,N_19805,N_19970);
and UO_1725 (O_1725,N_19944,N_19836);
nand UO_1726 (O_1726,N_19872,N_19882);
nor UO_1727 (O_1727,N_19913,N_19808);
nor UO_1728 (O_1728,N_19835,N_19821);
nand UO_1729 (O_1729,N_19893,N_19993);
and UO_1730 (O_1730,N_19840,N_19907);
or UO_1731 (O_1731,N_19810,N_19935);
or UO_1732 (O_1732,N_19820,N_19838);
nor UO_1733 (O_1733,N_19961,N_19976);
and UO_1734 (O_1734,N_19999,N_19806);
nand UO_1735 (O_1735,N_19883,N_19804);
or UO_1736 (O_1736,N_19997,N_19907);
or UO_1737 (O_1737,N_19869,N_19952);
and UO_1738 (O_1738,N_19820,N_19927);
nand UO_1739 (O_1739,N_19858,N_19916);
nor UO_1740 (O_1740,N_19962,N_19973);
and UO_1741 (O_1741,N_19959,N_19919);
nor UO_1742 (O_1742,N_19953,N_19857);
nand UO_1743 (O_1743,N_19979,N_19996);
nor UO_1744 (O_1744,N_19902,N_19982);
nor UO_1745 (O_1745,N_19949,N_19957);
and UO_1746 (O_1746,N_19876,N_19998);
nor UO_1747 (O_1747,N_19950,N_19935);
nor UO_1748 (O_1748,N_19848,N_19843);
nor UO_1749 (O_1749,N_19846,N_19886);
or UO_1750 (O_1750,N_19946,N_19964);
and UO_1751 (O_1751,N_19826,N_19965);
nor UO_1752 (O_1752,N_19977,N_19825);
or UO_1753 (O_1753,N_19985,N_19992);
or UO_1754 (O_1754,N_19881,N_19945);
and UO_1755 (O_1755,N_19915,N_19921);
nand UO_1756 (O_1756,N_19913,N_19957);
and UO_1757 (O_1757,N_19873,N_19849);
nor UO_1758 (O_1758,N_19816,N_19881);
nor UO_1759 (O_1759,N_19894,N_19958);
or UO_1760 (O_1760,N_19981,N_19930);
nand UO_1761 (O_1761,N_19928,N_19863);
or UO_1762 (O_1762,N_19967,N_19952);
or UO_1763 (O_1763,N_19835,N_19943);
nand UO_1764 (O_1764,N_19976,N_19875);
and UO_1765 (O_1765,N_19948,N_19925);
or UO_1766 (O_1766,N_19936,N_19822);
xor UO_1767 (O_1767,N_19873,N_19958);
or UO_1768 (O_1768,N_19972,N_19976);
and UO_1769 (O_1769,N_19959,N_19927);
nor UO_1770 (O_1770,N_19990,N_19911);
and UO_1771 (O_1771,N_19860,N_19831);
nor UO_1772 (O_1772,N_19879,N_19943);
nand UO_1773 (O_1773,N_19961,N_19990);
nor UO_1774 (O_1774,N_19873,N_19932);
nor UO_1775 (O_1775,N_19821,N_19990);
nand UO_1776 (O_1776,N_19988,N_19912);
nor UO_1777 (O_1777,N_19954,N_19804);
or UO_1778 (O_1778,N_19895,N_19857);
nand UO_1779 (O_1779,N_19979,N_19829);
and UO_1780 (O_1780,N_19873,N_19928);
xor UO_1781 (O_1781,N_19921,N_19880);
nor UO_1782 (O_1782,N_19862,N_19850);
nand UO_1783 (O_1783,N_19866,N_19821);
nor UO_1784 (O_1784,N_19899,N_19886);
nand UO_1785 (O_1785,N_19887,N_19903);
nor UO_1786 (O_1786,N_19856,N_19869);
nand UO_1787 (O_1787,N_19829,N_19843);
nand UO_1788 (O_1788,N_19940,N_19849);
or UO_1789 (O_1789,N_19892,N_19964);
or UO_1790 (O_1790,N_19878,N_19968);
and UO_1791 (O_1791,N_19865,N_19892);
nand UO_1792 (O_1792,N_19962,N_19866);
nor UO_1793 (O_1793,N_19891,N_19867);
nor UO_1794 (O_1794,N_19982,N_19966);
nor UO_1795 (O_1795,N_19997,N_19904);
nand UO_1796 (O_1796,N_19887,N_19873);
nand UO_1797 (O_1797,N_19926,N_19830);
nand UO_1798 (O_1798,N_19915,N_19924);
or UO_1799 (O_1799,N_19815,N_19955);
and UO_1800 (O_1800,N_19978,N_19867);
nand UO_1801 (O_1801,N_19993,N_19896);
and UO_1802 (O_1802,N_19812,N_19955);
or UO_1803 (O_1803,N_19874,N_19860);
or UO_1804 (O_1804,N_19924,N_19836);
xnor UO_1805 (O_1805,N_19802,N_19827);
and UO_1806 (O_1806,N_19974,N_19911);
nor UO_1807 (O_1807,N_19944,N_19923);
xnor UO_1808 (O_1808,N_19813,N_19914);
nand UO_1809 (O_1809,N_19834,N_19965);
and UO_1810 (O_1810,N_19837,N_19845);
or UO_1811 (O_1811,N_19920,N_19810);
and UO_1812 (O_1812,N_19993,N_19928);
nor UO_1813 (O_1813,N_19878,N_19957);
and UO_1814 (O_1814,N_19806,N_19996);
nand UO_1815 (O_1815,N_19860,N_19921);
nor UO_1816 (O_1816,N_19856,N_19885);
and UO_1817 (O_1817,N_19868,N_19846);
nand UO_1818 (O_1818,N_19906,N_19949);
nand UO_1819 (O_1819,N_19820,N_19871);
and UO_1820 (O_1820,N_19943,N_19839);
or UO_1821 (O_1821,N_19884,N_19887);
or UO_1822 (O_1822,N_19843,N_19808);
and UO_1823 (O_1823,N_19959,N_19823);
and UO_1824 (O_1824,N_19929,N_19942);
nand UO_1825 (O_1825,N_19888,N_19998);
nor UO_1826 (O_1826,N_19956,N_19958);
or UO_1827 (O_1827,N_19989,N_19886);
nor UO_1828 (O_1828,N_19870,N_19953);
nand UO_1829 (O_1829,N_19806,N_19997);
and UO_1830 (O_1830,N_19825,N_19996);
nand UO_1831 (O_1831,N_19939,N_19901);
nor UO_1832 (O_1832,N_19966,N_19881);
and UO_1833 (O_1833,N_19994,N_19872);
nand UO_1834 (O_1834,N_19947,N_19912);
nand UO_1835 (O_1835,N_19966,N_19835);
or UO_1836 (O_1836,N_19956,N_19983);
and UO_1837 (O_1837,N_19812,N_19929);
or UO_1838 (O_1838,N_19823,N_19955);
or UO_1839 (O_1839,N_19938,N_19904);
and UO_1840 (O_1840,N_19814,N_19880);
and UO_1841 (O_1841,N_19956,N_19823);
nand UO_1842 (O_1842,N_19813,N_19934);
nand UO_1843 (O_1843,N_19852,N_19807);
and UO_1844 (O_1844,N_19899,N_19966);
or UO_1845 (O_1845,N_19840,N_19977);
and UO_1846 (O_1846,N_19849,N_19878);
nand UO_1847 (O_1847,N_19869,N_19885);
and UO_1848 (O_1848,N_19989,N_19820);
nor UO_1849 (O_1849,N_19828,N_19937);
and UO_1850 (O_1850,N_19965,N_19862);
or UO_1851 (O_1851,N_19997,N_19908);
or UO_1852 (O_1852,N_19867,N_19906);
or UO_1853 (O_1853,N_19865,N_19850);
or UO_1854 (O_1854,N_19884,N_19935);
and UO_1855 (O_1855,N_19858,N_19997);
and UO_1856 (O_1856,N_19883,N_19933);
or UO_1857 (O_1857,N_19831,N_19901);
nand UO_1858 (O_1858,N_19899,N_19879);
and UO_1859 (O_1859,N_19809,N_19933);
nand UO_1860 (O_1860,N_19936,N_19977);
nor UO_1861 (O_1861,N_19833,N_19858);
nor UO_1862 (O_1862,N_19852,N_19963);
nand UO_1863 (O_1863,N_19947,N_19861);
or UO_1864 (O_1864,N_19879,N_19841);
nor UO_1865 (O_1865,N_19866,N_19901);
nand UO_1866 (O_1866,N_19934,N_19817);
or UO_1867 (O_1867,N_19877,N_19862);
nand UO_1868 (O_1868,N_19922,N_19932);
nand UO_1869 (O_1869,N_19941,N_19964);
or UO_1870 (O_1870,N_19883,N_19973);
nand UO_1871 (O_1871,N_19914,N_19933);
nor UO_1872 (O_1872,N_19860,N_19872);
or UO_1873 (O_1873,N_19913,N_19864);
or UO_1874 (O_1874,N_19945,N_19940);
nand UO_1875 (O_1875,N_19963,N_19901);
or UO_1876 (O_1876,N_19914,N_19877);
or UO_1877 (O_1877,N_19834,N_19981);
and UO_1878 (O_1878,N_19846,N_19851);
or UO_1879 (O_1879,N_19864,N_19962);
or UO_1880 (O_1880,N_19833,N_19927);
and UO_1881 (O_1881,N_19843,N_19952);
or UO_1882 (O_1882,N_19959,N_19848);
and UO_1883 (O_1883,N_19932,N_19862);
or UO_1884 (O_1884,N_19812,N_19842);
nor UO_1885 (O_1885,N_19852,N_19826);
or UO_1886 (O_1886,N_19996,N_19997);
or UO_1887 (O_1887,N_19886,N_19893);
nor UO_1888 (O_1888,N_19971,N_19834);
nand UO_1889 (O_1889,N_19858,N_19996);
or UO_1890 (O_1890,N_19979,N_19953);
nand UO_1891 (O_1891,N_19819,N_19832);
or UO_1892 (O_1892,N_19915,N_19866);
nor UO_1893 (O_1893,N_19885,N_19979);
nand UO_1894 (O_1894,N_19962,N_19808);
nor UO_1895 (O_1895,N_19938,N_19898);
or UO_1896 (O_1896,N_19924,N_19955);
and UO_1897 (O_1897,N_19820,N_19953);
or UO_1898 (O_1898,N_19978,N_19983);
nand UO_1899 (O_1899,N_19849,N_19923);
or UO_1900 (O_1900,N_19999,N_19967);
or UO_1901 (O_1901,N_19822,N_19992);
and UO_1902 (O_1902,N_19992,N_19934);
and UO_1903 (O_1903,N_19857,N_19823);
or UO_1904 (O_1904,N_19959,N_19935);
or UO_1905 (O_1905,N_19894,N_19879);
and UO_1906 (O_1906,N_19916,N_19851);
or UO_1907 (O_1907,N_19994,N_19946);
and UO_1908 (O_1908,N_19955,N_19808);
nand UO_1909 (O_1909,N_19957,N_19900);
or UO_1910 (O_1910,N_19977,N_19850);
and UO_1911 (O_1911,N_19847,N_19845);
or UO_1912 (O_1912,N_19901,N_19814);
and UO_1913 (O_1913,N_19959,N_19842);
or UO_1914 (O_1914,N_19807,N_19984);
nor UO_1915 (O_1915,N_19914,N_19839);
nor UO_1916 (O_1916,N_19903,N_19958);
nand UO_1917 (O_1917,N_19857,N_19851);
and UO_1918 (O_1918,N_19932,N_19813);
nand UO_1919 (O_1919,N_19958,N_19992);
nor UO_1920 (O_1920,N_19915,N_19868);
nor UO_1921 (O_1921,N_19983,N_19811);
nor UO_1922 (O_1922,N_19901,N_19927);
xnor UO_1923 (O_1923,N_19935,N_19836);
and UO_1924 (O_1924,N_19978,N_19928);
nand UO_1925 (O_1925,N_19809,N_19835);
nor UO_1926 (O_1926,N_19958,N_19891);
or UO_1927 (O_1927,N_19972,N_19850);
and UO_1928 (O_1928,N_19849,N_19963);
nor UO_1929 (O_1929,N_19932,N_19882);
or UO_1930 (O_1930,N_19871,N_19947);
and UO_1931 (O_1931,N_19993,N_19825);
nor UO_1932 (O_1932,N_19970,N_19813);
nor UO_1933 (O_1933,N_19849,N_19826);
nor UO_1934 (O_1934,N_19870,N_19941);
nor UO_1935 (O_1935,N_19968,N_19899);
nand UO_1936 (O_1936,N_19947,N_19970);
nor UO_1937 (O_1937,N_19944,N_19927);
and UO_1938 (O_1938,N_19819,N_19852);
or UO_1939 (O_1939,N_19955,N_19865);
or UO_1940 (O_1940,N_19914,N_19855);
and UO_1941 (O_1941,N_19892,N_19811);
nor UO_1942 (O_1942,N_19905,N_19976);
nor UO_1943 (O_1943,N_19952,N_19880);
nand UO_1944 (O_1944,N_19980,N_19878);
or UO_1945 (O_1945,N_19858,N_19940);
nand UO_1946 (O_1946,N_19802,N_19807);
nor UO_1947 (O_1947,N_19856,N_19992);
and UO_1948 (O_1948,N_19874,N_19989);
or UO_1949 (O_1949,N_19835,N_19847);
or UO_1950 (O_1950,N_19860,N_19847);
or UO_1951 (O_1951,N_19878,N_19931);
or UO_1952 (O_1952,N_19952,N_19890);
and UO_1953 (O_1953,N_19934,N_19960);
nor UO_1954 (O_1954,N_19985,N_19868);
nand UO_1955 (O_1955,N_19865,N_19946);
nand UO_1956 (O_1956,N_19814,N_19900);
and UO_1957 (O_1957,N_19883,N_19969);
nor UO_1958 (O_1958,N_19821,N_19945);
or UO_1959 (O_1959,N_19814,N_19953);
nand UO_1960 (O_1960,N_19923,N_19942);
nand UO_1961 (O_1961,N_19895,N_19970);
or UO_1962 (O_1962,N_19984,N_19960);
and UO_1963 (O_1963,N_19946,N_19923);
and UO_1964 (O_1964,N_19877,N_19972);
nor UO_1965 (O_1965,N_19965,N_19835);
or UO_1966 (O_1966,N_19944,N_19872);
or UO_1967 (O_1967,N_19988,N_19975);
nand UO_1968 (O_1968,N_19928,N_19914);
and UO_1969 (O_1969,N_19986,N_19811);
nand UO_1970 (O_1970,N_19944,N_19861);
nor UO_1971 (O_1971,N_19928,N_19817);
nand UO_1972 (O_1972,N_19809,N_19962);
and UO_1973 (O_1973,N_19801,N_19829);
nand UO_1974 (O_1974,N_19802,N_19990);
nand UO_1975 (O_1975,N_19808,N_19965);
nor UO_1976 (O_1976,N_19906,N_19872);
nand UO_1977 (O_1977,N_19844,N_19803);
nor UO_1978 (O_1978,N_19853,N_19923);
and UO_1979 (O_1979,N_19807,N_19883);
and UO_1980 (O_1980,N_19838,N_19845);
nand UO_1981 (O_1981,N_19832,N_19862);
nor UO_1982 (O_1982,N_19811,N_19860);
and UO_1983 (O_1983,N_19869,N_19881);
nor UO_1984 (O_1984,N_19826,N_19899);
and UO_1985 (O_1985,N_19977,N_19940);
and UO_1986 (O_1986,N_19809,N_19840);
or UO_1987 (O_1987,N_19907,N_19890);
nand UO_1988 (O_1988,N_19804,N_19917);
or UO_1989 (O_1989,N_19997,N_19825);
nor UO_1990 (O_1990,N_19818,N_19990);
or UO_1991 (O_1991,N_19946,N_19998);
or UO_1992 (O_1992,N_19888,N_19983);
nor UO_1993 (O_1993,N_19895,N_19893);
nand UO_1994 (O_1994,N_19940,N_19881);
nor UO_1995 (O_1995,N_19914,N_19905);
nand UO_1996 (O_1996,N_19990,N_19897);
nand UO_1997 (O_1997,N_19995,N_19819);
nand UO_1998 (O_1998,N_19971,N_19943);
and UO_1999 (O_1999,N_19828,N_19934);
nand UO_2000 (O_2000,N_19821,N_19889);
or UO_2001 (O_2001,N_19927,N_19844);
nor UO_2002 (O_2002,N_19926,N_19861);
nor UO_2003 (O_2003,N_19826,N_19912);
and UO_2004 (O_2004,N_19910,N_19888);
or UO_2005 (O_2005,N_19991,N_19911);
nor UO_2006 (O_2006,N_19800,N_19833);
and UO_2007 (O_2007,N_19921,N_19884);
and UO_2008 (O_2008,N_19833,N_19808);
xnor UO_2009 (O_2009,N_19915,N_19913);
or UO_2010 (O_2010,N_19858,N_19850);
and UO_2011 (O_2011,N_19934,N_19901);
nand UO_2012 (O_2012,N_19817,N_19952);
and UO_2013 (O_2013,N_19871,N_19908);
and UO_2014 (O_2014,N_19897,N_19835);
nand UO_2015 (O_2015,N_19971,N_19838);
nand UO_2016 (O_2016,N_19960,N_19896);
nand UO_2017 (O_2017,N_19819,N_19895);
or UO_2018 (O_2018,N_19942,N_19964);
nor UO_2019 (O_2019,N_19988,N_19822);
and UO_2020 (O_2020,N_19918,N_19926);
or UO_2021 (O_2021,N_19973,N_19929);
or UO_2022 (O_2022,N_19892,N_19927);
nand UO_2023 (O_2023,N_19877,N_19977);
nor UO_2024 (O_2024,N_19847,N_19934);
or UO_2025 (O_2025,N_19936,N_19910);
nor UO_2026 (O_2026,N_19994,N_19901);
nand UO_2027 (O_2027,N_19866,N_19865);
nor UO_2028 (O_2028,N_19826,N_19984);
nor UO_2029 (O_2029,N_19854,N_19806);
and UO_2030 (O_2030,N_19888,N_19964);
or UO_2031 (O_2031,N_19989,N_19970);
nor UO_2032 (O_2032,N_19804,N_19949);
and UO_2033 (O_2033,N_19987,N_19980);
or UO_2034 (O_2034,N_19998,N_19962);
or UO_2035 (O_2035,N_19942,N_19800);
nand UO_2036 (O_2036,N_19933,N_19983);
and UO_2037 (O_2037,N_19941,N_19878);
nand UO_2038 (O_2038,N_19978,N_19919);
or UO_2039 (O_2039,N_19950,N_19996);
or UO_2040 (O_2040,N_19886,N_19969);
nor UO_2041 (O_2041,N_19867,N_19922);
or UO_2042 (O_2042,N_19939,N_19825);
or UO_2043 (O_2043,N_19930,N_19916);
or UO_2044 (O_2044,N_19909,N_19940);
nor UO_2045 (O_2045,N_19903,N_19902);
nor UO_2046 (O_2046,N_19964,N_19873);
nor UO_2047 (O_2047,N_19845,N_19815);
and UO_2048 (O_2048,N_19833,N_19804);
and UO_2049 (O_2049,N_19997,N_19836);
or UO_2050 (O_2050,N_19935,N_19899);
nor UO_2051 (O_2051,N_19871,N_19950);
and UO_2052 (O_2052,N_19854,N_19852);
and UO_2053 (O_2053,N_19804,N_19838);
or UO_2054 (O_2054,N_19973,N_19909);
nand UO_2055 (O_2055,N_19845,N_19800);
or UO_2056 (O_2056,N_19911,N_19992);
nand UO_2057 (O_2057,N_19808,N_19845);
nor UO_2058 (O_2058,N_19879,N_19985);
nor UO_2059 (O_2059,N_19927,N_19996);
and UO_2060 (O_2060,N_19844,N_19997);
nand UO_2061 (O_2061,N_19946,N_19810);
nor UO_2062 (O_2062,N_19836,N_19908);
and UO_2063 (O_2063,N_19867,N_19981);
and UO_2064 (O_2064,N_19904,N_19907);
nand UO_2065 (O_2065,N_19970,N_19949);
xnor UO_2066 (O_2066,N_19966,N_19834);
nand UO_2067 (O_2067,N_19866,N_19951);
nand UO_2068 (O_2068,N_19803,N_19835);
nor UO_2069 (O_2069,N_19878,N_19961);
or UO_2070 (O_2070,N_19845,N_19877);
or UO_2071 (O_2071,N_19925,N_19833);
nor UO_2072 (O_2072,N_19814,N_19824);
nor UO_2073 (O_2073,N_19920,N_19815);
nor UO_2074 (O_2074,N_19860,N_19904);
or UO_2075 (O_2075,N_19806,N_19994);
and UO_2076 (O_2076,N_19878,N_19955);
and UO_2077 (O_2077,N_19923,N_19802);
and UO_2078 (O_2078,N_19909,N_19829);
or UO_2079 (O_2079,N_19912,N_19844);
nor UO_2080 (O_2080,N_19843,N_19909);
and UO_2081 (O_2081,N_19811,N_19920);
nand UO_2082 (O_2082,N_19873,N_19905);
and UO_2083 (O_2083,N_19888,N_19853);
nor UO_2084 (O_2084,N_19994,N_19899);
and UO_2085 (O_2085,N_19905,N_19822);
nor UO_2086 (O_2086,N_19852,N_19804);
and UO_2087 (O_2087,N_19846,N_19960);
and UO_2088 (O_2088,N_19872,N_19984);
nand UO_2089 (O_2089,N_19805,N_19967);
xor UO_2090 (O_2090,N_19940,N_19813);
or UO_2091 (O_2091,N_19893,N_19842);
or UO_2092 (O_2092,N_19825,N_19897);
nor UO_2093 (O_2093,N_19957,N_19999);
nor UO_2094 (O_2094,N_19835,N_19838);
nand UO_2095 (O_2095,N_19994,N_19945);
xnor UO_2096 (O_2096,N_19919,N_19975);
and UO_2097 (O_2097,N_19814,N_19940);
nand UO_2098 (O_2098,N_19955,N_19849);
and UO_2099 (O_2099,N_19958,N_19943);
nor UO_2100 (O_2100,N_19967,N_19995);
and UO_2101 (O_2101,N_19960,N_19892);
and UO_2102 (O_2102,N_19968,N_19823);
or UO_2103 (O_2103,N_19908,N_19863);
and UO_2104 (O_2104,N_19821,N_19930);
nand UO_2105 (O_2105,N_19865,N_19887);
or UO_2106 (O_2106,N_19951,N_19878);
nor UO_2107 (O_2107,N_19966,N_19913);
or UO_2108 (O_2108,N_19936,N_19853);
nand UO_2109 (O_2109,N_19956,N_19873);
or UO_2110 (O_2110,N_19966,N_19888);
nand UO_2111 (O_2111,N_19885,N_19966);
and UO_2112 (O_2112,N_19922,N_19993);
nand UO_2113 (O_2113,N_19855,N_19885);
and UO_2114 (O_2114,N_19935,N_19975);
xor UO_2115 (O_2115,N_19987,N_19935);
nand UO_2116 (O_2116,N_19953,N_19840);
nor UO_2117 (O_2117,N_19829,N_19936);
or UO_2118 (O_2118,N_19804,N_19995);
nand UO_2119 (O_2119,N_19915,N_19865);
nand UO_2120 (O_2120,N_19969,N_19887);
xnor UO_2121 (O_2121,N_19869,N_19998);
nand UO_2122 (O_2122,N_19809,N_19961);
nand UO_2123 (O_2123,N_19804,N_19945);
and UO_2124 (O_2124,N_19879,N_19858);
or UO_2125 (O_2125,N_19943,N_19856);
or UO_2126 (O_2126,N_19837,N_19870);
nor UO_2127 (O_2127,N_19815,N_19806);
and UO_2128 (O_2128,N_19951,N_19828);
nor UO_2129 (O_2129,N_19933,N_19906);
nor UO_2130 (O_2130,N_19945,N_19962);
nand UO_2131 (O_2131,N_19822,N_19831);
or UO_2132 (O_2132,N_19805,N_19988);
nor UO_2133 (O_2133,N_19898,N_19815);
or UO_2134 (O_2134,N_19954,N_19836);
nor UO_2135 (O_2135,N_19802,N_19907);
nand UO_2136 (O_2136,N_19894,N_19849);
nor UO_2137 (O_2137,N_19982,N_19925);
and UO_2138 (O_2138,N_19801,N_19990);
or UO_2139 (O_2139,N_19803,N_19908);
nor UO_2140 (O_2140,N_19866,N_19829);
nor UO_2141 (O_2141,N_19818,N_19811);
nor UO_2142 (O_2142,N_19907,N_19833);
and UO_2143 (O_2143,N_19892,N_19945);
nor UO_2144 (O_2144,N_19948,N_19991);
xnor UO_2145 (O_2145,N_19942,N_19826);
or UO_2146 (O_2146,N_19841,N_19995);
nor UO_2147 (O_2147,N_19921,N_19933);
and UO_2148 (O_2148,N_19856,N_19839);
nor UO_2149 (O_2149,N_19846,N_19867);
and UO_2150 (O_2150,N_19842,N_19912);
nor UO_2151 (O_2151,N_19995,N_19805);
nor UO_2152 (O_2152,N_19953,N_19852);
nor UO_2153 (O_2153,N_19893,N_19904);
nand UO_2154 (O_2154,N_19895,N_19983);
and UO_2155 (O_2155,N_19807,N_19803);
or UO_2156 (O_2156,N_19974,N_19948);
and UO_2157 (O_2157,N_19964,N_19924);
or UO_2158 (O_2158,N_19891,N_19983);
or UO_2159 (O_2159,N_19948,N_19985);
and UO_2160 (O_2160,N_19867,N_19838);
nor UO_2161 (O_2161,N_19898,N_19882);
and UO_2162 (O_2162,N_19843,N_19914);
nand UO_2163 (O_2163,N_19883,N_19853);
nor UO_2164 (O_2164,N_19858,N_19849);
nand UO_2165 (O_2165,N_19848,N_19986);
nand UO_2166 (O_2166,N_19899,N_19964);
nand UO_2167 (O_2167,N_19806,N_19953);
nand UO_2168 (O_2168,N_19961,N_19813);
nand UO_2169 (O_2169,N_19841,N_19918);
nand UO_2170 (O_2170,N_19919,N_19865);
and UO_2171 (O_2171,N_19846,N_19879);
and UO_2172 (O_2172,N_19820,N_19887);
nor UO_2173 (O_2173,N_19992,N_19953);
or UO_2174 (O_2174,N_19998,N_19877);
nor UO_2175 (O_2175,N_19959,N_19956);
nand UO_2176 (O_2176,N_19892,N_19872);
or UO_2177 (O_2177,N_19863,N_19909);
or UO_2178 (O_2178,N_19808,N_19876);
nand UO_2179 (O_2179,N_19883,N_19948);
nor UO_2180 (O_2180,N_19931,N_19804);
nor UO_2181 (O_2181,N_19986,N_19858);
nor UO_2182 (O_2182,N_19848,N_19861);
nand UO_2183 (O_2183,N_19925,N_19911);
nor UO_2184 (O_2184,N_19906,N_19808);
nand UO_2185 (O_2185,N_19858,N_19828);
or UO_2186 (O_2186,N_19904,N_19822);
or UO_2187 (O_2187,N_19967,N_19977);
or UO_2188 (O_2188,N_19850,N_19970);
and UO_2189 (O_2189,N_19933,N_19996);
and UO_2190 (O_2190,N_19992,N_19987);
and UO_2191 (O_2191,N_19920,N_19862);
and UO_2192 (O_2192,N_19882,N_19934);
nor UO_2193 (O_2193,N_19870,N_19970);
and UO_2194 (O_2194,N_19813,N_19856);
nor UO_2195 (O_2195,N_19955,N_19856);
and UO_2196 (O_2196,N_19954,N_19994);
nand UO_2197 (O_2197,N_19985,N_19823);
nor UO_2198 (O_2198,N_19953,N_19886);
and UO_2199 (O_2199,N_19836,N_19876);
or UO_2200 (O_2200,N_19975,N_19913);
or UO_2201 (O_2201,N_19800,N_19832);
or UO_2202 (O_2202,N_19875,N_19895);
or UO_2203 (O_2203,N_19922,N_19819);
or UO_2204 (O_2204,N_19850,N_19952);
nor UO_2205 (O_2205,N_19831,N_19971);
or UO_2206 (O_2206,N_19849,N_19961);
or UO_2207 (O_2207,N_19970,N_19976);
nor UO_2208 (O_2208,N_19842,N_19988);
and UO_2209 (O_2209,N_19852,N_19941);
nand UO_2210 (O_2210,N_19960,N_19870);
or UO_2211 (O_2211,N_19946,N_19999);
and UO_2212 (O_2212,N_19968,N_19862);
nand UO_2213 (O_2213,N_19989,N_19821);
or UO_2214 (O_2214,N_19993,N_19852);
and UO_2215 (O_2215,N_19949,N_19990);
and UO_2216 (O_2216,N_19989,N_19995);
or UO_2217 (O_2217,N_19898,N_19813);
nor UO_2218 (O_2218,N_19870,N_19899);
and UO_2219 (O_2219,N_19829,N_19937);
nor UO_2220 (O_2220,N_19979,N_19884);
or UO_2221 (O_2221,N_19971,N_19809);
and UO_2222 (O_2222,N_19859,N_19832);
or UO_2223 (O_2223,N_19838,N_19877);
nor UO_2224 (O_2224,N_19825,N_19823);
nand UO_2225 (O_2225,N_19946,N_19808);
or UO_2226 (O_2226,N_19879,N_19928);
or UO_2227 (O_2227,N_19991,N_19802);
nor UO_2228 (O_2228,N_19990,N_19973);
and UO_2229 (O_2229,N_19827,N_19865);
nor UO_2230 (O_2230,N_19853,N_19964);
or UO_2231 (O_2231,N_19855,N_19897);
nor UO_2232 (O_2232,N_19906,N_19891);
and UO_2233 (O_2233,N_19832,N_19955);
or UO_2234 (O_2234,N_19917,N_19852);
nand UO_2235 (O_2235,N_19910,N_19891);
and UO_2236 (O_2236,N_19804,N_19823);
nand UO_2237 (O_2237,N_19944,N_19910);
nor UO_2238 (O_2238,N_19862,N_19898);
and UO_2239 (O_2239,N_19800,N_19978);
nor UO_2240 (O_2240,N_19839,N_19826);
or UO_2241 (O_2241,N_19838,N_19878);
and UO_2242 (O_2242,N_19894,N_19839);
or UO_2243 (O_2243,N_19843,N_19907);
and UO_2244 (O_2244,N_19973,N_19847);
nand UO_2245 (O_2245,N_19971,N_19848);
nor UO_2246 (O_2246,N_19821,N_19871);
or UO_2247 (O_2247,N_19899,N_19992);
nor UO_2248 (O_2248,N_19925,N_19996);
or UO_2249 (O_2249,N_19954,N_19921);
and UO_2250 (O_2250,N_19965,N_19992);
or UO_2251 (O_2251,N_19937,N_19834);
nor UO_2252 (O_2252,N_19800,N_19980);
xor UO_2253 (O_2253,N_19971,N_19859);
and UO_2254 (O_2254,N_19961,N_19951);
or UO_2255 (O_2255,N_19935,N_19869);
nand UO_2256 (O_2256,N_19915,N_19979);
nand UO_2257 (O_2257,N_19965,N_19922);
nand UO_2258 (O_2258,N_19870,N_19883);
and UO_2259 (O_2259,N_19972,N_19885);
and UO_2260 (O_2260,N_19895,N_19848);
or UO_2261 (O_2261,N_19806,N_19850);
and UO_2262 (O_2262,N_19828,N_19917);
nor UO_2263 (O_2263,N_19927,N_19891);
nor UO_2264 (O_2264,N_19988,N_19867);
and UO_2265 (O_2265,N_19985,N_19833);
nor UO_2266 (O_2266,N_19873,N_19975);
nor UO_2267 (O_2267,N_19901,N_19896);
nor UO_2268 (O_2268,N_19859,N_19905);
nand UO_2269 (O_2269,N_19957,N_19830);
and UO_2270 (O_2270,N_19919,N_19861);
nor UO_2271 (O_2271,N_19870,N_19892);
or UO_2272 (O_2272,N_19903,N_19989);
nor UO_2273 (O_2273,N_19863,N_19893);
or UO_2274 (O_2274,N_19874,N_19950);
and UO_2275 (O_2275,N_19938,N_19979);
nand UO_2276 (O_2276,N_19825,N_19878);
nand UO_2277 (O_2277,N_19887,N_19819);
nand UO_2278 (O_2278,N_19854,N_19997);
nand UO_2279 (O_2279,N_19982,N_19815);
and UO_2280 (O_2280,N_19906,N_19849);
nand UO_2281 (O_2281,N_19953,N_19947);
nor UO_2282 (O_2282,N_19866,N_19820);
or UO_2283 (O_2283,N_19944,N_19809);
nor UO_2284 (O_2284,N_19845,N_19996);
nor UO_2285 (O_2285,N_19835,N_19845);
or UO_2286 (O_2286,N_19858,N_19825);
nand UO_2287 (O_2287,N_19952,N_19853);
nor UO_2288 (O_2288,N_19809,N_19811);
nor UO_2289 (O_2289,N_19850,N_19879);
and UO_2290 (O_2290,N_19864,N_19969);
or UO_2291 (O_2291,N_19841,N_19935);
nor UO_2292 (O_2292,N_19955,N_19998);
nand UO_2293 (O_2293,N_19849,N_19948);
nand UO_2294 (O_2294,N_19838,N_19898);
or UO_2295 (O_2295,N_19931,N_19805);
or UO_2296 (O_2296,N_19844,N_19992);
nor UO_2297 (O_2297,N_19886,N_19971);
nand UO_2298 (O_2298,N_19978,N_19841);
nand UO_2299 (O_2299,N_19881,N_19944);
or UO_2300 (O_2300,N_19853,N_19855);
and UO_2301 (O_2301,N_19896,N_19886);
nand UO_2302 (O_2302,N_19978,N_19824);
or UO_2303 (O_2303,N_19940,N_19893);
and UO_2304 (O_2304,N_19807,N_19985);
nand UO_2305 (O_2305,N_19994,N_19962);
nor UO_2306 (O_2306,N_19854,N_19875);
and UO_2307 (O_2307,N_19893,N_19830);
nand UO_2308 (O_2308,N_19962,N_19891);
nor UO_2309 (O_2309,N_19976,N_19963);
and UO_2310 (O_2310,N_19965,N_19852);
nor UO_2311 (O_2311,N_19883,N_19894);
and UO_2312 (O_2312,N_19984,N_19972);
and UO_2313 (O_2313,N_19843,N_19919);
nand UO_2314 (O_2314,N_19972,N_19847);
nand UO_2315 (O_2315,N_19892,N_19871);
and UO_2316 (O_2316,N_19963,N_19854);
and UO_2317 (O_2317,N_19876,N_19992);
nand UO_2318 (O_2318,N_19867,N_19946);
xor UO_2319 (O_2319,N_19906,N_19999);
or UO_2320 (O_2320,N_19935,N_19968);
nand UO_2321 (O_2321,N_19977,N_19965);
nor UO_2322 (O_2322,N_19847,N_19856);
nand UO_2323 (O_2323,N_19929,N_19998);
or UO_2324 (O_2324,N_19854,N_19929);
or UO_2325 (O_2325,N_19817,N_19957);
or UO_2326 (O_2326,N_19926,N_19858);
or UO_2327 (O_2327,N_19865,N_19812);
nor UO_2328 (O_2328,N_19939,N_19803);
nand UO_2329 (O_2329,N_19925,N_19819);
and UO_2330 (O_2330,N_19954,N_19899);
or UO_2331 (O_2331,N_19920,N_19884);
or UO_2332 (O_2332,N_19914,N_19937);
and UO_2333 (O_2333,N_19921,N_19898);
or UO_2334 (O_2334,N_19841,N_19985);
nor UO_2335 (O_2335,N_19996,N_19857);
nand UO_2336 (O_2336,N_19825,N_19832);
or UO_2337 (O_2337,N_19853,N_19974);
and UO_2338 (O_2338,N_19813,N_19971);
nor UO_2339 (O_2339,N_19970,N_19922);
nand UO_2340 (O_2340,N_19912,N_19837);
or UO_2341 (O_2341,N_19928,N_19991);
nor UO_2342 (O_2342,N_19888,N_19934);
or UO_2343 (O_2343,N_19896,N_19828);
and UO_2344 (O_2344,N_19936,N_19961);
nand UO_2345 (O_2345,N_19969,N_19902);
or UO_2346 (O_2346,N_19948,N_19829);
and UO_2347 (O_2347,N_19813,N_19920);
nand UO_2348 (O_2348,N_19880,N_19982);
or UO_2349 (O_2349,N_19955,N_19830);
nand UO_2350 (O_2350,N_19810,N_19892);
or UO_2351 (O_2351,N_19918,N_19847);
and UO_2352 (O_2352,N_19808,N_19903);
nor UO_2353 (O_2353,N_19806,N_19965);
nand UO_2354 (O_2354,N_19921,N_19941);
and UO_2355 (O_2355,N_19856,N_19919);
or UO_2356 (O_2356,N_19960,N_19916);
nor UO_2357 (O_2357,N_19869,N_19997);
or UO_2358 (O_2358,N_19814,N_19954);
nor UO_2359 (O_2359,N_19810,N_19893);
nor UO_2360 (O_2360,N_19972,N_19816);
nor UO_2361 (O_2361,N_19830,N_19809);
and UO_2362 (O_2362,N_19969,N_19981);
nor UO_2363 (O_2363,N_19936,N_19994);
and UO_2364 (O_2364,N_19817,N_19869);
nand UO_2365 (O_2365,N_19996,N_19802);
nor UO_2366 (O_2366,N_19934,N_19994);
or UO_2367 (O_2367,N_19947,N_19820);
and UO_2368 (O_2368,N_19935,N_19907);
nor UO_2369 (O_2369,N_19880,N_19847);
and UO_2370 (O_2370,N_19971,N_19862);
nor UO_2371 (O_2371,N_19822,N_19971);
nor UO_2372 (O_2372,N_19893,N_19968);
nand UO_2373 (O_2373,N_19954,N_19840);
nand UO_2374 (O_2374,N_19820,N_19873);
nand UO_2375 (O_2375,N_19903,N_19934);
nor UO_2376 (O_2376,N_19813,N_19929);
and UO_2377 (O_2377,N_19849,N_19839);
xor UO_2378 (O_2378,N_19879,N_19864);
and UO_2379 (O_2379,N_19853,N_19870);
nand UO_2380 (O_2380,N_19931,N_19966);
nand UO_2381 (O_2381,N_19834,N_19877);
nand UO_2382 (O_2382,N_19833,N_19842);
nand UO_2383 (O_2383,N_19823,N_19970);
nand UO_2384 (O_2384,N_19805,N_19969);
xnor UO_2385 (O_2385,N_19988,N_19835);
nand UO_2386 (O_2386,N_19980,N_19807);
nor UO_2387 (O_2387,N_19843,N_19812);
nand UO_2388 (O_2388,N_19890,N_19896);
nand UO_2389 (O_2389,N_19941,N_19966);
and UO_2390 (O_2390,N_19907,N_19810);
nand UO_2391 (O_2391,N_19985,N_19969);
nand UO_2392 (O_2392,N_19809,N_19917);
or UO_2393 (O_2393,N_19888,N_19913);
nor UO_2394 (O_2394,N_19876,N_19800);
or UO_2395 (O_2395,N_19801,N_19945);
nor UO_2396 (O_2396,N_19966,N_19965);
or UO_2397 (O_2397,N_19849,N_19845);
and UO_2398 (O_2398,N_19922,N_19931);
and UO_2399 (O_2399,N_19941,N_19970);
nand UO_2400 (O_2400,N_19979,N_19918);
nor UO_2401 (O_2401,N_19947,N_19967);
nor UO_2402 (O_2402,N_19943,N_19953);
nand UO_2403 (O_2403,N_19844,N_19833);
nor UO_2404 (O_2404,N_19990,N_19995);
nand UO_2405 (O_2405,N_19915,N_19805);
and UO_2406 (O_2406,N_19902,N_19937);
nor UO_2407 (O_2407,N_19954,N_19805);
or UO_2408 (O_2408,N_19804,N_19848);
or UO_2409 (O_2409,N_19835,N_19810);
and UO_2410 (O_2410,N_19801,N_19835);
and UO_2411 (O_2411,N_19976,N_19973);
and UO_2412 (O_2412,N_19987,N_19941);
or UO_2413 (O_2413,N_19841,N_19852);
nand UO_2414 (O_2414,N_19850,N_19979);
nor UO_2415 (O_2415,N_19932,N_19996);
nor UO_2416 (O_2416,N_19833,N_19977);
or UO_2417 (O_2417,N_19869,N_19872);
and UO_2418 (O_2418,N_19991,N_19875);
or UO_2419 (O_2419,N_19827,N_19996);
nand UO_2420 (O_2420,N_19923,N_19979);
or UO_2421 (O_2421,N_19838,N_19926);
or UO_2422 (O_2422,N_19927,N_19905);
and UO_2423 (O_2423,N_19954,N_19934);
nor UO_2424 (O_2424,N_19934,N_19970);
or UO_2425 (O_2425,N_19900,N_19880);
or UO_2426 (O_2426,N_19818,N_19943);
and UO_2427 (O_2427,N_19926,N_19884);
nand UO_2428 (O_2428,N_19863,N_19892);
nor UO_2429 (O_2429,N_19814,N_19963);
and UO_2430 (O_2430,N_19950,N_19993);
or UO_2431 (O_2431,N_19899,N_19863);
nor UO_2432 (O_2432,N_19888,N_19959);
nor UO_2433 (O_2433,N_19874,N_19827);
nor UO_2434 (O_2434,N_19987,N_19863);
nand UO_2435 (O_2435,N_19817,N_19973);
and UO_2436 (O_2436,N_19808,N_19807);
or UO_2437 (O_2437,N_19951,N_19945);
nand UO_2438 (O_2438,N_19905,N_19844);
or UO_2439 (O_2439,N_19849,N_19957);
or UO_2440 (O_2440,N_19857,N_19903);
nand UO_2441 (O_2441,N_19945,N_19954);
or UO_2442 (O_2442,N_19948,N_19964);
or UO_2443 (O_2443,N_19973,N_19899);
or UO_2444 (O_2444,N_19809,N_19898);
and UO_2445 (O_2445,N_19957,N_19973);
or UO_2446 (O_2446,N_19820,N_19971);
nor UO_2447 (O_2447,N_19968,N_19881);
nand UO_2448 (O_2448,N_19889,N_19828);
or UO_2449 (O_2449,N_19922,N_19947);
or UO_2450 (O_2450,N_19831,N_19927);
nand UO_2451 (O_2451,N_19886,N_19955);
or UO_2452 (O_2452,N_19903,N_19872);
and UO_2453 (O_2453,N_19875,N_19968);
and UO_2454 (O_2454,N_19912,N_19919);
nor UO_2455 (O_2455,N_19872,N_19846);
nand UO_2456 (O_2456,N_19887,N_19959);
nor UO_2457 (O_2457,N_19827,N_19985);
nor UO_2458 (O_2458,N_19856,N_19873);
nor UO_2459 (O_2459,N_19893,N_19958);
or UO_2460 (O_2460,N_19974,N_19984);
nand UO_2461 (O_2461,N_19954,N_19817);
nand UO_2462 (O_2462,N_19895,N_19805);
nand UO_2463 (O_2463,N_19935,N_19872);
and UO_2464 (O_2464,N_19993,N_19969);
or UO_2465 (O_2465,N_19899,N_19937);
nor UO_2466 (O_2466,N_19868,N_19906);
nand UO_2467 (O_2467,N_19920,N_19838);
nor UO_2468 (O_2468,N_19990,N_19852);
nor UO_2469 (O_2469,N_19930,N_19861);
xor UO_2470 (O_2470,N_19848,N_19916);
or UO_2471 (O_2471,N_19975,N_19876);
and UO_2472 (O_2472,N_19964,N_19823);
and UO_2473 (O_2473,N_19876,N_19820);
nor UO_2474 (O_2474,N_19995,N_19870);
nand UO_2475 (O_2475,N_19836,N_19962);
or UO_2476 (O_2476,N_19865,N_19974);
and UO_2477 (O_2477,N_19843,N_19980);
nand UO_2478 (O_2478,N_19844,N_19879);
nand UO_2479 (O_2479,N_19960,N_19821);
and UO_2480 (O_2480,N_19934,N_19875);
and UO_2481 (O_2481,N_19972,N_19889);
nor UO_2482 (O_2482,N_19973,N_19808);
or UO_2483 (O_2483,N_19933,N_19986);
nor UO_2484 (O_2484,N_19823,N_19877);
xor UO_2485 (O_2485,N_19991,N_19873);
nand UO_2486 (O_2486,N_19837,N_19813);
nand UO_2487 (O_2487,N_19984,N_19806);
nand UO_2488 (O_2488,N_19897,N_19961);
and UO_2489 (O_2489,N_19910,N_19940);
and UO_2490 (O_2490,N_19969,N_19865);
nand UO_2491 (O_2491,N_19899,N_19996);
xnor UO_2492 (O_2492,N_19873,N_19897);
nor UO_2493 (O_2493,N_19989,N_19838);
nor UO_2494 (O_2494,N_19826,N_19865);
nand UO_2495 (O_2495,N_19924,N_19849);
nand UO_2496 (O_2496,N_19986,N_19969);
nor UO_2497 (O_2497,N_19944,N_19806);
or UO_2498 (O_2498,N_19844,N_19954);
nand UO_2499 (O_2499,N_19801,N_19919);
endmodule