module basic_500_3000_500_6_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_398,In_73);
and U1 (N_1,In_239,In_63);
nor U2 (N_2,In_452,In_438);
xnor U3 (N_3,In_0,In_117);
nor U4 (N_4,In_275,In_406);
and U5 (N_5,In_171,In_399);
and U6 (N_6,In_187,In_363);
nor U7 (N_7,In_11,In_321);
or U8 (N_8,In_329,In_299);
or U9 (N_9,In_195,In_41);
nand U10 (N_10,In_220,In_269);
xnor U11 (N_11,In_394,In_383);
nor U12 (N_12,In_3,In_270);
nor U13 (N_13,In_144,In_379);
nor U14 (N_14,In_172,In_158);
nand U15 (N_15,In_473,In_96);
xor U16 (N_16,In_24,In_232);
and U17 (N_17,In_100,In_78);
xnor U18 (N_18,In_318,In_451);
or U19 (N_19,In_5,In_86);
nand U20 (N_20,In_273,In_164);
and U21 (N_21,In_392,In_221);
nand U22 (N_22,In_39,In_61);
and U23 (N_23,In_437,In_217);
xnor U24 (N_24,In_281,In_170);
nand U25 (N_25,In_129,In_336);
or U26 (N_26,In_479,In_296);
nand U27 (N_27,In_209,In_27);
xor U28 (N_28,In_223,In_368);
xor U29 (N_29,In_391,In_48);
nor U30 (N_30,In_25,In_372);
and U31 (N_31,In_22,In_405);
nor U32 (N_32,In_285,In_136);
xor U33 (N_33,In_457,In_107);
nor U34 (N_34,In_141,In_198);
nand U35 (N_35,In_415,In_19);
xnor U36 (N_36,In_287,In_252);
and U37 (N_37,In_76,In_454);
or U38 (N_38,In_115,In_23);
nand U39 (N_39,In_148,In_421);
nand U40 (N_40,In_265,In_409);
xor U41 (N_41,In_54,In_259);
xnor U42 (N_42,In_359,In_348);
and U43 (N_43,In_43,In_143);
xnor U44 (N_44,In_42,In_53);
or U45 (N_45,In_484,In_190);
nand U46 (N_46,In_343,In_88);
nand U47 (N_47,In_38,In_330);
xor U48 (N_48,In_207,In_465);
and U49 (N_49,In_137,In_213);
nor U50 (N_50,In_295,In_416);
and U51 (N_51,In_153,In_499);
xnor U52 (N_52,In_494,In_2);
nand U53 (N_53,In_331,In_430);
nor U54 (N_54,In_192,In_126);
xor U55 (N_55,In_342,In_133);
xnor U56 (N_56,In_442,In_112);
and U57 (N_57,In_49,In_305);
nand U58 (N_58,In_340,In_151);
and U59 (N_59,In_498,In_445);
or U60 (N_60,In_434,In_361);
or U61 (N_61,In_216,In_109);
xor U62 (N_62,In_357,In_358);
or U63 (N_63,In_8,In_150);
or U64 (N_64,In_453,In_227);
xnor U65 (N_65,In_108,In_243);
and U66 (N_66,In_196,In_201);
xor U67 (N_67,In_279,In_414);
nand U68 (N_68,In_166,In_180);
and U69 (N_69,In_244,In_118);
and U70 (N_70,In_74,In_104);
xor U71 (N_71,In_183,In_135);
or U72 (N_72,In_84,In_116);
nand U73 (N_73,In_215,In_450);
and U74 (N_74,In_225,In_175);
nor U75 (N_75,In_256,In_472);
or U76 (N_76,In_354,In_360);
nand U77 (N_77,In_30,In_300);
xnor U78 (N_78,In_492,In_206);
nor U79 (N_79,In_461,In_355);
and U80 (N_80,In_468,In_91);
and U81 (N_81,In_337,In_441);
or U82 (N_82,In_288,In_167);
or U83 (N_83,In_474,In_333);
nand U84 (N_84,In_145,In_9);
nor U85 (N_85,In_272,In_66);
xor U86 (N_86,In_419,In_245);
nand U87 (N_87,In_423,In_45);
and U88 (N_88,In_15,In_56);
nand U89 (N_89,In_212,In_369);
xor U90 (N_90,In_134,In_464);
and U91 (N_91,In_185,In_306);
and U92 (N_92,In_59,In_81);
or U93 (N_93,In_155,In_458);
nor U94 (N_94,In_93,In_493);
xor U95 (N_95,In_72,In_236);
and U96 (N_96,In_388,In_413);
nor U97 (N_97,In_482,In_335);
or U98 (N_98,In_101,In_427);
nor U99 (N_99,In_334,In_261);
nand U100 (N_100,In_55,In_204);
and U101 (N_101,In_268,In_124);
nor U102 (N_102,In_401,In_477);
or U103 (N_103,In_267,In_352);
nand U104 (N_104,In_467,In_50);
and U105 (N_105,In_407,In_481);
nor U106 (N_106,In_233,In_226);
nor U107 (N_107,In_478,In_142);
or U108 (N_108,In_40,In_283);
and U109 (N_109,In_436,In_266);
and U110 (N_110,In_77,In_312);
nand U111 (N_111,In_254,In_51);
and U112 (N_112,In_353,In_264);
and U113 (N_113,In_229,In_121);
and U114 (N_114,In_176,In_189);
xor U115 (N_115,In_128,In_122);
xnor U116 (N_116,In_263,In_29);
or U117 (N_117,In_292,In_486);
or U118 (N_118,In_160,In_370);
xnor U119 (N_119,In_130,In_242);
nand U120 (N_120,In_488,In_308);
nand U121 (N_121,In_120,In_483);
nor U122 (N_122,In_328,In_444);
nor U123 (N_123,In_293,In_320);
or U124 (N_124,In_18,In_106);
nor U125 (N_125,In_471,In_113);
nand U126 (N_126,In_98,In_378);
xor U127 (N_127,In_79,In_411);
or U128 (N_128,In_33,In_332);
and U129 (N_129,In_289,In_282);
nor U130 (N_130,In_297,In_278);
or U131 (N_131,In_140,In_314);
nand U132 (N_132,In_6,In_10);
xor U133 (N_133,In_230,In_410);
nand U134 (N_134,In_365,In_257);
xnor U135 (N_135,In_367,In_469);
nor U136 (N_136,In_31,In_179);
or U137 (N_137,In_208,In_377);
and U138 (N_138,In_324,In_322);
nor U139 (N_139,In_235,In_75);
or U140 (N_140,In_138,In_271);
xor U141 (N_141,In_13,In_374);
nand U142 (N_142,In_169,In_376);
nand U143 (N_143,In_119,In_114);
nor U144 (N_144,In_149,In_83);
nor U145 (N_145,In_184,In_203);
and U146 (N_146,In_339,In_253);
nand U147 (N_147,In_387,In_491);
or U148 (N_148,In_380,In_237);
nand U149 (N_149,In_487,In_85);
or U150 (N_150,In_17,In_131);
nor U151 (N_151,In_350,In_188);
nor U152 (N_152,In_302,In_90);
nand U153 (N_153,In_455,In_424);
and U154 (N_154,In_47,In_260);
or U155 (N_155,In_303,In_351);
nor U156 (N_156,In_349,In_480);
xor U157 (N_157,In_87,In_404);
or U158 (N_158,In_356,In_341);
and U159 (N_159,In_7,In_470);
or U160 (N_160,In_364,In_165);
or U161 (N_161,In_161,In_127);
or U162 (N_162,In_97,In_286);
and U163 (N_163,In_182,In_110);
or U164 (N_164,In_319,In_92);
and U165 (N_165,In_420,In_60);
xnor U166 (N_166,In_403,In_375);
xor U167 (N_167,In_178,In_386);
or U168 (N_168,In_238,In_428);
nor U169 (N_169,In_224,In_248);
nand U170 (N_170,In_4,In_62);
or U171 (N_171,In_280,In_80);
nand U172 (N_172,In_94,In_396);
xnor U173 (N_173,In_456,In_163);
nor U174 (N_174,In_389,In_234);
and U175 (N_175,In_439,In_57);
xor U176 (N_176,In_362,In_311);
xor U177 (N_177,In_466,In_146);
and U178 (N_178,In_313,In_397);
nand U179 (N_179,In_123,In_345);
nor U180 (N_180,In_307,In_46);
nand U181 (N_181,In_366,In_463);
nand U182 (N_182,In_174,In_301);
nand U183 (N_183,In_448,In_393);
xor U184 (N_184,In_181,In_347);
and U185 (N_185,In_426,In_385);
or U186 (N_186,In_459,In_422);
nand U187 (N_187,In_432,In_418);
and U188 (N_188,In_309,In_390);
or U189 (N_189,In_125,In_373);
and U190 (N_190,In_147,In_408);
nand U191 (N_191,In_139,In_460);
or U192 (N_192,In_241,In_310);
or U193 (N_193,In_70,In_496);
xnor U194 (N_194,In_250,In_315);
nand U195 (N_195,In_102,In_68);
nor U196 (N_196,In_298,In_440);
nor U197 (N_197,In_26,In_37);
nand U198 (N_198,In_475,In_326);
and U199 (N_199,In_371,In_52);
nand U200 (N_200,In_20,In_338);
xor U201 (N_201,In_284,In_489);
and U202 (N_202,In_67,In_327);
nand U203 (N_203,In_490,In_177);
nor U204 (N_204,In_417,In_159);
xnor U205 (N_205,In_497,In_476);
nand U206 (N_206,In_173,In_412);
and U207 (N_207,In_290,In_89);
or U208 (N_208,In_111,In_205);
and U209 (N_209,In_447,In_425);
xor U210 (N_210,In_211,In_395);
nor U211 (N_211,In_431,In_168);
or U212 (N_212,In_429,In_435);
or U213 (N_213,In_199,In_495);
nand U214 (N_214,In_197,In_246);
or U215 (N_215,In_154,In_462);
or U216 (N_216,In_218,In_44);
and U217 (N_217,In_382,In_202);
nor U218 (N_218,In_71,In_99);
or U219 (N_219,In_28,In_194);
xor U220 (N_220,In_291,In_162);
xor U221 (N_221,In_69,In_255);
and U222 (N_222,In_277,In_251);
xor U223 (N_223,In_485,In_449);
xnor U224 (N_224,In_384,In_258);
xnor U225 (N_225,In_193,In_1);
nand U226 (N_226,In_433,In_32);
and U227 (N_227,In_294,In_381);
nand U228 (N_228,In_219,In_240);
nand U229 (N_229,In_222,In_58);
xnor U230 (N_230,In_64,In_82);
nor U231 (N_231,In_16,In_247);
or U232 (N_232,In_346,In_316);
xnor U233 (N_233,In_344,In_14);
nand U234 (N_234,In_317,In_274);
nor U235 (N_235,In_156,In_105);
nand U236 (N_236,In_325,In_36);
xnor U237 (N_237,In_103,In_402);
nand U238 (N_238,In_446,In_231);
nand U239 (N_239,In_35,In_249);
xor U240 (N_240,In_262,In_443);
and U241 (N_241,In_214,In_210);
xor U242 (N_242,In_65,In_191);
and U243 (N_243,In_12,In_95);
nor U244 (N_244,In_132,In_276);
xnor U245 (N_245,In_228,In_200);
and U246 (N_246,In_34,In_323);
nor U247 (N_247,In_304,In_157);
xor U248 (N_248,In_152,In_21);
xnor U249 (N_249,In_400,In_186);
nor U250 (N_250,In_361,In_19);
or U251 (N_251,In_304,In_203);
xor U252 (N_252,In_142,In_151);
xnor U253 (N_253,In_439,In_360);
nor U254 (N_254,In_252,In_372);
xnor U255 (N_255,In_472,In_124);
nand U256 (N_256,In_399,In_49);
nand U257 (N_257,In_298,In_50);
or U258 (N_258,In_330,In_236);
and U259 (N_259,In_327,In_221);
and U260 (N_260,In_350,In_226);
nand U261 (N_261,In_254,In_446);
nand U262 (N_262,In_58,In_126);
nand U263 (N_263,In_409,In_106);
nand U264 (N_264,In_484,In_256);
or U265 (N_265,In_249,In_390);
or U266 (N_266,In_406,In_333);
nand U267 (N_267,In_108,In_411);
nor U268 (N_268,In_35,In_449);
nor U269 (N_269,In_105,In_329);
or U270 (N_270,In_171,In_324);
xnor U271 (N_271,In_350,In_186);
xor U272 (N_272,In_229,In_493);
nand U273 (N_273,In_46,In_392);
nand U274 (N_274,In_143,In_4);
xnor U275 (N_275,In_448,In_332);
xor U276 (N_276,In_181,In_53);
or U277 (N_277,In_460,In_197);
and U278 (N_278,In_187,In_298);
and U279 (N_279,In_173,In_40);
nand U280 (N_280,In_322,In_72);
and U281 (N_281,In_364,In_180);
or U282 (N_282,In_488,In_260);
xnor U283 (N_283,In_95,In_468);
nand U284 (N_284,In_119,In_85);
or U285 (N_285,In_5,In_227);
or U286 (N_286,In_251,In_68);
nor U287 (N_287,In_187,In_394);
nor U288 (N_288,In_161,In_373);
nor U289 (N_289,In_224,In_438);
or U290 (N_290,In_458,In_137);
xnor U291 (N_291,In_462,In_248);
and U292 (N_292,In_141,In_246);
nand U293 (N_293,In_232,In_171);
or U294 (N_294,In_140,In_268);
and U295 (N_295,In_213,In_133);
nand U296 (N_296,In_382,In_198);
xnor U297 (N_297,In_254,In_174);
and U298 (N_298,In_165,In_352);
xnor U299 (N_299,In_1,In_263);
nor U300 (N_300,In_337,In_135);
and U301 (N_301,In_197,In_290);
xor U302 (N_302,In_425,In_313);
or U303 (N_303,In_136,In_392);
and U304 (N_304,In_154,In_312);
or U305 (N_305,In_209,In_431);
and U306 (N_306,In_127,In_69);
nor U307 (N_307,In_405,In_213);
and U308 (N_308,In_163,In_371);
nor U309 (N_309,In_347,In_305);
or U310 (N_310,In_474,In_457);
xor U311 (N_311,In_397,In_42);
nor U312 (N_312,In_357,In_375);
nor U313 (N_313,In_95,In_32);
xnor U314 (N_314,In_352,In_0);
nor U315 (N_315,In_36,In_128);
xnor U316 (N_316,In_41,In_254);
or U317 (N_317,In_16,In_191);
nand U318 (N_318,In_104,In_18);
xnor U319 (N_319,In_164,In_251);
and U320 (N_320,In_28,In_37);
or U321 (N_321,In_7,In_101);
nor U322 (N_322,In_159,In_402);
and U323 (N_323,In_402,In_460);
and U324 (N_324,In_156,In_39);
xnor U325 (N_325,In_420,In_119);
nand U326 (N_326,In_78,In_405);
or U327 (N_327,In_276,In_101);
xnor U328 (N_328,In_454,In_4);
nand U329 (N_329,In_129,In_67);
nor U330 (N_330,In_419,In_50);
and U331 (N_331,In_255,In_108);
and U332 (N_332,In_224,In_244);
nor U333 (N_333,In_305,In_413);
or U334 (N_334,In_452,In_350);
nor U335 (N_335,In_326,In_172);
and U336 (N_336,In_211,In_404);
nand U337 (N_337,In_175,In_203);
nand U338 (N_338,In_245,In_115);
nor U339 (N_339,In_272,In_410);
and U340 (N_340,In_315,In_228);
or U341 (N_341,In_315,In_216);
and U342 (N_342,In_446,In_25);
and U343 (N_343,In_63,In_170);
xnor U344 (N_344,In_177,In_178);
and U345 (N_345,In_429,In_483);
nor U346 (N_346,In_228,In_235);
or U347 (N_347,In_428,In_224);
nor U348 (N_348,In_245,In_358);
or U349 (N_349,In_487,In_209);
xor U350 (N_350,In_330,In_234);
nand U351 (N_351,In_298,In_332);
and U352 (N_352,In_447,In_291);
nor U353 (N_353,In_46,In_417);
or U354 (N_354,In_439,In_377);
nand U355 (N_355,In_45,In_21);
nand U356 (N_356,In_258,In_214);
nor U357 (N_357,In_174,In_146);
xnor U358 (N_358,In_337,In_444);
xnor U359 (N_359,In_234,In_111);
xnor U360 (N_360,In_200,In_59);
xor U361 (N_361,In_48,In_63);
xor U362 (N_362,In_37,In_177);
or U363 (N_363,In_489,In_167);
nor U364 (N_364,In_287,In_403);
nand U365 (N_365,In_280,In_93);
xnor U366 (N_366,In_329,In_146);
and U367 (N_367,In_338,In_191);
and U368 (N_368,In_328,In_192);
nor U369 (N_369,In_365,In_395);
or U370 (N_370,In_5,In_412);
or U371 (N_371,In_377,In_142);
xnor U372 (N_372,In_214,In_185);
xor U373 (N_373,In_258,In_133);
xor U374 (N_374,In_59,In_380);
nand U375 (N_375,In_249,In_260);
nor U376 (N_376,In_114,In_177);
nor U377 (N_377,In_286,In_17);
xor U378 (N_378,In_94,In_318);
nor U379 (N_379,In_123,In_46);
xnor U380 (N_380,In_205,In_375);
and U381 (N_381,In_140,In_37);
or U382 (N_382,In_105,In_415);
or U383 (N_383,In_275,In_246);
and U384 (N_384,In_194,In_100);
nand U385 (N_385,In_17,In_273);
nand U386 (N_386,In_109,In_277);
and U387 (N_387,In_72,In_29);
or U388 (N_388,In_445,In_141);
nand U389 (N_389,In_227,In_135);
nor U390 (N_390,In_415,In_339);
nand U391 (N_391,In_354,In_496);
or U392 (N_392,In_468,In_52);
nor U393 (N_393,In_18,In_218);
nor U394 (N_394,In_336,In_144);
xnor U395 (N_395,In_190,In_68);
or U396 (N_396,In_454,In_436);
or U397 (N_397,In_127,In_420);
and U398 (N_398,In_74,In_233);
nor U399 (N_399,In_156,In_358);
nor U400 (N_400,In_52,In_147);
nor U401 (N_401,In_440,In_330);
or U402 (N_402,In_361,In_111);
or U403 (N_403,In_253,In_375);
nand U404 (N_404,In_79,In_314);
nor U405 (N_405,In_250,In_440);
or U406 (N_406,In_487,In_261);
and U407 (N_407,In_447,In_378);
xnor U408 (N_408,In_257,In_12);
or U409 (N_409,In_132,In_126);
xor U410 (N_410,In_396,In_359);
nand U411 (N_411,In_9,In_368);
nand U412 (N_412,In_205,In_121);
or U413 (N_413,In_17,In_210);
nand U414 (N_414,In_253,In_148);
xor U415 (N_415,In_191,In_91);
nand U416 (N_416,In_69,In_91);
nor U417 (N_417,In_78,In_34);
xnor U418 (N_418,In_36,In_225);
and U419 (N_419,In_495,In_200);
and U420 (N_420,In_243,In_256);
nor U421 (N_421,In_322,In_121);
nand U422 (N_422,In_476,In_120);
nand U423 (N_423,In_322,In_406);
nor U424 (N_424,In_395,In_311);
and U425 (N_425,In_178,In_436);
nor U426 (N_426,In_203,In_455);
nand U427 (N_427,In_106,In_39);
and U428 (N_428,In_7,In_310);
xor U429 (N_429,In_213,In_336);
nor U430 (N_430,In_278,In_205);
nand U431 (N_431,In_25,In_400);
nand U432 (N_432,In_434,In_454);
xnor U433 (N_433,In_51,In_305);
nand U434 (N_434,In_12,In_120);
and U435 (N_435,In_481,In_29);
or U436 (N_436,In_172,In_125);
nor U437 (N_437,In_43,In_313);
xor U438 (N_438,In_316,In_30);
nand U439 (N_439,In_490,In_296);
xor U440 (N_440,In_69,In_78);
or U441 (N_441,In_244,In_200);
nor U442 (N_442,In_208,In_110);
nand U443 (N_443,In_279,In_27);
and U444 (N_444,In_154,In_194);
xnor U445 (N_445,In_81,In_461);
nand U446 (N_446,In_301,In_105);
and U447 (N_447,In_195,In_439);
and U448 (N_448,In_394,In_428);
xor U449 (N_449,In_157,In_101);
nor U450 (N_450,In_125,In_30);
nor U451 (N_451,In_469,In_233);
nand U452 (N_452,In_268,In_146);
and U453 (N_453,In_103,In_211);
and U454 (N_454,In_1,In_452);
or U455 (N_455,In_411,In_451);
nor U456 (N_456,In_33,In_99);
and U457 (N_457,In_45,In_355);
xor U458 (N_458,In_473,In_329);
xnor U459 (N_459,In_327,In_487);
nand U460 (N_460,In_99,In_38);
or U461 (N_461,In_226,In_335);
nor U462 (N_462,In_237,In_141);
nand U463 (N_463,In_288,In_327);
and U464 (N_464,In_395,In_199);
xor U465 (N_465,In_73,In_228);
nor U466 (N_466,In_188,In_136);
and U467 (N_467,In_276,In_62);
xnor U468 (N_468,In_404,In_314);
and U469 (N_469,In_161,In_88);
nor U470 (N_470,In_269,In_498);
or U471 (N_471,In_274,In_132);
or U472 (N_472,In_492,In_368);
nand U473 (N_473,In_390,In_329);
xor U474 (N_474,In_323,In_12);
xnor U475 (N_475,In_145,In_153);
or U476 (N_476,In_473,In_35);
nand U477 (N_477,In_478,In_392);
nor U478 (N_478,In_8,In_0);
or U479 (N_479,In_296,In_258);
nand U480 (N_480,In_468,In_356);
xnor U481 (N_481,In_47,In_48);
or U482 (N_482,In_388,In_343);
nand U483 (N_483,In_414,In_372);
nor U484 (N_484,In_446,In_156);
or U485 (N_485,In_313,In_471);
nand U486 (N_486,In_41,In_272);
nand U487 (N_487,In_127,In_116);
nand U488 (N_488,In_335,In_469);
or U489 (N_489,In_390,In_308);
xnor U490 (N_490,In_291,In_442);
nand U491 (N_491,In_4,In_378);
or U492 (N_492,In_23,In_225);
or U493 (N_493,In_57,In_194);
or U494 (N_494,In_0,In_164);
nand U495 (N_495,In_457,In_39);
and U496 (N_496,In_116,In_145);
and U497 (N_497,In_258,In_270);
nand U498 (N_498,In_278,In_133);
nand U499 (N_499,In_139,In_312);
and U500 (N_500,N_364,N_10);
and U501 (N_501,N_391,N_446);
nor U502 (N_502,N_396,N_223);
nor U503 (N_503,N_186,N_188);
xor U504 (N_504,N_202,N_171);
xnor U505 (N_505,N_363,N_31);
xor U506 (N_506,N_329,N_442);
nor U507 (N_507,N_265,N_493);
or U508 (N_508,N_343,N_407);
and U509 (N_509,N_266,N_296);
xnor U510 (N_510,N_383,N_149);
xnor U511 (N_511,N_52,N_419);
nor U512 (N_512,N_77,N_244);
xor U513 (N_513,N_7,N_35);
and U514 (N_514,N_424,N_51);
xnor U515 (N_515,N_260,N_479);
or U516 (N_516,N_57,N_434);
and U517 (N_517,N_23,N_44);
and U518 (N_518,N_9,N_5);
or U519 (N_519,N_166,N_69);
nor U520 (N_520,N_106,N_298);
nor U521 (N_521,N_382,N_6);
xnor U522 (N_522,N_344,N_195);
or U523 (N_523,N_490,N_82);
nand U524 (N_524,N_468,N_164);
nor U525 (N_525,N_375,N_270);
or U526 (N_526,N_61,N_420);
nand U527 (N_527,N_181,N_127);
xnor U528 (N_528,N_183,N_222);
nor U529 (N_529,N_131,N_198);
xor U530 (N_530,N_261,N_279);
xor U531 (N_531,N_132,N_73);
and U532 (N_532,N_399,N_193);
and U533 (N_533,N_84,N_327);
nand U534 (N_534,N_154,N_20);
nand U535 (N_535,N_205,N_315);
xnor U536 (N_536,N_301,N_303);
or U537 (N_537,N_307,N_14);
and U538 (N_538,N_397,N_176);
nor U539 (N_539,N_240,N_226);
or U540 (N_540,N_458,N_254);
and U541 (N_541,N_477,N_384);
xor U542 (N_542,N_412,N_295);
and U543 (N_543,N_237,N_361);
or U544 (N_544,N_256,N_416);
nand U545 (N_545,N_174,N_64);
nand U546 (N_546,N_107,N_109);
or U547 (N_547,N_457,N_325);
nand U548 (N_548,N_232,N_247);
and U549 (N_549,N_321,N_406);
xnor U550 (N_550,N_264,N_98);
nor U551 (N_551,N_25,N_103);
nor U552 (N_552,N_337,N_322);
nor U553 (N_553,N_481,N_354);
nand U554 (N_554,N_297,N_410);
nand U555 (N_555,N_191,N_492);
nand U556 (N_556,N_385,N_86);
nand U557 (N_557,N_224,N_283);
nand U558 (N_558,N_165,N_341);
or U559 (N_559,N_444,N_114);
xnor U560 (N_560,N_0,N_189);
and U561 (N_561,N_314,N_259);
and U562 (N_562,N_138,N_429);
xor U563 (N_563,N_286,N_278);
or U564 (N_564,N_309,N_230);
nor U565 (N_565,N_48,N_452);
xor U566 (N_566,N_494,N_87);
nand U567 (N_567,N_275,N_245);
nor U568 (N_568,N_498,N_324);
nor U569 (N_569,N_117,N_2);
and U570 (N_570,N_367,N_92);
nand U571 (N_571,N_475,N_448);
xor U572 (N_572,N_394,N_499);
xnor U573 (N_573,N_285,N_376);
or U574 (N_574,N_172,N_58);
and U575 (N_575,N_66,N_306);
xor U576 (N_576,N_393,N_464);
and U577 (N_577,N_423,N_12);
xor U578 (N_578,N_357,N_22);
nand U579 (N_579,N_157,N_252);
and U580 (N_580,N_318,N_438);
xor U581 (N_581,N_453,N_459);
or U582 (N_582,N_120,N_41);
and U583 (N_583,N_373,N_436);
xnor U584 (N_584,N_110,N_36);
xor U585 (N_585,N_276,N_352);
or U586 (N_586,N_136,N_118);
xor U587 (N_587,N_471,N_108);
xnor U588 (N_588,N_305,N_68);
xnor U589 (N_589,N_34,N_451);
nor U590 (N_590,N_351,N_160);
nor U591 (N_591,N_94,N_227);
and U592 (N_592,N_379,N_330);
and U593 (N_593,N_435,N_210);
xor U594 (N_594,N_81,N_83);
nand U595 (N_595,N_496,N_173);
nor U596 (N_596,N_70,N_30);
and U597 (N_597,N_115,N_4);
nor U598 (N_598,N_26,N_112);
nand U599 (N_599,N_17,N_428);
or U600 (N_600,N_142,N_430);
nor U601 (N_601,N_484,N_483);
nor U602 (N_602,N_105,N_190);
or U603 (N_603,N_130,N_184);
or U604 (N_604,N_241,N_233);
nor U605 (N_605,N_273,N_388);
or U606 (N_606,N_178,N_338);
nor U607 (N_607,N_390,N_111);
or U608 (N_608,N_304,N_85);
or U609 (N_609,N_93,N_345);
xnor U610 (N_610,N_439,N_179);
nor U611 (N_611,N_217,N_443);
or U612 (N_612,N_1,N_15);
and U613 (N_613,N_347,N_162);
nand U614 (N_614,N_308,N_43);
and U615 (N_615,N_139,N_284);
and U616 (N_616,N_231,N_478);
xor U617 (N_617,N_380,N_476);
xnor U618 (N_618,N_311,N_40);
nand U619 (N_619,N_269,N_146);
nor U620 (N_620,N_74,N_128);
or U621 (N_621,N_370,N_371);
or U622 (N_622,N_249,N_365);
xor U623 (N_623,N_119,N_433);
and U624 (N_624,N_491,N_248);
xor U625 (N_625,N_46,N_404);
xnor U626 (N_626,N_134,N_258);
nand U627 (N_627,N_161,N_447);
and U628 (N_628,N_113,N_200);
and U629 (N_629,N_350,N_437);
nor U630 (N_630,N_16,N_328);
nand U631 (N_631,N_408,N_213);
or U632 (N_632,N_91,N_427);
xor U633 (N_633,N_239,N_387);
and U634 (N_634,N_389,N_121);
and U635 (N_635,N_194,N_60);
nand U636 (N_636,N_280,N_169);
nor U637 (N_637,N_418,N_197);
or U638 (N_638,N_487,N_317);
nor U639 (N_639,N_495,N_455);
or U640 (N_640,N_401,N_374);
nand U641 (N_641,N_372,N_413);
and U642 (N_642,N_449,N_225);
nor U643 (N_643,N_480,N_359);
nand U644 (N_644,N_421,N_294);
nand U645 (N_645,N_145,N_79);
or U646 (N_646,N_192,N_402);
or U647 (N_647,N_211,N_462);
nor U648 (N_648,N_137,N_167);
nand U649 (N_649,N_116,N_3);
nand U650 (N_650,N_47,N_212);
xnor U651 (N_651,N_353,N_300);
nor U652 (N_652,N_168,N_182);
nand U653 (N_653,N_348,N_355);
or U654 (N_654,N_319,N_201);
xnor U655 (N_655,N_257,N_340);
nor U656 (N_656,N_155,N_485);
xor U657 (N_657,N_126,N_398);
or U658 (N_658,N_378,N_150);
nor U659 (N_659,N_246,N_268);
nor U660 (N_660,N_49,N_177);
and U661 (N_661,N_80,N_271);
and U662 (N_662,N_152,N_432);
nor U663 (N_663,N_470,N_153);
or U664 (N_664,N_219,N_71);
or U665 (N_665,N_214,N_377);
or U666 (N_666,N_59,N_469);
xor U667 (N_667,N_253,N_358);
and U668 (N_668,N_431,N_133);
nor U669 (N_669,N_11,N_33);
nand U670 (N_670,N_334,N_262);
or U671 (N_671,N_274,N_368);
or U672 (N_672,N_450,N_332);
xnor U673 (N_673,N_95,N_331);
or U674 (N_674,N_381,N_96);
or U675 (N_675,N_482,N_218);
and U676 (N_676,N_175,N_147);
nand U677 (N_677,N_38,N_461);
nor U678 (N_678,N_187,N_422);
nand U679 (N_679,N_290,N_90);
nand U680 (N_680,N_208,N_21);
nor U681 (N_681,N_124,N_441);
and U682 (N_682,N_29,N_414);
or U683 (N_683,N_221,N_488);
or U684 (N_684,N_209,N_346);
xor U685 (N_685,N_89,N_88);
nor U686 (N_686,N_288,N_466);
or U687 (N_687,N_250,N_180);
nand U688 (N_688,N_203,N_158);
or U689 (N_689,N_235,N_460);
nand U690 (N_690,N_199,N_39);
xnor U691 (N_691,N_236,N_411);
nand U692 (N_692,N_292,N_251);
and U693 (N_693,N_267,N_125);
nand U694 (N_694,N_456,N_18);
nor U695 (N_695,N_349,N_170);
and U696 (N_696,N_140,N_122);
nand U697 (N_697,N_101,N_243);
nand U698 (N_698,N_24,N_360);
nand U699 (N_699,N_141,N_299);
xor U700 (N_700,N_13,N_425);
nor U701 (N_701,N_76,N_216);
xnor U702 (N_702,N_238,N_287);
xnor U703 (N_703,N_272,N_467);
nor U704 (N_704,N_28,N_67);
nand U705 (N_705,N_206,N_473);
and U706 (N_706,N_281,N_335);
nor U707 (N_707,N_472,N_97);
and U708 (N_708,N_497,N_163);
or U709 (N_709,N_342,N_313);
nand U710 (N_710,N_310,N_339);
or U711 (N_711,N_392,N_228);
and U712 (N_712,N_282,N_56);
xnor U713 (N_713,N_242,N_417);
nand U714 (N_714,N_27,N_323);
xor U715 (N_715,N_440,N_336);
and U716 (N_716,N_291,N_289);
or U717 (N_717,N_185,N_42);
or U718 (N_718,N_143,N_489);
and U719 (N_719,N_302,N_53);
and U720 (N_720,N_99,N_104);
and U721 (N_721,N_100,N_102);
xnor U722 (N_722,N_405,N_159);
nor U723 (N_723,N_72,N_486);
nor U724 (N_724,N_220,N_445);
and U725 (N_725,N_135,N_156);
or U726 (N_726,N_333,N_129);
xor U727 (N_727,N_8,N_293);
or U728 (N_728,N_54,N_234);
nand U729 (N_729,N_229,N_362);
nor U730 (N_730,N_400,N_123);
xor U731 (N_731,N_463,N_409);
nor U732 (N_732,N_78,N_454);
and U733 (N_733,N_37,N_207);
xnor U734 (N_734,N_263,N_63);
and U735 (N_735,N_65,N_366);
nand U736 (N_736,N_312,N_426);
and U737 (N_737,N_356,N_75);
nand U738 (N_738,N_465,N_215);
and U739 (N_739,N_474,N_395);
or U740 (N_740,N_320,N_277);
nand U741 (N_741,N_151,N_196);
and U742 (N_742,N_369,N_32);
xor U743 (N_743,N_255,N_204);
xor U744 (N_744,N_415,N_62);
or U745 (N_745,N_148,N_326);
or U746 (N_746,N_45,N_144);
xor U747 (N_747,N_386,N_403);
xnor U748 (N_748,N_316,N_55);
and U749 (N_749,N_19,N_50);
nor U750 (N_750,N_14,N_431);
nor U751 (N_751,N_374,N_15);
nor U752 (N_752,N_354,N_223);
nor U753 (N_753,N_379,N_291);
xor U754 (N_754,N_151,N_494);
nand U755 (N_755,N_60,N_149);
nor U756 (N_756,N_130,N_359);
nor U757 (N_757,N_188,N_419);
nand U758 (N_758,N_303,N_165);
or U759 (N_759,N_472,N_147);
nor U760 (N_760,N_108,N_310);
xor U761 (N_761,N_141,N_331);
or U762 (N_762,N_331,N_285);
nor U763 (N_763,N_381,N_210);
xor U764 (N_764,N_264,N_407);
or U765 (N_765,N_441,N_103);
or U766 (N_766,N_56,N_174);
nor U767 (N_767,N_197,N_465);
and U768 (N_768,N_173,N_353);
nand U769 (N_769,N_103,N_423);
nor U770 (N_770,N_11,N_343);
or U771 (N_771,N_144,N_124);
or U772 (N_772,N_242,N_403);
and U773 (N_773,N_398,N_88);
and U774 (N_774,N_230,N_17);
nand U775 (N_775,N_168,N_319);
or U776 (N_776,N_461,N_141);
nor U777 (N_777,N_302,N_463);
nor U778 (N_778,N_367,N_75);
and U779 (N_779,N_213,N_239);
nor U780 (N_780,N_106,N_332);
or U781 (N_781,N_314,N_450);
or U782 (N_782,N_107,N_309);
and U783 (N_783,N_325,N_227);
xnor U784 (N_784,N_79,N_85);
nor U785 (N_785,N_319,N_219);
or U786 (N_786,N_418,N_26);
and U787 (N_787,N_414,N_40);
nand U788 (N_788,N_271,N_9);
nor U789 (N_789,N_245,N_148);
nor U790 (N_790,N_317,N_486);
xnor U791 (N_791,N_48,N_223);
or U792 (N_792,N_74,N_340);
xor U793 (N_793,N_316,N_482);
or U794 (N_794,N_295,N_495);
nor U795 (N_795,N_131,N_139);
or U796 (N_796,N_204,N_129);
and U797 (N_797,N_452,N_15);
or U798 (N_798,N_112,N_456);
nor U799 (N_799,N_351,N_383);
xnor U800 (N_800,N_289,N_283);
nor U801 (N_801,N_363,N_459);
nand U802 (N_802,N_1,N_217);
or U803 (N_803,N_379,N_228);
or U804 (N_804,N_1,N_78);
and U805 (N_805,N_118,N_187);
or U806 (N_806,N_196,N_13);
nor U807 (N_807,N_168,N_21);
and U808 (N_808,N_155,N_488);
or U809 (N_809,N_464,N_171);
or U810 (N_810,N_171,N_294);
xor U811 (N_811,N_168,N_288);
xor U812 (N_812,N_464,N_443);
and U813 (N_813,N_318,N_417);
xor U814 (N_814,N_273,N_461);
nor U815 (N_815,N_100,N_160);
nand U816 (N_816,N_163,N_382);
nand U817 (N_817,N_252,N_303);
xnor U818 (N_818,N_231,N_56);
and U819 (N_819,N_204,N_343);
nor U820 (N_820,N_36,N_27);
nor U821 (N_821,N_28,N_323);
nand U822 (N_822,N_439,N_372);
xnor U823 (N_823,N_468,N_18);
nor U824 (N_824,N_126,N_414);
xnor U825 (N_825,N_51,N_189);
xnor U826 (N_826,N_341,N_460);
nor U827 (N_827,N_337,N_34);
or U828 (N_828,N_387,N_124);
nor U829 (N_829,N_306,N_458);
or U830 (N_830,N_316,N_401);
nand U831 (N_831,N_147,N_381);
nor U832 (N_832,N_11,N_123);
nand U833 (N_833,N_447,N_350);
nand U834 (N_834,N_8,N_64);
nor U835 (N_835,N_334,N_174);
or U836 (N_836,N_496,N_56);
or U837 (N_837,N_203,N_299);
and U838 (N_838,N_370,N_420);
nand U839 (N_839,N_57,N_382);
and U840 (N_840,N_406,N_430);
nor U841 (N_841,N_88,N_38);
and U842 (N_842,N_391,N_332);
nand U843 (N_843,N_439,N_72);
xor U844 (N_844,N_129,N_20);
nor U845 (N_845,N_489,N_334);
nor U846 (N_846,N_171,N_440);
nor U847 (N_847,N_104,N_90);
xnor U848 (N_848,N_7,N_56);
or U849 (N_849,N_313,N_355);
or U850 (N_850,N_38,N_242);
or U851 (N_851,N_420,N_293);
or U852 (N_852,N_259,N_165);
and U853 (N_853,N_145,N_315);
xor U854 (N_854,N_310,N_74);
and U855 (N_855,N_300,N_143);
xnor U856 (N_856,N_200,N_333);
or U857 (N_857,N_87,N_262);
nand U858 (N_858,N_233,N_206);
nor U859 (N_859,N_130,N_142);
and U860 (N_860,N_71,N_266);
nor U861 (N_861,N_160,N_147);
and U862 (N_862,N_61,N_370);
xor U863 (N_863,N_11,N_31);
nand U864 (N_864,N_447,N_81);
and U865 (N_865,N_338,N_381);
and U866 (N_866,N_436,N_96);
xor U867 (N_867,N_139,N_347);
xnor U868 (N_868,N_145,N_168);
and U869 (N_869,N_474,N_443);
and U870 (N_870,N_494,N_462);
nor U871 (N_871,N_209,N_158);
nor U872 (N_872,N_338,N_285);
and U873 (N_873,N_102,N_367);
or U874 (N_874,N_395,N_254);
or U875 (N_875,N_345,N_243);
or U876 (N_876,N_360,N_389);
xor U877 (N_877,N_427,N_333);
or U878 (N_878,N_417,N_415);
nand U879 (N_879,N_187,N_484);
nand U880 (N_880,N_250,N_305);
or U881 (N_881,N_275,N_174);
xnor U882 (N_882,N_193,N_456);
nand U883 (N_883,N_7,N_295);
or U884 (N_884,N_171,N_90);
nand U885 (N_885,N_352,N_1);
xnor U886 (N_886,N_1,N_269);
xor U887 (N_887,N_138,N_193);
nor U888 (N_888,N_100,N_64);
nand U889 (N_889,N_457,N_353);
or U890 (N_890,N_388,N_445);
and U891 (N_891,N_337,N_372);
nor U892 (N_892,N_344,N_461);
or U893 (N_893,N_399,N_64);
xnor U894 (N_894,N_418,N_303);
xnor U895 (N_895,N_108,N_313);
nor U896 (N_896,N_357,N_337);
xnor U897 (N_897,N_133,N_141);
or U898 (N_898,N_234,N_142);
or U899 (N_899,N_338,N_43);
nor U900 (N_900,N_371,N_259);
nand U901 (N_901,N_243,N_77);
nand U902 (N_902,N_455,N_376);
xor U903 (N_903,N_165,N_138);
and U904 (N_904,N_104,N_142);
nor U905 (N_905,N_278,N_478);
nor U906 (N_906,N_259,N_297);
xnor U907 (N_907,N_428,N_403);
or U908 (N_908,N_167,N_17);
nand U909 (N_909,N_17,N_128);
and U910 (N_910,N_222,N_409);
xor U911 (N_911,N_479,N_53);
nor U912 (N_912,N_187,N_258);
or U913 (N_913,N_136,N_490);
and U914 (N_914,N_480,N_467);
and U915 (N_915,N_40,N_477);
xor U916 (N_916,N_277,N_151);
xor U917 (N_917,N_168,N_77);
nor U918 (N_918,N_372,N_282);
nor U919 (N_919,N_380,N_141);
nand U920 (N_920,N_211,N_28);
nor U921 (N_921,N_156,N_139);
nor U922 (N_922,N_352,N_421);
xor U923 (N_923,N_323,N_376);
or U924 (N_924,N_413,N_437);
nor U925 (N_925,N_384,N_479);
or U926 (N_926,N_105,N_289);
nor U927 (N_927,N_156,N_112);
xnor U928 (N_928,N_270,N_154);
xor U929 (N_929,N_254,N_428);
xor U930 (N_930,N_448,N_408);
xnor U931 (N_931,N_431,N_480);
xnor U932 (N_932,N_480,N_269);
or U933 (N_933,N_411,N_484);
and U934 (N_934,N_360,N_86);
xor U935 (N_935,N_458,N_296);
and U936 (N_936,N_48,N_292);
nor U937 (N_937,N_168,N_10);
nand U938 (N_938,N_456,N_250);
and U939 (N_939,N_62,N_115);
or U940 (N_940,N_328,N_221);
nor U941 (N_941,N_446,N_273);
nand U942 (N_942,N_162,N_397);
nand U943 (N_943,N_485,N_171);
nand U944 (N_944,N_67,N_326);
nor U945 (N_945,N_328,N_330);
nand U946 (N_946,N_434,N_156);
or U947 (N_947,N_428,N_341);
nor U948 (N_948,N_231,N_70);
nand U949 (N_949,N_309,N_88);
and U950 (N_950,N_142,N_222);
or U951 (N_951,N_80,N_89);
and U952 (N_952,N_71,N_249);
xnor U953 (N_953,N_338,N_29);
or U954 (N_954,N_297,N_95);
xnor U955 (N_955,N_150,N_205);
nor U956 (N_956,N_318,N_224);
and U957 (N_957,N_310,N_497);
nor U958 (N_958,N_124,N_64);
xnor U959 (N_959,N_177,N_213);
or U960 (N_960,N_391,N_111);
and U961 (N_961,N_97,N_118);
nand U962 (N_962,N_264,N_358);
nand U963 (N_963,N_333,N_186);
xnor U964 (N_964,N_469,N_311);
nand U965 (N_965,N_443,N_359);
nand U966 (N_966,N_147,N_12);
xnor U967 (N_967,N_284,N_360);
or U968 (N_968,N_18,N_186);
or U969 (N_969,N_3,N_478);
or U970 (N_970,N_237,N_267);
nand U971 (N_971,N_70,N_296);
xnor U972 (N_972,N_70,N_415);
nand U973 (N_973,N_398,N_261);
nor U974 (N_974,N_322,N_198);
nand U975 (N_975,N_197,N_287);
nor U976 (N_976,N_154,N_481);
nor U977 (N_977,N_81,N_174);
xnor U978 (N_978,N_252,N_457);
xnor U979 (N_979,N_41,N_201);
nor U980 (N_980,N_132,N_399);
nand U981 (N_981,N_32,N_206);
nand U982 (N_982,N_426,N_77);
or U983 (N_983,N_226,N_324);
nor U984 (N_984,N_296,N_366);
xnor U985 (N_985,N_132,N_305);
and U986 (N_986,N_160,N_396);
or U987 (N_987,N_184,N_314);
xor U988 (N_988,N_471,N_143);
xor U989 (N_989,N_438,N_350);
and U990 (N_990,N_76,N_152);
or U991 (N_991,N_369,N_307);
nor U992 (N_992,N_348,N_11);
or U993 (N_993,N_123,N_266);
and U994 (N_994,N_313,N_20);
xor U995 (N_995,N_3,N_371);
and U996 (N_996,N_478,N_37);
nand U997 (N_997,N_34,N_93);
nor U998 (N_998,N_273,N_333);
and U999 (N_999,N_220,N_194);
and U1000 (N_1000,N_521,N_850);
nand U1001 (N_1001,N_687,N_979);
and U1002 (N_1002,N_572,N_792);
nor U1003 (N_1003,N_984,N_745);
and U1004 (N_1004,N_925,N_715);
nor U1005 (N_1005,N_772,N_778);
and U1006 (N_1006,N_777,N_693);
nand U1007 (N_1007,N_591,N_871);
xor U1008 (N_1008,N_712,N_844);
nand U1009 (N_1009,N_587,N_929);
nor U1010 (N_1010,N_617,N_906);
nand U1011 (N_1011,N_508,N_868);
or U1012 (N_1012,N_806,N_663);
xor U1013 (N_1013,N_574,N_797);
nor U1014 (N_1014,N_863,N_857);
and U1015 (N_1015,N_581,N_896);
nor U1016 (N_1016,N_530,N_600);
nand U1017 (N_1017,N_773,N_755);
nor U1018 (N_1018,N_924,N_500);
and U1019 (N_1019,N_575,N_951);
or U1020 (N_1020,N_762,N_598);
xor U1021 (N_1021,N_640,N_930);
nor U1022 (N_1022,N_610,N_991);
and U1023 (N_1023,N_803,N_515);
and U1024 (N_1024,N_845,N_887);
or U1025 (N_1025,N_890,N_717);
xnor U1026 (N_1026,N_722,N_684);
nor U1027 (N_1027,N_597,N_620);
nor U1028 (N_1028,N_697,N_823);
xnor U1029 (N_1029,N_932,N_696);
xor U1030 (N_1030,N_674,N_965);
nor U1031 (N_1031,N_593,N_959);
or U1032 (N_1032,N_752,N_732);
and U1033 (N_1033,N_634,N_997);
and U1034 (N_1034,N_649,N_630);
or U1035 (N_1035,N_604,N_669);
or U1036 (N_1036,N_730,N_765);
and U1037 (N_1037,N_822,N_662);
or U1038 (N_1038,N_567,N_812);
and U1039 (N_1039,N_829,N_690);
nand U1040 (N_1040,N_681,N_731);
xnor U1041 (N_1041,N_657,N_672);
xor U1042 (N_1042,N_908,N_518);
nand U1043 (N_1043,N_677,N_854);
or U1044 (N_1044,N_665,N_769);
nor U1045 (N_1045,N_815,N_711);
xor U1046 (N_1046,N_704,N_945);
and U1047 (N_1047,N_539,N_898);
or U1048 (N_1048,N_688,N_832);
or U1049 (N_1049,N_749,N_963);
or U1050 (N_1050,N_835,N_526);
and U1051 (N_1051,N_628,N_555);
nor U1052 (N_1052,N_816,N_541);
nor U1053 (N_1053,N_897,N_580);
and U1054 (N_1054,N_960,N_577);
xnor U1055 (N_1055,N_557,N_886);
xnor U1056 (N_1056,N_987,N_758);
or U1057 (N_1057,N_830,N_912);
nor U1058 (N_1058,N_742,N_876);
or U1059 (N_1059,N_952,N_913);
and U1060 (N_1060,N_970,N_904);
nor U1061 (N_1061,N_905,N_714);
or U1062 (N_1062,N_921,N_551);
and U1063 (N_1063,N_546,N_607);
nand U1064 (N_1064,N_700,N_909);
nor U1065 (N_1065,N_942,N_888);
and U1066 (N_1066,N_759,N_736);
and U1067 (N_1067,N_972,N_667);
or U1068 (N_1068,N_535,N_611);
or U1069 (N_1069,N_976,N_757);
nor U1070 (N_1070,N_743,N_827);
and U1071 (N_1071,N_614,N_892);
nand U1072 (N_1072,N_579,N_520);
xnor U1073 (N_1073,N_721,N_708);
or U1074 (N_1074,N_689,N_622);
and U1075 (N_1075,N_872,N_613);
nand U1076 (N_1076,N_955,N_642);
nand U1077 (N_1077,N_571,N_784);
and U1078 (N_1078,N_785,N_560);
nand U1079 (N_1079,N_549,N_540);
xnor U1080 (N_1080,N_615,N_795);
xor U1081 (N_1081,N_990,N_660);
nand U1082 (N_1082,N_719,N_514);
and U1083 (N_1083,N_817,N_875);
or U1084 (N_1084,N_939,N_561);
nor U1085 (N_1085,N_701,N_973);
nor U1086 (N_1086,N_893,N_847);
nor U1087 (N_1087,N_957,N_988);
nor U1088 (N_1088,N_703,N_918);
and U1089 (N_1089,N_527,N_603);
or U1090 (N_1090,N_788,N_879);
and U1091 (N_1091,N_922,N_566);
nor U1092 (N_1092,N_947,N_969);
or U1093 (N_1093,N_501,N_946);
xnor U1094 (N_1094,N_910,N_564);
nor U1095 (N_1095,N_670,N_519);
nor U1096 (N_1096,N_691,N_837);
xnor U1097 (N_1097,N_589,N_761);
nand U1098 (N_1098,N_650,N_992);
nor U1099 (N_1099,N_986,N_744);
xnor U1100 (N_1100,N_858,N_737);
nand U1101 (N_1101,N_899,N_855);
and U1102 (N_1102,N_569,N_861);
nor U1103 (N_1103,N_768,N_920);
nand U1104 (N_1104,N_584,N_609);
or U1105 (N_1105,N_631,N_638);
xor U1106 (N_1106,N_673,N_510);
and U1107 (N_1107,N_625,N_867);
xor U1108 (N_1108,N_851,N_935);
nand U1109 (N_1109,N_683,N_629);
nor U1110 (N_1110,N_651,N_654);
or U1111 (N_1111,N_919,N_864);
nand U1112 (N_1112,N_513,N_974);
xnor U1113 (N_1113,N_636,N_917);
nand U1114 (N_1114,N_779,N_776);
xnor U1115 (N_1115,N_559,N_928);
or U1116 (N_1116,N_543,N_528);
xor U1117 (N_1117,N_729,N_900);
nor U1118 (N_1118,N_975,N_971);
or U1119 (N_1119,N_804,N_764);
nand U1120 (N_1120,N_962,N_881);
nand U1121 (N_1121,N_668,N_766);
nor U1122 (N_1122,N_658,N_841);
nand U1123 (N_1123,N_915,N_907);
or U1124 (N_1124,N_632,N_727);
and U1125 (N_1125,N_627,N_588);
nand U1126 (N_1126,N_728,N_790);
xnor U1127 (N_1127,N_968,N_709);
or U1128 (N_1128,N_570,N_516);
or U1129 (N_1129,N_506,N_767);
or U1130 (N_1130,N_751,N_583);
or U1131 (N_1131,N_801,N_914);
or U1132 (N_1132,N_882,N_695);
nand U1133 (N_1133,N_573,N_671);
xor U1134 (N_1134,N_723,N_874);
nor U1135 (N_1135,N_825,N_994);
xor U1136 (N_1136,N_750,N_739);
nand U1137 (N_1137,N_891,N_621);
and U1138 (N_1138,N_808,N_582);
nand U1139 (N_1139,N_756,N_853);
nand U1140 (N_1140,N_648,N_655);
nor U1141 (N_1141,N_878,N_941);
xor U1142 (N_1142,N_562,N_894);
nand U1143 (N_1143,N_786,N_552);
and U1144 (N_1144,N_507,N_998);
nor U1145 (N_1145,N_565,N_512);
xor U1146 (N_1146,N_558,N_706);
or U1147 (N_1147,N_926,N_568);
xor U1148 (N_1148,N_511,N_978);
nand U1149 (N_1149,N_550,N_503);
nor U1150 (N_1150,N_852,N_753);
nand U1151 (N_1151,N_537,N_680);
and U1152 (N_1152,N_661,N_787);
and U1153 (N_1153,N_834,N_999);
xor U1154 (N_1154,N_846,N_576);
and U1155 (N_1155,N_838,N_783);
xnor U1156 (N_1156,N_967,N_641);
or U1157 (N_1157,N_828,N_980);
xor U1158 (N_1158,N_545,N_517);
and U1159 (N_1159,N_809,N_664);
and U1160 (N_1160,N_800,N_839);
or U1161 (N_1161,N_694,N_702);
xor U1162 (N_1162,N_843,N_760);
nand U1163 (N_1163,N_705,N_682);
nand U1164 (N_1164,N_596,N_870);
nand U1165 (N_1165,N_977,N_633);
and U1166 (N_1166,N_889,N_509);
xnor U1167 (N_1167,N_840,N_793);
nand U1168 (N_1168,N_869,N_954);
xnor U1169 (N_1169,N_811,N_623);
nand U1170 (N_1170,N_933,N_995);
nor U1171 (N_1171,N_563,N_956);
xor U1172 (N_1172,N_985,N_590);
and U1173 (N_1173,N_848,N_547);
nor U1174 (N_1174,N_612,N_849);
xor U1175 (N_1175,N_802,N_733);
and U1176 (N_1176,N_578,N_747);
nor U1177 (N_1177,N_532,N_548);
or U1178 (N_1178,N_780,N_740);
and U1179 (N_1179,N_524,N_505);
nand U1180 (N_1180,N_877,N_504);
and U1181 (N_1181,N_798,N_554);
or U1182 (N_1182,N_544,N_653);
nand U1183 (N_1183,N_943,N_964);
or U1184 (N_1184,N_923,N_819);
nor U1185 (N_1185,N_618,N_781);
xnor U1186 (N_1186,N_934,N_646);
xnor U1187 (N_1187,N_948,N_726);
xor U1188 (N_1188,N_754,N_707);
and U1189 (N_1189,N_901,N_824);
and U1190 (N_1190,N_884,N_710);
and U1191 (N_1191,N_679,N_525);
xor U1192 (N_1192,N_866,N_799);
or U1193 (N_1193,N_652,N_666);
nand U1194 (N_1194,N_937,N_938);
or U1195 (N_1195,N_675,N_599);
or U1196 (N_1196,N_686,N_865);
nand U1197 (N_1197,N_903,N_996);
or U1198 (N_1198,N_616,N_542);
xnor U1199 (N_1199,N_813,N_531);
nand U1200 (N_1200,N_927,N_608);
nand U1201 (N_1201,N_883,N_553);
xnor U1202 (N_1202,N_953,N_763);
nor U1203 (N_1203,N_601,N_647);
and U1204 (N_1204,N_873,N_724);
and U1205 (N_1205,N_856,N_602);
nor U1206 (N_1206,N_529,N_771);
xor U1207 (N_1207,N_595,N_916);
and U1208 (N_1208,N_738,N_966);
nor U1209 (N_1209,N_534,N_944);
xnor U1210 (N_1210,N_699,N_814);
nor U1211 (N_1211,N_656,N_810);
or U1212 (N_1212,N_961,N_796);
xnor U1213 (N_1213,N_592,N_605);
or U1214 (N_1214,N_775,N_789);
nor U1215 (N_1215,N_741,N_782);
xnor U1216 (N_1216,N_626,N_842);
xnor U1217 (N_1217,N_826,N_940);
nand U1218 (N_1218,N_821,N_911);
and U1219 (N_1219,N_862,N_958);
and U1220 (N_1220,N_993,N_594);
or U1221 (N_1221,N_936,N_950);
nand U1222 (N_1222,N_746,N_533);
and U1223 (N_1223,N_836,N_820);
nand U1224 (N_1224,N_606,N_676);
and U1225 (N_1225,N_982,N_716);
nor U1226 (N_1226,N_645,N_718);
xor U1227 (N_1227,N_831,N_735);
xnor U1228 (N_1228,N_523,N_692);
and U1229 (N_1229,N_734,N_585);
or U1230 (N_1230,N_536,N_774);
xnor U1231 (N_1231,N_502,N_713);
xnor U1232 (N_1232,N_659,N_833);
or U1233 (N_1233,N_791,N_644);
nand U1234 (N_1234,N_538,N_698);
and U1235 (N_1235,N_805,N_748);
nand U1236 (N_1236,N_983,N_770);
nor U1237 (N_1237,N_639,N_931);
nand U1238 (N_1238,N_902,N_895);
nor U1239 (N_1239,N_725,N_637);
xnor U1240 (N_1240,N_989,N_685);
or U1241 (N_1241,N_720,N_860);
or U1242 (N_1242,N_643,N_807);
or U1243 (N_1243,N_859,N_624);
nor U1244 (N_1244,N_619,N_556);
nand U1245 (N_1245,N_794,N_949);
or U1246 (N_1246,N_880,N_635);
xor U1247 (N_1247,N_885,N_678);
xor U1248 (N_1248,N_586,N_818);
or U1249 (N_1249,N_981,N_522);
or U1250 (N_1250,N_595,N_748);
nand U1251 (N_1251,N_894,N_840);
or U1252 (N_1252,N_752,N_963);
xor U1253 (N_1253,N_651,N_549);
nor U1254 (N_1254,N_570,N_767);
nand U1255 (N_1255,N_820,N_717);
and U1256 (N_1256,N_791,N_824);
and U1257 (N_1257,N_674,N_902);
and U1258 (N_1258,N_505,N_940);
and U1259 (N_1259,N_613,N_844);
or U1260 (N_1260,N_541,N_651);
nor U1261 (N_1261,N_531,N_755);
nor U1262 (N_1262,N_937,N_846);
xor U1263 (N_1263,N_714,N_799);
and U1264 (N_1264,N_815,N_798);
xnor U1265 (N_1265,N_529,N_569);
nor U1266 (N_1266,N_927,N_948);
or U1267 (N_1267,N_611,N_865);
nor U1268 (N_1268,N_624,N_875);
or U1269 (N_1269,N_862,N_954);
or U1270 (N_1270,N_691,N_707);
xnor U1271 (N_1271,N_796,N_635);
nand U1272 (N_1272,N_844,N_673);
xor U1273 (N_1273,N_758,N_654);
or U1274 (N_1274,N_543,N_638);
and U1275 (N_1275,N_571,N_814);
nor U1276 (N_1276,N_837,N_968);
and U1277 (N_1277,N_573,N_733);
nand U1278 (N_1278,N_595,N_578);
and U1279 (N_1279,N_985,N_914);
nand U1280 (N_1280,N_999,N_738);
xnor U1281 (N_1281,N_793,N_608);
nand U1282 (N_1282,N_861,N_707);
nor U1283 (N_1283,N_896,N_504);
nor U1284 (N_1284,N_733,N_601);
and U1285 (N_1285,N_707,N_899);
xnor U1286 (N_1286,N_776,N_892);
or U1287 (N_1287,N_972,N_665);
nand U1288 (N_1288,N_957,N_563);
xnor U1289 (N_1289,N_666,N_596);
xor U1290 (N_1290,N_937,N_652);
and U1291 (N_1291,N_645,N_742);
nand U1292 (N_1292,N_824,N_928);
nand U1293 (N_1293,N_738,N_699);
or U1294 (N_1294,N_569,N_658);
nand U1295 (N_1295,N_676,N_602);
nand U1296 (N_1296,N_548,N_920);
or U1297 (N_1297,N_613,N_556);
xor U1298 (N_1298,N_821,N_515);
xnor U1299 (N_1299,N_906,N_510);
and U1300 (N_1300,N_895,N_638);
nor U1301 (N_1301,N_503,N_841);
nand U1302 (N_1302,N_696,N_914);
or U1303 (N_1303,N_735,N_944);
and U1304 (N_1304,N_956,N_855);
xor U1305 (N_1305,N_692,N_744);
or U1306 (N_1306,N_836,N_567);
and U1307 (N_1307,N_947,N_787);
or U1308 (N_1308,N_615,N_987);
xor U1309 (N_1309,N_642,N_715);
nor U1310 (N_1310,N_600,N_936);
nor U1311 (N_1311,N_925,N_596);
nand U1312 (N_1312,N_948,N_799);
xor U1313 (N_1313,N_679,N_522);
xor U1314 (N_1314,N_710,N_782);
xor U1315 (N_1315,N_516,N_939);
xor U1316 (N_1316,N_968,N_755);
xor U1317 (N_1317,N_788,N_573);
and U1318 (N_1318,N_569,N_630);
xnor U1319 (N_1319,N_961,N_996);
nor U1320 (N_1320,N_740,N_509);
nor U1321 (N_1321,N_889,N_725);
nor U1322 (N_1322,N_662,N_771);
and U1323 (N_1323,N_996,N_623);
nand U1324 (N_1324,N_723,N_593);
and U1325 (N_1325,N_528,N_612);
nand U1326 (N_1326,N_903,N_594);
xor U1327 (N_1327,N_937,N_963);
and U1328 (N_1328,N_635,N_919);
and U1329 (N_1329,N_913,N_978);
and U1330 (N_1330,N_706,N_610);
and U1331 (N_1331,N_822,N_732);
xor U1332 (N_1332,N_718,N_661);
xnor U1333 (N_1333,N_726,N_851);
and U1334 (N_1334,N_679,N_834);
nor U1335 (N_1335,N_882,N_694);
nand U1336 (N_1336,N_725,N_514);
or U1337 (N_1337,N_654,N_971);
nand U1338 (N_1338,N_813,N_800);
xor U1339 (N_1339,N_996,N_705);
xnor U1340 (N_1340,N_519,N_623);
nor U1341 (N_1341,N_771,N_562);
nor U1342 (N_1342,N_657,N_513);
or U1343 (N_1343,N_886,N_975);
or U1344 (N_1344,N_553,N_652);
nor U1345 (N_1345,N_764,N_690);
nand U1346 (N_1346,N_714,N_912);
nor U1347 (N_1347,N_716,N_878);
nand U1348 (N_1348,N_789,N_648);
or U1349 (N_1349,N_867,N_596);
nand U1350 (N_1350,N_675,N_605);
xor U1351 (N_1351,N_545,N_603);
xor U1352 (N_1352,N_929,N_980);
nor U1353 (N_1353,N_689,N_713);
nor U1354 (N_1354,N_709,N_886);
nand U1355 (N_1355,N_869,N_996);
xnor U1356 (N_1356,N_637,N_545);
nor U1357 (N_1357,N_962,N_686);
nor U1358 (N_1358,N_869,N_595);
or U1359 (N_1359,N_571,N_835);
and U1360 (N_1360,N_894,N_985);
nand U1361 (N_1361,N_594,N_846);
or U1362 (N_1362,N_847,N_718);
xnor U1363 (N_1363,N_924,N_837);
xnor U1364 (N_1364,N_505,N_791);
or U1365 (N_1365,N_706,N_789);
xnor U1366 (N_1366,N_751,N_875);
and U1367 (N_1367,N_975,N_991);
nand U1368 (N_1368,N_944,N_686);
xnor U1369 (N_1369,N_817,N_828);
and U1370 (N_1370,N_818,N_823);
or U1371 (N_1371,N_671,N_528);
or U1372 (N_1372,N_937,N_677);
xnor U1373 (N_1373,N_888,N_524);
nand U1374 (N_1374,N_739,N_621);
and U1375 (N_1375,N_702,N_886);
nand U1376 (N_1376,N_781,N_880);
and U1377 (N_1377,N_914,N_821);
nand U1378 (N_1378,N_713,N_520);
and U1379 (N_1379,N_672,N_590);
xnor U1380 (N_1380,N_935,N_972);
or U1381 (N_1381,N_851,N_863);
or U1382 (N_1382,N_596,N_970);
nor U1383 (N_1383,N_655,N_884);
xnor U1384 (N_1384,N_960,N_664);
nor U1385 (N_1385,N_690,N_583);
nand U1386 (N_1386,N_785,N_573);
nand U1387 (N_1387,N_979,N_691);
nand U1388 (N_1388,N_747,N_813);
and U1389 (N_1389,N_542,N_732);
and U1390 (N_1390,N_871,N_750);
or U1391 (N_1391,N_939,N_615);
xor U1392 (N_1392,N_604,N_775);
and U1393 (N_1393,N_999,N_600);
and U1394 (N_1394,N_724,N_631);
xor U1395 (N_1395,N_965,N_713);
nand U1396 (N_1396,N_591,N_672);
nor U1397 (N_1397,N_790,N_995);
nor U1398 (N_1398,N_657,N_504);
and U1399 (N_1399,N_583,N_994);
nand U1400 (N_1400,N_782,N_943);
and U1401 (N_1401,N_510,N_789);
and U1402 (N_1402,N_524,N_892);
or U1403 (N_1403,N_887,N_548);
nor U1404 (N_1404,N_645,N_719);
and U1405 (N_1405,N_746,N_797);
xor U1406 (N_1406,N_767,N_632);
or U1407 (N_1407,N_684,N_740);
xor U1408 (N_1408,N_654,N_675);
nand U1409 (N_1409,N_920,N_636);
nor U1410 (N_1410,N_752,N_549);
and U1411 (N_1411,N_568,N_919);
xnor U1412 (N_1412,N_710,N_863);
nor U1413 (N_1413,N_537,N_608);
and U1414 (N_1414,N_983,N_818);
nor U1415 (N_1415,N_991,N_970);
xnor U1416 (N_1416,N_930,N_636);
and U1417 (N_1417,N_897,N_514);
or U1418 (N_1418,N_905,N_569);
and U1419 (N_1419,N_981,N_891);
and U1420 (N_1420,N_904,N_788);
or U1421 (N_1421,N_542,N_830);
nand U1422 (N_1422,N_984,N_670);
and U1423 (N_1423,N_728,N_681);
xor U1424 (N_1424,N_816,N_870);
xnor U1425 (N_1425,N_992,N_947);
nor U1426 (N_1426,N_786,N_923);
or U1427 (N_1427,N_839,N_810);
nand U1428 (N_1428,N_759,N_953);
nor U1429 (N_1429,N_787,N_590);
or U1430 (N_1430,N_988,N_605);
xor U1431 (N_1431,N_583,N_727);
nand U1432 (N_1432,N_525,N_589);
xor U1433 (N_1433,N_914,N_647);
and U1434 (N_1434,N_555,N_754);
xor U1435 (N_1435,N_714,N_926);
nor U1436 (N_1436,N_822,N_893);
nand U1437 (N_1437,N_757,N_604);
nand U1438 (N_1438,N_780,N_997);
and U1439 (N_1439,N_890,N_607);
and U1440 (N_1440,N_717,N_644);
nor U1441 (N_1441,N_862,N_698);
xor U1442 (N_1442,N_744,N_817);
xnor U1443 (N_1443,N_712,N_657);
and U1444 (N_1444,N_806,N_805);
xnor U1445 (N_1445,N_912,N_639);
nand U1446 (N_1446,N_901,N_781);
nor U1447 (N_1447,N_538,N_602);
and U1448 (N_1448,N_572,N_771);
and U1449 (N_1449,N_757,N_946);
nand U1450 (N_1450,N_953,N_632);
nand U1451 (N_1451,N_771,N_683);
xor U1452 (N_1452,N_908,N_507);
nor U1453 (N_1453,N_572,N_740);
xor U1454 (N_1454,N_885,N_652);
and U1455 (N_1455,N_529,N_680);
nand U1456 (N_1456,N_551,N_899);
xor U1457 (N_1457,N_726,N_774);
xnor U1458 (N_1458,N_714,N_979);
xor U1459 (N_1459,N_882,N_939);
nor U1460 (N_1460,N_795,N_902);
and U1461 (N_1461,N_646,N_949);
and U1462 (N_1462,N_911,N_935);
xor U1463 (N_1463,N_893,N_998);
xnor U1464 (N_1464,N_831,N_565);
xnor U1465 (N_1465,N_977,N_627);
and U1466 (N_1466,N_538,N_850);
or U1467 (N_1467,N_768,N_733);
xnor U1468 (N_1468,N_947,N_639);
and U1469 (N_1469,N_774,N_670);
and U1470 (N_1470,N_875,N_706);
nand U1471 (N_1471,N_974,N_934);
and U1472 (N_1472,N_717,N_641);
and U1473 (N_1473,N_531,N_684);
nand U1474 (N_1474,N_862,N_830);
nor U1475 (N_1475,N_799,N_926);
or U1476 (N_1476,N_583,N_895);
nand U1477 (N_1477,N_827,N_807);
nor U1478 (N_1478,N_995,N_834);
and U1479 (N_1479,N_976,N_912);
nor U1480 (N_1480,N_836,N_975);
nor U1481 (N_1481,N_693,N_514);
nor U1482 (N_1482,N_908,N_691);
and U1483 (N_1483,N_698,N_968);
nand U1484 (N_1484,N_700,N_503);
nand U1485 (N_1485,N_836,N_553);
nor U1486 (N_1486,N_820,N_509);
nand U1487 (N_1487,N_602,N_934);
xnor U1488 (N_1488,N_840,N_747);
or U1489 (N_1489,N_801,N_777);
or U1490 (N_1490,N_732,N_707);
xor U1491 (N_1491,N_997,N_688);
and U1492 (N_1492,N_657,N_503);
nand U1493 (N_1493,N_923,N_859);
and U1494 (N_1494,N_857,N_573);
nand U1495 (N_1495,N_842,N_885);
nor U1496 (N_1496,N_502,N_958);
and U1497 (N_1497,N_685,N_627);
xnor U1498 (N_1498,N_502,N_508);
xor U1499 (N_1499,N_602,N_746);
and U1500 (N_1500,N_1416,N_1215);
and U1501 (N_1501,N_1339,N_1028);
or U1502 (N_1502,N_1213,N_1033);
xor U1503 (N_1503,N_1048,N_1266);
nor U1504 (N_1504,N_1248,N_1024);
or U1505 (N_1505,N_1143,N_1447);
and U1506 (N_1506,N_1167,N_1351);
or U1507 (N_1507,N_1050,N_1274);
and U1508 (N_1508,N_1346,N_1265);
or U1509 (N_1509,N_1377,N_1180);
and U1510 (N_1510,N_1086,N_1078);
nand U1511 (N_1511,N_1343,N_1103);
nand U1512 (N_1512,N_1119,N_1304);
and U1513 (N_1513,N_1002,N_1275);
or U1514 (N_1514,N_1132,N_1185);
xor U1515 (N_1515,N_1127,N_1195);
xnor U1516 (N_1516,N_1191,N_1374);
or U1517 (N_1517,N_1146,N_1397);
or U1518 (N_1518,N_1294,N_1223);
nand U1519 (N_1519,N_1034,N_1417);
or U1520 (N_1520,N_1237,N_1403);
xnor U1521 (N_1521,N_1067,N_1053);
xor U1522 (N_1522,N_1211,N_1197);
or U1523 (N_1523,N_1329,N_1101);
nor U1524 (N_1524,N_1272,N_1220);
nor U1525 (N_1525,N_1059,N_1031);
nor U1526 (N_1526,N_1171,N_1254);
xnor U1527 (N_1527,N_1009,N_1462);
or U1528 (N_1528,N_1070,N_1268);
nand U1529 (N_1529,N_1432,N_1150);
nor U1530 (N_1530,N_1301,N_1169);
nand U1531 (N_1531,N_1423,N_1310);
or U1532 (N_1532,N_1194,N_1173);
and U1533 (N_1533,N_1300,N_1056);
xnor U1534 (N_1534,N_1141,N_1456);
nor U1535 (N_1535,N_1434,N_1362);
or U1536 (N_1536,N_1096,N_1198);
or U1537 (N_1537,N_1473,N_1044);
nor U1538 (N_1538,N_1262,N_1359);
nor U1539 (N_1539,N_1023,N_1499);
nand U1540 (N_1540,N_1270,N_1394);
nand U1541 (N_1541,N_1155,N_1179);
nand U1542 (N_1542,N_1085,N_1322);
nor U1543 (N_1543,N_1207,N_1235);
nand U1544 (N_1544,N_1095,N_1130);
nor U1545 (N_1545,N_1321,N_1226);
nand U1546 (N_1546,N_1421,N_1384);
or U1547 (N_1547,N_1071,N_1126);
or U1548 (N_1548,N_1001,N_1174);
and U1549 (N_1549,N_1135,N_1260);
xnor U1550 (N_1550,N_1381,N_1243);
nand U1551 (N_1551,N_1388,N_1252);
and U1552 (N_1552,N_1204,N_1413);
nand U1553 (N_1553,N_1344,N_1145);
nand U1554 (N_1554,N_1016,N_1396);
xnor U1555 (N_1555,N_1291,N_1478);
and U1556 (N_1556,N_1389,N_1225);
nand U1557 (N_1557,N_1057,N_1289);
xnor U1558 (N_1558,N_1458,N_1046);
nand U1559 (N_1559,N_1365,N_1232);
nor U1560 (N_1560,N_1054,N_1282);
or U1561 (N_1561,N_1350,N_1429);
or U1562 (N_1562,N_1228,N_1151);
or U1563 (N_1563,N_1172,N_1099);
nand U1564 (N_1564,N_1247,N_1315);
and U1565 (N_1565,N_1334,N_1401);
and U1566 (N_1566,N_1007,N_1214);
nand U1567 (N_1567,N_1476,N_1333);
xnor U1568 (N_1568,N_1387,N_1409);
and U1569 (N_1569,N_1457,N_1330);
and U1570 (N_1570,N_1287,N_1307);
nor U1571 (N_1571,N_1245,N_1349);
or U1572 (N_1572,N_1471,N_1088);
xnor U1573 (N_1573,N_1345,N_1355);
nor U1574 (N_1574,N_1182,N_1391);
or U1575 (N_1575,N_1039,N_1075);
or U1576 (N_1576,N_1133,N_1335);
nor U1577 (N_1577,N_1372,N_1368);
nor U1578 (N_1578,N_1443,N_1450);
xnor U1579 (N_1579,N_1393,N_1227);
nand U1580 (N_1580,N_1183,N_1414);
and U1581 (N_1581,N_1410,N_1159);
or U1582 (N_1582,N_1113,N_1149);
xnor U1583 (N_1583,N_1285,N_1255);
and U1584 (N_1584,N_1358,N_1115);
xnor U1585 (N_1585,N_1383,N_1461);
nor U1586 (N_1586,N_1200,N_1206);
or U1587 (N_1587,N_1222,N_1418);
and U1588 (N_1588,N_1470,N_1336);
or U1589 (N_1589,N_1292,N_1273);
xnor U1590 (N_1590,N_1297,N_1486);
nor U1591 (N_1591,N_1490,N_1382);
nand U1592 (N_1592,N_1010,N_1224);
and U1593 (N_1593,N_1452,N_1229);
xnor U1594 (N_1594,N_1128,N_1072);
nor U1595 (N_1595,N_1385,N_1323);
or U1596 (N_1596,N_1314,N_1079);
xnor U1597 (N_1597,N_1332,N_1316);
xnor U1598 (N_1598,N_1014,N_1110);
nor U1599 (N_1599,N_1481,N_1049);
xnor U1600 (N_1600,N_1459,N_1451);
nor U1601 (N_1601,N_1440,N_1152);
nor U1602 (N_1602,N_1188,N_1361);
nor U1603 (N_1603,N_1011,N_1186);
and U1604 (N_1604,N_1045,N_1123);
nand U1605 (N_1605,N_1318,N_1308);
or U1606 (N_1606,N_1295,N_1276);
and U1607 (N_1607,N_1106,N_1267);
nand U1608 (N_1608,N_1453,N_1463);
and U1609 (N_1609,N_1148,N_1497);
nor U1610 (N_1610,N_1092,N_1379);
and U1611 (N_1611,N_1455,N_1269);
nand U1612 (N_1612,N_1436,N_1375);
and U1613 (N_1613,N_1062,N_1153);
nand U1614 (N_1614,N_1217,N_1311);
xor U1615 (N_1615,N_1472,N_1154);
and U1616 (N_1616,N_1430,N_1063);
nand U1617 (N_1617,N_1138,N_1166);
nand U1618 (N_1618,N_1105,N_1129);
or U1619 (N_1619,N_1017,N_1058);
xnor U1620 (N_1620,N_1283,N_1352);
xnor U1621 (N_1621,N_1250,N_1040);
nor U1622 (N_1622,N_1124,N_1111);
nand U1623 (N_1623,N_1036,N_1491);
xor U1624 (N_1624,N_1264,N_1331);
nor U1625 (N_1625,N_1277,N_1077);
xnor U1626 (N_1626,N_1032,N_1395);
and U1627 (N_1627,N_1003,N_1425);
and U1628 (N_1628,N_1411,N_1064);
nand U1629 (N_1629,N_1437,N_1445);
xor U1630 (N_1630,N_1068,N_1464);
nor U1631 (N_1631,N_1249,N_1373);
nor U1632 (N_1632,N_1156,N_1340);
or U1633 (N_1633,N_1137,N_1134);
or U1634 (N_1634,N_1242,N_1390);
nor U1635 (N_1635,N_1469,N_1114);
xor U1636 (N_1636,N_1027,N_1366);
nand U1637 (N_1637,N_1427,N_1231);
and U1638 (N_1638,N_1378,N_1131);
or U1639 (N_1639,N_1326,N_1042);
nand U1640 (N_1640,N_1446,N_1082);
xnor U1641 (N_1641,N_1319,N_1238);
xor U1642 (N_1642,N_1158,N_1051);
or U1643 (N_1643,N_1348,N_1052);
and U1644 (N_1644,N_1439,N_1073);
xnor U1645 (N_1645,N_1369,N_1233);
and U1646 (N_1646,N_1426,N_1162);
xnor U1647 (N_1647,N_1398,N_1431);
nand U1648 (N_1648,N_1176,N_1196);
nor U1649 (N_1649,N_1354,N_1083);
or U1650 (N_1650,N_1177,N_1000);
nand U1651 (N_1651,N_1239,N_1121);
and U1652 (N_1652,N_1107,N_1263);
nand U1653 (N_1653,N_1454,N_1221);
or U1654 (N_1654,N_1407,N_1139);
xnor U1655 (N_1655,N_1018,N_1261);
and U1656 (N_1656,N_1097,N_1312);
and U1657 (N_1657,N_1192,N_1412);
or U1658 (N_1658,N_1386,N_1482);
nor U1659 (N_1659,N_1466,N_1256);
and U1660 (N_1660,N_1100,N_1371);
nor U1661 (N_1661,N_1306,N_1147);
or U1662 (N_1662,N_1399,N_1298);
xor U1663 (N_1663,N_1424,N_1120);
xor U1664 (N_1664,N_1030,N_1404);
and U1665 (N_1665,N_1029,N_1015);
and U1666 (N_1666,N_1420,N_1433);
or U1667 (N_1667,N_1234,N_1193);
nand U1668 (N_1668,N_1047,N_1157);
xor U1669 (N_1669,N_1109,N_1498);
and U1670 (N_1670,N_1244,N_1094);
nand U1671 (N_1671,N_1325,N_1069);
or U1672 (N_1672,N_1038,N_1025);
nand U1673 (N_1673,N_1118,N_1184);
or U1674 (N_1674,N_1376,N_1074);
or U1675 (N_1675,N_1091,N_1367);
nand U1676 (N_1676,N_1444,N_1286);
or U1677 (N_1677,N_1019,N_1483);
nor U1678 (N_1678,N_1468,N_1302);
nor U1679 (N_1679,N_1415,N_1013);
nand U1680 (N_1680,N_1202,N_1363);
nor U1681 (N_1681,N_1144,N_1303);
nor U1682 (N_1682,N_1380,N_1280);
xor U1683 (N_1683,N_1210,N_1278);
and U1684 (N_1684,N_1108,N_1093);
or U1685 (N_1685,N_1465,N_1102);
or U1686 (N_1686,N_1136,N_1435);
or U1687 (N_1687,N_1246,N_1161);
nand U1688 (N_1688,N_1008,N_1338);
and U1689 (N_1689,N_1125,N_1060);
or U1690 (N_1690,N_1405,N_1284);
nor U1691 (N_1691,N_1485,N_1087);
or U1692 (N_1692,N_1178,N_1496);
nor U1693 (N_1693,N_1089,N_1189);
nor U1694 (N_1694,N_1474,N_1449);
and U1695 (N_1695,N_1112,N_1020);
nor U1696 (N_1696,N_1309,N_1219);
and U1697 (N_1697,N_1342,N_1317);
and U1698 (N_1698,N_1104,N_1084);
nand U1699 (N_1699,N_1006,N_1324);
nor U1700 (N_1700,N_1035,N_1216);
or U1701 (N_1701,N_1203,N_1187);
and U1702 (N_1702,N_1175,N_1392);
and U1703 (N_1703,N_1259,N_1199);
or U1704 (N_1704,N_1477,N_1026);
xor U1705 (N_1705,N_1168,N_1037);
nand U1706 (N_1706,N_1438,N_1253);
xor U1707 (N_1707,N_1208,N_1489);
and U1708 (N_1708,N_1212,N_1021);
nand U1709 (N_1709,N_1328,N_1305);
nand U1710 (N_1710,N_1117,N_1061);
or U1711 (N_1711,N_1055,N_1364);
and U1712 (N_1712,N_1479,N_1041);
or U1713 (N_1713,N_1251,N_1043);
nand U1714 (N_1714,N_1205,N_1370);
nand U1715 (N_1715,N_1240,N_1460);
nor U1716 (N_1716,N_1288,N_1065);
or U1717 (N_1717,N_1441,N_1090);
or U1718 (N_1718,N_1442,N_1160);
nor U1719 (N_1719,N_1494,N_1492);
xnor U1720 (N_1720,N_1258,N_1209);
nor U1721 (N_1721,N_1004,N_1356);
nand U1722 (N_1722,N_1281,N_1066);
nand U1723 (N_1723,N_1290,N_1142);
xor U1724 (N_1724,N_1320,N_1122);
nor U1725 (N_1725,N_1279,N_1230);
xnor U1726 (N_1726,N_1293,N_1357);
or U1727 (N_1727,N_1487,N_1408);
nand U1728 (N_1728,N_1327,N_1012);
or U1729 (N_1729,N_1005,N_1428);
or U1730 (N_1730,N_1313,N_1218);
or U1731 (N_1731,N_1480,N_1257);
nand U1732 (N_1732,N_1341,N_1353);
and U1733 (N_1733,N_1022,N_1165);
nor U1734 (N_1734,N_1190,N_1406);
and U1735 (N_1735,N_1163,N_1495);
nand U1736 (N_1736,N_1181,N_1493);
nor U1737 (N_1737,N_1076,N_1241);
and U1738 (N_1738,N_1488,N_1337);
or U1739 (N_1739,N_1419,N_1271);
and U1740 (N_1740,N_1116,N_1484);
or U1741 (N_1741,N_1081,N_1140);
xnor U1742 (N_1742,N_1080,N_1448);
and U1743 (N_1743,N_1475,N_1299);
nor U1744 (N_1744,N_1170,N_1400);
nor U1745 (N_1745,N_1296,N_1347);
xor U1746 (N_1746,N_1164,N_1236);
nor U1747 (N_1747,N_1201,N_1402);
and U1748 (N_1748,N_1422,N_1098);
xnor U1749 (N_1749,N_1467,N_1360);
xnor U1750 (N_1750,N_1119,N_1483);
nand U1751 (N_1751,N_1462,N_1170);
nor U1752 (N_1752,N_1032,N_1088);
nand U1753 (N_1753,N_1359,N_1431);
or U1754 (N_1754,N_1075,N_1034);
nor U1755 (N_1755,N_1315,N_1431);
or U1756 (N_1756,N_1402,N_1432);
xor U1757 (N_1757,N_1467,N_1349);
or U1758 (N_1758,N_1440,N_1298);
and U1759 (N_1759,N_1369,N_1346);
or U1760 (N_1760,N_1071,N_1386);
nand U1761 (N_1761,N_1435,N_1059);
or U1762 (N_1762,N_1225,N_1388);
xor U1763 (N_1763,N_1118,N_1493);
nor U1764 (N_1764,N_1337,N_1046);
or U1765 (N_1765,N_1071,N_1329);
and U1766 (N_1766,N_1298,N_1028);
or U1767 (N_1767,N_1472,N_1192);
nand U1768 (N_1768,N_1172,N_1171);
nand U1769 (N_1769,N_1300,N_1304);
nand U1770 (N_1770,N_1389,N_1076);
nand U1771 (N_1771,N_1172,N_1070);
or U1772 (N_1772,N_1340,N_1138);
or U1773 (N_1773,N_1397,N_1494);
nor U1774 (N_1774,N_1254,N_1322);
nor U1775 (N_1775,N_1107,N_1308);
xnor U1776 (N_1776,N_1186,N_1018);
nor U1777 (N_1777,N_1422,N_1276);
or U1778 (N_1778,N_1270,N_1062);
or U1779 (N_1779,N_1203,N_1323);
xor U1780 (N_1780,N_1487,N_1407);
xnor U1781 (N_1781,N_1290,N_1321);
or U1782 (N_1782,N_1349,N_1017);
nor U1783 (N_1783,N_1179,N_1008);
nand U1784 (N_1784,N_1052,N_1147);
xor U1785 (N_1785,N_1239,N_1096);
nor U1786 (N_1786,N_1361,N_1145);
nand U1787 (N_1787,N_1356,N_1351);
and U1788 (N_1788,N_1196,N_1115);
and U1789 (N_1789,N_1394,N_1300);
or U1790 (N_1790,N_1489,N_1388);
or U1791 (N_1791,N_1269,N_1042);
xnor U1792 (N_1792,N_1464,N_1150);
nand U1793 (N_1793,N_1471,N_1001);
nor U1794 (N_1794,N_1394,N_1224);
or U1795 (N_1795,N_1323,N_1235);
xor U1796 (N_1796,N_1333,N_1202);
xor U1797 (N_1797,N_1166,N_1263);
nand U1798 (N_1798,N_1319,N_1425);
or U1799 (N_1799,N_1369,N_1300);
nand U1800 (N_1800,N_1142,N_1164);
and U1801 (N_1801,N_1374,N_1489);
xor U1802 (N_1802,N_1180,N_1032);
nor U1803 (N_1803,N_1285,N_1256);
or U1804 (N_1804,N_1177,N_1265);
nand U1805 (N_1805,N_1011,N_1090);
nor U1806 (N_1806,N_1376,N_1043);
nor U1807 (N_1807,N_1038,N_1099);
xnor U1808 (N_1808,N_1285,N_1455);
and U1809 (N_1809,N_1297,N_1275);
or U1810 (N_1810,N_1377,N_1294);
or U1811 (N_1811,N_1327,N_1137);
or U1812 (N_1812,N_1426,N_1002);
or U1813 (N_1813,N_1101,N_1481);
xor U1814 (N_1814,N_1447,N_1314);
nor U1815 (N_1815,N_1496,N_1481);
nor U1816 (N_1816,N_1193,N_1091);
and U1817 (N_1817,N_1308,N_1333);
nor U1818 (N_1818,N_1228,N_1054);
nor U1819 (N_1819,N_1295,N_1158);
xnor U1820 (N_1820,N_1495,N_1159);
and U1821 (N_1821,N_1448,N_1409);
xor U1822 (N_1822,N_1290,N_1224);
and U1823 (N_1823,N_1345,N_1105);
and U1824 (N_1824,N_1342,N_1050);
and U1825 (N_1825,N_1425,N_1158);
xor U1826 (N_1826,N_1386,N_1440);
and U1827 (N_1827,N_1451,N_1356);
nor U1828 (N_1828,N_1140,N_1390);
nand U1829 (N_1829,N_1047,N_1020);
and U1830 (N_1830,N_1150,N_1278);
and U1831 (N_1831,N_1127,N_1105);
or U1832 (N_1832,N_1159,N_1136);
xor U1833 (N_1833,N_1066,N_1063);
and U1834 (N_1834,N_1206,N_1231);
nand U1835 (N_1835,N_1074,N_1123);
or U1836 (N_1836,N_1414,N_1028);
nand U1837 (N_1837,N_1049,N_1047);
nand U1838 (N_1838,N_1252,N_1450);
and U1839 (N_1839,N_1137,N_1127);
nor U1840 (N_1840,N_1148,N_1345);
xnor U1841 (N_1841,N_1148,N_1177);
nor U1842 (N_1842,N_1022,N_1258);
and U1843 (N_1843,N_1203,N_1425);
nand U1844 (N_1844,N_1077,N_1437);
nor U1845 (N_1845,N_1186,N_1375);
or U1846 (N_1846,N_1464,N_1441);
nor U1847 (N_1847,N_1282,N_1345);
nor U1848 (N_1848,N_1255,N_1183);
xor U1849 (N_1849,N_1159,N_1225);
nand U1850 (N_1850,N_1361,N_1293);
xnor U1851 (N_1851,N_1216,N_1030);
and U1852 (N_1852,N_1497,N_1099);
or U1853 (N_1853,N_1043,N_1124);
nand U1854 (N_1854,N_1437,N_1289);
nor U1855 (N_1855,N_1181,N_1005);
xor U1856 (N_1856,N_1238,N_1146);
xnor U1857 (N_1857,N_1382,N_1424);
nand U1858 (N_1858,N_1429,N_1320);
nor U1859 (N_1859,N_1381,N_1285);
nand U1860 (N_1860,N_1120,N_1123);
or U1861 (N_1861,N_1144,N_1405);
or U1862 (N_1862,N_1463,N_1447);
nand U1863 (N_1863,N_1053,N_1058);
nor U1864 (N_1864,N_1199,N_1223);
xor U1865 (N_1865,N_1212,N_1165);
and U1866 (N_1866,N_1289,N_1083);
nand U1867 (N_1867,N_1366,N_1110);
nand U1868 (N_1868,N_1224,N_1428);
xnor U1869 (N_1869,N_1464,N_1020);
nand U1870 (N_1870,N_1338,N_1208);
and U1871 (N_1871,N_1047,N_1089);
or U1872 (N_1872,N_1382,N_1481);
nand U1873 (N_1873,N_1337,N_1412);
and U1874 (N_1874,N_1479,N_1362);
nor U1875 (N_1875,N_1211,N_1200);
xnor U1876 (N_1876,N_1232,N_1489);
nand U1877 (N_1877,N_1096,N_1067);
nor U1878 (N_1878,N_1270,N_1131);
nor U1879 (N_1879,N_1369,N_1382);
or U1880 (N_1880,N_1446,N_1309);
or U1881 (N_1881,N_1491,N_1449);
and U1882 (N_1882,N_1220,N_1494);
and U1883 (N_1883,N_1128,N_1426);
xor U1884 (N_1884,N_1187,N_1189);
or U1885 (N_1885,N_1326,N_1013);
or U1886 (N_1886,N_1100,N_1431);
xnor U1887 (N_1887,N_1280,N_1477);
nor U1888 (N_1888,N_1485,N_1044);
and U1889 (N_1889,N_1044,N_1460);
nor U1890 (N_1890,N_1423,N_1019);
or U1891 (N_1891,N_1369,N_1187);
nor U1892 (N_1892,N_1371,N_1214);
nand U1893 (N_1893,N_1324,N_1099);
xnor U1894 (N_1894,N_1022,N_1175);
nor U1895 (N_1895,N_1155,N_1234);
or U1896 (N_1896,N_1239,N_1080);
and U1897 (N_1897,N_1156,N_1231);
xor U1898 (N_1898,N_1093,N_1182);
xnor U1899 (N_1899,N_1451,N_1202);
or U1900 (N_1900,N_1366,N_1011);
and U1901 (N_1901,N_1322,N_1191);
xnor U1902 (N_1902,N_1022,N_1380);
nor U1903 (N_1903,N_1303,N_1433);
nand U1904 (N_1904,N_1078,N_1489);
nand U1905 (N_1905,N_1418,N_1057);
nor U1906 (N_1906,N_1113,N_1385);
xor U1907 (N_1907,N_1153,N_1276);
and U1908 (N_1908,N_1172,N_1187);
nor U1909 (N_1909,N_1312,N_1142);
nor U1910 (N_1910,N_1465,N_1371);
or U1911 (N_1911,N_1217,N_1168);
or U1912 (N_1912,N_1111,N_1478);
or U1913 (N_1913,N_1193,N_1485);
or U1914 (N_1914,N_1279,N_1412);
and U1915 (N_1915,N_1038,N_1441);
nand U1916 (N_1916,N_1025,N_1428);
xnor U1917 (N_1917,N_1010,N_1318);
xnor U1918 (N_1918,N_1488,N_1275);
or U1919 (N_1919,N_1104,N_1453);
and U1920 (N_1920,N_1014,N_1235);
nor U1921 (N_1921,N_1447,N_1096);
xor U1922 (N_1922,N_1001,N_1028);
nor U1923 (N_1923,N_1099,N_1069);
xnor U1924 (N_1924,N_1474,N_1304);
nand U1925 (N_1925,N_1367,N_1281);
nor U1926 (N_1926,N_1273,N_1073);
or U1927 (N_1927,N_1140,N_1263);
xnor U1928 (N_1928,N_1314,N_1393);
nor U1929 (N_1929,N_1203,N_1006);
nand U1930 (N_1930,N_1106,N_1351);
xnor U1931 (N_1931,N_1314,N_1117);
or U1932 (N_1932,N_1200,N_1281);
and U1933 (N_1933,N_1198,N_1166);
nand U1934 (N_1934,N_1322,N_1495);
xnor U1935 (N_1935,N_1246,N_1171);
xor U1936 (N_1936,N_1322,N_1050);
nor U1937 (N_1937,N_1131,N_1476);
and U1938 (N_1938,N_1432,N_1418);
or U1939 (N_1939,N_1451,N_1485);
nor U1940 (N_1940,N_1308,N_1031);
or U1941 (N_1941,N_1373,N_1155);
nor U1942 (N_1942,N_1211,N_1068);
nand U1943 (N_1943,N_1373,N_1487);
and U1944 (N_1944,N_1390,N_1144);
nor U1945 (N_1945,N_1331,N_1249);
and U1946 (N_1946,N_1393,N_1384);
xnor U1947 (N_1947,N_1103,N_1169);
or U1948 (N_1948,N_1022,N_1375);
nand U1949 (N_1949,N_1047,N_1084);
or U1950 (N_1950,N_1327,N_1337);
nor U1951 (N_1951,N_1309,N_1109);
nor U1952 (N_1952,N_1078,N_1092);
nor U1953 (N_1953,N_1484,N_1010);
xnor U1954 (N_1954,N_1452,N_1157);
nor U1955 (N_1955,N_1255,N_1153);
nor U1956 (N_1956,N_1130,N_1317);
nand U1957 (N_1957,N_1358,N_1367);
xnor U1958 (N_1958,N_1275,N_1293);
or U1959 (N_1959,N_1132,N_1247);
xnor U1960 (N_1960,N_1297,N_1449);
and U1961 (N_1961,N_1068,N_1438);
xnor U1962 (N_1962,N_1087,N_1351);
xnor U1963 (N_1963,N_1004,N_1310);
nor U1964 (N_1964,N_1053,N_1440);
nor U1965 (N_1965,N_1165,N_1100);
nand U1966 (N_1966,N_1024,N_1386);
nor U1967 (N_1967,N_1010,N_1258);
nand U1968 (N_1968,N_1480,N_1146);
and U1969 (N_1969,N_1313,N_1419);
nand U1970 (N_1970,N_1050,N_1306);
xnor U1971 (N_1971,N_1353,N_1061);
nor U1972 (N_1972,N_1205,N_1347);
nor U1973 (N_1973,N_1079,N_1343);
or U1974 (N_1974,N_1089,N_1353);
xor U1975 (N_1975,N_1136,N_1383);
nand U1976 (N_1976,N_1040,N_1492);
nand U1977 (N_1977,N_1348,N_1113);
nor U1978 (N_1978,N_1330,N_1140);
and U1979 (N_1979,N_1127,N_1223);
nand U1980 (N_1980,N_1394,N_1053);
and U1981 (N_1981,N_1175,N_1339);
xnor U1982 (N_1982,N_1436,N_1277);
or U1983 (N_1983,N_1239,N_1284);
and U1984 (N_1984,N_1415,N_1277);
nand U1985 (N_1985,N_1427,N_1165);
or U1986 (N_1986,N_1238,N_1214);
nor U1987 (N_1987,N_1255,N_1179);
nor U1988 (N_1988,N_1144,N_1177);
nand U1989 (N_1989,N_1425,N_1242);
xnor U1990 (N_1990,N_1487,N_1101);
or U1991 (N_1991,N_1341,N_1036);
nand U1992 (N_1992,N_1315,N_1181);
nand U1993 (N_1993,N_1487,N_1190);
nand U1994 (N_1994,N_1180,N_1482);
nand U1995 (N_1995,N_1053,N_1005);
nor U1996 (N_1996,N_1471,N_1145);
and U1997 (N_1997,N_1194,N_1388);
or U1998 (N_1998,N_1173,N_1124);
and U1999 (N_1999,N_1494,N_1240);
xnor U2000 (N_2000,N_1925,N_1856);
or U2001 (N_2001,N_1891,N_1559);
xor U2002 (N_2002,N_1930,N_1591);
or U2003 (N_2003,N_1870,N_1893);
and U2004 (N_2004,N_1763,N_1949);
xnor U2005 (N_2005,N_1954,N_1619);
or U2006 (N_2006,N_1741,N_1698);
nor U2007 (N_2007,N_1672,N_1509);
xnor U2008 (N_2008,N_1775,N_1734);
or U2009 (N_2009,N_1529,N_1759);
and U2010 (N_2010,N_1609,N_1620);
nor U2011 (N_2011,N_1952,N_1669);
xnor U2012 (N_2012,N_1661,N_1535);
and U2013 (N_2013,N_1504,N_1629);
or U2014 (N_2014,N_1543,N_1625);
xnor U2015 (N_2015,N_1566,N_1875);
nor U2016 (N_2016,N_1674,N_1912);
or U2017 (N_2017,N_1867,N_1686);
nand U2018 (N_2018,N_1809,N_1935);
or U2019 (N_2019,N_1712,N_1731);
nand U2020 (N_2020,N_1506,N_1719);
and U2021 (N_2021,N_1804,N_1917);
and U2022 (N_2022,N_1864,N_1755);
or U2023 (N_2023,N_1994,N_1993);
xor U2024 (N_2024,N_1924,N_1874);
and U2025 (N_2025,N_1563,N_1770);
nor U2026 (N_2026,N_1995,N_1682);
xnor U2027 (N_2027,N_1857,N_1542);
and U2028 (N_2028,N_1579,N_1983);
xnor U2029 (N_2029,N_1711,N_1733);
nand U2030 (N_2030,N_1773,N_1788);
or U2031 (N_2031,N_1806,N_1974);
or U2032 (N_2032,N_1704,N_1735);
xor U2033 (N_2033,N_1501,N_1821);
and U2034 (N_2034,N_1966,N_1915);
nand U2035 (N_2035,N_1636,N_1932);
nand U2036 (N_2036,N_1572,N_1665);
xor U2037 (N_2037,N_1789,N_1771);
xnor U2038 (N_2038,N_1650,N_1908);
xor U2039 (N_2039,N_1914,N_1889);
and U2040 (N_2040,N_1548,N_1802);
or U2041 (N_2041,N_1555,N_1573);
xnor U2042 (N_2042,N_1996,N_1517);
or U2043 (N_2043,N_1622,N_1919);
nand U2044 (N_2044,N_1703,N_1911);
and U2045 (N_2045,N_1670,N_1599);
xor U2046 (N_2046,N_1524,N_1987);
xnor U2047 (N_2047,N_1764,N_1793);
or U2048 (N_2048,N_1598,N_1737);
or U2049 (N_2049,N_1964,N_1520);
nor U2050 (N_2050,N_1798,N_1586);
xor U2051 (N_2051,N_1991,N_1971);
or U2052 (N_2052,N_1955,N_1904);
nand U2053 (N_2053,N_1651,N_1766);
or U2054 (N_2054,N_1722,N_1849);
and U2055 (N_2055,N_1505,N_1847);
and U2056 (N_2056,N_1745,N_1982);
and U2057 (N_2057,N_1929,N_1967);
xnor U2058 (N_2058,N_1962,N_1736);
nor U2059 (N_2059,N_1829,N_1600);
or U2060 (N_2060,N_1634,N_1618);
nand U2061 (N_2061,N_1880,N_1783);
or U2062 (N_2062,N_1762,N_1851);
nor U2063 (N_2063,N_1881,N_1948);
xor U2064 (N_2064,N_1842,N_1615);
and U2065 (N_2065,N_1754,N_1696);
or U2066 (N_2066,N_1892,N_1920);
nand U2067 (N_2067,N_1805,N_1637);
xor U2068 (N_2068,N_1845,N_1702);
nand U2069 (N_2069,N_1561,N_1989);
xor U2070 (N_2070,N_1981,N_1684);
nor U2071 (N_2071,N_1585,N_1776);
xor U2072 (N_2072,N_1990,N_1641);
and U2073 (N_2073,N_1862,N_1679);
xnor U2074 (N_2074,N_1588,N_1593);
nand U2075 (N_2075,N_1873,N_1888);
nor U2076 (N_2076,N_1581,N_1811);
and U2077 (N_2077,N_1723,N_1640);
nand U2078 (N_2078,N_1950,N_1694);
nor U2079 (N_2079,N_1608,N_1595);
nand U2080 (N_2080,N_1965,N_1512);
xnor U2081 (N_2081,N_1706,N_1639);
nand U2082 (N_2082,N_1905,N_1786);
nand U2083 (N_2083,N_1659,N_1508);
xor U2084 (N_2084,N_1791,N_1539);
or U2085 (N_2085,N_1886,N_1601);
xnor U2086 (N_2086,N_1503,N_1726);
and U2087 (N_2087,N_1516,N_1537);
nor U2088 (N_2088,N_1638,N_1869);
or U2089 (N_2089,N_1787,N_1700);
xor U2090 (N_2090,N_1848,N_1610);
xor U2091 (N_2091,N_1819,N_1947);
and U2092 (N_2092,N_1833,N_1744);
xnor U2093 (N_2093,N_1533,N_1541);
or U2094 (N_2094,N_1937,N_1569);
nor U2095 (N_2095,N_1837,N_1836);
xnor U2096 (N_2096,N_1902,N_1685);
xnor U2097 (N_2097,N_1826,N_1866);
or U2098 (N_2098,N_1526,N_1532);
or U2099 (N_2099,N_1655,N_1898);
nand U2100 (N_2100,N_1676,N_1876);
or U2101 (N_2101,N_1681,N_1827);
nor U2102 (N_2102,N_1590,N_1560);
nor U2103 (N_2103,N_1589,N_1872);
xnor U2104 (N_2104,N_1810,N_1680);
or U2105 (N_2105,N_1832,N_1969);
nor U2106 (N_2106,N_1714,N_1976);
nor U2107 (N_2107,N_1576,N_1612);
or U2108 (N_2108,N_1739,N_1528);
nand U2109 (N_2109,N_1753,N_1758);
and U2110 (N_2110,N_1545,N_1642);
or U2111 (N_2111,N_1689,N_1627);
xor U2112 (N_2112,N_1671,N_1584);
and U2113 (N_2113,N_1717,N_1603);
and U2114 (N_2114,N_1580,N_1594);
xnor U2115 (N_2115,N_1777,N_1792);
nand U2116 (N_2116,N_1668,N_1648);
nand U2117 (N_2117,N_1839,N_1887);
and U2118 (N_2118,N_1534,N_1913);
nor U2119 (N_2119,N_1772,N_1831);
nor U2120 (N_2120,N_1878,N_1796);
nand U2121 (N_2121,N_1746,N_1975);
and U2122 (N_2122,N_1607,N_1575);
nor U2123 (N_2123,N_1557,N_1664);
or U2124 (N_2124,N_1592,N_1656);
nor U2125 (N_2125,N_1514,N_1906);
or U2126 (N_2126,N_1883,N_1630);
and U2127 (N_2127,N_1749,N_1815);
or U2128 (N_2128,N_1646,N_1551);
xnor U2129 (N_2129,N_1556,N_1934);
xor U2130 (N_2130,N_1999,N_1818);
and U2131 (N_2131,N_1631,N_1901);
or U2132 (N_2132,N_1823,N_1743);
or U2133 (N_2133,N_1732,N_1748);
xnor U2134 (N_2134,N_1624,N_1979);
or U2135 (N_2135,N_1562,N_1752);
xnor U2136 (N_2136,N_1657,N_1647);
xnor U2137 (N_2137,N_1946,N_1747);
and U2138 (N_2138,N_1769,N_1918);
or U2139 (N_2139,N_1797,N_1790);
and U2140 (N_2140,N_1817,N_1840);
or U2141 (N_2141,N_1910,N_1997);
xnor U2142 (N_2142,N_1527,N_1709);
and U2143 (N_2143,N_1960,N_1718);
xnor U2144 (N_2144,N_1943,N_1899);
nand U2145 (N_2145,N_1568,N_1985);
or U2146 (N_2146,N_1574,N_1500);
nand U2147 (N_2147,N_1540,N_1701);
nand U2148 (N_2148,N_1662,N_1956);
xor U2149 (N_2149,N_1725,N_1895);
xnor U2150 (N_2150,N_1807,N_1523);
and U2151 (N_2151,N_1850,N_1884);
xor U2152 (N_2152,N_1614,N_1785);
and U2153 (N_2153,N_1571,N_1644);
or U2154 (N_2154,N_1939,N_1677);
xnor U2155 (N_2155,N_1604,N_1801);
or U2156 (N_2156,N_1705,N_1536);
or U2157 (N_2157,N_1626,N_1544);
xnor U2158 (N_2158,N_1959,N_1928);
nand U2159 (N_2159,N_1757,N_1998);
or U2160 (N_2160,N_1896,N_1666);
nor U2161 (N_2161,N_1643,N_1549);
nor U2162 (N_2162,N_1820,N_1903);
and U2163 (N_2163,N_1550,N_1660);
and U2164 (N_2164,N_1519,N_1861);
xor U2165 (N_2165,N_1940,N_1721);
and U2166 (N_2166,N_1742,N_1830);
xnor U2167 (N_2167,N_1961,N_1727);
and U2168 (N_2168,N_1938,N_1708);
and U2169 (N_2169,N_1605,N_1779);
or U2170 (N_2170,N_1795,N_1724);
nand U2171 (N_2171,N_1564,N_1835);
nand U2172 (N_2172,N_1781,N_1782);
and U2173 (N_2173,N_1623,N_1907);
xor U2174 (N_2174,N_1633,N_1558);
xnor U2175 (N_2175,N_1768,N_1690);
xor U2176 (N_2176,N_1877,N_1868);
nand U2177 (N_2177,N_1844,N_1538);
and U2178 (N_2178,N_1578,N_1926);
or U2179 (N_2179,N_1582,N_1728);
nand U2180 (N_2180,N_1658,N_1688);
nand U2181 (N_2181,N_1531,N_1813);
nand U2182 (N_2182,N_1695,N_1778);
nor U2183 (N_2183,N_1865,N_1678);
nor U2184 (N_2184,N_1583,N_1577);
nand U2185 (N_2185,N_1611,N_1632);
or U2186 (N_2186,N_1522,N_1780);
nor U2187 (N_2187,N_1936,N_1653);
xor U2188 (N_2188,N_1713,N_1963);
nor U2189 (N_2189,N_1909,N_1751);
nand U2190 (N_2190,N_1860,N_1518);
nor U2191 (N_2191,N_1968,N_1834);
xor U2192 (N_2192,N_1565,N_1953);
nor U2193 (N_2193,N_1921,N_1654);
nand U2194 (N_2194,N_1794,N_1931);
or U2195 (N_2195,N_1803,N_1635);
xnor U2196 (N_2196,N_1756,N_1855);
and U2197 (N_2197,N_1730,N_1970);
nand U2198 (N_2198,N_1977,N_1699);
or U2199 (N_2199,N_1942,N_1502);
xor U2200 (N_2200,N_1716,N_1941);
nor U2201 (N_2201,N_1628,N_1570);
nor U2202 (N_2202,N_1957,N_1825);
xnor U2203 (N_2203,N_1854,N_1916);
and U2204 (N_2204,N_1693,N_1675);
or U2205 (N_2205,N_1897,N_1663);
nand U2206 (N_2206,N_1944,N_1828);
or U2207 (N_2207,N_1507,N_1973);
or U2208 (N_2208,N_1738,N_1838);
nor U2209 (N_2209,N_1691,N_1707);
and U2210 (N_2210,N_1692,N_1513);
nor U2211 (N_2211,N_1510,N_1649);
or U2212 (N_2212,N_1822,N_1816);
nor U2213 (N_2213,N_1774,N_1871);
nor U2214 (N_2214,N_1846,N_1852);
and U2215 (N_2215,N_1687,N_1890);
or U2216 (N_2216,N_1927,N_1992);
nand U2217 (N_2217,N_1697,N_1984);
and U2218 (N_2218,N_1933,N_1552);
xor U2219 (N_2219,N_1740,N_1613);
nor U2220 (N_2220,N_1645,N_1546);
nor U2221 (N_2221,N_1547,N_1683);
or U2222 (N_2222,N_1812,N_1800);
xor U2223 (N_2223,N_1606,N_1885);
or U2224 (N_2224,N_1814,N_1894);
nand U2225 (N_2225,N_1616,N_1530);
and U2226 (N_2226,N_1567,N_1761);
and U2227 (N_2227,N_1841,N_1525);
xor U2228 (N_2228,N_1554,N_1765);
nor U2229 (N_2229,N_1853,N_1710);
nor U2230 (N_2230,N_1750,N_1843);
xor U2231 (N_2231,N_1980,N_1978);
nor U2232 (N_2232,N_1958,N_1945);
or U2233 (N_2233,N_1617,N_1988);
nor U2234 (N_2234,N_1900,N_1652);
or U2235 (N_2235,N_1767,N_1859);
nand U2236 (N_2236,N_1824,N_1951);
or U2237 (N_2237,N_1972,N_1882);
and U2238 (N_2238,N_1621,N_1799);
xnor U2239 (N_2239,N_1784,N_1729);
xnor U2240 (N_2240,N_1858,N_1879);
and U2241 (N_2241,N_1760,N_1521);
nand U2242 (N_2242,N_1720,N_1511);
nor U2243 (N_2243,N_1715,N_1553);
xnor U2244 (N_2244,N_1596,N_1986);
nor U2245 (N_2245,N_1923,N_1667);
xnor U2246 (N_2246,N_1673,N_1602);
or U2247 (N_2247,N_1587,N_1863);
or U2248 (N_2248,N_1597,N_1922);
nor U2249 (N_2249,N_1515,N_1808);
nand U2250 (N_2250,N_1740,N_1631);
or U2251 (N_2251,N_1970,N_1718);
nor U2252 (N_2252,N_1824,N_1570);
and U2253 (N_2253,N_1839,N_1796);
nand U2254 (N_2254,N_1771,N_1932);
xnor U2255 (N_2255,N_1532,N_1651);
nand U2256 (N_2256,N_1894,N_1509);
nand U2257 (N_2257,N_1862,N_1703);
and U2258 (N_2258,N_1753,N_1657);
nor U2259 (N_2259,N_1700,N_1581);
or U2260 (N_2260,N_1689,N_1560);
nor U2261 (N_2261,N_1920,N_1758);
nor U2262 (N_2262,N_1793,N_1537);
and U2263 (N_2263,N_1778,N_1939);
nor U2264 (N_2264,N_1939,N_1625);
nand U2265 (N_2265,N_1616,N_1989);
nor U2266 (N_2266,N_1501,N_1845);
nor U2267 (N_2267,N_1997,N_1734);
and U2268 (N_2268,N_1552,N_1780);
xor U2269 (N_2269,N_1973,N_1783);
nor U2270 (N_2270,N_1722,N_1629);
or U2271 (N_2271,N_1628,N_1932);
or U2272 (N_2272,N_1687,N_1938);
or U2273 (N_2273,N_1704,N_1532);
or U2274 (N_2274,N_1737,N_1761);
and U2275 (N_2275,N_1760,N_1594);
nand U2276 (N_2276,N_1910,N_1907);
and U2277 (N_2277,N_1740,N_1753);
and U2278 (N_2278,N_1503,N_1677);
xor U2279 (N_2279,N_1583,N_1596);
nand U2280 (N_2280,N_1607,N_1719);
nand U2281 (N_2281,N_1813,N_1500);
xnor U2282 (N_2282,N_1763,N_1721);
and U2283 (N_2283,N_1575,N_1959);
nor U2284 (N_2284,N_1832,N_1841);
nand U2285 (N_2285,N_1946,N_1547);
xnor U2286 (N_2286,N_1810,N_1570);
nand U2287 (N_2287,N_1552,N_1653);
xnor U2288 (N_2288,N_1790,N_1650);
and U2289 (N_2289,N_1626,N_1976);
nand U2290 (N_2290,N_1897,N_1747);
xor U2291 (N_2291,N_1648,N_1831);
xnor U2292 (N_2292,N_1828,N_1527);
and U2293 (N_2293,N_1770,N_1633);
xnor U2294 (N_2294,N_1884,N_1762);
xnor U2295 (N_2295,N_1665,N_1960);
and U2296 (N_2296,N_1763,N_1896);
and U2297 (N_2297,N_1529,N_1965);
nand U2298 (N_2298,N_1588,N_1979);
nor U2299 (N_2299,N_1822,N_1931);
xor U2300 (N_2300,N_1610,N_1872);
and U2301 (N_2301,N_1653,N_1857);
xnor U2302 (N_2302,N_1647,N_1604);
xor U2303 (N_2303,N_1634,N_1748);
nor U2304 (N_2304,N_1920,N_1941);
nand U2305 (N_2305,N_1587,N_1948);
xnor U2306 (N_2306,N_1706,N_1773);
nor U2307 (N_2307,N_1887,N_1957);
nand U2308 (N_2308,N_1769,N_1723);
and U2309 (N_2309,N_1854,N_1717);
nor U2310 (N_2310,N_1754,N_1542);
nor U2311 (N_2311,N_1908,N_1681);
nand U2312 (N_2312,N_1804,N_1913);
or U2313 (N_2313,N_1678,N_1923);
or U2314 (N_2314,N_1682,N_1935);
nor U2315 (N_2315,N_1786,N_1838);
nor U2316 (N_2316,N_1920,N_1768);
and U2317 (N_2317,N_1789,N_1974);
or U2318 (N_2318,N_1803,N_1703);
xor U2319 (N_2319,N_1868,N_1594);
and U2320 (N_2320,N_1637,N_1731);
nand U2321 (N_2321,N_1734,N_1697);
or U2322 (N_2322,N_1529,N_1985);
nand U2323 (N_2323,N_1532,N_1571);
xor U2324 (N_2324,N_1648,N_1842);
nand U2325 (N_2325,N_1865,N_1975);
nor U2326 (N_2326,N_1608,N_1542);
nand U2327 (N_2327,N_1955,N_1514);
or U2328 (N_2328,N_1624,N_1622);
nor U2329 (N_2329,N_1798,N_1993);
xor U2330 (N_2330,N_1522,N_1955);
or U2331 (N_2331,N_1652,N_1669);
nor U2332 (N_2332,N_1929,N_1526);
nand U2333 (N_2333,N_1857,N_1641);
and U2334 (N_2334,N_1901,N_1772);
nand U2335 (N_2335,N_1537,N_1797);
and U2336 (N_2336,N_1819,N_1825);
or U2337 (N_2337,N_1526,N_1936);
nor U2338 (N_2338,N_1806,N_1970);
xor U2339 (N_2339,N_1808,N_1889);
nor U2340 (N_2340,N_1958,N_1746);
and U2341 (N_2341,N_1731,N_1971);
and U2342 (N_2342,N_1861,N_1691);
nor U2343 (N_2343,N_1874,N_1827);
nand U2344 (N_2344,N_1563,N_1554);
or U2345 (N_2345,N_1715,N_1718);
and U2346 (N_2346,N_1812,N_1550);
and U2347 (N_2347,N_1500,N_1612);
or U2348 (N_2348,N_1826,N_1882);
or U2349 (N_2349,N_1591,N_1623);
nand U2350 (N_2350,N_1506,N_1741);
or U2351 (N_2351,N_1612,N_1563);
and U2352 (N_2352,N_1585,N_1502);
and U2353 (N_2353,N_1937,N_1995);
nand U2354 (N_2354,N_1884,N_1521);
nand U2355 (N_2355,N_1739,N_1563);
xnor U2356 (N_2356,N_1802,N_1924);
nand U2357 (N_2357,N_1922,N_1810);
nand U2358 (N_2358,N_1960,N_1805);
nand U2359 (N_2359,N_1686,N_1721);
xor U2360 (N_2360,N_1715,N_1711);
xnor U2361 (N_2361,N_1507,N_1717);
or U2362 (N_2362,N_1529,N_1614);
xnor U2363 (N_2363,N_1959,N_1918);
nand U2364 (N_2364,N_1627,N_1847);
nand U2365 (N_2365,N_1590,N_1647);
and U2366 (N_2366,N_1622,N_1618);
and U2367 (N_2367,N_1865,N_1833);
and U2368 (N_2368,N_1670,N_1557);
xnor U2369 (N_2369,N_1794,N_1954);
and U2370 (N_2370,N_1974,N_1845);
nor U2371 (N_2371,N_1619,N_1932);
xor U2372 (N_2372,N_1532,N_1541);
nand U2373 (N_2373,N_1871,N_1864);
or U2374 (N_2374,N_1512,N_1889);
xnor U2375 (N_2375,N_1551,N_1830);
nor U2376 (N_2376,N_1720,N_1991);
xnor U2377 (N_2377,N_1788,N_1759);
and U2378 (N_2378,N_1641,N_1777);
nand U2379 (N_2379,N_1837,N_1921);
or U2380 (N_2380,N_1885,N_1585);
nor U2381 (N_2381,N_1897,N_1573);
nand U2382 (N_2382,N_1798,N_1904);
or U2383 (N_2383,N_1686,N_1860);
and U2384 (N_2384,N_1692,N_1709);
nand U2385 (N_2385,N_1865,N_1534);
nand U2386 (N_2386,N_1846,N_1697);
and U2387 (N_2387,N_1824,N_1697);
xor U2388 (N_2388,N_1822,N_1769);
xnor U2389 (N_2389,N_1657,N_1998);
xor U2390 (N_2390,N_1748,N_1534);
and U2391 (N_2391,N_1636,N_1808);
xnor U2392 (N_2392,N_1691,N_1695);
nor U2393 (N_2393,N_1794,N_1787);
and U2394 (N_2394,N_1892,N_1554);
xnor U2395 (N_2395,N_1561,N_1881);
xor U2396 (N_2396,N_1900,N_1927);
nand U2397 (N_2397,N_1675,N_1657);
xnor U2398 (N_2398,N_1917,N_1844);
xor U2399 (N_2399,N_1960,N_1954);
xnor U2400 (N_2400,N_1974,N_1818);
nor U2401 (N_2401,N_1665,N_1511);
nor U2402 (N_2402,N_1766,N_1852);
xnor U2403 (N_2403,N_1626,N_1556);
or U2404 (N_2404,N_1608,N_1731);
xnor U2405 (N_2405,N_1812,N_1752);
xnor U2406 (N_2406,N_1783,N_1526);
and U2407 (N_2407,N_1613,N_1992);
nor U2408 (N_2408,N_1728,N_1604);
and U2409 (N_2409,N_1847,N_1754);
xor U2410 (N_2410,N_1948,N_1798);
and U2411 (N_2411,N_1593,N_1660);
nand U2412 (N_2412,N_1962,N_1835);
nor U2413 (N_2413,N_1727,N_1929);
or U2414 (N_2414,N_1996,N_1721);
nor U2415 (N_2415,N_1642,N_1940);
nor U2416 (N_2416,N_1937,N_1988);
xor U2417 (N_2417,N_1543,N_1705);
and U2418 (N_2418,N_1771,N_1996);
nor U2419 (N_2419,N_1789,N_1871);
xnor U2420 (N_2420,N_1783,N_1649);
nor U2421 (N_2421,N_1592,N_1636);
xor U2422 (N_2422,N_1846,N_1937);
nand U2423 (N_2423,N_1775,N_1742);
nand U2424 (N_2424,N_1553,N_1787);
xor U2425 (N_2425,N_1797,N_1996);
or U2426 (N_2426,N_1545,N_1584);
and U2427 (N_2427,N_1724,N_1904);
nand U2428 (N_2428,N_1925,N_1534);
nand U2429 (N_2429,N_1603,N_1799);
or U2430 (N_2430,N_1955,N_1693);
nand U2431 (N_2431,N_1767,N_1938);
nand U2432 (N_2432,N_1826,N_1601);
nand U2433 (N_2433,N_1542,N_1578);
nor U2434 (N_2434,N_1692,N_1586);
or U2435 (N_2435,N_1551,N_1794);
xor U2436 (N_2436,N_1651,N_1751);
or U2437 (N_2437,N_1828,N_1923);
nand U2438 (N_2438,N_1701,N_1862);
or U2439 (N_2439,N_1721,N_1523);
nand U2440 (N_2440,N_1828,N_1744);
nor U2441 (N_2441,N_1883,N_1757);
and U2442 (N_2442,N_1657,N_1799);
xnor U2443 (N_2443,N_1753,N_1782);
nand U2444 (N_2444,N_1546,N_1738);
xnor U2445 (N_2445,N_1614,N_1887);
nor U2446 (N_2446,N_1879,N_1562);
nand U2447 (N_2447,N_1722,N_1976);
nand U2448 (N_2448,N_1770,N_1528);
xnor U2449 (N_2449,N_1793,N_1971);
xnor U2450 (N_2450,N_1710,N_1824);
xor U2451 (N_2451,N_1740,N_1950);
nand U2452 (N_2452,N_1593,N_1861);
nor U2453 (N_2453,N_1911,N_1522);
nand U2454 (N_2454,N_1846,N_1968);
nor U2455 (N_2455,N_1600,N_1720);
or U2456 (N_2456,N_1769,N_1895);
nor U2457 (N_2457,N_1779,N_1910);
or U2458 (N_2458,N_1672,N_1957);
nor U2459 (N_2459,N_1905,N_1813);
nand U2460 (N_2460,N_1651,N_1739);
xor U2461 (N_2461,N_1539,N_1559);
xor U2462 (N_2462,N_1504,N_1507);
xnor U2463 (N_2463,N_1930,N_1750);
nor U2464 (N_2464,N_1856,N_1594);
xnor U2465 (N_2465,N_1757,N_1944);
or U2466 (N_2466,N_1799,N_1848);
nor U2467 (N_2467,N_1998,N_1670);
nor U2468 (N_2468,N_1570,N_1569);
nor U2469 (N_2469,N_1546,N_1821);
and U2470 (N_2470,N_1871,N_1867);
nand U2471 (N_2471,N_1714,N_1530);
nor U2472 (N_2472,N_1753,N_1815);
nand U2473 (N_2473,N_1650,N_1688);
xnor U2474 (N_2474,N_1505,N_1985);
or U2475 (N_2475,N_1894,N_1798);
and U2476 (N_2476,N_1633,N_1590);
and U2477 (N_2477,N_1959,N_1962);
xor U2478 (N_2478,N_1616,N_1979);
nor U2479 (N_2479,N_1659,N_1585);
and U2480 (N_2480,N_1960,N_1783);
or U2481 (N_2481,N_1811,N_1630);
xnor U2482 (N_2482,N_1861,N_1797);
nand U2483 (N_2483,N_1800,N_1755);
nor U2484 (N_2484,N_1708,N_1906);
and U2485 (N_2485,N_1547,N_1588);
xor U2486 (N_2486,N_1713,N_1604);
and U2487 (N_2487,N_1633,N_1584);
and U2488 (N_2488,N_1858,N_1784);
and U2489 (N_2489,N_1627,N_1706);
and U2490 (N_2490,N_1821,N_1773);
nor U2491 (N_2491,N_1643,N_1590);
and U2492 (N_2492,N_1598,N_1896);
nand U2493 (N_2493,N_1907,N_1758);
xor U2494 (N_2494,N_1849,N_1504);
and U2495 (N_2495,N_1618,N_1582);
nor U2496 (N_2496,N_1528,N_1714);
nor U2497 (N_2497,N_1586,N_1739);
xor U2498 (N_2498,N_1871,N_1685);
nand U2499 (N_2499,N_1738,N_1573);
nand U2500 (N_2500,N_2371,N_2472);
nor U2501 (N_2501,N_2110,N_2437);
nor U2502 (N_2502,N_2406,N_2132);
xor U2503 (N_2503,N_2191,N_2359);
nand U2504 (N_2504,N_2459,N_2360);
xnor U2505 (N_2505,N_2423,N_2023);
nor U2506 (N_2506,N_2282,N_2452);
or U2507 (N_2507,N_2442,N_2245);
xor U2508 (N_2508,N_2238,N_2131);
nand U2509 (N_2509,N_2012,N_2017);
and U2510 (N_2510,N_2106,N_2060);
or U2511 (N_2511,N_2397,N_2021);
and U2512 (N_2512,N_2408,N_2253);
xor U2513 (N_2513,N_2281,N_2162);
xor U2514 (N_2514,N_2388,N_2016);
nand U2515 (N_2515,N_2159,N_2204);
nand U2516 (N_2516,N_2321,N_2476);
nor U2517 (N_2517,N_2052,N_2010);
and U2518 (N_2518,N_2491,N_2414);
nor U2519 (N_2519,N_2415,N_2305);
xor U2520 (N_2520,N_2381,N_2148);
or U2521 (N_2521,N_2498,N_2308);
and U2522 (N_2522,N_2180,N_2461);
xor U2523 (N_2523,N_2424,N_2404);
xnor U2524 (N_2524,N_2128,N_2145);
and U2525 (N_2525,N_2441,N_2272);
xnor U2526 (N_2526,N_2002,N_2140);
nand U2527 (N_2527,N_2050,N_2146);
nor U2528 (N_2528,N_2113,N_2264);
nor U2529 (N_2529,N_2174,N_2008);
xnor U2530 (N_2530,N_2446,N_2109);
nand U2531 (N_2531,N_2161,N_2116);
and U2532 (N_2532,N_2209,N_2088);
nand U2533 (N_2533,N_2107,N_2073);
nor U2534 (N_2534,N_2483,N_2463);
nor U2535 (N_2535,N_2158,N_2470);
or U2536 (N_2536,N_2176,N_2197);
nand U2537 (N_2537,N_2320,N_2056);
nor U2538 (N_2538,N_2066,N_2494);
or U2539 (N_2539,N_2306,N_2293);
and U2540 (N_2540,N_2297,N_2436);
xor U2541 (N_2541,N_2172,N_2059);
nor U2542 (N_2542,N_2137,N_2339);
or U2543 (N_2543,N_2098,N_2227);
nor U2544 (N_2544,N_2150,N_2263);
and U2545 (N_2545,N_2244,N_2118);
and U2546 (N_2546,N_2211,N_2228);
or U2547 (N_2547,N_2215,N_2223);
and U2548 (N_2548,N_2327,N_2328);
or U2549 (N_2549,N_2280,N_2235);
nand U2550 (N_2550,N_2286,N_2045);
nor U2551 (N_2551,N_2468,N_2323);
nor U2552 (N_2552,N_2011,N_2481);
xor U2553 (N_2553,N_2038,N_2487);
nand U2554 (N_2554,N_2034,N_2234);
xor U2555 (N_2555,N_2399,N_2333);
nand U2556 (N_2556,N_2499,N_2094);
xor U2557 (N_2557,N_2347,N_2037);
nand U2558 (N_2558,N_2004,N_2267);
xnor U2559 (N_2559,N_2389,N_2425);
xor U2560 (N_2560,N_2292,N_2385);
nor U2561 (N_2561,N_2458,N_2496);
xnor U2562 (N_2562,N_2111,N_2495);
xnor U2563 (N_2563,N_2091,N_2251);
xor U2564 (N_2564,N_2341,N_2394);
nor U2565 (N_2565,N_2236,N_2299);
xor U2566 (N_2566,N_2455,N_2284);
nand U2567 (N_2567,N_2497,N_2075);
nor U2568 (N_2568,N_2257,N_2068);
and U2569 (N_2569,N_2265,N_2322);
or U2570 (N_2570,N_2212,N_2445);
xnor U2571 (N_2571,N_2310,N_2188);
nor U2572 (N_2572,N_2474,N_2230);
and U2573 (N_2573,N_2307,N_2022);
xnor U2574 (N_2574,N_2168,N_2380);
xor U2575 (N_2575,N_2478,N_2165);
or U2576 (N_2576,N_2271,N_2024);
nor U2577 (N_2577,N_2312,N_2342);
xnor U2578 (N_2578,N_2001,N_2489);
and U2579 (N_2579,N_2029,N_2040);
and U2580 (N_2580,N_2170,N_2260);
xnor U2581 (N_2581,N_2413,N_2213);
nand U2582 (N_2582,N_2490,N_2199);
or U2583 (N_2583,N_2203,N_2138);
or U2584 (N_2584,N_2332,N_2324);
xor U2585 (N_2585,N_2080,N_2447);
nand U2586 (N_2586,N_2258,N_2384);
or U2587 (N_2587,N_2355,N_2096);
nor U2588 (N_2588,N_2007,N_2421);
or U2589 (N_2589,N_2041,N_2229);
xnor U2590 (N_2590,N_2104,N_2061);
nor U2591 (N_2591,N_2195,N_2467);
or U2592 (N_2592,N_2396,N_2157);
nor U2593 (N_2593,N_2405,N_2175);
xor U2594 (N_2594,N_2039,N_2124);
xnor U2595 (N_2595,N_2015,N_2062);
and U2596 (N_2596,N_2337,N_2390);
xor U2597 (N_2597,N_2419,N_2454);
and U2598 (N_2598,N_2147,N_2363);
nor U2599 (N_2599,N_2285,N_2208);
nand U2600 (N_2600,N_2361,N_2407);
or U2601 (N_2601,N_2439,N_2484);
or U2602 (N_2602,N_2448,N_2125);
nor U2603 (N_2603,N_2063,N_2471);
and U2604 (N_2604,N_2298,N_2398);
and U2605 (N_2605,N_2351,N_2087);
or U2606 (N_2606,N_2274,N_2067);
nand U2607 (N_2607,N_2089,N_2090);
nor U2608 (N_2608,N_2336,N_2185);
nand U2609 (N_2609,N_2451,N_2231);
or U2610 (N_2610,N_2233,N_2444);
and U2611 (N_2611,N_2289,N_2279);
xor U2612 (N_2612,N_2036,N_2477);
nor U2613 (N_2613,N_2095,N_2329);
nand U2614 (N_2614,N_2400,N_2275);
nor U2615 (N_2615,N_2206,N_2373);
xor U2616 (N_2616,N_2026,N_2276);
and U2617 (N_2617,N_2278,N_2457);
or U2618 (N_2618,N_2144,N_2134);
and U2619 (N_2619,N_2420,N_2009);
nand U2620 (N_2620,N_2184,N_2469);
xnor U2621 (N_2621,N_2325,N_2435);
and U2622 (N_2622,N_2316,N_2013);
xnor U2623 (N_2623,N_2123,N_2261);
and U2624 (N_2624,N_2345,N_2177);
and U2625 (N_2625,N_2295,N_2377);
xor U2626 (N_2626,N_2338,N_2365);
xnor U2627 (N_2627,N_2099,N_2273);
and U2628 (N_2628,N_2256,N_2205);
or U2629 (N_2629,N_2376,N_2250);
nand U2630 (N_2630,N_2422,N_2084);
or U2631 (N_2631,N_2243,N_2375);
and U2632 (N_2632,N_2102,N_2129);
and U2633 (N_2633,N_2190,N_2222);
xor U2634 (N_2634,N_2402,N_2353);
and U2635 (N_2635,N_2178,N_2220);
and U2636 (N_2636,N_2051,N_2302);
nand U2637 (N_2637,N_2058,N_2464);
and U2638 (N_2638,N_2268,N_2319);
xor U2639 (N_2639,N_2440,N_2462);
or U2640 (N_2640,N_2315,N_2081);
or U2641 (N_2641,N_2028,N_2014);
or U2642 (N_2642,N_2167,N_2006);
xor U2643 (N_2643,N_2266,N_2072);
xnor U2644 (N_2644,N_2382,N_2126);
nand U2645 (N_2645,N_2317,N_2169);
nor U2646 (N_2646,N_2386,N_2097);
xor U2647 (N_2647,N_2114,N_2300);
and U2648 (N_2648,N_2369,N_2427);
nand U2649 (N_2649,N_2112,N_2183);
xnor U2650 (N_2650,N_2093,N_2149);
nor U2651 (N_2651,N_2348,N_2370);
nand U2652 (N_2652,N_2069,N_2249);
and U2653 (N_2653,N_2432,N_2456);
xor U2654 (N_2654,N_2493,N_2117);
xnor U2655 (N_2655,N_2433,N_2240);
nor U2656 (N_2656,N_2130,N_2387);
or U2657 (N_2657,N_2076,N_2255);
or U2658 (N_2658,N_2179,N_2460);
or U2659 (N_2659,N_2480,N_2374);
nor U2660 (N_2660,N_2296,N_2163);
and U2661 (N_2661,N_2127,N_2226);
and U2662 (N_2662,N_2003,N_2173);
or U2663 (N_2663,N_2120,N_2330);
nor U2664 (N_2664,N_2473,N_2005);
and U2665 (N_2665,N_2194,N_2290);
or U2666 (N_2666,N_2362,N_2350);
and U2667 (N_2667,N_2262,N_2311);
nand U2668 (N_2668,N_2103,N_2486);
nor U2669 (N_2669,N_2378,N_2364);
nand U2670 (N_2670,N_2270,N_2071);
and U2671 (N_2671,N_2343,N_2152);
nand U2672 (N_2672,N_2313,N_2239);
nand U2673 (N_2673,N_2426,N_2367);
xor U2674 (N_2674,N_2142,N_2242);
xor U2675 (N_2675,N_2078,N_2492);
and U2676 (N_2676,N_2434,N_2331);
nor U2677 (N_2677,N_2122,N_2277);
nand U2678 (N_2678,N_2181,N_2064);
or U2679 (N_2679,N_2032,N_2189);
xor U2680 (N_2680,N_2200,N_2100);
nor U2681 (N_2681,N_2115,N_2366);
xor U2682 (N_2682,N_2031,N_2418);
nand U2683 (N_2683,N_2417,N_2340);
and U2684 (N_2684,N_2309,N_2135);
nor U2685 (N_2685,N_2372,N_2475);
and U2686 (N_2686,N_2139,N_2065);
nor U2687 (N_2687,N_2287,N_2030);
and U2688 (N_2688,N_2141,N_2153);
or U2689 (N_2689,N_2196,N_2193);
and U2690 (N_2690,N_2049,N_2121);
xor U2691 (N_2691,N_2237,N_2086);
nand U2692 (N_2692,N_2054,N_2335);
xnor U2693 (N_2693,N_2438,N_2154);
nor U2694 (N_2694,N_2465,N_2395);
or U2695 (N_2695,N_2042,N_2379);
nor U2696 (N_2696,N_2416,N_2217);
nand U2697 (N_2697,N_2357,N_2354);
or U2698 (N_2698,N_2079,N_2187);
or U2699 (N_2699,N_2083,N_2254);
or U2700 (N_2700,N_2352,N_2232);
nand U2701 (N_2701,N_2428,N_2156);
and U2702 (N_2702,N_2085,N_2027);
nor U2703 (N_2703,N_2207,N_2344);
nor U2704 (N_2704,N_2186,N_2247);
and U2705 (N_2705,N_2025,N_2000);
xor U2706 (N_2706,N_2119,N_2403);
and U2707 (N_2707,N_2092,N_2057);
or U2708 (N_2708,N_2252,N_2151);
nor U2709 (N_2709,N_2401,N_2383);
nand U2710 (N_2710,N_2346,N_2166);
xor U2711 (N_2711,N_2449,N_2409);
xnor U2712 (N_2712,N_2070,N_2019);
nand U2713 (N_2713,N_2259,N_2288);
nor U2714 (N_2714,N_2283,N_2466);
nor U2715 (N_2715,N_2431,N_2301);
or U2716 (N_2716,N_2160,N_2044);
nand U2717 (N_2717,N_2074,N_2429);
xor U2718 (N_2718,N_2430,N_2485);
xnor U2719 (N_2719,N_2241,N_2368);
nor U2720 (N_2720,N_2210,N_2294);
or U2721 (N_2721,N_2246,N_2055);
nor U2722 (N_2722,N_2047,N_2269);
xor U2723 (N_2723,N_2488,N_2077);
and U2724 (N_2724,N_2479,N_2410);
xnor U2725 (N_2725,N_2219,N_2216);
nor U2726 (N_2726,N_2326,N_2198);
nor U2727 (N_2727,N_2101,N_2391);
and U2728 (N_2728,N_2043,N_2453);
and U2729 (N_2729,N_2171,N_2318);
or U2730 (N_2730,N_2221,N_2133);
nor U2731 (N_2731,N_2482,N_2443);
xnor U2732 (N_2732,N_2349,N_2411);
nor U2733 (N_2733,N_2164,N_2450);
xor U2734 (N_2734,N_2224,N_2392);
xnor U2735 (N_2735,N_2201,N_2393);
and U2736 (N_2736,N_2020,N_2018);
nor U2737 (N_2737,N_2356,N_2053);
nand U2738 (N_2738,N_2304,N_2218);
nand U2739 (N_2739,N_2248,N_2082);
xnor U2740 (N_2740,N_2314,N_2035);
xnor U2741 (N_2741,N_2303,N_2143);
nor U2742 (N_2742,N_2046,N_2291);
or U2743 (N_2743,N_2225,N_2334);
and U2744 (N_2744,N_2033,N_2155);
or U2745 (N_2745,N_2048,N_2192);
or U2746 (N_2746,N_2182,N_2202);
or U2747 (N_2747,N_2136,N_2105);
or U2748 (N_2748,N_2358,N_2214);
xor U2749 (N_2749,N_2412,N_2108);
or U2750 (N_2750,N_2046,N_2197);
xnor U2751 (N_2751,N_2120,N_2147);
and U2752 (N_2752,N_2147,N_2005);
and U2753 (N_2753,N_2112,N_2009);
and U2754 (N_2754,N_2342,N_2058);
nand U2755 (N_2755,N_2356,N_2076);
xor U2756 (N_2756,N_2399,N_2090);
and U2757 (N_2757,N_2063,N_2358);
or U2758 (N_2758,N_2410,N_2027);
nor U2759 (N_2759,N_2362,N_2179);
nor U2760 (N_2760,N_2111,N_2060);
and U2761 (N_2761,N_2488,N_2311);
nand U2762 (N_2762,N_2483,N_2077);
xor U2763 (N_2763,N_2254,N_2414);
and U2764 (N_2764,N_2087,N_2206);
or U2765 (N_2765,N_2256,N_2411);
nor U2766 (N_2766,N_2401,N_2134);
nor U2767 (N_2767,N_2255,N_2169);
nor U2768 (N_2768,N_2009,N_2036);
xnor U2769 (N_2769,N_2166,N_2039);
and U2770 (N_2770,N_2225,N_2023);
nor U2771 (N_2771,N_2141,N_2064);
xor U2772 (N_2772,N_2056,N_2310);
nor U2773 (N_2773,N_2388,N_2159);
nor U2774 (N_2774,N_2033,N_2166);
nand U2775 (N_2775,N_2483,N_2301);
nor U2776 (N_2776,N_2143,N_2287);
xor U2777 (N_2777,N_2257,N_2284);
nor U2778 (N_2778,N_2138,N_2188);
nor U2779 (N_2779,N_2147,N_2433);
or U2780 (N_2780,N_2012,N_2196);
nand U2781 (N_2781,N_2407,N_2323);
nor U2782 (N_2782,N_2252,N_2050);
or U2783 (N_2783,N_2265,N_2445);
nor U2784 (N_2784,N_2324,N_2010);
nand U2785 (N_2785,N_2213,N_2390);
nor U2786 (N_2786,N_2183,N_2159);
nor U2787 (N_2787,N_2093,N_2080);
nand U2788 (N_2788,N_2459,N_2406);
nor U2789 (N_2789,N_2369,N_2164);
nand U2790 (N_2790,N_2467,N_2481);
nand U2791 (N_2791,N_2167,N_2269);
nor U2792 (N_2792,N_2456,N_2392);
nor U2793 (N_2793,N_2221,N_2247);
nor U2794 (N_2794,N_2032,N_2350);
and U2795 (N_2795,N_2016,N_2306);
and U2796 (N_2796,N_2028,N_2440);
xor U2797 (N_2797,N_2265,N_2465);
and U2798 (N_2798,N_2153,N_2447);
or U2799 (N_2799,N_2440,N_2053);
xor U2800 (N_2800,N_2096,N_2372);
nor U2801 (N_2801,N_2369,N_2321);
xnor U2802 (N_2802,N_2192,N_2181);
xnor U2803 (N_2803,N_2465,N_2176);
xor U2804 (N_2804,N_2419,N_2184);
nand U2805 (N_2805,N_2483,N_2281);
nand U2806 (N_2806,N_2101,N_2354);
xor U2807 (N_2807,N_2419,N_2138);
nor U2808 (N_2808,N_2291,N_2078);
xnor U2809 (N_2809,N_2064,N_2026);
and U2810 (N_2810,N_2254,N_2210);
nor U2811 (N_2811,N_2411,N_2113);
nand U2812 (N_2812,N_2326,N_2376);
nand U2813 (N_2813,N_2348,N_2232);
xnor U2814 (N_2814,N_2221,N_2406);
xnor U2815 (N_2815,N_2240,N_2377);
xnor U2816 (N_2816,N_2379,N_2426);
nand U2817 (N_2817,N_2049,N_2052);
and U2818 (N_2818,N_2254,N_2481);
nor U2819 (N_2819,N_2181,N_2044);
nand U2820 (N_2820,N_2257,N_2208);
nor U2821 (N_2821,N_2193,N_2413);
or U2822 (N_2822,N_2251,N_2354);
xor U2823 (N_2823,N_2185,N_2241);
nor U2824 (N_2824,N_2303,N_2497);
or U2825 (N_2825,N_2315,N_2209);
or U2826 (N_2826,N_2129,N_2131);
xor U2827 (N_2827,N_2330,N_2336);
nor U2828 (N_2828,N_2008,N_2424);
or U2829 (N_2829,N_2110,N_2150);
or U2830 (N_2830,N_2078,N_2489);
nand U2831 (N_2831,N_2259,N_2462);
nor U2832 (N_2832,N_2154,N_2138);
nand U2833 (N_2833,N_2159,N_2218);
nor U2834 (N_2834,N_2381,N_2229);
or U2835 (N_2835,N_2383,N_2476);
nand U2836 (N_2836,N_2273,N_2171);
or U2837 (N_2837,N_2194,N_2122);
xnor U2838 (N_2838,N_2222,N_2279);
and U2839 (N_2839,N_2081,N_2172);
xnor U2840 (N_2840,N_2475,N_2330);
nor U2841 (N_2841,N_2452,N_2124);
nor U2842 (N_2842,N_2211,N_2199);
nor U2843 (N_2843,N_2177,N_2235);
xnor U2844 (N_2844,N_2134,N_2438);
or U2845 (N_2845,N_2496,N_2003);
or U2846 (N_2846,N_2079,N_2337);
xnor U2847 (N_2847,N_2214,N_2275);
and U2848 (N_2848,N_2359,N_2362);
and U2849 (N_2849,N_2434,N_2147);
xor U2850 (N_2850,N_2186,N_2385);
xnor U2851 (N_2851,N_2005,N_2048);
and U2852 (N_2852,N_2499,N_2163);
nor U2853 (N_2853,N_2303,N_2245);
and U2854 (N_2854,N_2251,N_2246);
and U2855 (N_2855,N_2221,N_2279);
or U2856 (N_2856,N_2418,N_2181);
nand U2857 (N_2857,N_2239,N_2067);
and U2858 (N_2858,N_2027,N_2420);
nor U2859 (N_2859,N_2495,N_2409);
xnor U2860 (N_2860,N_2265,N_2250);
xor U2861 (N_2861,N_2139,N_2041);
nand U2862 (N_2862,N_2408,N_2212);
nor U2863 (N_2863,N_2434,N_2100);
xor U2864 (N_2864,N_2448,N_2300);
nand U2865 (N_2865,N_2490,N_2016);
xnor U2866 (N_2866,N_2498,N_2030);
nor U2867 (N_2867,N_2485,N_2346);
nand U2868 (N_2868,N_2207,N_2185);
nor U2869 (N_2869,N_2453,N_2279);
nand U2870 (N_2870,N_2462,N_2041);
nand U2871 (N_2871,N_2448,N_2227);
or U2872 (N_2872,N_2443,N_2158);
and U2873 (N_2873,N_2088,N_2153);
and U2874 (N_2874,N_2453,N_2187);
and U2875 (N_2875,N_2333,N_2227);
nor U2876 (N_2876,N_2451,N_2371);
or U2877 (N_2877,N_2136,N_2293);
xor U2878 (N_2878,N_2149,N_2176);
and U2879 (N_2879,N_2253,N_2456);
xnor U2880 (N_2880,N_2476,N_2296);
nor U2881 (N_2881,N_2046,N_2303);
and U2882 (N_2882,N_2229,N_2117);
xor U2883 (N_2883,N_2060,N_2247);
nor U2884 (N_2884,N_2411,N_2390);
or U2885 (N_2885,N_2057,N_2098);
and U2886 (N_2886,N_2192,N_2089);
xnor U2887 (N_2887,N_2321,N_2426);
nor U2888 (N_2888,N_2102,N_2278);
and U2889 (N_2889,N_2112,N_2289);
and U2890 (N_2890,N_2413,N_2076);
xnor U2891 (N_2891,N_2051,N_2430);
xnor U2892 (N_2892,N_2437,N_2299);
nor U2893 (N_2893,N_2293,N_2078);
nor U2894 (N_2894,N_2169,N_2360);
and U2895 (N_2895,N_2292,N_2137);
xnor U2896 (N_2896,N_2430,N_2464);
or U2897 (N_2897,N_2337,N_2055);
and U2898 (N_2898,N_2178,N_2020);
nor U2899 (N_2899,N_2387,N_2378);
xor U2900 (N_2900,N_2477,N_2251);
xor U2901 (N_2901,N_2042,N_2436);
or U2902 (N_2902,N_2159,N_2279);
nand U2903 (N_2903,N_2309,N_2214);
xor U2904 (N_2904,N_2284,N_2380);
nor U2905 (N_2905,N_2255,N_2139);
and U2906 (N_2906,N_2071,N_2420);
xor U2907 (N_2907,N_2467,N_2182);
xor U2908 (N_2908,N_2256,N_2366);
xor U2909 (N_2909,N_2141,N_2259);
and U2910 (N_2910,N_2315,N_2326);
nor U2911 (N_2911,N_2378,N_2049);
or U2912 (N_2912,N_2122,N_2360);
or U2913 (N_2913,N_2331,N_2411);
xnor U2914 (N_2914,N_2297,N_2276);
or U2915 (N_2915,N_2113,N_2167);
nand U2916 (N_2916,N_2065,N_2328);
nor U2917 (N_2917,N_2213,N_2342);
or U2918 (N_2918,N_2425,N_2483);
and U2919 (N_2919,N_2373,N_2473);
and U2920 (N_2920,N_2068,N_2046);
or U2921 (N_2921,N_2218,N_2341);
nand U2922 (N_2922,N_2451,N_2094);
and U2923 (N_2923,N_2031,N_2034);
and U2924 (N_2924,N_2341,N_2372);
nor U2925 (N_2925,N_2000,N_2303);
xor U2926 (N_2926,N_2242,N_2455);
nor U2927 (N_2927,N_2365,N_2072);
and U2928 (N_2928,N_2000,N_2150);
xnor U2929 (N_2929,N_2359,N_2451);
xnor U2930 (N_2930,N_2168,N_2253);
nand U2931 (N_2931,N_2494,N_2146);
and U2932 (N_2932,N_2179,N_2395);
and U2933 (N_2933,N_2003,N_2167);
xor U2934 (N_2934,N_2305,N_2022);
or U2935 (N_2935,N_2439,N_2022);
xnor U2936 (N_2936,N_2066,N_2419);
or U2937 (N_2937,N_2366,N_2069);
nor U2938 (N_2938,N_2333,N_2113);
nor U2939 (N_2939,N_2454,N_2382);
or U2940 (N_2940,N_2179,N_2064);
and U2941 (N_2941,N_2400,N_2194);
or U2942 (N_2942,N_2051,N_2410);
nor U2943 (N_2943,N_2323,N_2493);
xnor U2944 (N_2944,N_2373,N_2472);
nor U2945 (N_2945,N_2031,N_2276);
nand U2946 (N_2946,N_2131,N_2470);
nand U2947 (N_2947,N_2409,N_2446);
or U2948 (N_2948,N_2312,N_2253);
xor U2949 (N_2949,N_2081,N_2023);
xnor U2950 (N_2950,N_2078,N_2026);
or U2951 (N_2951,N_2327,N_2283);
xnor U2952 (N_2952,N_2227,N_2492);
nor U2953 (N_2953,N_2087,N_2235);
nor U2954 (N_2954,N_2029,N_2368);
and U2955 (N_2955,N_2003,N_2227);
or U2956 (N_2956,N_2085,N_2005);
and U2957 (N_2957,N_2108,N_2006);
nor U2958 (N_2958,N_2037,N_2493);
nand U2959 (N_2959,N_2290,N_2473);
nand U2960 (N_2960,N_2093,N_2377);
nor U2961 (N_2961,N_2454,N_2135);
or U2962 (N_2962,N_2236,N_2386);
or U2963 (N_2963,N_2190,N_2278);
and U2964 (N_2964,N_2420,N_2316);
nor U2965 (N_2965,N_2004,N_2455);
nand U2966 (N_2966,N_2391,N_2027);
nand U2967 (N_2967,N_2098,N_2082);
or U2968 (N_2968,N_2016,N_2223);
nand U2969 (N_2969,N_2372,N_2477);
or U2970 (N_2970,N_2354,N_2371);
nor U2971 (N_2971,N_2404,N_2055);
xnor U2972 (N_2972,N_2267,N_2447);
and U2973 (N_2973,N_2468,N_2321);
nand U2974 (N_2974,N_2255,N_2153);
nand U2975 (N_2975,N_2128,N_2107);
or U2976 (N_2976,N_2009,N_2309);
or U2977 (N_2977,N_2079,N_2111);
nor U2978 (N_2978,N_2103,N_2407);
and U2979 (N_2979,N_2031,N_2409);
nand U2980 (N_2980,N_2156,N_2303);
xor U2981 (N_2981,N_2040,N_2225);
nor U2982 (N_2982,N_2286,N_2122);
or U2983 (N_2983,N_2339,N_2095);
and U2984 (N_2984,N_2165,N_2103);
nand U2985 (N_2985,N_2181,N_2052);
and U2986 (N_2986,N_2424,N_2167);
xnor U2987 (N_2987,N_2242,N_2399);
nor U2988 (N_2988,N_2240,N_2272);
or U2989 (N_2989,N_2329,N_2029);
and U2990 (N_2990,N_2015,N_2048);
xnor U2991 (N_2991,N_2047,N_2114);
nor U2992 (N_2992,N_2164,N_2176);
nor U2993 (N_2993,N_2238,N_2249);
xnor U2994 (N_2994,N_2176,N_2367);
or U2995 (N_2995,N_2109,N_2110);
or U2996 (N_2996,N_2448,N_2179);
or U2997 (N_2997,N_2397,N_2488);
nand U2998 (N_2998,N_2138,N_2351);
and U2999 (N_2999,N_2401,N_2320);
xnor UO_0 (O_0,N_2840,N_2847);
nand UO_1 (O_1,N_2773,N_2671);
or UO_2 (O_2,N_2538,N_2843);
xnor UO_3 (O_3,N_2756,N_2804);
and UO_4 (O_4,N_2883,N_2642);
nor UO_5 (O_5,N_2566,N_2586);
nor UO_6 (O_6,N_2984,N_2914);
and UO_7 (O_7,N_2946,N_2514);
nand UO_8 (O_8,N_2599,N_2604);
and UO_9 (O_9,N_2725,N_2881);
nor UO_10 (O_10,N_2697,N_2991);
and UO_11 (O_11,N_2698,N_2995);
and UO_12 (O_12,N_2973,N_2859);
xnor UO_13 (O_13,N_2627,N_2791);
or UO_14 (O_14,N_2659,N_2755);
xor UO_15 (O_15,N_2633,N_2649);
nand UO_16 (O_16,N_2759,N_2987);
or UO_17 (O_17,N_2726,N_2715);
xnor UO_18 (O_18,N_2714,N_2570);
nand UO_19 (O_19,N_2529,N_2929);
nor UO_20 (O_20,N_2508,N_2636);
and UO_21 (O_21,N_2862,N_2864);
or UO_22 (O_22,N_2788,N_2970);
and UO_23 (O_23,N_2936,N_2863);
and UO_24 (O_24,N_2886,N_2763);
or UO_25 (O_25,N_2744,N_2823);
xor UO_26 (O_26,N_2792,N_2776);
and UO_27 (O_27,N_2975,N_2727);
or UO_28 (O_28,N_2805,N_2800);
and UO_29 (O_29,N_2880,N_2923);
nand UO_30 (O_30,N_2562,N_2907);
xor UO_31 (O_31,N_2783,N_2898);
or UO_32 (O_32,N_2739,N_2640);
nand UO_33 (O_33,N_2913,N_2996);
and UO_34 (O_34,N_2748,N_2705);
or UO_35 (O_35,N_2510,N_2769);
nand UO_36 (O_36,N_2962,N_2968);
nand UO_37 (O_37,N_2612,N_2850);
and UO_38 (O_38,N_2641,N_2741);
or UO_39 (O_39,N_2596,N_2543);
nand UO_40 (O_40,N_2650,N_2573);
or UO_41 (O_41,N_2515,N_2990);
and UO_42 (O_42,N_2896,N_2935);
and UO_43 (O_43,N_2723,N_2849);
nor UO_44 (O_44,N_2554,N_2799);
or UO_45 (O_45,N_2717,N_2735);
or UO_46 (O_46,N_2889,N_2597);
nor UO_47 (O_47,N_2789,N_2801);
or UO_48 (O_48,N_2572,N_2977);
nand UO_49 (O_49,N_2525,N_2887);
nand UO_50 (O_50,N_2796,N_2590);
nand UO_51 (O_51,N_2643,N_2501);
and UO_52 (O_52,N_2874,N_2775);
nand UO_53 (O_53,N_2895,N_2951);
or UO_54 (O_54,N_2561,N_2629);
xor UO_55 (O_55,N_2552,N_2948);
nor UO_56 (O_56,N_2678,N_2931);
xnor UO_57 (O_57,N_2702,N_2736);
nand UO_58 (O_58,N_2782,N_2871);
and UO_59 (O_59,N_2712,N_2952);
nand UO_60 (O_60,N_2595,N_2567);
nor UO_61 (O_61,N_2879,N_2966);
nor UO_62 (O_62,N_2555,N_2527);
or UO_63 (O_63,N_2528,N_2814);
and UO_64 (O_64,N_2797,N_2954);
nand UO_65 (O_65,N_2908,N_2689);
or UO_66 (O_66,N_2956,N_2787);
nand UO_67 (O_67,N_2638,N_2507);
or UO_68 (O_68,N_2713,N_2553);
and UO_69 (O_69,N_2606,N_2536);
nand UO_70 (O_70,N_2682,N_2925);
xnor UO_71 (O_71,N_2794,N_2544);
or UO_72 (O_72,N_2818,N_2560);
and UO_73 (O_73,N_2729,N_2877);
or UO_74 (O_74,N_2746,N_2551);
nand UO_75 (O_75,N_2575,N_2967);
nand UO_76 (O_76,N_2778,N_2731);
nand UO_77 (O_77,N_2774,N_2518);
xor UO_78 (O_78,N_2686,N_2696);
xor UO_79 (O_79,N_2989,N_2845);
xnor UO_80 (O_80,N_2500,N_2601);
or UO_81 (O_81,N_2998,N_2542);
or UO_82 (O_82,N_2706,N_2583);
xor UO_83 (O_83,N_2988,N_2777);
or UO_84 (O_84,N_2982,N_2812);
and UO_85 (O_85,N_2878,N_2904);
nand UO_86 (O_86,N_2837,N_2709);
nand UO_87 (O_87,N_2738,N_2512);
nor UO_88 (O_88,N_2733,N_2826);
and UO_89 (O_89,N_2732,N_2912);
and UO_90 (O_90,N_2669,N_2683);
nand UO_91 (O_91,N_2622,N_2838);
xnor UO_92 (O_92,N_2835,N_2891);
nor UO_93 (O_93,N_2607,N_2858);
nand UO_94 (O_94,N_2532,N_2978);
xor UO_95 (O_95,N_2993,N_2822);
or UO_96 (O_96,N_2885,N_2541);
and UO_97 (O_97,N_2593,N_2588);
nand UO_98 (O_98,N_2917,N_2721);
nor UO_99 (O_99,N_2634,N_2861);
nor UO_100 (O_100,N_2911,N_2548);
xor UO_101 (O_101,N_2747,N_2694);
or UO_102 (O_102,N_2716,N_2563);
nor UO_103 (O_103,N_2992,N_2829);
and UO_104 (O_104,N_2621,N_2585);
nand UO_105 (O_105,N_2519,N_2663);
nor UO_106 (O_106,N_2930,N_2517);
nand UO_107 (O_107,N_2944,N_2730);
and UO_108 (O_108,N_2937,N_2608);
or UO_109 (O_109,N_2785,N_2524);
nand UO_110 (O_110,N_2701,N_2979);
xnor UO_111 (O_111,N_2577,N_2584);
or UO_112 (O_112,N_2509,N_2708);
xor UO_113 (O_113,N_2947,N_2916);
nor UO_114 (O_114,N_2520,N_2860);
nand UO_115 (O_115,N_2919,N_2790);
nor UO_116 (O_116,N_2971,N_2617);
xnor UO_117 (O_117,N_2893,N_2869);
and UO_118 (O_118,N_2758,N_2894);
nand UO_119 (O_119,N_2626,N_2511);
or UO_120 (O_120,N_2784,N_2546);
or UO_121 (O_121,N_2579,N_2892);
nor UO_122 (O_122,N_2976,N_2753);
and UO_123 (O_123,N_2559,N_2668);
or UO_124 (O_124,N_2737,N_2700);
and UO_125 (O_125,N_2873,N_2899);
nor UO_126 (O_126,N_2594,N_2506);
or UO_127 (O_127,N_2592,N_2587);
and UO_128 (O_128,N_2964,N_2603);
nand UO_129 (O_129,N_2628,N_2934);
nand UO_130 (O_130,N_2631,N_2693);
nor UO_131 (O_131,N_2672,N_2902);
nand UO_132 (O_132,N_2531,N_2945);
or UO_133 (O_133,N_2820,N_2695);
or UO_134 (O_134,N_2957,N_2651);
and UO_135 (O_135,N_2928,N_2870);
nand UO_136 (O_136,N_2866,N_2802);
or UO_137 (O_137,N_2811,N_2969);
and UO_138 (O_138,N_2656,N_2939);
nand UO_139 (O_139,N_2900,N_2997);
and UO_140 (O_140,N_2503,N_2819);
and UO_141 (O_141,N_2722,N_2537);
or UO_142 (O_142,N_2679,N_2620);
and UO_143 (O_143,N_2614,N_2724);
nor UO_144 (O_144,N_2950,N_2574);
nand UO_145 (O_145,N_2685,N_2830);
nor UO_146 (O_146,N_2922,N_2576);
xnor UO_147 (O_147,N_2750,N_2666);
nand UO_148 (O_148,N_2875,N_2605);
or UO_149 (O_149,N_2619,N_2994);
or UO_150 (O_150,N_2901,N_2591);
and UO_151 (O_151,N_2646,N_2854);
or UO_152 (O_152,N_2882,N_2851);
or UO_153 (O_153,N_2921,N_2852);
and UO_154 (O_154,N_2942,N_2924);
nor UO_155 (O_155,N_2781,N_2960);
nor UO_156 (O_156,N_2910,N_2676);
and UO_157 (O_157,N_2578,N_2751);
and UO_158 (O_158,N_2827,N_2813);
nor UO_159 (O_159,N_2557,N_2985);
and UO_160 (O_160,N_2760,N_2568);
nor UO_161 (O_161,N_2652,N_2807);
or UO_162 (O_162,N_2855,N_2965);
nor UO_163 (O_163,N_2692,N_2865);
xor UO_164 (O_164,N_2580,N_2999);
nor UO_165 (O_165,N_2662,N_2623);
and UO_166 (O_166,N_2961,N_2540);
and UO_167 (O_167,N_2770,N_2857);
or UO_168 (O_168,N_2534,N_2581);
xor UO_169 (O_169,N_2740,N_2728);
nor UO_170 (O_170,N_2615,N_2876);
nor UO_171 (O_171,N_2856,N_2571);
or UO_172 (O_172,N_2981,N_2719);
or UO_173 (O_173,N_2611,N_2765);
xnor UO_174 (O_174,N_2890,N_2779);
nand UO_175 (O_175,N_2909,N_2691);
or UO_176 (O_176,N_2675,N_2644);
or UO_177 (O_177,N_2806,N_2647);
nor UO_178 (O_178,N_2953,N_2833);
nor UO_179 (O_179,N_2824,N_2545);
or UO_180 (O_180,N_2761,N_2842);
nand UO_181 (O_181,N_2793,N_2920);
and UO_182 (O_182,N_2613,N_2609);
nand UO_183 (O_183,N_2711,N_2625);
nand UO_184 (O_184,N_2959,N_2762);
or UO_185 (O_185,N_2905,N_2927);
xor UO_186 (O_186,N_2598,N_2754);
nand UO_187 (O_187,N_2718,N_2817);
nor UO_188 (O_188,N_2955,N_2624);
xnor UO_189 (O_189,N_2600,N_2828);
nor UO_190 (O_190,N_2771,N_2556);
nor UO_191 (O_191,N_2690,N_2795);
xnor UO_192 (O_192,N_2926,N_2958);
and UO_193 (O_193,N_2523,N_2549);
and UO_194 (O_194,N_2639,N_2550);
xnor UO_195 (O_195,N_2505,N_2767);
xnor UO_196 (O_196,N_2749,N_2667);
xor UO_197 (O_197,N_2834,N_2846);
nand UO_198 (O_198,N_2680,N_2618);
and UO_199 (O_199,N_2832,N_2582);
or UO_200 (O_200,N_2853,N_2972);
and UO_201 (O_201,N_2745,N_2815);
xor UO_202 (O_202,N_2915,N_2938);
xor UO_203 (O_203,N_2764,N_2809);
or UO_204 (O_204,N_2825,N_2918);
nand UO_205 (O_205,N_2674,N_2848);
nor UO_206 (O_206,N_2710,N_2547);
nand UO_207 (O_207,N_2707,N_2704);
nand UO_208 (O_208,N_2533,N_2963);
and UO_209 (O_209,N_2661,N_2980);
and UO_210 (O_210,N_2743,N_2699);
and UO_211 (O_211,N_2808,N_2836);
or UO_212 (O_212,N_2630,N_2844);
nor UO_213 (O_213,N_2868,N_2903);
xor UO_214 (O_214,N_2949,N_2897);
and UO_215 (O_215,N_2665,N_2648);
and UO_216 (O_216,N_2637,N_2657);
nand UO_217 (O_217,N_2831,N_2504);
nor UO_218 (O_218,N_2752,N_2821);
xnor UO_219 (O_219,N_2816,N_2610);
and UO_220 (O_220,N_2786,N_2670);
xor UO_221 (O_221,N_2703,N_2673);
and UO_222 (O_222,N_2940,N_2780);
nor UO_223 (O_223,N_2645,N_2635);
xnor UO_224 (O_224,N_2720,N_2803);
nand UO_225 (O_225,N_2888,N_2526);
nand UO_226 (O_226,N_2933,N_2602);
and UO_227 (O_227,N_2558,N_2810);
and UO_228 (O_228,N_2502,N_2766);
nor UO_229 (O_229,N_2932,N_2632);
nor UO_230 (O_230,N_2757,N_2664);
xor UO_231 (O_231,N_2768,N_2522);
nor UO_232 (O_232,N_2564,N_2734);
and UO_233 (O_233,N_2535,N_2616);
and UO_234 (O_234,N_2677,N_2841);
nand UO_235 (O_235,N_2516,N_2798);
and UO_236 (O_236,N_2772,N_2521);
or UO_237 (O_237,N_2589,N_2565);
or UO_238 (O_238,N_2654,N_2530);
nand UO_239 (O_239,N_2943,N_2684);
xnor UO_240 (O_240,N_2872,N_2660);
nor UO_241 (O_241,N_2513,N_2653);
and UO_242 (O_242,N_2906,N_2884);
or UO_243 (O_243,N_2658,N_2839);
nor UO_244 (O_244,N_2941,N_2655);
nand UO_245 (O_245,N_2867,N_2681);
xnor UO_246 (O_246,N_2688,N_2569);
nor UO_247 (O_247,N_2986,N_2983);
nor UO_248 (O_248,N_2742,N_2687);
or UO_249 (O_249,N_2539,N_2974);
xor UO_250 (O_250,N_2547,N_2944);
xnor UO_251 (O_251,N_2507,N_2953);
nor UO_252 (O_252,N_2755,N_2697);
xor UO_253 (O_253,N_2617,N_2858);
nor UO_254 (O_254,N_2748,N_2843);
nand UO_255 (O_255,N_2826,N_2667);
xnor UO_256 (O_256,N_2604,N_2957);
xnor UO_257 (O_257,N_2581,N_2566);
nor UO_258 (O_258,N_2784,N_2665);
and UO_259 (O_259,N_2629,N_2909);
or UO_260 (O_260,N_2547,N_2968);
nor UO_261 (O_261,N_2898,N_2837);
and UO_262 (O_262,N_2535,N_2972);
and UO_263 (O_263,N_2852,N_2916);
and UO_264 (O_264,N_2877,N_2589);
or UO_265 (O_265,N_2964,N_2812);
and UO_266 (O_266,N_2630,N_2853);
nand UO_267 (O_267,N_2901,N_2736);
xnor UO_268 (O_268,N_2842,N_2794);
and UO_269 (O_269,N_2714,N_2591);
xor UO_270 (O_270,N_2593,N_2761);
and UO_271 (O_271,N_2884,N_2620);
and UO_272 (O_272,N_2917,N_2663);
and UO_273 (O_273,N_2843,N_2757);
nor UO_274 (O_274,N_2842,N_2607);
nand UO_275 (O_275,N_2700,N_2772);
or UO_276 (O_276,N_2736,N_2856);
nor UO_277 (O_277,N_2747,N_2738);
nand UO_278 (O_278,N_2940,N_2539);
xor UO_279 (O_279,N_2867,N_2609);
or UO_280 (O_280,N_2958,N_2547);
xnor UO_281 (O_281,N_2516,N_2962);
nand UO_282 (O_282,N_2640,N_2994);
or UO_283 (O_283,N_2586,N_2801);
and UO_284 (O_284,N_2612,N_2672);
nand UO_285 (O_285,N_2624,N_2759);
or UO_286 (O_286,N_2579,N_2835);
or UO_287 (O_287,N_2712,N_2824);
nand UO_288 (O_288,N_2800,N_2854);
nand UO_289 (O_289,N_2623,N_2708);
nand UO_290 (O_290,N_2793,N_2751);
nand UO_291 (O_291,N_2774,N_2601);
nor UO_292 (O_292,N_2583,N_2746);
xnor UO_293 (O_293,N_2839,N_2588);
nand UO_294 (O_294,N_2922,N_2758);
and UO_295 (O_295,N_2681,N_2696);
nand UO_296 (O_296,N_2970,N_2895);
and UO_297 (O_297,N_2632,N_2875);
or UO_298 (O_298,N_2742,N_2739);
xnor UO_299 (O_299,N_2544,N_2667);
and UO_300 (O_300,N_2959,N_2552);
nand UO_301 (O_301,N_2764,N_2603);
and UO_302 (O_302,N_2745,N_2702);
nand UO_303 (O_303,N_2848,N_2609);
and UO_304 (O_304,N_2679,N_2974);
and UO_305 (O_305,N_2527,N_2557);
xnor UO_306 (O_306,N_2757,N_2569);
xnor UO_307 (O_307,N_2825,N_2796);
nand UO_308 (O_308,N_2917,N_2852);
and UO_309 (O_309,N_2681,N_2825);
nand UO_310 (O_310,N_2663,N_2927);
and UO_311 (O_311,N_2894,N_2860);
xnor UO_312 (O_312,N_2919,N_2708);
nor UO_313 (O_313,N_2512,N_2811);
or UO_314 (O_314,N_2990,N_2731);
xor UO_315 (O_315,N_2573,N_2965);
or UO_316 (O_316,N_2934,N_2912);
nand UO_317 (O_317,N_2683,N_2988);
or UO_318 (O_318,N_2814,N_2679);
or UO_319 (O_319,N_2636,N_2806);
and UO_320 (O_320,N_2704,N_2629);
or UO_321 (O_321,N_2525,N_2697);
xor UO_322 (O_322,N_2673,N_2817);
nand UO_323 (O_323,N_2857,N_2629);
nor UO_324 (O_324,N_2824,N_2516);
or UO_325 (O_325,N_2544,N_2580);
and UO_326 (O_326,N_2619,N_2685);
or UO_327 (O_327,N_2864,N_2911);
xor UO_328 (O_328,N_2762,N_2615);
and UO_329 (O_329,N_2993,N_2769);
nor UO_330 (O_330,N_2645,N_2582);
nand UO_331 (O_331,N_2747,N_2920);
and UO_332 (O_332,N_2703,N_2932);
and UO_333 (O_333,N_2797,N_2546);
and UO_334 (O_334,N_2752,N_2824);
or UO_335 (O_335,N_2768,N_2843);
nand UO_336 (O_336,N_2685,N_2558);
or UO_337 (O_337,N_2705,N_2808);
nor UO_338 (O_338,N_2772,N_2801);
nor UO_339 (O_339,N_2598,N_2699);
or UO_340 (O_340,N_2774,N_2941);
or UO_341 (O_341,N_2964,N_2913);
and UO_342 (O_342,N_2891,N_2604);
nand UO_343 (O_343,N_2797,N_2650);
nand UO_344 (O_344,N_2848,N_2577);
nand UO_345 (O_345,N_2808,N_2915);
or UO_346 (O_346,N_2937,N_2777);
xor UO_347 (O_347,N_2607,N_2623);
nor UO_348 (O_348,N_2833,N_2716);
nor UO_349 (O_349,N_2852,N_2910);
or UO_350 (O_350,N_2735,N_2908);
and UO_351 (O_351,N_2893,N_2885);
and UO_352 (O_352,N_2876,N_2991);
and UO_353 (O_353,N_2860,N_2522);
nand UO_354 (O_354,N_2654,N_2668);
xnor UO_355 (O_355,N_2708,N_2621);
nor UO_356 (O_356,N_2855,N_2925);
and UO_357 (O_357,N_2663,N_2817);
nand UO_358 (O_358,N_2903,N_2890);
or UO_359 (O_359,N_2805,N_2929);
nand UO_360 (O_360,N_2868,N_2838);
nor UO_361 (O_361,N_2569,N_2737);
and UO_362 (O_362,N_2743,N_2579);
and UO_363 (O_363,N_2551,N_2571);
or UO_364 (O_364,N_2955,N_2763);
and UO_365 (O_365,N_2576,N_2734);
nand UO_366 (O_366,N_2851,N_2649);
nor UO_367 (O_367,N_2614,N_2895);
and UO_368 (O_368,N_2610,N_2868);
nand UO_369 (O_369,N_2656,N_2668);
or UO_370 (O_370,N_2563,N_2893);
and UO_371 (O_371,N_2798,N_2837);
nor UO_372 (O_372,N_2809,N_2983);
or UO_373 (O_373,N_2868,N_2716);
and UO_374 (O_374,N_2716,N_2933);
or UO_375 (O_375,N_2595,N_2773);
or UO_376 (O_376,N_2890,N_2653);
or UO_377 (O_377,N_2758,N_2506);
nand UO_378 (O_378,N_2679,N_2560);
nand UO_379 (O_379,N_2884,N_2797);
xnor UO_380 (O_380,N_2908,N_2520);
or UO_381 (O_381,N_2692,N_2585);
nor UO_382 (O_382,N_2701,N_2910);
nand UO_383 (O_383,N_2673,N_2856);
and UO_384 (O_384,N_2914,N_2831);
or UO_385 (O_385,N_2543,N_2917);
nor UO_386 (O_386,N_2915,N_2650);
or UO_387 (O_387,N_2972,N_2888);
nor UO_388 (O_388,N_2836,N_2842);
xnor UO_389 (O_389,N_2875,N_2575);
nor UO_390 (O_390,N_2971,N_2696);
nor UO_391 (O_391,N_2650,N_2779);
xor UO_392 (O_392,N_2749,N_2727);
nor UO_393 (O_393,N_2731,N_2791);
xnor UO_394 (O_394,N_2858,N_2628);
and UO_395 (O_395,N_2737,N_2773);
nand UO_396 (O_396,N_2961,N_2646);
and UO_397 (O_397,N_2748,N_2754);
and UO_398 (O_398,N_2976,N_2577);
xor UO_399 (O_399,N_2761,N_2887);
and UO_400 (O_400,N_2683,N_2815);
xor UO_401 (O_401,N_2661,N_2642);
nor UO_402 (O_402,N_2784,N_2580);
or UO_403 (O_403,N_2921,N_2965);
nor UO_404 (O_404,N_2625,N_2926);
nand UO_405 (O_405,N_2974,N_2693);
xor UO_406 (O_406,N_2703,N_2519);
nor UO_407 (O_407,N_2727,N_2718);
or UO_408 (O_408,N_2729,N_2595);
and UO_409 (O_409,N_2653,N_2560);
and UO_410 (O_410,N_2822,N_2817);
and UO_411 (O_411,N_2962,N_2775);
and UO_412 (O_412,N_2979,N_2596);
nor UO_413 (O_413,N_2602,N_2905);
nor UO_414 (O_414,N_2511,N_2870);
nand UO_415 (O_415,N_2902,N_2970);
xnor UO_416 (O_416,N_2642,N_2631);
or UO_417 (O_417,N_2996,N_2884);
xnor UO_418 (O_418,N_2607,N_2555);
nand UO_419 (O_419,N_2995,N_2876);
nand UO_420 (O_420,N_2775,N_2960);
xor UO_421 (O_421,N_2885,N_2877);
xor UO_422 (O_422,N_2904,N_2937);
nor UO_423 (O_423,N_2990,N_2811);
xnor UO_424 (O_424,N_2636,N_2997);
and UO_425 (O_425,N_2688,N_2756);
nor UO_426 (O_426,N_2703,N_2577);
nand UO_427 (O_427,N_2982,N_2741);
and UO_428 (O_428,N_2706,N_2742);
and UO_429 (O_429,N_2934,N_2780);
or UO_430 (O_430,N_2624,N_2974);
nand UO_431 (O_431,N_2933,N_2561);
nand UO_432 (O_432,N_2736,N_2780);
xnor UO_433 (O_433,N_2904,N_2959);
nand UO_434 (O_434,N_2766,N_2518);
and UO_435 (O_435,N_2665,N_2738);
nand UO_436 (O_436,N_2934,N_2804);
or UO_437 (O_437,N_2976,N_2764);
and UO_438 (O_438,N_2688,N_2898);
and UO_439 (O_439,N_2991,N_2655);
and UO_440 (O_440,N_2537,N_2832);
or UO_441 (O_441,N_2939,N_2997);
nor UO_442 (O_442,N_2568,N_2534);
or UO_443 (O_443,N_2698,N_2776);
or UO_444 (O_444,N_2727,N_2674);
xor UO_445 (O_445,N_2606,N_2558);
or UO_446 (O_446,N_2770,N_2826);
nand UO_447 (O_447,N_2577,N_2661);
or UO_448 (O_448,N_2859,N_2633);
xor UO_449 (O_449,N_2504,N_2885);
xnor UO_450 (O_450,N_2538,N_2726);
and UO_451 (O_451,N_2779,N_2551);
and UO_452 (O_452,N_2619,N_2514);
xnor UO_453 (O_453,N_2662,N_2665);
xnor UO_454 (O_454,N_2999,N_2564);
and UO_455 (O_455,N_2625,N_2564);
nand UO_456 (O_456,N_2960,N_2975);
or UO_457 (O_457,N_2808,N_2913);
xor UO_458 (O_458,N_2815,N_2997);
and UO_459 (O_459,N_2642,N_2875);
or UO_460 (O_460,N_2674,N_2794);
and UO_461 (O_461,N_2725,N_2606);
nand UO_462 (O_462,N_2709,N_2945);
xnor UO_463 (O_463,N_2683,N_2760);
and UO_464 (O_464,N_2932,N_2990);
and UO_465 (O_465,N_2555,N_2997);
and UO_466 (O_466,N_2718,N_2843);
and UO_467 (O_467,N_2599,N_2701);
or UO_468 (O_468,N_2718,N_2778);
nor UO_469 (O_469,N_2794,N_2653);
xnor UO_470 (O_470,N_2602,N_2809);
or UO_471 (O_471,N_2810,N_2754);
nand UO_472 (O_472,N_2999,N_2774);
or UO_473 (O_473,N_2778,N_2661);
and UO_474 (O_474,N_2939,N_2717);
xnor UO_475 (O_475,N_2702,N_2696);
nand UO_476 (O_476,N_2800,N_2870);
and UO_477 (O_477,N_2680,N_2910);
nand UO_478 (O_478,N_2792,N_2822);
nor UO_479 (O_479,N_2901,N_2841);
xor UO_480 (O_480,N_2772,N_2637);
xnor UO_481 (O_481,N_2736,N_2790);
and UO_482 (O_482,N_2925,N_2829);
xnor UO_483 (O_483,N_2605,N_2703);
xnor UO_484 (O_484,N_2783,N_2543);
and UO_485 (O_485,N_2607,N_2633);
or UO_486 (O_486,N_2754,N_2734);
or UO_487 (O_487,N_2974,N_2943);
or UO_488 (O_488,N_2550,N_2846);
and UO_489 (O_489,N_2871,N_2551);
nand UO_490 (O_490,N_2679,N_2895);
nand UO_491 (O_491,N_2901,N_2597);
or UO_492 (O_492,N_2563,N_2956);
or UO_493 (O_493,N_2726,N_2928);
nor UO_494 (O_494,N_2840,N_2658);
nand UO_495 (O_495,N_2768,N_2905);
nand UO_496 (O_496,N_2555,N_2784);
xor UO_497 (O_497,N_2711,N_2706);
and UO_498 (O_498,N_2670,N_2601);
or UO_499 (O_499,N_2512,N_2940);
endmodule