module basic_2000_20000_2500_4_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_693,In_261);
and U1 (N_1,In_1310,In_1022);
xnor U2 (N_2,In_1340,In_1183);
or U3 (N_3,In_43,In_126);
and U4 (N_4,In_710,In_1087);
xor U5 (N_5,In_1979,In_677);
and U6 (N_6,In_567,In_1698);
nand U7 (N_7,In_1684,In_599);
xnor U8 (N_8,In_990,In_1637);
xor U9 (N_9,In_799,In_946);
xor U10 (N_10,In_912,In_795);
nand U11 (N_11,In_88,In_974);
xor U12 (N_12,In_582,In_1890);
nand U13 (N_13,In_123,In_1256);
nor U14 (N_14,In_897,In_505);
xnor U15 (N_15,In_153,In_1642);
and U16 (N_16,In_933,In_1804);
or U17 (N_17,In_102,In_1156);
nand U18 (N_18,In_1289,In_943);
and U19 (N_19,In_371,In_321);
nor U20 (N_20,In_1522,In_1826);
nor U21 (N_21,In_1753,In_213);
nor U22 (N_22,In_275,In_1773);
or U23 (N_23,In_1580,In_1261);
nor U24 (N_24,In_56,In_1357);
nor U25 (N_25,In_818,In_10);
or U26 (N_26,In_1540,In_1665);
nand U27 (N_27,In_924,In_381);
nor U28 (N_28,In_966,In_875);
and U29 (N_29,In_728,In_1696);
nor U30 (N_30,In_1635,In_1094);
nand U31 (N_31,In_4,In_1300);
or U32 (N_32,In_1863,In_1039);
xnor U33 (N_33,In_394,In_40);
nand U34 (N_34,In_197,In_1502);
or U35 (N_35,In_607,In_490);
nor U36 (N_36,In_141,In_923);
nand U37 (N_37,In_1151,In_1566);
xnor U38 (N_38,In_781,In_1251);
and U39 (N_39,In_1085,In_691);
nor U40 (N_40,In_545,In_904);
and U41 (N_41,In_867,In_31);
or U42 (N_42,In_30,In_753);
nand U43 (N_43,In_1672,In_1601);
or U44 (N_44,In_532,In_1434);
nor U45 (N_45,In_1180,In_942);
and U46 (N_46,In_898,In_1099);
or U47 (N_47,In_257,In_733);
xor U48 (N_48,In_1649,In_1072);
xnor U49 (N_49,In_313,In_354);
nand U50 (N_50,In_651,In_214);
xnor U51 (N_51,In_33,In_1882);
xnor U52 (N_52,In_209,In_439);
nor U53 (N_53,In_806,In_1402);
and U54 (N_54,In_1438,In_212);
or U55 (N_55,In_909,In_1046);
xor U56 (N_56,In_750,In_422);
nand U57 (N_57,In_235,In_1073);
and U58 (N_58,In_1596,In_1206);
and U59 (N_59,In_1880,In_1314);
and U60 (N_60,In_850,In_1062);
or U61 (N_61,In_1417,In_1690);
or U62 (N_62,In_177,In_879);
xnor U63 (N_63,In_1556,In_1608);
nor U64 (N_64,In_1510,In_1762);
or U65 (N_65,In_1348,In_1155);
or U66 (N_66,In_715,In_1385);
nand U67 (N_67,In_264,In_903);
and U68 (N_68,In_1000,In_719);
nand U69 (N_69,In_1888,In_657);
nor U70 (N_70,In_736,In_1021);
nor U71 (N_71,In_1600,In_117);
xnor U72 (N_72,In_411,In_1875);
nand U73 (N_73,In_253,In_999);
xnor U74 (N_74,In_1767,In_470);
and U75 (N_75,In_1704,In_805);
or U76 (N_76,In_198,In_1053);
nand U77 (N_77,In_1104,In_992);
xnor U78 (N_78,In_62,In_1164);
and U79 (N_79,In_959,In_154);
nor U80 (N_80,In_695,In_383);
xnor U81 (N_81,In_1306,In_618);
xor U82 (N_82,In_1913,In_1865);
nand U83 (N_83,In_1627,In_796);
nor U84 (N_84,In_1236,In_1924);
and U85 (N_85,In_1383,In_1332);
and U86 (N_86,In_614,In_1598);
xnor U87 (N_87,In_466,In_1778);
and U88 (N_88,In_1214,In_108);
or U89 (N_89,In_45,In_399);
nor U90 (N_90,In_522,In_1508);
or U91 (N_91,In_1721,In_1080);
nand U92 (N_92,In_165,In_1195);
or U93 (N_93,In_889,In_940);
nand U94 (N_94,In_143,In_670);
xnor U95 (N_95,In_1377,In_1070);
nor U96 (N_96,In_1802,In_1136);
nor U97 (N_97,In_191,In_1747);
nor U98 (N_98,In_1602,In_1727);
nand U99 (N_99,In_1414,In_229);
and U100 (N_100,In_487,In_1892);
nor U101 (N_101,In_1234,In_1707);
xnor U102 (N_102,In_449,In_1049);
and U103 (N_103,In_1037,In_134);
and U104 (N_104,In_1106,In_969);
xnor U105 (N_105,In_506,In_1638);
nand U106 (N_106,In_1551,In_1681);
or U107 (N_107,In_916,In_1650);
xor U108 (N_108,In_574,In_975);
or U109 (N_109,In_544,In_1130);
nor U110 (N_110,In_1683,In_1565);
xnor U111 (N_111,In_888,In_914);
nor U112 (N_112,In_420,In_1969);
nor U113 (N_113,In_1008,In_1299);
nor U114 (N_114,In_666,In_1670);
xnor U115 (N_115,In_442,In_1339);
nor U116 (N_116,In_260,In_1862);
and U117 (N_117,In_1978,In_484);
and U118 (N_118,In_745,In_1581);
nand U119 (N_119,In_1280,In_1504);
nand U120 (N_120,In_917,In_39);
xor U121 (N_121,In_1571,In_1895);
nand U122 (N_122,In_1125,In_1856);
xnor U123 (N_123,In_182,In_678);
nor U124 (N_124,In_1382,In_1176);
nor U125 (N_125,In_1415,In_519);
and U126 (N_126,In_1406,In_1217);
or U127 (N_127,In_389,In_118);
xor U128 (N_128,In_1379,In_921);
and U129 (N_129,In_823,In_90);
xnor U130 (N_130,In_479,In_988);
and U131 (N_131,In_1906,In_638);
and U132 (N_132,In_436,In_1981);
and U133 (N_133,In_396,In_1883);
nand U134 (N_134,In_1931,In_1497);
and U135 (N_135,In_288,In_1606);
nor U136 (N_136,In_873,In_619);
nor U137 (N_137,In_1149,In_1735);
nor U138 (N_138,In_1868,In_107);
nor U139 (N_139,In_534,In_902);
or U140 (N_140,In_830,In_747);
and U141 (N_141,In_206,In_1347);
and U142 (N_142,In_149,In_1489);
and U143 (N_143,In_148,In_1536);
nand U144 (N_144,In_1264,In_1364);
nand U145 (N_145,In_1367,In_308);
and U146 (N_146,In_970,In_1060);
or U147 (N_147,In_652,In_1419);
and U148 (N_148,In_299,In_832);
xor U149 (N_149,In_485,In_878);
nor U150 (N_150,In_391,In_1610);
xor U151 (N_151,In_1171,In_1576);
xnor U152 (N_152,In_1129,In_663);
or U153 (N_153,In_1173,In_502);
nand U154 (N_154,In_1886,In_103);
nor U155 (N_155,In_1829,In_827);
nand U156 (N_156,In_1474,In_406);
xnor U157 (N_157,In_312,In_233);
xor U158 (N_158,In_1421,In_1559);
xnor U159 (N_159,In_293,In_1546);
nor U160 (N_160,In_1639,In_1718);
and U161 (N_161,In_981,In_160);
or U162 (N_162,In_512,In_549);
nand U163 (N_163,In_530,In_1273);
and U164 (N_164,In_1059,In_855);
and U165 (N_165,In_106,In_1607);
and U166 (N_166,In_709,In_1633);
and U167 (N_167,In_221,In_847);
or U168 (N_168,In_460,In_964);
xor U169 (N_169,In_611,In_468);
or U170 (N_170,In_1496,In_1617);
xnor U171 (N_171,In_415,In_155);
xnor U172 (N_172,In_1398,In_1745);
nor U173 (N_173,In_23,In_1561);
or U174 (N_174,In_1462,In_1801);
nor U175 (N_175,In_1492,In_1507);
or U176 (N_176,In_244,In_1354);
xor U177 (N_177,In_1433,In_1957);
nor U178 (N_178,In_1679,In_1884);
xor U179 (N_179,In_132,In_989);
xnor U180 (N_180,In_1488,In_1248);
nor U181 (N_181,In_1994,In_12);
or U182 (N_182,In_962,In_448);
nand U183 (N_183,In_1612,In_1946);
or U184 (N_184,In_334,In_782);
nand U185 (N_185,In_294,In_1734);
nor U186 (N_186,In_1452,In_410);
and U187 (N_187,In_1772,In_324);
and U188 (N_188,In_29,In_471);
and U189 (N_189,In_386,In_1834);
xnor U190 (N_190,In_729,In_1041);
and U191 (N_191,In_1618,In_1160);
nand U192 (N_192,In_1418,In_1036);
xor U193 (N_193,In_584,In_1885);
nor U194 (N_194,In_105,In_227);
xnor U195 (N_195,In_1876,In_1515);
and U196 (N_196,In_1451,In_1756);
and U197 (N_197,In_248,In_413);
or U198 (N_198,In_373,In_1476);
xor U199 (N_199,In_707,In_403);
or U200 (N_200,In_204,In_284);
or U201 (N_201,In_626,In_359);
and U202 (N_202,In_1102,In_1014);
xnor U203 (N_203,In_1475,In_16);
and U204 (N_204,In_1032,In_402);
and U205 (N_205,In_1712,In_857);
xor U206 (N_206,In_79,In_292);
xor U207 (N_207,In_97,In_1442);
or U208 (N_208,In_1467,In_1643);
xnor U209 (N_209,In_1737,In_1222);
and U210 (N_210,In_690,In_899);
and U211 (N_211,In_3,In_412);
and U212 (N_212,In_535,In_537);
nand U213 (N_213,In_667,In_110);
and U214 (N_214,In_780,In_1907);
nand U215 (N_215,In_1320,In_1422);
and U216 (N_216,In_891,In_127);
xnor U217 (N_217,In_1569,In_1653);
or U218 (N_218,In_846,In_1594);
nor U219 (N_219,In_1221,In_685);
or U220 (N_220,In_527,In_1345);
nor U221 (N_221,In_1168,In_1803);
nor U222 (N_222,In_800,In_1274);
xnor U223 (N_223,In_147,In_1212);
or U224 (N_224,In_83,In_1544);
nor U225 (N_225,In_1460,In_301);
nand U226 (N_226,In_1832,In_1524);
nand U227 (N_227,In_1459,In_556);
xnor U228 (N_228,In_557,In_886);
nor U229 (N_229,In_1381,In_1064);
nor U230 (N_230,In_428,In_1901);
nor U231 (N_231,In_1330,In_1947);
and U232 (N_232,In_372,In_408);
nand U233 (N_233,In_600,In_392);
xor U234 (N_234,In_590,In_0);
and U235 (N_235,In_189,In_1407);
xor U236 (N_236,In_1687,In_1484);
and U237 (N_237,In_978,In_1131);
and U238 (N_238,In_1575,In_342);
and U239 (N_239,In_1268,In_1847);
nand U240 (N_240,In_1819,In_765);
xnor U241 (N_241,In_1035,In_347);
nand U242 (N_242,In_1004,In_13);
or U243 (N_243,In_1031,In_1447);
nor U244 (N_244,In_1799,In_673);
nand U245 (N_245,In_85,In_1584);
and U246 (N_246,In_605,In_1470);
xnor U247 (N_247,In_1403,In_186);
xnor U248 (N_248,In_36,In_896);
xor U249 (N_249,In_1355,In_1420);
nand U250 (N_250,In_151,In_1291);
nor U251 (N_251,In_499,In_700);
and U252 (N_252,In_1161,In_547);
xor U253 (N_253,In_936,In_1239);
nand U254 (N_254,In_508,In_880);
nand U255 (N_255,In_825,In_1869);
nand U256 (N_256,In_1919,In_1597);
xor U257 (N_257,In_711,In_998);
and U258 (N_258,In_98,In_1716);
nor U259 (N_259,In_1976,In_1245);
xor U260 (N_260,In_1686,In_675);
nor U261 (N_261,In_1086,In_792);
and U262 (N_262,In_1954,In_205);
xor U263 (N_263,In_1333,In_318);
nor U264 (N_264,In_60,In_735);
and U265 (N_265,In_188,In_1172);
xnor U266 (N_266,In_1817,In_1674);
or U267 (N_267,In_456,In_330);
and U268 (N_268,In_1654,In_200);
or U269 (N_269,In_1843,In_554);
xor U270 (N_270,In_1232,In_616);
nand U271 (N_271,In_384,In_1401);
or U272 (N_272,In_349,In_1436);
nand U273 (N_273,In_525,In_1108);
xnor U274 (N_274,In_1793,In_784);
nand U275 (N_275,In_844,In_791);
xor U276 (N_276,In_9,In_174);
nand U277 (N_277,In_1162,In_459);
and U278 (N_278,In_250,In_280);
nand U279 (N_279,In_1917,In_247);
nand U280 (N_280,In_941,In_1067);
nand U281 (N_281,In_314,In_1092);
or U282 (N_282,In_374,In_404);
nand U283 (N_283,In_1481,In_1193);
and U284 (N_284,In_524,In_1450);
and U285 (N_285,In_375,In_445);
nand U286 (N_286,In_698,In_734);
nor U287 (N_287,In_1996,In_1246);
nor U288 (N_288,In_885,In_669);
xor U289 (N_289,In_409,In_1900);
xor U290 (N_290,In_96,In_1916);
and U291 (N_291,In_538,In_1873);
xor U292 (N_292,In_895,In_104);
nand U293 (N_293,In_1061,In_1084);
and U294 (N_294,In_1758,In_653);
nor U295 (N_295,In_682,In_778);
nor U296 (N_296,In_1097,In_232);
nor U297 (N_297,In_272,In_1257);
and U298 (N_298,In_1995,In_357);
or U299 (N_299,In_1609,In_1122);
and U300 (N_300,In_637,In_430);
and U301 (N_301,In_124,In_71);
nor U302 (N_302,In_571,In_274);
xor U303 (N_303,In_376,In_401);
or U304 (N_304,In_1150,In_1668);
nand U305 (N_305,In_911,In_1361);
or U306 (N_306,In_1628,In_1350);
nor U307 (N_307,In_1018,In_730);
nor U308 (N_308,In_1558,In_1203);
nand U309 (N_309,In_1837,In_1187);
or U310 (N_310,In_564,In_771);
nand U311 (N_311,In_1430,In_1867);
nor U312 (N_312,In_1293,In_1741);
nand U313 (N_313,In_1529,In_370);
nor U314 (N_314,In_683,In_1990);
nor U315 (N_315,In_1237,In_737);
nand U316 (N_316,In_1482,In_196);
nand U317 (N_317,In_146,In_89);
xnor U318 (N_318,In_424,In_202);
nand U319 (N_319,In_433,In_54);
nand U320 (N_320,In_1325,In_1063);
nand U321 (N_321,In_1233,In_749);
xnor U322 (N_322,In_822,In_1848);
xnor U323 (N_323,In_1667,In_469);
and U324 (N_324,In_491,In_1375);
xnor U325 (N_325,In_1748,In_1523);
nor U326 (N_326,In_1960,In_1751);
nor U327 (N_327,In_230,In_379);
nor U328 (N_328,In_1699,In_594);
and U329 (N_329,In_720,In_22);
and U330 (N_330,In_1531,In_1912);
nand U331 (N_331,In_176,In_1999);
nor U332 (N_332,In_788,In_915);
nor U333 (N_333,In_608,In_1105);
or U334 (N_334,In_440,In_1042);
xor U335 (N_335,In_1077,In_851);
xor U336 (N_336,In_1213,In_1055);
or U337 (N_337,In_503,In_1505);
and U338 (N_338,In_1045,In_1872);
or U339 (N_339,In_1956,In_829);
or U340 (N_340,In_131,In_723);
xnor U341 (N_341,In_526,In_1316);
and U342 (N_342,In_1694,In_533);
or U343 (N_343,In_363,In_659);
and U344 (N_344,In_1644,In_1360);
and U345 (N_345,In_759,In_1208);
xor U346 (N_346,In_355,In_963);
or U347 (N_347,In_1790,In_1537);
and U348 (N_348,In_388,In_1615);
and U349 (N_349,In_1849,In_1705);
or U350 (N_350,In_1166,In_872);
or U351 (N_351,In_1645,In_518);
nand U352 (N_352,In_658,In_493);
or U353 (N_353,In_234,In_344);
nor U354 (N_354,In_699,In_377);
and U355 (N_355,In_1216,In_1282);
or U356 (N_356,In_1223,In_511);
nand U357 (N_357,In_1701,In_1689);
nand U358 (N_358,In_152,In_1307);
xor U359 (N_359,In_612,In_425);
or U360 (N_360,In_335,In_1851);
nand U361 (N_361,In_429,In_70);
nor U362 (N_362,In_310,In_1089);
or U363 (N_363,In_953,In_1044);
or U364 (N_364,In_713,In_92);
nor U365 (N_365,In_1939,In_708);
nand U366 (N_366,In_1542,In_1011);
nor U367 (N_367,In_1958,In_853);
or U368 (N_368,In_1308,In_1614);
nor U369 (N_369,In_803,In_874);
and U370 (N_370,In_239,In_671);
nor U371 (N_371,In_722,In_1368);
xor U372 (N_372,In_520,In_842);
nor U373 (N_373,In_368,In_282);
or U374 (N_374,In_1528,In_1292);
nor U375 (N_375,In_1201,In_1750);
and U376 (N_376,In_934,In_835);
and U377 (N_377,In_919,In_1968);
xnor U378 (N_378,In_1238,In_1113);
nand U379 (N_379,In_1514,In_1324);
and U380 (N_380,In_365,In_304);
and U381 (N_381,In_1365,In_1048);
nor U382 (N_382,In_1940,In_810);
xnor U383 (N_383,In_1950,In_1478);
nand U384 (N_384,In_1126,In_591);
xnor U385 (N_385,In_1530,In_1552);
nor U386 (N_386,In_37,In_461);
and U387 (N_387,In_441,In_732);
xor U388 (N_388,In_1980,In_1013);
nor U389 (N_389,In_15,In_1853);
nor U390 (N_390,In_325,In_987);
nor U391 (N_391,In_1592,In_1091);
or U392 (N_392,In_1527,In_1294);
xor U393 (N_393,In_854,In_315);
and U394 (N_394,In_680,In_965);
xor U395 (N_395,In_483,In_967);
nand U396 (N_396,In_1296,In_1855);
xor U397 (N_397,In_1792,In_341);
xor U398 (N_398,In_1319,In_1736);
nand U399 (N_399,In_225,In_138);
and U400 (N_400,In_812,In_1586);
nand U401 (N_401,In_418,In_985);
xor U402 (N_402,In_1518,In_1194);
or U403 (N_403,In_1432,In_1386);
and U404 (N_404,In_1700,In_38);
nor U405 (N_405,In_305,In_639);
and U406 (N_406,In_701,In_845);
and U407 (N_407,In_1871,In_1656);
nor U408 (N_408,In_64,In_297);
xnor U409 (N_409,In_817,In_1866);
nand U410 (N_410,In_1850,In_1831);
nand U411 (N_411,In_1394,In_979);
nand U412 (N_412,In_1797,In_1074);
or U413 (N_413,In_434,In_1358);
nand U414 (N_414,In_774,In_1798);
or U415 (N_415,In_1119,In_1247);
and U416 (N_416,In_119,In_164);
and U417 (N_417,In_1148,In_190);
and U418 (N_418,In_1275,In_553);
and U419 (N_419,In_1265,In_1971);
xnor U420 (N_420,In_361,In_1229);
or U421 (N_421,In_1134,In_358);
or U422 (N_422,In_661,In_1854);
xor U423 (N_423,In_517,In_1154);
xnor U424 (N_424,In_1153,In_1163);
xnor U425 (N_425,In_770,In_1657);
xor U426 (N_426,In_1408,In_1362);
nor U427 (N_427,In_1814,In_793);
or U428 (N_428,In_597,In_1137);
or U429 (N_429,In_566,In_1413);
or U430 (N_430,In_416,In_50);
or U431 (N_431,In_1393,In_339);
nor U432 (N_432,In_871,In_210);
and U433 (N_433,In_907,In_5);
nand U434 (N_434,In_1953,In_478);
and U435 (N_435,In_776,In_1192);
or U436 (N_436,In_203,In_926);
xor U437 (N_437,In_1336,In_1186);
xor U438 (N_438,In_1346,In_1692);
nand U439 (N_439,In_258,In_1342);
nor U440 (N_440,In_704,In_1260);
and U441 (N_441,In_1219,In_1374);
and U442 (N_442,In_1915,In_906);
nand U443 (N_443,In_928,In_382);
and U444 (N_444,In_1746,In_565);
nor U445 (N_445,In_684,In_801);
nand U446 (N_446,In_1123,In_1709);
or U447 (N_447,In_1006,In_1779);
nand U448 (N_448,In_760,In_1555);
xnor U449 (N_449,In_1152,In_1241);
xnor U450 (N_450,In_1791,In_86);
or U451 (N_451,In_1483,In_1052);
nor U452 (N_452,In_496,In_217);
and U453 (N_453,In_1982,In_681);
nor U454 (N_454,In_1807,In_6);
nor U455 (N_455,In_1144,In_1664);
xor U456 (N_456,In_580,In_1749);
nand U457 (N_457,In_350,In_1646);
nor U458 (N_458,In_884,In_465);
and U459 (N_459,In_971,In_1965);
nor U460 (N_460,In_1519,In_1846);
or U461 (N_461,In_259,In_1179);
nor U462 (N_462,In_1998,In_1839);
nand U463 (N_463,In_1114,In_834);
nor U464 (N_464,In_621,In_1881);
xor U465 (N_465,In_1455,In_668);
nor U466 (N_466,In_289,In_562);
nor U467 (N_467,In_647,In_1605);
and U468 (N_468,In_929,In_1424);
and U469 (N_469,In_1103,In_1720);
nand U470 (N_470,In_1286,In_457);
nor U471 (N_471,In_1509,In_369);
nand U472 (N_472,In_52,In_378);
or U473 (N_473,In_1763,In_474);
and U474 (N_474,In_109,In_61);
and U475 (N_475,In_1396,In_1050);
nand U476 (N_476,In_1445,In_1812);
or U477 (N_477,In_1526,In_492);
nor U478 (N_478,In_1040,In_169);
and U479 (N_479,In_1399,In_498);
or U480 (N_480,In_727,In_1794);
or U481 (N_481,In_1541,In_1285);
or U482 (N_482,In_150,In_1276);
nand U483 (N_483,In_1677,In_1202);
xnor U484 (N_484,In_655,In_1949);
or U485 (N_485,In_1927,In_1648);
and U486 (N_486,In_1242,In_262);
xor U487 (N_487,In_1093,In_1057);
nand U488 (N_488,In_72,In_1047);
xor U489 (N_489,In_1189,In_996);
nor U490 (N_490,In_620,In_757);
or U491 (N_491,In_1457,In_636);
or U492 (N_492,In_601,In_1659);
xor U493 (N_493,In_219,In_306);
or U494 (N_494,In_20,In_1009);
nand U495 (N_495,In_1412,In_1107);
nand U496 (N_496,In_346,In_1444);
and U497 (N_497,In_552,In_397);
xnor U498 (N_498,In_1120,In_41);
nand U499 (N_499,In_954,In_1963);
and U500 (N_500,In_1977,In_1503);
or U501 (N_501,In_26,In_746);
nand U502 (N_502,In_320,In_161);
and U503 (N_503,In_1570,In_432);
or U504 (N_504,In_278,In_837);
and U505 (N_505,In_1005,In_101);
xor U506 (N_506,In_180,In_1277);
or U507 (N_507,In_362,In_1992);
nor U508 (N_508,In_1955,In_208);
nor U509 (N_509,In_598,In_1015);
and U510 (N_510,In_1535,In_1376);
and U511 (N_511,In_265,In_1328);
xor U512 (N_512,In_163,In_631);
nand U513 (N_513,In_1641,In_192);
nand U514 (N_514,In_19,In_863);
and U515 (N_515,In_1454,In_252);
and U516 (N_516,In_431,In_311);
xor U517 (N_517,In_489,In_218);
nor U518 (N_518,In_625,In_1538);
nor U519 (N_519,In_380,In_650);
nor U520 (N_520,In_516,In_694);
and U521 (N_521,In_504,In_1490);
nand U522 (N_522,In_1288,In_319);
or U523 (N_523,In_215,In_1711);
xor U524 (N_524,In_649,In_1076);
or U525 (N_525,In_1822,In_1796);
nand U526 (N_526,In_513,In_34);
or U527 (N_527,In_665,In_944);
nor U528 (N_528,In_1572,In_1338);
and U529 (N_529,In_78,In_283);
nand U530 (N_530,In_951,In_1770);
nor U531 (N_531,In_73,In_849);
nor U532 (N_532,In_287,In_1170);
nand U533 (N_533,In_1599,In_798);
nand U534 (N_534,In_1722,In_1910);
xor U535 (N_535,In_277,In_1431);
nand U536 (N_536,In_1781,In_1972);
and U537 (N_537,In_1027,In_1185);
and U538 (N_538,In_1929,In_866);
xor U539 (N_539,In_1833,In_1337);
or U540 (N_540,In_1416,In_1962);
nand U541 (N_541,In_1409,In_576);
and U542 (N_542,In_762,In_838);
nand U543 (N_543,In_1210,In_1010);
xnor U544 (N_544,In_1662,In_142);
nand U545 (N_545,In_1279,In_1761);
nand U546 (N_546,In_1859,In_1682);
nor U547 (N_547,In_1620,In_558);
nor U548 (N_548,In_1673,In_360);
or U549 (N_549,In_1302,In_1456);
nand U550 (N_550,In_686,In_1001);
nor U551 (N_551,In_1808,In_1397);
nand U552 (N_552,In_1651,In_761);
xor U553 (N_553,In_1564,In_1738);
nand U554 (N_554,In_1220,In_1717);
xor U555 (N_555,In_1908,In_99);
xnor U556 (N_556,In_1071,In_414);
and U557 (N_557,In_642,In_1218);
nand U558 (N_558,In_602,In_581);
nor U559 (N_559,In_1007,In_1016);
nor U560 (N_560,In_1023,In_44);
and U561 (N_561,In_1487,In_551);
nand U562 (N_562,In_1317,In_758);
and U563 (N_563,In_270,In_949);
and U564 (N_564,In_1623,In_1587);
nor U565 (N_565,In_569,In_1780);
xor U566 (N_566,In_1743,In_1577);
or U567 (N_567,In_1054,In_1889);
nand U568 (N_568,In_1028,In_843);
or U569 (N_569,In_688,In_1318);
and U570 (N_570,In_158,In_268);
nor U571 (N_571,In_1928,In_646);
xor U572 (N_572,In_450,In_1935);
nor U573 (N_573,In_1771,In_839);
xnor U574 (N_574,In_1197,In_568);
nand U575 (N_575,In_1078,In_931);
xor U576 (N_576,In_57,In_323);
nor U577 (N_577,In_1585,In_1404);
xor U578 (N_578,In_1811,In_859);
xor U579 (N_579,In_982,In_1621);
nor U580 (N_580,In_955,In_592);
nor U581 (N_581,In_922,In_1616);
nor U582 (N_582,In_1553,In_1517);
nor U583 (N_583,In_1765,In_1661);
or U584 (N_584,In_162,In_1539);
nand U585 (N_585,In_1930,In_819);
and U586 (N_586,In_634,In_135);
and U587 (N_587,In_1026,In_286);
and U588 (N_588,In_1343,In_193);
xnor U589 (N_589,In_240,In_47);
xor U590 (N_590,In_632,In_331);
xor U591 (N_591,In_595,In_1703);
or U592 (N_592,In_1098,In_1205);
nand U593 (N_593,In_276,In_654);
nor U594 (N_594,In_702,In_112);
xnor U595 (N_595,In_1469,In_1961);
or U596 (N_596,In_629,In_1550);
nand U597 (N_597,In_1691,In_583);
xor U598 (N_598,In_1845,In_351);
nand U599 (N_599,In_1353,In_1352);
and U600 (N_600,In_1991,In_560);
xnor U601 (N_601,In_236,In_766);
nand U602 (N_602,In_273,In_712);
and U603 (N_603,In_285,In_263);
xnor U604 (N_604,In_1341,In_1904);
nor U605 (N_605,In_453,In_1934);
nand U606 (N_606,In_1909,In_811);
or U607 (N_607,In_1278,In_1730);
and U608 (N_608,In_1012,In_1858);
or U609 (N_609,In_24,In_387);
nor U610 (N_610,In_1787,In_1427);
nand U611 (N_611,In_643,In_184);
nor U612 (N_612,In_1334,In_11);
and U613 (N_613,In_1259,In_1918);
nor U614 (N_614,In_1878,In_175);
or U615 (N_615,In_1169,In_495);
nand U616 (N_616,In_271,In_500);
and U617 (N_617,In_1100,In_81);
nand U618 (N_618,In_1461,In_773);
nand U619 (N_619,In_1088,In_220);
xnor U620 (N_620,In_1464,In_1877);
nor U621 (N_621,In_14,In_366);
nand U622 (N_622,In_692,In_1243);
xor U623 (N_623,In_1574,In_1254);
or U624 (N_624,In_748,In_231);
nor U625 (N_625,In_816,In_1157);
and U626 (N_626,In_1384,In_1902);
and U627 (N_627,In_333,In_84);
or U628 (N_628,In_1760,In_932);
and U629 (N_629,In_1270,In_1304);
xor U630 (N_630,In_145,In_1477);
nor U631 (N_631,In_1019,In_94);
xor U632 (N_632,In_400,In_1740);
and U633 (N_633,In_1312,In_622);
nand U634 (N_634,In_443,In_332);
xor U635 (N_635,In_51,In_458);
xnor U636 (N_636,In_281,In_993);
and U637 (N_637,In_645,In_473);
and U638 (N_638,In_1321,In_266);
nand U639 (N_639,In_840,In_905);
xnor U640 (N_640,In_1135,In_1733);
nand U641 (N_641,In_223,In_1159);
nand U642 (N_642,In_35,In_1754);
xor U643 (N_643,In_1786,In_435);
nor U644 (N_644,In_1498,In_1744);
and U645 (N_645,In_744,In_1305);
nand U646 (N_646,In_1175,In_984);
or U647 (N_647,In_1590,In_115);
nand U648 (N_648,In_1471,In_438);
and U649 (N_649,In_1486,In_676);
nor U650 (N_650,In_648,In_1117);
and U651 (N_651,In_1631,In_1174);
nand U652 (N_652,In_1723,In_706);
and U653 (N_653,In_507,In_1548);
xnor U654 (N_654,In_1993,In_578);
nand U655 (N_655,In_1491,In_1267);
or U656 (N_656,In_848,In_201);
nor U657 (N_657,In_785,In_199);
or U658 (N_658,In_1782,In_937);
or U659 (N_659,In_353,In_893);
and U660 (N_660,In_405,In_1387);
nor U661 (N_661,In_714,In_166);
xor U662 (N_662,In_797,In_1380);
and U663 (N_663,In_58,In_1922);
xnor U664 (N_664,In_1271,In_1521);
nand U665 (N_665,In_1287,In_555);
nand U666 (N_666,In_1516,In_452);
nand U667 (N_667,In_1611,In_1116);
and U668 (N_668,In_997,In_1784);
xor U669 (N_669,In_1426,In_786);
nor U670 (N_670,In_444,In_1051);
xnor U671 (N_671,In_1813,In_1997);
nand U672 (N_672,In_738,In_587);
nor U673 (N_673,In_1678,In_1143);
xnor U674 (N_674,In_1636,In_1309);
nand U675 (N_675,In_1188,In_1920);
and U676 (N_676,In_1942,In_925);
nor U677 (N_677,In_1959,In_881);
nor U678 (N_678,In_187,In_1369);
or U679 (N_679,In_1827,In_423);
xor U680 (N_680,In_1788,In_588);
nor U681 (N_681,In_664,In_1405);
nor U682 (N_682,In_808,In_1675);
xnor U683 (N_683,In_497,In_1002);
nor U684 (N_684,In_628,In_1830);
and U685 (N_685,In_716,In_877);
nor U686 (N_686,In_1595,In_1485);
or U687 (N_687,In_17,In_920);
xor U688 (N_688,In_1435,In_865);
xor U689 (N_689,In_575,In_1588);
and U690 (N_690,In_1842,In_279);
nor U691 (N_691,In_935,In_1715);
nand U692 (N_692,In_1020,In_129);
xor U693 (N_693,In_585,In_1759);
or U694 (N_694,In_858,In_1764);
xor U695 (N_695,In_1634,In_1140);
and U696 (N_696,In_1964,In_1914);
nor U697 (N_697,In_1583,In_1446);
and U698 (N_698,In_1766,In_367);
or U699 (N_699,In_1728,In_972);
nor U700 (N_700,In_211,In_296);
xor U701 (N_701,In_894,In_833);
and U702 (N_702,In_1768,In_345);
nand U703 (N_703,In_1591,In_1472);
xnor U704 (N_704,In_860,In_245);
nor U705 (N_705,In_1861,In_65);
and U706 (N_706,In_222,In_957);
xor U707 (N_707,In_1563,In_1178);
nand U708 (N_708,In_1056,In_1816);
nor U709 (N_709,In_156,In_1025);
or U710 (N_710,In_789,In_1923);
or U711 (N_711,In_1899,In_1165);
or U712 (N_712,In_1984,In_1331);
nand U713 (N_713,In_1543,In_1757);
and U714 (N_714,In_828,In_1896);
nand U715 (N_715,In_1702,In_462);
or U716 (N_716,In_831,In_1640);
nand U717 (N_717,In_820,In_1303);
xnor U718 (N_718,In_1501,In_1695);
xnor U719 (N_719,In_116,In_1755);
or U720 (N_720,In_113,In_1809);
nand U721 (N_721,In_1685,In_1810);
or U722 (N_722,In_139,In_1520);
nand U723 (N_723,In_1295,In_224);
and U724 (N_724,In_1731,In_291);
nand U725 (N_725,In_624,In_1262);
nand U726 (N_726,In_824,In_1970);
xnor U727 (N_727,In_1603,In_1789);
xor U728 (N_728,In_317,In_892);
nand U729 (N_729,In_251,In_1506);
nand U730 (N_730,In_168,In_1824);
xnor U731 (N_731,In_1207,In_751);
xor U732 (N_732,In_53,In_821);
nand U733 (N_733,In_772,In_804);
nand U734 (N_734,In_76,In_1429);
and U735 (N_735,In_322,In_703);
nand U736 (N_736,In_1622,In_1582);
nor U737 (N_737,In_1857,In_1676);
or U738 (N_738,In_1196,In_1775);
nand U739 (N_739,In_1619,In_973);
xnor U740 (N_740,In_510,In_900);
nor U741 (N_741,In_1370,In_364);
nor U742 (N_742,In_242,In_337);
or U743 (N_743,In_1141,In_307);
xor U744 (N_744,In_977,In_1647);
and U745 (N_745,In_1142,In_994);
and U746 (N_746,In_1921,In_1167);
nor U747 (N_747,In_300,In_1652);
xnor U748 (N_748,In_521,In_1579);
and U749 (N_749,In_1986,In_1785);
nand U750 (N_750,In_1458,In_48);
xnor U751 (N_751,In_1800,In_329);
or U752 (N_752,In_1512,In_559);
nor U753 (N_753,In_1311,In_1693);
nand U754 (N_754,In_1395,In_1392);
or U755 (N_755,In_69,In_918);
nand U756 (N_756,In_1688,In_178);
nor U757 (N_757,In_130,In_514);
nor U758 (N_758,In_1821,In_144);
or U759 (N_759,In_1335,In_1448);
nor U760 (N_760,In_159,In_1573);
nand U761 (N_761,In_488,In_1425);
xor U762 (N_762,In_1893,In_1250);
xnor U763 (N_763,In_49,In_303);
or U764 (N_764,In_1281,In_572);
nand U765 (N_765,In_1658,In_216);
nand U766 (N_766,In_1589,In_1604);
or U767 (N_767,In_633,In_1371);
xor U768 (N_768,In_950,In_528);
nor U769 (N_769,In_1315,In_890);
nand U770 (N_770,In_1666,In_1776);
nand U771 (N_771,In_91,In_627);
xnor U772 (N_772,In_74,In_195);
nand U773 (N_773,In_726,In_596);
xnor U774 (N_774,In_267,In_769);
nand U775 (N_775,In_672,In_1329);
or U776 (N_776,In_1453,In_952);
nand U777 (N_777,In_869,In_764);
nor U778 (N_778,In_437,In_980);
nand U779 (N_779,In_1897,In_1437);
nor U780 (N_780,In_1937,In_515);
nor U781 (N_781,In_1874,In_509);
xor U782 (N_782,In_1891,In_939);
xnor U783 (N_783,In_27,In_1441);
nor U784 (N_784,In_1209,In_783);
or U785 (N_785,In_755,In_687);
nor U786 (N_786,In_908,In_1255);
and U787 (N_787,In_1752,In_1410);
nor U788 (N_788,In_1714,In_326);
or U789 (N_789,In_172,In_604);
nor U790 (N_790,In_1043,In_609);
nand U791 (N_791,In_739,In_756);
nand U792 (N_792,In_1400,In_1146);
nor U793 (N_793,In_913,In_1297);
or U794 (N_794,In_1841,In_1083);
or U795 (N_795,In_1578,In_641);
nor U796 (N_796,In_1269,In_1121);
nor U797 (N_797,In_1198,In_1708);
and U798 (N_798,In_183,In_1989);
nand U799 (N_799,In_1323,In_1836);
nand U800 (N_800,In_238,In_1145);
nor U801 (N_801,In_991,In_1356);
nand U802 (N_802,In_1795,In_948);
and U803 (N_803,In_170,In_1133);
and U804 (N_804,In_1112,In_1096);
and U805 (N_805,In_87,In_546);
nand U806 (N_806,In_1283,In_1465);
nor U807 (N_807,In_1974,In_167);
and U808 (N_808,In_1066,In_309);
xor U809 (N_809,In_1327,In_67);
nor U810 (N_810,In_1228,In_856);
or U811 (N_811,In_1805,In_813);
or U812 (N_812,In_269,In_185);
and U813 (N_813,In_1069,In_419);
xor U814 (N_814,In_133,In_660);
or U815 (N_815,In_336,In_523);
nor U816 (N_816,In_1128,In_1284);
nand U817 (N_817,In_960,In_1118);
or U818 (N_818,In_910,In_802);
or U819 (N_819,In_752,In_128);
xor U820 (N_820,In_1391,In_1494);
xnor U821 (N_821,In_80,In_237);
nand U822 (N_822,In_28,In_1545);
or U823 (N_823,In_956,In_539);
and U824 (N_824,In_476,In_407);
and U825 (N_825,In_947,In_1200);
nor U826 (N_826,In_1363,In_995);
or U827 (N_827,In_486,In_298);
or U828 (N_828,In_1630,In_927);
xor U829 (N_829,In_1898,In_1249);
and U830 (N_830,In_815,In_1499);
and U831 (N_831,In_328,In_1230);
xor U832 (N_832,In_1838,In_548);
nand U833 (N_833,In_1177,In_1428);
xnor U834 (N_834,In_1351,In_1253);
xor U835 (N_835,In_1388,In_1806);
and U836 (N_836,In_25,In_529);
or U837 (N_837,In_1065,In_1879);
or U838 (N_838,In_1127,In_356);
or U839 (N_839,In_1769,In_451);
nand U840 (N_840,In_1547,In_1562);
nand U841 (N_841,In_343,In_968);
and U842 (N_842,In_1549,In_1068);
xor U843 (N_843,In_644,In_1366);
nand U844 (N_844,In_1975,In_316);
and U845 (N_845,In_1864,In_1557);
or U846 (N_846,In_1725,In_741);
and U847 (N_847,In_1894,In_1033);
or U848 (N_848,In_724,In_1184);
xor U849 (N_849,In_1138,In_983);
nand U850 (N_850,In_1945,In_531);
nor U851 (N_851,In_181,In_125);
xor U852 (N_852,In_226,In_82);
nor U853 (N_853,In_1115,In_656);
or U854 (N_854,In_194,In_1967);
nand U855 (N_855,In_1227,In_137);
and U856 (N_856,In_1739,In_1500);
nand U857 (N_857,In_1532,In_1003);
or U858 (N_858,In_1240,In_348);
or U859 (N_859,In_586,In_852);
nor U860 (N_860,In_2,In_18);
nor U861 (N_861,In_1034,In_754);
xnor U862 (N_862,In_1655,In_114);
nor U863 (N_863,In_256,In_21);
xnor U864 (N_864,In_1493,In_887);
and U865 (N_865,In_464,In_1181);
and U866 (N_866,In_1663,In_1110);
xor U867 (N_867,In_1344,In_787);
nand U868 (N_868,In_1525,In_615);
nor U869 (N_869,In_1480,In_1389);
xor U870 (N_870,In_1625,In_1903);
nor U871 (N_871,In_543,In_731);
and U872 (N_872,In_1511,In_228);
or U873 (N_873,In_613,In_790);
nand U874 (N_874,In_1985,In_725);
nor U875 (N_875,In_179,In_717);
nand U876 (N_876,In_1777,In_340);
nand U877 (N_877,In_930,In_426);
nand U878 (N_878,In_207,In_1936);
or U879 (N_879,In_870,In_1081);
xnor U880 (N_880,In_100,In_1925);
xnor U881 (N_881,In_1624,In_1373);
nand U882 (N_882,In_1423,In_883);
or U883 (N_883,In_1870,In_542);
or U884 (N_884,In_1479,In_623);
or U885 (N_885,In_63,In_1298);
and U886 (N_886,In_1190,In_570);
nand U887 (N_887,In_136,In_1567);
xnor U888 (N_888,In_1732,In_171);
and U889 (N_889,In_740,In_1593);
or U890 (N_890,In_640,In_1533);
or U891 (N_891,In_617,In_1966);
nand U892 (N_892,In_1090,In_779);
and U893 (N_893,In_1823,In_603);
nor U894 (N_894,In_1079,In_1719);
nand U895 (N_895,In_463,In_826);
nor U896 (N_896,In_1139,In_501);
nand U897 (N_897,In_1411,In_1513);
and U898 (N_898,In_1211,In_1263);
xor U899 (N_899,In_807,In_1473);
or U900 (N_900,In_1244,In_579);
xnor U901 (N_901,In_1905,In_1326);
nor U902 (N_902,In_1322,In_255);
and U903 (N_903,In_7,In_338);
and U904 (N_904,In_1075,In_1669);
and U905 (N_905,In_697,In_561);
nor U906 (N_906,In_1941,In_836);
xor U907 (N_907,In_1926,In_290);
nor U908 (N_908,In_1710,In_679);
nor U909 (N_909,In_1182,In_1840);
nor U910 (N_910,In_1835,In_1815);
xor U911 (N_911,In_1390,In_1252);
or U912 (N_912,In_1726,In_1225);
nand U913 (N_913,In_1724,In_32);
and U914 (N_914,In_446,In_390);
nand U915 (N_915,In_1029,In_1449);
nor U916 (N_916,In_976,In_763);
nand U917 (N_917,In_1887,In_1231);
and U918 (N_918,In_563,In_1671);
and U919 (N_919,In_1132,In_1554);
and U920 (N_920,In_1204,In_1258);
and U921 (N_921,In_241,In_75);
nand U922 (N_922,In_398,In_541);
nand U923 (N_923,In_447,In_494);
nand U924 (N_924,In_1820,In_876);
nand U925 (N_925,In_630,In_901);
nor U926 (N_926,In_42,In_246);
xnor U927 (N_927,In_254,In_1774);
or U928 (N_928,In_1,In_1199);
and U929 (N_929,In_59,In_841);
nor U930 (N_930,In_295,In_1783);
nor U931 (N_931,In_1440,In_589);
or U932 (N_932,In_1860,In_1948);
or U933 (N_933,In_421,In_610);
nand U934 (N_934,In_696,In_1943);
nand U935 (N_935,In_475,In_1534);
or U936 (N_936,In_1266,In_1301);
or U937 (N_937,In_1713,In_1030);
xor U938 (N_938,In_718,In_352);
or U939 (N_939,In_606,In_1680);
or U940 (N_940,In_1944,In_1313);
nand U941 (N_941,In_1988,In_861);
and U942 (N_942,In_814,In_68);
and U943 (N_943,In_573,In_882);
xnor U944 (N_944,In_122,In_635);
nand U945 (N_945,In_593,In_1495);
nor U946 (N_946,In_1952,In_864);
nand U947 (N_947,In_455,In_1818);
xor U948 (N_948,In_1111,In_243);
nand U949 (N_949,In_1911,In_1095);
and U950 (N_950,In_467,In_1828);
or U951 (N_951,In_417,In_121);
or U952 (N_952,In_674,In_1742);
and U953 (N_953,In_1468,In_1101);
or U954 (N_954,In_742,In_1938);
and U955 (N_955,In_775,In_1568);
and U956 (N_956,In_862,In_1706);
nor U957 (N_957,In_482,In_8);
and U958 (N_958,In_961,In_868);
and U959 (N_959,In_93,In_1158);
or U960 (N_960,In_1235,In_938);
nand U961 (N_961,In_1983,In_1466);
or U962 (N_962,In_140,In_662);
nand U963 (N_963,In_777,In_536);
or U964 (N_964,In_481,In_95);
nand U965 (N_965,In_1191,In_1215);
nand U966 (N_966,In_249,In_1443);
nand U967 (N_967,In_705,In_1024);
nor U968 (N_968,In_1933,In_1951);
and U969 (N_969,In_986,In_1844);
nand U970 (N_970,In_1290,In_472);
and U971 (N_971,In_1660,In_809);
xor U972 (N_972,In_794,In_768);
and U973 (N_973,In_1272,In_157);
nand U974 (N_974,In_1852,In_77);
or U975 (N_975,In_393,In_1932);
xnor U976 (N_976,In_577,In_1825);
nor U977 (N_977,In_1226,In_1629);
or U978 (N_978,In_1973,In_46);
xnor U979 (N_979,In_1038,In_302);
or U980 (N_980,In_454,In_1147);
or U981 (N_981,In_385,In_395);
nand U982 (N_982,In_111,In_1626);
nand U983 (N_983,In_327,In_767);
nand U984 (N_984,In_1124,In_477);
nor U985 (N_985,In_540,In_958);
and U986 (N_986,In_55,In_427);
and U987 (N_987,In_1224,In_1560);
nand U988 (N_988,In_1109,In_743);
nor U989 (N_989,In_66,In_1058);
nor U990 (N_990,In_721,In_1613);
nand U991 (N_991,In_173,In_550);
or U992 (N_992,In_120,In_1359);
xnor U993 (N_993,In_1372,In_945);
or U994 (N_994,In_480,In_1697);
nor U995 (N_995,In_1349,In_1439);
and U996 (N_996,In_1463,In_1082);
nand U997 (N_997,In_1378,In_1017);
or U998 (N_998,In_1632,In_1987);
and U999 (N_999,In_689,In_1729);
nand U1000 (N_1000,In_461,In_1083);
nand U1001 (N_1001,In_357,In_1305);
xnor U1002 (N_1002,In_1035,In_814);
or U1003 (N_1003,In_1089,In_348);
or U1004 (N_1004,In_499,In_664);
nor U1005 (N_1005,In_1227,In_1373);
and U1006 (N_1006,In_259,In_46);
xor U1007 (N_1007,In_664,In_1160);
nor U1008 (N_1008,In_339,In_1543);
and U1009 (N_1009,In_1884,In_1621);
or U1010 (N_1010,In_1626,In_117);
and U1011 (N_1011,In_1732,In_1414);
or U1012 (N_1012,In_171,In_1182);
nand U1013 (N_1013,In_1057,In_1265);
and U1014 (N_1014,In_421,In_1591);
nand U1015 (N_1015,In_524,In_107);
or U1016 (N_1016,In_166,In_1770);
nand U1017 (N_1017,In_745,In_1158);
nor U1018 (N_1018,In_1323,In_810);
or U1019 (N_1019,In_337,In_1778);
and U1020 (N_1020,In_854,In_1637);
nand U1021 (N_1021,In_1291,In_709);
nand U1022 (N_1022,In_1608,In_404);
nand U1023 (N_1023,In_484,In_20);
and U1024 (N_1024,In_497,In_59);
xnor U1025 (N_1025,In_311,In_1864);
nand U1026 (N_1026,In_1893,In_1541);
xor U1027 (N_1027,In_1743,In_1985);
or U1028 (N_1028,In_16,In_463);
or U1029 (N_1029,In_1284,In_1746);
xor U1030 (N_1030,In_1259,In_1954);
xor U1031 (N_1031,In_1853,In_1817);
xnor U1032 (N_1032,In_1778,In_518);
and U1033 (N_1033,In_704,In_1781);
and U1034 (N_1034,In_821,In_1513);
nand U1035 (N_1035,In_1534,In_628);
or U1036 (N_1036,In_663,In_73);
and U1037 (N_1037,In_551,In_169);
or U1038 (N_1038,In_235,In_1976);
nor U1039 (N_1039,In_14,In_1220);
nor U1040 (N_1040,In_1763,In_1654);
nand U1041 (N_1041,In_429,In_869);
and U1042 (N_1042,In_1053,In_1379);
nor U1043 (N_1043,In_1701,In_926);
nand U1044 (N_1044,In_1003,In_267);
and U1045 (N_1045,In_862,In_1521);
and U1046 (N_1046,In_1214,In_1409);
nor U1047 (N_1047,In_1301,In_1606);
and U1048 (N_1048,In_796,In_1700);
nand U1049 (N_1049,In_1731,In_1328);
or U1050 (N_1050,In_1657,In_928);
xor U1051 (N_1051,In_878,In_1516);
nor U1052 (N_1052,In_1013,In_1463);
or U1053 (N_1053,In_174,In_1223);
or U1054 (N_1054,In_1789,In_216);
nand U1055 (N_1055,In_1581,In_1022);
nor U1056 (N_1056,In_930,In_42);
or U1057 (N_1057,In_143,In_1624);
or U1058 (N_1058,In_963,In_1239);
nand U1059 (N_1059,In_1046,In_129);
xor U1060 (N_1060,In_196,In_77);
nor U1061 (N_1061,In_1264,In_1302);
and U1062 (N_1062,In_1033,In_1849);
nand U1063 (N_1063,In_289,In_994);
nand U1064 (N_1064,In_527,In_1363);
nand U1065 (N_1065,In_845,In_1317);
or U1066 (N_1066,In_292,In_1081);
or U1067 (N_1067,In_1424,In_971);
nand U1068 (N_1068,In_155,In_744);
and U1069 (N_1069,In_477,In_52);
xor U1070 (N_1070,In_327,In_1777);
nand U1071 (N_1071,In_1138,In_558);
and U1072 (N_1072,In_1037,In_1005);
nand U1073 (N_1073,In_1648,In_525);
nor U1074 (N_1074,In_782,In_813);
xor U1075 (N_1075,In_385,In_696);
and U1076 (N_1076,In_558,In_446);
and U1077 (N_1077,In_1857,In_364);
and U1078 (N_1078,In_183,In_896);
and U1079 (N_1079,In_1857,In_1790);
xor U1080 (N_1080,In_1821,In_517);
nand U1081 (N_1081,In_1666,In_1318);
xor U1082 (N_1082,In_1469,In_247);
nor U1083 (N_1083,In_1201,In_1542);
xor U1084 (N_1084,In_1045,In_1065);
or U1085 (N_1085,In_477,In_1606);
and U1086 (N_1086,In_493,In_923);
and U1087 (N_1087,In_1706,In_1737);
or U1088 (N_1088,In_1378,In_269);
or U1089 (N_1089,In_1735,In_1517);
or U1090 (N_1090,In_1592,In_1967);
nor U1091 (N_1091,In_1571,In_1499);
or U1092 (N_1092,In_1472,In_1279);
xnor U1093 (N_1093,In_983,In_883);
nand U1094 (N_1094,In_800,In_1377);
nand U1095 (N_1095,In_458,In_1373);
nand U1096 (N_1096,In_28,In_482);
xnor U1097 (N_1097,In_245,In_818);
and U1098 (N_1098,In_1680,In_617);
xnor U1099 (N_1099,In_229,In_1990);
nor U1100 (N_1100,In_579,In_362);
or U1101 (N_1101,In_1745,In_475);
nand U1102 (N_1102,In_874,In_1090);
nand U1103 (N_1103,In_1480,In_175);
xnor U1104 (N_1104,In_632,In_345);
nor U1105 (N_1105,In_1495,In_1349);
nand U1106 (N_1106,In_377,In_1989);
nand U1107 (N_1107,In_668,In_1261);
or U1108 (N_1108,In_665,In_386);
nand U1109 (N_1109,In_437,In_25);
xor U1110 (N_1110,In_1625,In_1134);
and U1111 (N_1111,In_657,In_800);
and U1112 (N_1112,In_1177,In_929);
xnor U1113 (N_1113,In_306,In_945);
or U1114 (N_1114,In_1578,In_1463);
nor U1115 (N_1115,In_425,In_1542);
nor U1116 (N_1116,In_601,In_1378);
or U1117 (N_1117,In_425,In_1410);
xor U1118 (N_1118,In_1065,In_503);
and U1119 (N_1119,In_1054,In_756);
nand U1120 (N_1120,In_81,In_1263);
nor U1121 (N_1121,In_616,In_8);
xnor U1122 (N_1122,In_1140,In_4);
nor U1123 (N_1123,In_891,In_768);
xor U1124 (N_1124,In_520,In_1471);
xor U1125 (N_1125,In_246,In_347);
xor U1126 (N_1126,In_912,In_1809);
nand U1127 (N_1127,In_400,In_1170);
nand U1128 (N_1128,In_1796,In_1116);
and U1129 (N_1129,In_1998,In_1530);
or U1130 (N_1130,In_402,In_1659);
and U1131 (N_1131,In_845,In_110);
xor U1132 (N_1132,In_330,In_1545);
and U1133 (N_1133,In_561,In_445);
nor U1134 (N_1134,In_962,In_1497);
xor U1135 (N_1135,In_1606,In_187);
or U1136 (N_1136,In_1970,In_479);
nor U1137 (N_1137,In_922,In_139);
nand U1138 (N_1138,In_792,In_1826);
nand U1139 (N_1139,In_1078,In_1937);
xor U1140 (N_1140,In_213,In_1836);
xor U1141 (N_1141,In_459,In_1431);
or U1142 (N_1142,In_1724,In_1009);
xor U1143 (N_1143,In_228,In_1116);
xnor U1144 (N_1144,In_1067,In_325);
nand U1145 (N_1145,In_1298,In_386);
and U1146 (N_1146,In_1578,In_1731);
xnor U1147 (N_1147,In_1787,In_1587);
xor U1148 (N_1148,In_1407,In_1486);
nor U1149 (N_1149,In_1394,In_1440);
xnor U1150 (N_1150,In_993,In_1717);
or U1151 (N_1151,In_1047,In_1305);
or U1152 (N_1152,In_1890,In_244);
nand U1153 (N_1153,In_48,In_940);
nor U1154 (N_1154,In_1981,In_390);
nor U1155 (N_1155,In_1466,In_1217);
nand U1156 (N_1156,In_1879,In_1840);
and U1157 (N_1157,In_646,In_773);
nor U1158 (N_1158,In_196,In_300);
and U1159 (N_1159,In_176,In_1298);
nor U1160 (N_1160,In_631,In_1323);
nand U1161 (N_1161,In_1530,In_1031);
nor U1162 (N_1162,In_748,In_72);
or U1163 (N_1163,In_1738,In_299);
and U1164 (N_1164,In_552,In_266);
xor U1165 (N_1165,In_972,In_1616);
xnor U1166 (N_1166,In_1588,In_623);
nand U1167 (N_1167,In_737,In_1047);
and U1168 (N_1168,In_726,In_612);
or U1169 (N_1169,In_423,In_1599);
nor U1170 (N_1170,In_522,In_1774);
nand U1171 (N_1171,In_378,In_1066);
or U1172 (N_1172,In_519,In_186);
or U1173 (N_1173,In_1856,In_404);
or U1174 (N_1174,In_445,In_1213);
nor U1175 (N_1175,In_797,In_683);
nand U1176 (N_1176,In_1464,In_596);
nor U1177 (N_1177,In_365,In_744);
and U1178 (N_1178,In_1219,In_1046);
and U1179 (N_1179,In_1701,In_1134);
nor U1180 (N_1180,In_679,In_138);
or U1181 (N_1181,In_641,In_1289);
nor U1182 (N_1182,In_13,In_908);
nand U1183 (N_1183,In_1067,In_1167);
xnor U1184 (N_1184,In_1994,In_787);
or U1185 (N_1185,In_300,In_1061);
xnor U1186 (N_1186,In_144,In_1492);
xor U1187 (N_1187,In_375,In_829);
nor U1188 (N_1188,In_1941,In_1656);
xnor U1189 (N_1189,In_50,In_390);
xnor U1190 (N_1190,In_958,In_1795);
nor U1191 (N_1191,In_891,In_1761);
nor U1192 (N_1192,In_580,In_132);
nor U1193 (N_1193,In_473,In_1060);
xnor U1194 (N_1194,In_989,In_142);
xor U1195 (N_1195,In_1029,In_1987);
nor U1196 (N_1196,In_1546,In_229);
xnor U1197 (N_1197,In_1366,In_1220);
and U1198 (N_1198,In_1696,In_862);
or U1199 (N_1199,In_2,In_1987);
and U1200 (N_1200,In_486,In_356);
nand U1201 (N_1201,In_729,In_1099);
nor U1202 (N_1202,In_1786,In_145);
and U1203 (N_1203,In_1313,In_165);
and U1204 (N_1204,In_1457,In_390);
nand U1205 (N_1205,In_1940,In_476);
and U1206 (N_1206,In_338,In_1448);
nor U1207 (N_1207,In_1083,In_512);
and U1208 (N_1208,In_601,In_1227);
and U1209 (N_1209,In_1420,In_1338);
xnor U1210 (N_1210,In_1773,In_1300);
and U1211 (N_1211,In_114,In_1467);
nor U1212 (N_1212,In_679,In_847);
or U1213 (N_1213,In_610,In_988);
or U1214 (N_1214,In_1456,In_176);
nand U1215 (N_1215,In_1242,In_1103);
xor U1216 (N_1216,In_97,In_1368);
or U1217 (N_1217,In_1552,In_721);
or U1218 (N_1218,In_1080,In_1067);
nor U1219 (N_1219,In_486,In_1094);
nor U1220 (N_1220,In_1588,In_1628);
and U1221 (N_1221,In_739,In_37);
and U1222 (N_1222,In_398,In_191);
and U1223 (N_1223,In_1386,In_318);
or U1224 (N_1224,In_1773,In_1660);
nand U1225 (N_1225,In_437,In_890);
xnor U1226 (N_1226,In_1478,In_1521);
nand U1227 (N_1227,In_248,In_1281);
and U1228 (N_1228,In_988,In_1026);
nand U1229 (N_1229,In_1976,In_284);
nand U1230 (N_1230,In_1299,In_470);
and U1231 (N_1231,In_244,In_1196);
nor U1232 (N_1232,In_657,In_446);
nand U1233 (N_1233,In_523,In_365);
or U1234 (N_1234,In_853,In_691);
or U1235 (N_1235,In_1688,In_644);
nor U1236 (N_1236,In_1697,In_1500);
xnor U1237 (N_1237,In_1512,In_2);
and U1238 (N_1238,In_394,In_376);
and U1239 (N_1239,In_50,In_499);
or U1240 (N_1240,In_68,In_178);
nor U1241 (N_1241,In_749,In_983);
nand U1242 (N_1242,In_1186,In_248);
xor U1243 (N_1243,In_515,In_1896);
nor U1244 (N_1244,In_822,In_1203);
xor U1245 (N_1245,In_403,In_251);
xnor U1246 (N_1246,In_510,In_134);
nand U1247 (N_1247,In_296,In_279);
xor U1248 (N_1248,In_1838,In_1226);
or U1249 (N_1249,In_1375,In_1934);
or U1250 (N_1250,In_1484,In_978);
and U1251 (N_1251,In_1659,In_351);
xor U1252 (N_1252,In_796,In_1074);
nand U1253 (N_1253,In_523,In_693);
nand U1254 (N_1254,In_1570,In_251);
xnor U1255 (N_1255,In_1899,In_1078);
and U1256 (N_1256,In_1439,In_958);
and U1257 (N_1257,In_497,In_96);
or U1258 (N_1258,In_8,In_620);
nand U1259 (N_1259,In_1669,In_1203);
and U1260 (N_1260,In_306,In_1500);
nor U1261 (N_1261,In_1771,In_1216);
nor U1262 (N_1262,In_994,In_838);
xnor U1263 (N_1263,In_392,In_109);
nor U1264 (N_1264,In_355,In_1994);
xnor U1265 (N_1265,In_1222,In_1872);
nand U1266 (N_1266,In_1665,In_1081);
nand U1267 (N_1267,In_503,In_1438);
xor U1268 (N_1268,In_771,In_654);
xor U1269 (N_1269,In_1017,In_1476);
or U1270 (N_1270,In_1519,In_1036);
nor U1271 (N_1271,In_720,In_1325);
or U1272 (N_1272,In_1950,In_306);
and U1273 (N_1273,In_348,In_238);
nand U1274 (N_1274,In_1324,In_1582);
nand U1275 (N_1275,In_1454,In_667);
or U1276 (N_1276,In_1328,In_307);
nand U1277 (N_1277,In_1712,In_1154);
or U1278 (N_1278,In_106,In_59);
and U1279 (N_1279,In_786,In_24);
or U1280 (N_1280,In_1450,In_1618);
or U1281 (N_1281,In_72,In_101);
nand U1282 (N_1282,In_1991,In_685);
nor U1283 (N_1283,In_690,In_1693);
nor U1284 (N_1284,In_995,In_444);
xor U1285 (N_1285,In_200,In_454);
nand U1286 (N_1286,In_236,In_1961);
and U1287 (N_1287,In_1010,In_1541);
xor U1288 (N_1288,In_552,In_380);
nand U1289 (N_1289,In_727,In_1585);
nor U1290 (N_1290,In_663,In_1601);
or U1291 (N_1291,In_852,In_1539);
and U1292 (N_1292,In_724,In_1243);
nor U1293 (N_1293,In_1248,In_331);
nand U1294 (N_1294,In_1177,In_1376);
xnor U1295 (N_1295,In_289,In_621);
and U1296 (N_1296,In_1830,In_683);
nor U1297 (N_1297,In_1167,In_786);
and U1298 (N_1298,In_1974,In_1961);
and U1299 (N_1299,In_95,In_633);
and U1300 (N_1300,In_190,In_1847);
nand U1301 (N_1301,In_847,In_1419);
nor U1302 (N_1302,In_1436,In_950);
xnor U1303 (N_1303,In_1388,In_1152);
xnor U1304 (N_1304,In_1552,In_236);
and U1305 (N_1305,In_849,In_1243);
and U1306 (N_1306,In_575,In_1803);
nand U1307 (N_1307,In_1739,In_594);
or U1308 (N_1308,In_1459,In_1180);
or U1309 (N_1309,In_427,In_113);
nor U1310 (N_1310,In_787,In_1099);
nand U1311 (N_1311,In_508,In_992);
and U1312 (N_1312,In_176,In_1092);
xnor U1313 (N_1313,In_1784,In_826);
nor U1314 (N_1314,In_411,In_1223);
and U1315 (N_1315,In_356,In_551);
and U1316 (N_1316,In_1890,In_1730);
nand U1317 (N_1317,In_1146,In_800);
nor U1318 (N_1318,In_942,In_1754);
xor U1319 (N_1319,In_1979,In_353);
nor U1320 (N_1320,In_250,In_839);
and U1321 (N_1321,In_940,In_149);
nor U1322 (N_1322,In_1893,In_1906);
and U1323 (N_1323,In_1917,In_116);
nor U1324 (N_1324,In_1205,In_1751);
and U1325 (N_1325,In_804,In_569);
and U1326 (N_1326,In_188,In_1252);
or U1327 (N_1327,In_140,In_8);
xnor U1328 (N_1328,In_1169,In_787);
nand U1329 (N_1329,In_313,In_1623);
or U1330 (N_1330,In_1228,In_450);
nand U1331 (N_1331,In_663,In_337);
nand U1332 (N_1332,In_1915,In_178);
nor U1333 (N_1333,In_445,In_70);
or U1334 (N_1334,In_346,In_1829);
nand U1335 (N_1335,In_1816,In_472);
nand U1336 (N_1336,In_670,In_1177);
or U1337 (N_1337,In_1241,In_608);
nand U1338 (N_1338,In_651,In_491);
nor U1339 (N_1339,In_1904,In_1754);
and U1340 (N_1340,In_1999,In_25);
or U1341 (N_1341,In_1034,In_1170);
or U1342 (N_1342,In_164,In_214);
nor U1343 (N_1343,In_39,In_201);
and U1344 (N_1344,In_749,In_1759);
nand U1345 (N_1345,In_1094,In_626);
nand U1346 (N_1346,In_858,In_547);
or U1347 (N_1347,In_1702,In_317);
xor U1348 (N_1348,In_1017,In_994);
and U1349 (N_1349,In_1908,In_771);
nor U1350 (N_1350,In_48,In_426);
nand U1351 (N_1351,In_1861,In_485);
and U1352 (N_1352,In_895,In_1253);
nor U1353 (N_1353,In_1210,In_783);
and U1354 (N_1354,In_1852,In_804);
or U1355 (N_1355,In_796,In_412);
xor U1356 (N_1356,In_627,In_1077);
nor U1357 (N_1357,In_629,In_1272);
xor U1358 (N_1358,In_590,In_845);
xnor U1359 (N_1359,In_1367,In_1677);
or U1360 (N_1360,In_107,In_1132);
xor U1361 (N_1361,In_1981,In_951);
nand U1362 (N_1362,In_333,In_179);
xor U1363 (N_1363,In_676,In_501);
nor U1364 (N_1364,In_718,In_1521);
xnor U1365 (N_1365,In_51,In_53);
nor U1366 (N_1366,In_1962,In_267);
xor U1367 (N_1367,In_698,In_609);
and U1368 (N_1368,In_1629,In_1130);
xor U1369 (N_1369,In_627,In_1829);
nor U1370 (N_1370,In_1806,In_440);
xnor U1371 (N_1371,In_442,In_482);
xnor U1372 (N_1372,In_992,In_1622);
or U1373 (N_1373,In_1619,In_1260);
xor U1374 (N_1374,In_1095,In_1276);
nand U1375 (N_1375,In_1931,In_564);
nor U1376 (N_1376,In_235,In_1977);
and U1377 (N_1377,In_1982,In_131);
nor U1378 (N_1378,In_733,In_1400);
nor U1379 (N_1379,In_1398,In_1427);
and U1380 (N_1380,In_736,In_1240);
xor U1381 (N_1381,In_1554,In_1122);
nor U1382 (N_1382,In_1814,In_1678);
nor U1383 (N_1383,In_1542,In_1066);
nand U1384 (N_1384,In_863,In_1480);
xor U1385 (N_1385,In_108,In_971);
xor U1386 (N_1386,In_461,In_622);
and U1387 (N_1387,In_185,In_591);
or U1388 (N_1388,In_1143,In_1561);
xor U1389 (N_1389,In_1099,In_1270);
and U1390 (N_1390,In_1508,In_898);
and U1391 (N_1391,In_164,In_492);
xnor U1392 (N_1392,In_1306,In_1424);
nand U1393 (N_1393,In_1775,In_206);
nor U1394 (N_1394,In_726,In_51);
or U1395 (N_1395,In_1368,In_82);
nor U1396 (N_1396,In_697,In_850);
or U1397 (N_1397,In_147,In_1997);
nand U1398 (N_1398,In_277,In_1247);
xnor U1399 (N_1399,In_1674,In_1556);
nor U1400 (N_1400,In_655,In_1232);
and U1401 (N_1401,In_285,In_1292);
nand U1402 (N_1402,In_1005,In_116);
or U1403 (N_1403,In_1400,In_531);
and U1404 (N_1404,In_376,In_192);
xor U1405 (N_1405,In_136,In_1716);
or U1406 (N_1406,In_1212,In_1982);
nor U1407 (N_1407,In_726,In_1905);
xor U1408 (N_1408,In_187,In_806);
xnor U1409 (N_1409,In_1418,In_1391);
or U1410 (N_1410,In_327,In_1183);
and U1411 (N_1411,In_533,In_1173);
nand U1412 (N_1412,In_952,In_508);
nand U1413 (N_1413,In_140,In_1600);
nand U1414 (N_1414,In_348,In_1540);
nor U1415 (N_1415,In_1159,In_221);
and U1416 (N_1416,In_1363,In_1301);
nand U1417 (N_1417,In_1413,In_1937);
xnor U1418 (N_1418,In_886,In_294);
nor U1419 (N_1419,In_1898,In_1073);
and U1420 (N_1420,In_1227,In_1506);
and U1421 (N_1421,In_1674,In_1259);
xnor U1422 (N_1422,In_1258,In_1038);
xnor U1423 (N_1423,In_1673,In_1571);
xnor U1424 (N_1424,In_26,In_576);
or U1425 (N_1425,In_1456,In_981);
xor U1426 (N_1426,In_327,In_796);
nor U1427 (N_1427,In_1575,In_424);
nor U1428 (N_1428,In_1234,In_1573);
nor U1429 (N_1429,In_557,In_1197);
and U1430 (N_1430,In_1169,In_1380);
or U1431 (N_1431,In_1272,In_585);
and U1432 (N_1432,In_1641,In_1261);
nor U1433 (N_1433,In_405,In_1202);
nor U1434 (N_1434,In_1406,In_361);
xor U1435 (N_1435,In_103,In_1729);
xor U1436 (N_1436,In_63,In_1507);
xor U1437 (N_1437,In_926,In_1128);
nand U1438 (N_1438,In_706,In_1960);
nor U1439 (N_1439,In_1137,In_123);
xor U1440 (N_1440,In_76,In_1811);
xor U1441 (N_1441,In_602,In_145);
or U1442 (N_1442,In_1930,In_808);
nor U1443 (N_1443,In_775,In_866);
xnor U1444 (N_1444,In_757,In_1809);
and U1445 (N_1445,In_1584,In_1375);
or U1446 (N_1446,In_930,In_201);
and U1447 (N_1447,In_189,In_226);
nor U1448 (N_1448,In_774,In_1733);
or U1449 (N_1449,In_1103,In_47);
and U1450 (N_1450,In_15,In_1131);
xnor U1451 (N_1451,In_839,In_1975);
and U1452 (N_1452,In_21,In_1898);
xor U1453 (N_1453,In_1543,In_1014);
nand U1454 (N_1454,In_1174,In_965);
nand U1455 (N_1455,In_1912,In_1938);
and U1456 (N_1456,In_1480,In_684);
or U1457 (N_1457,In_1759,In_1418);
nand U1458 (N_1458,In_926,In_1210);
or U1459 (N_1459,In_1641,In_972);
nor U1460 (N_1460,In_1460,In_1682);
or U1461 (N_1461,In_1818,In_1775);
nor U1462 (N_1462,In_1098,In_1246);
or U1463 (N_1463,In_890,In_668);
nand U1464 (N_1464,In_1459,In_288);
or U1465 (N_1465,In_360,In_307);
or U1466 (N_1466,In_14,In_1675);
xnor U1467 (N_1467,In_1449,In_1374);
nor U1468 (N_1468,In_1570,In_1450);
nor U1469 (N_1469,In_1086,In_1534);
or U1470 (N_1470,In_1304,In_361);
nor U1471 (N_1471,In_658,In_682);
xor U1472 (N_1472,In_745,In_958);
nand U1473 (N_1473,In_1392,In_639);
xor U1474 (N_1474,In_1735,In_1758);
nor U1475 (N_1475,In_585,In_1550);
and U1476 (N_1476,In_1302,In_675);
xor U1477 (N_1477,In_648,In_1004);
nor U1478 (N_1478,In_1602,In_956);
xor U1479 (N_1479,In_1206,In_382);
nand U1480 (N_1480,In_1058,In_1109);
xnor U1481 (N_1481,In_916,In_1929);
xor U1482 (N_1482,In_589,In_615);
and U1483 (N_1483,In_145,In_1599);
or U1484 (N_1484,In_1094,In_1059);
nand U1485 (N_1485,In_169,In_115);
nor U1486 (N_1486,In_1557,In_293);
or U1487 (N_1487,In_310,In_113);
and U1488 (N_1488,In_1785,In_494);
and U1489 (N_1489,In_222,In_442);
and U1490 (N_1490,In_1735,In_882);
and U1491 (N_1491,In_1512,In_929);
nor U1492 (N_1492,In_1886,In_936);
nor U1493 (N_1493,In_1242,In_1957);
xor U1494 (N_1494,In_1561,In_417);
nand U1495 (N_1495,In_1070,In_246);
or U1496 (N_1496,In_946,In_655);
nand U1497 (N_1497,In_1933,In_339);
and U1498 (N_1498,In_178,In_56);
nand U1499 (N_1499,In_631,In_1249);
xnor U1500 (N_1500,In_14,In_895);
xnor U1501 (N_1501,In_598,In_1268);
or U1502 (N_1502,In_1927,In_1032);
nand U1503 (N_1503,In_8,In_958);
and U1504 (N_1504,In_1324,In_13);
xor U1505 (N_1505,In_1478,In_575);
and U1506 (N_1506,In_1678,In_45);
or U1507 (N_1507,In_1039,In_1561);
xnor U1508 (N_1508,In_583,In_535);
and U1509 (N_1509,In_274,In_1933);
and U1510 (N_1510,In_1725,In_1492);
and U1511 (N_1511,In_1942,In_153);
xor U1512 (N_1512,In_391,In_1069);
nor U1513 (N_1513,In_1269,In_1763);
xor U1514 (N_1514,In_1543,In_1062);
and U1515 (N_1515,In_278,In_1592);
or U1516 (N_1516,In_1659,In_1673);
nor U1517 (N_1517,In_1671,In_567);
or U1518 (N_1518,In_1083,In_1539);
or U1519 (N_1519,In_1523,In_1986);
or U1520 (N_1520,In_1395,In_804);
and U1521 (N_1521,In_1333,In_718);
and U1522 (N_1522,In_834,In_1180);
and U1523 (N_1523,In_1380,In_1067);
xnor U1524 (N_1524,In_1860,In_1621);
or U1525 (N_1525,In_1011,In_166);
xnor U1526 (N_1526,In_1293,In_207);
and U1527 (N_1527,In_432,In_485);
xor U1528 (N_1528,In_916,In_684);
and U1529 (N_1529,In_1283,In_375);
nor U1530 (N_1530,In_138,In_556);
nor U1531 (N_1531,In_1113,In_966);
xor U1532 (N_1532,In_1481,In_1527);
nor U1533 (N_1533,In_822,In_1517);
xnor U1534 (N_1534,In_1585,In_1573);
xor U1535 (N_1535,In_185,In_679);
or U1536 (N_1536,In_102,In_1373);
or U1537 (N_1537,In_576,In_1084);
xor U1538 (N_1538,In_355,In_1695);
nor U1539 (N_1539,In_1154,In_1529);
xnor U1540 (N_1540,In_1111,In_1371);
xnor U1541 (N_1541,In_854,In_515);
nand U1542 (N_1542,In_1322,In_1536);
xnor U1543 (N_1543,In_400,In_28);
xnor U1544 (N_1544,In_1430,In_1259);
nor U1545 (N_1545,In_1799,In_1079);
or U1546 (N_1546,In_1142,In_1593);
nor U1547 (N_1547,In_697,In_547);
or U1548 (N_1548,In_1348,In_127);
or U1549 (N_1549,In_749,In_803);
xor U1550 (N_1550,In_1273,In_1857);
or U1551 (N_1551,In_92,In_479);
or U1552 (N_1552,In_806,In_1507);
or U1553 (N_1553,In_1557,In_249);
xor U1554 (N_1554,In_631,In_574);
xor U1555 (N_1555,In_1234,In_1192);
and U1556 (N_1556,In_906,In_1823);
nand U1557 (N_1557,In_1631,In_1672);
or U1558 (N_1558,In_1159,In_663);
nor U1559 (N_1559,In_745,In_206);
and U1560 (N_1560,In_726,In_1377);
or U1561 (N_1561,In_1939,In_1560);
and U1562 (N_1562,In_1814,In_978);
and U1563 (N_1563,In_901,In_451);
nand U1564 (N_1564,In_801,In_1777);
xnor U1565 (N_1565,In_1576,In_39);
or U1566 (N_1566,In_1173,In_780);
nor U1567 (N_1567,In_1697,In_436);
nor U1568 (N_1568,In_1540,In_507);
or U1569 (N_1569,In_1405,In_641);
or U1570 (N_1570,In_1122,In_1989);
or U1571 (N_1571,In_1348,In_310);
nand U1572 (N_1572,In_1129,In_772);
nand U1573 (N_1573,In_276,In_1512);
or U1574 (N_1574,In_1591,In_1700);
nor U1575 (N_1575,In_87,In_520);
nor U1576 (N_1576,In_1915,In_1531);
nand U1577 (N_1577,In_202,In_1705);
and U1578 (N_1578,In_1812,In_272);
and U1579 (N_1579,In_933,In_101);
nor U1580 (N_1580,In_1520,In_954);
or U1581 (N_1581,In_1789,In_980);
nand U1582 (N_1582,In_791,In_1968);
nor U1583 (N_1583,In_1283,In_280);
xor U1584 (N_1584,In_1271,In_643);
nand U1585 (N_1585,In_802,In_268);
or U1586 (N_1586,In_574,In_700);
or U1587 (N_1587,In_549,In_941);
xor U1588 (N_1588,In_994,In_1536);
nand U1589 (N_1589,In_1536,In_1033);
and U1590 (N_1590,In_1040,In_726);
nor U1591 (N_1591,In_1734,In_599);
xnor U1592 (N_1592,In_706,In_1733);
xor U1593 (N_1593,In_1495,In_1895);
and U1594 (N_1594,In_1344,In_200);
xnor U1595 (N_1595,In_1277,In_893);
xnor U1596 (N_1596,In_102,In_1582);
or U1597 (N_1597,In_353,In_308);
nor U1598 (N_1598,In_1573,In_1112);
and U1599 (N_1599,In_1656,In_1766);
and U1600 (N_1600,In_1654,In_620);
or U1601 (N_1601,In_834,In_961);
and U1602 (N_1602,In_661,In_480);
or U1603 (N_1603,In_1466,In_110);
or U1604 (N_1604,In_1769,In_1262);
nand U1605 (N_1605,In_876,In_1749);
and U1606 (N_1606,In_466,In_1921);
or U1607 (N_1607,In_12,In_1819);
nor U1608 (N_1608,In_317,In_1227);
nand U1609 (N_1609,In_1354,In_899);
or U1610 (N_1610,In_1951,In_1780);
nor U1611 (N_1611,In_1583,In_1413);
xnor U1612 (N_1612,In_1887,In_1546);
nor U1613 (N_1613,In_1808,In_1968);
xor U1614 (N_1614,In_1581,In_1595);
nor U1615 (N_1615,In_1467,In_744);
or U1616 (N_1616,In_1329,In_1238);
xor U1617 (N_1617,In_1169,In_1106);
nand U1618 (N_1618,In_739,In_117);
or U1619 (N_1619,In_473,In_70);
and U1620 (N_1620,In_1596,In_463);
nor U1621 (N_1621,In_140,In_431);
or U1622 (N_1622,In_609,In_1342);
or U1623 (N_1623,In_811,In_471);
xor U1624 (N_1624,In_299,In_267);
and U1625 (N_1625,In_737,In_1121);
xor U1626 (N_1626,In_1380,In_1800);
and U1627 (N_1627,In_991,In_1987);
xor U1628 (N_1628,In_1386,In_116);
xor U1629 (N_1629,In_311,In_9);
nand U1630 (N_1630,In_1287,In_1329);
and U1631 (N_1631,In_639,In_1403);
nand U1632 (N_1632,In_817,In_1086);
or U1633 (N_1633,In_472,In_825);
or U1634 (N_1634,In_1054,In_1550);
xnor U1635 (N_1635,In_1157,In_551);
xnor U1636 (N_1636,In_464,In_1918);
xor U1637 (N_1637,In_786,In_1547);
or U1638 (N_1638,In_1138,In_1094);
or U1639 (N_1639,In_1711,In_1378);
nor U1640 (N_1640,In_1164,In_1256);
nand U1641 (N_1641,In_593,In_1390);
nand U1642 (N_1642,In_1825,In_81);
xnor U1643 (N_1643,In_1843,In_71);
xor U1644 (N_1644,In_1820,In_1167);
nand U1645 (N_1645,In_1518,In_674);
and U1646 (N_1646,In_1207,In_41);
and U1647 (N_1647,In_7,In_1127);
or U1648 (N_1648,In_174,In_1970);
nand U1649 (N_1649,In_81,In_1265);
and U1650 (N_1650,In_426,In_1368);
nand U1651 (N_1651,In_466,In_916);
and U1652 (N_1652,In_707,In_1566);
nand U1653 (N_1653,In_1018,In_587);
nand U1654 (N_1654,In_997,In_1192);
and U1655 (N_1655,In_1955,In_924);
xor U1656 (N_1656,In_659,In_996);
and U1657 (N_1657,In_487,In_1950);
and U1658 (N_1658,In_1508,In_944);
nor U1659 (N_1659,In_1194,In_944);
nand U1660 (N_1660,In_593,In_1478);
or U1661 (N_1661,In_1654,In_622);
and U1662 (N_1662,In_331,In_1289);
xnor U1663 (N_1663,In_811,In_957);
or U1664 (N_1664,In_1863,In_164);
and U1665 (N_1665,In_959,In_626);
and U1666 (N_1666,In_1334,In_550);
nand U1667 (N_1667,In_452,In_1625);
xor U1668 (N_1668,In_56,In_405);
nor U1669 (N_1669,In_291,In_257);
and U1670 (N_1670,In_540,In_1516);
nor U1671 (N_1671,In_1119,In_1842);
xor U1672 (N_1672,In_1128,In_1747);
and U1673 (N_1673,In_1192,In_1650);
xnor U1674 (N_1674,In_110,In_841);
or U1675 (N_1675,In_649,In_1609);
or U1676 (N_1676,In_364,In_1214);
nor U1677 (N_1677,In_1376,In_1644);
or U1678 (N_1678,In_416,In_411);
and U1679 (N_1679,In_459,In_1160);
nand U1680 (N_1680,In_468,In_1334);
nor U1681 (N_1681,In_645,In_1378);
nand U1682 (N_1682,In_1985,In_983);
xor U1683 (N_1683,In_233,In_551);
nand U1684 (N_1684,In_1288,In_415);
or U1685 (N_1685,In_1685,In_1247);
or U1686 (N_1686,In_1945,In_1557);
xnor U1687 (N_1687,In_1867,In_1731);
nor U1688 (N_1688,In_897,In_801);
nor U1689 (N_1689,In_1762,In_1062);
nor U1690 (N_1690,In_1950,In_1236);
and U1691 (N_1691,In_1054,In_554);
or U1692 (N_1692,In_45,In_1672);
and U1693 (N_1693,In_980,In_1651);
xor U1694 (N_1694,In_84,In_1858);
nand U1695 (N_1695,In_831,In_800);
or U1696 (N_1696,In_1082,In_773);
xnor U1697 (N_1697,In_1191,In_310);
nor U1698 (N_1698,In_803,In_922);
xor U1699 (N_1699,In_787,In_310);
xnor U1700 (N_1700,In_778,In_865);
xnor U1701 (N_1701,In_766,In_898);
nor U1702 (N_1702,In_404,In_686);
nand U1703 (N_1703,In_1980,In_31);
nor U1704 (N_1704,In_1019,In_1408);
and U1705 (N_1705,In_1320,In_1300);
nand U1706 (N_1706,In_229,In_824);
or U1707 (N_1707,In_615,In_133);
or U1708 (N_1708,In_1338,In_1599);
xor U1709 (N_1709,In_1665,In_433);
nand U1710 (N_1710,In_219,In_1950);
xor U1711 (N_1711,In_1644,In_291);
nor U1712 (N_1712,In_90,In_374);
nand U1713 (N_1713,In_133,In_793);
or U1714 (N_1714,In_1562,In_1601);
xnor U1715 (N_1715,In_1327,In_906);
nand U1716 (N_1716,In_764,In_1309);
or U1717 (N_1717,In_1637,In_761);
nand U1718 (N_1718,In_502,In_814);
nand U1719 (N_1719,In_974,In_1129);
and U1720 (N_1720,In_607,In_877);
xnor U1721 (N_1721,In_1394,In_1260);
xnor U1722 (N_1722,In_704,In_302);
nor U1723 (N_1723,In_234,In_1935);
xor U1724 (N_1724,In_877,In_1368);
nor U1725 (N_1725,In_897,In_286);
xnor U1726 (N_1726,In_581,In_369);
nand U1727 (N_1727,In_225,In_1624);
and U1728 (N_1728,In_1427,In_1011);
and U1729 (N_1729,In_201,In_1269);
or U1730 (N_1730,In_1929,In_1765);
nor U1731 (N_1731,In_208,In_496);
and U1732 (N_1732,In_405,In_652);
nor U1733 (N_1733,In_471,In_374);
xnor U1734 (N_1734,In_1874,In_1679);
and U1735 (N_1735,In_1779,In_892);
and U1736 (N_1736,In_1108,In_690);
xnor U1737 (N_1737,In_92,In_983);
nor U1738 (N_1738,In_1178,In_1673);
nor U1739 (N_1739,In_433,In_154);
or U1740 (N_1740,In_1073,In_198);
nand U1741 (N_1741,In_737,In_1066);
xnor U1742 (N_1742,In_661,In_870);
and U1743 (N_1743,In_854,In_982);
and U1744 (N_1744,In_1329,In_440);
nor U1745 (N_1745,In_1660,In_18);
nand U1746 (N_1746,In_1751,In_1351);
nand U1747 (N_1747,In_1206,In_217);
or U1748 (N_1748,In_1790,In_1043);
xor U1749 (N_1749,In_190,In_176);
nand U1750 (N_1750,In_1486,In_1618);
xor U1751 (N_1751,In_737,In_1131);
and U1752 (N_1752,In_346,In_633);
nand U1753 (N_1753,In_93,In_748);
or U1754 (N_1754,In_1404,In_471);
nand U1755 (N_1755,In_1291,In_1241);
and U1756 (N_1756,In_541,In_849);
xnor U1757 (N_1757,In_691,In_549);
or U1758 (N_1758,In_586,In_838);
nor U1759 (N_1759,In_1930,In_705);
xor U1760 (N_1760,In_838,In_220);
nor U1761 (N_1761,In_1770,In_1914);
nand U1762 (N_1762,In_1555,In_674);
xnor U1763 (N_1763,In_1984,In_1379);
nand U1764 (N_1764,In_672,In_1819);
nor U1765 (N_1765,In_1910,In_587);
xnor U1766 (N_1766,In_1787,In_640);
or U1767 (N_1767,In_1018,In_726);
nand U1768 (N_1768,In_30,In_1367);
nand U1769 (N_1769,In_305,In_1362);
nand U1770 (N_1770,In_1470,In_1556);
or U1771 (N_1771,In_1690,In_606);
and U1772 (N_1772,In_911,In_839);
xnor U1773 (N_1773,In_267,In_1996);
or U1774 (N_1774,In_1763,In_1388);
nor U1775 (N_1775,In_362,In_1126);
or U1776 (N_1776,In_1592,In_1837);
xnor U1777 (N_1777,In_475,In_1946);
nor U1778 (N_1778,In_464,In_846);
nor U1779 (N_1779,In_671,In_1680);
and U1780 (N_1780,In_86,In_1267);
xnor U1781 (N_1781,In_463,In_1311);
or U1782 (N_1782,In_1255,In_554);
nor U1783 (N_1783,In_117,In_1794);
and U1784 (N_1784,In_1289,In_291);
xnor U1785 (N_1785,In_1292,In_405);
nand U1786 (N_1786,In_1824,In_988);
or U1787 (N_1787,In_978,In_1896);
and U1788 (N_1788,In_282,In_514);
and U1789 (N_1789,In_606,In_1284);
and U1790 (N_1790,In_1955,In_573);
and U1791 (N_1791,In_682,In_19);
or U1792 (N_1792,In_679,In_1914);
xor U1793 (N_1793,In_979,In_1664);
and U1794 (N_1794,In_38,In_152);
nand U1795 (N_1795,In_885,In_1319);
or U1796 (N_1796,In_1711,In_1292);
xnor U1797 (N_1797,In_760,In_1294);
xnor U1798 (N_1798,In_1158,In_867);
xor U1799 (N_1799,In_647,In_1659);
nand U1800 (N_1800,In_1838,In_1060);
xor U1801 (N_1801,In_1579,In_179);
or U1802 (N_1802,In_373,In_1464);
or U1803 (N_1803,In_1377,In_634);
or U1804 (N_1804,In_1618,In_1811);
and U1805 (N_1805,In_1789,In_101);
nand U1806 (N_1806,In_1068,In_627);
or U1807 (N_1807,In_478,In_522);
and U1808 (N_1808,In_1291,In_1038);
xor U1809 (N_1809,In_880,In_688);
or U1810 (N_1810,In_68,In_503);
or U1811 (N_1811,In_1291,In_4);
xor U1812 (N_1812,In_366,In_305);
xor U1813 (N_1813,In_1563,In_1336);
and U1814 (N_1814,In_1169,In_530);
nor U1815 (N_1815,In_1309,In_1560);
xnor U1816 (N_1816,In_524,In_906);
nand U1817 (N_1817,In_1859,In_744);
or U1818 (N_1818,In_431,In_671);
and U1819 (N_1819,In_958,In_835);
and U1820 (N_1820,In_1909,In_1186);
and U1821 (N_1821,In_257,In_45);
or U1822 (N_1822,In_254,In_498);
nor U1823 (N_1823,In_209,In_1042);
nor U1824 (N_1824,In_1878,In_748);
xnor U1825 (N_1825,In_192,In_114);
nor U1826 (N_1826,In_470,In_436);
nand U1827 (N_1827,In_1439,In_571);
xnor U1828 (N_1828,In_681,In_1499);
nand U1829 (N_1829,In_154,In_897);
and U1830 (N_1830,In_749,In_479);
and U1831 (N_1831,In_1075,In_670);
or U1832 (N_1832,In_808,In_1332);
xor U1833 (N_1833,In_1936,In_1392);
nor U1834 (N_1834,In_1651,In_563);
nor U1835 (N_1835,In_198,In_1549);
and U1836 (N_1836,In_1524,In_1885);
nand U1837 (N_1837,In_1190,In_1845);
xor U1838 (N_1838,In_1188,In_435);
xor U1839 (N_1839,In_105,In_1558);
or U1840 (N_1840,In_989,In_968);
nand U1841 (N_1841,In_1524,In_1346);
nand U1842 (N_1842,In_1780,In_1164);
nor U1843 (N_1843,In_208,In_1364);
and U1844 (N_1844,In_455,In_204);
nor U1845 (N_1845,In_438,In_157);
nand U1846 (N_1846,In_1146,In_590);
or U1847 (N_1847,In_28,In_16);
or U1848 (N_1848,In_1105,In_1915);
nand U1849 (N_1849,In_1642,In_1115);
xnor U1850 (N_1850,In_493,In_1762);
and U1851 (N_1851,In_590,In_1290);
nand U1852 (N_1852,In_326,In_1584);
xnor U1853 (N_1853,In_718,In_40);
nor U1854 (N_1854,In_1871,In_1353);
xor U1855 (N_1855,In_1102,In_452);
and U1856 (N_1856,In_478,In_1854);
nor U1857 (N_1857,In_1279,In_717);
nor U1858 (N_1858,In_90,In_36);
nor U1859 (N_1859,In_1831,In_291);
xnor U1860 (N_1860,In_1692,In_1897);
or U1861 (N_1861,In_1956,In_1023);
nor U1862 (N_1862,In_1557,In_613);
xnor U1863 (N_1863,In_988,In_413);
nand U1864 (N_1864,In_1587,In_1185);
xor U1865 (N_1865,In_637,In_1415);
nor U1866 (N_1866,In_720,In_669);
or U1867 (N_1867,In_1019,In_673);
nand U1868 (N_1868,In_194,In_962);
xnor U1869 (N_1869,In_347,In_718);
and U1870 (N_1870,In_1904,In_90);
nand U1871 (N_1871,In_1599,In_799);
nor U1872 (N_1872,In_264,In_425);
nor U1873 (N_1873,In_1949,In_1930);
xnor U1874 (N_1874,In_1220,In_1300);
nand U1875 (N_1875,In_247,In_1467);
and U1876 (N_1876,In_1111,In_922);
xnor U1877 (N_1877,In_1953,In_1023);
or U1878 (N_1878,In_140,In_1134);
nor U1879 (N_1879,In_1751,In_832);
nor U1880 (N_1880,In_1039,In_470);
nor U1881 (N_1881,In_864,In_1246);
and U1882 (N_1882,In_1014,In_1321);
nand U1883 (N_1883,In_1741,In_654);
nand U1884 (N_1884,In_1680,In_1867);
or U1885 (N_1885,In_106,In_1944);
xnor U1886 (N_1886,In_1490,In_1483);
or U1887 (N_1887,In_211,In_1835);
nor U1888 (N_1888,In_213,In_231);
xor U1889 (N_1889,In_460,In_1675);
and U1890 (N_1890,In_1411,In_192);
xnor U1891 (N_1891,In_1973,In_929);
nor U1892 (N_1892,In_841,In_700);
nand U1893 (N_1893,In_464,In_750);
nor U1894 (N_1894,In_1605,In_381);
and U1895 (N_1895,In_992,In_313);
nand U1896 (N_1896,In_191,In_81);
nand U1897 (N_1897,In_1865,In_1094);
and U1898 (N_1898,In_1528,In_1578);
or U1899 (N_1899,In_954,In_813);
and U1900 (N_1900,In_812,In_738);
and U1901 (N_1901,In_1500,In_1699);
xnor U1902 (N_1902,In_163,In_1282);
nor U1903 (N_1903,In_706,In_1239);
and U1904 (N_1904,In_167,In_1629);
and U1905 (N_1905,In_151,In_1564);
and U1906 (N_1906,In_1791,In_322);
xnor U1907 (N_1907,In_1644,In_752);
or U1908 (N_1908,In_1225,In_503);
and U1909 (N_1909,In_1005,In_1923);
or U1910 (N_1910,In_1968,In_1572);
nor U1911 (N_1911,In_1726,In_778);
or U1912 (N_1912,In_207,In_1819);
xnor U1913 (N_1913,In_68,In_1756);
xor U1914 (N_1914,In_747,In_118);
xor U1915 (N_1915,In_1117,In_624);
nand U1916 (N_1916,In_1096,In_585);
and U1917 (N_1917,In_1587,In_923);
or U1918 (N_1918,In_75,In_1075);
and U1919 (N_1919,In_70,In_1416);
xnor U1920 (N_1920,In_424,In_1629);
and U1921 (N_1921,In_1439,In_1331);
xnor U1922 (N_1922,In_1912,In_32);
or U1923 (N_1923,In_158,In_881);
or U1924 (N_1924,In_178,In_121);
and U1925 (N_1925,In_332,In_1904);
and U1926 (N_1926,In_722,In_1402);
nand U1927 (N_1927,In_1246,In_1379);
and U1928 (N_1928,In_1579,In_799);
or U1929 (N_1929,In_1668,In_1376);
xnor U1930 (N_1930,In_1186,In_1968);
and U1931 (N_1931,In_1566,In_1877);
or U1932 (N_1932,In_833,In_1260);
or U1933 (N_1933,In_1351,In_1549);
xnor U1934 (N_1934,In_719,In_580);
xnor U1935 (N_1935,In_416,In_1945);
or U1936 (N_1936,In_1063,In_1509);
or U1937 (N_1937,In_520,In_253);
nand U1938 (N_1938,In_811,In_12);
and U1939 (N_1939,In_1558,In_1139);
nand U1940 (N_1940,In_1597,In_567);
or U1941 (N_1941,In_614,In_165);
and U1942 (N_1942,In_1556,In_345);
or U1943 (N_1943,In_1583,In_1064);
nor U1944 (N_1944,In_976,In_1032);
nand U1945 (N_1945,In_247,In_837);
and U1946 (N_1946,In_949,In_549);
and U1947 (N_1947,In_162,In_1966);
nor U1948 (N_1948,In_1479,In_1540);
nor U1949 (N_1949,In_458,In_1924);
xnor U1950 (N_1950,In_1023,In_1846);
or U1951 (N_1951,In_1948,In_790);
nand U1952 (N_1952,In_498,In_1385);
or U1953 (N_1953,In_1770,In_1251);
nand U1954 (N_1954,In_892,In_798);
nor U1955 (N_1955,In_1117,In_1700);
nand U1956 (N_1956,In_1902,In_1253);
xnor U1957 (N_1957,In_846,In_71);
and U1958 (N_1958,In_418,In_111);
nand U1959 (N_1959,In_876,In_1029);
or U1960 (N_1960,In_1667,In_1024);
or U1961 (N_1961,In_1014,In_101);
xnor U1962 (N_1962,In_1242,In_1657);
or U1963 (N_1963,In_1409,In_1567);
or U1964 (N_1964,In_712,In_630);
xnor U1965 (N_1965,In_1371,In_1437);
nand U1966 (N_1966,In_1856,In_115);
and U1967 (N_1967,In_456,In_1749);
or U1968 (N_1968,In_105,In_365);
and U1969 (N_1969,In_674,In_517);
and U1970 (N_1970,In_465,In_460);
nand U1971 (N_1971,In_479,In_990);
nand U1972 (N_1972,In_757,In_823);
nor U1973 (N_1973,In_1949,In_1495);
nor U1974 (N_1974,In_1495,In_1360);
or U1975 (N_1975,In_1008,In_1418);
or U1976 (N_1976,In_1910,In_1757);
or U1977 (N_1977,In_1017,In_1629);
xnor U1978 (N_1978,In_9,In_1953);
nor U1979 (N_1979,In_1730,In_1437);
nor U1980 (N_1980,In_1119,In_737);
nor U1981 (N_1981,In_1577,In_105);
and U1982 (N_1982,In_856,In_1182);
and U1983 (N_1983,In_479,In_367);
nor U1984 (N_1984,In_479,In_508);
nor U1985 (N_1985,In_48,In_1932);
and U1986 (N_1986,In_1165,In_1267);
or U1987 (N_1987,In_1342,In_1857);
nand U1988 (N_1988,In_1366,In_816);
and U1989 (N_1989,In_1967,In_1045);
or U1990 (N_1990,In_1915,In_783);
nand U1991 (N_1991,In_130,In_481);
xor U1992 (N_1992,In_788,In_856);
nand U1993 (N_1993,In_719,In_287);
or U1994 (N_1994,In_392,In_1781);
or U1995 (N_1995,In_964,In_1624);
nor U1996 (N_1996,In_939,In_21);
nor U1997 (N_1997,In_1851,In_219);
nor U1998 (N_1998,In_1440,In_761);
nand U1999 (N_1999,In_694,In_1912);
nand U2000 (N_2000,In_1410,In_1424);
xnor U2001 (N_2001,In_352,In_894);
xnor U2002 (N_2002,In_1715,In_1080);
or U2003 (N_2003,In_1530,In_1680);
and U2004 (N_2004,In_33,In_238);
nand U2005 (N_2005,In_321,In_740);
nor U2006 (N_2006,In_862,In_1257);
and U2007 (N_2007,In_573,In_1872);
and U2008 (N_2008,In_1680,In_1053);
and U2009 (N_2009,In_1920,In_985);
nand U2010 (N_2010,In_900,In_1727);
xor U2011 (N_2011,In_638,In_517);
nand U2012 (N_2012,In_152,In_1114);
nand U2013 (N_2013,In_1079,In_1264);
nor U2014 (N_2014,In_1441,In_1985);
nor U2015 (N_2015,In_553,In_260);
and U2016 (N_2016,In_867,In_948);
xor U2017 (N_2017,In_45,In_395);
or U2018 (N_2018,In_1847,In_1063);
and U2019 (N_2019,In_1297,In_1334);
xor U2020 (N_2020,In_1932,In_1008);
xor U2021 (N_2021,In_1875,In_9);
nor U2022 (N_2022,In_638,In_1993);
xnor U2023 (N_2023,In_1821,In_1410);
nand U2024 (N_2024,In_1933,In_1360);
nand U2025 (N_2025,In_1370,In_1713);
nand U2026 (N_2026,In_508,In_333);
nor U2027 (N_2027,In_830,In_127);
or U2028 (N_2028,In_388,In_68);
or U2029 (N_2029,In_1769,In_411);
or U2030 (N_2030,In_1257,In_1012);
xnor U2031 (N_2031,In_493,In_1239);
xor U2032 (N_2032,In_976,In_832);
nand U2033 (N_2033,In_935,In_1944);
and U2034 (N_2034,In_752,In_821);
xor U2035 (N_2035,In_394,In_206);
xor U2036 (N_2036,In_205,In_645);
xor U2037 (N_2037,In_1121,In_227);
or U2038 (N_2038,In_1135,In_1243);
xnor U2039 (N_2039,In_353,In_315);
nor U2040 (N_2040,In_1023,In_563);
xor U2041 (N_2041,In_225,In_536);
xor U2042 (N_2042,In_371,In_417);
or U2043 (N_2043,In_982,In_796);
and U2044 (N_2044,In_454,In_1424);
nor U2045 (N_2045,In_1179,In_384);
and U2046 (N_2046,In_128,In_1268);
xnor U2047 (N_2047,In_437,In_1562);
nand U2048 (N_2048,In_1216,In_888);
nor U2049 (N_2049,In_1869,In_1667);
xnor U2050 (N_2050,In_60,In_1218);
nand U2051 (N_2051,In_1571,In_780);
xor U2052 (N_2052,In_422,In_1657);
nand U2053 (N_2053,In_83,In_1453);
or U2054 (N_2054,In_1132,In_1761);
nor U2055 (N_2055,In_1534,In_269);
and U2056 (N_2056,In_1230,In_287);
xor U2057 (N_2057,In_770,In_398);
xor U2058 (N_2058,In_193,In_1448);
nor U2059 (N_2059,In_736,In_1143);
xnor U2060 (N_2060,In_1210,In_996);
nor U2061 (N_2061,In_70,In_41);
or U2062 (N_2062,In_1395,In_1747);
nor U2063 (N_2063,In_917,In_325);
or U2064 (N_2064,In_1886,In_1593);
or U2065 (N_2065,In_1789,In_430);
or U2066 (N_2066,In_196,In_1649);
or U2067 (N_2067,In_1749,In_323);
nor U2068 (N_2068,In_1696,In_858);
and U2069 (N_2069,In_53,In_353);
xnor U2070 (N_2070,In_918,In_45);
xnor U2071 (N_2071,In_906,In_572);
nand U2072 (N_2072,In_737,In_1429);
xnor U2073 (N_2073,In_1344,In_635);
nand U2074 (N_2074,In_299,In_822);
and U2075 (N_2075,In_1372,In_923);
nor U2076 (N_2076,In_1602,In_795);
nor U2077 (N_2077,In_1833,In_1062);
or U2078 (N_2078,In_572,In_446);
or U2079 (N_2079,In_1865,In_1857);
nor U2080 (N_2080,In_1186,In_961);
or U2081 (N_2081,In_837,In_495);
xnor U2082 (N_2082,In_190,In_1483);
or U2083 (N_2083,In_1184,In_348);
nand U2084 (N_2084,In_890,In_1799);
xor U2085 (N_2085,In_1939,In_1948);
xnor U2086 (N_2086,In_962,In_1128);
nor U2087 (N_2087,In_111,In_1599);
xor U2088 (N_2088,In_470,In_524);
xnor U2089 (N_2089,In_1173,In_549);
nor U2090 (N_2090,In_1688,In_395);
xnor U2091 (N_2091,In_717,In_1429);
nand U2092 (N_2092,In_884,In_254);
xnor U2093 (N_2093,In_1865,In_1350);
or U2094 (N_2094,In_243,In_1154);
or U2095 (N_2095,In_666,In_235);
or U2096 (N_2096,In_171,In_1815);
or U2097 (N_2097,In_1113,In_1271);
xnor U2098 (N_2098,In_1867,In_1142);
nor U2099 (N_2099,In_1419,In_1855);
nor U2100 (N_2100,In_1677,In_1660);
and U2101 (N_2101,In_45,In_327);
and U2102 (N_2102,In_1411,In_637);
and U2103 (N_2103,In_1533,In_425);
xor U2104 (N_2104,In_686,In_322);
or U2105 (N_2105,In_632,In_82);
xor U2106 (N_2106,In_239,In_1365);
xor U2107 (N_2107,In_709,In_1431);
nor U2108 (N_2108,In_1443,In_1859);
and U2109 (N_2109,In_72,In_711);
xor U2110 (N_2110,In_324,In_1185);
and U2111 (N_2111,In_1426,In_832);
or U2112 (N_2112,In_467,In_81);
or U2113 (N_2113,In_1735,In_727);
nor U2114 (N_2114,In_1936,In_414);
nand U2115 (N_2115,In_1628,In_219);
xnor U2116 (N_2116,In_1941,In_942);
xnor U2117 (N_2117,In_1853,In_692);
or U2118 (N_2118,In_1718,In_370);
xnor U2119 (N_2119,In_700,In_296);
nand U2120 (N_2120,In_733,In_1951);
nand U2121 (N_2121,In_1537,In_1630);
and U2122 (N_2122,In_1283,In_1718);
nand U2123 (N_2123,In_985,In_592);
and U2124 (N_2124,In_1917,In_988);
nand U2125 (N_2125,In_1954,In_370);
or U2126 (N_2126,In_1663,In_1747);
xnor U2127 (N_2127,In_1098,In_1907);
xnor U2128 (N_2128,In_389,In_737);
xnor U2129 (N_2129,In_1899,In_273);
nor U2130 (N_2130,In_57,In_1950);
nand U2131 (N_2131,In_809,In_366);
and U2132 (N_2132,In_431,In_1301);
xnor U2133 (N_2133,In_1250,In_1918);
nand U2134 (N_2134,In_571,In_884);
and U2135 (N_2135,In_1930,In_957);
nand U2136 (N_2136,In_928,In_1629);
nand U2137 (N_2137,In_1631,In_481);
nor U2138 (N_2138,In_1820,In_1361);
nand U2139 (N_2139,In_1703,In_1983);
xnor U2140 (N_2140,In_1718,In_502);
nor U2141 (N_2141,In_1809,In_1926);
and U2142 (N_2142,In_1135,In_1904);
nand U2143 (N_2143,In_130,In_1804);
or U2144 (N_2144,In_1736,In_788);
or U2145 (N_2145,In_111,In_630);
and U2146 (N_2146,In_1057,In_484);
nor U2147 (N_2147,In_922,In_21);
xor U2148 (N_2148,In_1699,In_1279);
or U2149 (N_2149,In_671,In_1107);
nor U2150 (N_2150,In_1998,In_910);
nand U2151 (N_2151,In_1115,In_688);
xor U2152 (N_2152,In_375,In_1636);
and U2153 (N_2153,In_893,In_290);
nand U2154 (N_2154,In_1250,In_1943);
xnor U2155 (N_2155,In_803,In_1889);
and U2156 (N_2156,In_1924,In_1938);
xor U2157 (N_2157,In_1471,In_577);
xnor U2158 (N_2158,In_1293,In_847);
nor U2159 (N_2159,In_233,In_1145);
nor U2160 (N_2160,In_1757,In_1238);
xor U2161 (N_2161,In_1020,In_973);
nand U2162 (N_2162,In_1448,In_1422);
xnor U2163 (N_2163,In_186,In_1901);
or U2164 (N_2164,In_499,In_169);
and U2165 (N_2165,In_1026,In_82);
and U2166 (N_2166,In_1595,In_22);
xnor U2167 (N_2167,In_1026,In_1342);
xor U2168 (N_2168,In_1488,In_1508);
nand U2169 (N_2169,In_1384,In_1455);
and U2170 (N_2170,In_327,In_1963);
xnor U2171 (N_2171,In_500,In_727);
or U2172 (N_2172,In_710,In_1523);
or U2173 (N_2173,In_616,In_1188);
or U2174 (N_2174,In_1609,In_1903);
and U2175 (N_2175,In_1571,In_1700);
and U2176 (N_2176,In_1537,In_894);
or U2177 (N_2177,In_335,In_989);
xnor U2178 (N_2178,In_409,In_394);
or U2179 (N_2179,In_1980,In_1783);
or U2180 (N_2180,In_15,In_642);
xnor U2181 (N_2181,In_1934,In_1371);
or U2182 (N_2182,In_179,In_551);
nor U2183 (N_2183,In_508,In_318);
nor U2184 (N_2184,In_1242,In_1141);
or U2185 (N_2185,In_1681,In_1510);
nor U2186 (N_2186,In_1251,In_1176);
and U2187 (N_2187,In_1983,In_54);
nand U2188 (N_2188,In_1851,In_389);
nand U2189 (N_2189,In_1079,In_1926);
xor U2190 (N_2190,In_1917,In_902);
or U2191 (N_2191,In_1031,In_44);
xor U2192 (N_2192,In_923,In_673);
nand U2193 (N_2193,In_955,In_990);
or U2194 (N_2194,In_518,In_767);
nand U2195 (N_2195,In_1089,In_314);
and U2196 (N_2196,In_1405,In_1154);
nor U2197 (N_2197,In_1170,In_1471);
nor U2198 (N_2198,In_956,In_1590);
and U2199 (N_2199,In_1476,In_1062);
or U2200 (N_2200,In_937,In_1754);
nor U2201 (N_2201,In_696,In_1848);
xnor U2202 (N_2202,In_677,In_1546);
or U2203 (N_2203,In_243,In_1920);
and U2204 (N_2204,In_1600,In_198);
and U2205 (N_2205,In_788,In_1738);
xor U2206 (N_2206,In_181,In_581);
and U2207 (N_2207,In_915,In_106);
or U2208 (N_2208,In_919,In_1217);
and U2209 (N_2209,In_845,In_1874);
nor U2210 (N_2210,In_117,In_698);
or U2211 (N_2211,In_741,In_1663);
and U2212 (N_2212,In_809,In_367);
and U2213 (N_2213,In_862,In_676);
nand U2214 (N_2214,In_461,In_1528);
or U2215 (N_2215,In_1746,In_1370);
or U2216 (N_2216,In_1474,In_927);
and U2217 (N_2217,In_948,In_698);
or U2218 (N_2218,In_692,In_1812);
or U2219 (N_2219,In_232,In_1182);
or U2220 (N_2220,In_1900,In_1155);
nand U2221 (N_2221,In_1432,In_129);
and U2222 (N_2222,In_1912,In_531);
and U2223 (N_2223,In_1314,In_894);
or U2224 (N_2224,In_437,In_987);
xor U2225 (N_2225,In_1808,In_884);
nand U2226 (N_2226,In_658,In_71);
nor U2227 (N_2227,In_755,In_123);
nand U2228 (N_2228,In_686,In_1627);
nor U2229 (N_2229,In_433,In_646);
nor U2230 (N_2230,In_593,In_1761);
xnor U2231 (N_2231,In_121,In_640);
and U2232 (N_2232,In_876,In_1165);
and U2233 (N_2233,In_1325,In_961);
and U2234 (N_2234,In_172,In_1541);
or U2235 (N_2235,In_363,In_1129);
and U2236 (N_2236,In_422,In_1228);
xnor U2237 (N_2237,In_1390,In_70);
xor U2238 (N_2238,In_44,In_1435);
and U2239 (N_2239,In_794,In_1157);
xor U2240 (N_2240,In_1719,In_1914);
nor U2241 (N_2241,In_1587,In_1010);
or U2242 (N_2242,In_1646,In_451);
or U2243 (N_2243,In_58,In_602);
nand U2244 (N_2244,In_982,In_117);
nor U2245 (N_2245,In_309,In_1273);
nand U2246 (N_2246,In_1874,In_825);
nor U2247 (N_2247,In_1428,In_243);
or U2248 (N_2248,In_121,In_1999);
nand U2249 (N_2249,In_843,In_680);
and U2250 (N_2250,In_1868,In_1370);
and U2251 (N_2251,In_133,In_122);
and U2252 (N_2252,In_1762,In_840);
xor U2253 (N_2253,In_274,In_1530);
nand U2254 (N_2254,In_1711,In_1636);
nor U2255 (N_2255,In_930,In_358);
xor U2256 (N_2256,In_806,In_146);
or U2257 (N_2257,In_88,In_488);
and U2258 (N_2258,In_1295,In_1930);
and U2259 (N_2259,In_1116,In_870);
xor U2260 (N_2260,In_87,In_1869);
nor U2261 (N_2261,In_1563,In_14);
or U2262 (N_2262,In_578,In_1090);
nand U2263 (N_2263,In_1647,In_971);
or U2264 (N_2264,In_285,In_1952);
xnor U2265 (N_2265,In_1188,In_345);
nor U2266 (N_2266,In_1606,In_648);
and U2267 (N_2267,In_1115,In_1747);
xor U2268 (N_2268,In_48,In_1552);
and U2269 (N_2269,In_1233,In_256);
nand U2270 (N_2270,In_8,In_66);
or U2271 (N_2271,In_608,In_1612);
nor U2272 (N_2272,In_700,In_729);
and U2273 (N_2273,In_868,In_1699);
xor U2274 (N_2274,In_1059,In_759);
xnor U2275 (N_2275,In_1693,In_798);
xnor U2276 (N_2276,In_435,In_1331);
xnor U2277 (N_2277,In_71,In_1199);
nor U2278 (N_2278,In_1975,In_256);
and U2279 (N_2279,In_851,In_890);
xor U2280 (N_2280,In_158,In_218);
or U2281 (N_2281,In_226,In_1339);
or U2282 (N_2282,In_1885,In_807);
nand U2283 (N_2283,In_1170,In_512);
and U2284 (N_2284,In_695,In_1231);
xor U2285 (N_2285,In_785,In_810);
nand U2286 (N_2286,In_404,In_763);
nand U2287 (N_2287,In_355,In_1715);
nand U2288 (N_2288,In_1691,In_1417);
or U2289 (N_2289,In_407,In_596);
xor U2290 (N_2290,In_698,In_1582);
nand U2291 (N_2291,In_1407,In_326);
and U2292 (N_2292,In_1758,In_715);
xor U2293 (N_2293,In_419,In_260);
nand U2294 (N_2294,In_1042,In_524);
and U2295 (N_2295,In_1320,In_1030);
nand U2296 (N_2296,In_269,In_429);
and U2297 (N_2297,In_443,In_1697);
xor U2298 (N_2298,In_1785,In_1572);
and U2299 (N_2299,In_1560,In_1416);
nor U2300 (N_2300,In_76,In_470);
xnor U2301 (N_2301,In_1809,In_1658);
nor U2302 (N_2302,In_142,In_1176);
and U2303 (N_2303,In_522,In_1693);
nand U2304 (N_2304,In_1656,In_152);
nor U2305 (N_2305,In_1154,In_44);
nand U2306 (N_2306,In_1009,In_192);
xnor U2307 (N_2307,In_321,In_276);
or U2308 (N_2308,In_240,In_645);
or U2309 (N_2309,In_604,In_1877);
or U2310 (N_2310,In_1195,In_1008);
nor U2311 (N_2311,In_785,In_668);
nand U2312 (N_2312,In_1417,In_1245);
or U2313 (N_2313,In_1984,In_326);
xor U2314 (N_2314,In_1540,In_1573);
nor U2315 (N_2315,In_496,In_1615);
xor U2316 (N_2316,In_1882,In_80);
nor U2317 (N_2317,In_1821,In_565);
xor U2318 (N_2318,In_1447,In_1122);
xnor U2319 (N_2319,In_681,In_561);
xor U2320 (N_2320,In_1598,In_1138);
or U2321 (N_2321,In_949,In_911);
nor U2322 (N_2322,In_395,In_698);
nor U2323 (N_2323,In_1947,In_296);
nand U2324 (N_2324,In_1388,In_1097);
and U2325 (N_2325,In_1572,In_1009);
nand U2326 (N_2326,In_900,In_1492);
nor U2327 (N_2327,In_502,In_1527);
nor U2328 (N_2328,In_814,In_1922);
nand U2329 (N_2329,In_1074,In_1248);
xor U2330 (N_2330,In_240,In_1493);
nor U2331 (N_2331,In_1479,In_1343);
and U2332 (N_2332,In_1363,In_1997);
and U2333 (N_2333,In_1378,In_1202);
or U2334 (N_2334,In_1789,In_1314);
nand U2335 (N_2335,In_1100,In_1642);
xnor U2336 (N_2336,In_264,In_1535);
nand U2337 (N_2337,In_1970,In_1255);
xor U2338 (N_2338,In_1703,In_1919);
nand U2339 (N_2339,In_592,In_1515);
nor U2340 (N_2340,In_292,In_1348);
nand U2341 (N_2341,In_73,In_121);
nor U2342 (N_2342,In_1110,In_617);
nor U2343 (N_2343,In_409,In_1835);
and U2344 (N_2344,In_1433,In_624);
nand U2345 (N_2345,In_709,In_306);
xor U2346 (N_2346,In_1172,In_1342);
or U2347 (N_2347,In_572,In_1623);
nand U2348 (N_2348,In_566,In_1485);
nand U2349 (N_2349,In_937,In_1260);
and U2350 (N_2350,In_1412,In_1878);
and U2351 (N_2351,In_1434,In_1273);
nand U2352 (N_2352,In_1627,In_933);
and U2353 (N_2353,In_1083,In_1278);
or U2354 (N_2354,In_951,In_1995);
and U2355 (N_2355,In_337,In_449);
xor U2356 (N_2356,In_1979,In_1388);
or U2357 (N_2357,In_781,In_984);
nand U2358 (N_2358,In_871,In_1670);
and U2359 (N_2359,In_533,In_540);
xnor U2360 (N_2360,In_1779,In_1533);
xnor U2361 (N_2361,In_637,In_962);
nand U2362 (N_2362,In_11,In_105);
or U2363 (N_2363,In_1741,In_984);
nor U2364 (N_2364,In_687,In_432);
nand U2365 (N_2365,In_1745,In_1009);
xor U2366 (N_2366,In_1264,In_79);
nand U2367 (N_2367,In_1407,In_737);
nor U2368 (N_2368,In_332,In_594);
nand U2369 (N_2369,In_331,In_1056);
nand U2370 (N_2370,In_1866,In_870);
and U2371 (N_2371,In_1910,In_66);
and U2372 (N_2372,In_58,In_1636);
xnor U2373 (N_2373,In_1158,In_443);
and U2374 (N_2374,In_1048,In_780);
nor U2375 (N_2375,In_972,In_1691);
or U2376 (N_2376,In_1718,In_1999);
or U2377 (N_2377,In_1628,In_383);
and U2378 (N_2378,In_1913,In_1635);
nand U2379 (N_2379,In_1997,In_1889);
nor U2380 (N_2380,In_1341,In_1909);
and U2381 (N_2381,In_961,In_1858);
nor U2382 (N_2382,In_1763,In_744);
or U2383 (N_2383,In_469,In_554);
xor U2384 (N_2384,In_514,In_1688);
nor U2385 (N_2385,In_1808,In_969);
or U2386 (N_2386,In_877,In_1111);
nand U2387 (N_2387,In_1596,In_1718);
nor U2388 (N_2388,In_1408,In_1327);
xor U2389 (N_2389,In_489,In_1110);
or U2390 (N_2390,In_1879,In_428);
nand U2391 (N_2391,In_970,In_883);
or U2392 (N_2392,In_1201,In_721);
or U2393 (N_2393,In_1541,In_584);
nand U2394 (N_2394,In_1114,In_633);
xnor U2395 (N_2395,In_1480,In_234);
xnor U2396 (N_2396,In_480,In_1733);
nor U2397 (N_2397,In_720,In_368);
or U2398 (N_2398,In_1070,In_899);
and U2399 (N_2399,In_195,In_1597);
or U2400 (N_2400,In_907,In_1855);
nor U2401 (N_2401,In_1606,In_468);
and U2402 (N_2402,In_588,In_584);
nor U2403 (N_2403,In_648,In_1150);
and U2404 (N_2404,In_1807,In_1627);
and U2405 (N_2405,In_1994,In_1996);
nand U2406 (N_2406,In_632,In_398);
or U2407 (N_2407,In_83,In_942);
and U2408 (N_2408,In_609,In_1553);
xnor U2409 (N_2409,In_1368,In_442);
nor U2410 (N_2410,In_96,In_643);
and U2411 (N_2411,In_780,In_885);
and U2412 (N_2412,In_1916,In_768);
xor U2413 (N_2413,In_1658,In_1101);
nand U2414 (N_2414,In_942,In_683);
nand U2415 (N_2415,In_732,In_142);
xor U2416 (N_2416,In_763,In_282);
and U2417 (N_2417,In_1392,In_1618);
or U2418 (N_2418,In_783,In_1987);
or U2419 (N_2419,In_685,In_479);
xnor U2420 (N_2420,In_71,In_653);
or U2421 (N_2421,In_1837,In_225);
nand U2422 (N_2422,In_695,In_385);
nor U2423 (N_2423,In_852,In_1310);
or U2424 (N_2424,In_1908,In_1824);
nor U2425 (N_2425,In_1876,In_1418);
nand U2426 (N_2426,In_791,In_558);
nor U2427 (N_2427,In_679,In_1896);
and U2428 (N_2428,In_1266,In_720);
xor U2429 (N_2429,In_1297,In_996);
xor U2430 (N_2430,In_1293,In_1760);
xor U2431 (N_2431,In_720,In_683);
or U2432 (N_2432,In_306,In_932);
nand U2433 (N_2433,In_854,In_896);
or U2434 (N_2434,In_88,In_1634);
and U2435 (N_2435,In_1313,In_1841);
nor U2436 (N_2436,In_1488,In_226);
or U2437 (N_2437,In_38,In_1199);
and U2438 (N_2438,In_735,In_349);
nor U2439 (N_2439,In_1526,In_91);
and U2440 (N_2440,In_97,In_779);
xnor U2441 (N_2441,In_1073,In_1193);
and U2442 (N_2442,In_1919,In_1246);
nor U2443 (N_2443,In_224,In_473);
nand U2444 (N_2444,In_1423,In_471);
and U2445 (N_2445,In_1647,In_1609);
and U2446 (N_2446,In_141,In_286);
xor U2447 (N_2447,In_1712,In_1011);
and U2448 (N_2448,In_209,In_887);
or U2449 (N_2449,In_276,In_109);
nor U2450 (N_2450,In_712,In_1064);
xnor U2451 (N_2451,In_1798,In_1957);
xnor U2452 (N_2452,In_480,In_1468);
or U2453 (N_2453,In_1048,In_380);
and U2454 (N_2454,In_1493,In_557);
and U2455 (N_2455,In_443,In_1262);
nor U2456 (N_2456,In_656,In_1390);
or U2457 (N_2457,In_1696,In_2);
nand U2458 (N_2458,In_1811,In_611);
nor U2459 (N_2459,In_1707,In_1182);
and U2460 (N_2460,In_1379,In_705);
nor U2461 (N_2461,In_912,In_1221);
nand U2462 (N_2462,In_812,In_181);
and U2463 (N_2463,In_428,In_741);
nand U2464 (N_2464,In_823,In_1442);
xor U2465 (N_2465,In_1558,In_955);
xnor U2466 (N_2466,In_1266,In_1452);
and U2467 (N_2467,In_614,In_27);
xnor U2468 (N_2468,In_76,In_500);
and U2469 (N_2469,In_1722,In_1860);
or U2470 (N_2470,In_1394,In_551);
nand U2471 (N_2471,In_640,In_1646);
nand U2472 (N_2472,In_1197,In_509);
or U2473 (N_2473,In_247,In_302);
nand U2474 (N_2474,In_314,In_1665);
xor U2475 (N_2475,In_472,In_1432);
or U2476 (N_2476,In_26,In_1094);
nor U2477 (N_2477,In_833,In_231);
xnor U2478 (N_2478,In_1813,In_1809);
nor U2479 (N_2479,In_1936,In_309);
nor U2480 (N_2480,In_999,In_1634);
nand U2481 (N_2481,In_714,In_1581);
or U2482 (N_2482,In_1291,In_696);
and U2483 (N_2483,In_538,In_736);
xor U2484 (N_2484,In_753,In_1085);
xor U2485 (N_2485,In_1652,In_1456);
or U2486 (N_2486,In_619,In_1288);
xor U2487 (N_2487,In_1785,In_220);
and U2488 (N_2488,In_1849,In_279);
xnor U2489 (N_2489,In_272,In_766);
xnor U2490 (N_2490,In_1530,In_542);
xor U2491 (N_2491,In_497,In_1534);
xnor U2492 (N_2492,In_1378,In_1638);
nor U2493 (N_2493,In_1366,In_823);
and U2494 (N_2494,In_1860,In_95);
and U2495 (N_2495,In_353,In_1421);
nand U2496 (N_2496,In_1965,In_918);
nand U2497 (N_2497,In_1418,In_1377);
nand U2498 (N_2498,In_866,In_1811);
nand U2499 (N_2499,In_1793,In_1633);
nor U2500 (N_2500,In_817,In_884);
xnor U2501 (N_2501,In_146,In_1548);
or U2502 (N_2502,In_674,In_1689);
and U2503 (N_2503,In_131,In_1684);
nand U2504 (N_2504,In_1120,In_920);
nand U2505 (N_2505,In_1560,In_1127);
nor U2506 (N_2506,In_1789,In_1982);
nand U2507 (N_2507,In_312,In_1662);
nor U2508 (N_2508,In_931,In_1979);
or U2509 (N_2509,In_1110,In_21);
or U2510 (N_2510,In_441,In_24);
nor U2511 (N_2511,In_104,In_1357);
nand U2512 (N_2512,In_1461,In_206);
nor U2513 (N_2513,In_724,In_212);
nand U2514 (N_2514,In_710,In_543);
xnor U2515 (N_2515,In_254,In_1247);
or U2516 (N_2516,In_1432,In_335);
or U2517 (N_2517,In_1127,In_972);
nor U2518 (N_2518,In_1846,In_1323);
or U2519 (N_2519,In_292,In_1600);
nor U2520 (N_2520,In_1978,In_173);
nand U2521 (N_2521,In_289,In_343);
xor U2522 (N_2522,In_1596,In_1743);
or U2523 (N_2523,In_1711,In_1943);
and U2524 (N_2524,In_1008,In_83);
nand U2525 (N_2525,In_1700,In_336);
nor U2526 (N_2526,In_600,In_1795);
and U2527 (N_2527,In_1853,In_837);
nor U2528 (N_2528,In_1894,In_577);
or U2529 (N_2529,In_808,In_803);
nor U2530 (N_2530,In_1250,In_97);
nor U2531 (N_2531,In_600,In_1606);
nand U2532 (N_2532,In_1681,In_971);
nor U2533 (N_2533,In_1340,In_822);
nand U2534 (N_2534,In_530,In_1253);
nand U2535 (N_2535,In_805,In_1585);
nand U2536 (N_2536,In_734,In_966);
nor U2537 (N_2537,In_563,In_1380);
nor U2538 (N_2538,In_1517,In_832);
and U2539 (N_2539,In_654,In_1294);
nand U2540 (N_2540,In_1685,In_491);
xor U2541 (N_2541,In_1057,In_1938);
nand U2542 (N_2542,In_70,In_1205);
nor U2543 (N_2543,In_1804,In_986);
and U2544 (N_2544,In_1744,In_709);
xnor U2545 (N_2545,In_677,In_1368);
nand U2546 (N_2546,In_1096,In_1372);
nand U2547 (N_2547,In_229,In_248);
nand U2548 (N_2548,In_1499,In_81);
or U2549 (N_2549,In_428,In_634);
or U2550 (N_2550,In_1821,In_1947);
nor U2551 (N_2551,In_1952,In_1016);
nor U2552 (N_2552,In_682,In_1532);
and U2553 (N_2553,In_515,In_687);
or U2554 (N_2554,In_1353,In_1662);
nand U2555 (N_2555,In_486,In_648);
xnor U2556 (N_2556,In_1036,In_591);
xnor U2557 (N_2557,In_491,In_18);
xor U2558 (N_2558,In_1543,In_1728);
nand U2559 (N_2559,In_33,In_311);
nor U2560 (N_2560,In_728,In_932);
nand U2561 (N_2561,In_744,In_320);
or U2562 (N_2562,In_1165,In_618);
or U2563 (N_2563,In_1772,In_1645);
or U2564 (N_2564,In_1693,In_35);
nor U2565 (N_2565,In_336,In_414);
or U2566 (N_2566,In_1829,In_235);
nand U2567 (N_2567,In_1431,In_23);
nand U2568 (N_2568,In_1743,In_1917);
nor U2569 (N_2569,In_1444,In_19);
or U2570 (N_2570,In_77,In_1634);
or U2571 (N_2571,In_953,In_1111);
or U2572 (N_2572,In_1871,In_1787);
or U2573 (N_2573,In_1704,In_1002);
xor U2574 (N_2574,In_276,In_478);
xnor U2575 (N_2575,In_1001,In_1809);
xor U2576 (N_2576,In_222,In_403);
xor U2577 (N_2577,In_1114,In_1771);
nand U2578 (N_2578,In_1557,In_1865);
nor U2579 (N_2579,In_1318,In_1416);
xnor U2580 (N_2580,In_923,In_1311);
nand U2581 (N_2581,In_12,In_715);
nor U2582 (N_2582,In_1431,In_125);
and U2583 (N_2583,In_478,In_1688);
or U2584 (N_2584,In_1784,In_1329);
xor U2585 (N_2585,In_26,In_1487);
and U2586 (N_2586,In_1340,In_411);
nand U2587 (N_2587,In_1376,In_1059);
xor U2588 (N_2588,In_1341,In_1115);
xor U2589 (N_2589,In_1281,In_1151);
or U2590 (N_2590,In_1680,In_1454);
and U2591 (N_2591,In_769,In_696);
and U2592 (N_2592,In_1138,In_337);
nor U2593 (N_2593,In_1433,In_165);
xor U2594 (N_2594,In_760,In_1496);
or U2595 (N_2595,In_576,In_1068);
xor U2596 (N_2596,In_388,In_1960);
or U2597 (N_2597,In_237,In_931);
nand U2598 (N_2598,In_1574,In_1634);
or U2599 (N_2599,In_464,In_839);
and U2600 (N_2600,In_114,In_375);
or U2601 (N_2601,In_953,In_47);
and U2602 (N_2602,In_1117,In_286);
nand U2603 (N_2603,In_1075,In_1337);
nor U2604 (N_2604,In_1932,In_436);
xor U2605 (N_2605,In_982,In_64);
or U2606 (N_2606,In_1856,In_1019);
nand U2607 (N_2607,In_1826,In_1918);
and U2608 (N_2608,In_802,In_816);
or U2609 (N_2609,In_53,In_1917);
or U2610 (N_2610,In_220,In_1936);
or U2611 (N_2611,In_1241,In_1879);
nor U2612 (N_2612,In_997,In_1693);
and U2613 (N_2613,In_1303,In_1914);
nor U2614 (N_2614,In_761,In_1275);
or U2615 (N_2615,In_135,In_511);
nor U2616 (N_2616,In_521,In_84);
nor U2617 (N_2617,In_497,In_248);
nand U2618 (N_2618,In_594,In_1573);
and U2619 (N_2619,In_1199,In_1107);
or U2620 (N_2620,In_161,In_591);
xnor U2621 (N_2621,In_634,In_1197);
and U2622 (N_2622,In_1064,In_1416);
nor U2623 (N_2623,In_107,In_1276);
nand U2624 (N_2624,In_1071,In_777);
or U2625 (N_2625,In_1612,In_57);
xnor U2626 (N_2626,In_575,In_245);
and U2627 (N_2627,In_528,In_1030);
xnor U2628 (N_2628,In_1836,In_408);
and U2629 (N_2629,In_1048,In_1442);
or U2630 (N_2630,In_1892,In_1386);
and U2631 (N_2631,In_972,In_795);
xor U2632 (N_2632,In_989,In_223);
xor U2633 (N_2633,In_48,In_343);
and U2634 (N_2634,In_627,In_1101);
xnor U2635 (N_2635,In_1584,In_1843);
and U2636 (N_2636,In_1295,In_70);
xnor U2637 (N_2637,In_242,In_1125);
nor U2638 (N_2638,In_1160,In_1792);
or U2639 (N_2639,In_35,In_394);
xnor U2640 (N_2640,In_1862,In_1299);
xnor U2641 (N_2641,In_1902,In_698);
or U2642 (N_2642,In_110,In_56);
nand U2643 (N_2643,In_1162,In_641);
or U2644 (N_2644,In_1426,In_11);
xnor U2645 (N_2645,In_413,In_381);
and U2646 (N_2646,In_159,In_887);
nor U2647 (N_2647,In_1260,In_1177);
and U2648 (N_2648,In_1301,In_1755);
and U2649 (N_2649,In_541,In_221);
nor U2650 (N_2650,In_523,In_794);
or U2651 (N_2651,In_103,In_721);
nand U2652 (N_2652,In_722,In_1473);
xor U2653 (N_2653,In_1312,In_153);
nand U2654 (N_2654,In_1809,In_1748);
and U2655 (N_2655,In_588,In_1810);
and U2656 (N_2656,In_1850,In_1394);
nand U2657 (N_2657,In_192,In_1098);
nor U2658 (N_2658,In_182,In_1873);
or U2659 (N_2659,In_356,In_1875);
nor U2660 (N_2660,In_441,In_1097);
nand U2661 (N_2661,In_1282,In_1443);
nand U2662 (N_2662,In_484,In_415);
nor U2663 (N_2663,In_1497,In_1583);
xor U2664 (N_2664,In_1460,In_1600);
xnor U2665 (N_2665,In_1739,In_204);
and U2666 (N_2666,In_1445,In_426);
nand U2667 (N_2667,In_1915,In_1546);
nor U2668 (N_2668,In_1849,In_1679);
nand U2669 (N_2669,In_92,In_1107);
or U2670 (N_2670,In_1744,In_638);
and U2671 (N_2671,In_585,In_152);
xnor U2672 (N_2672,In_673,In_938);
xnor U2673 (N_2673,In_1283,In_827);
nand U2674 (N_2674,In_308,In_126);
and U2675 (N_2675,In_1403,In_673);
nand U2676 (N_2676,In_189,In_1133);
nor U2677 (N_2677,In_70,In_792);
nor U2678 (N_2678,In_1998,In_1787);
and U2679 (N_2679,In_137,In_217);
xnor U2680 (N_2680,In_395,In_1361);
nand U2681 (N_2681,In_1152,In_1325);
nor U2682 (N_2682,In_284,In_940);
and U2683 (N_2683,In_299,In_1576);
or U2684 (N_2684,In_1781,In_1884);
xnor U2685 (N_2685,In_426,In_953);
xor U2686 (N_2686,In_513,In_657);
xnor U2687 (N_2687,In_140,In_1513);
nor U2688 (N_2688,In_1509,In_117);
xor U2689 (N_2689,In_1605,In_1808);
xnor U2690 (N_2690,In_1940,In_236);
or U2691 (N_2691,In_196,In_1770);
xnor U2692 (N_2692,In_541,In_557);
and U2693 (N_2693,In_393,In_644);
nand U2694 (N_2694,In_1573,In_609);
xor U2695 (N_2695,In_678,In_48);
and U2696 (N_2696,In_976,In_1829);
nor U2697 (N_2697,In_636,In_1461);
and U2698 (N_2698,In_926,In_1240);
xor U2699 (N_2699,In_485,In_332);
or U2700 (N_2700,In_1010,In_386);
xor U2701 (N_2701,In_227,In_1823);
or U2702 (N_2702,In_693,In_121);
xor U2703 (N_2703,In_8,In_388);
nand U2704 (N_2704,In_1176,In_681);
and U2705 (N_2705,In_1867,In_1896);
nor U2706 (N_2706,In_349,In_545);
nor U2707 (N_2707,In_1349,In_1739);
nand U2708 (N_2708,In_513,In_1940);
xnor U2709 (N_2709,In_1411,In_833);
or U2710 (N_2710,In_306,In_1436);
nand U2711 (N_2711,In_1198,In_1447);
nor U2712 (N_2712,In_1091,In_533);
nand U2713 (N_2713,In_485,In_1854);
xor U2714 (N_2714,In_82,In_223);
and U2715 (N_2715,In_1986,In_967);
xor U2716 (N_2716,In_965,In_562);
and U2717 (N_2717,In_1398,In_141);
nor U2718 (N_2718,In_246,In_230);
nand U2719 (N_2719,In_1523,In_86);
nand U2720 (N_2720,In_1642,In_369);
xnor U2721 (N_2721,In_7,In_655);
nand U2722 (N_2722,In_534,In_136);
and U2723 (N_2723,In_1802,In_648);
xnor U2724 (N_2724,In_1529,In_1735);
or U2725 (N_2725,In_1054,In_1194);
nor U2726 (N_2726,In_107,In_1646);
or U2727 (N_2727,In_1465,In_664);
xnor U2728 (N_2728,In_950,In_217);
nand U2729 (N_2729,In_192,In_928);
nor U2730 (N_2730,In_757,In_1346);
and U2731 (N_2731,In_582,In_956);
nor U2732 (N_2732,In_535,In_684);
or U2733 (N_2733,In_1166,In_897);
nand U2734 (N_2734,In_1626,In_1409);
xnor U2735 (N_2735,In_1133,In_359);
or U2736 (N_2736,In_1639,In_1756);
xor U2737 (N_2737,In_18,In_52);
nand U2738 (N_2738,In_200,In_1774);
xnor U2739 (N_2739,In_112,In_255);
nor U2740 (N_2740,In_1673,In_1396);
xor U2741 (N_2741,In_1526,In_1049);
nor U2742 (N_2742,In_1384,In_1679);
and U2743 (N_2743,In_1220,In_1454);
xor U2744 (N_2744,In_1149,In_1343);
and U2745 (N_2745,In_1419,In_1599);
or U2746 (N_2746,In_25,In_1014);
and U2747 (N_2747,In_1130,In_1452);
nand U2748 (N_2748,In_1725,In_1153);
xor U2749 (N_2749,In_943,In_1949);
and U2750 (N_2750,In_1417,In_1354);
or U2751 (N_2751,In_987,In_1530);
nand U2752 (N_2752,In_1728,In_834);
nor U2753 (N_2753,In_493,In_1982);
nor U2754 (N_2754,In_1751,In_1914);
and U2755 (N_2755,In_1919,In_362);
xor U2756 (N_2756,In_115,In_202);
or U2757 (N_2757,In_1178,In_578);
and U2758 (N_2758,In_251,In_276);
nor U2759 (N_2759,In_1877,In_729);
xor U2760 (N_2760,In_328,In_1898);
and U2761 (N_2761,In_381,In_1190);
nor U2762 (N_2762,In_291,In_681);
nand U2763 (N_2763,In_613,In_1105);
nor U2764 (N_2764,In_546,In_984);
xnor U2765 (N_2765,In_768,In_1407);
and U2766 (N_2766,In_1994,In_424);
or U2767 (N_2767,In_1579,In_1619);
nand U2768 (N_2768,In_1512,In_1500);
xor U2769 (N_2769,In_1869,In_646);
nor U2770 (N_2770,In_753,In_161);
nor U2771 (N_2771,In_102,In_759);
nor U2772 (N_2772,In_1270,In_450);
or U2773 (N_2773,In_518,In_157);
and U2774 (N_2774,In_1817,In_1772);
or U2775 (N_2775,In_1271,In_1817);
xnor U2776 (N_2776,In_1029,In_348);
or U2777 (N_2777,In_96,In_1568);
xnor U2778 (N_2778,In_1273,In_1514);
xnor U2779 (N_2779,In_712,In_1743);
nor U2780 (N_2780,In_1760,In_680);
xnor U2781 (N_2781,In_216,In_1256);
and U2782 (N_2782,In_474,In_1164);
or U2783 (N_2783,In_610,In_818);
nor U2784 (N_2784,In_732,In_1336);
xnor U2785 (N_2785,In_1960,In_398);
nand U2786 (N_2786,In_912,In_1079);
nor U2787 (N_2787,In_663,In_1592);
or U2788 (N_2788,In_1157,In_273);
xnor U2789 (N_2789,In_1438,In_1367);
and U2790 (N_2790,In_414,In_440);
nor U2791 (N_2791,In_315,In_1528);
or U2792 (N_2792,In_22,In_1651);
or U2793 (N_2793,In_132,In_867);
and U2794 (N_2794,In_1739,In_1095);
nand U2795 (N_2795,In_1252,In_1649);
or U2796 (N_2796,In_1003,In_1510);
or U2797 (N_2797,In_734,In_75);
xnor U2798 (N_2798,In_128,In_726);
nor U2799 (N_2799,In_285,In_979);
and U2800 (N_2800,In_1510,In_1293);
nand U2801 (N_2801,In_539,In_1449);
or U2802 (N_2802,In_513,In_10);
xnor U2803 (N_2803,In_196,In_406);
or U2804 (N_2804,In_1693,In_12);
xor U2805 (N_2805,In_1040,In_46);
nor U2806 (N_2806,In_137,In_1082);
xor U2807 (N_2807,In_11,In_1543);
and U2808 (N_2808,In_1617,In_1810);
nor U2809 (N_2809,In_1536,In_1679);
or U2810 (N_2810,In_1489,In_1682);
nand U2811 (N_2811,In_1852,In_1348);
nor U2812 (N_2812,In_461,In_1590);
or U2813 (N_2813,In_374,In_1827);
nor U2814 (N_2814,In_296,In_70);
nand U2815 (N_2815,In_652,In_263);
and U2816 (N_2816,In_775,In_741);
and U2817 (N_2817,In_1495,In_473);
xor U2818 (N_2818,In_391,In_1639);
nor U2819 (N_2819,In_503,In_176);
xnor U2820 (N_2820,In_306,In_166);
nor U2821 (N_2821,In_347,In_1765);
or U2822 (N_2822,In_1516,In_1128);
and U2823 (N_2823,In_1759,In_828);
and U2824 (N_2824,In_714,In_1052);
and U2825 (N_2825,In_412,In_1347);
or U2826 (N_2826,In_1793,In_519);
xnor U2827 (N_2827,In_160,In_507);
nand U2828 (N_2828,In_1468,In_592);
or U2829 (N_2829,In_1556,In_924);
nand U2830 (N_2830,In_1781,In_1058);
xnor U2831 (N_2831,In_1085,In_559);
xor U2832 (N_2832,In_285,In_1522);
or U2833 (N_2833,In_1246,In_892);
nor U2834 (N_2834,In_648,In_1315);
and U2835 (N_2835,In_131,In_1784);
nor U2836 (N_2836,In_561,In_928);
xnor U2837 (N_2837,In_476,In_1630);
nand U2838 (N_2838,In_779,In_1591);
and U2839 (N_2839,In_1415,In_444);
and U2840 (N_2840,In_1605,In_1634);
xor U2841 (N_2841,In_300,In_1150);
nor U2842 (N_2842,In_1250,In_490);
or U2843 (N_2843,In_1289,In_1545);
xnor U2844 (N_2844,In_1245,In_1892);
or U2845 (N_2845,In_1652,In_1200);
or U2846 (N_2846,In_1454,In_1415);
xor U2847 (N_2847,In_1210,In_795);
nand U2848 (N_2848,In_405,In_730);
or U2849 (N_2849,In_1627,In_158);
or U2850 (N_2850,In_645,In_1296);
nor U2851 (N_2851,In_1957,In_485);
nand U2852 (N_2852,In_1507,In_689);
nor U2853 (N_2853,In_1573,In_29);
nor U2854 (N_2854,In_1438,In_572);
nand U2855 (N_2855,In_610,In_1491);
or U2856 (N_2856,In_1306,In_763);
and U2857 (N_2857,In_1659,In_1426);
and U2858 (N_2858,In_1885,In_414);
or U2859 (N_2859,In_773,In_598);
xnor U2860 (N_2860,In_1456,In_1183);
xnor U2861 (N_2861,In_1060,In_769);
nand U2862 (N_2862,In_7,In_1750);
nor U2863 (N_2863,In_401,In_1928);
and U2864 (N_2864,In_697,In_1543);
and U2865 (N_2865,In_1710,In_1956);
nand U2866 (N_2866,In_436,In_353);
nor U2867 (N_2867,In_1132,In_276);
and U2868 (N_2868,In_926,In_269);
nand U2869 (N_2869,In_1960,In_193);
xnor U2870 (N_2870,In_1160,In_1973);
nand U2871 (N_2871,In_1969,In_4);
xnor U2872 (N_2872,In_663,In_622);
and U2873 (N_2873,In_859,In_1063);
nor U2874 (N_2874,In_491,In_526);
nor U2875 (N_2875,In_629,In_1883);
nand U2876 (N_2876,In_1044,In_1415);
xor U2877 (N_2877,In_1168,In_1271);
xnor U2878 (N_2878,In_614,In_1626);
nor U2879 (N_2879,In_311,In_1131);
nand U2880 (N_2880,In_1759,In_1604);
or U2881 (N_2881,In_1413,In_1106);
xor U2882 (N_2882,In_1529,In_862);
nand U2883 (N_2883,In_966,In_507);
xor U2884 (N_2884,In_457,In_862);
nor U2885 (N_2885,In_1427,In_1884);
and U2886 (N_2886,In_1586,In_851);
nor U2887 (N_2887,In_851,In_724);
nor U2888 (N_2888,In_1985,In_1726);
and U2889 (N_2889,In_1432,In_1852);
xor U2890 (N_2890,In_1016,In_509);
or U2891 (N_2891,In_1853,In_27);
and U2892 (N_2892,In_969,In_1892);
nor U2893 (N_2893,In_1888,In_592);
nand U2894 (N_2894,In_1939,In_737);
and U2895 (N_2895,In_1358,In_1414);
nand U2896 (N_2896,In_966,In_1110);
nand U2897 (N_2897,In_501,In_216);
nor U2898 (N_2898,In_1303,In_1913);
nor U2899 (N_2899,In_263,In_1896);
nor U2900 (N_2900,In_1530,In_594);
and U2901 (N_2901,In_1744,In_1685);
and U2902 (N_2902,In_1976,In_1439);
nand U2903 (N_2903,In_608,In_1570);
xor U2904 (N_2904,In_1230,In_172);
nor U2905 (N_2905,In_41,In_269);
nand U2906 (N_2906,In_1770,In_896);
xnor U2907 (N_2907,In_621,In_1860);
nor U2908 (N_2908,In_431,In_193);
nand U2909 (N_2909,In_1355,In_353);
and U2910 (N_2910,In_676,In_975);
and U2911 (N_2911,In_1785,In_84);
xor U2912 (N_2912,In_1139,In_1199);
nor U2913 (N_2913,In_178,In_1524);
xor U2914 (N_2914,In_238,In_1660);
xnor U2915 (N_2915,In_1312,In_1999);
xor U2916 (N_2916,In_506,In_565);
or U2917 (N_2917,In_718,In_654);
xnor U2918 (N_2918,In_932,In_1030);
nor U2919 (N_2919,In_371,In_1891);
xor U2920 (N_2920,In_1082,In_1689);
and U2921 (N_2921,In_601,In_918);
and U2922 (N_2922,In_1213,In_1370);
or U2923 (N_2923,In_762,In_682);
or U2924 (N_2924,In_905,In_1610);
and U2925 (N_2925,In_755,In_1479);
xnor U2926 (N_2926,In_1044,In_815);
and U2927 (N_2927,In_206,In_556);
nor U2928 (N_2928,In_911,In_9);
nor U2929 (N_2929,In_300,In_1773);
and U2930 (N_2930,In_1198,In_289);
xor U2931 (N_2931,In_1075,In_470);
xnor U2932 (N_2932,In_35,In_1708);
xnor U2933 (N_2933,In_837,In_1083);
or U2934 (N_2934,In_1110,In_1655);
nor U2935 (N_2935,In_827,In_1212);
xnor U2936 (N_2936,In_928,In_1541);
or U2937 (N_2937,In_26,In_756);
nor U2938 (N_2938,In_1981,In_1748);
and U2939 (N_2939,In_1756,In_1582);
and U2940 (N_2940,In_1810,In_1222);
xor U2941 (N_2941,In_761,In_1100);
nand U2942 (N_2942,In_626,In_1027);
and U2943 (N_2943,In_1727,In_619);
xnor U2944 (N_2944,In_430,In_1816);
xnor U2945 (N_2945,In_602,In_126);
nand U2946 (N_2946,In_95,In_252);
nor U2947 (N_2947,In_1479,In_10);
nand U2948 (N_2948,In_1279,In_246);
xor U2949 (N_2949,In_655,In_1709);
and U2950 (N_2950,In_206,In_1113);
or U2951 (N_2951,In_858,In_1566);
and U2952 (N_2952,In_733,In_683);
and U2953 (N_2953,In_1718,In_1198);
nand U2954 (N_2954,In_681,In_1762);
nor U2955 (N_2955,In_1903,In_446);
or U2956 (N_2956,In_468,In_629);
and U2957 (N_2957,In_399,In_1981);
or U2958 (N_2958,In_389,In_801);
and U2959 (N_2959,In_1403,In_883);
nand U2960 (N_2960,In_125,In_1989);
nor U2961 (N_2961,In_1580,In_1886);
or U2962 (N_2962,In_661,In_110);
nor U2963 (N_2963,In_1841,In_996);
nand U2964 (N_2964,In_1362,In_108);
and U2965 (N_2965,In_1503,In_1892);
xor U2966 (N_2966,In_1156,In_1995);
and U2967 (N_2967,In_91,In_967);
nand U2968 (N_2968,In_190,In_1817);
nor U2969 (N_2969,In_555,In_745);
or U2970 (N_2970,In_367,In_217);
and U2971 (N_2971,In_602,In_741);
and U2972 (N_2972,In_899,In_1970);
or U2973 (N_2973,In_997,In_761);
nand U2974 (N_2974,In_1675,In_261);
xor U2975 (N_2975,In_1027,In_598);
nor U2976 (N_2976,In_948,In_1594);
nand U2977 (N_2977,In_1736,In_1573);
nor U2978 (N_2978,In_1391,In_1237);
nand U2979 (N_2979,In_238,In_414);
nor U2980 (N_2980,In_1263,In_1230);
or U2981 (N_2981,In_803,In_1507);
and U2982 (N_2982,In_1468,In_575);
and U2983 (N_2983,In_768,In_1713);
nand U2984 (N_2984,In_890,In_1329);
and U2985 (N_2985,In_1415,In_1968);
or U2986 (N_2986,In_1393,In_1630);
or U2987 (N_2987,In_1272,In_1762);
nor U2988 (N_2988,In_657,In_818);
xnor U2989 (N_2989,In_1741,In_1012);
and U2990 (N_2990,In_1856,In_163);
nor U2991 (N_2991,In_1626,In_131);
and U2992 (N_2992,In_242,In_1094);
and U2993 (N_2993,In_1359,In_1947);
nand U2994 (N_2994,In_682,In_1513);
or U2995 (N_2995,In_1361,In_1415);
xnor U2996 (N_2996,In_99,In_382);
nand U2997 (N_2997,In_1583,In_378);
nand U2998 (N_2998,In_754,In_701);
nor U2999 (N_2999,In_1134,In_198);
nor U3000 (N_3000,In_518,In_564);
and U3001 (N_3001,In_1232,In_1115);
nand U3002 (N_3002,In_1777,In_1716);
nand U3003 (N_3003,In_1646,In_1634);
nand U3004 (N_3004,In_928,In_1327);
and U3005 (N_3005,In_636,In_764);
xor U3006 (N_3006,In_1076,In_1815);
or U3007 (N_3007,In_1596,In_1986);
xor U3008 (N_3008,In_467,In_1633);
and U3009 (N_3009,In_1583,In_1441);
xnor U3010 (N_3010,In_76,In_1437);
or U3011 (N_3011,In_1339,In_1301);
nand U3012 (N_3012,In_807,In_972);
nand U3013 (N_3013,In_1742,In_579);
and U3014 (N_3014,In_1093,In_1336);
xnor U3015 (N_3015,In_197,In_278);
xnor U3016 (N_3016,In_106,In_614);
xor U3017 (N_3017,In_1672,In_647);
nor U3018 (N_3018,In_1790,In_1208);
and U3019 (N_3019,In_1629,In_1840);
xnor U3020 (N_3020,In_1237,In_1549);
xnor U3021 (N_3021,In_829,In_976);
and U3022 (N_3022,In_492,In_128);
and U3023 (N_3023,In_1743,In_1939);
xnor U3024 (N_3024,In_1103,In_1071);
and U3025 (N_3025,In_692,In_851);
and U3026 (N_3026,In_1501,In_1118);
and U3027 (N_3027,In_1028,In_716);
xor U3028 (N_3028,In_1112,In_924);
nand U3029 (N_3029,In_449,In_800);
or U3030 (N_3030,In_939,In_1489);
xor U3031 (N_3031,In_1072,In_355);
nand U3032 (N_3032,In_1024,In_480);
xor U3033 (N_3033,In_1257,In_487);
nand U3034 (N_3034,In_56,In_1075);
nand U3035 (N_3035,In_1122,In_848);
and U3036 (N_3036,In_1899,In_1257);
xnor U3037 (N_3037,In_827,In_86);
xnor U3038 (N_3038,In_59,In_517);
and U3039 (N_3039,In_1750,In_21);
nand U3040 (N_3040,In_567,In_837);
or U3041 (N_3041,In_1534,In_1736);
or U3042 (N_3042,In_1769,In_606);
xnor U3043 (N_3043,In_1232,In_528);
xnor U3044 (N_3044,In_1080,In_230);
xnor U3045 (N_3045,In_1803,In_919);
nor U3046 (N_3046,In_1839,In_583);
nor U3047 (N_3047,In_1548,In_1852);
or U3048 (N_3048,In_748,In_995);
and U3049 (N_3049,In_638,In_629);
or U3050 (N_3050,In_1968,In_525);
nand U3051 (N_3051,In_763,In_1082);
or U3052 (N_3052,In_532,In_910);
xor U3053 (N_3053,In_61,In_8);
nor U3054 (N_3054,In_689,In_1688);
and U3055 (N_3055,In_616,In_153);
xnor U3056 (N_3056,In_410,In_1425);
nand U3057 (N_3057,In_1186,In_646);
xnor U3058 (N_3058,In_1549,In_1867);
and U3059 (N_3059,In_383,In_797);
or U3060 (N_3060,In_472,In_1234);
nor U3061 (N_3061,In_832,In_204);
or U3062 (N_3062,In_450,In_1789);
nand U3063 (N_3063,In_1461,In_783);
xor U3064 (N_3064,In_347,In_129);
or U3065 (N_3065,In_1112,In_631);
nor U3066 (N_3066,In_280,In_223);
nand U3067 (N_3067,In_1965,In_1712);
nor U3068 (N_3068,In_990,In_600);
and U3069 (N_3069,In_232,In_752);
nor U3070 (N_3070,In_384,In_76);
xnor U3071 (N_3071,In_697,In_51);
nand U3072 (N_3072,In_1426,In_868);
and U3073 (N_3073,In_1809,In_1447);
and U3074 (N_3074,In_854,In_454);
and U3075 (N_3075,In_1846,In_806);
nor U3076 (N_3076,In_833,In_1769);
or U3077 (N_3077,In_807,In_1992);
xor U3078 (N_3078,In_132,In_1632);
or U3079 (N_3079,In_1482,In_1215);
nand U3080 (N_3080,In_1137,In_156);
nand U3081 (N_3081,In_209,In_50);
xnor U3082 (N_3082,In_1635,In_707);
nor U3083 (N_3083,In_1070,In_1202);
and U3084 (N_3084,In_558,In_228);
nor U3085 (N_3085,In_1117,In_656);
or U3086 (N_3086,In_412,In_103);
and U3087 (N_3087,In_1460,In_673);
nand U3088 (N_3088,In_1857,In_1707);
nor U3089 (N_3089,In_1775,In_1879);
and U3090 (N_3090,In_549,In_213);
or U3091 (N_3091,In_1066,In_1872);
or U3092 (N_3092,In_804,In_1169);
or U3093 (N_3093,In_62,In_339);
and U3094 (N_3094,In_219,In_1875);
or U3095 (N_3095,In_593,In_1831);
or U3096 (N_3096,In_1731,In_1688);
or U3097 (N_3097,In_1256,In_335);
nand U3098 (N_3098,In_1267,In_1101);
nor U3099 (N_3099,In_1919,In_1537);
xnor U3100 (N_3100,In_1377,In_603);
xnor U3101 (N_3101,In_1378,In_1801);
nand U3102 (N_3102,In_951,In_1756);
nand U3103 (N_3103,In_472,In_676);
or U3104 (N_3104,In_1494,In_881);
nand U3105 (N_3105,In_1354,In_1323);
or U3106 (N_3106,In_1737,In_1484);
xnor U3107 (N_3107,In_48,In_1507);
or U3108 (N_3108,In_1173,In_103);
nand U3109 (N_3109,In_1216,In_356);
and U3110 (N_3110,In_1281,In_620);
and U3111 (N_3111,In_1172,In_1964);
and U3112 (N_3112,In_966,In_1348);
xor U3113 (N_3113,In_1513,In_437);
and U3114 (N_3114,In_1017,In_830);
and U3115 (N_3115,In_824,In_236);
nor U3116 (N_3116,In_316,In_1798);
or U3117 (N_3117,In_1243,In_47);
nor U3118 (N_3118,In_267,In_154);
and U3119 (N_3119,In_1818,In_723);
nor U3120 (N_3120,In_925,In_1046);
nor U3121 (N_3121,In_1983,In_950);
nand U3122 (N_3122,In_64,In_1796);
xnor U3123 (N_3123,In_574,In_90);
nor U3124 (N_3124,In_1838,In_186);
xor U3125 (N_3125,In_1639,In_1948);
xnor U3126 (N_3126,In_1871,In_1370);
or U3127 (N_3127,In_1877,In_1289);
or U3128 (N_3128,In_231,In_951);
and U3129 (N_3129,In_1914,In_775);
nor U3130 (N_3130,In_1182,In_1658);
nor U3131 (N_3131,In_1331,In_1903);
nor U3132 (N_3132,In_151,In_1161);
nor U3133 (N_3133,In_1772,In_1131);
xor U3134 (N_3134,In_1558,In_1936);
and U3135 (N_3135,In_1299,In_232);
nand U3136 (N_3136,In_1883,In_923);
xnor U3137 (N_3137,In_156,In_649);
and U3138 (N_3138,In_210,In_906);
or U3139 (N_3139,In_975,In_1129);
nor U3140 (N_3140,In_1072,In_1263);
xnor U3141 (N_3141,In_1165,In_1236);
nor U3142 (N_3142,In_156,In_1323);
or U3143 (N_3143,In_834,In_30);
nand U3144 (N_3144,In_1358,In_289);
and U3145 (N_3145,In_553,In_1056);
or U3146 (N_3146,In_1004,In_319);
nor U3147 (N_3147,In_1747,In_1243);
or U3148 (N_3148,In_608,In_1921);
xnor U3149 (N_3149,In_504,In_1688);
xnor U3150 (N_3150,In_48,In_1034);
and U3151 (N_3151,In_1954,In_268);
or U3152 (N_3152,In_728,In_901);
or U3153 (N_3153,In_236,In_494);
or U3154 (N_3154,In_1991,In_910);
nand U3155 (N_3155,In_1496,In_46);
nand U3156 (N_3156,In_1739,In_910);
nand U3157 (N_3157,In_874,In_1449);
and U3158 (N_3158,In_323,In_343);
nand U3159 (N_3159,In_341,In_12);
or U3160 (N_3160,In_1913,In_1626);
xnor U3161 (N_3161,In_1754,In_1636);
nor U3162 (N_3162,In_1015,In_2);
nor U3163 (N_3163,In_1630,In_137);
or U3164 (N_3164,In_1549,In_829);
xor U3165 (N_3165,In_892,In_129);
nand U3166 (N_3166,In_1678,In_1093);
or U3167 (N_3167,In_771,In_485);
nand U3168 (N_3168,In_705,In_1319);
xor U3169 (N_3169,In_729,In_1998);
xnor U3170 (N_3170,In_238,In_933);
xnor U3171 (N_3171,In_663,In_1459);
and U3172 (N_3172,In_1097,In_1969);
or U3173 (N_3173,In_359,In_471);
or U3174 (N_3174,In_1751,In_879);
xor U3175 (N_3175,In_1043,In_1003);
nor U3176 (N_3176,In_618,In_22);
or U3177 (N_3177,In_178,In_1636);
nor U3178 (N_3178,In_271,In_127);
xor U3179 (N_3179,In_1417,In_94);
xnor U3180 (N_3180,In_1582,In_1380);
nand U3181 (N_3181,In_581,In_29);
or U3182 (N_3182,In_905,In_251);
and U3183 (N_3183,In_1664,In_739);
xor U3184 (N_3184,In_1674,In_40);
or U3185 (N_3185,In_651,In_460);
xor U3186 (N_3186,In_1542,In_1204);
and U3187 (N_3187,In_1955,In_89);
or U3188 (N_3188,In_1489,In_850);
nor U3189 (N_3189,In_1817,In_784);
and U3190 (N_3190,In_1055,In_1666);
nand U3191 (N_3191,In_884,In_715);
nand U3192 (N_3192,In_819,In_1726);
xor U3193 (N_3193,In_897,In_1995);
nand U3194 (N_3194,In_1418,In_322);
nand U3195 (N_3195,In_1363,In_1931);
nand U3196 (N_3196,In_1180,In_713);
xnor U3197 (N_3197,In_1165,In_925);
xor U3198 (N_3198,In_1577,In_1558);
and U3199 (N_3199,In_778,In_1321);
or U3200 (N_3200,In_158,In_1238);
or U3201 (N_3201,In_6,In_261);
and U3202 (N_3202,In_82,In_1686);
or U3203 (N_3203,In_424,In_845);
or U3204 (N_3204,In_502,In_1048);
and U3205 (N_3205,In_23,In_86);
nand U3206 (N_3206,In_373,In_1541);
xor U3207 (N_3207,In_383,In_319);
nand U3208 (N_3208,In_467,In_1923);
nor U3209 (N_3209,In_363,In_464);
xnor U3210 (N_3210,In_85,In_1022);
nor U3211 (N_3211,In_197,In_880);
or U3212 (N_3212,In_606,In_232);
nor U3213 (N_3213,In_1084,In_915);
xor U3214 (N_3214,In_1216,In_1067);
nor U3215 (N_3215,In_70,In_1857);
or U3216 (N_3216,In_952,In_1473);
or U3217 (N_3217,In_1994,In_421);
nand U3218 (N_3218,In_992,In_1704);
or U3219 (N_3219,In_1505,In_1232);
and U3220 (N_3220,In_1194,In_822);
and U3221 (N_3221,In_674,In_841);
xor U3222 (N_3222,In_1467,In_1808);
or U3223 (N_3223,In_1726,In_843);
nand U3224 (N_3224,In_852,In_1384);
nor U3225 (N_3225,In_882,In_1646);
xor U3226 (N_3226,In_1160,In_258);
nor U3227 (N_3227,In_749,In_1213);
xor U3228 (N_3228,In_111,In_41);
nor U3229 (N_3229,In_813,In_152);
xor U3230 (N_3230,In_1163,In_509);
and U3231 (N_3231,In_624,In_378);
and U3232 (N_3232,In_677,In_786);
xnor U3233 (N_3233,In_1388,In_227);
xnor U3234 (N_3234,In_1993,In_1483);
nor U3235 (N_3235,In_1159,In_1880);
or U3236 (N_3236,In_1725,In_62);
or U3237 (N_3237,In_376,In_917);
xor U3238 (N_3238,In_780,In_208);
xnor U3239 (N_3239,In_503,In_1352);
nand U3240 (N_3240,In_1979,In_1642);
nor U3241 (N_3241,In_1086,In_296);
and U3242 (N_3242,In_1832,In_1047);
and U3243 (N_3243,In_659,In_172);
nor U3244 (N_3244,In_179,In_1743);
xor U3245 (N_3245,In_826,In_149);
or U3246 (N_3246,In_696,In_933);
and U3247 (N_3247,In_855,In_250);
nand U3248 (N_3248,In_1213,In_1388);
nor U3249 (N_3249,In_1391,In_238);
and U3250 (N_3250,In_1643,In_447);
nor U3251 (N_3251,In_967,In_398);
and U3252 (N_3252,In_567,In_359);
xor U3253 (N_3253,In_1516,In_297);
or U3254 (N_3254,In_820,In_1045);
xnor U3255 (N_3255,In_745,In_1324);
nor U3256 (N_3256,In_1629,In_712);
nor U3257 (N_3257,In_996,In_957);
xnor U3258 (N_3258,In_1433,In_1602);
nand U3259 (N_3259,In_1347,In_1159);
nor U3260 (N_3260,In_1942,In_371);
and U3261 (N_3261,In_441,In_1854);
or U3262 (N_3262,In_1007,In_394);
nand U3263 (N_3263,In_495,In_1627);
nor U3264 (N_3264,In_1380,In_353);
or U3265 (N_3265,In_824,In_441);
and U3266 (N_3266,In_1140,In_1950);
xor U3267 (N_3267,In_131,In_1640);
xor U3268 (N_3268,In_1426,In_884);
nand U3269 (N_3269,In_1695,In_1929);
and U3270 (N_3270,In_10,In_283);
nand U3271 (N_3271,In_375,In_749);
or U3272 (N_3272,In_1753,In_811);
or U3273 (N_3273,In_1175,In_1018);
or U3274 (N_3274,In_513,In_1049);
or U3275 (N_3275,In_715,In_953);
or U3276 (N_3276,In_1713,In_1942);
and U3277 (N_3277,In_598,In_908);
or U3278 (N_3278,In_1459,In_1302);
or U3279 (N_3279,In_370,In_937);
and U3280 (N_3280,In_1345,In_1598);
nand U3281 (N_3281,In_246,In_457);
xor U3282 (N_3282,In_1830,In_1481);
and U3283 (N_3283,In_1454,In_157);
and U3284 (N_3284,In_94,In_52);
nor U3285 (N_3285,In_821,In_1612);
or U3286 (N_3286,In_352,In_1602);
or U3287 (N_3287,In_867,In_1467);
and U3288 (N_3288,In_400,In_1970);
nor U3289 (N_3289,In_1871,In_343);
nand U3290 (N_3290,In_580,In_1454);
nand U3291 (N_3291,In_1361,In_105);
xnor U3292 (N_3292,In_798,In_976);
or U3293 (N_3293,In_1597,In_1901);
and U3294 (N_3294,In_1031,In_800);
and U3295 (N_3295,In_1934,In_1854);
or U3296 (N_3296,In_1552,In_1383);
nand U3297 (N_3297,In_197,In_1087);
xor U3298 (N_3298,In_1075,In_94);
and U3299 (N_3299,In_1863,In_1074);
nor U3300 (N_3300,In_707,In_1961);
and U3301 (N_3301,In_636,In_164);
nor U3302 (N_3302,In_1451,In_192);
and U3303 (N_3303,In_1690,In_1941);
or U3304 (N_3304,In_1986,In_741);
nor U3305 (N_3305,In_328,In_763);
nand U3306 (N_3306,In_1414,In_890);
nor U3307 (N_3307,In_582,In_26);
and U3308 (N_3308,In_829,In_1753);
nor U3309 (N_3309,In_1272,In_534);
and U3310 (N_3310,In_1025,In_1919);
or U3311 (N_3311,In_1385,In_204);
nand U3312 (N_3312,In_368,In_13);
or U3313 (N_3313,In_1275,In_477);
and U3314 (N_3314,In_1551,In_609);
xor U3315 (N_3315,In_986,In_696);
or U3316 (N_3316,In_738,In_1120);
xnor U3317 (N_3317,In_60,In_1684);
and U3318 (N_3318,In_1032,In_1299);
nor U3319 (N_3319,In_980,In_1556);
nand U3320 (N_3320,In_246,In_314);
nor U3321 (N_3321,In_484,In_820);
nor U3322 (N_3322,In_722,In_1245);
xor U3323 (N_3323,In_653,In_1113);
xor U3324 (N_3324,In_938,In_1895);
or U3325 (N_3325,In_1449,In_652);
or U3326 (N_3326,In_1072,In_734);
xor U3327 (N_3327,In_1515,In_1105);
nand U3328 (N_3328,In_1389,In_1409);
nor U3329 (N_3329,In_63,In_1501);
xor U3330 (N_3330,In_779,In_1002);
nor U3331 (N_3331,In_403,In_337);
nor U3332 (N_3332,In_854,In_202);
and U3333 (N_3333,In_1950,In_1986);
nor U3334 (N_3334,In_1199,In_645);
or U3335 (N_3335,In_4,In_1773);
nand U3336 (N_3336,In_129,In_639);
xor U3337 (N_3337,In_415,In_1984);
or U3338 (N_3338,In_876,In_234);
or U3339 (N_3339,In_733,In_526);
xnor U3340 (N_3340,In_25,In_116);
xor U3341 (N_3341,In_434,In_1236);
and U3342 (N_3342,In_113,In_1861);
and U3343 (N_3343,In_769,In_1604);
nand U3344 (N_3344,In_1913,In_1581);
nor U3345 (N_3345,In_289,In_1141);
nor U3346 (N_3346,In_1997,In_1478);
and U3347 (N_3347,In_629,In_563);
xor U3348 (N_3348,In_1979,In_905);
xor U3349 (N_3349,In_1225,In_1921);
nand U3350 (N_3350,In_1736,In_974);
xnor U3351 (N_3351,In_1149,In_1409);
nand U3352 (N_3352,In_501,In_1045);
xnor U3353 (N_3353,In_138,In_883);
nand U3354 (N_3354,In_1349,In_502);
xor U3355 (N_3355,In_902,In_1885);
xnor U3356 (N_3356,In_450,In_1765);
nor U3357 (N_3357,In_1873,In_1744);
or U3358 (N_3358,In_1354,In_119);
nor U3359 (N_3359,In_697,In_877);
nand U3360 (N_3360,In_1473,In_1698);
and U3361 (N_3361,In_637,In_566);
and U3362 (N_3362,In_1877,In_1530);
xor U3363 (N_3363,In_1550,In_1983);
nor U3364 (N_3364,In_295,In_1036);
nand U3365 (N_3365,In_419,In_400);
nand U3366 (N_3366,In_1007,In_779);
nand U3367 (N_3367,In_1512,In_1614);
nor U3368 (N_3368,In_1282,In_967);
and U3369 (N_3369,In_1383,In_203);
xor U3370 (N_3370,In_1786,In_1339);
and U3371 (N_3371,In_1318,In_1538);
or U3372 (N_3372,In_84,In_309);
or U3373 (N_3373,In_962,In_1291);
nor U3374 (N_3374,In_723,In_514);
xnor U3375 (N_3375,In_1064,In_241);
xnor U3376 (N_3376,In_1550,In_1159);
and U3377 (N_3377,In_443,In_938);
and U3378 (N_3378,In_259,In_1426);
or U3379 (N_3379,In_928,In_77);
and U3380 (N_3380,In_1330,In_1090);
and U3381 (N_3381,In_1961,In_1570);
nand U3382 (N_3382,In_1351,In_676);
xnor U3383 (N_3383,In_973,In_624);
xor U3384 (N_3384,In_326,In_1121);
and U3385 (N_3385,In_850,In_667);
xor U3386 (N_3386,In_1305,In_240);
or U3387 (N_3387,In_53,In_669);
nor U3388 (N_3388,In_572,In_247);
or U3389 (N_3389,In_1129,In_471);
nand U3390 (N_3390,In_1335,In_575);
nand U3391 (N_3391,In_1220,In_365);
nor U3392 (N_3392,In_238,In_1691);
nand U3393 (N_3393,In_378,In_396);
nor U3394 (N_3394,In_538,In_547);
nand U3395 (N_3395,In_270,In_770);
xnor U3396 (N_3396,In_1620,In_1798);
xor U3397 (N_3397,In_289,In_1554);
nand U3398 (N_3398,In_479,In_1785);
nor U3399 (N_3399,In_538,In_1521);
nor U3400 (N_3400,In_1560,In_1722);
and U3401 (N_3401,In_1178,In_1477);
xor U3402 (N_3402,In_1725,In_319);
and U3403 (N_3403,In_595,In_1110);
and U3404 (N_3404,In_1893,In_1180);
nand U3405 (N_3405,In_598,In_1272);
or U3406 (N_3406,In_906,In_775);
and U3407 (N_3407,In_376,In_139);
or U3408 (N_3408,In_1261,In_1726);
and U3409 (N_3409,In_1352,In_1665);
nor U3410 (N_3410,In_1357,In_1059);
or U3411 (N_3411,In_1937,In_983);
and U3412 (N_3412,In_1927,In_1100);
nand U3413 (N_3413,In_1853,In_1679);
or U3414 (N_3414,In_1267,In_338);
xnor U3415 (N_3415,In_513,In_1656);
or U3416 (N_3416,In_1486,In_88);
nand U3417 (N_3417,In_323,In_73);
and U3418 (N_3418,In_66,In_1142);
xnor U3419 (N_3419,In_117,In_1489);
nand U3420 (N_3420,In_1804,In_1516);
nand U3421 (N_3421,In_889,In_1906);
and U3422 (N_3422,In_1054,In_1945);
nor U3423 (N_3423,In_106,In_1741);
xor U3424 (N_3424,In_29,In_6);
or U3425 (N_3425,In_43,In_1415);
or U3426 (N_3426,In_343,In_519);
and U3427 (N_3427,In_876,In_1720);
and U3428 (N_3428,In_1613,In_62);
xnor U3429 (N_3429,In_1904,In_1608);
xnor U3430 (N_3430,In_1221,In_72);
nor U3431 (N_3431,In_1473,In_1629);
nand U3432 (N_3432,In_1783,In_1639);
xor U3433 (N_3433,In_854,In_636);
and U3434 (N_3434,In_1387,In_1323);
nand U3435 (N_3435,In_214,In_1929);
or U3436 (N_3436,In_1800,In_256);
nor U3437 (N_3437,In_719,In_1346);
nand U3438 (N_3438,In_124,In_1693);
nor U3439 (N_3439,In_1075,In_650);
nand U3440 (N_3440,In_972,In_1647);
xnor U3441 (N_3441,In_157,In_1599);
xnor U3442 (N_3442,In_1588,In_1054);
xnor U3443 (N_3443,In_1009,In_763);
or U3444 (N_3444,In_1350,In_36);
nand U3445 (N_3445,In_1348,In_1857);
or U3446 (N_3446,In_109,In_1978);
and U3447 (N_3447,In_560,In_1520);
xnor U3448 (N_3448,In_265,In_986);
or U3449 (N_3449,In_1374,In_1598);
and U3450 (N_3450,In_1568,In_993);
xor U3451 (N_3451,In_483,In_1433);
or U3452 (N_3452,In_281,In_738);
or U3453 (N_3453,In_923,In_93);
and U3454 (N_3454,In_1569,In_436);
and U3455 (N_3455,In_1478,In_83);
nand U3456 (N_3456,In_169,In_1087);
nand U3457 (N_3457,In_841,In_1784);
or U3458 (N_3458,In_1680,In_444);
nand U3459 (N_3459,In_76,In_1046);
nand U3460 (N_3460,In_1429,In_1444);
nand U3461 (N_3461,In_1214,In_1029);
and U3462 (N_3462,In_376,In_633);
and U3463 (N_3463,In_1597,In_367);
and U3464 (N_3464,In_903,In_1458);
nor U3465 (N_3465,In_1430,In_1456);
and U3466 (N_3466,In_114,In_617);
and U3467 (N_3467,In_1219,In_1475);
or U3468 (N_3468,In_1971,In_109);
nand U3469 (N_3469,In_285,In_450);
xnor U3470 (N_3470,In_1472,In_983);
nand U3471 (N_3471,In_619,In_1521);
and U3472 (N_3472,In_1087,In_1198);
and U3473 (N_3473,In_1853,In_207);
nand U3474 (N_3474,In_1788,In_1211);
xor U3475 (N_3475,In_1147,In_1207);
xor U3476 (N_3476,In_214,In_1295);
or U3477 (N_3477,In_264,In_936);
xnor U3478 (N_3478,In_1326,In_1044);
xnor U3479 (N_3479,In_1730,In_476);
nor U3480 (N_3480,In_1595,In_1801);
nor U3481 (N_3481,In_92,In_384);
xnor U3482 (N_3482,In_1009,In_1316);
nand U3483 (N_3483,In_570,In_275);
xor U3484 (N_3484,In_1401,In_1918);
nand U3485 (N_3485,In_896,In_116);
nand U3486 (N_3486,In_1826,In_478);
or U3487 (N_3487,In_936,In_428);
nand U3488 (N_3488,In_59,In_880);
and U3489 (N_3489,In_1863,In_473);
or U3490 (N_3490,In_477,In_718);
nor U3491 (N_3491,In_1740,In_1229);
or U3492 (N_3492,In_741,In_1460);
nor U3493 (N_3493,In_493,In_1515);
or U3494 (N_3494,In_767,In_247);
and U3495 (N_3495,In_1629,In_958);
or U3496 (N_3496,In_395,In_940);
and U3497 (N_3497,In_1253,In_1103);
nand U3498 (N_3498,In_575,In_851);
and U3499 (N_3499,In_1523,In_1875);
nor U3500 (N_3500,In_551,In_576);
nor U3501 (N_3501,In_1420,In_772);
or U3502 (N_3502,In_1895,In_1092);
nor U3503 (N_3503,In_1137,In_1147);
or U3504 (N_3504,In_1974,In_1109);
or U3505 (N_3505,In_1635,In_816);
or U3506 (N_3506,In_1182,In_174);
nand U3507 (N_3507,In_385,In_661);
xor U3508 (N_3508,In_1320,In_569);
or U3509 (N_3509,In_1756,In_731);
nand U3510 (N_3510,In_1716,In_1851);
nor U3511 (N_3511,In_736,In_1382);
xnor U3512 (N_3512,In_1219,In_77);
xor U3513 (N_3513,In_1497,In_1820);
nor U3514 (N_3514,In_317,In_1958);
or U3515 (N_3515,In_903,In_230);
nand U3516 (N_3516,In_1411,In_1332);
nand U3517 (N_3517,In_1557,In_1602);
and U3518 (N_3518,In_1426,In_1494);
or U3519 (N_3519,In_337,In_842);
or U3520 (N_3520,In_1256,In_583);
nor U3521 (N_3521,In_606,In_548);
and U3522 (N_3522,In_1879,In_759);
nor U3523 (N_3523,In_245,In_652);
or U3524 (N_3524,In_1295,In_1964);
xnor U3525 (N_3525,In_366,In_724);
or U3526 (N_3526,In_799,In_1666);
and U3527 (N_3527,In_419,In_979);
xor U3528 (N_3528,In_1917,In_1853);
and U3529 (N_3529,In_1385,In_807);
or U3530 (N_3530,In_1523,In_152);
nor U3531 (N_3531,In_175,In_464);
nor U3532 (N_3532,In_1365,In_831);
and U3533 (N_3533,In_1287,In_679);
nor U3534 (N_3534,In_684,In_575);
or U3535 (N_3535,In_1767,In_1844);
or U3536 (N_3536,In_987,In_1345);
nand U3537 (N_3537,In_895,In_1416);
nand U3538 (N_3538,In_405,In_1495);
nand U3539 (N_3539,In_1135,In_365);
and U3540 (N_3540,In_1576,In_916);
or U3541 (N_3541,In_1050,In_1799);
or U3542 (N_3542,In_1275,In_1939);
or U3543 (N_3543,In_1747,In_930);
nand U3544 (N_3544,In_1120,In_403);
and U3545 (N_3545,In_1869,In_584);
nand U3546 (N_3546,In_1725,In_464);
and U3547 (N_3547,In_493,In_1166);
nand U3548 (N_3548,In_679,In_1645);
nand U3549 (N_3549,In_1159,In_687);
and U3550 (N_3550,In_1014,In_1383);
or U3551 (N_3551,In_367,In_1564);
and U3552 (N_3552,In_1062,In_504);
nor U3553 (N_3553,In_1613,In_1136);
and U3554 (N_3554,In_1103,In_260);
xor U3555 (N_3555,In_186,In_884);
and U3556 (N_3556,In_823,In_1902);
nand U3557 (N_3557,In_1206,In_347);
and U3558 (N_3558,In_272,In_1336);
or U3559 (N_3559,In_1683,In_290);
and U3560 (N_3560,In_391,In_1841);
or U3561 (N_3561,In_1398,In_1275);
xnor U3562 (N_3562,In_1028,In_825);
or U3563 (N_3563,In_151,In_289);
nor U3564 (N_3564,In_358,In_1933);
and U3565 (N_3565,In_1366,In_1116);
nand U3566 (N_3566,In_1579,In_1529);
or U3567 (N_3567,In_1822,In_444);
nand U3568 (N_3568,In_613,In_1268);
nand U3569 (N_3569,In_560,In_510);
xnor U3570 (N_3570,In_1611,In_551);
nor U3571 (N_3571,In_1958,In_1611);
and U3572 (N_3572,In_1650,In_1302);
or U3573 (N_3573,In_1728,In_1973);
xnor U3574 (N_3574,In_1421,In_601);
nor U3575 (N_3575,In_1226,In_819);
and U3576 (N_3576,In_1319,In_1249);
or U3577 (N_3577,In_1575,In_519);
nor U3578 (N_3578,In_1007,In_1864);
xnor U3579 (N_3579,In_1030,In_211);
xor U3580 (N_3580,In_1317,In_149);
nor U3581 (N_3581,In_431,In_1686);
xnor U3582 (N_3582,In_644,In_1298);
or U3583 (N_3583,In_1176,In_943);
nand U3584 (N_3584,In_595,In_1779);
nand U3585 (N_3585,In_556,In_34);
xnor U3586 (N_3586,In_765,In_1162);
nor U3587 (N_3587,In_1462,In_573);
xnor U3588 (N_3588,In_815,In_931);
xor U3589 (N_3589,In_232,In_1242);
and U3590 (N_3590,In_917,In_172);
or U3591 (N_3591,In_1042,In_309);
and U3592 (N_3592,In_415,In_1763);
nand U3593 (N_3593,In_1957,In_1081);
nand U3594 (N_3594,In_680,In_1242);
nand U3595 (N_3595,In_1938,In_568);
or U3596 (N_3596,In_963,In_1086);
nor U3597 (N_3597,In_491,In_365);
xor U3598 (N_3598,In_238,In_1677);
and U3599 (N_3599,In_967,In_573);
and U3600 (N_3600,In_1838,In_460);
xor U3601 (N_3601,In_419,In_415);
nor U3602 (N_3602,In_1132,In_848);
or U3603 (N_3603,In_1723,In_550);
xor U3604 (N_3604,In_745,In_1203);
nor U3605 (N_3605,In_648,In_71);
nor U3606 (N_3606,In_1048,In_769);
nor U3607 (N_3607,In_128,In_457);
nor U3608 (N_3608,In_1817,In_1096);
and U3609 (N_3609,In_864,In_1208);
nor U3610 (N_3610,In_868,In_1708);
or U3611 (N_3611,In_656,In_125);
xnor U3612 (N_3612,In_632,In_1168);
and U3613 (N_3613,In_1368,In_1269);
or U3614 (N_3614,In_198,In_1044);
and U3615 (N_3615,In_812,In_737);
nand U3616 (N_3616,In_27,In_221);
and U3617 (N_3617,In_1464,In_1425);
xnor U3618 (N_3618,In_556,In_763);
nand U3619 (N_3619,In_1553,In_710);
or U3620 (N_3620,In_1762,In_845);
xor U3621 (N_3621,In_355,In_903);
and U3622 (N_3622,In_1924,In_704);
or U3623 (N_3623,In_231,In_762);
or U3624 (N_3624,In_913,In_1422);
nor U3625 (N_3625,In_1114,In_1312);
or U3626 (N_3626,In_1831,In_95);
nand U3627 (N_3627,In_281,In_1211);
nor U3628 (N_3628,In_1584,In_1077);
or U3629 (N_3629,In_1217,In_1300);
nand U3630 (N_3630,In_51,In_1060);
nand U3631 (N_3631,In_1347,In_1058);
nor U3632 (N_3632,In_171,In_725);
or U3633 (N_3633,In_1653,In_984);
nor U3634 (N_3634,In_1622,In_311);
and U3635 (N_3635,In_315,In_1349);
xor U3636 (N_3636,In_484,In_8);
or U3637 (N_3637,In_724,In_215);
and U3638 (N_3638,In_906,In_1501);
xor U3639 (N_3639,In_1820,In_180);
nor U3640 (N_3640,In_659,In_1804);
and U3641 (N_3641,In_1130,In_1508);
nor U3642 (N_3642,In_1553,In_29);
and U3643 (N_3643,In_294,In_1314);
or U3644 (N_3644,In_1912,In_884);
nand U3645 (N_3645,In_677,In_1626);
nand U3646 (N_3646,In_257,In_413);
nor U3647 (N_3647,In_167,In_1834);
nor U3648 (N_3648,In_1621,In_1386);
xnor U3649 (N_3649,In_368,In_1388);
nor U3650 (N_3650,In_1537,In_693);
and U3651 (N_3651,In_684,In_1868);
xor U3652 (N_3652,In_1660,In_1735);
xnor U3653 (N_3653,In_1632,In_329);
xnor U3654 (N_3654,In_538,In_1920);
and U3655 (N_3655,In_1867,In_1531);
xnor U3656 (N_3656,In_1864,In_1594);
and U3657 (N_3657,In_1988,In_914);
xnor U3658 (N_3658,In_114,In_1646);
or U3659 (N_3659,In_382,In_153);
or U3660 (N_3660,In_1778,In_748);
nand U3661 (N_3661,In_190,In_608);
nor U3662 (N_3662,In_890,In_1559);
nand U3663 (N_3663,In_31,In_1807);
or U3664 (N_3664,In_104,In_1464);
or U3665 (N_3665,In_956,In_1586);
nor U3666 (N_3666,In_1909,In_624);
nor U3667 (N_3667,In_1929,In_1251);
nand U3668 (N_3668,In_1228,In_870);
or U3669 (N_3669,In_1040,In_615);
xnor U3670 (N_3670,In_457,In_1512);
nor U3671 (N_3671,In_1002,In_228);
and U3672 (N_3672,In_820,In_515);
nor U3673 (N_3673,In_1295,In_1220);
or U3674 (N_3674,In_800,In_1247);
and U3675 (N_3675,In_695,In_713);
nand U3676 (N_3676,In_54,In_14);
nand U3677 (N_3677,In_1466,In_594);
nand U3678 (N_3678,In_1911,In_761);
nor U3679 (N_3679,In_1120,In_180);
nand U3680 (N_3680,In_1449,In_43);
nor U3681 (N_3681,In_863,In_66);
and U3682 (N_3682,In_726,In_1276);
nor U3683 (N_3683,In_1503,In_479);
and U3684 (N_3684,In_1449,In_173);
and U3685 (N_3685,In_1946,In_597);
xnor U3686 (N_3686,In_99,In_421);
and U3687 (N_3687,In_1007,In_1745);
nand U3688 (N_3688,In_1344,In_1048);
xnor U3689 (N_3689,In_1853,In_407);
and U3690 (N_3690,In_1956,In_1792);
nor U3691 (N_3691,In_635,In_1307);
or U3692 (N_3692,In_1578,In_1630);
nand U3693 (N_3693,In_1127,In_71);
nor U3694 (N_3694,In_470,In_1120);
and U3695 (N_3695,In_1404,In_1011);
and U3696 (N_3696,In_1944,In_706);
nand U3697 (N_3697,In_838,In_370);
xor U3698 (N_3698,In_766,In_740);
or U3699 (N_3699,In_560,In_1235);
or U3700 (N_3700,In_1779,In_1762);
nor U3701 (N_3701,In_776,In_16);
and U3702 (N_3702,In_230,In_197);
or U3703 (N_3703,In_5,In_720);
xnor U3704 (N_3704,In_86,In_856);
or U3705 (N_3705,In_1147,In_1350);
nand U3706 (N_3706,In_46,In_1719);
xnor U3707 (N_3707,In_402,In_395);
xnor U3708 (N_3708,In_264,In_1758);
nand U3709 (N_3709,In_748,In_1892);
nor U3710 (N_3710,In_1091,In_1292);
or U3711 (N_3711,In_440,In_748);
xor U3712 (N_3712,In_1263,In_52);
nand U3713 (N_3713,In_1462,In_231);
xor U3714 (N_3714,In_592,In_279);
or U3715 (N_3715,In_772,In_1845);
nor U3716 (N_3716,In_1789,In_53);
nand U3717 (N_3717,In_942,In_792);
nor U3718 (N_3718,In_1936,In_1039);
nor U3719 (N_3719,In_256,In_1916);
or U3720 (N_3720,In_191,In_1789);
and U3721 (N_3721,In_1788,In_610);
xor U3722 (N_3722,In_872,In_1910);
xor U3723 (N_3723,In_1628,In_1069);
xor U3724 (N_3724,In_1237,In_294);
or U3725 (N_3725,In_1055,In_135);
nor U3726 (N_3726,In_99,In_1978);
or U3727 (N_3727,In_202,In_1729);
and U3728 (N_3728,In_442,In_79);
and U3729 (N_3729,In_803,In_297);
nor U3730 (N_3730,In_1982,In_987);
and U3731 (N_3731,In_1259,In_1369);
xor U3732 (N_3732,In_1533,In_368);
nand U3733 (N_3733,In_924,In_91);
or U3734 (N_3734,In_838,In_815);
and U3735 (N_3735,In_1612,In_240);
nor U3736 (N_3736,In_1476,In_1955);
nor U3737 (N_3737,In_1665,In_1244);
and U3738 (N_3738,In_1193,In_1967);
and U3739 (N_3739,In_1339,In_1783);
xnor U3740 (N_3740,In_33,In_1851);
or U3741 (N_3741,In_1325,In_1626);
nand U3742 (N_3742,In_1136,In_881);
or U3743 (N_3743,In_1877,In_1558);
or U3744 (N_3744,In_440,In_1202);
and U3745 (N_3745,In_246,In_174);
xnor U3746 (N_3746,In_897,In_1882);
and U3747 (N_3747,In_1138,In_722);
and U3748 (N_3748,In_432,In_1510);
or U3749 (N_3749,In_564,In_555);
nor U3750 (N_3750,In_1384,In_339);
nand U3751 (N_3751,In_388,In_1743);
xor U3752 (N_3752,In_614,In_15);
nor U3753 (N_3753,In_1797,In_84);
nand U3754 (N_3754,In_1873,In_586);
xor U3755 (N_3755,In_246,In_1630);
and U3756 (N_3756,In_62,In_1203);
nand U3757 (N_3757,In_809,In_1524);
xnor U3758 (N_3758,In_1465,In_885);
and U3759 (N_3759,In_731,In_1029);
nor U3760 (N_3760,In_172,In_1485);
nor U3761 (N_3761,In_1208,In_1954);
and U3762 (N_3762,In_656,In_152);
nand U3763 (N_3763,In_769,In_306);
and U3764 (N_3764,In_1189,In_1696);
and U3765 (N_3765,In_1156,In_1198);
and U3766 (N_3766,In_1829,In_1451);
xnor U3767 (N_3767,In_693,In_1742);
and U3768 (N_3768,In_1237,In_275);
xnor U3769 (N_3769,In_1109,In_305);
or U3770 (N_3770,In_634,In_279);
nand U3771 (N_3771,In_1995,In_738);
nand U3772 (N_3772,In_158,In_744);
nor U3773 (N_3773,In_1478,In_1135);
and U3774 (N_3774,In_249,In_1894);
xnor U3775 (N_3775,In_633,In_1020);
or U3776 (N_3776,In_1654,In_1927);
xnor U3777 (N_3777,In_594,In_179);
nor U3778 (N_3778,In_152,In_1195);
nor U3779 (N_3779,In_671,In_174);
or U3780 (N_3780,In_683,In_1441);
nor U3781 (N_3781,In_497,In_1732);
nor U3782 (N_3782,In_1078,In_340);
and U3783 (N_3783,In_405,In_1490);
and U3784 (N_3784,In_596,In_1745);
xor U3785 (N_3785,In_1750,In_1092);
nand U3786 (N_3786,In_894,In_1844);
nand U3787 (N_3787,In_1149,In_1197);
or U3788 (N_3788,In_6,In_1519);
or U3789 (N_3789,In_1433,In_612);
xor U3790 (N_3790,In_1348,In_996);
xor U3791 (N_3791,In_557,In_1992);
nor U3792 (N_3792,In_1293,In_1747);
nand U3793 (N_3793,In_883,In_529);
and U3794 (N_3794,In_43,In_585);
and U3795 (N_3795,In_1885,In_1707);
nand U3796 (N_3796,In_695,In_1188);
nor U3797 (N_3797,In_1519,In_1623);
xor U3798 (N_3798,In_1489,In_548);
or U3799 (N_3799,In_1719,In_459);
xor U3800 (N_3800,In_1547,In_1024);
nor U3801 (N_3801,In_1959,In_832);
xor U3802 (N_3802,In_888,In_1618);
xnor U3803 (N_3803,In_1620,In_144);
xor U3804 (N_3804,In_921,In_381);
nand U3805 (N_3805,In_284,In_820);
nand U3806 (N_3806,In_1245,In_89);
and U3807 (N_3807,In_1489,In_104);
xor U3808 (N_3808,In_1751,In_1245);
and U3809 (N_3809,In_1081,In_1650);
or U3810 (N_3810,In_244,In_847);
nand U3811 (N_3811,In_500,In_1830);
nand U3812 (N_3812,In_1409,In_1356);
and U3813 (N_3813,In_474,In_1688);
nand U3814 (N_3814,In_471,In_1075);
xor U3815 (N_3815,In_1355,In_101);
nand U3816 (N_3816,In_557,In_1542);
xnor U3817 (N_3817,In_1423,In_1793);
nand U3818 (N_3818,In_258,In_1517);
nor U3819 (N_3819,In_716,In_915);
and U3820 (N_3820,In_1158,In_1857);
nand U3821 (N_3821,In_1867,In_1332);
nor U3822 (N_3822,In_70,In_1591);
nor U3823 (N_3823,In_175,In_657);
xnor U3824 (N_3824,In_477,In_1077);
and U3825 (N_3825,In_88,In_8);
and U3826 (N_3826,In_919,In_1007);
nor U3827 (N_3827,In_523,In_574);
or U3828 (N_3828,In_866,In_466);
xor U3829 (N_3829,In_1752,In_772);
xnor U3830 (N_3830,In_132,In_40);
and U3831 (N_3831,In_1013,In_897);
nor U3832 (N_3832,In_290,In_1274);
and U3833 (N_3833,In_1306,In_1617);
nor U3834 (N_3834,In_613,In_118);
nor U3835 (N_3835,In_842,In_454);
xor U3836 (N_3836,In_691,In_1626);
xnor U3837 (N_3837,In_680,In_693);
nor U3838 (N_3838,In_1799,In_161);
xor U3839 (N_3839,In_1552,In_1550);
or U3840 (N_3840,In_1720,In_481);
nor U3841 (N_3841,In_1222,In_1069);
nor U3842 (N_3842,In_1919,In_130);
or U3843 (N_3843,In_705,In_931);
nor U3844 (N_3844,In_24,In_1607);
xnor U3845 (N_3845,In_996,In_1860);
nor U3846 (N_3846,In_451,In_1189);
or U3847 (N_3847,In_1320,In_1182);
or U3848 (N_3848,In_480,In_243);
xnor U3849 (N_3849,In_407,In_830);
nor U3850 (N_3850,In_1646,In_1655);
or U3851 (N_3851,In_1544,In_992);
nor U3852 (N_3852,In_1343,In_26);
or U3853 (N_3853,In_1576,In_1910);
or U3854 (N_3854,In_1766,In_1942);
nand U3855 (N_3855,In_919,In_379);
nand U3856 (N_3856,In_690,In_747);
nor U3857 (N_3857,In_952,In_1305);
nand U3858 (N_3858,In_162,In_527);
nor U3859 (N_3859,In_558,In_1553);
nand U3860 (N_3860,In_1446,In_1895);
and U3861 (N_3861,In_60,In_1021);
and U3862 (N_3862,In_242,In_633);
nand U3863 (N_3863,In_1129,In_1896);
and U3864 (N_3864,In_739,In_1015);
or U3865 (N_3865,In_270,In_1831);
and U3866 (N_3866,In_1487,In_892);
and U3867 (N_3867,In_399,In_1068);
or U3868 (N_3868,In_1166,In_1443);
nand U3869 (N_3869,In_1915,In_1772);
nor U3870 (N_3870,In_352,In_1951);
nand U3871 (N_3871,In_1198,In_1911);
nand U3872 (N_3872,In_1323,In_299);
xor U3873 (N_3873,In_1771,In_1598);
nor U3874 (N_3874,In_429,In_689);
nand U3875 (N_3875,In_1611,In_900);
and U3876 (N_3876,In_734,In_1931);
nor U3877 (N_3877,In_888,In_181);
or U3878 (N_3878,In_1818,In_650);
or U3879 (N_3879,In_870,In_653);
and U3880 (N_3880,In_109,In_862);
nand U3881 (N_3881,In_1040,In_1636);
nand U3882 (N_3882,In_1704,In_1274);
and U3883 (N_3883,In_173,In_1041);
nand U3884 (N_3884,In_732,In_589);
xor U3885 (N_3885,In_1887,In_1535);
nor U3886 (N_3886,In_158,In_114);
xor U3887 (N_3887,In_1574,In_569);
xor U3888 (N_3888,In_1512,In_1671);
nor U3889 (N_3889,In_1293,In_287);
nand U3890 (N_3890,In_140,In_584);
xor U3891 (N_3891,In_1258,In_1867);
xor U3892 (N_3892,In_734,In_1582);
nand U3893 (N_3893,In_834,In_1024);
and U3894 (N_3894,In_1438,In_103);
or U3895 (N_3895,In_1887,In_943);
nor U3896 (N_3896,In_1758,In_614);
nand U3897 (N_3897,In_1404,In_1789);
nor U3898 (N_3898,In_598,In_335);
nand U3899 (N_3899,In_1246,In_1244);
nor U3900 (N_3900,In_1502,In_258);
nor U3901 (N_3901,In_1849,In_380);
and U3902 (N_3902,In_1077,In_576);
nor U3903 (N_3903,In_859,In_839);
and U3904 (N_3904,In_555,In_322);
xor U3905 (N_3905,In_1898,In_1589);
nand U3906 (N_3906,In_1009,In_666);
xnor U3907 (N_3907,In_188,In_1216);
and U3908 (N_3908,In_1674,In_1924);
xor U3909 (N_3909,In_1095,In_1558);
nor U3910 (N_3910,In_855,In_201);
xnor U3911 (N_3911,In_1019,In_1095);
and U3912 (N_3912,In_1318,In_1492);
xor U3913 (N_3913,In_809,In_1080);
nand U3914 (N_3914,In_1315,In_1655);
nand U3915 (N_3915,In_404,In_1709);
xnor U3916 (N_3916,In_222,In_1020);
or U3917 (N_3917,In_495,In_777);
nand U3918 (N_3918,In_1678,In_212);
nor U3919 (N_3919,In_1136,In_1179);
and U3920 (N_3920,In_1913,In_131);
nand U3921 (N_3921,In_695,In_633);
nand U3922 (N_3922,In_166,In_285);
nand U3923 (N_3923,In_613,In_1662);
nand U3924 (N_3924,In_1949,In_526);
nor U3925 (N_3925,In_1716,In_1261);
and U3926 (N_3926,In_147,In_366);
and U3927 (N_3927,In_1883,In_1863);
nand U3928 (N_3928,In_1949,In_208);
nor U3929 (N_3929,In_826,In_492);
nand U3930 (N_3930,In_1442,In_1065);
and U3931 (N_3931,In_1071,In_128);
or U3932 (N_3932,In_741,In_950);
xnor U3933 (N_3933,In_1774,In_1831);
xor U3934 (N_3934,In_1167,In_1828);
and U3935 (N_3935,In_1144,In_400);
nor U3936 (N_3936,In_1685,In_575);
nor U3937 (N_3937,In_693,In_1212);
nor U3938 (N_3938,In_721,In_1535);
or U3939 (N_3939,In_1889,In_1963);
nand U3940 (N_3940,In_1317,In_559);
nor U3941 (N_3941,In_432,In_1888);
xor U3942 (N_3942,In_104,In_164);
nand U3943 (N_3943,In_156,In_1211);
nor U3944 (N_3944,In_383,In_1201);
xor U3945 (N_3945,In_90,In_1583);
nand U3946 (N_3946,In_1953,In_1704);
nor U3947 (N_3947,In_559,In_1654);
nor U3948 (N_3948,In_788,In_1060);
xnor U3949 (N_3949,In_1715,In_1079);
or U3950 (N_3950,In_1891,In_222);
xor U3951 (N_3951,In_491,In_85);
or U3952 (N_3952,In_1168,In_1966);
xor U3953 (N_3953,In_1638,In_223);
or U3954 (N_3954,In_1744,In_1930);
or U3955 (N_3955,In_110,In_26);
xnor U3956 (N_3956,In_1323,In_181);
or U3957 (N_3957,In_337,In_960);
and U3958 (N_3958,In_1476,In_116);
or U3959 (N_3959,In_539,In_1364);
xor U3960 (N_3960,In_285,In_1152);
xnor U3961 (N_3961,In_1748,In_701);
nand U3962 (N_3962,In_237,In_154);
or U3963 (N_3963,In_1170,In_95);
nor U3964 (N_3964,In_1670,In_1560);
or U3965 (N_3965,In_668,In_163);
or U3966 (N_3966,In_1762,In_417);
nand U3967 (N_3967,In_1145,In_111);
nand U3968 (N_3968,In_1799,In_1997);
xor U3969 (N_3969,In_1368,In_1793);
and U3970 (N_3970,In_959,In_1855);
or U3971 (N_3971,In_1038,In_1212);
nor U3972 (N_3972,In_1934,In_1449);
and U3973 (N_3973,In_1760,In_1214);
or U3974 (N_3974,In_1045,In_33);
and U3975 (N_3975,In_1700,In_1783);
nor U3976 (N_3976,In_1898,In_1046);
nor U3977 (N_3977,In_1001,In_1298);
nand U3978 (N_3978,In_149,In_362);
xnor U3979 (N_3979,In_1953,In_1125);
nand U3980 (N_3980,In_1557,In_1104);
or U3981 (N_3981,In_1111,In_136);
and U3982 (N_3982,In_424,In_456);
or U3983 (N_3983,In_1289,In_363);
nand U3984 (N_3984,In_864,In_1168);
and U3985 (N_3985,In_1071,In_317);
nor U3986 (N_3986,In_424,In_1864);
nor U3987 (N_3987,In_1096,In_1364);
nor U3988 (N_3988,In_1710,In_1536);
nand U3989 (N_3989,In_1940,In_442);
nand U3990 (N_3990,In_213,In_1725);
nand U3991 (N_3991,In_1174,In_1753);
and U3992 (N_3992,In_1165,In_813);
nor U3993 (N_3993,In_468,In_1184);
xor U3994 (N_3994,In_1221,In_641);
nand U3995 (N_3995,In_1841,In_1104);
nand U3996 (N_3996,In_147,In_123);
and U3997 (N_3997,In_349,In_1087);
xnor U3998 (N_3998,In_1801,In_1890);
nand U3999 (N_3999,In_1252,In_1145);
xor U4000 (N_4000,In_1076,In_1624);
or U4001 (N_4001,In_109,In_272);
and U4002 (N_4002,In_1924,In_927);
nand U4003 (N_4003,In_1087,In_215);
and U4004 (N_4004,In_1503,In_1013);
nand U4005 (N_4005,In_628,In_1163);
xor U4006 (N_4006,In_415,In_1124);
and U4007 (N_4007,In_1060,In_351);
or U4008 (N_4008,In_1331,In_1445);
nor U4009 (N_4009,In_19,In_1494);
nand U4010 (N_4010,In_1328,In_188);
and U4011 (N_4011,In_1202,In_878);
nor U4012 (N_4012,In_1722,In_1859);
nand U4013 (N_4013,In_168,In_654);
nand U4014 (N_4014,In_1089,In_776);
nor U4015 (N_4015,In_0,In_1096);
nand U4016 (N_4016,In_1201,In_418);
nand U4017 (N_4017,In_1149,In_502);
and U4018 (N_4018,In_592,In_46);
nor U4019 (N_4019,In_685,In_196);
xnor U4020 (N_4020,In_750,In_622);
and U4021 (N_4021,In_569,In_1323);
nand U4022 (N_4022,In_863,In_428);
and U4023 (N_4023,In_399,In_1915);
nand U4024 (N_4024,In_1451,In_499);
or U4025 (N_4025,In_1520,In_1623);
and U4026 (N_4026,In_436,In_340);
xnor U4027 (N_4027,In_1874,In_1098);
nand U4028 (N_4028,In_469,In_13);
or U4029 (N_4029,In_1588,In_1996);
xor U4030 (N_4030,In_1098,In_1636);
nand U4031 (N_4031,In_1297,In_961);
or U4032 (N_4032,In_987,In_792);
nand U4033 (N_4033,In_260,In_163);
nand U4034 (N_4034,In_1049,In_1876);
nand U4035 (N_4035,In_803,In_1086);
nor U4036 (N_4036,In_1912,In_251);
nor U4037 (N_4037,In_635,In_745);
and U4038 (N_4038,In_1878,In_1051);
xor U4039 (N_4039,In_865,In_701);
xor U4040 (N_4040,In_1411,In_1461);
or U4041 (N_4041,In_961,In_1033);
or U4042 (N_4042,In_503,In_1265);
nor U4043 (N_4043,In_361,In_1812);
or U4044 (N_4044,In_96,In_985);
and U4045 (N_4045,In_1733,In_703);
nand U4046 (N_4046,In_575,In_932);
xnor U4047 (N_4047,In_216,In_1184);
or U4048 (N_4048,In_1543,In_1287);
nand U4049 (N_4049,In_840,In_1179);
and U4050 (N_4050,In_450,In_733);
and U4051 (N_4051,In_767,In_439);
or U4052 (N_4052,In_1043,In_693);
xnor U4053 (N_4053,In_766,In_1484);
nor U4054 (N_4054,In_937,In_138);
or U4055 (N_4055,In_1613,In_1413);
and U4056 (N_4056,In_1747,In_222);
nand U4057 (N_4057,In_1964,In_378);
and U4058 (N_4058,In_592,In_418);
xor U4059 (N_4059,In_1715,In_759);
xnor U4060 (N_4060,In_437,In_1060);
nor U4061 (N_4061,In_1347,In_184);
nor U4062 (N_4062,In_651,In_740);
nor U4063 (N_4063,In_1856,In_821);
nand U4064 (N_4064,In_1631,In_1685);
xnor U4065 (N_4065,In_274,In_1929);
or U4066 (N_4066,In_1198,In_1784);
nand U4067 (N_4067,In_240,In_118);
and U4068 (N_4068,In_1335,In_1342);
nand U4069 (N_4069,In_1352,In_792);
or U4070 (N_4070,In_1531,In_1609);
xnor U4071 (N_4071,In_1586,In_173);
nor U4072 (N_4072,In_1864,In_463);
nand U4073 (N_4073,In_358,In_1562);
nand U4074 (N_4074,In_1229,In_1190);
xnor U4075 (N_4075,In_487,In_518);
xnor U4076 (N_4076,In_854,In_1869);
nor U4077 (N_4077,In_422,In_1445);
nand U4078 (N_4078,In_1490,In_397);
or U4079 (N_4079,In_700,In_24);
nor U4080 (N_4080,In_765,In_156);
or U4081 (N_4081,In_420,In_424);
xor U4082 (N_4082,In_583,In_1688);
nor U4083 (N_4083,In_521,In_1263);
nor U4084 (N_4084,In_894,In_1082);
or U4085 (N_4085,In_504,In_115);
nand U4086 (N_4086,In_1313,In_89);
nor U4087 (N_4087,In_1821,In_1459);
or U4088 (N_4088,In_60,In_1327);
nor U4089 (N_4089,In_1769,In_727);
nor U4090 (N_4090,In_1238,In_1009);
nor U4091 (N_4091,In_1805,In_1921);
xor U4092 (N_4092,In_1770,In_1843);
and U4093 (N_4093,In_602,In_1899);
and U4094 (N_4094,In_1924,In_15);
nand U4095 (N_4095,In_876,In_1572);
and U4096 (N_4096,In_491,In_98);
or U4097 (N_4097,In_309,In_1124);
or U4098 (N_4098,In_836,In_1964);
nand U4099 (N_4099,In_701,In_655);
nor U4100 (N_4100,In_461,In_239);
nand U4101 (N_4101,In_510,In_1930);
and U4102 (N_4102,In_607,In_908);
xnor U4103 (N_4103,In_1209,In_1364);
or U4104 (N_4104,In_788,In_1045);
and U4105 (N_4105,In_1776,In_1074);
or U4106 (N_4106,In_1990,In_979);
nor U4107 (N_4107,In_1656,In_587);
nand U4108 (N_4108,In_1673,In_1757);
and U4109 (N_4109,In_1587,In_162);
nor U4110 (N_4110,In_1532,In_1033);
and U4111 (N_4111,In_1899,In_254);
and U4112 (N_4112,In_1091,In_474);
xnor U4113 (N_4113,In_1095,In_130);
and U4114 (N_4114,In_1377,In_1720);
or U4115 (N_4115,In_1301,In_342);
nor U4116 (N_4116,In_1547,In_101);
nand U4117 (N_4117,In_1556,In_1831);
and U4118 (N_4118,In_938,In_1131);
and U4119 (N_4119,In_1473,In_832);
or U4120 (N_4120,In_630,In_622);
nand U4121 (N_4121,In_1412,In_1788);
xnor U4122 (N_4122,In_1442,In_879);
nand U4123 (N_4123,In_1444,In_1598);
nand U4124 (N_4124,In_215,In_40);
and U4125 (N_4125,In_765,In_1136);
nand U4126 (N_4126,In_659,In_1162);
nor U4127 (N_4127,In_1763,In_1835);
nor U4128 (N_4128,In_823,In_350);
nor U4129 (N_4129,In_535,In_581);
nand U4130 (N_4130,In_606,In_216);
nand U4131 (N_4131,In_1968,In_1284);
or U4132 (N_4132,In_1178,In_1490);
xnor U4133 (N_4133,In_1461,In_740);
or U4134 (N_4134,In_988,In_1320);
and U4135 (N_4135,In_1740,In_1325);
xor U4136 (N_4136,In_429,In_318);
nand U4137 (N_4137,In_427,In_1720);
nand U4138 (N_4138,In_1042,In_635);
and U4139 (N_4139,In_1748,In_1228);
or U4140 (N_4140,In_1955,In_1246);
xnor U4141 (N_4141,In_218,In_1951);
or U4142 (N_4142,In_1609,In_1417);
xor U4143 (N_4143,In_1557,In_1600);
nand U4144 (N_4144,In_1436,In_350);
and U4145 (N_4145,In_1389,In_644);
nand U4146 (N_4146,In_263,In_1764);
or U4147 (N_4147,In_1505,In_281);
nor U4148 (N_4148,In_1345,In_1430);
and U4149 (N_4149,In_1124,In_515);
nand U4150 (N_4150,In_678,In_1749);
xor U4151 (N_4151,In_1028,In_444);
nand U4152 (N_4152,In_1064,In_1198);
or U4153 (N_4153,In_790,In_1626);
nand U4154 (N_4154,In_329,In_1951);
nor U4155 (N_4155,In_1142,In_929);
or U4156 (N_4156,In_1305,In_1346);
xor U4157 (N_4157,In_1416,In_1084);
xnor U4158 (N_4158,In_753,In_324);
xor U4159 (N_4159,In_867,In_385);
nand U4160 (N_4160,In_1134,In_417);
or U4161 (N_4161,In_1984,In_1902);
nand U4162 (N_4162,In_1388,In_543);
xor U4163 (N_4163,In_680,In_1439);
or U4164 (N_4164,In_1981,In_386);
xnor U4165 (N_4165,In_124,In_180);
xor U4166 (N_4166,In_382,In_1797);
nand U4167 (N_4167,In_1972,In_673);
xnor U4168 (N_4168,In_1377,In_1036);
nand U4169 (N_4169,In_832,In_1609);
or U4170 (N_4170,In_1602,In_659);
nand U4171 (N_4171,In_1519,In_1516);
nor U4172 (N_4172,In_389,In_1790);
xor U4173 (N_4173,In_1160,In_36);
nand U4174 (N_4174,In_1561,In_1952);
or U4175 (N_4175,In_1896,In_437);
xor U4176 (N_4176,In_238,In_789);
nor U4177 (N_4177,In_355,In_787);
nor U4178 (N_4178,In_766,In_507);
or U4179 (N_4179,In_515,In_767);
or U4180 (N_4180,In_1684,In_1482);
and U4181 (N_4181,In_1775,In_1332);
nor U4182 (N_4182,In_46,In_894);
nand U4183 (N_4183,In_547,In_1910);
xor U4184 (N_4184,In_416,In_785);
nand U4185 (N_4185,In_62,In_490);
or U4186 (N_4186,In_722,In_647);
or U4187 (N_4187,In_1239,In_605);
or U4188 (N_4188,In_1846,In_1355);
nor U4189 (N_4189,In_1504,In_247);
xor U4190 (N_4190,In_885,In_123);
nand U4191 (N_4191,In_1150,In_449);
and U4192 (N_4192,In_1591,In_1237);
nor U4193 (N_4193,In_1977,In_1099);
or U4194 (N_4194,In_563,In_1705);
and U4195 (N_4195,In_854,In_964);
xor U4196 (N_4196,In_220,In_1573);
xnor U4197 (N_4197,In_873,In_886);
or U4198 (N_4198,In_1152,In_1712);
xnor U4199 (N_4199,In_467,In_1148);
and U4200 (N_4200,In_954,In_141);
nor U4201 (N_4201,In_1808,In_1715);
or U4202 (N_4202,In_1474,In_1012);
nand U4203 (N_4203,In_140,In_189);
nand U4204 (N_4204,In_581,In_322);
and U4205 (N_4205,In_1539,In_1582);
nand U4206 (N_4206,In_340,In_1943);
nor U4207 (N_4207,In_964,In_1777);
and U4208 (N_4208,In_1310,In_1986);
nor U4209 (N_4209,In_1664,In_1235);
or U4210 (N_4210,In_1947,In_991);
xnor U4211 (N_4211,In_548,In_1381);
xor U4212 (N_4212,In_656,In_1617);
and U4213 (N_4213,In_1007,In_223);
or U4214 (N_4214,In_1590,In_35);
xor U4215 (N_4215,In_1381,In_581);
and U4216 (N_4216,In_54,In_1375);
nand U4217 (N_4217,In_410,In_869);
nor U4218 (N_4218,In_1897,In_1394);
and U4219 (N_4219,In_704,In_435);
nor U4220 (N_4220,In_948,In_1169);
and U4221 (N_4221,In_1254,In_1540);
nand U4222 (N_4222,In_805,In_1106);
or U4223 (N_4223,In_505,In_1915);
nand U4224 (N_4224,In_822,In_741);
nor U4225 (N_4225,In_1359,In_1819);
nand U4226 (N_4226,In_173,In_1972);
nand U4227 (N_4227,In_1679,In_1106);
nand U4228 (N_4228,In_584,In_750);
and U4229 (N_4229,In_566,In_1766);
nor U4230 (N_4230,In_1737,In_1460);
or U4231 (N_4231,In_782,In_234);
and U4232 (N_4232,In_1398,In_1372);
and U4233 (N_4233,In_1826,In_597);
and U4234 (N_4234,In_1523,In_1352);
and U4235 (N_4235,In_1658,In_935);
or U4236 (N_4236,In_1324,In_613);
and U4237 (N_4237,In_612,In_1264);
nor U4238 (N_4238,In_1659,In_424);
and U4239 (N_4239,In_253,In_1943);
or U4240 (N_4240,In_100,In_141);
and U4241 (N_4241,In_1360,In_1274);
nor U4242 (N_4242,In_914,In_1976);
and U4243 (N_4243,In_1288,In_877);
or U4244 (N_4244,In_1160,In_1219);
nor U4245 (N_4245,In_1924,In_1508);
and U4246 (N_4246,In_1977,In_804);
nor U4247 (N_4247,In_1943,In_1690);
or U4248 (N_4248,In_302,In_427);
or U4249 (N_4249,In_1512,In_1250);
or U4250 (N_4250,In_1405,In_113);
nor U4251 (N_4251,In_943,In_1373);
nor U4252 (N_4252,In_174,In_1425);
and U4253 (N_4253,In_1864,In_1252);
nor U4254 (N_4254,In_1579,In_1640);
or U4255 (N_4255,In_5,In_260);
nor U4256 (N_4256,In_1690,In_307);
xnor U4257 (N_4257,In_1462,In_1830);
xor U4258 (N_4258,In_322,In_916);
nor U4259 (N_4259,In_1547,In_860);
nand U4260 (N_4260,In_151,In_1103);
xor U4261 (N_4261,In_843,In_1918);
xor U4262 (N_4262,In_1078,In_1319);
or U4263 (N_4263,In_361,In_849);
nor U4264 (N_4264,In_796,In_24);
and U4265 (N_4265,In_1741,In_817);
and U4266 (N_4266,In_1482,In_823);
nand U4267 (N_4267,In_582,In_1693);
and U4268 (N_4268,In_1922,In_242);
nand U4269 (N_4269,In_1868,In_116);
nor U4270 (N_4270,In_235,In_1125);
nand U4271 (N_4271,In_588,In_1122);
xnor U4272 (N_4272,In_627,In_296);
xor U4273 (N_4273,In_436,In_1730);
nor U4274 (N_4274,In_985,In_110);
or U4275 (N_4275,In_1698,In_299);
or U4276 (N_4276,In_1345,In_1582);
and U4277 (N_4277,In_966,In_1477);
xor U4278 (N_4278,In_1743,In_886);
nor U4279 (N_4279,In_1801,In_78);
xnor U4280 (N_4280,In_1319,In_328);
nor U4281 (N_4281,In_1091,In_1202);
xnor U4282 (N_4282,In_292,In_907);
or U4283 (N_4283,In_123,In_29);
nand U4284 (N_4284,In_1946,In_256);
nor U4285 (N_4285,In_1592,In_238);
xor U4286 (N_4286,In_815,In_46);
xnor U4287 (N_4287,In_372,In_1421);
xor U4288 (N_4288,In_1601,In_1767);
xnor U4289 (N_4289,In_295,In_1045);
nor U4290 (N_4290,In_1759,In_1305);
and U4291 (N_4291,In_1042,In_1867);
xor U4292 (N_4292,In_1169,In_942);
or U4293 (N_4293,In_430,In_1825);
xor U4294 (N_4294,In_800,In_1392);
nand U4295 (N_4295,In_1241,In_1965);
and U4296 (N_4296,In_1131,In_1636);
or U4297 (N_4297,In_689,In_1782);
or U4298 (N_4298,In_455,In_896);
xor U4299 (N_4299,In_1856,In_1965);
xor U4300 (N_4300,In_743,In_346);
or U4301 (N_4301,In_564,In_480);
nor U4302 (N_4302,In_1437,In_627);
and U4303 (N_4303,In_1630,In_1531);
nor U4304 (N_4304,In_757,In_682);
nor U4305 (N_4305,In_1881,In_1374);
xor U4306 (N_4306,In_1446,In_1749);
or U4307 (N_4307,In_1940,In_342);
nor U4308 (N_4308,In_621,In_1918);
or U4309 (N_4309,In_694,In_1563);
nand U4310 (N_4310,In_98,In_1728);
and U4311 (N_4311,In_446,In_1583);
nor U4312 (N_4312,In_1934,In_920);
nor U4313 (N_4313,In_555,In_707);
and U4314 (N_4314,In_62,In_599);
nor U4315 (N_4315,In_534,In_235);
nor U4316 (N_4316,In_1975,In_778);
nand U4317 (N_4317,In_296,In_1528);
xor U4318 (N_4318,In_1280,In_862);
nand U4319 (N_4319,In_377,In_1110);
nand U4320 (N_4320,In_593,In_1068);
xnor U4321 (N_4321,In_1061,In_1066);
and U4322 (N_4322,In_1277,In_649);
nor U4323 (N_4323,In_1318,In_784);
nor U4324 (N_4324,In_826,In_994);
and U4325 (N_4325,In_31,In_1422);
nor U4326 (N_4326,In_1532,In_719);
nor U4327 (N_4327,In_983,In_1490);
and U4328 (N_4328,In_1954,In_303);
and U4329 (N_4329,In_44,In_1248);
nand U4330 (N_4330,In_1254,In_1636);
and U4331 (N_4331,In_1775,In_545);
nor U4332 (N_4332,In_282,In_1548);
nand U4333 (N_4333,In_1305,In_1270);
nor U4334 (N_4334,In_28,In_1071);
and U4335 (N_4335,In_1275,In_1879);
and U4336 (N_4336,In_43,In_746);
nand U4337 (N_4337,In_194,In_46);
xnor U4338 (N_4338,In_424,In_1917);
xor U4339 (N_4339,In_236,In_1217);
xnor U4340 (N_4340,In_1990,In_364);
and U4341 (N_4341,In_1203,In_1023);
or U4342 (N_4342,In_17,In_1892);
nand U4343 (N_4343,In_1476,In_407);
xnor U4344 (N_4344,In_752,In_1791);
or U4345 (N_4345,In_1951,In_1117);
nor U4346 (N_4346,In_120,In_1495);
nand U4347 (N_4347,In_959,In_1402);
xor U4348 (N_4348,In_823,In_410);
xor U4349 (N_4349,In_1031,In_889);
nor U4350 (N_4350,In_124,In_1003);
xor U4351 (N_4351,In_1608,In_1552);
nand U4352 (N_4352,In_1208,In_70);
or U4353 (N_4353,In_780,In_1909);
xnor U4354 (N_4354,In_1652,In_705);
or U4355 (N_4355,In_149,In_1662);
and U4356 (N_4356,In_860,In_1976);
or U4357 (N_4357,In_1942,In_1051);
xor U4358 (N_4358,In_47,In_620);
and U4359 (N_4359,In_1729,In_285);
or U4360 (N_4360,In_370,In_770);
nand U4361 (N_4361,In_922,In_1839);
and U4362 (N_4362,In_862,In_863);
nor U4363 (N_4363,In_357,In_708);
and U4364 (N_4364,In_733,In_787);
or U4365 (N_4365,In_626,In_1958);
or U4366 (N_4366,In_444,In_127);
and U4367 (N_4367,In_34,In_252);
xnor U4368 (N_4368,In_243,In_1566);
nand U4369 (N_4369,In_1990,In_1980);
or U4370 (N_4370,In_258,In_642);
nand U4371 (N_4371,In_1338,In_1664);
xor U4372 (N_4372,In_1761,In_1602);
nor U4373 (N_4373,In_175,In_1873);
or U4374 (N_4374,In_613,In_1248);
or U4375 (N_4375,In_587,In_1051);
or U4376 (N_4376,In_95,In_958);
xor U4377 (N_4377,In_1076,In_1545);
nor U4378 (N_4378,In_1170,In_15);
xor U4379 (N_4379,In_1221,In_974);
nand U4380 (N_4380,In_372,In_580);
nand U4381 (N_4381,In_494,In_899);
xnor U4382 (N_4382,In_1710,In_956);
nor U4383 (N_4383,In_71,In_1573);
nand U4384 (N_4384,In_738,In_1977);
nor U4385 (N_4385,In_331,In_978);
nor U4386 (N_4386,In_1700,In_1436);
nand U4387 (N_4387,In_1419,In_924);
or U4388 (N_4388,In_745,In_1918);
or U4389 (N_4389,In_661,In_363);
xnor U4390 (N_4390,In_1988,In_506);
and U4391 (N_4391,In_666,In_1893);
nor U4392 (N_4392,In_528,In_1708);
and U4393 (N_4393,In_687,In_1474);
nand U4394 (N_4394,In_44,In_433);
and U4395 (N_4395,In_693,In_964);
and U4396 (N_4396,In_410,In_982);
and U4397 (N_4397,In_1966,In_1644);
and U4398 (N_4398,In_1809,In_593);
xnor U4399 (N_4399,In_924,In_1447);
nand U4400 (N_4400,In_267,In_57);
and U4401 (N_4401,In_1997,In_1651);
nor U4402 (N_4402,In_1218,In_678);
xnor U4403 (N_4403,In_476,In_276);
nand U4404 (N_4404,In_544,In_1063);
or U4405 (N_4405,In_1917,In_1070);
or U4406 (N_4406,In_438,In_426);
nand U4407 (N_4407,In_1444,In_834);
nand U4408 (N_4408,In_899,In_161);
and U4409 (N_4409,In_1277,In_916);
xor U4410 (N_4410,In_876,In_1759);
and U4411 (N_4411,In_651,In_1468);
nor U4412 (N_4412,In_1908,In_1589);
nand U4413 (N_4413,In_1075,In_828);
nand U4414 (N_4414,In_600,In_1537);
and U4415 (N_4415,In_66,In_428);
or U4416 (N_4416,In_1379,In_478);
nor U4417 (N_4417,In_854,In_803);
or U4418 (N_4418,In_1310,In_309);
and U4419 (N_4419,In_891,In_990);
xor U4420 (N_4420,In_1282,In_522);
and U4421 (N_4421,In_1719,In_126);
nor U4422 (N_4422,In_1574,In_760);
or U4423 (N_4423,In_1716,In_1871);
xnor U4424 (N_4424,In_276,In_366);
nand U4425 (N_4425,In_511,In_933);
or U4426 (N_4426,In_208,In_605);
and U4427 (N_4427,In_758,In_1025);
and U4428 (N_4428,In_808,In_1437);
and U4429 (N_4429,In_1772,In_567);
nand U4430 (N_4430,In_1308,In_1554);
xnor U4431 (N_4431,In_596,In_1194);
nand U4432 (N_4432,In_198,In_598);
or U4433 (N_4433,In_1012,In_28);
and U4434 (N_4434,In_1432,In_1474);
nand U4435 (N_4435,In_1734,In_1211);
xor U4436 (N_4436,In_147,In_29);
and U4437 (N_4437,In_1145,In_1986);
and U4438 (N_4438,In_1669,In_1897);
xor U4439 (N_4439,In_1267,In_554);
xor U4440 (N_4440,In_133,In_190);
nand U4441 (N_4441,In_1963,In_64);
and U4442 (N_4442,In_394,In_1174);
or U4443 (N_4443,In_1086,In_1118);
nand U4444 (N_4444,In_1871,In_763);
and U4445 (N_4445,In_338,In_1011);
nor U4446 (N_4446,In_630,In_309);
nand U4447 (N_4447,In_44,In_1411);
xor U4448 (N_4448,In_1414,In_1072);
or U4449 (N_4449,In_6,In_1010);
and U4450 (N_4450,In_1068,In_1462);
or U4451 (N_4451,In_13,In_531);
nand U4452 (N_4452,In_1289,In_1233);
or U4453 (N_4453,In_995,In_480);
nor U4454 (N_4454,In_295,In_283);
nor U4455 (N_4455,In_1166,In_1061);
nor U4456 (N_4456,In_635,In_1337);
nand U4457 (N_4457,In_650,In_386);
xor U4458 (N_4458,In_1606,In_678);
nor U4459 (N_4459,In_730,In_1498);
nand U4460 (N_4460,In_1945,In_1529);
or U4461 (N_4461,In_1714,In_1731);
nand U4462 (N_4462,In_1698,In_1388);
xor U4463 (N_4463,In_1555,In_1866);
nor U4464 (N_4464,In_1826,In_1718);
nand U4465 (N_4465,In_1846,In_383);
or U4466 (N_4466,In_1034,In_1224);
and U4467 (N_4467,In_1387,In_1320);
nor U4468 (N_4468,In_1355,In_778);
nor U4469 (N_4469,In_1024,In_1681);
xor U4470 (N_4470,In_741,In_811);
nand U4471 (N_4471,In_1148,In_466);
or U4472 (N_4472,In_1369,In_1327);
or U4473 (N_4473,In_569,In_1285);
xnor U4474 (N_4474,In_1390,In_975);
or U4475 (N_4475,In_1729,In_1400);
or U4476 (N_4476,In_460,In_1889);
nand U4477 (N_4477,In_1848,In_1948);
nand U4478 (N_4478,In_1491,In_1724);
and U4479 (N_4479,In_1571,In_1279);
and U4480 (N_4480,In_1287,In_1723);
and U4481 (N_4481,In_1042,In_523);
nor U4482 (N_4482,In_726,In_1928);
or U4483 (N_4483,In_1112,In_1352);
and U4484 (N_4484,In_1011,In_534);
xnor U4485 (N_4485,In_1048,In_404);
nand U4486 (N_4486,In_193,In_615);
nor U4487 (N_4487,In_856,In_178);
xor U4488 (N_4488,In_906,In_454);
nor U4489 (N_4489,In_267,In_835);
or U4490 (N_4490,In_1570,In_1745);
nor U4491 (N_4491,In_1615,In_271);
nor U4492 (N_4492,In_469,In_940);
nor U4493 (N_4493,In_639,In_275);
nand U4494 (N_4494,In_1685,In_1521);
or U4495 (N_4495,In_909,In_616);
and U4496 (N_4496,In_346,In_1774);
or U4497 (N_4497,In_1149,In_195);
nand U4498 (N_4498,In_548,In_54);
and U4499 (N_4499,In_764,In_1179);
xor U4500 (N_4500,In_599,In_1903);
nor U4501 (N_4501,In_1743,In_1027);
xor U4502 (N_4502,In_1361,In_1151);
xor U4503 (N_4503,In_592,In_647);
and U4504 (N_4504,In_1385,In_222);
nand U4505 (N_4505,In_299,In_1308);
nor U4506 (N_4506,In_120,In_688);
or U4507 (N_4507,In_64,In_1886);
xnor U4508 (N_4508,In_1996,In_90);
and U4509 (N_4509,In_1540,In_1409);
and U4510 (N_4510,In_1348,In_341);
or U4511 (N_4511,In_1388,In_1675);
nor U4512 (N_4512,In_1684,In_1068);
or U4513 (N_4513,In_281,In_439);
nand U4514 (N_4514,In_1320,In_673);
or U4515 (N_4515,In_851,In_622);
or U4516 (N_4516,In_959,In_51);
nor U4517 (N_4517,In_1143,In_107);
nor U4518 (N_4518,In_1338,In_206);
xnor U4519 (N_4519,In_930,In_1295);
or U4520 (N_4520,In_805,In_1929);
nand U4521 (N_4521,In_912,In_428);
nor U4522 (N_4522,In_432,In_1580);
nor U4523 (N_4523,In_379,In_310);
nor U4524 (N_4524,In_1645,In_182);
or U4525 (N_4525,In_1205,In_264);
nor U4526 (N_4526,In_1204,In_1205);
nand U4527 (N_4527,In_270,In_1209);
nand U4528 (N_4528,In_1982,In_509);
xor U4529 (N_4529,In_1765,In_1163);
nor U4530 (N_4530,In_1759,In_549);
and U4531 (N_4531,In_1524,In_716);
nand U4532 (N_4532,In_1173,In_1111);
nor U4533 (N_4533,In_1164,In_1807);
nand U4534 (N_4534,In_907,In_1961);
xor U4535 (N_4535,In_1890,In_174);
or U4536 (N_4536,In_1502,In_1660);
and U4537 (N_4537,In_1579,In_1854);
or U4538 (N_4538,In_479,In_54);
nor U4539 (N_4539,In_1659,In_743);
nor U4540 (N_4540,In_1196,In_858);
xor U4541 (N_4541,In_1977,In_1774);
nor U4542 (N_4542,In_1438,In_26);
nand U4543 (N_4543,In_1909,In_1977);
nor U4544 (N_4544,In_930,In_418);
nand U4545 (N_4545,In_1088,In_447);
xor U4546 (N_4546,In_1682,In_64);
nand U4547 (N_4547,In_1622,In_1879);
nor U4548 (N_4548,In_1415,In_1605);
nand U4549 (N_4549,In_486,In_809);
xor U4550 (N_4550,In_1926,In_1247);
nor U4551 (N_4551,In_66,In_1945);
or U4552 (N_4552,In_1990,In_297);
nand U4553 (N_4553,In_1209,In_61);
and U4554 (N_4554,In_1526,In_1833);
xor U4555 (N_4555,In_1152,In_1762);
nand U4556 (N_4556,In_1847,In_626);
nand U4557 (N_4557,In_1838,In_1529);
nor U4558 (N_4558,In_1473,In_1677);
xor U4559 (N_4559,In_1665,In_1633);
xor U4560 (N_4560,In_1413,In_420);
nor U4561 (N_4561,In_217,In_140);
nand U4562 (N_4562,In_1918,In_1438);
xor U4563 (N_4563,In_839,In_1339);
and U4564 (N_4564,In_1736,In_517);
or U4565 (N_4565,In_1502,In_398);
and U4566 (N_4566,In_1747,In_1508);
nand U4567 (N_4567,In_415,In_1090);
or U4568 (N_4568,In_1009,In_27);
nand U4569 (N_4569,In_969,In_1633);
and U4570 (N_4570,In_1257,In_1000);
xnor U4571 (N_4571,In_359,In_1817);
and U4572 (N_4572,In_1582,In_665);
and U4573 (N_4573,In_1506,In_873);
or U4574 (N_4574,In_984,In_1912);
nand U4575 (N_4575,In_1241,In_1769);
and U4576 (N_4576,In_1252,In_850);
or U4577 (N_4577,In_1500,In_379);
and U4578 (N_4578,In_658,In_1666);
xor U4579 (N_4579,In_947,In_1838);
and U4580 (N_4580,In_1849,In_1153);
or U4581 (N_4581,In_1921,In_461);
nand U4582 (N_4582,In_1071,In_191);
nor U4583 (N_4583,In_883,In_1686);
or U4584 (N_4584,In_480,In_1114);
and U4585 (N_4585,In_568,In_46);
xor U4586 (N_4586,In_583,In_1416);
nand U4587 (N_4587,In_407,In_154);
nand U4588 (N_4588,In_584,In_330);
xnor U4589 (N_4589,In_578,In_1448);
nand U4590 (N_4590,In_307,In_835);
and U4591 (N_4591,In_1286,In_1620);
xnor U4592 (N_4592,In_588,In_1591);
and U4593 (N_4593,In_1739,In_1907);
nand U4594 (N_4594,In_385,In_980);
or U4595 (N_4595,In_1399,In_1736);
nor U4596 (N_4596,In_1976,In_1870);
nand U4597 (N_4597,In_1656,In_223);
and U4598 (N_4598,In_91,In_219);
xor U4599 (N_4599,In_1624,In_1211);
nor U4600 (N_4600,In_1001,In_1660);
nand U4601 (N_4601,In_648,In_383);
and U4602 (N_4602,In_1615,In_1774);
nor U4603 (N_4603,In_1579,In_109);
nand U4604 (N_4604,In_1299,In_913);
xor U4605 (N_4605,In_1425,In_1917);
nor U4606 (N_4606,In_688,In_161);
and U4607 (N_4607,In_367,In_76);
and U4608 (N_4608,In_803,In_670);
nand U4609 (N_4609,In_445,In_550);
nor U4610 (N_4610,In_939,In_1971);
or U4611 (N_4611,In_956,In_626);
nor U4612 (N_4612,In_351,In_855);
or U4613 (N_4613,In_132,In_1739);
or U4614 (N_4614,In_1990,In_1743);
nor U4615 (N_4615,In_1997,In_501);
xnor U4616 (N_4616,In_76,In_1377);
or U4617 (N_4617,In_1339,In_503);
and U4618 (N_4618,In_1755,In_1886);
and U4619 (N_4619,In_162,In_828);
xor U4620 (N_4620,In_1971,In_1632);
or U4621 (N_4621,In_199,In_1372);
and U4622 (N_4622,In_1024,In_1244);
nor U4623 (N_4623,In_1676,In_1767);
or U4624 (N_4624,In_1688,In_1858);
and U4625 (N_4625,In_227,In_0);
nor U4626 (N_4626,In_1990,In_1703);
nor U4627 (N_4627,In_722,In_540);
nor U4628 (N_4628,In_540,In_1014);
nand U4629 (N_4629,In_1096,In_788);
nand U4630 (N_4630,In_1012,In_689);
xor U4631 (N_4631,In_1923,In_798);
xnor U4632 (N_4632,In_1954,In_1561);
xnor U4633 (N_4633,In_403,In_1998);
xor U4634 (N_4634,In_307,In_1333);
nor U4635 (N_4635,In_1413,In_1370);
and U4636 (N_4636,In_1057,In_465);
or U4637 (N_4637,In_1424,In_427);
or U4638 (N_4638,In_408,In_278);
and U4639 (N_4639,In_764,In_1782);
nand U4640 (N_4640,In_754,In_988);
nand U4641 (N_4641,In_1065,In_7);
nor U4642 (N_4642,In_1374,In_1131);
nor U4643 (N_4643,In_1596,In_200);
nor U4644 (N_4644,In_103,In_941);
nand U4645 (N_4645,In_415,In_1600);
nand U4646 (N_4646,In_189,In_228);
nand U4647 (N_4647,In_675,In_1708);
and U4648 (N_4648,In_102,In_52);
and U4649 (N_4649,In_1329,In_1042);
xnor U4650 (N_4650,In_1028,In_871);
nand U4651 (N_4651,In_995,In_0);
nor U4652 (N_4652,In_279,In_1289);
xor U4653 (N_4653,In_515,In_1965);
nor U4654 (N_4654,In_861,In_465);
and U4655 (N_4655,In_1365,In_1846);
nor U4656 (N_4656,In_1190,In_1128);
or U4657 (N_4657,In_1120,In_1178);
nand U4658 (N_4658,In_869,In_1833);
xnor U4659 (N_4659,In_1197,In_814);
xnor U4660 (N_4660,In_1626,In_589);
and U4661 (N_4661,In_782,In_721);
nor U4662 (N_4662,In_1239,In_1425);
nand U4663 (N_4663,In_1640,In_1831);
xor U4664 (N_4664,In_1603,In_824);
nor U4665 (N_4665,In_998,In_1721);
xor U4666 (N_4666,In_1953,In_452);
or U4667 (N_4667,In_945,In_45);
and U4668 (N_4668,In_563,In_706);
xor U4669 (N_4669,In_1999,In_1536);
xnor U4670 (N_4670,In_1238,In_235);
nand U4671 (N_4671,In_298,In_77);
nor U4672 (N_4672,In_871,In_1677);
and U4673 (N_4673,In_221,In_522);
nand U4674 (N_4674,In_1464,In_1159);
nor U4675 (N_4675,In_1278,In_993);
or U4676 (N_4676,In_1046,In_934);
or U4677 (N_4677,In_377,In_971);
and U4678 (N_4678,In_1753,In_1627);
nand U4679 (N_4679,In_209,In_205);
nand U4680 (N_4680,In_1242,In_787);
xnor U4681 (N_4681,In_1900,In_616);
or U4682 (N_4682,In_1437,In_1434);
or U4683 (N_4683,In_448,In_88);
or U4684 (N_4684,In_395,In_1201);
or U4685 (N_4685,In_1168,In_1735);
nand U4686 (N_4686,In_1176,In_90);
or U4687 (N_4687,In_1643,In_1918);
or U4688 (N_4688,In_573,In_1021);
nor U4689 (N_4689,In_652,In_569);
xor U4690 (N_4690,In_1991,In_1344);
or U4691 (N_4691,In_763,In_668);
xor U4692 (N_4692,In_39,In_143);
and U4693 (N_4693,In_1462,In_1420);
xor U4694 (N_4694,In_1067,In_469);
and U4695 (N_4695,In_568,In_318);
nor U4696 (N_4696,In_1866,In_309);
nor U4697 (N_4697,In_1910,In_174);
or U4698 (N_4698,In_1380,In_1397);
and U4699 (N_4699,In_44,In_315);
nand U4700 (N_4700,In_1913,In_757);
or U4701 (N_4701,In_636,In_855);
or U4702 (N_4702,In_158,In_387);
nor U4703 (N_4703,In_1838,In_1232);
nor U4704 (N_4704,In_197,In_1370);
nor U4705 (N_4705,In_415,In_1543);
xnor U4706 (N_4706,In_1783,In_1534);
nor U4707 (N_4707,In_227,In_1638);
and U4708 (N_4708,In_418,In_510);
nor U4709 (N_4709,In_1861,In_345);
or U4710 (N_4710,In_1968,In_649);
xor U4711 (N_4711,In_1910,In_149);
nor U4712 (N_4712,In_1175,In_802);
xnor U4713 (N_4713,In_1147,In_699);
nor U4714 (N_4714,In_1979,In_1594);
nand U4715 (N_4715,In_1107,In_1909);
and U4716 (N_4716,In_1334,In_421);
nor U4717 (N_4717,In_1339,In_266);
or U4718 (N_4718,In_454,In_519);
xnor U4719 (N_4719,In_520,In_1601);
xnor U4720 (N_4720,In_1302,In_402);
nand U4721 (N_4721,In_788,In_1031);
nor U4722 (N_4722,In_887,In_1882);
nor U4723 (N_4723,In_485,In_1150);
xor U4724 (N_4724,In_1688,In_1783);
xnor U4725 (N_4725,In_1380,In_1874);
or U4726 (N_4726,In_1054,In_842);
and U4727 (N_4727,In_1978,In_1050);
xnor U4728 (N_4728,In_1806,In_1681);
or U4729 (N_4729,In_1661,In_634);
and U4730 (N_4730,In_250,In_1316);
or U4731 (N_4731,In_864,In_239);
or U4732 (N_4732,In_711,In_1383);
nand U4733 (N_4733,In_767,In_623);
nand U4734 (N_4734,In_623,In_1875);
and U4735 (N_4735,In_556,In_242);
nand U4736 (N_4736,In_1380,In_881);
nor U4737 (N_4737,In_1255,In_719);
or U4738 (N_4738,In_817,In_213);
or U4739 (N_4739,In_165,In_127);
and U4740 (N_4740,In_1314,In_1668);
xnor U4741 (N_4741,In_1485,In_1656);
or U4742 (N_4742,In_1243,In_214);
nand U4743 (N_4743,In_1459,In_1133);
or U4744 (N_4744,In_1022,In_999);
or U4745 (N_4745,In_1196,In_644);
or U4746 (N_4746,In_468,In_938);
nor U4747 (N_4747,In_1917,In_389);
nand U4748 (N_4748,In_1868,In_1934);
nand U4749 (N_4749,In_885,In_603);
nand U4750 (N_4750,In_1387,In_1554);
or U4751 (N_4751,In_1282,In_309);
and U4752 (N_4752,In_1690,In_1616);
or U4753 (N_4753,In_1880,In_1200);
xnor U4754 (N_4754,In_1073,In_1933);
xnor U4755 (N_4755,In_1974,In_174);
nand U4756 (N_4756,In_759,In_895);
or U4757 (N_4757,In_388,In_1051);
or U4758 (N_4758,In_1030,In_1747);
and U4759 (N_4759,In_1973,In_162);
nand U4760 (N_4760,In_1597,In_889);
nor U4761 (N_4761,In_506,In_156);
xor U4762 (N_4762,In_106,In_1464);
nor U4763 (N_4763,In_696,In_920);
nand U4764 (N_4764,In_1730,In_1986);
nand U4765 (N_4765,In_40,In_1663);
and U4766 (N_4766,In_1247,In_393);
and U4767 (N_4767,In_544,In_1051);
nand U4768 (N_4768,In_506,In_886);
and U4769 (N_4769,In_1745,In_1614);
xor U4770 (N_4770,In_725,In_1864);
nand U4771 (N_4771,In_569,In_255);
xnor U4772 (N_4772,In_767,In_87);
and U4773 (N_4773,In_1183,In_294);
or U4774 (N_4774,In_1410,In_1025);
xnor U4775 (N_4775,In_492,In_96);
or U4776 (N_4776,In_1696,In_193);
or U4777 (N_4777,In_935,In_1288);
nor U4778 (N_4778,In_1775,In_1281);
nand U4779 (N_4779,In_1442,In_696);
nand U4780 (N_4780,In_1485,In_1228);
and U4781 (N_4781,In_1287,In_1974);
and U4782 (N_4782,In_94,In_1155);
nor U4783 (N_4783,In_958,In_822);
nor U4784 (N_4784,In_730,In_1131);
or U4785 (N_4785,In_1066,In_344);
xor U4786 (N_4786,In_1130,In_174);
nor U4787 (N_4787,In_905,In_1573);
xnor U4788 (N_4788,In_930,In_507);
and U4789 (N_4789,In_1417,In_1519);
xnor U4790 (N_4790,In_1330,In_414);
xor U4791 (N_4791,In_43,In_1844);
and U4792 (N_4792,In_1638,In_750);
or U4793 (N_4793,In_1649,In_1696);
xnor U4794 (N_4794,In_1214,In_1416);
nand U4795 (N_4795,In_299,In_138);
and U4796 (N_4796,In_1651,In_250);
nand U4797 (N_4797,In_83,In_44);
nor U4798 (N_4798,In_1270,In_1138);
xor U4799 (N_4799,In_795,In_1759);
nand U4800 (N_4800,In_1505,In_1006);
xnor U4801 (N_4801,In_752,In_351);
xor U4802 (N_4802,In_591,In_1512);
or U4803 (N_4803,In_1623,In_1476);
nor U4804 (N_4804,In_508,In_1787);
and U4805 (N_4805,In_1032,In_1289);
xnor U4806 (N_4806,In_541,In_1154);
nor U4807 (N_4807,In_1841,In_673);
xor U4808 (N_4808,In_204,In_377);
nand U4809 (N_4809,In_1830,In_671);
xor U4810 (N_4810,In_1593,In_213);
or U4811 (N_4811,In_1987,In_289);
nand U4812 (N_4812,In_220,In_1130);
nor U4813 (N_4813,In_809,In_1011);
and U4814 (N_4814,In_1103,In_545);
nor U4815 (N_4815,In_1143,In_1887);
or U4816 (N_4816,In_1301,In_820);
or U4817 (N_4817,In_1643,In_638);
or U4818 (N_4818,In_313,In_362);
and U4819 (N_4819,In_1045,In_1057);
or U4820 (N_4820,In_383,In_169);
nor U4821 (N_4821,In_950,In_1904);
xnor U4822 (N_4822,In_155,In_1576);
nand U4823 (N_4823,In_1856,In_209);
and U4824 (N_4824,In_1218,In_127);
nand U4825 (N_4825,In_1507,In_1105);
or U4826 (N_4826,In_1915,In_479);
or U4827 (N_4827,In_1213,In_1664);
or U4828 (N_4828,In_1315,In_1351);
xor U4829 (N_4829,In_923,In_1414);
nand U4830 (N_4830,In_1989,In_154);
nand U4831 (N_4831,In_953,In_487);
nor U4832 (N_4832,In_1290,In_553);
nor U4833 (N_4833,In_746,In_464);
nor U4834 (N_4834,In_1098,In_27);
nand U4835 (N_4835,In_1968,In_516);
nor U4836 (N_4836,In_708,In_359);
nand U4837 (N_4837,In_127,In_26);
nor U4838 (N_4838,In_1574,In_98);
or U4839 (N_4839,In_1551,In_1988);
and U4840 (N_4840,In_526,In_291);
nand U4841 (N_4841,In_317,In_344);
nand U4842 (N_4842,In_197,In_1398);
or U4843 (N_4843,In_1033,In_1741);
or U4844 (N_4844,In_1770,In_720);
xnor U4845 (N_4845,In_263,In_1742);
nand U4846 (N_4846,In_899,In_1060);
and U4847 (N_4847,In_625,In_761);
and U4848 (N_4848,In_1641,In_1662);
nor U4849 (N_4849,In_681,In_687);
or U4850 (N_4850,In_1553,In_677);
xor U4851 (N_4851,In_474,In_85);
nor U4852 (N_4852,In_218,In_1870);
nor U4853 (N_4853,In_1240,In_1738);
xnor U4854 (N_4854,In_706,In_1312);
and U4855 (N_4855,In_428,In_725);
and U4856 (N_4856,In_29,In_1775);
nor U4857 (N_4857,In_1125,In_1441);
xor U4858 (N_4858,In_1018,In_1291);
xor U4859 (N_4859,In_1566,In_1269);
nor U4860 (N_4860,In_1123,In_1025);
and U4861 (N_4861,In_1591,In_1376);
xnor U4862 (N_4862,In_357,In_1198);
and U4863 (N_4863,In_1842,In_1635);
or U4864 (N_4864,In_581,In_1747);
xor U4865 (N_4865,In_121,In_1185);
nor U4866 (N_4866,In_1405,In_1993);
and U4867 (N_4867,In_1946,In_1822);
nand U4868 (N_4868,In_421,In_1131);
nor U4869 (N_4869,In_267,In_76);
or U4870 (N_4870,In_1245,In_854);
and U4871 (N_4871,In_1078,In_244);
nand U4872 (N_4872,In_1512,In_1176);
nor U4873 (N_4873,In_893,In_1561);
and U4874 (N_4874,In_733,In_1245);
nand U4875 (N_4875,In_1366,In_90);
xnor U4876 (N_4876,In_209,In_1488);
nor U4877 (N_4877,In_1756,In_261);
and U4878 (N_4878,In_1165,In_937);
and U4879 (N_4879,In_1142,In_265);
xnor U4880 (N_4880,In_917,In_921);
nand U4881 (N_4881,In_1897,In_1636);
nand U4882 (N_4882,In_1803,In_1373);
nand U4883 (N_4883,In_343,In_1114);
nand U4884 (N_4884,In_1146,In_1738);
or U4885 (N_4885,In_1603,In_1136);
nand U4886 (N_4886,In_123,In_368);
nand U4887 (N_4887,In_1477,In_1468);
and U4888 (N_4888,In_685,In_180);
and U4889 (N_4889,In_890,In_1934);
nand U4890 (N_4890,In_538,In_713);
nand U4891 (N_4891,In_909,In_1174);
nor U4892 (N_4892,In_747,In_538);
or U4893 (N_4893,In_1169,In_941);
and U4894 (N_4894,In_725,In_1781);
nand U4895 (N_4895,In_1570,In_972);
and U4896 (N_4896,In_262,In_1656);
or U4897 (N_4897,In_497,In_780);
xor U4898 (N_4898,In_456,In_1329);
xnor U4899 (N_4899,In_608,In_1966);
and U4900 (N_4900,In_1994,In_9);
nor U4901 (N_4901,In_1489,In_991);
xor U4902 (N_4902,In_1244,In_342);
and U4903 (N_4903,In_1164,In_512);
xnor U4904 (N_4904,In_653,In_1741);
xnor U4905 (N_4905,In_1448,In_1950);
xor U4906 (N_4906,In_622,In_1924);
nor U4907 (N_4907,In_890,In_1665);
nor U4908 (N_4908,In_184,In_157);
or U4909 (N_4909,In_831,In_55);
xnor U4910 (N_4910,In_1815,In_657);
xnor U4911 (N_4911,In_1156,In_533);
or U4912 (N_4912,In_360,In_1865);
nor U4913 (N_4913,In_793,In_1705);
nand U4914 (N_4914,In_936,In_1386);
or U4915 (N_4915,In_1321,In_1348);
xor U4916 (N_4916,In_198,In_451);
nor U4917 (N_4917,In_1662,In_179);
nor U4918 (N_4918,In_1363,In_274);
nor U4919 (N_4919,In_1177,In_684);
xor U4920 (N_4920,In_1723,In_1887);
or U4921 (N_4921,In_883,In_1182);
nor U4922 (N_4922,In_309,In_1069);
nor U4923 (N_4923,In_1851,In_924);
or U4924 (N_4924,In_1256,In_1857);
or U4925 (N_4925,In_1411,In_397);
nand U4926 (N_4926,In_1561,In_1960);
and U4927 (N_4927,In_869,In_1109);
or U4928 (N_4928,In_78,In_1970);
xor U4929 (N_4929,In_1576,In_481);
and U4930 (N_4930,In_1828,In_1056);
or U4931 (N_4931,In_1107,In_306);
and U4932 (N_4932,In_1739,In_376);
nor U4933 (N_4933,In_574,In_113);
or U4934 (N_4934,In_34,In_735);
nor U4935 (N_4935,In_13,In_523);
or U4936 (N_4936,In_46,In_39);
and U4937 (N_4937,In_1195,In_1696);
nor U4938 (N_4938,In_1997,In_1917);
nor U4939 (N_4939,In_1896,In_379);
or U4940 (N_4940,In_1249,In_894);
or U4941 (N_4941,In_704,In_1633);
nor U4942 (N_4942,In_827,In_1415);
nand U4943 (N_4943,In_560,In_1717);
xor U4944 (N_4944,In_1782,In_1057);
and U4945 (N_4945,In_1897,In_1785);
nor U4946 (N_4946,In_1270,In_1386);
and U4947 (N_4947,In_1532,In_1294);
nand U4948 (N_4948,In_1730,In_1015);
or U4949 (N_4949,In_1441,In_72);
nor U4950 (N_4950,In_1635,In_832);
or U4951 (N_4951,In_1488,In_776);
or U4952 (N_4952,In_1727,In_1753);
nand U4953 (N_4953,In_1065,In_1981);
xor U4954 (N_4954,In_37,In_1751);
or U4955 (N_4955,In_46,In_204);
xnor U4956 (N_4956,In_1558,In_1373);
and U4957 (N_4957,In_95,In_677);
xnor U4958 (N_4958,In_1984,In_744);
or U4959 (N_4959,In_244,In_1211);
or U4960 (N_4960,In_705,In_292);
or U4961 (N_4961,In_658,In_1865);
or U4962 (N_4962,In_1513,In_491);
nand U4963 (N_4963,In_1430,In_1474);
nand U4964 (N_4964,In_1805,In_198);
nand U4965 (N_4965,In_1726,In_1233);
or U4966 (N_4966,In_293,In_441);
and U4967 (N_4967,In_1742,In_367);
nand U4968 (N_4968,In_1888,In_730);
nor U4969 (N_4969,In_308,In_1705);
nand U4970 (N_4970,In_988,In_77);
xor U4971 (N_4971,In_1524,In_308);
nand U4972 (N_4972,In_1965,In_1780);
or U4973 (N_4973,In_1607,In_324);
nand U4974 (N_4974,In_1074,In_1099);
xor U4975 (N_4975,In_589,In_556);
xnor U4976 (N_4976,In_138,In_12);
or U4977 (N_4977,In_1112,In_328);
nor U4978 (N_4978,In_1340,In_1296);
xor U4979 (N_4979,In_709,In_702);
nor U4980 (N_4980,In_1439,In_1798);
xnor U4981 (N_4981,In_179,In_840);
or U4982 (N_4982,In_1161,In_109);
and U4983 (N_4983,In_1362,In_552);
xor U4984 (N_4984,In_1285,In_388);
nand U4985 (N_4985,In_425,In_1485);
nor U4986 (N_4986,In_1057,In_1134);
or U4987 (N_4987,In_1229,In_445);
xnor U4988 (N_4988,In_1781,In_795);
and U4989 (N_4989,In_445,In_160);
or U4990 (N_4990,In_1806,In_1617);
nor U4991 (N_4991,In_984,In_1104);
nor U4992 (N_4992,In_396,In_1747);
nor U4993 (N_4993,In_1557,In_1037);
nor U4994 (N_4994,In_1622,In_749);
nor U4995 (N_4995,In_463,In_1417);
and U4996 (N_4996,In_847,In_1931);
or U4997 (N_4997,In_1254,In_1879);
nand U4998 (N_4998,In_1062,In_1193);
nand U4999 (N_4999,In_1670,In_1585);
nand U5000 (N_5000,N_2136,N_1818);
nor U5001 (N_5001,N_1794,N_4327);
nand U5002 (N_5002,N_3330,N_4113);
xor U5003 (N_5003,N_1123,N_616);
and U5004 (N_5004,N_3966,N_2854);
nor U5005 (N_5005,N_3210,N_4886);
and U5006 (N_5006,N_3826,N_4084);
or U5007 (N_5007,N_519,N_3683);
or U5008 (N_5008,N_1457,N_3470);
xor U5009 (N_5009,N_2964,N_2418);
xor U5010 (N_5010,N_1115,N_4805);
nor U5011 (N_5011,N_922,N_1541);
or U5012 (N_5012,N_3660,N_1645);
nand U5013 (N_5013,N_3334,N_4118);
and U5014 (N_5014,N_2923,N_1079);
and U5015 (N_5015,N_681,N_2844);
or U5016 (N_5016,N_4640,N_4900);
xor U5017 (N_5017,N_908,N_4937);
and U5018 (N_5018,N_1395,N_3746);
xnor U5019 (N_5019,N_3578,N_1742);
xor U5020 (N_5020,N_2201,N_4442);
and U5021 (N_5021,N_2540,N_714);
and U5022 (N_5022,N_2877,N_1705);
nor U5023 (N_5023,N_206,N_1325);
nand U5024 (N_5024,N_234,N_4148);
nor U5025 (N_5025,N_3739,N_2238);
and U5026 (N_5026,N_1548,N_831);
nand U5027 (N_5027,N_3290,N_4379);
and U5028 (N_5028,N_3544,N_770);
or U5029 (N_5029,N_4976,N_3878);
and U5030 (N_5030,N_1148,N_2782);
or U5031 (N_5031,N_1721,N_3235);
and U5032 (N_5032,N_4581,N_2938);
xnor U5033 (N_5033,N_2525,N_2465);
xnor U5034 (N_5034,N_3644,N_2118);
or U5035 (N_5035,N_2441,N_2889);
nor U5036 (N_5036,N_574,N_2348);
or U5037 (N_5037,N_703,N_1108);
or U5038 (N_5038,N_1062,N_940);
and U5039 (N_5039,N_1257,N_2448);
nor U5040 (N_5040,N_4866,N_4566);
or U5041 (N_5041,N_2506,N_3575);
or U5042 (N_5042,N_4445,N_3383);
or U5043 (N_5043,N_3159,N_4396);
nand U5044 (N_5044,N_59,N_1194);
and U5045 (N_5045,N_3521,N_466);
xor U5046 (N_5046,N_1241,N_285);
xor U5047 (N_5047,N_4429,N_4486);
and U5048 (N_5048,N_2994,N_2583);
nor U5049 (N_5049,N_1909,N_634);
and U5050 (N_5050,N_2934,N_4249);
xnor U5051 (N_5051,N_4035,N_1475);
xor U5052 (N_5052,N_540,N_1055);
or U5053 (N_5053,N_1432,N_3526);
xnor U5054 (N_5054,N_2288,N_926);
nand U5055 (N_5055,N_3753,N_807);
nand U5056 (N_5056,N_4018,N_1379);
and U5057 (N_5057,N_3111,N_687);
or U5058 (N_5058,N_1571,N_4220);
nand U5059 (N_5059,N_3052,N_4408);
or U5060 (N_5060,N_1380,N_3907);
or U5061 (N_5061,N_4724,N_788);
nor U5062 (N_5062,N_4876,N_3423);
nor U5063 (N_5063,N_1514,N_3310);
nand U5064 (N_5064,N_1833,N_4114);
and U5065 (N_5065,N_1303,N_638);
nor U5066 (N_5066,N_839,N_512);
and U5067 (N_5067,N_4940,N_2237);
xnor U5068 (N_5068,N_4434,N_643);
and U5069 (N_5069,N_546,N_2191);
or U5070 (N_5070,N_2622,N_1993);
or U5071 (N_5071,N_2295,N_580);
or U5072 (N_5072,N_2900,N_1799);
or U5073 (N_5073,N_3469,N_538);
xor U5074 (N_5074,N_4037,N_2912);
nand U5075 (N_5075,N_2235,N_4490);
or U5076 (N_5076,N_463,N_2343);
nand U5077 (N_5077,N_828,N_259);
nand U5078 (N_5078,N_1785,N_1586);
nand U5079 (N_5079,N_2204,N_2944);
and U5080 (N_5080,N_1052,N_3938);
xnor U5081 (N_5081,N_2513,N_3172);
or U5082 (N_5082,N_452,N_1805);
nor U5083 (N_5083,N_31,N_4013);
nor U5084 (N_5084,N_3054,N_2231);
nor U5085 (N_5085,N_1838,N_2217);
nor U5086 (N_5086,N_3463,N_3563);
xnor U5087 (N_5087,N_2268,N_1498);
xor U5088 (N_5088,N_4304,N_4675);
xor U5089 (N_5089,N_3695,N_2323);
or U5090 (N_5090,N_1458,N_2248);
nand U5091 (N_5091,N_3078,N_371);
or U5092 (N_5092,N_1916,N_1998);
xor U5093 (N_5093,N_2797,N_1627);
and U5094 (N_5094,N_2134,N_1864);
or U5095 (N_5095,N_3097,N_4115);
or U5096 (N_5096,N_3299,N_4131);
and U5097 (N_5097,N_1210,N_2765);
and U5098 (N_5098,N_2063,N_146);
or U5099 (N_5099,N_360,N_4927);
nor U5100 (N_5100,N_1015,N_4189);
or U5101 (N_5101,N_4286,N_786);
or U5102 (N_5102,N_1246,N_4687);
xor U5103 (N_5103,N_3253,N_3029);
xnor U5104 (N_5104,N_2753,N_559);
xnor U5105 (N_5105,N_3934,N_3178);
or U5106 (N_5106,N_484,N_2332);
nand U5107 (N_5107,N_3741,N_4748);
nor U5108 (N_5108,N_3760,N_3239);
xnor U5109 (N_5109,N_4266,N_1016);
and U5110 (N_5110,N_809,N_3967);
or U5111 (N_5111,N_2074,N_3522);
xor U5112 (N_5112,N_4596,N_1206);
nand U5113 (N_5113,N_3602,N_3217);
nand U5114 (N_5114,N_2549,N_384);
or U5115 (N_5115,N_2858,N_2747);
nand U5116 (N_5116,N_261,N_232);
and U5117 (N_5117,N_4849,N_305);
or U5118 (N_5118,N_4673,N_2030);
or U5119 (N_5119,N_4419,N_4955);
and U5120 (N_5120,N_986,N_2672);
xor U5121 (N_5121,N_4850,N_3059);
nand U5122 (N_5122,N_3020,N_3140);
and U5123 (N_5123,N_2031,N_4345);
or U5124 (N_5124,N_4284,N_4425);
and U5125 (N_5125,N_674,N_4941);
and U5126 (N_5126,N_17,N_1463);
xnor U5127 (N_5127,N_622,N_1328);
nand U5128 (N_5128,N_4470,N_4781);
nor U5129 (N_5129,N_980,N_4293);
and U5130 (N_5130,N_2629,N_4219);
xor U5131 (N_5131,N_2094,N_605);
nand U5132 (N_5132,N_2957,N_3603);
xnor U5133 (N_5133,N_3839,N_999);
nor U5134 (N_5134,N_2654,N_298);
and U5135 (N_5135,N_74,N_260);
nor U5136 (N_5136,N_2645,N_3809);
nor U5137 (N_5137,N_2636,N_101);
xor U5138 (N_5138,N_1099,N_3361);
and U5139 (N_5139,N_4819,N_4611);
and U5140 (N_5140,N_887,N_2628);
or U5141 (N_5141,N_4183,N_600);
xor U5142 (N_5142,N_2970,N_3411);
nor U5143 (N_5143,N_3884,N_2649);
nor U5144 (N_5144,N_2452,N_725);
nand U5145 (N_5145,N_2499,N_1740);
nor U5146 (N_5146,N_3388,N_2675);
nor U5147 (N_5147,N_856,N_4202);
or U5148 (N_5148,N_2868,N_207);
nand U5149 (N_5149,N_2001,N_675);
or U5150 (N_5150,N_2907,N_2976);
or U5151 (N_5151,N_416,N_3498);
xor U5152 (N_5152,N_3674,N_1832);
xnor U5153 (N_5153,N_3297,N_453);
nand U5154 (N_5154,N_2692,N_1130);
xnor U5155 (N_5155,N_4593,N_1327);
and U5156 (N_5156,N_3780,N_4815);
nor U5157 (N_5157,N_2977,N_4760);
nand U5158 (N_5158,N_2402,N_3721);
and U5159 (N_5159,N_2334,N_2808);
nand U5160 (N_5160,N_1543,N_3110);
nand U5161 (N_5161,N_4936,N_4125);
nand U5162 (N_5162,N_239,N_1215);
xor U5163 (N_5163,N_3833,N_276);
nor U5164 (N_5164,N_1531,N_3138);
xnor U5165 (N_5165,N_4464,N_404);
or U5166 (N_5166,N_3853,N_156);
nand U5167 (N_5167,N_2006,N_1193);
nand U5168 (N_5168,N_1101,N_2515);
nand U5169 (N_5169,N_2177,N_3616);
nand U5170 (N_5170,N_4973,N_4375);
or U5171 (N_5171,N_721,N_2982);
nor U5172 (N_5172,N_1520,N_93);
xnor U5173 (N_5173,N_4367,N_1390);
and U5174 (N_5174,N_3195,N_2487);
and U5175 (N_5175,N_248,N_625);
or U5176 (N_5176,N_1716,N_4440);
nor U5177 (N_5177,N_222,N_3272);
nand U5178 (N_5178,N_2014,N_4845);
nor U5179 (N_5179,N_3656,N_3148);
nand U5180 (N_5180,N_2953,N_2059);
or U5181 (N_5181,N_1105,N_3992);
nand U5182 (N_5182,N_1988,N_1782);
or U5183 (N_5183,N_3363,N_3598);
or U5184 (N_5184,N_1985,N_1124);
nor U5185 (N_5185,N_3803,N_3911);
xor U5186 (N_5186,N_1885,N_1011);
nand U5187 (N_5187,N_1027,N_79);
xnor U5188 (N_5188,N_697,N_428);
xor U5189 (N_5189,N_3731,N_746);
and U5190 (N_5190,N_1230,N_4101);
xor U5191 (N_5191,N_4280,N_907);
or U5192 (N_5192,N_2149,N_4506);
xor U5193 (N_5193,N_70,N_1237);
nor U5194 (N_5194,N_2872,N_845);
nor U5195 (N_5195,N_1147,N_2038);
xor U5196 (N_5196,N_1787,N_4315);
and U5197 (N_5197,N_4816,N_1236);
nor U5198 (N_5198,N_2621,N_1508);
xor U5199 (N_5199,N_2123,N_4086);
xnor U5200 (N_5200,N_4311,N_2971);
nand U5201 (N_5201,N_602,N_4128);
and U5202 (N_5202,N_4667,N_4617);
nor U5203 (N_5203,N_1707,N_2545);
or U5204 (N_5204,N_4601,N_2918);
nand U5205 (N_5205,N_628,N_1069);
and U5206 (N_5206,N_2202,N_1876);
or U5207 (N_5207,N_3662,N_1681);
xnor U5208 (N_5208,N_4205,N_1150);
nand U5209 (N_5209,N_2531,N_2043);
or U5210 (N_5210,N_2798,N_3390);
xor U5211 (N_5211,N_1001,N_2406);
xor U5212 (N_5212,N_383,N_571);
and U5213 (N_5213,N_4503,N_797);
nand U5214 (N_5214,N_2679,N_1023);
nor U5215 (N_5215,N_1720,N_1933);
nor U5216 (N_5216,N_1638,N_3023);
xnor U5217 (N_5217,N_4420,N_2085);
nor U5218 (N_5218,N_1251,N_3407);
nor U5219 (N_5219,N_4576,N_3086);
nand U5220 (N_5220,N_4481,N_1595);
xor U5221 (N_5221,N_724,N_537);
nand U5222 (N_5222,N_2389,N_3332);
nor U5223 (N_5223,N_2641,N_4435);
nor U5224 (N_5224,N_4550,N_4681);
or U5225 (N_5225,N_3730,N_249);
nand U5226 (N_5226,N_4625,N_4599);
and U5227 (N_5227,N_3800,N_2005);
nor U5228 (N_5228,N_4789,N_4061);
and U5229 (N_5229,N_1316,N_4361);
or U5230 (N_5230,N_1704,N_4378);
and U5231 (N_5231,N_491,N_1051);
xnor U5232 (N_5232,N_796,N_4144);
nor U5233 (N_5233,N_561,N_1481);
nand U5234 (N_5234,N_2646,N_3315);
xnor U5235 (N_5235,N_4334,N_2607);
xor U5236 (N_5236,N_4338,N_4465);
xor U5237 (N_5237,N_4364,N_1323);
xor U5238 (N_5238,N_3693,N_1986);
nand U5239 (N_5239,N_753,N_3336);
or U5240 (N_5240,N_1228,N_567);
or U5241 (N_5241,N_4331,N_4431);
nor U5242 (N_5242,N_2785,N_526);
xnor U5243 (N_5243,N_4691,N_1609);
xnor U5244 (N_5244,N_3251,N_2392);
nand U5245 (N_5245,N_1250,N_3894);
nand U5246 (N_5246,N_1753,N_1593);
nor U5247 (N_5247,N_765,N_3179);
or U5248 (N_5248,N_800,N_1533);
nor U5249 (N_5249,N_1219,N_495);
or U5250 (N_5250,N_541,N_1830);
or U5251 (N_5251,N_3948,N_4105);
and U5252 (N_5252,N_1562,N_1668);
xnor U5253 (N_5253,N_1343,N_2486);
nor U5254 (N_5254,N_3200,N_2444);
xnor U5255 (N_5255,N_2779,N_2829);
and U5256 (N_5256,N_4081,N_3044);
or U5257 (N_5257,N_4902,N_1601);
and U5258 (N_5258,N_3050,N_2309);
and U5259 (N_5259,N_2055,N_4723);
nor U5260 (N_5260,N_3830,N_2774);
and U5261 (N_5261,N_4042,N_2256);
nor U5262 (N_5262,N_2065,N_2954);
nor U5263 (N_5263,N_3512,N_1085);
nand U5264 (N_5264,N_3011,N_3220);
nand U5265 (N_5265,N_3331,N_668);
nor U5266 (N_5266,N_3565,N_711);
xor U5267 (N_5267,N_326,N_1403);
or U5268 (N_5268,N_1300,N_1112);
nand U5269 (N_5269,N_492,N_439);
xnor U5270 (N_5270,N_4837,N_465);
xor U5271 (N_5271,N_2521,N_565);
nor U5272 (N_5272,N_4256,N_3633);
or U5273 (N_5273,N_197,N_792);
and U5274 (N_5274,N_1033,N_60);
or U5275 (N_5275,N_2058,N_3484);
and U5276 (N_5276,N_784,N_1731);
xor U5277 (N_5277,N_2351,N_252);
or U5278 (N_5278,N_3122,N_4136);
nand U5279 (N_5279,N_3196,N_472);
nand U5280 (N_5280,N_1895,N_3678);
xor U5281 (N_5281,N_3751,N_1911);
or U5282 (N_5282,N_3728,N_505);
nand U5283 (N_5283,N_4689,N_3124);
nor U5284 (N_5284,N_4762,N_1470);
nor U5285 (N_5285,N_504,N_3344);
nand U5286 (N_5286,N_1817,N_1814);
xnor U5287 (N_5287,N_2956,N_544);
xor U5288 (N_5288,N_2220,N_587);
nand U5289 (N_5289,N_3924,N_4478);
nand U5290 (N_5290,N_2955,N_3065);
nand U5291 (N_5291,N_22,N_368);
and U5292 (N_5292,N_3556,N_296);
or U5293 (N_5293,N_4127,N_506);
nor U5294 (N_5294,N_2875,N_4180);
nand U5295 (N_5295,N_1734,N_4967);
and U5296 (N_5296,N_3087,N_4926);
and U5297 (N_5297,N_2169,N_3600);
and U5298 (N_5298,N_3379,N_240);
xnor U5299 (N_5299,N_4143,N_1955);
nand U5300 (N_5300,N_4444,N_3520);
and U5301 (N_5301,N_1169,N_4476);
nor U5302 (N_5302,N_4836,N_4264);
nand U5303 (N_5303,N_2437,N_3726);
xor U5304 (N_5304,N_2674,N_4177);
nor U5305 (N_5305,N_852,N_362);
nand U5306 (N_5306,N_4300,N_1862);
and U5307 (N_5307,N_4810,N_2473);
xnor U5308 (N_5308,N_3434,N_1413);
and U5309 (N_5309,N_3776,N_695);
nor U5310 (N_5310,N_3748,N_3798);
nor U5311 (N_5311,N_755,N_3108);
nor U5312 (N_5312,N_4366,N_2575);
xor U5313 (N_5313,N_2130,N_2847);
or U5314 (N_5314,N_94,N_2713);
nor U5315 (N_5315,N_2544,N_4226);
nand U5316 (N_5316,N_3387,N_2366);
nand U5317 (N_5317,N_402,N_757);
nand U5318 (N_5318,N_4620,N_2377);
nand U5319 (N_5319,N_1559,N_2972);
and U5320 (N_5320,N_3533,N_1240);
or U5321 (N_5321,N_4775,N_2383);
or U5322 (N_5322,N_2456,N_3652);
xnor U5323 (N_5323,N_2269,N_4504);
nand U5324 (N_5324,N_1155,N_2120);
xnor U5325 (N_5325,N_4879,N_1837);
and U5326 (N_5326,N_1198,N_564);
xnor U5327 (N_5327,N_4947,N_1329);
or U5328 (N_5328,N_434,N_814);
or U5329 (N_5329,N_4371,N_886);
nand U5330 (N_5330,N_3278,N_4090);
and U5331 (N_5331,N_3669,N_4210);
nor U5332 (N_5332,N_773,N_2990);
xor U5333 (N_5333,N_1987,N_2585);
and U5334 (N_5334,N_4492,N_352);
nand U5335 (N_5335,N_900,N_1089);
or U5336 (N_5336,N_4817,N_2436);
nand U5337 (N_5337,N_1423,N_3064);
and U5338 (N_5338,N_3041,N_2812);
or U5339 (N_5339,N_1965,N_3567);
nor U5340 (N_5340,N_467,N_3441);
xnor U5341 (N_5341,N_4795,N_861);
xor U5342 (N_5342,N_1715,N_4227);
or U5343 (N_5343,N_1450,N_1293);
or U5344 (N_5344,N_586,N_1968);
nor U5345 (N_5345,N_461,N_3864);
and U5346 (N_5346,N_915,N_2037);
or U5347 (N_5347,N_1188,N_3818);
nand U5348 (N_5348,N_2440,N_336);
nand U5349 (N_5349,N_3127,N_767);
and U5350 (N_5350,N_2686,N_89);
nand U5351 (N_5351,N_1451,N_4875);
nand U5352 (N_5352,N_826,N_3827);
xor U5353 (N_5353,N_4905,N_4911);
and U5354 (N_5354,N_2589,N_2292);
or U5355 (N_5355,N_4642,N_4979);
nor U5356 (N_5356,N_1739,N_719);
xnor U5357 (N_5357,N_2767,N_737);
xnor U5358 (N_5358,N_1798,N_1920);
xnor U5359 (N_5359,N_1407,N_4864);
nor U5360 (N_5360,N_1331,N_3506);
or U5361 (N_5361,N_4708,N_2310);
nor U5362 (N_5362,N_3625,N_3175);
or U5363 (N_5363,N_14,N_3569);
nor U5364 (N_5364,N_859,N_40);
and U5365 (N_5365,N_2626,N_679);
and U5366 (N_5366,N_4600,N_3893);
or U5367 (N_5367,N_1262,N_2601);
nand U5368 (N_5368,N_4421,N_2624);
nor U5369 (N_5369,N_3141,N_1603);
and U5370 (N_5370,N_3667,N_3339);
xnor U5371 (N_5371,N_3237,N_3984);
xnor U5372 (N_5372,N_851,N_1845);
nor U5373 (N_5373,N_983,N_2229);
and U5374 (N_5374,N_245,N_1274);
nor U5375 (N_5375,N_392,N_4904);
xnor U5376 (N_5376,N_1696,N_3790);
nand U5377 (N_5377,N_2443,N_4551);
nand U5378 (N_5378,N_202,N_3550);
and U5379 (N_5379,N_573,N_995);
nor U5380 (N_5380,N_2153,N_2532);
nand U5381 (N_5381,N_3416,N_1127);
or U5382 (N_5382,N_1633,N_1644);
or U5383 (N_5383,N_2261,N_1733);
or U5384 (N_5384,N_3996,N_1528);
xnor U5385 (N_5385,N_902,N_4591);
or U5386 (N_5386,N_4910,N_3534);
xor U5387 (N_5387,N_2281,N_3362);
xor U5388 (N_5388,N_1133,N_3255);
nand U5389 (N_5389,N_2744,N_1128);
or U5390 (N_5390,N_2635,N_4323);
xor U5391 (N_5391,N_4228,N_1036);
nand U5392 (N_5392,N_1984,N_3910);
or U5393 (N_5393,N_3002,N_2565);
nor U5394 (N_5394,N_4867,N_2018);
and U5395 (N_5395,N_2145,N_1999);
xor U5396 (N_5396,N_297,N_3164);
nand U5397 (N_5397,N_386,N_3295);
xnor U5398 (N_5398,N_4637,N_4363);
xnor U5399 (N_5399,N_2630,N_2394);
or U5400 (N_5400,N_4075,N_2299);
and U5401 (N_5401,N_2080,N_4531);
or U5402 (N_5402,N_4423,N_4702);
xnor U5403 (N_5403,N_1442,N_3129);
nand U5404 (N_5404,N_819,N_2328);
and U5405 (N_5405,N_1482,N_4071);
or U5406 (N_5406,N_3980,N_4843);
xor U5407 (N_5407,N_3004,N_2225);
nand U5408 (N_5408,N_4489,N_4062);
or U5409 (N_5409,N_4052,N_1936);
and U5410 (N_5410,N_1095,N_1340);
nor U5411 (N_5411,N_3326,N_4703);
and U5412 (N_5412,N_2340,N_4610);
or U5413 (N_5413,N_3048,N_1163);
xnor U5414 (N_5414,N_1378,N_1007);
xnor U5415 (N_5415,N_2042,N_2083);
nand U5416 (N_5416,N_609,N_3703);
nand U5417 (N_5417,N_4627,N_4415);
and U5418 (N_5418,N_2886,N_3347);
nand U5419 (N_5419,N_1118,N_3187);
nor U5420 (N_5420,N_1302,N_4178);
or U5421 (N_5421,N_3529,N_3382);
nand U5422 (N_5422,N_3699,N_1225);
or U5423 (N_5423,N_2246,N_637);
nand U5424 (N_5424,N_3262,N_4651);
nand U5425 (N_5425,N_2947,N_2416);
xnor U5426 (N_5426,N_4840,N_2690);
xor U5427 (N_5427,N_3051,N_2572);
nand U5428 (N_5428,N_4368,N_1973);
or U5429 (N_5429,N_3579,N_947);
and U5430 (N_5430,N_2073,N_4253);
nor U5431 (N_5431,N_1354,N_4006);
nand U5432 (N_5432,N_2845,N_3228);
xnor U5433 (N_5433,N_2039,N_656);
nor U5434 (N_5434,N_1088,N_3213);
nand U5435 (N_5435,N_3482,N_2285);
and U5436 (N_5436,N_4729,N_4482);
nand U5437 (N_5437,N_2175,N_1960);
or U5438 (N_5438,N_2514,N_4682);
and U5439 (N_5439,N_821,N_1426);
and U5440 (N_5440,N_2656,N_3045);
xnor U5441 (N_5441,N_718,N_4669);
and U5442 (N_5442,N_1978,N_2324);
and U5443 (N_5443,N_1264,N_4523);
and U5444 (N_5444,N_3063,N_2099);
and U5445 (N_5445,N_4484,N_3510);
nand U5446 (N_5446,N_1848,N_361);
or U5447 (N_5447,N_2391,N_4285);
or U5448 (N_5448,N_4138,N_1077);
nand U5449 (N_5449,N_2476,N_589);
nor U5450 (N_5450,N_335,N_1856);
nor U5451 (N_5451,N_4170,N_4332);
nor U5452 (N_5452,N_2438,N_3926);
nand U5453 (N_5453,N_33,N_647);
or U5454 (N_5454,N_2325,N_575);
nor U5455 (N_5455,N_1653,N_3345);
nor U5456 (N_5456,N_3152,N_4535);
and U5457 (N_5457,N_80,N_3821);
or U5458 (N_5458,N_1614,N_179);
xnor U5459 (N_5459,N_3929,N_2403);
nand U5460 (N_5460,N_4545,N_401);
or U5461 (N_5461,N_3904,N_4918);
xor U5462 (N_5462,N_3585,N_3712);
or U5463 (N_5463,N_910,N_3873);
nor U5464 (N_5464,N_568,N_3994);
nand U5465 (N_5465,N_1345,N_2909);
xnor U5466 (N_5466,N_1672,N_2313);
xor U5467 (N_5467,N_1440,N_177);
nand U5468 (N_5468,N_3875,N_2411);
xor U5469 (N_5469,N_4389,N_4142);
xnor U5470 (N_5470,N_3626,N_4383);
nand U5471 (N_5471,N_1892,N_3426);
and U5472 (N_5472,N_4337,N_2801);
nor U5473 (N_5473,N_1290,N_3915);
and U5474 (N_5474,N_2122,N_698);
nor U5475 (N_5475,N_268,N_1822);
xor U5476 (N_5476,N_3927,N_2528);
and U5477 (N_5477,N_1552,N_1493);
and U5478 (N_5478,N_4255,N_2148);
or U5479 (N_5479,N_1752,N_112);
xnor U5480 (N_5480,N_1454,N_1282);
nor U5481 (N_5481,N_3692,N_4381);
nor U5482 (N_5482,N_3499,N_4290);
or U5483 (N_5483,N_794,N_2932);
nand U5484 (N_5484,N_4921,N_2358);
or U5485 (N_5485,N_1092,N_3083);
xor U5486 (N_5486,N_1082,N_516);
xor U5487 (N_5487,N_3198,N_144);
nor U5488 (N_5488,N_3930,N_4044);
nor U5489 (N_5489,N_3885,N_2570);
and U5490 (N_5490,N_3012,N_3612);
and U5491 (N_5491,N_1630,N_2210);
nand U5492 (N_5492,N_131,N_2578);
nor U5493 (N_5493,N_3010,N_3417);
or U5494 (N_5494,N_2454,N_929);
xnor U5495 (N_5495,N_2236,N_2103);
and U5496 (N_5496,N_2825,N_1900);
xnor U5497 (N_5497,N_2260,N_3158);
nor U5498 (N_5498,N_1622,N_2710);
and U5499 (N_5499,N_1268,N_1438);
or U5500 (N_5500,N_4742,N_1466);
xor U5501 (N_5501,N_1418,N_766);
and U5502 (N_5502,N_665,N_3707);
or U5503 (N_5503,N_4158,N_1065);
nand U5504 (N_5504,N_2209,N_1244);
nand U5505 (N_5505,N_4318,N_229);
xor U5506 (N_5506,N_1640,N_2963);
nor U5507 (N_5507,N_3778,N_1298);
and U5508 (N_5508,N_2208,N_4680);
nand U5509 (N_5509,N_1979,N_3524);
and U5510 (N_5510,N_633,N_1485);
nor U5511 (N_5511,N_1540,N_2523);
and U5512 (N_5512,N_3370,N_1137);
xnor U5513 (N_5513,N_1373,N_1249);
xor U5514 (N_5514,N_3306,N_3337);
xor U5515 (N_5515,N_4353,N_2771);
xnor U5516 (N_5516,N_1151,N_4741);
or U5517 (N_5517,N_2841,N_832);
and U5518 (N_5518,N_1404,N_458);
nor U5519 (N_5519,N_3348,N_646);
xor U5520 (N_5520,N_4961,N_4502);
nand U5521 (N_5521,N_1326,N_1879);
xor U5522 (N_5522,N_3130,N_1878);
or U5523 (N_5523,N_3705,N_497);
xnor U5524 (N_5524,N_918,N_167);
nand U5525 (N_5525,N_1256,N_2051);
nand U5526 (N_5526,N_1589,N_2067);
nor U5527 (N_5527,N_4073,N_4661);
or U5528 (N_5528,N_4913,N_3562);
or U5529 (N_5529,N_210,N_263);
and U5530 (N_5530,N_549,N_3225);
nand U5531 (N_5531,N_606,N_4467);
and U5532 (N_5532,N_3385,N_1171);
nor U5533 (N_5533,N_1714,N_115);
and U5534 (N_5534,N_2471,N_4494);
and U5535 (N_5535,N_4069,N_196);
xor U5536 (N_5536,N_2161,N_1098);
xor U5537 (N_5537,N_4639,N_812);
xor U5538 (N_5538,N_288,N_4515);
nor U5539 (N_5539,N_2106,N_4152);
and U5540 (N_5540,N_4761,N_295);
nor U5541 (N_5541,N_2985,N_141);
xor U5542 (N_5542,N_3824,N_4313);
or U5543 (N_5543,N_1170,N_4861);
and U5544 (N_5544,N_653,N_1229);
and U5545 (N_5545,N_328,N_1060);
nand U5546 (N_5546,N_2722,N_3836);
xor U5547 (N_5547,N_1392,N_4046);
nand U5548 (N_5548,N_3651,N_2553);
nand U5549 (N_5549,N_464,N_1405);
and U5550 (N_5550,N_1565,N_4995);
and U5551 (N_5551,N_2772,N_2180);
nor U5552 (N_5552,N_1063,N_318);
xnor U5553 (N_5553,N_3874,N_2640);
and U5554 (N_5554,N_2509,N_496);
xor U5555 (N_5555,N_2386,N_4745);
nor U5556 (N_5556,N_28,N_4088);
xnor U5557 (N_5557,N_837,N_3223);
and U5558 (N_5558,N_3089,N_1834);
and U5559 (N_5559,N_3160,N_2759);
nand U5560 (N_5560,N_787,N_1859);
and U5561 (N_5561,N_3287,N_1336);
and U5562 (N_5562,N_3723,N_2791);
xnor U5563 (N_5563,N_91,N_3823);
and U5564 (N_5564,N_2969,N_2850);
nand U5565 (N_5565,N_1026,N_2593);
and U5566 (N_5566,N_2302,N_2962);
xnor U5567 (N_5567,N_4856,N_4471);
or U5568 (N_5568,N_3664,N_289);
or U5569 (N_5569,N_4700,N_3869);
or U5570 (N_5570,N_4824,N_4335);
nor U5571 (N_5571,N_3744,N_3954);
and U5572 (N_5572,N_4278,N_2387);
xnor U5573 (N_5573,N_3952,N_1573);
nand U5574 (N_5574,N_2836,N_4823);
and U5575 (N_5575,N_4908,N_2614);
nor U5576 (N_5576,N_3219,N_98);
nor U5577 (N_5577,N_2318,N_4507);
xnor U5578 (N_5578,N_1521,N_3451);
nand U5579 (N_5579,N_3149,N_2355);
and U5580 (N_5580,N_4070,N_1996);
or U5581 (N_5581,N_2211,N_3921);
nand U5582 (N_5582,N_836,N_1261);
xnor U5583 (N_5583,N_1529,N_170);
or U5584 (N_5584,N_3335,N_1471);
xor U5585 (N_5585,N_4384,N_1104);
nand U5586 (N_5586,N_990,N_716);
nand U5587 (N_5587,N_710,N_2587);
or U5588 (N_5588,N_4009,N_2110);
nor U5589 (N_5589,N_2735,N_1808);
and U5590 (N_5590,N_4533,N_3756);
and U5591 (N_5591,N_1365,N_2749);
or U5592 (N_5592,N_1538,N_3324);
or U5593 (N_5593,N_3338,N_1078);
and U5594 (N_5594,N_534,N_3207);
xnor U5595 (N_5595,N_4387,N_2495);
nor U5596 (N_5596,N_3489,N_3783);
nand U5597 (N_5597,N_3177,N_644);
or U5598 (N_5598,N_1263,N_2044);
xor U5599 (N_5599,N_1160,N_1929);
xnor U5600 (N_5600,N_4041,N_1969);
and U5601 (N_5601,N_3852,N_4130);
xor U5602 (N_5602,N_1967,N_2457);
nor U5603 (N_5603,N_3835,N_57);
nor U5604 (N_5604,N_1553,N_481);
or U5605 (N_5605,N_768,N_3151);
xor U5606 (N_5606,N_103,N_1692);
nand U5607 (N_5607,N_4261,N_2135);
xor U5608 (N_5608,N_3427,N_3635);
xnor U5609 (N_5609,N_2943,N_3364);
xor U5610 (N_5610,N_924,N_3995);
nor U5611 (N_5611,N_1791,N_4320);
xnor U5612 (N_5612,N_414,N_4590);
and U5613 (N_5613,N_3881,N_3504);
nor U5614 (N_5614,N_966,N_4528);
xnor U5615 (N_5615,N_551,N_1971);
xor U5616 (N_5616,N_3473,N_2516);
nor U5617 (N_5617,N_2725,N_1071);
nor U5618 (N_5618,N_585,N_331);
and U5619 (N_5619,N_2802,N_610);
nor U5620 (N_5620,N_3057,N_3000);
nor U5621 (N_5621,N_2676,N_1663);
or U5622 (N_5622,N_3845,N_4891);
nand U5623 (N_5623,N_2991,N_3190);
xor U5624 (N_5624,N_3391,N_4725);
and U5625 (N_5625,N_511,N_1810);
xnor U5626 (N_5626,N_2342,N_1361);
or U5627 (N_5627,N_1038,N_3675);
xor U5628 (N_5628,N_1804,N_2921);
nor U5629 (N_5629,N_1068,N_2093);
nand U5630 (N_5630,N_2089,N_4939);
xor U5631 (N_5631,N_3505,N_4583);
nor U5632 (N_5632,N_143,N_2517);
or U5633 (N_5633,N_3240,N_317);
xor U5634 (N_5634,N_704,N_2468);
or U5635 (N_5635,N_950,N_1578);
or U5636 (N_5636,N_1433,N_2114);
or U5637 (N_5637,N_394,N_3580);
nand U5638 (N_5638,N_3098,N_2033);
xor U5639 (N_5639,N_3284,N_1172);
or U5640 (N_5640,N_3677,N_1386);
and U5641 (N_5641,N_4848,N_4897);
nor U5642 (N_5642,N_4390,N_1939);
nor U5643 (N_5643,N_3729,N_4704);
or U5644 (N_5644,N_3947,N_1358);
nand U5645 (N_5645,N_3905,N_3525);
xnor U5646 (N_5646,N_1769,N_134);
nor U5647 (N_5647,N_3856,N_1989);
xor U5648 (N_5648,N_4514,N_2989);
and U5649 (N_5649,N_3890,N_3170);
nor U5650 (N_5650,N_1890,N_242);
xnor U5651 (N_5651,N_4530,N_2270);
xor U5652 (N_5652,N_4040,N_1469);
or U5653 (N_5653,N_3258,N_844);
xor U5654 (N_5654,N_4638,N_2760);
and U5655 (N_5655,N_3542,N_2069);
nor U5656 (N_5656,N_330,N_2866);
or U5657 (N_5657,N_225,N_880);
or U5658 (N_5658,N_2395,N_271);
nor U5659 (N_5659,N_4853,N_4912);
nand U5660 (N_5660,N_2158,N_919);
nor U5661 (N_5661,N_4965,N_378);
nand U5662 (N_5662,N_741,N_4922);
xnor U5663 (N_5663,N_2752,N_854);
xor U5664 (N_5664,N_3280,N_1192);
xor U5665 (N_5665,N_2190,N_4827);
xnor U5666 (N_5666,N_3858,N_2727);
and U5667 (N_5667,N_1736,N_4031);
and U5668 (N_5668,N_65,N_104);
xor U5669 (N_5669,N_4977,N_3714);
nand U5670 (N_5670,N_2584,N_4250);
nand U5671 (N_5671,N_642,N_1227);
and U5672 (N_5672,N_3819,N_4287);
nand U5673 (N_5673,N_860,N_303);
and U5674 (N_5674,N_4655,N_4968);
xnor U5675 (N_5675,N_2396,N_2247);
and U5676 (N_5676,N_344,N_2602);
nor U5677 (N_5677,N_4555,N_411);
and U5678 (N_5678,N_4771,N_435);
nand U5679 (N_5679,N_3991,N_294);
nand U5680 (N_5680,N_4426,N_178);
xor U5681 (N_5681,N_1394,N_1385);
nand U5682 (N_5682,N_1330,N_3913);
and U5683 (N_5683,N_3487,N_3766);
nand U5684 (N_5684,N_399,N_4239);
nor U5685 (N_5685,N_4841,N_3107);
and U5686 (N_5686,N_522,N_4929);
or U5687 (N_5687,N_412,N_238);
nor U5688 (N_5688,N_4738,N_2315);
or U5689 (N_5689,N_441,N_132);
or U5690 (N_5690,N_2420,N_3496);
nand U5691 (N_5691,N_2306,N_429);
or U5692 (N_5692,N_556,N_4559);
or U5693 (N_5693,N_3458,N_2661);
and U5694 (N_5694,N_4746,N_201);
or U5695 (N_5695,N_4350,N_4665);
xor U5696 (N_5696,N_1387,N_2398);
nand U5697 (N_5697,N_4764,N_256);
xnor U5698 (N_5698,N_3820,N_1779);
nand U5699 (N_5699,N_3492,N_2693);
nor U5700 (N_5700,N_1846,N_1216);
nand U5701 (N_5701,N_4059,N_2049);
nand U5702 (N_5702,N_430,N_158);
xnor U5703 (N_5703,N_311,N_3249);
nor U5704 (N_5704,N_989,N_4401);
nand U5705 (N_5705,N_1686,N_678);
nor U5706 (N_5706,N_2142,N_2447);
xor U5707 (N_5707,N_4699,N_2363);
nor U5708 (N_5708,N_4107,N_1319);
and U5709 (N_5709,N_3493,N_798);
nor U5710 (N_5710,N_2818,N_1143);
or U5711 (N_5711,N_142,N_3945);
or U5712 (N_5712,N_4244,N_3920);
or U5713 (N_5713,N_1995,N_2421);
and U5714 (N_5714,N_1519,N_1927);
nand U5715 (N_5715,N_1530,N_2314);
nor U5716 (N_5716,N_4829,N_3680);
nor U5717 (N_5717,N_3155,N_4398);
nand U5718 (N_5718,N_909,N_2497);
or U5719 (N_5719,N_4393,N_4433);
nand U5720 (N_5720,N_180,N_4721);
nand U5721 (N_5721,N_1534,N_3259);
nand U5722 (N_5722,N_1523,N_120);
nand U5723 (N_5723,N_2415,N_4706);
nor U5724 (N_5724,N_2748,N_4790);
nor U5725 (N_5725,N_4223,N_3745);
nand U5726 (N_5726,N_3979,N_4882);
or U5727 (N_5727,N_2880,N_272);
or U5728 (N_5728,N_2655,N_1546);
xnor U5729 (N_5729,N_3468,N_811);
or U5730 (N_5730,N_2763,N_1456);
and U5731 (N_5731,N_4151,N_1318);
xnor U5732 (N_5732,N_2155,N_4776);
or U5733 (N_5733,N_660,N_4191);
or U5734 (N_5734,N_3061,N_4728);
nand U5735 (N_5735,N_2755,N_4339);
and U5736 (N_5736,N_483,N_1976);
nand U5737 (N_5737,N_4298,N_4358);
nand U5738 (N_5738,N_4720,N_2718);
nand U5739 (N_5739,N_2401,N_4295);
or U5740 (N_5740,N_3075,N_3015);
nor U5741 (N_5741,N_164,N_3865);
and U5742 (N_5742,N_2696,N_1497);
xor U5743 (N_5743,N_2071,N_356);
nand U5744 (N_5744,N_2370,N_1179);
nor U5745 (N_5745,N_1694,N_2301);
nor U5746 (N_5746,N_4055,N_2160);
or U5747 (N_5747,N_4271,N_751);
nor U5748 (N_5748,N_3294,N_2839);
nand U5749 (N_5749,N_1308,N_1500);
and U5750 (N_5750,N_2653,N_3263);
xor U5751 (N_5751,N_2368,N_1332);
nand U5752 (N_5752,N_4449,N_4888);
and U5753 (N_5753,N_4167,N_2060);
and U5754 (N_5754,N_623,N_4446);
xnor U5755 (N_5755,N_3437,N_991);
and U5756 (N_5756,N_186,N_38);
xor U5757 (N_5757,N_4011,N_396);
nor U5758 (N_5758,N_3166,N_652);
nand U5759 (N_5759,N_494,N_3577);
or U5760 (N_5760,N_3619,N_3953);
xnor U5761 (N_5761,N_3857,N_4192);
or U5762 (N_5762,N_4996,N_897);
or U5763 (N_5763,N_645,N_1132);
nand U5764 (N_5764,N_3156,N_670);
nand U5765 (N_5765,N_608,N_4087);
or U5766 (N_5766,N_4053,N_865);
nor U5767 (N_5767,N_872,N_4262);
or U5768 (N_5768,N_2975,N_4303);
or U5769 (N_5769,N_667,N_2573);
xnor U5770 (N_5770,N_1090,N_1294);
or U5771 (N_5771,N_4564,N_3357);
or U5772 (N_5772,N_1517,N_4224);
and U5773 (N_5773,N_1221,N_4175);
nand U5774 (N_5774,N_2303,N_3768);
and U5775 (N_5775,N_1189,N_3665);
or U5776 (N_5776,N_3058,N_1258);
nand U5777 (N_5777,N_415,N_3145);
xnor U5778 (N_5778,N_4666,N_669);
and U5779 (N_5779,N_267,N_4993);
nor U5780 (N_5780,N_967,N_572);
and U5781 (N_5781,N_2960,N_4305);
nand U5782 (N_5782,N_1551,N_4459);
nor U5783 (N_5783,N_1886,N_1510);
and U5784 (N_5784,N_651,N_1877);
and U5785 (N_5785,N_4586,N_2293);
and U5786 (N_5786,N_1428,N_4754);
xnor U5787 (N_5787,N_2393,N_2009);
nand U5788 (N_5788,N_1919,N_3467);
or U5789 (N_5789,N_3474,N_1435);
xnor U5790 (N_5790,N_1676,N_4139);
and U5791 (N_5791,N_3486,N_601);
nor U5792 (N_5792,N_2683,N_2855);
nand U5793 (N_5793,N_3566,N_3131);
and U5794 (N_5794,N_1870,N_736);
xnor U5795 (N_5795,N_2305,N_3939);
xor U5796 (N_5796,N_3848,N_3409);
xnor U5797 (N_5797,N_124,N_4809);
and U5798 (N_5798,N_3784,N_763);
xnor U5799 (N_5799,N_2087,N_3188);
nor U5800 (N_5800,N_3402,N_2092);
or U5801 (N_5801,N_1030,N_3301);
or U5802 (N_5802,N_2547,N_3925);
nand U5803 (N_5803,N_4207,N_446);
nor U5804 (N_5804,N_4359,N_760);
nor U5805 (N_5805,N_4215,N_1623);
nand U5806 (N_5806,N_2959,N_2034);
or U5807 (N_5807,N_3537,N_1058);
nand U5808 (N_5808,N_1045,N_485);
or U5809 (N_5809,N_1812,N_1284);
or U5810 (N_5810,N_1159,N_655);
and U5811 (N_5811,N_4094,N_2884);
nor U5812 (N_5812,N_1688,N_47);
xor U5813 (N_5813,N_3392,N_818);
nand U5814 (N_5814,N_3084,N_2445);
and U5815 (N_5815,N_2397,N_1773);
xor U5816 (N_5816,N_140,N_3648);
nand U5817 (N_5817,N_2967,N_2478);
xnor U5818 (N_5818,N_4732,N_1117);
nor U5819 (N_5819,N_4644,N_2703);
and U5820 (N_5820,N_3772,N_4717);
xnor U5821 (N_5821,N_3530,N_2048);
or U5822 (N_5822,N_3557,N_2076);
nor U5823 (N_5823,N_3318,N_2367);
and U5824 (N_5824,N_997,N_3007);
nor U5825 (N_5825,N_4438,N_2814);
and U5826 (N_5826,N_2508,N_4240);
or U5827 (N_5827,N_193,N_4857);
and U5828 (N_5828,N_1096,N_3658);
nor U5829 (N_5829,N_3116,N_199);
and U5830 (N_5830,N_536,N_482);
and U5831 (N_5831,N_913,N_1613);
nor U5832 (N_5832,N_1367,N_1043);
nand U5833 (N_5833,N_3515,N_2891);
or U5834 (N_5834,N_2086,N_533);
nor U5835 (N_5835,N_322,N_4842);
nand U5836 (N_5836,N_1844,N_3570);
and U5837 (N_5837,N_3366,N_2778);
or U5838 (N_5838,N_1643,N_3799);
or U5839 (N_5839,N_4966,N_708);
and U5840 (N_5840,N_1374,N_4212);
xor U5841 (N_5841,N_942,N_3327);
xnor U5842 (N_5842,N_4735,N_1190);
and U5843 (N_5843,N_2978,N_4058);
xor U5844 (N_5844,N_3919,N_925);
xnor U5845 (N_5845,N_4184,N_3001);
and U5846 (N_5846,N_1047,N_3747);
and U5847 (N_5847,N_1288,N_899);
nor U5848 (N_5848,N_2029,N_3999);
and U5849 (N_5849,N_1924,N_4736);
and U5850 (N_5850,N_4737,N_1922);
nand U5851 (N_5851,N_3604,N_3475);
nor U5852 (N_5852,N_1310,N_474);
and U5853 (N_5853,N_4020,N_948);
xnor U5854 (N_5854,N_1841,N_1307);
xor U5855 (N_5855,N_1880,N_4844);
nand U5856 (N_5856,N_4710,N_2183);
and U5857 (N_5857,N_290,N_1453);
nand U5858 (N_5858,N_2036,N_2388);
nor U5859 (N_5859,N_3137,N_2434);
nand U5860 (N_5860,N_938,N_3901);
xnor U5861 (N_5861,N_713,N_3481);
nor U5862 (N_5862,N_3055,N_3169);
or U5863 (N_5863,N_2529,N_2322);
nand U5864 (N_5864,N_1254,N_372);
nand U5865 (N_5865,N_314,N_594);
or U5866 (N_5866,N_2493,N_2003);
or U5867 (N_5867,N_4034,N_3274);
xor U5868 (N_5868,N_2789,N_1382);
xor U5869 (N_5869,N_955,N_3773);
and U5870 (N_5870,N_2027,N_1144);
nor U5871 (N_5871,N_1474,N_1765);
and U5872 (N_5872,N_2706,N_3374);
or U5873 (N_5873,N_1756,N_2543);
and U5874 (N_5874,N_3880,N_3548);
or U5875 (N_5875,N_4067,N_154);
and U5876 (N_5876,N_1964,N_2171);
nand U5877 (N_5877,N_3789,N_1164);
nor U5878 (N_5878,N_1646,N_2198);
nand U5879 (N_5879,N_1362,N_857);
and U5880 (N_5880,N_820,N_3940);
nand U5881 (N_5881,N_801,N_2422);
xor U5882 (N_5882,N_2417,N_2218);
or U5883 (N_5883,N_3650,N_4102);
and U5884 (N_5884,N_2537,N_2127);
nor U5885 (N_5885,N_13,N_2806);
xor U5886 (N_5886,N_1902,N_3877);
nand U5887 (N_5887,N_3960,N_3121);
or U5888 (N_5888,N_3854,N_694);
and U5889 (N_5889,N_2151,N_578);
nand U5890 (N_5890,N_2867,N_4124);
nand U5891 (N_5891,N_3700,N_1377);
or U5892 (N_5892,N_1444,N_2412);
nand U5893 (N_5893,N_592,N_1461);
xnor U5894 (N_5894,N_2139,N_502);
and U5895 (N_5895,N_1191,N_1391);
and U5896 (N_5896,N_1728,N_3671);
or U5897 (N_5897,N_2084,N_4399);
xor U5898 (N_5898,N_370,N_2916);
or U5899 (N_5899,N_3226,N_4452);
and U5900 (N_5900,N_4214,N_2108);
and U5901 (N_5901,N_1778,N_2373);
nor U5902 (N_5902,N_964,N_1443);
and U5903 (N_5903,N_3457,N_3701);
or U5904 (N_5904,N_2463,N_312);
or U5905 (N_5905,N_777,N_3404);
xnor U5906 (N_5906,N_4302,N_457);
and U5907 (N_5907,N_4326,N_3174);
nand U5908 (N_5908,N_4063,N_4833);
or U5909 (N_5909,N_309,N_2714);
nor U5910 (N_5910,N_4536,N_2284);
nor U5911 (N_5911,N_3949,N_689);
xnor U5912 (N_5912,N_1858,N_4659);
nand U5913 (N_5913,N_847,N_2425);
nor U5914 (N_5914,N_123,N_3655);
nand U5915 (N_5915,N_4048,N_1334);
and U5916 (N_5916,N_4257,N_358);
nand U5917 (N_5917,N_1044,N_2096);
or U5918 (N_5918,N_3077,N_971);
nand U5919 (N_5919,N_1566,N_1437);
nand U5920 (N_5920,N_3807,N_2786);
xor U5921 (N_5921,N_46,N_4082);
nor U5922 (N_5922,N_4646,N_162);
or U5923 (N_5923,N_3194,N_1940);
or U5924 (N_5924,N_4989,N_4279);
nand U5925 (N_5925,N_3168,N_2946);
or U5926 (N_5926,N_2287,N_2908);
and U5927 (N_5927,N_1496,N_2253);
nor U5928 (N_5928,N_2813,N_2730);
nand U5929 (N_5929,N_2375,N_27);
nor U5930 (N_5930,N_3341,N_4356);
nor U5931 (N_5931,N_4237,N_75);
xnor U5932 (N_5932,N_3672,N_3480);
xnor U5933 (N_5933,N_11,N_1629);
xor U5934 (N_5934,N_4539,N_3369);
nor U5935 (N_5935,N_4715,N_1730);
or U5936 (N_5936,N_2477,N_3531);
nand U5937 (N_5937,N_4685,N_3613);
and U5938 (N_5938,N_1356,N_1295);
or U5939 (N_5939,N_1353,N_871);
and U5940 (N_5940,N_1218,N_4668);
nand U5941 (N_5941,N_1152,N_1906);
nand U5942 (N_5942,N_4060,N_2888);
xnor U5943 (N_5943,N_2372,N_2833);
and U5944 (N_5944,N_2466,N_3267);
or U5945 (N_5945,N_2736,N_354);
nor U5946 (N_5946,N_621,N_1723);
xnor U5947 (N_5947,N_139,N_3229);
or U5948 (N_5948,N_427,N_3444);
nor U5949 (N_5949,N_4970,N_2484);
or U5950 (N_5950,N_1611,N_3622);
nor U5951 (N_5951,N_1711,N_3476);
nand U5952 (N_5952,N_1398,N_3988);
or U5953 (N_5953,N_4162,N_1217);
or U5954 (N_5954,N_2599,N_4865);
nand U5955 (N_5955,N_3989,N_1828);
and U5956 (N_5956,N_774,N_1002);
nand U5957 (N_5957,N_509,N_1792);
xor U5958 (N_5958,N_3135,N_269);
nand U5959 (N_5959,N_745,N_649);
nand U5960 (N_5960,N_108,N_1746);
or U5961 (N_5961,N_614,N_1591);
and U5962 (N_5962,N_1337,N_2605);
nand U5963 (N_5963,N_3443,N_709);
or U5964 (N_5964,N_223,N_4768);
xor U5965 (N_5965,N_418,N_3973);
nand U5966 (N_5966,N_3264,N_4803);
xnor U5967 (N_5967,N_3452,N_3628);
or U5968 (N_5968,N_1816,N_228);
xor U5969 (N_5969,N_1869,N_2604);
nand U5970 (N_5970,N_4416,N_3899);
nor U5971 (N_5971,N_1934,N_2929);
nor U5972 (N_5972,N_3970,N_2203);
xor U5973 (N_5973,N_2853,N_3720);
xnor U5974 (N_5974,N_1780,N_722);
and U5975 (N_5975,N_351,N_3139);
xnor U5976 (N_5976,N_4901,N_892);
xnor U5977 (N_5977,N_4362,N_42);
nor U5978 (N_5978,N_758,N_4933);
and U5979 (N_5979,N_4039,N_4773);
xnor U5980 (N_5980,N_1383,N_3424);
xor U5981 (N_5981,N_376,N_1590);
nor U5982 (N_5982,N_1706,N_2167);
or U5983 (N_5983,N_4238,N_3356);
xor U5984 (N_5984,N_3102,N_1597);
nand U5985 (N_5985,N_3408,N_1761);
nand U5986 (N_5986,N_4099,N_2878);
and U5987 (N_5987,N_4928,N_4553);
xnor U5988 (N_5988,N_2166,N_2639);
or U5989 (N_5989,N_1827,N_4005);
nor U5990 (N_5990,N_4352,N_3256);
nor U5991 (N_5991,N_1783,N_785);
or U5992 (N_5992,N_1675,N_4618);
and U5993 (N_5993,N_1835,N_3353);
and U5994 (N_5994,N_4153,N_3734);
nand U5995 (N_5995,N_4365,N_4263);
nand U5996 (N_5996,N_2615,N_515);
and U5997 (N_5997,N_3986,N_612);
nor U5998 (N_5998,N_2197,N_2339);
nand U5999 (N_5999,N_3903,N_996);
and U6000 (N_6000,N_4333,N_419);
xnor U6001 (N_6001,N_479,N_4701);
and U6002 (N_6002,N_4983,N_2491);
xnor U6003 (N_6003,N_566,N_583);
and U6004 (N_6004,N_3384,N_2399);
nand U6005 (N_6005,N_4195,N_1656);
or U6006 (N_6006,N_4281,N_1097);
nor U6007 (N_6007,N_4801,N_76);
nor U6008 (N_6008,N_894,N_1156);
or U6009 (N_6009,N_4571,N_539);
xor U6010 (N_6010,N_4050,N_1991);
or U6011 (N_6011,N_1954,N_3862);
xor U6012 (N_6012,N_1650,N_1139);
and U6013 (N_6013,N_2053,N_3816);
or U6014 (N_6014,N_2409,N_4150);
and U6015 (N_6015,N_1824,N_4314);
nor U6016 (N_6016,N_1793,N_2337);
nor U6017 (N_6017,N_2873,N_1806);
nor U6018 (N_6018,N_2914,N_4372);
xor U6019 (N_6019,N_2899,N_3405);
and U6020 (N_6020,N_2939,N_3153);
and U6021 (N_6021,N_1131,N_215);
nand U6022 (N_6022,N_3277,N_3112);
xor U6023 (N_6023,N_438,N_2280);
nand U6024 (N_6024,N_3822,N_175);
and U6025 (N_6025,N_2439,N_395);
xor U6026 (N_6026,N_4999,N_4510);
xor U6027 (N_6027,N_3211,N_1401);
and U6028 (N_6028,N_993,N_476);
and U6029 (N_6029,N_55,N_1901);
and U6030 (N_6030,N_715,N_1866);
nor U6031 (N_6031,N_171,N_2600);
xnor U6032 (N_6032,N_2199,N_1464);
xnor U6033 (N_6033,N_1154,N_1434);
or U6034 (N_6034,N_4294,N_1871);
or U6035 (N_6035,N_2382,N_635);
and U6036 (N_6036,N_2128,N_4194);
nand U6037 (N_6037,N_1355,N_1350);
nor U6038 (N_6038,N_4552,N_2079);
or U6039 (N_6039,N_2896,N_4095);
nor U6040 (N_6040,N_4217,N_1882);
nand U6041 (N_6041,N_490,N_1207);
and U6042 (N_6042,N_1925,N_3053);
nor U6043 (N_6043,N_2184,N_726);
nand U6044 (N_6044,N_4649,N_3046);
nand U6045 (N_6045,N_3230,N_4163);
nand U6046 (N_6046,N_3101,N_2726);
and U6047 (N_6047,N_1182,N_96);
nand U6048 (N_6048,N_1056,N_2784);
or U6049 (N_6049,N_3896,N_1851);
or U6050 (N_6050,N_813,N_1592);
nand U6051 (N_6051,N_3922,N_604);
or U6052 (N_6052,N_4418,N_2091);
and U6053 (N_6053,N_4382,N_3191);
or U6054 (N_6054,N_3981,N_2739);
xnor U6055 (N_6055,N_3205,N_2156);
xnor U6056 (N_6056,N_1893,N_444);
nand U6057 (N_6057,N_3509,N_795);
xor U6058 (N_6058,N_4834,N_4511);
nand U6059 (N_6059,N_2795,N_1121);
and U6060 (N_6060,N_4181,N_3812);
or U6061 (N_6061,N_3410,N_1484);
or U6062 (N_6062,N_198,N_3814);
nor U6063 (N_6063,N_4549,N_2554);
nand U6064 (N_6064,N_4623,N_1048);
nand U6065 (N_6065,N_1100,N_2556);
nor U6066 (N_6066,N_1477,N_4800);
or U6067 (N_6067,N_2659,N_2068);
nand U6068 (N_6068,N_2926,N_1019);
and U6069 (N_6069,N_369,N_3583);
or U6070 (N_6070,N_4505,N_4808);
nor U6071 (N_6071,N_2937,N_3897);
and U6072 (N_6072,N_901,N_2979);
nand U6073 (N_6073,N_4868,N_883);
and U6074 (N_6074,N_1269,N_398);
and U6075 (N_6075,N_3645,N_1320);
nand U6076 (N_6076,N_4024,N_2488);
xnor U6077 (N_6077,N_870,N_3134);
or U6078 (N_6078,N_26,N_1567);
or U6079 (N_6079,N_1596,N_1935);
and U6080 (N_6080,N_4733,N_4982);
nor U6081 (N_6081,N_1324,N_304);
nor U6082 (N_6082,N_4917,N_1177);
nor U6083 (N_6083,N_2563,N_3815);
and U6084 (N_6084,N_931,N_3373);
nor U6085 (N_6085,N_4247,N_2222);
xnor U6086 (N_6086,N_3906,N_1046);
or U6087 (N_6087,N_4677,N_1990);
xnor U6088 (N_6088,N_2958,N_1974);
or U6089 (N_6089,N_3040,N_1375);
or U6090 (N_6090,N_4348,N_4126);
nand U6091 (N_6091,N_3133,N_1141);
nand U6092 (N_6092,N_863,N_3754);
xnor U6093 (N_6093,N_1569,N_3847);
nor U6094 (N_6094,N_2997,N_4543);
xnor U6095 (N_6095,N_216,N_4954);
nor U6096 (N_6096,N_2143,N_1018);
and U6097 (N_6097,N_4767,N_3208);
or U6098 (N_6098,N_1480,N_3342);
and U6099 (N_6099,N_1699,N_3245);
nand U6100 (N_6100,N_308,N_315);
and U6101 (N_6101,N_4985,N_1953);
xnor U6102 (N_6102,N_3535,N_664);
nand U6103 (N_6103,N_3381,N_4716);
or U6104 (N_6104,N_3555,N_963);
nor U6105 (N_6105,N_2272,N_2147);
and U6106 (N_6106,N_3755,N_413);
nand U6107 (N_6107,N_3244,N_2594);
xor U6108 (N_6108,N_945,N_68);
and U6109 (N_6109,N_3378,N_1560);
nor U6110 (N_6110,N_3686,N_4045);
nor U6111 (N_6111,N_3900,N_2574);
or U6112 (N_6112,N_4292,N_4664);
nand U6113 (N_6113,N_2424,N_2482);
or U6114 (N_6114,N_2408,N_442);
xor U6115 (N_6115,N_3690,N_421);
nor U6116 (N_6116,N_4632,N_2354);
or U6117 (N_6117,N_4778,N_2695);
and U6118 (N_6118,N_3808,N_1655);
or U6119 (N_6119,N_2721,N_1564);
nand U6120 (N_6120,N_1662,N_4516);
and U6121 (N_6121,N_4360,N_1712);
xor U6122 (N_6122,N_2524,N_691);
xnor U6123 (N_6123,N_4881,N_1966);
and U6124 (N_6124,N_2764,N_3302);
or U6125 (N_6125,N_2327,N_4693);
nor U6126 (N_6126,N_4930,N_4019);
xnor U6127 (N_6127,N_3840,N_4321);
or U6128 (N_6128,N_2775,N_2637);
and U6129 (N_6129,N_251,N_4705);
and U6130 (N_6130,N_4832,N_340);
and U6131 (N_6131,N_932,N_2265);
and U6132 (N_6132,N_122,N_1255);
nand U6133 (N_6133,N_95,N_3659);
nand U6134 (N_6134,N_1624,N_302);
and U6135 (N_6135,N_2510,N_2154);
nand U6136 (N_6136,N_4981,N_1700);
nor U6137 (N_6137,N_500,N_1297);
xor U6138 (N_6138,N_1421,N_3460);
nor U6139 (N_6139,N_4209,N_3183);
nand U6140 (N_6140,N_3609,N_3367);
nand U6141 (N_6141,N_2691,N_1691);
nor U6142 (N_6142,N_684,N_2965);
nand U6143 (N_6143,N_4001,N_4919);
nor U6144 (N_6144,N_4641,N_527);
nand U6145 (N_6145,N_2428,N_4235);
nor U6146 (N_6146,N_3231,N_4630);
and U6147 (N_6147,N_2152,N_4174);
xnor U6148 (N_6148,N_4615,N_3222);
or U6149 (N_6149,N_3073,N_247);
xor U6150 (N_6150,N_1944,N_4952);
and U6151 (N_6151,N_2826,N_2883);
and U6152 (N_6152,N_3975,N_2330);
nand U6153 (N_6153,N_3401,N_1685);
xnor U6154 (N_6154,N_4974,N_1505);
nand U6155 (N_6155,N_4546,N_3039);
xnor U6156 (N_6156,N_400,N_58);
nand U6157 (N_6157,N_611,N_1679);
nand U6158 (N_6158,N_2992,N_4828);
or U6159 (N_6159,N_1196,N_1669);
nor U6160 (N_6160,N_4038,N_2856);
and U6161 (N_6161,N_2530,N_3464);
nor U6162 (N_6162,N_4653,N_930);
xnor U6163 (N_6163,N_2163,N_100);
nand U6164 (N_6164,N_2518,N_2095);
nand U6165 (N_6165,N_3964,N_3181);
nor U6166 (N_6166,N_3673,N_4258);
or U6167 (N_6167,N_3455,N_4121);
xor U6168 (N_6168,N_4786,N_1826);
nand U6169 (N_6169,N_350,N_2762);
nor U6170 (N_6170,N_106,N_2407);
and U6171 (N_6171,N_4787,N_4959);
nand U6172 (N_6172,N_2689,N_3681);
xor U6173 (N_6173,N_2756,N_960);
xnor U6174 (N_6174,N_3599,N_3792);
nor U6175 (N_6175,N_3252,N_3459);
and U6176 (N_6176,N_4946,N_3796);
xnor U6177 (N_6177,N_4347,N_10);
nor U6178 (N_6178,N_2319,N_4783);
nor U6179 (N_6179,N_1422,N_2564);
or U6180 (N_6180,N_1894,N_4597);
nor U6181 (N_6181,N_1158,N_4455);
nor U6182 (N_6182,N_3421,N_393);
nand U6183 (N_6183,N_1738,N_3025);
xnor U6184 (N_6184,N_3541,N_3043);
xnor U6185 (N_6185,N_4002,N_1473);
and U6186 (N_6186,N_4274,N_173);
nand U6187 (N_6187,N_4521,N_4297);
xnor U6188 (N_6188,N_2980,N_307);
nand U6189 (N_6189,N_4674,N_961);
or U6190 (N_6190,N_275,N_4855);
and U6191 (N_6191,N_1600,N_417);
xor U6192 (N_6192,N_172,N_4785);
or U6193 (N_6193,N_2020,N_1959);
and U6194 (N_6194,N_3261,N_3511);
nand U6195 (N_6195,N_3128,N_2298);
xor U6196 (N_6196,N_2249,N_4588);
or U6197 (N_6197,N_1301,N_4734);
xor U6198 (N_6198,N_4920,N_99);
xor U6199 (N_6199,N_4770,N_1947);
nand U6200 (N_6200,N_1980,N_4906);
and U6201 (N_6201,N_283,N_4877);
nand U6202 (N_6202,N_3931,N_1080);
xnor U6203 (N_6203,N_1145,N_4146);
or U6204 (N_6204,N_250,N_1759);
and U6205 (N_6205,N_2336,N_2609);
xnor U6206 (N_6206,N_4574,N_508);
nor U6207 (N_6207,N_2291,N_4582);
nand U6208 (N_6208,N_4089,N_2851);
nand U6209 (N_6209,N_2054,N_2863);
nand U6210 (N_6210,N_1086,N_2737);
and U6211 (N_6211,N_3916,N_3944);
nor U6212 (N_6212,N_214,N_806);
or U6213 (N_6213,N_1938,N_3126);
nand U6214 (N_6214,N_4892,N_2423);
xnor U6215 (N_6215,N_4608,N_3618);
or U6216 (N_6216,N_1153,N_3019);
nor U6217 (N_6217,N_2378,N_1344);
nand U6218 (N_6218,N_4513,N_1915);
xor U6219 (N_6219,N_4199,N_3100);
xor U6220 (N_6220,N_4878,N_241);
or U6221 (N_6221,N_1896,N_4299);
or U6222 (N_6222,N_2663,N_4547);
or U6223 (N_6223,N_3495,N_4080);
nor U6224 (N_6224,N_3419,N_671);
xnor U6225 (N_6225,N_2685,N_3425);
nand U6226 (N_6226,N_4351,N_1425);
xor U6227 (N_6227,N_119,N_137);
nand U6228 (N_6228,N_3605,N_64);
and U6229 (N_6229,N_3694,N_3998);
nand U6230 (N_6230,N_174,N_525);
and U6231 (N_6231,N_3376,N_959);
and U6232 (N_6232,N_1912,N_3968);
and U6233 (N_6233,N_518,N_3418);
nor U6234 (N_6234,N_510,N_1803);
or U6235 (N_6235,N_630,N_1000);
or U6236 (N_6236,N_4245,N_3371);
and U6237 (N_6237,N_355,N_4182);
and U6238 (N_6238,N_1253,N_3641);
xor U6239 (N_6239,N_4417,N_552);
or U6240 (N_6240,N_4652,N_1223);
xnor U6241 (N_6241,N_1972,N_4769);
and U6242 (N_6242,N_3234,N_2887);
nor U6243 (N_6243,N_1185,N_804);
nand U6244 (N_6244,N_301,N_1370);
nand U6245 (N_6245,N_1125,N_1659);
and U6246 (N_6246,N_2224,N_3794);
and U6247 (N_6247,N_962,N_4893);
nor U6248 (N_6248,N_2728,N_1735);
xnor U6249 (N_6249,N_1932,N_4288);
nor U6250 (N_6250,N_917,N_1010);
xor U6251 (N_6251,N_2490,N_3883);
and U6252 (N_6252,N_3718,N_3691);
nand U6253 (N_6253,N_2019,N_2671);
nor U6254 (N_6254,N_2062,N_1744);
xnor U6255 (N_6255,N_4949,N_3113);
nand U6256 (N_6256,N_2874,N_4629);
nand U6257 (N_6257,N_1741,N_4695);
and U6258 (N_6258,N_4943,N_776);
and U6259 (N_6259,N_4462,N_2016);
nor U6260 (N_6260,N_4568,N_2250);
and U6261 (N_6261,N_3774,N_3513);
nor U6262 (N_6262,N_1073,N_3028);
or U6263 (N_6263,N_125,N_1665);
or U6264 (N_6264,N_3154,N_4054);
and U6265 (N_6265,N_2431,N_576);
nand U6266 (N_6266,N_4565,N_2405);
xor U6267 (N_6267,N_3976,N_2241);
xor U6268 (N_6268,N_982,N_3197);
or U6269 (N_6269,N_4140,N_1847);
nor U6270 (N_6270,N_1488,N_4234);
and U6271 (N_6271,N_4898,N_357);
or U6272 (N_6272,N_1606,N_1014);
nor U6273 (N_6273,N_35,N_1024);
or U6274 (N_6274,N_3066,N_2519);
nor U6275 (N_6275,N_4168,N_1187);
nand U6276 (N_6276,N_2021,N_4860);
xor U6277 (N_6277,N_885,N_4852);
or U6278 (N_6278,N_1618,N_2731);
xor U6279 (N_6279,N_2616,N_279);
nand U6280 (N_6280,N_4460,N_3247);
and U6281 (N_6281,N_1059,N_563);
nand U6282 (N_6282,N_2449,N_890);
xor U6283 (N_6283,N_2917,N_631);
or U6284 (N_6284,N_1635,N_3350);
nor U6285 (N_6285,N_2638,N_2119);
or U6286 (N_6286,N_4945,N_3879);
xor U6287 (N_6287,N_1903,N_1491);
and U6288 (N_6288,N_531,N_3785);
or U6289 (N_6289,N_1535,N_78);
and U6290 (N_6290,N_4341,N_4684);
or U6291 (N_6291,N_4395,N_1338);
and U6292 (N_6292,N_4612,N_789);
nor U6293 (N_6293,N_4584,N_650);
xor U6294 (N_6294,N_3270,N_1758);
nor U6295 (N_6295,N_3488,N_1608);
nand U6296 (N_6296,N_2859,N_3283);
xnor U6297 (N_6297,N_3666,N_4007);
xor U6298 (N_6298,N_3298,N_3553);
or U6299 (N_6299,N_4799,N_3634);
and U6300 (N_6300,N_4755,N_2193);
nand U6301 (N_6301,N_4475,N_2660);
xnor U6302 (N_6302,N_4157,N_701);
nor U6303 (N_6303,N_1369,N_881);
nand U6304 (N_6304,N_4187,N_3573);
and U6305 (N_6305,N_2650,N_3453);
and U6306 (N_6306,N_4432,N_542);
or U6307 (N_6307,N_4517,N_2112);
xor U6308 (N_6308,N_1512,N_359);
and U6309 (N_6309,N_1126,N_19);
or U6310 (N_6310,N_707,N_976);
and U6311 (N_6311,N_1279,N_2362);
nand U6312 (N_6312,N_4916,N_3850);
xor U6313 (N_6313,N_1050,N_3035);
xor U6314 (N_6314,N_4196,N_3312);
nand U6315 (N_6315,N_4686,N_4887);
or U6316 (N_6316,N_4657,N_1286);
nor U6317 (N_6317,N_4149,N_2790);
nor U6318 (N_6318,N_2981,N_332);
nor U6319 (N_6319,N_2381,N_3793);
nor U6320 (N_6320,N_4863,N_4443);
xor U6321 (N_6321,N_4122,N_4233);
nand U6322 (N_6322,N_2182,N_4036);
nor U6323 (N_6323,N_4759,N_233);
or U6324 (N_6324,N_1786,N_3501);
and U6325 (N_6325,N_118,N_4561);
xnor U6326 (N_6326,N_2125,N_443);
or U6327 (N_6327,N_2333,N_2861);
and U6328 (N_6328,N_1950,N_3096);
xor U6329 (N_6329,N_2385,N_3321);
nor U6330 (N_6330,N_1970,N_2464);
nor U6331 (N_6331,N_168,N_803);
or U6332 (N_6332,N_1430,N_3115);
or U6333 (N_6333,N_4296,N_2536);
and U6334 (N_6334,N_54,N_66);
nand U6335 (N_6335,N_3323,N_769);
xor U6336 (N_6336,N_3069,N_4458);
nor U6337 (N_6337,N_2173,N_4806);
xnor U6338 (N_6338,N_3103,N_4474);
xnor U6339 (N_6339,N_4589,N_1448);
and U6340 (N_6340,N_3632,N_2911);
nor U6341 (N_6341,N_4096,N_2432);
and U6342 (N_6342,N_3494,N_3546);
and U6343 (N_6343,N_939,N_20);
xnor U6344 (N_6344,N_2369,N_1183);
nor U6345 (N_6345,N_636,N_1499);
or U6346 (N_6346,N_3094,N_4951);
nand U6347 (N_6347,N_3192,N_4825);
nor U6348 (N_6348,N_236,N_875);
nor U6349 (N_6349,N_1654,N_903);
and U6350 (N_6350,N_1416,N_1397);
xor U6351 (N_6351,N_3176,N_2678);
xor U6352 (N_6352,N_2504,N_3547);
and U6353 (N_6353,N_2901,N_1272);
and U6354 (N_6354,N_2832,N_1366);
nand U6355 (N_6355,N_3647,N_4537);
and U6356 (N_6356,N_1436,N_2787);
nand U6357 (N_6357,N_884,N_4726);
or U6358 (N_6358,N_1883,N_1626);
or U6359 (N_6359,N_4373,N_2028);
xnor U6360 (N_6360,N_2002,N_2376);
and U6361 (N_6361,N_943,N_2329);
xor U6362 (N_6362,N_2185,N_3932);
nor U6363 (N_6363,N_717,N_2715);
nor U6364 (N_6364,N_3017,N_4780);
nor U6365 (N_6365,N_67,N_584);
or U6366 (N_6366,N_3125,N_3810);
nand U6367 (N_6367,N_842,N_1478);
and U6368 (N_6368,N_2987,N_213);
or U6369 (N_6369,N_3144,N_1825);
nand U6370 (N_6370,N_954,N_1208);
nor U6371 (N_6371,N_4896,N_4609);
xnor U6372 (N_6372,N_2754,N_4962);
or U6373 (N_6373,N_4160,N_2255);
nor U6374 (N_6374,N_3340,N_1053);
nor U6375 (N_6375,N_3958,N_1094);
or U6376 (N_6376,N_493,N_528);
nor U6377 (N_6377,N_1544,N_4111);
and U6378 (N_6378,N_562,N_3449);
or U6379 (N_6379,N_4097,N_1106);
or U6380 (N_6380,N_2010,N_624);
xor U6381 (N_6381,N_4469,N_2435);
nand U6382 (N_6382,N_1119,N_4740);
nand U6383 (N_6383,N_1138,N_3202);
or U6384 (N_6384,N_639,N_4707);
or U6385 (N_6385,N_2311,N_1695);
and U6386 (N_6386,N_2681,N_3889);
xnor U6387 (N_6387,N_1317,N_4802);
nor U6388 (N_6388,N_658,N_2107);
nand U6389 (N_6389,N_456,N_1994);
nor U6390 (N_6390,N_1313,N_1459);
xor U6391 (N_6391,N_3386,N_1677);
xnor U6392 (N_6392,N_4972,N_4777);
and U6393 (N_6393,N_827,N_4500);
and U6394 (N_6394,N_2799,N_270);
xnor U6395 (N_6395,N_316,N_4796);
or U6396 (N_6396,N_2700,N_188);
or U6397 (N_6397,N_874,N_3333);
xnor U6398 (N_6398,N_2780,N_16);
and U6399 (N_6399,N_742,N_346);
and U6400 (N_6400,N_2040,N_4594);
nand U6401 (N_6401,N_4694,N_2275);
nor U6402 (N_6402,N_873,N_4807);
xnor U6403 (N_6403,N_2501,N_743);
nor U6404 (N_6404,N_2619,N_2586);
xor U6405 (N_6405,N_4772,N_4508);
and U6406 (N_6406,N_2259,N_1790);
and U6407 (N_6407,N_4676,N_2732);
and U6408 (N_6408,N_4232,N_2252);
nand U6409 (N_6409,N_1502,N_3733);
nor U6410 (N_6410,N_2061,N_3742);
xnor U6411 (N_6411,N_284,N_2170);
nand U6412 (N_6412,N_1214,N_77);
nand U6413 (N_6413,N_4948,N_3624);
nand U6414 (N_6414,N_3805,N_953);
xnor U6415 (N_6415,N_448,N_2262);
nor U6416 (N_6416,N_2961,N_136);
xor U6417 (N_6417,N_1745,N_407);
or U6418 (N_6418,N_107,N_1291);
or U6419 (N_6419,N_1958,N_3060);
nand U6420 (N_6420,N_44,N_3849);
nor U6421 (N_6421,N_4727,N_3769);
xor U6422 (N_6422,N_3685,N_4851);
xor U6423 (N_6423,N_2777,N_3978);
or U6424 (N_6424,N_4526,N_1420);
nor U6425 (N_6425,N_1076,N_720);
nand U6426 (N_6426,N_424,N_345);
and U6427 (N_6427,N_4956,N_3317);
xor U6428 (N_6428,N_3917,N_3629);
and U6429 (N_6429,N_4165,N_514);
nand U6430 (N_6430,N_729,N_2750);
or U6431 (N_6431,N_138,N_3936);
xor U6432 (N_6432,N_3143,N_3123);
xnor U6433 (N_6433,N_4112,N_3095);
nor U6434 (N_6434,N_342,N_2591);
and U6435 (N_6435,N_4021,N_1698);
and U6436 (N_6436,N_3642,N_4259);
or U6437 (N_6437,N_615,N_2669);
and U6438 (N_6438,N_799,N_981);
and U6439 (N_6439,N_4023,N_25);
and U6440 (N_6440,N_985,N_2566);
and U6441 (N_6441,N_3022,N_850);
and U6442 (N_6442,N_2379,N_447);
xnor U6443 (N_6443,N_2881,N_169);
nand U6444 (N_6444,N_3834,N_3933);
nand U6445 (N_6445,N_750,N_1857);
nor U6446 (N_6446,N_1492,N_550);
and U6447 (N_6447,N_3851,N_1226);
or U6448 (N_6448,N_1238,N_204);
nor U6449 (N_6449,N_4894,N_951);
nor U6450 (N_6450,N_4477,N_3398);
nor U6451 (N_6451,N_1299,N_2172);
xnor U6452 (N_6452,N_626,N_3582);
nand U6453 (N_6453,N_2000,N_3643);
and U6454 (N_6454,N_3269,N_2557);
or U6455 (N_6455,N_731,N_293);
nand U6456 (N_6456,N_3591,N_2579);
nor U6457 (N_6457,N_673,N_702);
or U6458 (N_6458,N_1772,N_2057);
nand U6459 (N_6459,N_161,N_553);
nor U6460 (N_6460,N_4621,N_2652);
xor U6461 (N_6461,N_3786,N_2569);
nand U6462 (N_6462,N_2215,N_2761);
or U6463 (N_6463,N_1872,N_2317);
xnor U6464 (N_6464,N_3554,N_3985);
nand U6465 (N_6465,N_3081,N_1399);
nor U6466 (N_6466,N_1061,N_4119);
xnor U6467 (N_6467,N_4172,N_86);
nand U6468 (N_6468,N_366,N_3891);
xor U6469 (N_6469,N_4466,N_1040);
nor U6470 (N_6470,N_3576,N_4242);
or U6471 (N_6471,N_1372,N_343);
xnor U6472 (N_6472,N_4752,N_489);
nand U6473 (N_6473,N_2890,N_205);
xnor U6474 (N_6474,N_4145,N_2993);
and U6475 (N_6475,N_1545,N_217);
nand U6476 (N_6476,N_4883,N_3832);
xor U6477 (N_6477,N_1649,N_4750);
and U6478 (N_6478,N_1424,N_4436);
xor U6479 (N_6479,N_1339,N_4672);
and U6480 (N_6480,N_779,N_85);
xor U6481 (N_6481,N_4791,N_2590);
or U6482 (N_6482,N_2297,N_2746);
nand U6483 (N_6483,N_1898,N_4106);
nor U6484 (N_6484,N_2353,N_2410);
xnor U6485 (N_6485,N_1371,N_1174);
nand U6486 (N_6486,N_2673,N_4043);
xnor U6487 (N_6487,N_3454,N_2046);
nand U6488 (N_6488,N_4862,N_149);
xnor U6489 (N_6489,N_3092,N_3767);
and U6490 (N_6490,N_3090,N_3422);
nor U6491 (N_6491,N_6,N_182);
xor U6492 (N_6492,N_7,N_2824);
and U6493 (N_6493,N_2984,N_4029);
and U6494 (N_6494,N_1719,N_373);
xnor U6495 (N_6495,N_4056,N_1511);
xnor U6496 (N_6496,N_1952,N_3485);
xor U6497 (N_6497,N_4380,N_4104);
nor U6498 (N_6498,N_1142,N_4000);
and U6499 (N_6499,N_3855,N_730);
and U6500 (N_6500,N_1277,N_2882);
nand U6501 (N_6501,N_4998,N_4643);
xnor U6502 (N_6502,N_2304,N_2453);
xor U6503 (N_6503,N_2483,N_3611);
nor U6504 (N_6504,N_2835,N_3132);
xnor U6505 (N_6505,N_1495,N_2708);
or U6506 (N_6506,N_4598,N_2526);
nor U6507 (N_6507,N_4847,N_1709);
and U6508 (N_6508,N_4570,N_390);
nor U6509 (N_6509,N_3186,N_1801);
nor U6510 (N_6510,N_4487,N_672);
or U6511 (N_6511,N_90,N_3961);
or U6512 (N_6512,N_4645,N_2948);
nor U6513 (N_6513,N_1928,N_1829);
or U6514 (N_6514,N_153,N_43);
or U6515 (N_6515,N_3831,N_4765);
xnor U6516 (N_6516,N_1908,N_4456);
or U6517 (N_6517,N_4798,N_3396);
xnor U6518 (N_6518,N_165,N_3497);
or U6519 (N_6519,N_3461,N_1836);
nand U6520 (N_6520,N_952,N_2360);
nand U6521 (N_6521,N_4110,N_4731);
nor U6522 (N_6522,N_2945,N_2603);
nor U6523 (N_6523,N_3201,N_3106);
nand U6524 (N_6524,N_1667,N_2188);
xor U6525 (N_6525,N_4792,N_3478);
and U6526 (N_6526,N_133,N_1634);
xnor U6527 (N_6527,N_3719,N_2194);
nor U6528 (N_6528,N_475,N_3);
or U6529 (N_6529,N_2704,N_1022);
nor U6530 (N_6530,N_62,N_3471);
nor U6531 (N_6531,N_2117,N_830);
nor U6532 (N_6532,N_1702,N_1619);
xnor U6533 (N_6533,N_1617,N_914);
and U6534 (N_6534,N_1648,N_3757);
nor U6535 (N_6535,N_4935,N_2688);
or U6536 (N_6536,N_2915,N_3142);
and U6537 (N_6537,N_4997,N_680);
or U6538 (N_6538,N_440,N_4322);
and U6539 (N_6539,N_3018,N_1636);
xor U6540 (N_6540,N_4563,N_1281);
and U6541 (N_6541,N_3465,N_1400);
nor U6542 (N_6542,N_3006,N_3552);
or U6543 (N_6543,N_4133,N_1006);
xnor U6544 (N_6544,N_739,N_4);
or U6545 (N_6545,N_829,N_2555);
and U6546 (N_6546,N_4386,N_3466);
nand U6547 (N_6547,N_2520,N_1943);
nor U6548 (N_6548,N_4899,N_2857);
and U6549 (N_6549,N_520,N_1066);
or U6550 (N_6550,N_2734,N_648);
nand U6551 (N_6551,N_1881,N_1917);
nor U6552 (N_6552,N_2928,N_4839);
or U6553 (N_6553,N_4120,N_2870);
xnor U6554 (N_6554,N_52,N_2741);
and U6555 (N_6555,N_2380,N_4343);
nand U6556 (N_6556,N_1103,N_2986);
and U6557 (N_6557,N_4265,N_4647);
xnor U6558 (N_6558,N_3436,N_454);
and U6559 (N_6559,N_1914,N_4683);
and U6560 (N_6560,N_3761,N_2090);
or U6561 (N_6561,N_3571,N_824);
nand U6562 (N_6562,N_3038,N_3162);
nor U6563 (N_6563,N_1232,N_3303);
nand U6564 (N_6564,N_2804,N_1075);
or U6565 (N_6565,N_944,N_1203);
and U6566 (N_6566,N_3762,N_389);
or U6567 (N_6567,N_191,N_1364);
nor U6568 (N_6568,N_2588,N_3282);
and U6569 (N_6569,N_4656,N_1231);
or U6570 (N_6570,N_1064,N_3199);
or U6571 (N_6571,N_607,N_3750);
nand U6572 (N_6572,N_2195,N_1693);
nor U6573 (N_6573,N_4994,N_1280);
xor U6574 (N_6574,N_409,N_1781);
or U6575 (N_6575,N_50,N_3037);
nor U6576 (N_6576,N_4229,N_2433);
and U6577 (N_6577,N_3882,N_2390);
nand U6578 (N_6578,N_3412,N_1167);
nand U6579 (N_6579,N_450,N_4992);
or U6580 (N_6580,N_3395,N_2503);
xor U6581 (N_6581,N_4098,N_1084);
nor U6582 (N_6582,N_1931,N_4774);
nor U6583 (N_6583,N_4944,N_3500);
or U6584 (N_6584,N_4562,N_3559);
nand U6585 (N_6585,N_934,N_4527);
nor U6586 (N_6586,N_324,N_4766);
nor U6587 (N_6587,N_3093,N_3743);
xnor U6588 (N_6588,N_1427,N_2910);
nand U6589 (N_6589,N_2371,N_775);
or U6590 (N_6590,N_4557,N_2179);
and U6591 (N_6591,N_1602,N_3564);
nor U6592 (N_6592,N_2558,N_436);
nor U6593 (N_6593,N_683,N_4991);
or U6594 (N_6594,N_4480,N_1178);
or U6595 (N_6595,N_974,N_1388);
xor U6596 (N_6596,N_2047,N_761);
or U6597 (N_6597,N_3867,N_1292);
nand U6598 (N_6598,N_4077,N_3214);
and U6599 (N_6599,N_4134,N_965);
nor U6600 (N_6600,N_37,N_4934);
nand U6601 (N_6601,N_3070,N_1275);
nand U6602 (N_6602,N_1632,N_2597);
xor U6603 (N_6603,N_3351,N_686);
xnor U6604 (N_6604,N_603,N_4556);
nand U6605 (N_6605,N_4051,N_4522);
and U6606 (N_6606,N_333,N_2817);
nor U6607 (N_6607,N_3983,N_84);
xor U6608 (N_6608,N_3031,N_1554);
and U6609 (N_6609,N_157,N_2178);
nor U6610 (N_6610,N_2745,N_2951);
nand U6611 (N_6611,N_1821,N_4869);
nand U6612 (N_6612,N_4203,N_740);
xor U6613 (N_6613,N_1852,N_2876);
nor U6614 (N_6614,N_3704,N_3034);
and U6615 (N_6615,N_34,N_1008);
xnor U6616 (N_6616,N_4779,N_1823);
xnor U6617 (N_6617,N_3636,N_2903);
xor U6618 (N_6618,N_1220,N_3289);
and U6619 (N_6619,N_994,N_437);
nor U6620 (N_6620,N_4743,N_4218);
nor U6621 (N_6621,N_661,N_1849);
xor U6622 (N_6622,N_2132,N_375);
xnor U6623 (N_6623,N_1537,N_1913);
or U6624 (N_6624,N_3813,N_2187);
xor U6625 (N_6625,N_51,N_1594);
or U6626 (N_6626,N_4749,N_2576);
nand U6627 (N_6627,N_1674,N_365);
nor U6628 (N_6628,N_1070,N_3447);
nand U6629 (N_6629,N_4885,N_977);
and U6630 (N_6630,N_4497,N_4402);
xnor U6631 (N_6631,N_2647,N_888);
and U6632 (N_6632,N_2560,N_4461);
nand U6633 (N_6633,N_3668,N_1689);
or U6634 (N_6634,N_3026,N_3545);
or U6635 (N_6635,N_2687,N_1576);
or U6636 (N_6636,N_4524,N_3663);
xnor U6637 (N_6637,N_3895,N_1199);
nor U6638 (N_6638,N_4858,N_3646);
xor U6639 (N_6639,N_18,N_805);
xor U6640 (N_6640,N_1683,N_4222);
nand U6641 (N_6641,N_3993,N_692);
nor U6642 (N_6642,N_2843,N_3696);
nand U6643 (N_6643,N_3620,N_1074);
nand U6644 (N_6644,N_3062,N_449);
or U6645 (N_6645,N_4156,N_3286);
nand U6646 (N_6646,N_4822,N_3372);
xnor U6647 (N_6647,N_2666,N_1921);
or U6648 (N_6648,N_3036,N_184);
and U6649 (N_6649,N_2541,N_3965);
xor U6650 (N_6650,N_3088,N_337);
nor U6651 (N_6651,N_3997,N_1311);
or U6652 (N_6652,N_3724,N_3584);
and U6653 (N_6653,N_727,N_2240);
or U6654 (N_6654,N_2680,N_641);
and U6655 (N_6655,N_4316,N_3182);
nor U6656 (N_6656,N_3030,N_3033);
or U6657 (N_6657,N_532,N_4324);
nand U6658 (N_6658,N_4532,N_4697);
nor U6659 (N_6659,N_1134,N_4573);
nor U6660 (N_6660,N_4670,N_3687);
and U6661 (N_6661,N_2216,N_3732);
and U6662 (N_6662,N_543,N_4079);
and U6663 (N_6663,N_4277,N_2206);
nand U6664 (N_6664,N_406,N_3654);
or U6665 (N_6665,N_2023,N_4633);
xor U6666 (N_6666,N_1414,N_2041);
and U6667 (N_6667,N_969,N_1680);
and U6668 (N_6668,N_4782,N_1525);
or U6669 (N_6669,N_3866,N_599);
nor U6670 (N_6670,N_3319,N_0);
nor U6671 (N_6671,N_292,N_2500);
nor U6672 (N_6672,N_738,N_48);
or U6673 (N_6673,N_858,N_3859);
nand U6674 (N_6674,N_127,N_3246);
nand U6675 (N_6675,N_2913,N_3715);
nand U6676 (N_6676,N_4678,N_3977);
or U6677 (N_6677,N_946,N_187);
nor U6678 (N_6678,N_1749,N_1489);
nor U6679 (N_6679,N_1760,N_1270);
nand U6680 (N_6680,N_1737,N_2788);
and U6681 (N_6681,N_3435,N_1992);
or U6682 (N_6682,N_928,N_1717);
nand U6683 (N_6683,N_1768,N_1360);
nor U6684 (N_6684,N_1907,N_1173);
or U6685 (N_6685,N_1670,N_4166);
xnor U6686 (N_6686,N_1587,N_2613);
nand U6687 (N_6687,N_3016,N_190);
and U6688 (N_6688,N_1157,N_2286);
or U6689 (N_6689,N_1727,N_911);
or U6690 (N_6690,N_2848,N_4577);
nand U6691 (N_6691,N_3828,N_3119);
xnor U6692 (N_6692,N_109,N_63);
xnor U6693 (N_6693,N_3079,N_778);
and U6694 (N_6694,N_110,N_2022);
or U6695 (N_6695,N_2610,N_1962);
xnor U6696 (N_6696,N_1122,N_3639);
or U6697 (N_6697,N_1129,N_244);
xor U6698 (N_6698,N_1774,N_1615);
and U6699 (N_6699,N_4354,N_1315);
nor U6700 (N_6700,N_203,N_1777);
or U6701 (N_6701,N_486,N_1631);
nor U6702 (N_6702,N_1503,N_1767);
xor U6703 (N_6703,N_282,N_5);
nand U6704 (N_6704,N_3204,N_4635);
and U6705 (N_6705,N_2442,N_2684);
and U6706 (N_6706,N_243,N_2294);
xnor U6707 (N_6707,N_1114,N_4033);
xnor U6708 (N_6708,N_4587,N_306);
or U6709 (N_6709,N_4216,N_1419);
or U6710 (N_6710,N_1642,N_185);
nand U6711 (N_6711,N_2892,N_1555);
nor U6712 (N_6712,N_425,N_2830);
xnor U6713 (N_6713,N_987,N_477);
nand U6714 (N_6714,N_4308,N_3242);
and U6715 (N_6715,N_2658,N_2078);
or U6716 (N_6716,N_3519,N_1109);
and U6717 (N_6717,N_979,N_4117);
xnor U6718 (N_6718,N_1863,N_1651);
xor U6719 (N_6719,N_632,N_3490);
xnor U6720 (N_6720,N_1266,N_3067);
and U6721 (N_6721,N_166,N_2207);
nor U6722 (N_6722,N_4030,N_783);
and U6723 (N_6723,N_2966,N_3586);
nor U6724 (N_6724,N_220,N_4344);
xnor U6725 (N_6725,N_1584,N_4330);
nand U6726 (N_6726,N_848,N_4873);
and U6727 (N_6727,N_2278,N_3727);
nor U6728 (N_6728,N_4310,N_4014);
and U6729 (N_6729,N_1467,N_2919);
or U6730 (N_6730,N_338,N_4548);
or U6731 (N_6731,N_2770,N_2467);
nor U6732 (N_6732,N_513,N_3514);
or U6733 (N_6733,N_627,N_3871);
and U6734 (N_6734,N_1579,N_4377);
and U6735 (N_6735,N_1346,N_2279);
nand U6736 (N_6736,N_1349,N_105);
nand U6737 (N_6737,N_577,N_4137);
xnor U6738 (N_6738,N_4092,N_1532);
nor U6739 (N_6739,N_2542,N_3502);
xnor U6740 (N_6740,N_2245,N_2056);
xor U6741 (N_6741,N_4925,N_1671);
and U6742 (N_6742,N_1840,N_4439);
nor U6743 (N_6743,N_4428,N_2113);
nand U6744 (N_6744,N_3311,N_949);
nand U6745 (N_6745,N_3593,N_3193);
nand U6746 (N_6746,N_617,N_3136);
nor U6747 (N_6747,N_129,N_554);
nor U6748 (N_6748,N_2705,N_2794);
or U6749 (N_6749,N_1678,N_771);
xor U6750 (N_6750,N_2800,N_570);
nor U6751 (N_6751,N_1515,N_3536);
and U6752 (N_6752,N_2562,N_3203);
nand U6753 (N_6753,N_3091,N_2827);
or U6754 (N_6754,N_262,N_2936);
xor U6755 (N_6755,N_4624,N_4468);
or U6756 (N_6756,N_923,N_160);
nor U6757 (N_6757,N_1775,N_2895);
xor U6758 (N_6758,N_69,N_397);
nor U6759 (N_6759,N_3806,N_3265);
nor U6760 (N_6760,N_1574,N_3610);
and U6761 (N_6761,N_3266,N_3923);
xor U6762 (N_6762,N_3971,N_895);
xnor U6763 (N_6763,N_2338,N_71);
or U6764 (N_6764,N_3518,N_3013);
nor U6765 (N_6765,N_310,N_1788);
or U6766 (N_6766,N_4132,N_4870);
xor U6767 (N_6767,N_613,N_2550);
nor U6768 (N_6768,N_1725,N_4990);
nand U6769 (N_6769,N_3462,N_2935);
xnor U6770 (N_6770,N_1524,N_1710);
xnor U6771 (N_6771,N_1800,N_4176);
nor U6772 (N_6772,N_3804,N_3309);
and U6773 (N_6773,N_530,N_4711);
and U6774 (N_6774,N_1017,N_2475);
nor U6775 (N_6775,N_1393,N_2740);
or U6776 (N_6776,N_4147,N_4753);
nor U6777 (N_6777,N_2081,N_3080);
nand U6778 (N_6778,N_3574,N_4493);
or U6779 (N_6779,N_3503,N_4821);
xnor U6780 (N_6780,N_3601,N_582);
nand U6781 (N_6781,N_321,N_363);
and U6782 (N_6782,N_3951,N_4859);
nor U6783 (N_6783,N_4307,N_9);
nor U6784 (N_6784,N_237,N_2840);
nor U6785 (N_6785,N_426,N_3561);
or U6786 (N_6786,N_3307,N_1202);
and U6787 (N_6787,N_2242,N_3491);
nor U6788 (N_6788,N_957,N_3972);
nand U6789 (N_6789,N_329,N_2766);
or U6790 (N_6790,N_555,N_150);
xnor U6791 (N_6791,N_4251,N_377);
or U6792 (N_6792,N_3403,N_2667);
or U6793 (N_6793,N_3005,N_2254);
and U6794 (N_6794,N_2729,N_1452);
and U6795 (N_6795,N_1175,N_2905);
or U6796 (N_6796,N_2361,N_2595);
nand U6797 (N_6797,N_1410,N_385);
xnor U6798 (N_6798,N_2264,N_2498);
and U6799 (N_6799,N_4722,N_2642);
and U6800 (N_6800,N_1197,N_3365);
nor U6801 (N_6801,N_1113,N_121);
xnor U6802 (N_6802,N_2008,N_3250);
and U6803 (N_6803,N_4838,N_1860);
xor U6804 (N_6804,N_278,N_1625);
nand U6805 (N_6805,N_277,N_3281);
xor U6806 (N_6806,N_4712,N_2592);
or U6807 (N_6807,N_4017,N_257);
nor U6808 (N_6808,N_754,N_3329);
nor U6809 (N_6809,N_4412,N_4575);
or U6810 (N_6810,N_1260,N_2496);
or U6811 (N_6811,N_73,N_3887);
nand U6812 (N_6812,N_4169,N_2522);
xnor U6813 (N_6813,N_4835,N_4135);
nor U6814 (N_6814,N_1542,N_1948);
and U6815 (N_6815,N_3254,N_3763);
or U6816 (N_6816,N_2559,N_2581);
nor U6817 (N_6817,N_1479,N_1165);
nor U6818 (N_6818,N_1607,N_2862);
nor U6819 (N_6819,N_2308,N_3679);
nand U6820 (N_6820,N_4658,N_4820);
xor U6821 (N_6821,N_3540,N_2052);
and U6822 (N_6822,N_3027,N_2469);
nand U6823 (N_6823,N_3623,N_1813);
or U6824 (N_6824,N_3689,N_1797);
or U6825 (N_6825,N_4100,N_4730);
or U6826 (N_6826,N_3688,N_2852);
nor U6827 (N_6827,N_1351,N_3517);
nor U6828 (N_6828,N_4427,N_2232);
nor U6829 (N_6829,N_4709,N_1755);
nor U6830 (N_6830,N_3777,N_735);
xor U6831 (N_6831,N_1285,N_1472);
and U6832 (N_6832,N_1415,N_3117);
or U6833 (N_6833,N_3946,N_4797);
nor U6834 (N_6834,N_1184,N_498);
nand U6835 (N_6835,N_4376,N_148);
xor U6836 (N_6836,N_2227,N_3275);
or U6837 (N_6837,N_968,N_379);
nand U6838 (N_6838,N_1384,N_1982);
nor U6839 (N_6839,N_3074,N_560);
and U6840 (N_6840,N_3120,N_898);
nand U6841 (N_6841,N_2429,N_3590);
xnor U6842 (N_6842,N_3837,N_700);
and U6843 (N_6843,N_4273,N_1747);
and U6844 (N_6844,N_2596,N_3568);
nor U6845 (N_6845,N_2643,N_2296);
or U6846 (N_6846,N_2657,N_867);
or U6847 (N_6847,N_4592,N_3206);
nand U6848 (N_6848,N_4542,N_1083);
nand U6849 (N_6849,N_733,N_1887);
and U6850 (N_6850,N_1012,N_4179);
nor U6851 (N_6851,N_666,N_732);
or U6852 (N_6852,N_1265,N_4236);
nand U6853 (N_6853,N_790,N_3713);
or U6854 (N_6854,N_4671,N_4064);
or U6855 (N_6855,N_2450,N_3549);
nor U6856 (N_6856,N_291,N_840);
and U6857 (N_6857,N_4248,N_1754);
nand U6858 (N_6858,N_4010,N_348);
nand U6859 (N_6859,N_1091,N_2174);
or U6860 (N_6860,N_501,N_1899);
nor U6861 (N_6861,N_2277,N_1639);
nor U6862 (N_6862,N_2212,N_1396);
xnor U6863 (N_6863,N_1946,N_2941);
nand U6864 (N_6864,N_503,N_2580);
or U6865 (N_6865,N_3393,N_3021);
nand U6866 (N_6866,N_4329,N_1494);
nand U6867 (N_6867,N_3898,N_677);
and U6868 (N_6868,N_2571,N_4814);
xor U6869 (N_6869,N_300,N_3171);
and U6870 (N_6870,N_2577,N_2176);
and U6871 (N_6871,N_2860,N_211);
and U6872 (N_6872,N_3346,N_3735);
xor U6873 (N_6873,N_1363,N_3846);
and U6874 (N_6874,N_2233,N_2838);
nor U6875 (N_6875,N_2150,N_4987);
xnor U6876 (N_6876,N_4572,N_937);
nor U6877 (N_6877,N_3349,N_629);
or U6878 (N_6878,N_2842,N_1748);
xnor U6879 (N_6879,N_1637,N_471);
nor U6880 (N_6880,N_4355,N_3380);
or U6881 (N_6881,N_3440,N_4411);
or U6882 (N_6882,N_4495,N_1588);
xor U6883 (N_6883,N_3477,N_970);
nor U6884 (N_6884,N_1222,N_3630);
nor U6885 (N_6885,N_4246,N_2664);
and U6886 (N_6886,N_2885,N_2894);
xor U6887 (N_6887,N_2809,N_111);
nor U6888 (N_6888,N_896,N_3450);
and U6889 (N_6889,N_3817,N_3430);
nand U6890 (N_6890,N_1652,N_258);
nor U6891 (N_6891,N_2623,N_2717);
nor U6892 (N_6892,N_3829,N_4252);
and U6893 (N_6893,N_1897,N_3775);
nand U6894 (N_6894,N_2283,N_4931);
and U6895 (N_6895,N_3749,N_2821);
and U6896 (N_6896,N_1795,N_793);
nand U6897 (N_6897,N_4275,N_802);
xnor U6898 (N_6898,N_2157,N_4485);
and U6899 (N_6899,N_39,N_2244);
or U6900 (N_6900,N_1949,N_4975);
and U6901 (N_6901,N_3868,N_3163);
xnor U6902 (N_6902,N_4758,N_3355);
or U6903 (N_6903,N_2070,N_1342);
and U6904 (N_6904,N_3389,N_1462);
and U6905 (N_6905,N_1888,N_3682);
or U6906 (N_6906,N_1809,N_1441);
and U6907 (N_6907,N_2257,N_529);
and U6908 (N_6908,N_1776,N_2940);
xor U6909 (N_6909,N_2326,N_3709);
or U6910 (N_6910,N_114,N_3657);
and U6911 (N_6911,N_274,N_3791);
nor U6912 (N_6912,N_61,N_2974);
nand U6913 (N_6913,N_2925,N_487);
or U6914 (N_6914,N_868,N_21);
and U6915 (N_6915,N_2632,N_2144);
xor U6916 (N_6916,N_1815,N_2968);
or U6917 (N_6917,N_1612,N_3725);
or U6918 (N_6918,N_4544,N_4602);
and U6919 (N_6919,N_3291,N_53);
xor U6920 (N_6920,N_2489,N_2131);
xor U6921 (N_6921,N_705,N_4269);
xor U6922 (N_6922,N_2606,N_3432);
nand U6923 (N_6923,N_1072,N_1168);
nand U6924 (N_6924,N_935,N_1195);
xor U6925 (N_6925,N_4688,N_4204);
nand U6926 (N_6926,N_1107,N_218);
xnor U6927 (N_6927,N_1572,N_1789);
and U6928 (N_6928,N_597,N_4230);
nand U6929 (N_6929,N_4747,N_253);
or U6930 (N_6930,N_507,N_4254);
nand U6931 (N_6931,N_4986,N_4404);
nor U6932 (N_6932,N_4569,N_936);
nor U6933 (N_6933,N_1802,N_2568);
and U6934 (N_6934,N_152,N_4580);
nor U6935 (N_6935,N_744,N_4057);
nand U6936 (N_6936,N_759,N_834);
or U6937 (N_6937,N_4942,N_3649);
nand U6938 (N_6938,N_1306,N_4306);
nor U6939 (N_6939,N_3305,N_1556);
xnor U6940 (N_6940,N_882,N_3969);
xnor U6941 (N_6941,N_2263,N_4025);
nor U6942 (N_6942,N_347,N_1942);
and U6943 (N_6943,N_2930,N_4282);
nand U6944 (N_6944,N_2129,N_3257);
xor U6945 (N_6945,N_973,N_4826);
nand U6946 (N_6946,N_4541,N_1146);
nor U6947 (N_6947,N_4312,N_2738);
nor U6948 (N_6948,N_4696,N_445);
nor U6949 (N_6949,N_2,N_2455);
xor U6950 (N_6950,N_473,N_1575);
nand U6951 (N_6951,N_2533,N_4028);
xnor U6952 (N_6952,N_4529,N_2651);
xnor U6953 (N_6953,N_488,N_3802);
or U6954 (N_6954,N_878,N_846);
and U6955 (N_6955,N_3221,N_1918);
and U6956 (N_6956,N_1647,N_45);
and U6957 (N_6957,N_4291,N_2702);
xnor U6958 (N_6958,N_4890,N_4501);
nand U6959 (N_6959,N_2472,N_2300);
xnor U6960 (N_6960,N_3722,N_3024);
xnor U6961 (N_6961,N_1321,N_1417);
and U6962 (N_6962,N_4003,N_1509);
nand U6963 (N_6963,N_2146,N_1041);
xor U6964 (N_6964,N_2582,N_135);
or U6965 (N_6965,N_1724,N_4385);
or U6966 (N_6966,N_2864,N_524);
and U6967 (N_6967,N_23,N_4793);
nand U6968 (N_6968,N_2927,N_4984);
nor U6969 (N_6969,N_4813,N_1004);
nand U6970 (N_6970,N_2267,N_2461);
nor U6971 (N_6971,N_3428,N_4186);
nand U6972 (N_6972,N_3516,N_3354);
xor U6973 (N_6973,N_1487,N_1296);
xnor U6974 (N_6974,N_688,N_1402);
and U6975 (N_6975,N_2617,N_3165);
nand U6976 (N_6976,N_4208,N_1868);
nor U6977 (N_6977,N_825,N_36);
nand U6978 (N_6978,N_3359,N_194);
and U6979 (N_6979,N_2312,N_4403);
xnor U6980 (N_6980,N_2869,N_2699);
nand U6981 (N_6981,N_4276,N_3400);
nand U6982 (N_6982,N_3684,N_904);
nor U6983 (N_6983,N_4963,N_4161);
xor U6984 (N_6984,N_1376,N_1359);
nor U6985 (N_6985,N_869,N_3375);
or U6986 (N_6986,N_1020,N_3587);
xor U6987 (N_6987,N_2192,N_3736);
and U6988 (N_6988,N_4026,N_3446);
or U6989 (N_6989,N_2828,N_4698);
nand U6990 (N_6990,N_3316,N_1975);
nand U6991 (N_6991,N_1243,N_226);
nand U6992 (N_6992,N_227,N_200);
nor U6993 (N_6993,N_2773,N_782);
nand U6994 (N_6994,N_657,N_1181);
and U6995 (N_6995,N_3706,N_4289);
and U6996 (N_6996,N_3071,N_3072);
nand U6997 (N_6997,N_1513,N_2025);
nand U6998 (N_6998,N_1660,N_4744);
or U6999 (N_6999,N_3232,N_2007);
or U7000 (N_7000,N_1981,N_4457);
xnor U7001 (N_7001,N_4049,N_3698);
nand U7002 (N_7002,N_3236,N_2618);
or U7003 (N_7003,N_380,N_2627);
nor U7004 (N_7004,N_1547,N_3982);
nand U7005 (N_7005,N_2316,N_3241);
nand U7006 (N_7006,N_2810,N_3928);
and U7007 (N_7007,N_1429,N_3180);
or U7008 (N_7008,N_4410,N_2223);
and U7009 (N_7009,N_4319,N_4400);
nor U7010 (N_7010,N_1110,N_208);
or U7011 (N_7011,N_364,N_3420);
or U7012 (N_7012,N_3770,N_3076);
and U7013 (N_7013,N_2527,N_1029);
or U7014 (N_7014,N_3296,N_1604);
nor U7015 (N_7015,N_1501,N_1204);
nand U7016 (N_7016,N_4496,N_3787);
nand U7017 (N_7017,N_2427,N_3990);
and U7018 (N_7018,N_2716,N_163);
xnor U7019 (N_7019,N_3589,N_2349);
xnor U7020 (N_7020,N_2346,N_3558);
and U7021 (N_7021,N_4964,N_2243);
or U7022 (N_7022,N_4093,N_1259);
and U7023 (N_7023,N_772,N_4116);
xor U7024 (N_7024,N_3708,N_810);
or U7025 (N_7025,N_1526,N_4960);
nor U7026 (N_7026,N_4520,N_3937);
and U7027 (N_7027,N_2552,N_3438);
or U7028 (N_7028,N_3941,N_2004);
and U7029 (N_7029,N_4155,N_4719);
nand U7030 (N_7030,N_4613,N_2831);
nand U7031 (N_7031,N_1289,N_3607);
and U7032 (N_7032,N_1977,N_128);
nor U7033 (N_7033,N_1411,N_3581);
xnor U7034 (N_7034,N_752,N_374);
nor U7035 (N_7035,N_1577,N_1620);
or U7036 (N_7036,N_82,N_2013);
xor U7037 (N_7037,N_3173,N_4971);
nand U7038 (N_7038,N_2221,N_4915);
nand U7039 (N_7039,N_2213,N_591);
or U7040 (N_7040,N_619,N_4211);
nand U7041 (N_7041,N_3042,N_3507);
and U7042 (N_7042,N_1743,N_548);
nand U7043 (N_7043,N_2289,N_838);
nand U7044 (N_7044,N_4340,N_816);
nor U7045 (N_7045,N_1961,N_313);
and U7046 (N_7046,N_2271,N_3670);
and U7047 (N_7047,N_1248,N_835);
nand U7048 (N_7048,N_4078,N_3797);
nand U7049 (N_7049,N_1468,N_2709);
xnor U7050 (N_7050,N_3702,N_4325);
and U7051 (N_7051,N_231,N_287);
and U7052 (N_7052,N_286,N_3711);
nand U7053 (N_7053,N_517,N_4907);
xnor U7054 (N_7054,N_189,N_4260);
xnor U7055 (N_7055,N_1930,N_1910);
nand U7056 (N_7056,N_235,N_319);
and U7057 (N_7057,N_1205,N_3987);
and U7058 (N_7058,N_325,N_4662);
nand U7059 (N_7059,N_1766,N_4714);
and U7060 (N_7060,N_4193,N_2783);
xnor U7061 (N_7061,N_4108,N_4567);
and U7062 (N_7062,N_2480,N_2140);
xnor U7063 (N_7063,N_2485,N_921);
xnor U7064 (N_7064,N_654,N_4924);
xnor U7065 (N_7065,N_1983,N_833);
nand U7066 (N_7066,N_155,N_590);
or U7067 (N_7067,N_280,N_2995);
nand U7068 (N_7068,N_3697,N_451);
or U7069 (N_7069,N_2942,N_2404);
xor U7070 (N_7070,N_3414,N_327);
nand U7071 (N_7071,N_1684,N_3448);
or U7072 (N_7072,N_1926,N_4109);
and U7073 (N_7073,N_24,N_2625);
or U7074 (N_7074,N_3260,N_1003);
and U7075 (N_7075,N_1140,N_1028);
nor U7076 (N_7076,N_3397,N_126);
xor U7077 (N_7077,N_4874,N_2751);
and U7078 (N_7078,N_3638,N_791);
or U7079 (N_7079,N_2644,N_4872);
and U7080 (N_7080,N_1035,N_1242);
xor U7081 (N_7081,N_4022,N_2266);
nand U7082 (N_7082,N_3886,N_4634);
or U7083 (N_7083,N_3343,N_2502);
nor U7084 (N_7084,N_1561,N_521);
xnor U7085 (N_7085,N_1616,N_4309);
or U7086 (N_7086,N_2988,N_3243);
or U7087 (N_7087,N_4473,N_3764);
or U7088 (N_7088,N_2733,N_4560);
or U7089 (N_7089,N_3943,N_2871);
nor U7090 (N_7090,N_1120,N_2015);
xnor U7091 (N_7091,N_1446,N_3843);
nand U7092 (N_7092,N_3320,N_3844);
nand U7093 (N_7093,N_3167,N_4164);
and U7094 (N_7094,N_1449,N_4606);
or U7095 (N_7095,N_2511,N_1031);
nor U7096 (N_7096,N_3811,N_975);
or U7097 (N_7097,N_88,N_2757);
nor U7098 (N_7098,N_1087,N_3595);
nor U7099 (N_7099,N_1333,N_662);
nor U7100 (N_7100,N_130,N_2697);
nand U7101 (N_7101,N_1161,N_4206);
nor U7102 (N_7102,N_2230,N_2364);
nor U7103 (N_7103,N_4370,N_4488);
xor U7104 (N_7104,N_1267,N_3653);
and U7105 (N_7105,N_4047,N_3956);
xor U7106 (N_7106,N_4784,N_3352);
or U7107 (N_7107,N_893,N_3528);
nand U7108 (N_7108,N_3209,N_984);
nor U7109 (N_7109,N_2100,N_4072);
or U7110 (N_7110,N_2347,N_151);
and U7111 (N_7111,N_273,N_4950);
and U7112 (N_7112,N_2102,N_1005);
xor U7113 (N_7113,N_2321,N_3876);
nand U7114 (N_7114,N_2539,N_3147);
or U7115 (N_7115,N_3360,N_2234);
nor U7116 (N_7116,N_2017,N_4818);
and U7117 (N_7117,N_2138,N_1224);
and U7118 (N_7118,N_4447,N_843);
xor U7119 (N_7119,N_468,N_3592);
and U7120 (N_7120,N_1312,N_1032);
nor U7121 (N_7121,N_3962,N_4660);
and U7122 (N_7122,N_3527,N_4636);
and U7123 (N_7123,N_1176,N_3912);
nand U7124 (N_7124,N_2492,N_353);
or U7125 (N_7125,N_2430,N_3637);
or U7126 (N_7126,N_4884,N_4953);
and U7127 (N_7127,N_2677,N_1718);
xnor U7128 (N_7128,N_4016,N_4938);
and U7129 (N_7129,N_2459,N_2239);
nand U7130 (N_7130,N_2137,N_676);
or U7131 (N_7131,N_879,N_3627);
or U7132 (N_7132,N_4650,N_1904);
xor U7133 (N_7133,N_4648,N_264);
nor U7134 (N_7134,N_1957,N_1701);
and U7135 (N_7135,N_3328,N_4437);
nor U7136 (N_7136,N_1661,N_2356);
xor U7137 (N_7137,N_1757,N_87);
nor U7138 (N_7138,N_2611,N_2999);
nor U7139 (N_7139,N_2612,N_1136);
and U7140 (N_7140,N_2792,N_2141);
nand U7141 (N_7141,N_1807,N_958);
nor U7142 (N_7142,N_3014,N_1764);
nor U7143 (N_7143,N_2534,N_4454);
xnor U7144 (N_7144,N_4076,N_3009);
nor U7145 (N_7145,N_4914,N_281);
or U7146 (N_7146,N_159,N_4903);
or U7147 (N_7147,N_1081,N_3308);
xnor U7148 (N_7148,N_2050,N_992);
and U7149 (N_7149,N_4198,N_877);
nor U7150 (N_7150,N_2126,N_2898);
and U7151 (N_7151,N_4654,N_1951);
nand U7152 (N_7152,N_2282,N_4499);
and U7153 (N_7153,N_4554,N_998);
and U7154 (N_7154,N_1460,N_4004);
nor U7155 (N_7155,N_815,N_588);
and U7156 (N_7156,N_183,N_4405);
or U7157 (N_7157,N_1486,N_3049);
or U7158 (N_7158,N_41,N_557);
nor U7159 (N_7159,N_3631,N_3293);
xor U7160 (N_7160,N_1149,N_3105);
and U7161 (N_7161,N_1093,N_1347);
and U7162 (N_7162,N_663,N_3676);
nor U7163 (N_7163,N_4008,N_3902);
nor U7164 (N_7164,N_1628,N_862);
or U7165 (N_7165,N_2551,N_1252);
or U7166 (N_7166,N_341,N_762);
or U7167 (N_7167,N_3588,N_49);
and U7168 (N_7168,N_912,N_4066);
nor U7169 (N_7169,N_2374,N_1839);
xnor U7170 (N_7170,N_1465,N_3157);
nand U7171 (N_7171,N_4757,N_1233);
xor U7172 (N_7172,N_3216,N_2546);
nand U7173 (N_7173,N_459,N_3551);
or U7174 (N_7174,N_147,N_1997);
and U7175 (N_7175,N_3288,N_1235);
nor U7176 (N_7176,N_1409,N_246);
nor U7177 (N_7177,N_4123,N_2823);
xnor U7178 (N_7178,N_4988,N_4607);
nor U7179 (N_7179,N_4622,N_4301);
nor U7180 (N_7180,N_1583,N_1682);
nor U7181 (N_7181,N_4346,N_1843);
xnor U7182 (N_7182,N_2104,N_1476);
xnor U7183 (N_7183,N_470,N_2413);
or U7184 (N_7184,N_3957,N_2307);
and U7185 (N_7185,N_2474,N_4201);
nor U7186 (N_7186,N_2335,N_1796);
xor U7187 (N_7187,N_3872,N_3640);
xor U7188 (N_7188,N_1234,N_4830);
nand U7189 (N_7189,N_2274,N_1135);
or U7190 (N_7190,N_2846,N_3433);
nand U7191 (N_7191,N_4424,N_4188);
nand U7192 (N_7192,N_3594,N_723);
or U7193 (N_7193,N_4491,N_420);
and U7194 (N_7194,N_387,N_176);
or U7195 (N_7195,N_1439,N_4512);
nand U7196 (N_7196,N_102,N_224);
or U7197 (N_7197,N_2365,N_1357);
nand U7198 (N_7198,N_2064,N_2538);
nor U7199 (N_7199,N_3543,N_1945);
or U7200 (N_7200,N_706,N_4012);
nor U7201 (N_7201,N_3538,N_1201);
xnor U7202 (N_7202,N_1598,N_4595);
xnor U7203 (N_7203,N_4690,N_4713);
and U7204 (N_7204,N_3532,N_2879);
xor U7205 (N_7205,N_618,N_2045);
nor U7206 (N_7206,N_4173,N_764);
nor U7207 (N_7207,N_1209,N_4190);
or U7208 (N_7208,N_1610,N_2682);
nor U7209 (N_7209,N_2816,N_1341);
or U7210 (N_7210,N_2111,N_480);
nand U7211 (N_7211,N_3955,N_3740);
xnor U7212 (N_7212,N_3752,N_4628);
and U7213 (N_7213,N_2758,N_3661);
or U7214 (N_7214,N_2743,N_4032);
or U7215 (N_7215,N_2115,N_3841);
nand U7216 (N_7216,N_2811,N_2712);
and U7217 (N_7217,N_988,N_4558);
nand U7218 (N_7218,N_3146,N_1352);
nand U7219 (N_7219,N_469,N_1854);
nor U7220 (N_7220,N_3292,N_3313);
nand U7221 (N_7221,N_2897,N_876);
xnor U7222 (N_7222,N_117,N_1522);
or U7223 (N_7223,N_2849,N_1568);
nor U7224 (N_7224,N_2097,N_116);
nor U7225 (N_7225,N_1889,N_4407);
nor U7226 (N_7226,N_3539,N_3596);
nor U7227 (N_7227,N_3322,N_4718);
and U7228 (N_7228,N_1490,N_432);
or U7229 (N_7229,N_2350,N_1506);
and U7230 (N_7230,N_2200,N_2719);
nor U7231 (N_7231,N_1057,N_3795);
xor U7232 (N_7232,N_685,N_1621);
and U7233 (N_7233,N_4422,N_4909);
and U7234 (N_7234,N_3782,N_455);
nor U7235 (N_7235,N_72,N_1762);
nor U7236 (N_7236,N_1278,N_3104);
or U7237 (N_7237,N_3268,N_699);
nor U7238 (N_7238,N_1305,N_4388);
xor U7239 (N_7239,N_2837,N_2933);
nor U7240 (N_7240,N_3560,N_3325);
or U7241 (N_7241,N_1180,N_2196);
xnor U7242 (N_7242,N_2711,N_2088);
nor U7243 (N_7243,N_1287,N_1923);
and U7244 (N_7244,N_4614,N_3621);
and U7245 (N_7245,N_4958,N_4270);
and U7246 (N_7246,N_3892,N_4619);
xnor U7247 (N_7247,N_4463,N_3483);
xnor U7248 (N_7248,N_1213,N_3479);
nand U7249 (N_7249,N_4794,N_3099);
xor U7250 (N_7250,N_2066,N_4336);
and U7251 (N_7251,N_2101,N_4889);
nor U7252 (N_7252,N_3406,N_1455);
xnor U7253 (N_7253,N_4430,N_3150);
nor U7254 (N_7254,N_4923,N_4392);
nand U7255 (N_7255,N_4171,N_4349);
nor U7256 (N_7256,N_1111,N_1867);
and U7257 (N_7257,N_1116,N_2032);
or U7258 (N_7258,N_2273,N_1853);
or U7259 (N_7259,N_2331,N_1874);
or U7260 (N_7260,N_2133,N_410);
nor U7261 (N_7261,N_4328,N_927);
nor U7262 (N_7262,N_2164,N_905);
nor U7263 (N_7263,N_1732,N_3279);
xor U7264 (N_7264,N_460,N_1708);
or U7265 (N_7265,N_4854,N_3271);
and U7266 (N_7266,N_1865,N_1021);
xnor U7267 (N_7267,N_1322,N_1504);
or U7268 (N_7268,N_1239,N_29);
or U7269 (N_7269,N_391,N_3738);
nand U7270 (N_7270,N_2426,N_1536);
xor U7271 (N_7271,N_2186,N_941);
nand U7272 (N_7272,N_4221,N_1431);
or U7273 (N_7273,N_690,N_4692);
or U7274 (N_7274,N_3950,N_749);
and U7275 (N_7275,N_1368,N_4788);
xnor U7276 (N_7276,N_1599,N_4159);
or U7277 (N_7277,N_266,N_4498);
nand U7278 (N_7278,N_1905,N_2567);
xor U7279 (N_7279,N_30,N_2904);
nand U7280 (N_7280,N_4751,N_3863);
or U7281 (N_7281,N_2983,N_334);
nand U7282 (N_7282,N_1666,N_3801);
and U7283 (N_7283,N_1,N_1941);
and U7284 (N_7284,N_2548,N_620);
or U7285 (N_7285,N_4129,N_2694);
nand U7286 (N_7286,N_3779,N_3304);
and U7287 (N_7287,N_864,N_4068);
or U7288 (N_7288,N_2620,N_956);
and U7289 (N_7289,N_4957,N_4197);
or U7290 (N_7290,N_2996,N_523);
nor U7291 (N_7291,N_2698,N_1570);
or U7292 (N_7292,N_972,N_1200);
or U7293 (N_7293,N_2793,N_3161);
nor U7294 (N_7294,N_2906,N_4739);
nand U7295 (N_7295,N_2077,N_4272);
nand U7296 (N_7296,N_3788,N_408);
nor U7297 (N_7297,N_1162,N_2665);
or U7298 (N_7298,N_558,N_4091);
or U7299 (N_7299,N_4213,N_2345);
xnor U7300 (N_7300,N_3918,N_2105);
or U7301 (N_7301,N_4812,N_367);
xnor U7302 (N_7302,N_2384,N_3273);
xor U7303 (N_7303,N_4663,N_83);
nor U7304 (N_7304,N_3314,N_2344);
xor U7305 (N_7305,N_4880,N_3909);
xor U7306 (N_7306,N_1309,N_1550);
nor U7307 (N_7307,N_1314,N_3415);
xnor U7308 (N_7308,N_2902,N_906);
or U7309 (N_7309,N_2228,N_2769);
nand U7310 (N_7310,N_3233,N_2116);
xnor U7311 (N_7311,N_4932,N_1273);
and U7312 (N_7312,N_535,N_4103);
or U7313 (N_7313,N_4406,N_1516);
or U7314 (N_7314,N_4756,N_2670);
xnor U7315 (N_7315,N_4268,N_3842);
and U7316 (N_7316,N_1850,N_4534);
or U7317 (N_7317,N_3442,N_1873);
and U7318 (N_7318,N_422,N_2494);
or U7319 (N_7319,N_2507,N_4450);
or U7320 (N_7320,N_2458,N_403);
nand U7321 (N_7321,N_423,N_2598);
nor U7322 (N_7322,N_1335,N_4895);
nor U7323 (N_7323,N_1750,N_230);
or U7324 (N_7324,N_4317,N_3825);
and U7325 (N_7325,N_2470,N_593);
xor U7326 (N_7326,N_3963,N_1763);
and U7327 (N_7327,N_2214,N_2796);
xor U7328 (N_7328,N_2931,N_1819);
xor U7329 (N_7329,N_212,N_15);
nand U7330 (N_7330,N_2024,N_3368);
xnor U7331 (N_7331,N_1102,N_920);
nor U7332 (N_7332,N_3472,N_2924);
nor U7333 (N_7333,N_2803,N_349);
xor U7334 (N_7334,N_2481,N_2720);
or U7335 (N_7335,N_2460,N_3215);
xor U7336 (N_7336,N_3838,N_1445);
nand U7337 (N_7337,N_4804,N_2451);
nand U7338 (N_7338,N_4074,N_4225);
nor U7339 (N_7339,N_712,N_3285);
and U7340 (N_7340,N_823,N_2634);
nor U7341 (N_7341,N_2446,N_1582);
and U7342 (N_7342,N_2819,N_1518);
nor U7343 (N_7343,N_1558,N_299);
nor U7344 (N_7344,N_1713,N_1585);
and U7345 (N_7345,N_3118,N_4448);
or U7346 (N_7346,N_1703,N_2608);
and U7347 (N_7347,N_2815,N_2109);
nor U7348 (N_7348,N_916,N_3781);
nand U7349 (N_7349,N_1408,N_3914);
xor U7350 (N_7350,N_1025,N_1729);
nor U7351 (N_7351,N_4453,N_4616);
and U7352 (N_7352,N_4538,N_2419);
nor U7353 (N_7353,N_1557,N_3935);
and U7354 (N_7354,N_113,N_3358);
and U7355 (N_7355,N_1186,N_4578);
and U7356 (N_7356,N_4085,N_3032);
nand U7357 (N_7357,N_2633,N_3238);
and U7358 (N_7358,N_780,N_2768);
nor U7359 (N_7359,N_2072,N_2026);
nand U7360 (N_7360,N_3431,N_4579);
nor U7361 (N_7361,N_4679,N_2648);
nand U7362 (N_7362,N_2834,N_2631);
and U7363 (N_7363,N_781,N_1687);
nand U7364 (N_7364,N_4518,N_3114);
xnor U7365 (N_7365,N_2949,N_978);
nand U7366 (N_7366,N_2701,N_3765);
nand U7367 (N_7367,N_3184,N_4414);
xnor U7368 (N_7368,N_3974,N_3888);
and U7369 (N_7369,N_3456,N_1039);
nand U7370 (N_7370,N_545,N_4369);
and U7371 (N_7371,N_2165,N_219);
or U7372 (N_7372,N_431,N_4394);
or U7373 (N_7373,N_4231,N_3716);
nand U7374 (N_7374,N_1580,N_320);
nor U7375 (N_7375,N_3614,N_4065);
xnor U7376 (N_7376,N_2462,N_4083);
nand U7377 (N_7377,N_3276,N_2973);
or U7378 (N_7378,N_1245,N_2320);
nand U7379 (N_7379,N_3212,N_3047);
nor U7380 (N_7380,N_1657,N_2820);
and U7381 (N_7381,N_581,N_2011);
and U7382 (N_7382,N_598,N_2742);
xor U7383 (N_7383,N_192,N_2950);
and U7384 (N_7384,N_1406,N_4342);
nor U7385 (N_7385,N_4978,N_2479);
nor U7386 (N_7386,N_4241,N_195);
nand U7387 (N_7387,N_2662,N_3523);
nor U7388 (N_7388,N_640,N_1875);
nor U7389 (N_7389,N_56,N_3300);
or U7390 (N_7390,N_3185,N_3224);
and U7391 (N_7391,N_4200,N_2258);
nor U7392 (N_7392,N_2012,N_2205);
xor U7393 (N_7393,N_1605,N_2168);
nor U7394 (N_7394,N_3429,N_323);
and U7395 (N_7395,N_462,N_2505);
nor U7396 (N_7396,N_2781,N_4626);
and U7397 (N_7397,N_1891,N_596);
and U7398 (N_7398,N_4763,N_2807);
or U7399 (N_7399,N_4391,N_3189);
and U7400 (N_7400,N_433,N_1784);
xnor U7401 (N_7401,N_499,N_3942);
or U7402 (N_7402,N_3109,N_4483);
xor U7403 (N_7403,N_3068,N_3003);
xor U7404 (N_7404,N_4871,N_2668);
or U7405 (N_7405,N_254,N_849);
or U7406 (N_7406,N_1820,N_2357);
and U7407 (N_7407,N_4441,N_1963);
nand U7408 (N_7408,N_8,N_1067);
nor U7409 (N_7409,N_3771,N_1166);
nand U7410 (N_7410,N_3248,N_579);
nor U7411 (N_7411,N_1483,N_933);
or U7412 (N_7412,N_4969,N_696);
nand U7413 (N_7413,N_4243,N_2276);
nand U7414 (N_7414,N_1271,N_1283);
and U7415 (N_7415,N_595,N_3861);
and U7416 (N_7416,N_1539,N_81);
and U7417 (N_7417,N_4409,N_4980);
and U7418 (N_7418,N_682,N_2952);
xnor U7419 (N_7419,N_1861,N_3710);
or U7420 (N_7420,N_2251,N_2082);
and U7421 (N_7421,N_1581,N_3717);
and U7422 (N_7422,N_1842,N_4283);
and U7423 (N_7423,N_547,N_3218);
or U7424 (N_7424,N_3908,N_1447);
or U7425 (N_7425,N_4519,N_4846);
nor U7426 (N_7426,N_3056,N_2865);
nor U7427 (N_7427,N_2121,N_209);
nor U7428 (N_7428,N_2162,N_2035);
and U7429 (N_7429,N_2707,N_339);
nand U7430 (N_7430,N_1527,N_1412);
nor U7431 (N_7431,N_4185,N_1726);
and U7432 (N_7432,N_1009,N_2341);
and U7433 (N_7433,N_3227,N_4451);
xor U7434 (N_7434,N_2414,N_145);
xor U7435 (N_7435,N_4397,N_2893);
and U7436 (N_7436,N_2776,N_4413);
nor U7437 (N_7437,N_855,N_756);
nand U7438 (N_7438,N_1937,N_808);
nand U7439 (N_7439,N_2920,N_4374);
and U7440 (N_7440,N_4525,N_1381);
nor U7441 (N_7441,N_1751,N_4472);
xnor U7442 (N_7442,N_891,N_4509);
nor U7443 (N_7443,N_817,N_1884);
and U7444 (N_7444,N_2352,N_4479);
nor U7445 (N_7445,N_4141,N_2400);
or U7446 (N_7446,N_1042,N_1697);
nor U7447 (N_7447,N_478,N_734);
xor U7448 (N_7448,N_3959,N_2359);
nor U7449 (N_7449,N_3758,N_4604);
nand U7450 (N_7450,N_748,N_2075);
and U7451 (N_7451,N_92,N_3860);
nand U7452 (N_7452,N_3439,N_2723);
nand U7453 (N_7453,N_2535,N_388);
nor U7454 (N_7454,N_2512,N_265);
nor U7455 (N_7455,N_4585,N_2219);
nand U7456 (N_7456,N_3608,N_221);
xor U7457 (N_7457,N_1673,N_4631);
or U7458 (N_7458,N_3870,N_1037);
nand U7459 (N_7459,N_728,N_1855);
xor U7460 (N_7460,N_4357,N_569);
nor U7461 (N_7461,N_405,N_1771);
nand U7462 (N_7462,N_1049,N_32);
nor U7463 (N_7463,N_889,N_1722);
nor U7464 (N_7464,N_4027,N_2226);
nand U7465 (N_7465,N_3597,N_1641);
nor U7466 (N_7466,N_1811,N_747);
or U7467 (N_7467,N_3445,N_255);
and U7468 (N_7468,N_4015,N_1690);
or U7469 (N_7469,N_382,N_4154);
xor U7470 (N_7470,N_1247,N_1664);
or U7471 (N_7471,N_4811,N_1276);
nor U7472 (N_7472,N_2805,N_822);
nor U7473 (N_7473,N_1034,N_1348);
xnor U7474 (N_7474,N_3759,N_1389);
nand U7475 (N_7475,N_2189,N_3413);
and U7476 (N_7476,N_4831,N_2290);
nor U7477 (N_7477,N_1658,N_3085);
nand U7478 (N_7478,N_381,N_2561);
and U7479 (N_7479,N_3615,N_693);
xnor U7480 (N_7480,N_2822,N_1563);
and U7481 (N_7481,N_1212,N_2724);
or U7482 (N_7482,N_181,N_3617);
nand U7483 (N_7483,N_3606,N_1956);
and U7484 (N_7484,N_4603,N_2098);
and U7485 (N_7485,N_1549,N_1770);
or U7486 (N_7486,N_4605,N_3399);
or U7487 (N_7487,N_3008,N_1304);
and U7488 (N_7488,N_2124,N_659);
and U7489 (N_7489,N_3394,N_3377);
nor U7490 (N_7490,N_2998,N_3082);
or U7491 (N_7491,N_1054,N_2159);
and U7492 (N_7492,N_1507,N_841);
or U7493 (N_7493,N_3572,N_12);
nor U7494 (N_7494,N_853,N_1211);
nand U7495 (N_7495,N_97,N_3508);
nor U7496 (N_7496,N_866,N_2922);
or U7497 (N_7497,N_1013,N_3737);
and U7498 (N_7498,N_1831,N_4540);
xnor U7499 (N_7499,N_4267,N_2181);
nor U7500 (N_7500,N_2448,N_2565);
or U7501 (N_7501,N_2676,N_2196);
or U7502 (N_7502,N_1709,N_4826);
or U7503 (N_7503,N_881,N_3104);
or U7504 (N_7504,N_1903,N_3649);
or U7505 (N_7505,N_1296,N_2412);
and U7506 (N_7506,N_1726,N_1504);
nor U7507 (N_7507,N_2179,N_1028);
nor U7508 (N_7508,N_3093,N_2493);
nand U7509 (N_7509,N_1181,N_695);
nand U7510 (N_7510,N_817,N_2517);
nor U7511 (N_7511,N_157,N_522);
or U7512 (N_7512,N_4585,N_3223);
nor U7513 (N_7513,N_3605,N_220);
nor U7514 (N_7514,N_3556,N_2483);
nor U7515 (N_7515,N_1019,N_2628);
nor U7516 (N_7516,N_1916,N_1172);
and U7517 (N_7517,N_4805,N_2423);
nor U7518 (N_7518,N_841,N_4602);
nand U7519 (N_7519,N_32,N_1080);
nor U7520 (N_7520,N_3135,N_1032);
nor U7521 (N_7521,N_1182,N_4736);
nor U7522 (N_7522,N_211,N_3213);
xnor U7523 (N_7523,N_2151,N_4218);
or U7524 (N_7524,N_1313,N_761);
xor U7525 (N_7525,N_2078,N_3660);
nor U7526 (N_7526,N_1988,N_2057);
or U7527 (N_7527,N_2148,N_802);
nor U7528 (N_7528,N_3792,N_3655);
nor U7529 (N_7529,N_2732,N_384);
nor U7530 (N_7530,N_3638,N_4294);
xnor U7531 (N_7531,N_3839,N_1676);
xnor U7532 (N_7532,N_3839,N_659);
and U7533 (N_7533,N_3564,N_1419);
or U7534 (N_7534,N_1055,N_2516);
or U7535 (N_7535,N_65,N_3979);
or U7536 (N_7536,N_1889,N_1117);
xnor U7537 (N_7537,N_3830,N_3972);
nor U7538 (N_7538,N_1550,N_4271);
xnor U7539 (N_7539,N_3272,N_4863);
nor U7540 (N_7540,N_4539,N_2051);
or U7541 (N_7541,N_399,N_3865);
or U7542 (N_7542,N_184,N_3361);
nor U7543 (N_7543,N_3020,N_2741);
and U7544 (N_7544,N_1271,N_4071);
or U7545 (N_7545,N_2507,N_4822);
nand U7546 (N_7546,N_3232,N_1220);
nor U7547 (N_7547,N_4689,N_3521);
and U7548 (N_7548,N_2107,N_2560);
nand U7549 (N_7549,N_2692,N_1945);
xor U7550 (N_7550,N_1400,N_291);
xnor U7551 (N_7551,N_1713,N_1117);
xnor U7552 (N_7552,N_1885,N_767);
or U7553 (N_7553,N_2352,N_2237);
nand U7554 (N_7554,N_3784,N_1209);
and U7555 (N_7555,N_2320,N_2511);
xor U7556 (N_7556,N_4426,N_837);
xnor U7557 (N_7557,N_3103,N_3821);
and U7558 (N_7558,N_3978,N_4406);
nor U7559 (N_7559,N_4358,N_3530);
nand U7560 (N_7560,N_4414,N_2185);
xnor U7561 (N_7561,N_2033,N_3111);
and U7562 (N_7562,N_3635,N_4956);
xor U7563 (N_7563,N_1664,N_2185);
xor U7564 (N_7564,N_4396,N_2601);
and U7565 (N_7565,N_2096,N_2361);
nand U7566 (N_7566,N_2219,N_1886);
nor U7567 (N_7567,N_4116,N_2642);
nand U7568 (N_7568,N_1437,N_534);
nand U7569 (N_7569,N_1187,N_2724);
nor U7570 (N_7570,N_4426,N_864);
nand U7571 (N_7571,N_2605,N_3298);
nor U7572 (N_7572,N_2079,N_373);
or U7573 (N_7573,N_2149,N_2150);
nor U7574 (N_7574,N_1007,N_3340);
nor U7575 (N_7575,N_2696,N_4050);
xnor U7576 (N_7576,N_1255,N_4032);
or U7577 (N_7577,N_4381,N_4522);
or U7578 (N_7578,N_4534,N_3438);
or U7579 (N_7579,N_2364,N_3824);
and U7580 (N_7580,N_25,N_1647);
nand U7581 (N_7581,N_1161,N_3607);
xor U7582 (N_7582,N_152,N_4184);
nand U7583 (N_7583,N_1413,N_757);
nor U7584 (N_7584,N_966,N_1836);
and U7585 (N_7585,N_4188,N_2700);
and U7586 (N_7586,N_3970,N_4634);
and U7587 (N_7587,N_983,N_3216);
xnor U7588 (N_7588,N_3749,N_4535);
nand U7589 (N_7589,N_3087,N_2378);
and U7590 (N_7590,N_2307,N_1939);
and U7591 (N_7591,N_4211,N_2768);
xor U7592 (N_7592,N_929,N_4485);
or U7593 (N_7593,N_3071,N_2478);
or U7594 (N_7594,N_1722,N_3549);
xor U7595 (N_7595,N_1959,N_1534);
or U7596 (N_7596,N_943,N_4004);
and U7597 (N_7597,N_2797,N_3834);
nand U7598 (N_7598,N_4900,N_4801);
nand U7599 (N_7599,N_3478,N_3461);
or U7600 (N_7600,N_1669,N_3765);
or U7601 (N_7601,N_734,N_530);
or U7602 (N_7602,N_1605,N_69);
nor U7603 (N_7603,N_3789,N_1487);
nand U7604 (N_7604,N_1152,N_4323);
and U7605 (N_7605,N_3848,N_195);
nor U7606 (N_7606,N_1152,N_4830);
nor U7607 (N_7607,N_3844,N_231);
or U7608 (N_7608,N_369,N_1375);
or U7609 (N_7609,N_833,N_4837);
xnor U7610 (N_7610,N_4823,N_4826);
nor U7611 (N_7611,N_4160,N_1511);
xor U7612 (N_7612,N_4432,N_390);
or U7613 (N_7613,N_1886,N_1178);
nor U7614 (N_7614,N_2714,N_1615);
and U7615 (N_7615,N_3511,N_4878);
xor U7616 (N_7616,N_2220,N_1069);
or U7617 (N_7617,N_1844,N_4802);
nand U7618 (N_7618,N_2313,N_270);
nor U7619 (N_7619,N_3933,N_170);
or U7620 (N_7620,N_3240,N_2429);
xnor U7621 (N_7621,N_4835,N_2076);
and U7622 (N_7622,N_3469,N_4829);
nor U7623 (N_7623,N_2529,N_1948);
xor U7624 (N_7624,N_4234,N_4553);
nor U7625 (N_7625,N_3522,N_4146);
xor U7626 (N_7626,N_2159,N_1772);
or U7627 (N_7627,N_1659,N_4914);
xnor U7628 (N_7628,N_4992,N_2765);
xor U7629 (N_7629,N_3654,N_2825);
or U7630 (N_7630,N_3439,N_1028);
or U7631 (N_7631,N_4528,N_3792);
nor U7632 (N_7632,N_1821,N_3188);
xor U7633 (N_7633,N_2430,N_2383);
nand U7634 (N_7634,N_1049,N_2500);
nor U7635 (N_7635,N_3936,N_1962);
nand U7636 (N_7636,N_1984,N_4733);
and U7637 (N_7637,N_664,N_1538);
and U7638 (N_7638,N_2371,N_4148);
and U7639 (N_7639,N_2544,N_1702);
nand U7640 (N_7640,N_2864,N_4923);
or U7641 (N_7641,N_3193,N_1314);
nor U7642 (N_7642,N_4882,N_971);
and U7643 (N_7643,N_2530,N_1953);
nand U7644 (N_7644,N_33,N_207);
xnor U7645 (N_7645,N_278,N_360);
and U7646 (N_7646,N_764,N_3646);
or U7647 (N_7647,N_1553,N_1383);
and U7648 (N_7648,N_3781,N_2196);
or U7649 (N_7649,N_4196,N_3102);
nor U7650 (N_7650,N_4086,N_335);
or U7651 (N_7651,N_2868,N_2415);
nor U7652 (N_7652,N_1356,N_3399);
nor U7653 (N_7653,N_4095,N_1366);
xor U7654 (N_7654,N_4678,N_3389);
and U7655 (N_7655,N_494,N_430);
nor U7656 (N_7656,N_3996,N_4480);
nor U7657 (N_7657,N_3362,N_228);
and U7658 (N_7658,N_4755,N_3986);
xor U7659 (N_7659,N_2190,N_3138);
nand U7660 (N_7660,N_3056,N_2431);
and U7661 (N_7661,N_321,N_598);
and U7662 (N_7662,N_294,N_4100);
xor U7663 (N_7663,N_4052,N_4601);
or U7664 (N_7664,N_4932,N_120);
or U7665 (N_7665,N_535,N_476);
nor U7666 (N_7666,N_2781,N_4508);
or U7667 (N_7667,N_1933,N_974);
or U7668 (N_7668,N_4108,N_1218);
and U7669 (N_7669,N_756,N_4635);
nor U7670 (N_7670,N_2433,N_3389);
and U7671 (N_7671,N_1850,N_2073);
or U7672 (N_7672,N_507,N_504);
xor U7673 (N_7673,N_2379,N_4029);
xnor U7674 (N_7674,N_4043,N_3134);
and U7675 (N_7675,N_2319,N_3671);
xnor U7676 (N_7676,N_2058,N_1514);
nand U7677 (N_7677,N_4439,N_4347);
xor U7678 (N_7678,N_3867,N_4919);
nand U7679 (N_7679,N_3296,N_4120);
nand U7680 (N_7680,N_4675,N_434);
and U7681 (N_7681,N_3267,N_1595);
or U7682 (N_7682,N_2716,N_3174);
and U7683 (N_7683,N_2832,N_3827);
xnor U7684 (N_7684,N_2074,N_2684);
nor U7685 (N_7685,N_2590,N_24);
or U7686 (N_7686,N_2793,N_2972);
or U7687 (N_7687,N_4862,N_3436);
xnor U7688 (N_7688,N_926,N_2404);
nand U7689 (N_7689,N_3282,N_3020);
or U7690 (N_7690,N_2566,N_1513);
xor U7691 (N_7691,N_3290,N_1119);
nand U7692 (N_7692,N_897,N_627);
nor U7693 (N_7693,N_1476,N_4185);
or U7694 (N_7694,N_1188,N_1291);
nor U7695 (N_7695,N_3032,N_572);
xnor U7696 (N_7696,N_3218,N_2960);
or U7697 (N_7697,N_1431,N_2295);
xor U7698 (N_7698,N_556,N_1411);
and U7699 (N_7699,N_2710,N_2518);
or U7700 (N_7700,N_1010,N_1074);
nor U7701 (N_7701,N_4019,N_489);
xor U7702 (N_7702,N_3135,N_3278);
nand U7703 (N_7703,N_3295,N_4663);
or U7704 (N_7704,N_310,N_384);
nor U7705 (N_7705,N_495,N_2063);
and U7706 (N_7706,N_3362,N_4884);
xor U7707 (N_7707,N_2060,N_3270);
and U7708 (N_7708,N_363,N_2289);
xor U7709 (N_7709,N_698,N_4298);
nand U7710 (N_7710,N_3555,N_2896);
and U7711 (N_7711,N_1100,N_2940);
xnor U7712 (N_7712,N_1580,N_2418);
xor U7713 (N_7713,N_1369,N_2155);
or U7714 (N_7714,N_104,N_393);
or U7715 (N_7715,N_3006,N_1811);
and U7716 (N_7716,N_2123,N_3445);
nor U7717 (N_7717,N_1611,N_3362);
or U7718 (N_7718,N_532,N_1270);
xor U7719 (N_7719,N_3625,N_4607);
or U7720 (N_7720,N_4169,N_4171);
or U7721 (N_7721,N_1335,N_997);
and U7722 (N_7722,N_1209,N_3623);
or U7723 (N_7723,N_1563,N_2746);
xnor U7724 (N_7724,N_1751,N_1973);
xnor U7725 (N_7725,N_744,N_2271);
nor U7726 (N_7726,N_324,N_1110);
xor U7727 (N_7727,N_1234,N_18);
nor U7728 (N_7728,N_2794,N_4917);
or U7729 (N_7729,N_657,N_209);
and U7730 (N_7730,N_1026,N_3622);
nand U7731 (N_7731,N_4547,N_483);
nand U7732 (N_7732,N_4596,N_1088);
xnor U7733 (N_7733,N_3489,N_3670);
nor U7734 (N_7734,N_1671,N_3935);
nand U7735 (N_7735,N_4747,N_3682);
and U7736 (N_7736,N_47,N_43);
and U7737 (N_7737,N_363,N_2535);
or U7738 (N_7738,N_4537,N_3015);
xnor U7739 (N_7739,N_176,N_2540);
xnor U7740 (N_7740,N_354,N_4476);
nand U7741 (N_7741,N_1959,N_366);
nand U7742 (N_7742,N_3827,N_3266);
or U7743 (N_7743,N_3236,N_3290);
and U7744 (N_7744,N_770,N_4960);
xnor U7745 (N_7745,N_3714,N_3313);
or U7746 (N_7746,N_3828,N_1904);
nand U7747 (N_7747,N_4429,N_4845);
nor U7748 (N_7748,N_4279,N_3448);
and U7749 (N_7749,N_2242,N_636);
or U7750 (N_7750,N_4071,N_1633);
and U7751 (N_7751,N_3011,N_3243);
and U7752 (N_7752,N_224,N_1520);
nand U7753 (N_7753,N_2713,N_489);
and U7754 (N_7754,N_51,N_4332);
and U7755 (N_7755,N_2325,N_1162);
or U7756 (N_7756,N_3218,N_3222);
nor U7757 (N_7757,N_1627,N_3044);
nand U7758 (N_7758,N_2128,N_2191);
or U7759 (N_7759,N_166,N_4007);
xor U7760 (N_7760,N_1757,N_2575);
nor U7761 (N_7761,N_2576,N_2090);
xor U7762 (N_7762,N_609,N_2443);
nand U7763 (N_7763,N_4355,N_1290);
or U7764 (N_7764,N_4519,N_2267);
and U7765 (N_7765,N_1708,N_4466);
xnor U7766 (N_7766,N_4828,N_4832);
nand U7767 (N_7767,N_1766,N_4731);
xnor U7768 (N_7768,N_1792,N_4122);
nand U7769 (N_7769,N_1212,N_2220);
and U7770 (N_7770,N_3223,N_2453);
or U7771 (N_7771,N_2566,N_1364);
and U7772 (N_7772,N_371,N_1038);
and U7773 (N_7773,N_4972,N_713);
or U7774 (N_7774,N_3886,N_3569);
or U7775 (N_7775,N_3069,N_1071);
or U7776 (N_7776,N_2905,N_2811);
and U7777 (N_7777,N_2740,N_4204);
nor U7778 (N_7778,N_3070,N_3383);
xnor U7779 (N_7779,N_265,N_3788);
nor U7780 (N_7780,N_1121,N_2663);
nand U7781 (N_7781,N_3396,N_183);
nor U7782 (N_7782,N_1195,N_4338);
or U7783 (N_7783,N_4142,N_4245);
nand U7784 (N_7784,N_562,N_2830);
and U7785 (N_7785,N_3543,N_1549);
nand U7786 (N_7786,N_1369,N_2740);
or U7787 (N_7787,N_4759,N_1553);
and U7788 (N_7788,N_230,N_773);
xor U7789 (N_7789,N_1452,N_4774);
and U7790 (N_7790,N_4319,N_65);
and U7791 (N_7791,N_691,N_3519);
xor U7792 (N_7792,N_4943,N_2338);
or U7793 (N_7793,N_3736,N_2300);
nor U7794 (N_7794,N_4503,N_233);
and U7795 (N_7795,N_1538,N_4217);
and U7796 (N_7796,N_2680,N_2561);
nand U7797 (N_7797,N_3906,N_3527);
and U7798 (N_7798,N_3960,N_2423);
nor U7799 (N_7799,N_3131,N_2196);
or U7800 (N_7800,N_4039,N_725);
nand U7801 (N_7801,N_3510,N_143);
and U7802 (N_7802,N_4687,N_2506);
and U7803 (N_7803,N_3336,N_3711);
nor U7804 (N_7804,N_936,N_3373);
nand U7805 (N_7805,N_1355,N_4062);
nand U7806 (N_7806,N_3383,N_1809);
xor U7807 (N_7807,N_4887,N_3999);
nand U7808 (N_7808,N_778,N_3911);
xnor U7809 (N_7809,N_237,N_4704);
xnor U7810 (N_7810,N_1841,N_3367);
and U7811 (N_7811,N_4037,N_2332);
nor U7812 (N_7812,N_4233,N_3773);
xor U7813 (N_7813,N_4375,N_2958);
nor U7814 (N_7814,N_3487,N_4105);
nand U7815 (N_7815,N_449,N_1738);
nand U7816 (N_7816,N_4285,N_2905);
nand U7817 (N_7817,N_2600,N_4565);
nand U7818 (N_7818,N_594,N_230);
nand U7819 (N_7819,N_4407,N_203);
or U7820 (N_7820,N_884,N_759);
nor U7821 (N_7821,N_1765,N_1078);
xnor U7822 (N_7822,N_3078,N_4441);
and U7823 (N_7823,N_2822,N_2466);
nand U7824 (N_7824,N_4896,N_2962);
nor U7825 (N_7825,N_2953,N_3553);
nor U7826 (N_7826,N_478,N_148);
xnor U7827 (N_7827,N_1219,N_1955);
and U7828 (N_7828,N_1568,N_4297);
nand U7829 (N_7829,N_1710,N_4084);
nor U7830 (N_7830,N_2659,N_3589);
and U7831 (N_7831,N_3267,N_1902);
and U7832 (N_7832,N_320,N_1958);
xor U7833 (N_7833,N_4778,N_2294);
nand U7834 (N_7834,N_2652,N_4936);
xor U7835 (N_7835,N_3456,N_2905);
nor U7836 (N_7836,N_2660,N_4759);
xnor U7837 (N_7837,N_1290,N_4076);
nor U7838 (N_7838,N_492,N_2395);
nand U7839 (N_7839,N_2838,N_1637);
xnor U7840 (N_7840,N_2604,N_1464);
xor U7841 (N_7841,N_2383,N_3141);
or U7842 (N_7842,N_387,N_574);
and U7843 (N_7843,N_260,N_1168);
and U7844 (N_7844,N_4588,N_4229);
nor U7845 (N_7845,N_489,N_3797);
and U7846 (N_7846,N_55,N_4829);
or U7847 (N_7847,N_3139,N_3816);
nand U7848 (N_7848,N_627,N_4629);
or U7849 (N_7849,N_1846,N_1360);
nor U7850 (N_7850,N_3675,N_3974);
nand U7851 (N_7851,N_2762,N_4039);
or U7852 (N_7852,N_2384,N_4791);
or U7853 (N_7853,N_1015,N_312);
nor U7854 (N_7854,N_871,N_1713);
nand U7855 (N_7855,N_2923,N_4181);
and U7856 (N_7856,N_4354,N_4062);
nand U7857 (N_7857,N_633,N_3122);
nand U7858 (N_7858,N_862,N_1558);
nand U7859 (N_7859,N_2651,N_2185);
and U7860 (N_7860,N_4742,N_3230);
nor U7861 (N_7861,N_256,N_4497);
and U7862 (N_7862,N_4249,N_4755);
nor U7863 (N_7863,N_4722,N_3029);
or U7864 (N_7864,N_2245,N_1494);
and U7865 (N_7865,N_1268,N_3832);
nand U7866 (N_7866,N_1586,N_3295);
nand U7867 (N_7867,N_4691,N_305);
nand U7868 (N_7868,N_2958,N_4477);
xor U7869 (N_7869,N_973,N_415);
and U7870 (N_7870,N_4389,N_4206);
nand U7871 (N_7871,N_368,N_1120);
nand U7872 (N_7872,N_408,N_1905);
and U7873 (N_7873,N_1620,N_2301);
or U7874 (N_7874,N_2541,N_2880);
and U7875 (N_7875,N_1670,N_2087);
nand U7876 (N_7876,N_1343,N_1211);
or U7877 (N_7877,N_73,N_990);
xor U7878 (N_7878,N_4752,N_2991);
and U7879 (N_7879,N_2143,N_3146);
nand U7880 (N_7880,N_4086,N_4099);
nand U7881 (N_7881,N_1332,N_3440);
or U7882 (N_7882,N_3596,N_2224);
and U7883 (N_7883,N_4741,N_125);
xnor U7884 (N_7884,N_574,N_2081);
or U7885 (N_7885,N_4876,N_3180);
xnor U7886 (N_7886,N_2599,N_2864);
and U7887 (N_7887,N_1914,N_2418);
nand U7888 (N_7888,N_122,N_1737);
or U7889 (N_7889,N_1837,N_2748);
nand U7890 (N_7890,N_4289,N_4695);
nor U7891 (N_7891,N_561,N_1220);
xnor U7892 (N_7892,N_2821,N_939);
nor U7893 (N_7893,N_2192,N_522);
or U7894 (N_7894,N_823,N_1220);
and U7895 (N_7895,N_2861,N_591);
nor U7896 (N_7896,N_2827,N_4023);
nand U7897 (N_7897,N_1938,N_2869);
nor U7898 (N_7898,N_4064,N_3480);
and U7899 (N_7899,N_245,N_699);
or U7900 (N_7900,N_935,N_398);
or U7901 (N_7901,N_4638,N_4012);
nor U7902 (N_7902,N_1590,N_4735);
or U7903 (N_7903,N_1861,N_2741);
and U7904 (N_7904,N_76,N_3288);
xor U7905 (N_7905,N_4784,N_4252);
nor U7906 (N_7906,N_3971,N_1704);
nor U7907 (N_7907,N_2630,N_2651);
nand U7908 (N_7908,N_920,N_2850);
and U7909 (N_7909,N_1473,N_4325);
or U7910 (N_7910,N_3170,N_457);
xor U7911 (N_7911,N_2394,N_1192);
nand U7912 (N_7912,N_3924,N_1122);
and U7913 (N_7913,N_736,N_3721);
and U7914 (N_7914,N_265,N_755);
xnor U7915 (N_7915,N_2769,N_2254);
nor U7916 (N_7916,N_3581,N_843);
nor U7917 (N_7917,N_1839,N_2136);
or U7918 (N_7918,N_2119,N_3538);
xor U7919 (N_7919,N_2685,N_1035);
nor U7920 (N_7920,N_4991,N_734);
and U7921 (N_7921,N_3831,N_2938);
nor U7922 (N_7922,N_606,N_2707);
nor U7923 (N_7923,N_3072,N_3513);
and U7924 (N_7924,N_959,N_3113);
nor U7925 (N_7925,N_4197,N_2680);
and U7926 (N_7926,N_1858,N_1472);
nand U7927 (N_7927,N_1953,N_3552);
and U7928 (N_7928,N_1789,N_912);
nor U7929 (N_7929,N_1557,N_3657);
nand U7930 (N_7930,N_218,N_2225);
xnor U7931 (N_7931,N_4806,N_4642);
xor U7932 (N_7932,N_3147,N_4767);
nand U7933 (N_7933,N_1048,N_3531);
nor U7934 (N_7934,N_2880,N_3656);
and U7935 (N_7935,N_2544,N_838);
or U7936 (N_7936,N_3173,N_3561);
nand U7937 (N_7937,N_997,N_2693);
and U7938 (N_7938,N_1981,N_4129);
or U7939 (N_7939,N_3981,N_2445);
nor U7940 (N_7940,N_818,N_2950);
nor U7941 (N_7941,N_3782,N_3629);
or U7942 (N_7942,N_3218,N_4322);
and U7943 (N_7943,N_2798,N_3183);
or U7944 (N_7944,N_140,N_4558);
xor U7945 (N_7945,N_3098,N_4842);
nand U7946 (N_7946,N_137,N_1081);
and U7947 (N_7947,N_56,N_1383);
or U7948 (N_7948,N_490,N_1813);
or U7949 (N_7949,N_3116,N_4157);
and U7950 (N_7950,N_382,N_1971);
or U7951 (N_7951,N_1305,N_119);
and U7952 (N_7952,N_721,N_497);
and U7953 (N_7953,N_1283,N_3944);
and U7954 (N_7954,N_1608,N_156);
or U7955 (N_7955,N_3967,N_2008);
and U7956 (N_7956,N_1326,N_941);
nand U7957 (N_7957,N_470,N_2125);
xor U7958 (N_7958,N_1552,N_3275);
xor U7959 (N_7959,N_4258,N_2183);
nand U7960 (N_7960,N_1278,N_2839);
xnor U7961 (N_7961,N_1357,N_414);
nor U7962 (N_7962,N_223,N_1646);
nand U7963 (N_7963,N_4510,N_2095);
nor U7964 (N_7964,N_4777,N_3764);
and U7965 (N_7965,N_1825,N_219);
nand U7966 (N_7966,N_2624,N_1818);
nand U7967 (N_7967,N_88,N_2378);
nand U7968 (N_7968,N_299,N_2001);
and U7969 (N_7969,N_2387,N_3138);
nand U7970 (N_7970,N_1926,N_1580);
xnor U7971 (N_7971,N_191,N_94);
and U7972 (N_7972,N_3927,N_3196);
nor U7973 (N_7973,N_3021,N_4105);
nor U7974 (N_7974,N_4054,N_2681);
or U7975 (N_7975,N_591,N_1700);
nand U7976 (N_7976,N_1233,N_3339);
nand U7977 (N_7977,N_3821,N_2646);
nand U7978 (N_7978,N_2110,N_2279);
or U7979 (N_7979,N_37,N_133);
nand U7980 (N_7980,N_550,N_892);
or U7981 (N_7981,N_1793,N_4397);
nand U7982 (N_7982,N_3231,N_3166);
and U7983 (N_7983,N_2498,N_2850);
and U7984 (N_7984,N_4716,N_2862);
xor U7985 (N_7985,N_1345,N_4092);
nor U7986 (N_7986,N_2148,N_792);
xor U7987 (N_7987,N_3245,N_2331);
nor U7988 (N_7988,N_2541,N_1760);
nor U7989 (N_7989,N_2001,N_3639);
and U7990 (N_7990,N_3215,N_4416);
nand U7991 (N_7991,N_1081,N_1782);
and U7992 (N_7992,N_1406,N_1176);
or U7993 (N_7993,N_2132,N_475);
nand U7994 (N_7994,N_4445,N_1763);
or U7995 (N_7995,N_2835,N_4713);
nand U7996 (N_7996,N_445,N_4371);
nand U7997 (N_7997,N_230,N_3900);
nor U7998 (N_7998,N_1433,N_868);
or U7999 (N_7999,N_2164,N_3712);
or U8000 (N_8000,N_3355,N_2580);
nand U8001 (N_8001,N_3831,N_112);
or U8002 (N_8002,N_2037,N_4142);
nor U8003 (N_8003,N_1775,N_4129);
or U8004 (N_8004,N_1096,N_2675);
or U8005 (N_8005,N_3230,N_4141);
and U8006 (N_8006,N_4738,N_3700);
or U8007 (N_8007,N_182,N_3562);
nor U8008 (N_8008,N_3094,N_757);
and U8009 (N_8009,N_4535,N_2869);
and U8010 (N_8010,N_4849,N_2023);
and U8011 (N_8011,N_4338,N_1193);
nand U8012 (N_8012,N_3154,N_3170);
and U8013 (N_8013,N_700,N_3225);
nor U8014 (N_8014,N_2792,N_2579);
or U8015 (N_8015,N_2151,N_4577);
nor U8016 (N_8016,N_1988,N_3234);
nand U8017 (N_8017,N_4203,N_4706);
or U8018 (N_8018,N_3619,N_2625);
nand U8019 (N_8019,N_353,N_3777);
xor U8020 (N_8020,N_3086,N_2393);
nor U8021 (N_8021,N_721,N_968);
nand U8022 (N_8022,N_2442,N_1311);
or U8023 (N_8023,N_4104,N_982);
and U8024 (N_8024,N_4420,N_2207);
or U8025 (N_8025,N_1030,N_3930);
or U8026 (N_8026,N_3857,N_4798);
or U8027 (N_8027,N_150,N_3807);
and U8028 (N_8028,N_2467,N_2744);
nor U8029 (N_8029,N_4618,N_2031);
or U8030 (N_8030,N_4017,N_3760);
and U8031 (N_8031,N_4693,N_1071);
nand U8032 (N_8032,N_4994,N_189);
or U8033 (N_8033,N_930,N_2515);
and U8034 (N_8034,N_2174,N_1459);
or U8035 (N_8035,N_3567,N_593);
xnor U8036 (N_8036,N_27,N_1641);
nand U8037 (N_8037,N_323,N_1231);
nand U8038 (N_8038,N_147,N_3013);
xor U8039 (N_8039,N_279,N_4117);
xnor U8040 (N_8040,N_1830,N_3333);
xnor U8041 (N_8041,N_2792,N_1615);
nor U8042 (N_8042,N_3626,N_1194);
and U8043 (N_8043,N_1809,N_1567);
and U8044 (N_8044,N_3991,N_15);
xor U8045 (N_8045,N_3886,N_1378);
nand U8046 (N_8046,N_1911,N_4101);
nor U8047 (N_8047,N_4066,N_661);
and U8048 (N_8048,N_3639,N_1137);
xor U8049 (N_8049,N_4169,N_3984);
nand U8050 (N_8050,N_1133,N_4966);
xnor U8051 (N_8051,N_1099,N_3515);
xor U8052 (N_8052,N_4212,N_2604);
xnor U8053 (N_8053,N_2069,N_2719);
nand U8054 (N_8054,N_4119,N_3999);
or U8055 (N_8055,N_692,N_920);
and U8056 (N_8056,N_1577,N_5);
nand U8057 (N_8057,N_870,N_3740);
nand U8058 (N_8058,N_4116,N_354);
nand U8059 (N_8059,N_1316,N_2229);
nand U8060 (N_8060,N_4888,N_3234);
or U8061 (N_8061,N_3143,N_4242);
or U8062 (N_8062,N_2675,N_2114);
and U8063 (N_8063,N_221,N_1138);
xor U8064 (N_8064,N_410,N_2580);
or U8065 (N_8065,N_2406,N_3470);
or U8066 (N_8066,N_3984,N_2307);
nand U8067 (N_8067,N_293,N_2160);
and U8068 (N_8068,N_1317,N_4777);
or U8069 (N_8069,N_4462,N_2386);
nand U8070 (N_8070,N_1246,N_3586);
and U8071 (N_8071,N_4182,N_1234);
nor U8072 (N_8072,N_2741,N_2001);
xor U8073 (N_8073,N_3897,N_1373);
nand U8074 (N_8074,N_2661,N_662);
and U8075 (N_8075,N_3537,N_4350);
or U8076 (N_8076,N_1589,N_1093);
and U8077 (N_8077,N_4831,N_4109);
nor U8078 (N_8078,N_3168,N_1970);
xor U8079 (N_8079,N_3457,N_4446);
xor U8080 (N_8080,N_991,N_3284);
xnor U8081 (N_8081,N_1782,N_1204);
xor U8082 (N_8082,N_3968,N_4890);
xnor U8083 (N_8083,N_2684,N_519);
or U8084 (N_8084,N_4251,N_4977);
xor U8085 (N_8085,N_3995,N_558);
nor U8086 (N_8086,N_584,N_1448);
and U8087 (N_8087,N_1776,N_2603);
and U8088 (N_8088,N_1131,N_1496);
xnor U8089 (N_8089,N_4530,N_1637);
nor U8090 (N_8090,N_2901,N_4268);
and U8091 (N_8091,N_445,N_4968);
xnor U8092 (N_8092,N_4396,N_3229);
xor U8093 (N_8093,N_4290,N_4596);
nand U8094 (N_8094,N_4650,N_4027);
and U8095 (N_8095,N_4434,N_3442);
nand U8096 (N_8096,N_939,N_1751);
nor U8097 (N_8097,N_2756,N_4147);
or U8098 (N_8098,N_3719,N_4976);
nor U8099 (N_8099,N_3373,N_2438);
nor U8100 (N_8100,N_234,N_4813);
nand U8101 (N_8101,N_2818,N_2152);
nand U8102 (N_8102,N_1079,N_4505);
and U8103 (N_8103,N_709,N_1926);
and U8104 (N_8104,N_696,N_4166);
and U8105 (N_8105,N_888,N_964);
or U8106 (N_8106,N_1497,N_4762);
and U8107 (N_8107,N_2950,N_308);
nor U8108 (N_8108,N_1274,N_4598);
or U8109 (N_8109,N_323,N_2675);
nor U8110 (N_8110,N_116,N_4497);
xnor U8111 (N_8111,N_3927,N_1583);
or U8112 (N_8112,N_4050,N_2648);
nand U8113 (N_8113,N_3750,N_3676);
xnor U8114 (N_8114,N_448,N_2385);
nor U8115 (N_8115,N_3091,N_2158);
xor U8116 (N_8116,N_3079,N_3645);
nand U8117 (N_8117,N_4065,N_1967);
nand U8118 (N_8118,N_2374,N_584);
or U8119 (N_8119,N_534,N_1493);
or U8120 (N_8120,N_3819,N_1551);
or U8121 (N_8121,N_4648,N_4971);
or U8122 (N_8122,N_1812,N_655);
nor U8123 (N_8123,N_3905,N_3172);
and U8124 (N_8124,N_697,N_3931);
xnor U8125 (N_8125,N_2147,N_3596);
nand U8126 (N_8126,N_3020,N_4345);
or U8127 (N_8127,N_1439,N_571);
or U8128 (N_8128,N_4038,N_1276);
or U8129 (N_8129,N_2154,N_2281);
or U8130 (N_8130,N_489,N_1897);
or U8131 (N_8131,N_2724,N_1392);
xnor U8132 (N_8132,N_394,N_3609);
xor U8133 (N_8133,N_1546,N_2523);
or U8134 (N_8134,N_984,N_4504);
and U8135 (N_8135,N_1119,N_2514);
and U8136 (N_8136,N_2932,N_1936);
and U8137 (N_8137,N_3021,N_2292);
or U8138 (N_8138,N_494,N_4021);
nor U8139 (N_8139,N_4777,N_1727);
and U8140 (N_8140,N_3603,N_975);
nor U8141 (N_8141,N_1468,N_1458);
and U8142 (N_8142,N_329,N_3599);
nor U8143 (N_8143,N_4212,N_4339);
nand U8144 (N_8144,N_4376,N_1285);
xor U8145 (N_8145,N_4306,N_1387);
or U8146 (N_8146,N_2841,N_4387);
xnor U8147 (N_8147,N_129,N_1872);
xnor U8148 (N_8148,N_1074,N_1980);
xnor U8149 (N_8149,N_3960,N_3903);
nor U8150 (N_8150,N_3769,N_3156);
nand U8151 (N_8151,N_1703,N_725);
nor U8152 (N_8152,N_2483,N_163);
xnor U8153 (N_8153,N_2893,N_1934);
and U8154 (N_8154,N_1313,N_390);
and U8155 (N_8155,N_4192,N_3654);
or U8156 (N_8156,N_1843,N_4668);
xnor U8157 (N_8157,N_4610,N_4332);
nand U8158 (N_8158,N_358,N_4537);
nand U8159 (N_8159,N_3307,N_3341);
xnor U8160 (N_8160,N_2312,N_455);
and U8161 (N_8161,N_2607,N_503);
xnor U8162 (N_8162,N_3065,N_736);
and U8163 (N_8163,N_1899,N_2954);
nor U8164 (N_8164,N_4877,N_4092);
or U8165 (N_8165,N_446,N_4530);
xor U8166 (N_8166,N_4905,N_3106);
or U8167 (N_8167,N_3153,N_2062);
xnor U8168 (N_8168,N_215,N_2960);
and U8169 (N_8169,N_1984,N_4606);
xnor U8170 (N_8170,N_3252,N_3937);
nand U8171 (N_8171,N_1168,N_2607);
nand U8172 (N_8172,N_2785,N_18);
nand U8173 (N_8173,N_1477,N_4593);
or U8174 (N_8174,N_2995,N_3537);
and U8175 (N_8175,N_3610,N_2054);
xor U8176 (N_8176,N_2924,N_567);
nor U8177 (N_8177,N_3342,N_961);
or U8178 (N_8178,N_1348,N_3146);
or U8179 (N_8179,N_2959,N_4165);
xor U8180 (N_8180,N_684,N_957);
or U8181 (N_8181,N_2081,N_3951);
or U8182 (N_8182,N_3836,N_2119);
and U8183 (N_8183,N_239,N_800);
nand U8184 (N_8184,N_2826,N_2644);
xnor U8185 (N_8185,N_4295,N_3560);
xnor U8186 (N_8186,N_2182,N_3688);
and U8187 (N_8187,N_410,N_4150);
nand U8188 (N_8188,N_1992,N_1899);
and U8189 (N_8189,N_1647,N_3364);
nor U8190 (N_8190,N_2117,N_3903);
nand U8191 (N_8191,N_4462,N_1388);
and U8192 (N_8192,N_2389,N_1100);
xor U8193 (N_8193,N_3805,N_3621);
xor U8194 (N_8194,N_2332,N_2905);
nor U8195 (N_8195,N_374,N_2839);
xnor U8196 (N_8196,N_1173,N_4469);
and U8197 (N_8197,N_1165,N_185);
nor U8198 (N_8198,N_3646,N_2191);
xnor U8199 (N_8199,N_4250,N_3468);
nand U8200 (N_8200,N_3246,N_1042);
or U8201 (N_8201,N_1115,N_388);
xor U8202 (N_8202,N_3622,N_4515);
and U8203 (N_8203,N_2091,N_1824);
and U8204 (N_8204,N_2594,N_700);
nand U8205 (N_8205,N_3723,N_3320);
nor U8206 (N_8206,N_2799,N_3723);
or U8207 (N_8207,N_3001,N_3234);
and U8208 (N_8208,N_2768,N_2828);
xnor U8209 (N_8209,N_890,N_800);
nor U8210 (N_8210,N_1030,N_4407);
xor U8211 (N_8211,N_1408,N_2593);
and U8212 (N_8212,N_4101,N_2934);
nand U8213 (N_8213,N_3886,N_881);
or U8214 (N_8214,N_341,N_1798);
nor U8215 (N_8215,N_869,N_65);
nor U8216 (N_8216,N_4401,N_4986);
and U8217 (N_8217,N_4261,N_4829);
nand U8218 (N_8218,N_2546,N_2767);
or U8219 (N_8219,N_3,N_1291);
xor U8220 (N_8220,N_954,N_1990);
and U8221 (N_8221,N_1097,N_1871);
or U8222 (N_8222,N_3479,N_1850);
xnor U8223 (N_8223,N_921,N_924);
or U8224 (N_8224,N_4961,N_1209);
or U8225 (N_8225,N_1604,N_2710);
nor U8226 (N_8226,N_2067,N_299);
or U8227 (N_8227,N_736,N_3307);
xor U8228 (N_8228,N_4776,N_919);
and U8229 (N_8229,N_4879,N_3928);
nor U8230 (N_8230,N_2190,N_502);
nand U8231 (N_8231,N_1444,N_2533);
and U8232 (N_8232,N_2447,N_4347);
xor U8233 (N_8233,N_4812,N_3218);
or U8234 (N_8234,N_1672,N_20);
or U8235 (N_8235,N_63,N_3028);
and U8236 (N_8236,N_1148,N_4101);
nor U8237 (N_8237,N_1775,N_4105);
nand U8238 (N_8238,N_4102,N_2036);
nor U8239 (N_8239,N_4183,N_1349);
nand U8240 (N_8240,N_2668,N_2302);
and U8241 (N_8241,N_2184,N_3508);
and U8242 (N_8242,N_4136,N_1562);
or U8243 (N_8243,N_2500,N_2802);
or U8244 (N_8244,N_1571,N_4172);
xor U8245 (N_8245,N_2904,N_4476);
and U8246 (N_8246,N_3944,N_3461);
and U8247 (N_8247,N_2358,N_4057);
and U8248 (N_8248,N_40,N_3728);
nor U8249 (N_8249,N_2856,N_685);
and U8250 (N_8250,N_4369,N_4129);
and U8251 (N_8251,N_4795,N_2116);
and U8252 (N_8252,N_3354,N_1589);
or U8253 (N_8253,N_1189,N_2701);
xor U8254 (N_8254,N_3569,N_1942);
nand U8255 (N_8255,N_3333,N_814);
and U8256 (N_8256,N_1110,N_494);
nand U8257 (N_8257,N_683,N_1326);
or U8258 (N_8258,N_1663,N_1284);
xor U8259 (N_8259,N_3039,N_31);
or U8260 (N_8260,N_893,N_4027);
or U8261 (N_8261,N_2942,N_2948);
or U8262 (N_8262,N_2086,N_2638);
or U8263 (N_8263,N_769,N_1321);
nor U8264 (N_8264,N_4670,N_3352);
nor U8265 (N_8265,N_2767,N_2558);
xor U8266 (N_8266,N_795,N_2460);
or U8267 (N_8267,N_2643,N_3246);
nand U8268 (N_8268,N_4886,N_1570);
or U8269 (N_8269,N_479,N_2780);
and U8270 (N_8270,N_2477,N_1020);
nor U8271 (N_8271,N_4025,N_4410);
and U8272 (N_8272,N_307,N_1695);
xor U8273 (N_8273,N_4935,N_4254);
nor U8274 (N_8274,N_523,N_1013);
xnor U8275 (N_8275,N_2465,N_4828);
xnor U8276 (N_8276,N_3729,N_1585);
nand U8277 (N_8277,N_2997,N_4237);
and U8278 (N_8278,N_770,N_2403);
xor U8279 (N_8279,N_2507,N_3515);
nand U8280 (N_8280,N_2491,N_2605);
and U8281 (N_8281,N_3146,N_100);
nor U8282 (N_8282,N_986,N_4656);
nor U8283 (N_8283,N_1063,N_1995);
and U8284 (N_8284,N_3272,N_8);
and U8285 (N_8285,N_3202,N_399);
nor U8286 (N_8286,N_3380,N_4728);
nand U8287 (N_8287,N_4609,N_2638);
and U8288 (N_8288,N_3937,N_2637);
nand U8289 (N_8289,N_2666,N_3654);
xnor U8290 (N_8290,N_2277,N_404);
and U8291 (N_8291,N_1320,N_4543);
or U8292 (N_8292,N_4626,N_346);
nand U8293 (N_8293,N_4198,N_1269);
and U8294 (N_8294,N_3916,N_3881);
xor U8295 (N_8295,N_559,N_2306);
xnor U8296 (N_8296,N_3476,N_911);
nor U8297 (N_8297,N_2053,N_785);
nand U8298 (N_8298,N_1452,N_3582);
xor U8299 (N_8299,N_604,N_559);
nor U8300 (N_8300,N_3117,N_3786);
or U8301 (N_8301,N_103,N_2686);
xnor U8302 (N_8302,N_182,N_3227);
nand U8303 (N_8303,N_155,N_732);
nand U8304 (N_8304,N_1990,N_1437);
xor U8305 (N_8305,N_8,N_4745);
or U8306 (N_8306,N_1808,N_2979);
nand U8307 (N_8307,N_1808,N_2736);
or U8308 (N_8308,N_781,N_1168);
xor U8309 (N_8309,N_4850,N_4114);
nor U8310 (N_8310,N_1648,N_4119);
nor U8311 (N_8311,N_2964,N_975);
xor U8312 (N_8312,N_4961,N_29);
and U8313 (N_8313,N_4583,N_1518);
nor U8314 (N_8314,N_413,N_2804);
or U8315 (N_8315,N_4167,N_3273);
xor U8316 (N_8316,N_4265,N_2659);
nand U8317 (N_8317,N_1356,N_2962);
and U8318 (N_8318,N_3072,N_1956);
nor U8319 (N_8319,N_133,N_1518);
or U8320 (N_8320,N_3513,N_4483);
and U8321 (N_8321,N_4170,N_3456);
or U8322 (N_8322,N_4493,N_3122);
and U8323 (N_8323,N_3511,N_3077);
xnor U8324 (N_8324,N_2577,N_4045);
nand U8325 (N_8325,N_4561,N_1377);
nand U8326 (N_8326,N_4297,N_1459);
nor U8327 (N_8327,N_2057,N_382);
nand U8328 (N_8328,N_702,N_716);
nand U8329 (N_8329,N_1899,N_1662);
nand U8330 (N_8330,N_4085,N_4353);
or U8331 (N_8331,N_2851,N_2672);
and U8332 (N_8332,N_2247,N_1659);
and U8333 (N_8333,N_859,N_154);
nand U8334 (N_8334,N_737,N_4551);
xnor U8335 (N_8335,N_4661,N_316);
xor U8336 (N_8336,N_391,N_2382);
and U8337 (N_8337,N_4869,N_1684);
nand U8338 (N_8338,N_3421,N_88);
or U8339 (N_8339,N_1373,N_3140);
or U8340 (N_8340,N_130,N_2517);
nor U8341 (N_8341,N_719,N_1474);
or U8342 (N_8342,N_3502,N_975);
xor U8343 (N_8343,N_4284,N_4489);
and U8344 (N_8344,N_2807,N_1840);
xor U8345 (N_8345,N_3943,N_1078);
and U8346 (N_8346,N_395,N_4992);
xor U8347 (N_8347,N_4952,N_2935);
and U8348 (N_8348,N_407,N_2015);
and U8349 (N_8349,N_1756,N_2067);
xnor U8350 (N_8350,N_166,N_815);
nand U8351 (N_8351,N_3925,N_2704);
or U8352 (N_8352,N_4848,N_553);
nand U8353 (N_8353,N_479,N_4760);
xor U8354 (N_8354,N_3060,N_4544);
nor U8355 (N_8355,N_4503,N_4350);
or U8356 (N_8356,N_2231,N_854);
nand U8357 (N_8357,N_996,N_4594);
nor U8358 (N_8358,N_2339,N_4181);
and U8359 (N_8359,N_1190,N_2133);
nor U8360 (N_8360,N_1916,N_1495);
xor U8361 (N_8361,N_3692,N_71);
nand U8362 (N_8362,N_1508,N_3756);
xor U8363 (N_8363,N_3749,N_2135);
nor U8364 (N_8364,N_3452,N_4147);
and U8365 (N_8365,N_4882,N_660);
and U8366 (N_8366,N_4053,N_464);
and U8367 (N_8367,N_3311,N_2444);
or U8368 (N_8368,N_3202,N_4237);
xnor U8369 (N_8369,N_4849,N_3437);
or U8370 (N_8370,N_1178,N_2141);
nor U8371 (N_8371,N_4298,N_3088);
or U8372 (N_8372,N_212,N_4019);
xnor U8373 (N_8373,N_681,N_4769);
and U8374 (N_8374,N_4551,N_674);
xnor U8375 (N_8375,N_418,N_4685);
xnor U8376 (N_8376,N_4818,N_1046);
or U8377 (N_8377,N_2977,N_2130);
and U8378 (N_8378,N_1175,N_470);
nand U8379 (N_8379,N_258,N_3210);
or U8380 (N_8380,N_3200,N_1529);
and U8381 (N_8381,N_526,N_681);
and U8382 (N_8382,N_397,N_862);
and U8383 (N_8383,N_3654,N_2502);
nor U8384 (N_8384,N_4030,N_4477);
nor U8385 (N_8385,N_3382,N_224);
or U8386 (N_8386,N_835,N_2068);
xnor U8387 (N_8387,N_4029,N_993);
and U8388 (N_8388,N_3638,N_3456);
or U8389 (N_8389,N_3718,N_4232);
nor U8390 (N_8390,N_4816,N_92);
xnor U8391 (N_8391,N_2021,N_4469);
xnor U8392 (N_8392,N_3782,N_3182);
xnor U8393 (N_8393,N_3996,N_1093);
xnor U8394 (N_8394,N_3621,N_2087);
or U8395 (N_8395,N_1968,N_273);
nor U8396 (N_8396,N_2989,N_3378);
and U8397 (N_8397,N_3492,N_816);
and U8398 (N_8398,N_2022,N_4489);
nand U8399 (N_8399,N_176,N_2643);
and U8400 (N_8400,N_1359,N_2997);
nand U8401 (N_8401,N_3033,N_2501);
nor U8402 (N_8402,N_740,N_385);
or U8403 (N_8403,N_2652,N_2184);
and U8404 (N_8404,N_1720,N_1732);
and U8405 (N_8405,N_3563,N_3355);
or U8406 (N_8406,N_2242,N_2559);
nand U8407 (N_8407,N_1623,N_4095);
or U8408 (N_8408,N_1603,N_2860);
nand U8409 (N_8409,N_721,N_2477);
xor U8410 (N_8410,N_2566,N_275);
xor U8411 (N_8411,N_3689,N_3042);
nor U8412 (N_8412,N_3291,N_16);
and U8413 (N_8413,N_512,N_1644);
or U8414 (N_8414,N_3497,N_1103);
nand U8415 (N_8415,N_350,N_817);
nand U8416 (N_8416,N_100,N_2106);
or U8417 (N_8417,N_4913,N_4436);
or U8418 (N_8418,N_2422,N_789);
nor U8419 (N_8419,N_206,N_2637);
nor U8420 (N_8420,N_1582,N_4507);
or U8421 (N_8421,N_922,N_3539);
xor U8422 (N_8422,N_4687,N_3316);
and U8423 (N_8423,N_2522,N_2077);
and U8424 (N_8424,N_1439,N_550);
or U8425 (N_8425,N_4593,N_4223);
nand U8426 (N_8426,N_1459,N_2201);
xor U8427 (N_8427,N_4360,N_718);
xnor U8428 (N_8428,N_2983,N_434);
xor U8429 (N_8429,N_3245,N_1852);
nor U8430 (N_8430,N_65,N_4843);
nor U8431 (N_8431,N_3405,N_2646);
xnor U8432 (N_8432,N_2545,N_2254);
nor U8433 (N_8433,N_889,N_3075);
or U8434 (N_8434,N_4860,N_4020);
xnor U8435 (N_8435,N_4286,N_2225);
or U8436 (N_8436,N_270,N_3773);
nor U8437 (N_8437,N_4208,N_436);
and U8438 (N_8438,N_1475,N_3517);
and U8439 (N_8439,N_2244,N_1066);
or U8440 (N_8440,N_4374,N_2441);
and U8441 (N_8441,N_2272,N_1022);
xnor U8442 (N_8442,N_4919,N_147);
nand U8443 (N_8443,N_141,N_1534);
or U8444 (N_8444,N_2852,N_4899);
or U8445 (N_8445,N_745,N_3216);
nor U8446 (N_8446,N_4180,N_2229);
xnor U8447 (N_8447,N_1377,N_4027);
and U8448 (N_8448,N_1396,N_1145);
and U8449 (N_8449,N_802,N_4850);
and U8450 (N_8450,N_2157,N_1673);
xor U8451 (N_8451,N_261,N_2364);
nor U8452 (N_8452,N_1214,N_1198);
and U8453 (N_8453,N_229,N_4138);
xor U8454 (N_8454,N_1302,N_4944);
nor U8455 (N_8455,N_2024,N_4249);
xnor U8456 (N_8456,N_1140,N_4039);
nor U8457 (N_8457,N_3837,N_1134);
and U8458 (N_8458,N_660,N_1017);
nand U8459 (N_8459,N_1723,N_2059);
xor U8460 (N_8460,N_2428,N_3928);
nand U8461 (N_8461,N_3991,N_4563);
and U8462 (N_8462,N_171,N_2643);
or U8463 (N_8463,N_2059,N_527);
nor U8464 (N_8464,N_491,N_3898);
or U8465 (N_8465,N_4585,N_2876);
nor U8466 (N_8466,N_46,N_3785);
and U8467 (N_8467,N_960,N_4305);
nor U8468 (N_8468,N_3023,N_3085);
nor U8469 (N_8469,N_4650,N_3565);
nor U8470 (N_8470,N_2030,N_4033);
xor U8471 (N_8471,N_830,N_2137);
or U8472 (N_8472,N_4993,N_479);
or U8473 (N_8473,N_3701,N_2026);
nor U8474 (N_8474,N_2761,N_1983);
xor U8475 (N_8475,N_2585,N_2439);
xnor U8476 (N_8476,N_569,N_4571);
nor U8477 (N_8477,N_16,N_535);
xor U8478 (N_8478,N_3394,N_1995);
xnor U8479 (N_8479,N_3221,N_1133);
or U8480 (N_8480,N_3230,N_2532);
or U8481 (N_8481,N_333,N_3863);
nand U8482 (N_8482,N_2360,N_2678);
nand U8483 (N_8483,N_4970,N_49);
or U8484 (N_8484,N_2082,N_4672);
nor U8485 (N_8485,N_2487,N_1297);
or U8486 (N_8486,N_1806,N_2665);
xor U8487 (N_8487,N_2493,N_4198);
or U8488 (N_8488,N_284,N_3426);
nor U8489 (N_8489,N_993,N_4236);
or U8490 (N_8490,N_2741,N_3561);
nor U8491 (N_8491,N_2621,N_3015);
or U8492 (N_8492,N_224,N_3745);
and U8493 (N_8493,N_4094,N_2958);
nor U8494 (N_8494,N_1276,N_2687);
and U8495 (N_8495,N_3184,N_4346);
or U8496 (N_8496,N_3604,N_2796);
and U8497 (N_8497,N_2579,N_3217);
or U8498 (N_8498,N_4876,N_3868);
xnor U8499 (N_8499,N_1198,N_4737);
and U8500 (N_8500,N_2747,N_3438);
nand U8501 (N_8501,N_3094,N_3467);
xor U8502 (N_8502,N_2991,N_80);
xnor U8503 (N_8503,N_4979,N_1350);
and U8504 (N_8504,N_107,N_1189);
xor U8505 (N_8505,N_4211,N_3272);
xnor U8506 (N_8506,N_3831,N_1011);
nand U8507 (N_8507,N_4309,N_1730);
xor U8508 (N_8508,N_3378,N_1086);
nand U8509 (N_8509,N_3120,N_3898);
xor U8510 (N_8510,N_2638,N_2162);
and U8511 (N_8511,N_1043,N_2458);
nand U8512 (N_8512,N_4860,N_4197);
or U8513 (N_8513,N_4224,N_622);
nand U8514 (N_8514,N_3342,N_3780);
or U8515 (N_8515,N_4063,N_1931);
and U8516 (N_8516,N_2489,N_2626);
or U8517 (N_8517,N_861,N_4188);
nand U8518 (N_8518,N_3040,N_2742);
nand U8519 (N_8519,N_222,N_1665);
or U8520 (N_8520,N_1914,N_3422);
nand U8521 (N_8521,N_3748,N_3002);
or U8522 (N_8522,N_1993,N_171);
xnor U8523 (N_8523,N_313,N_4049);
xor U8524 (N_8524,N_2785,N_547);
or U8525 (N_8525,N_1491,N_232);
nand U8526 (N_8526,N_2117,N_4190);
nor U8527 (N_8527,N_4432,N_1877);
nor U8528 (N_8528,N_1145,N_4813);
nor U8529 (N_8529,N_2181,N_1262);
xor U8530 (N_8530,N_4839,N_2339);
and U8531 (N_8531,N_2448,N_1857);
nor U8532 (N_8532,N_2618,N_3937);
or U8533 (N_8533,N_4610,N_1896);
nand U8534 (N_8534,N_2874,N_2531);
nand U8535 (N_8535,N_1190,N_281);
nor U8536 (N_8536,N_252,N_61);
xor U8537 (N_8537,N_93,N_4826);
nand U8538 (N_8538,N_3501,N_3332);
nor U8539 (N_8539,N_311,N_865);
or U8540 (N_8540,N_2730,N_3872);
or U8541 (N_8541,N_4078,N_1126);
and U8542 (N_8542,N_2429,N_234);
nand U8543 (N_8543,N_4654,N_4674);
nand U8544 (N_8544,N_2279,N_2958);
nand U8545 (N_8545,N_2980,N_588);
and U8546 (N_8546,N_3080,N_3919);
and U8547 (N_8547,N_4148,N_3144);
xor U8548 (N_8548,N_129,N_2596);
and U8549 (N_8549,N_845,N_3912);
or U8550 (N_8550,N_472,N_2830);
nand U8551 (N_8551,N_2493,N_399);
and U8552 (N_8552,N_2532,N_2008);
nand U8553 (N_8553,N_1563,N_779);
and U8554 (N_8554,N_3091,N_2004);
or U8555 (N_8555,N_3810,N_4184);
or U8556 (N_8556,N_1148,N_209);
nor U8557 (N_8557,N_3635,N_605);
and U8558 (N_8558,N_997,N_2107);
and U8559 (N_8559,N_4519,N_179);
xor U8560 (N_8560,N_1666,N_29);
nand U8561 (N_8561,N_1630,N_556);
or U8562 (N_8562,N_353,N_2353);
or U8563 (N_8563,N_2996,N_741);
xor U8564 (N_8564,N_3820,N_2017);
nand U8565 (N_8565,N_1518,N_1171);
and U8566 (N_8566,N_1667,N_3886);
xor U8567 (N_8567,N_143,N_3314);
or U8568 (N_8568,N_923,N_2097);
or U8569 (N_8569,N_2,N_1888);
nand U8570 (N_8570,N_2214,N_3618);
nor U8571 (N_8571,N_1904,N_2517);
nor U8572 (N_8572,N_3320,N_2100);
nand U8573 (N_8573,N_3740,N_1659);
or U8574 (N_8574,N_4392,N_2968);
xor U8575 (N_8575,N_1366,N_4913);
or U8576 (N_8576,N_4055,N_1922);
and U8577 (N_8577,N_3375,N_4073);
and U8578 (N_8578,N_3328,N_296);
nor U8579 (N_8579,N_3221,N_424);
nor U8580 (N_8580,N_3568,N_3314);
nor U8581 (N_8581,N_3156,N_1117);
nand U8582 (N_8582,N_3158,N_4431);
or U8583 (N_8583,N_4676,N_3327);
xnor U8584 (N_8584,N_2622,N_4473);
and U8585 (N_8585,N_3674,N_4934);
xnor U8586 (N_8586,N_4988,N_325);
or U8587 (N_8587,N_3430,N_2874);
nor U8588 (N_8588,N_3816,N_2123);
xor U8589 (N_8589,N_623,N_1820);
or U8590 (N_8590,N_806,N_4427);
nand U8591 (N_8591,N_1362,N_2859);
xor U8592 (N_8592,N_1755,N_3669);
xor U8593 (N_8593,N_3830,N_3167);
or U8594 (N_8594,N_4103,N_2778);
or U8595 (N_8595,N_4716,N_3731);
xnor U8596 (N_8596,N_674,N_4454);
xnor U8597 (N_8597,N_497,N_3840);
nand U8598 (N_8598,N_1605,N_3928);
nand U8599 (N_8599,N_4360,N_2874);
nand U8600 (N_8600,N_1348,N_4934);
nand U8601 (N_8601,N_2733,N_2378);
nor U8602 (N_8602,N_3083,N_466);
and U8603 (N_8603,N_2219,N_4193);
or U8604 (N_8604,N_768,N_920);
nand U8605 (N_8605,N_3845,N_3592);
and U8606 (N_8606,N_1736,N_3322);
or U8607 (N_8607,N_3971,N_2467);
nor U8608 (N_8608,N_3428,N_4382);
or U8609 (N_8609,N_1529,N_3825);
and U8610 (N_8610,N_3433,N_3815);
nand U8611 (N_8611,N_4224,N_4095);
and U8612 (N_8612,N_4538,N_4183);
xor U8613 (N_8613,N_2352,N_2433);
nor U8614 (N_8614,N_1066,N_2038);
nand U8615 (N_8615,N_2503,N_2182);
nor U8616 (N_8616,N_3327,N_1447);
and U8617 (N_8617,N_1726,N_4884);
nor U8618 (N_8618,N_3224,N_2001);
nand U8619 (N_8619,N_2178,N_4612);
xor U8620 (N_8620,N_3263,N_979);
or U8621 (N_8621,N_1390,N_475);
and U8622 (N_8622,N_4356,N_1769);
nor U8623 (N_8623,N_3624,N_4411);
and U8624 (N_8624,N_2625,N_4245);
nand U8625 (N_8625,N_3745,N_3208);
or U8626 (N_8626,N_967,N_1824);
and U8627 (N_8627,N_4066,N_4541);
xnor U8628 (N_8628,N_2108,N_4967);
and U8629 (N_8629,N_4686,N_1389);
nand U8630 (N_8630,N_3915,N_1073);
nor U8631 (N_8631,N_2402,N_819);
xor U8632 (N_8632,N_1587,N_415);
xor U8633 (N_8633,N_2235,N_3776);
or U8634 (N_8634,N_59,N_689);
and U8635 (N_8635,N_1245,N_4388);
nand U8636 (N_8636,N_4942,N_4213);
and U8637 (N_8637,N_406,N_1959);
nor U8638 (N_8638,N_699,N_2361);
and U8639 (N_8639,N_3354,N_3162);
and U8640 (N_8640,N_1666,N_1570);
nand U8641 (N_8641,N_3629,N_1462);
and U8642 (N_8642,N_3805,N_3808);
or U8643 (N_8643,N_3363,N_3674);
nor U8644 (N_8644,N_1726,N_288);
nor U8645 (N_8645,N_464,N_247);
nor U8646 (N_8646,N_1993,N_3980);
and U8647 (N_8647,N_1059,N_2790);
nor U8648 (N_8648,N_2469,N_1029);
xnor U8649 (N_8649,N_1608,N_1579);
nor U8650 (N_8650,N_1195,N_3708);
xnor U8651 (N_8651,N_318,N_4625);
and U8652 (N_8652,N_1676,N_4122);
xnor U8653 (N_8653,N_293,N_4721);
nor U8654 (N_8654,N_685,N_1655);
nor U8655 (N_8655,N_4561,N_3633);
nor U8656 (N_8656,N_4855,N_2814);
nand U8657 (N_8657,N_3222,N_4467);
or U8658 (N_8658,N_2711,N_2247);
or U8659 (N_8659,N_362,N_4249);
nor U8660 (N_8660,N_2729,N_3215);
or U8661 (N_8661,N_1903,N_747);
or U8662 (N_8662,N_2105,N_1666);
or U8663 (N_8663,N_2385,N_1468);
xor U8664 (N_8664,N_3165,N_4029);
nor U8665 (N_8665,N_2667,N_2093);
and U8666 (N_8666,N_2164,N_4776);
xnor U8667 (N_8667,N_718,N_2164);
and U8668 (N_8668,N_1720,N_1243);
xnor U8669 (N_8669,N_1772,N_3426);
nor U8670 (N_8670,N_4007,N_1556);
xnor U8671 (N_8671,N_2960,N_356);
nand U8672 (N_8672,N_603,N_2838);
nor U8673 (N_8673,N_2561,N_2580);
or U8674 (N_8674,N_3816,N_311);
or U8675 (N_8675,N_2274,N_2078);
nand U8676 (N_8676,N_4592,N_4380);
or U8677 (N_8677,N_4273,N_3789);
nor U8678 (N_8678,N_3865,N_4131);
xnor U8679 (N_8679,N_4135,N_2690);
or U8680 (N_8680,N_204,N_703);
nor U8681 (N_8681,N_3069,N_1658);
nor U8682 (N_8682,N_197,N_2266);
or U8683 (N_8683,N_3780,N_4729);
and U8684 (N_8684,N_2405,N_1981);
nor U8685 (N_8685,N_1054,N_2340);
or U8686 (N_8686,N_737,N_1138);
xor U8687 (N_8687,N_2,N_3223);
xor U8688 (N_8688,N_3260,N_4145);
and U8689 (N_8689,N_4925,N_4327);
and U8690 (N_8690,N_1913,N_3080);
and U8691 (N_8691,N_1204,N_4956);
or U8692 (N_8692,N_2604,N_4646);
and U8693 (N_8693,N_4485,N_82);
nand U8694 (N_8694,N_2986,N_3865);
or U8695 (N_8695,N_1289,N_2161);
nor U8696 (N_8696,N_3301,N_4825);
nand U8697 (N_8697,N_4279,N_1057);
nand U8698 (N_8698,N_1304,N_4336);
xnor U8699 (N_8699,N_2266,N_1159);
nand U8700 (N_8700,N_1502,N_420);
and U8701 (N_8701,N_3586,N_2109);
xor U8702 (N_8702,N_4112,N_2683);
or U8703 (N_8703,N_404,N_4705);
xor U8704 (N_8704,N_3305,N_1079);
and U8705 (N_8705,N_3379,N_3099);
and U8706 (N_8706,N_54,N_4244);
xnor U8707 (N_8707,N_4541,N_2324);
and U8708 (N_8708,N_51,N_1638);
xnor U8709 (N_8709,N_3661,N_2621);
nor U8710 (N_8710,N_4124,N_3133);
or U8711 (N_8711,N_4029,N_2318);
nor U8712 (N_8712,N_3313,N_1664);
nor U8713 (N_8713,N_1587,N_889);
nor U8714 (N_8714,N_4508,N_3639);
and U8715 (N_8715,N_2429,N_1412);
and U8716 (N_8716,N_4899,N_214);
and U8717 (N_8717,N_251,N_4788);
and U8718 (N_8718,N_1776,N_2838);
or U8719 (N_8719,N_4811,N_3344);
nand U8720 (N_8720,N_977,N_3502);
nor U8721 (N_8721,N_687,N_1026);
nor U8722 (N_8722,N_2494,N_77);
or U8723 (N_8723,N_1342,N_2576);
nand U8724 (N_8724,N_941,N_1362);
nor U8725 (N_8725,N_2033,N_2525);
nand U8726 (N_8726,N_2979,N_2136);
or U8727 (N_8727,N_2042,N_1066);
and U8728 (N_8728,N_2296,N_1469);
and U8729 (N_8729,N_1778,N_419);
and U8730 (N_8730,N_2540,N_3709);
and U8731 (N_8731,N_4512,N_588);
or U8732 (N_8732,N_4399,N_881);
xor U8733 (N_8733,N_558,N_2152);
or U8734 (N_8734,N_2851,N_2015);
xor U8735 (N_8735,N_4750,N_2676);
nand U8736 (N_8736,N_3160,N_4902);
and U8737 (N_8737,N_684,N_186);
and U8738 (N_8738,N_4679,N_1266);
nor U8739 (N_8739,N_350,N_1107);
nor U8740 (N_8740,N_479,N_1559);
or U8741 (N_8741,N_2799,N_1135);
xor U8742 (N_8742,N_1169,N_2071);
and U8743 (N_8743,N_1074,N_3885);
xor U8744 (N_8744,N_4914,N_3933);
and U8745 (N_8745,N_3442,N_295);
or U8746 (N_8746,N_3860,N_2371);
or U8747 (N_8747,N_4018,N_718);
xor U8748 (N_8748,N_1573,N_2086);
or U8749 (N_8749,N_20,N_2836);
and U8750 (N_8750,N_4734,N_3475);
and U8751 (N_8751,N_881,N_1831);
nor U8752 (N_8752,N_4345,N_1975);
nor U8753 (N_8753,N_3906,N_4371);
or U8754 (N_8754,N_2636,N_443);
nor U8755 (N_8755,N_1741,N_1996);
or U8756 (N_8756,N_3714,N_3301);
xor U8757 (N_8757,N_2617,N_2879);
and U8758 (N_8758,N_3882,N_4725);
xnor U8759 (N_8759,N_343,N_1490);
xor U8760 (N_8760,N_1936,N_4507);
or U8761 (N_8761,N_3696,N_4067);
nor U8762 (N_8762,N_350,N_3483);
or U8763 (N_8763,N_1199,N_4408);
and U8764 (N_8764,N_2163,N_3509);
or U8765 (N_8765,N_573,N_2170);
nand U8766 (N_8766,N_976,N_15);
or U8767 (N_8767,N_2453,N_1562);
nor U8768 (N_8768,N_420,N_63);
nand U8769 (N_8769,N_1677,N_3762);
or U8770 (N_8770,N_721,N_1475);
and U8771 (N_8771,N_2352,N_1261);
xnor U8772 (N_8772,N_4711,N_1114);
xor U8773 (N_8773,N_1600,N_2951);
or U8774 (N_8774,N_366,N_2866);
xnor U8775 (N_8775,N_3945,N_2430);
nand U8776 (N_8776,N_391,N_663);
and U8777 (N_8777,N_938,N_186);
nand U8778 (N_8778,N_51,N_1409);
xnor U8779 (N_8779,N_3436,N_2454);
nand U8780 (N_8780,N_4271,N_1000);
nand U8781 (N_8781,N_2577,N_773);
and U8782 (N_8782,N_1546,N_67);
nor U8783 (N_8783,N_4170,N_4137);
nor U8784 (N_8784,N_4303,N_967);
or U8785 (N_8785,N_3059,N_319);
nand U8786 (N_8786,N_2697,N_2684);
nand U8787 (N_8787,N_2932,N_522);
and U8788 (N_8788,N_3982,N_3078);
nor U8789 (N_8789,N_1985,N_2644);
nor U8790 (N_8790,N_26,N_4895);
or U8791 (N_8791,N_4924,N_4798);
nand U8792 (N_8792,N_4547,N_3721);
nand U8793 (N_8793,N_2614,N_3471);
and U8794 (N_8794,N_3775,N_457);
nor U8795 (N_8795,N_3867,N_183);
nand U8796 (N_8796,N_1271,N_2322);
nor U8797 (N_8797,N_3559,N_527);
and U8798 (N_8798,N_1037,N_2913);
xor U8799 (N_8799,N_619,N_32);
nor U8800 (N_8800,N_4483,N_3531);
or U8801 (N_8801,N_1106,N_315);
and U8802 (N_8802,N_1684,N_2727);
xnor U8803 (N_8803,N_4164,N_4718);
xnor U8804 (N_8804,N_1475,N_529);
and U8805 (N_8805,N_4785,N_4878);
and U8806 (N_8806,N_1851,N_418);
and U8807 (N_8807,N_1984,N_4674);
xnor U8808 (N_8808,N_3259,N_4880);
or U8809 (N_8809,N_2595,N_3979);
and U8810 (N_8810,N_219,N_1134);
xnor U8811 (N_8811,N_3638,N_2823);
and U8812 (N_8812,N_2159,N_774);
nand U8813 (N_8813,N_357,N_600);
nor U8814 (N_8814,N_190,N_2752);
nand U8815 (N_8815,N_2831,N_29);
nor U8816 (N_8816,N_1181,N_1543);
and U8817 (N_8817,N_2615,N_2487);
and U8818 (N_8818,N_14,N_1623);
xnor U8819 (N_8819,N_935,N_3338);
and U8820 (N_8820,N_435,N_3104);
or U8821 (N_8821,N_469,N_4200);
nor U8822 (N_8822,N_4466,N_4612);
nand U8823 (N_8823,N_378,N_1509);
or U8824 (N_8824,N_3621,N_609);
nand U8825 (N_8825,N_1039,N_3469);
nand U8826 (N_8826,N_3413,N_223);
xnor U8827 (N_8827,N_4943,N_909);
or U8828 (N_8828,N_2677,N_1068);
nor U8829 (N_8829,N_3110,N_2278);
and U8830 (N_8830,N_2316,N_3697);
nand U8831 (N_8831,N_2925,N_2027);
and U8832 (N_8832,N_2600,N_3128);
nand U8833 (N_8833,N_1000,N_2579);
xnor U8834 (N_8834,N_4217,N_1056);
nand U8835 (N_8835,N_4859,N_4799);
xnor U8836 (N_8836,N_3475,N_36);
xor U8837 (N_8837,N_4252,N_1980);
and U8838 (N_8838,N_3398,N_3554);
nand U8839 (N_8839,N_3563,N_2392);
xor U8840 (N_8840,N_2487,N_4141);
xor U8841 (N_8841,N_3318,N_2212);
and U8842 (N_8842,N_3507,N_532);
and U8843 (N_8843,N_4497,N_1107);
xnor U8844 (N_8844,N_4268,N_4442);
xor U8845 (N_8845,N_4317,N_1630);
nor U8846 (N_8846,N_3216,N_1634);
and U8847 (N_8847,N_1268,N_766);
nor U8848 (N_8848,N_2303,N_1379);
or U8849 (N_8849,N_1074,N_1635);
nor U8850 (N_8850,N_1120,N_2760);
xnor U8851 (N_8851,N_2356,N_317);
xor U8852 (N_8852,N_3525,N_2071);
nor U8853 (N_8853,N_4629,N_4342);
or U8854 (N_8854,N_350,N_1725);
and U8855 (N_8855,N_2991,N_1095);
nand U8856 (N_8856,N_1802,N_4896);
and U8857 (N_8857,N_4529,N_1084);
or U8858 (N_8858,N_3592,N_4259);
nand U8859 (N_8859,N_868,N_3283);
and U8860 (N_8860,N_2013,N_1836);
or U8861 (N_8861,N_4875,N_546);
xor U8862 (N_8862,N_1692,N_2025);
xor U8863 (N_8863,N_1800,N_2742);
xor U8864 (N_8864,N_2115,N_3289);
nor U8865 (N_8865,N_926,N_4497);
nor U8866 (N_8866,N_1881,N_4328);
nand U8867 (N_8867,N_4314,N_4481);
xnor U8868 (N_8868,N_3456,N_1480);
nor U8869 (N_8869,N_206,N_1239);
and U8870 (N_8870,N_3375,N_2506);
or U8871 (N_8871,N_3734,N_2714);
or U8872 (N_8872,N_3179,N_724);
xnor U8873 (N_8873,N_998,N_1059);
nand U8874 (N_8874,N_3335,N_3989);
nor U8875 (N_8875,N_1445,N_2294);
nor U8876 (N_8876,N_3378,N_4799);
or U8877 (N_8877,N_4352,N_510);
and U8878 (N_8878,N_679,N_1518);
and U8879 (N_8879,N_684,N_1972);
nand U8880 (N_8880,N_796,N_2354);
and U8881 (N_8881,N_2512,N_2958);
xor U8882 (N_8882,N_275,N_2316);
nor U8883 (N_8883,N_426,N_3622);
or U8884 (N_8884,N_725,N_2166);
or U8885 (N_8885,N_346,N_2077);
or U8886 (N_8886,N_913,N_4161);
nand U8887 (N_8887,N_162,N_3840);
nand U8888 (N_8888,N_619,N_4415);
xor U8889 (N_8889,N_3143,N_1837);
nand U8890 (N_8890,N_765,N_2679);
or U8891 (N_8891,N_3286,N_1519);
xnor U8892 (N_8892,N_185,N_981);
xnor U8893 (N_8893,N_3987,N_2362);
xnor U8894 (N_8894,N_2629,N_3976);
nor U8895 (N_8895,N_3894,N_1793);
nor U8896 (N_8896,N_4684,N_3556);
xnor U8897 (N_8897,N_2460,N_3616);
nor U8898 (N_8898,N_1721,N_3240);
nor U8899 (N_8899,N_1899,N_2322);
xor U8900 (N_8900,N_3266,N_4195);
or U8901 (N_8901,N_642,N_3736);
and U8902 (N_8902,N_1089,N_673);
nor U8903 (N_8903,N_1894,N_1453);
and U8904 (N_8904,N_3589,N_4920);
or U8905 (N_8905,N_2463,N_759);
nand U8906 (N_8906,N_1673,N_915);
and U8907 (N_8907,N_2561,N_3490);
and U8908 (N_8908,N_4963,N_1968);
xnor U8909 (N_8909,N_350,N_4835);
xor U8910 (N_8910,N_3286,N_356);
nor U8911 (N_8911,N_882,N_2776);
nand U8912 (N_8912,N_1942,N_151);
nand U8913 (N_8913,N_1881,N_1432);
or U8914 (N_8914,N_4688,N_1318);
xor U8915 (N_8915,N_3659,N_3660);
nor U8916 (N_8916,N_4104,N_3026);
and U8917 (N_8917,N_4928,N_2037);
or U8918 (N_8918,N_330,N_4966);
xnor U8919 (N_8919,N_933,N_3659);
xnor U8920 (N_8920,N_4247,N_4669);
nand U8921 (N_8921,N_3017,N_4610);
nor U8922 (N_8922,N_1747,N_3016);
or U8923 (N_8923,N_1552,N_1526);
nand U8924 (N_8924,N_2735,N_4352);
nor U8925 (N_8925,N_3889,N_157);
or U8926 (N_8926,N_4113,N_3502);
xnor U8927 (N_8927,N_798,N_326);
and U8928 (N_8928,N_2482,N_2818);
nand U8929 (N_8929,N_3093,N_543);
nand U8930 (N_8930,N_4817,N_1947);
or U8931 (N_8931,N_2674,N_1004);
and U8932 (N_8932,N_1208,N_1337);
nand U8933 (N_8933,N_2686,N_2986);
nor U8934 (N_8934,N_319,N_272);
and U8935 (N_8935,N_2912,N_1103);
nor U8936 (N_8936,N_4616,N_4835);
nor U8937 (N_8937,N_4417,N_1683);
nor U8938 (N_8938,N_2394,N_1310);
nand U8939 (N_8939,N_591,N_4463);
nand U8940 (N_8940,N_3260,N_840);
and U8941 (N_8941,N_391,N_1151);
nand U8942 (N_8942,N_3061,N_2084);
xor U8943 (N_8943,N_3151,N_4355);
nand U8944 (N_8944,N_4865,N_729);
xnor U8945 (N_8945,N_4798,N_4083);
nand U8946 (N_8946,N_704,N_4022);
xor U8947 (N_8947,N_3752,N_1520);
nand U8948 (N_8948,N_2249,N_2749);
or U8949 (N_8949,N_2953,N_597);
and U8950 (N_8950,N_1232,N_358);
and U8951 (N_8951,N_1744,N_141);
xor U8952 (N_8952,N_3060,N_4964);
xnor U8953 (N_8953,N_4627,N_114);
or U8954 (N_8954,N_561,N_3164);
and U8955 (N_8955,N_4919,N_2136);
nand U8956 (N_8956,N_1311,N_3401);
nand U8957 (N_8957,N_4194,N_2147);
nor U8958 (N_8958,N_4957,N_3515);
or U8959 (N_8959,N_1797,N_3103);
nand U8960 (N_8960,N_4947,N_947);
and U8961 (N_8961,N_1966,N_1003);
nor U8962 (N_8962,N_4278,N_1159);
xnor U8963 (N_8963,N_1808,N_3469);
nand U8964 (N_8964,N_2915,N_3820);
and U8965 (N_8965,N_891,N_3043);
xnor U8966 (N_8966,N_1516,N_2123);
or U8967 (N_8967,N_3745,N_2897);
xor U8968 (N_8968,N_4379,N_1880);
nand U8969 (N_8969,N_3210,N_4355);
nand U8970 (N_8970,N_483,N_1727);
nor U8971 (N_8971,N_4000,N_3136);
nand U8972 (N_8972,N_2821,N_3190);
nor U8973 (N_8973,N_1069,N_3564);
nor U8974 (N_8974,N_3613,N_1419);
nand U8975 (N_8975,N_2713,N_4590);
nor U8976 (N_8976,N_2191,N_1063);
or U8977 (N_8977,N_1405,N_4629);
nor U8978 (N_8978,N_289,N_2398);
xnor U8979 (N_8979,N_156,N_3669);
nand U8980 (N_8980,N_1525,N_4735);
nand U8981 (N_8981,N_1859,N_3154);
or U8982 (N_8982,N_560,N_394);
and U8983 (N_8983,N_1874,N_2162);
nor U8984 (N_8984,N_3533,N_4854);
nor U8985 (N_8985,N_2077,N_466);
or U8986 (N_8986,N_4859,N_1210);
nor U8987 (N_8987,N_3566,N_2184);
and U8988 (N_8988,N_3831,N_4834);
and U8989 (N_8989,N_2085,N_4107);
nand U8990 (N_8990,N_527,N_2602);
xor U8991 (N_8991,N_3878,N_1803);
nor U8992 (N_8992,N_3084,N_4359);
or U8993 (N_8993,N_111,N_2385);
or U8994 (N_8994,N_2258,N_2260);
nand U8995 (N_8995,N_435,N_60);
nand U8996 (N_8996,N_4199,N_4487);
and U8997 (N_8997,N_4125,N_3856);
nand U8998 (N_8998,N_2536,N_719);
xnor U8999 (N_8999,N_2456,N_487);
nand U9000 (N_9000,N_613,N_1385);
nand U9001 (N_9001,N_2370,N_1357);
and U9002 (N_9002,N_2885,N_4569);
and U9003 (N_9003,N_3451,N_4846);
and U9004 (N_9004,N_4460,N_4207);
and U9005 (N_9005,N_2569,N_690);
xor U9006 (N_9006,N_3916,N_113);
or U9007 (N_9007,N_4440,N_1576);
and U9008 (N_9008,N_4161,N_809);
or U9009 (N_9009,N_2485,N_2087);
and U9010 (N_9010,N_4816,N_463);
xor U9011 (N_9011,N_2757,N_1362);
nor U9012 (N_9012,N_996,N_866);
nor U9013 (N_9013,N_4816,N_690);
xnor U9014 (N_9014,N_1014,N_2184);
xnor U9015 (N_9015,N_4067,N_1118);
nor U9016 (N_9016,N_521,N_1644);
nor U9017 (N_9017,N_956,N_3436);
nand U9018 (N_9018,N_424,N_1620);
nor U9019 (N_9019,N_2960,N_486);
nor U9020 (N_9020,N_580,N_2443);
nand U9021 (N_9021,N_3773,N_3822);
nor U9022 (N_9022,N_2381,N_3869);
or U9023 (N_9023,N_870,N_1797);
xnor U9024 (N_9024,N_1706,N_4503);
nor U9025 (N_9025,N_3717,N_4593);
or U9026 (N_9026,N_2388,N_942);
or U9027 (N_9027,N_2761,N_4923);
nor U9028 (N_9028,N_1232,N_2789);
xor U9029 (N_9029,N_2195,N_2697);
nor U9030 (N_9030,N_4085,N_1173);
and U9031 (N_9031,N_39,N_3478);
or U9032 (N_9032,N_4681,N_2235);
and U9033 (N_9033,N_518,N_498);
or U9034 (N_9034,N_2506,N_692);
and U9035 (N_9035,N_1731,N_3485);
or U9036 (N_9036,N_3472,N_4290);
xnor U9037 (N_9037,N_2344,N_875);
or U9038 (N_9038,N_378,N_2144);
and U9039 (N_9039,N_747,N_3366);
xnor U9040 (N_9040,N_3325,N_2912);
nand U9041 (N_9041,N_200,N_1078);
and U9042 (N_9042,N_3499,N_2743);
nand U9043 (N_9043,N_3829,N_2919);
xor U9044 (N_9044,N_3663,N_55);
nor U9045 (N_9045,N_1312,N_3522);
nor U9046 (N_9046,N_100,N_2922);
xor U9047 (N_9047,N_4346,N_4690);
nor U9048 (N_9048,N_343,N_4227);
nand U9049 (N_9049,N_1094,N_1864);
xnor U9050 (N_9050,N_3800,N_4138);
or U9051 (N_9051,N_236,N_2029);
xor U9052 (N_9052,N_444,N_58);
and U9053 (N_9053,N_2845,N_853);
or U9054 (N_9054,N_3489,N_2191);
nand U9055 (N_9055,N_4999,N_998);
and U9056 (N_9056,N_3523,N_1324);
nor U9057 (N_9057,N_422,N_3489);
nand U9058 (N_9058,N_3092,N_997);
nand U9059 (N_9059,N_2434,N_742);
or U9060 (N_9060,N_1751,N_4611);
xor U9061 (N_9061,N_1248,N_3577);
nand U9062 (N_9062,N_2091,N_1706);
xor U9063 (N_9063,N_1933,N_4618);
and U9064 (N_9064,N_51,N_4576);
and U9065 (N_9065,N_4578,N_4703);
or U9066 (N_9066,N_4959,N_3867);
or U9067 (N_9067,N_3370,N_1337);
nand U9068 (N_9068,N_4840,N_348);
nand U9069 (N_9069,N_1443,N_4448);
and U9070 (N_9070,N_105,N_156);
and U9071 (N_9071,N_287,N_1867);
nor U9072 (N_9072,N_4175,N_2566);
or U9073 (N_9073,N_1201,N_2982);
nor U9074 (N_9074,N_1972,N_260);
or U9075 (N_9075,N_4374,N_4093);
nand U9076 (N_9076,N_4132,N_3864);
nand U9077 (N_9077,N_126,N_1553);
nand U9078 (N_9078,N_2393,N_482);
xor U9079 (N_9079,N_137,N_4634);
xnor U9080 (N_9080,N_4392,N_2521);
nor U9081 (N_9081,N_3854,N_4927);
xnor U9082 (N_9082,N_849,N_302);
or U9083 (N_9083,N_3895,N_4756);
xnor U9084 (N_9084,N_3047,N_1212);
or U9085 (N_9085,N_1352,N_1544);
and U9086 (N_9086,N_2171,N_1628);
nor U9087 (N_9087,N_331,N_1669);
nand U9088 (N_9088,N_3794,N_4520);
nor U9089 (N_9089,N_2968,N_1226);
nor U9090 (N_9090,N_3388,N_4374);
xor U9091 (N_9091,N_2522,N_3904);
nand U9092 (N_9092,N_674,N_4522);
or U9093 (N_9093,N_1852,N_950);
nor U9094 (N_9094,N_644,N_427);
nand U9095 (N_9095,N_1438,N_2118);
and U9096 (N_9096,N_91,N_2021);
nor U9097 (N_9097,N_5,N_153);
or U9098 (N_9098,N_4982,N_1742);
or U9099 (N_9099,N_2396,N_1453);
nand U9100 (N_9100,N_170,N_829);
and U9101 (N_9101,N_4317,N_3572);
nand U9102 (N_9102,N_1806,N_4451);
xor U9103 (N_9103,N_4069,N_1742);
or U9104 (N_9104,N_2762,N_247);
xor U9105 (N_9105,N_418,N_2939);
or U9106 (N_9106,N_4756,N_3665);
nor U9107 (N_9107,N_2594,N_1744);
xor U9108 (N_9108,N_2254,N_2776);
nor U9109 (N_9109,N_1721,N_2631);
and U9110 (N_9110,N_4175,N_3761);
nor U9111 (N_9111,N_4393,N_4043);
nand U9112 (N_9112,N_4485,N_492);
and U9113 (N_9113,N_4618,N_2269);
nor U9114 (N_9114,N_4652,N_1033);
nand U9115 (N_9115,N_1105,N_3553);
or U9116 (N_9116,N_319,N_1461);
or U9117 (N_9117,N_4605,N_2796);
xor U9118 (N_9118,N_4572,N_3091);
nand U9119 (N_9119,N_1572,N_4512);
or U9120 (N_9120,N_1746,N_428);
or U9121 (N_9121,N_1952,N_2422);
nand U9122 (N_9122,N_3265,N_2952);
nand U9123 (N_9123,N_174,N_2094);
xor U9124 (N_9124,N_972,N_1461);
and U9125 (N_9125,N_2357,N_1557);
or U9126 (N_9126,N_2532,N_298);
or U9127 (N_9127,N_86,N_3448);
and U9128 (N_9128,N_3901,N_3337);
nor U9129 (N_9129,N_2217,N_57);
and U9130 (N_9130,N_3265,N_4125);
nor U9131 (N_9131,N_1992,N_4670);
nand U9132 (N_9132,N_4912,N_988);
nand U9133 (N_9133,N_273,N_4924);
and U9134 (N_9134,N_737,N_1994);
nor U9135 (N_9135,N_3056,N_657);
xor U9136 (N_9136,N_193,N_1534);
nand U9137 (N_9137,N_1518,N_4156);
nand U9138 (N_9138,N_372,N_3990);
and U9139 (N_9139,N_549,N_4483);
nand U9140 (N_9140,N_1719,N_4092);
or U9141 (N_9141,N_1146,N_4221);
or U9142 (N_9142,N_1802,N_4829);
or U9143 (N_9143,N_958,N_1914);
nor U9144 (N_9144,N_2393,N_761);
nor U9145 (N_9145,N_1863,N_2578);
nor U9146 (N_9146,N_3344,N_3825);
nand U9147 (N_9147,N_2082,N_982);
or U9148 (N_9148,N_4576,N_1967);
xnor U9149 (N_9149,N_3659,N_3372);
or U9150 (N_9150,N_1295,N_704);
nand U9151 (N_9151,N_4612,N_1643);
nand U9152 (N_9152,N_1591,N_3869);
nand U9153 (N_9153,N_3161,N_1481);
and U9154 (N_9154,N_880,N_3978);
nand U9155 (N_9155,N_136,N_4293);
xnor U9156 (N_9156,N_97,N_3668);
or U9157 (N_9157,N_2972,N_394);
xnor U9158 (N_9158,N_3522,N_2636);
and U9159 (N_9159,N_1224,N_4808);
nand U9160 (N_9160,N_3789,N_3901);
nand U9161 (N_9161,N_30,N_4179);
xnor U9162 (N_9162,N_3855,N_3206);
or U9163 (N_9163,N_3017,N_3840);
and U9164 (N_9164,N_3129,N_4024);
and U9165 (N_9165,N_3060,N_200);
or U9166 (N_9166,N_2109,N_4745);
and U9167 (N_9167,N_796,N_2418);
nor U9168 (N_9168,N_3910,N_329);
nor U9169 (N_9169,N_2923,N_523);
xor U9170 (N_9170,N_936,N_3070);
or U9171 (N_9171,N_606,N_2791);
nor U9172 (N_9172,N_2219,N_2135);
xnor U9173 (N_9173,N_4912,N_794);
and U9174 (N_9174,N_1819,N_1138);
nor U9175 (N_9175,N_454,N_1119);
or U9176 (N_9176,N_916,N_3258);
nand U9177 (N_9177,N_2289,N_3214);
and U9178 (N_9178,N_4873,N_3182);
or U9179 (N_9179,N_11,N_574);
and U9180 (N_9180,N_3924,N_925);
nand U9181 (N_9181,N_3899,N_4887);
and U9182 (N_9182,N_1976,N_989);
and U9183 (N_9183,N_4502,N_353);
nor U9184 (N_9184,N_1389,N_3817);
xnor U9185 (N_9185,N_1329,N_2425);
or U9186 (N_9186,N_1473,N_2713);
or U9187 (N_9187,N_3776,N_987);
nor U9188 (N_9188,N_4685,N_2854);
and U9189 (N_9189,N_1017,N_1982);
nor U9190 (N_9190,N_3480,N_1852);
and U9191 (N_9191,N_4082,N_311);
nor U9192 (N_9192,N_2247,N_2231);
and U9193 (N_9193,N_80,N_850);
and U9194 (N_9194,N_3321,N_3858);
nor U9195 (N_9195,N_1420,N_4506);
nand U9196 (N_9196,N_1873,N_606);
nor U9197 (N_9197,N_281,N_4947);
nand U9198 (N_9198,N_4897,N_2673);
nand U9199 (N_9199,N_2901,N_1644);
nor U9200 (N_9200,N_3724,N_4657);
or U9201 (N_9201,N_896,N_129);
or U9202 (N_9202,N_1456,N_2350);
and U9203 (N_9203,N_3769,N_1499);
xor U9204 (N_9204,N_40,N_4773);
and U9205 (N_9205,N_3923,N_3799);
or U9206 (N_9206,N_4438,N_4655);
and U9207 (N_9207,N_1661,N_561);
or U9208 (N_9208,N_1518,N_4227);
nand U9209 (N_9209,N_2696,N_546);
nor U9210 (N_9210,N_591,N_1349);
xor U9211 (N_9211,N_4727,N_1690);
nand U9212 (N_9212,N_2398,N_2151);
nor U9213 (N_9213,N_1079,N_4277);
and U9214 (N_9214,N_2518,N_2343);
nand U9215 (N_9215,N_456,N_2898);
xor U9216 (N_9216,N_3411,N_4768);
xnor U9217 (N_9217,N_3681,N_4188);
nand U9218 (N_9218,N_3457,N_46);
nor U9219 (N_9219,N_4768,N_784);
nand U9220 (N_9220,N_3480,N_3426);
and U9221 (N_9221,N_2122,N_4022);
nor U9222 (N_9222,N_3463,N_1399);
or U9223 (N_9223,N_3129,N_4500);
and U9224 (N_9224,N_4393,N_4293);
nor U9225 (N_9225,N_4585,N_1950);
xnor U9226 (N_9226,N_187,N_1974);
nor U9227 (N_9227,N_2669,N_2573);
nand U9228 (N_9228,N_2804,N_133);
and U9229 (N_9229,N_4896,N_3818);
xnor U9230 (N_9230,N_2945,N_1615);
nor U9231 (N_9231,N_1684,N_3727);
and U9232 (N_9232,N_3947,N_568);
or U9233 (N_9233,N_3498,N_4664);
or U9234 (N_9234,N_1779,N_2173);
nand U9235 (N_9235,N_4949,N_835);
xnor U9236 (N_9236,N_4802,N_740);
nor U9237 (N_9237,N_2978,N_32);
and U9238 (N_9238,N_2599,N_1364);
xor U9239 (N_9239,N_693,N_4905);
and U9240 (N_9240,N_2587,N_3638);
nor U9241 (N_9241,N_1788,N_99);
or U9242 (N_9242,N_989,N_4400);
and U9243 (N_9243,N_969,N_4732);
or U9244 (N_9244,N_1028,N_1703);
xnor U9245 (N_9245,N_2378,N_569);
or U9246 (N_9246,N_1545,N_3359);
and U9247 (N_9247,N_4022,N_1167);
nor U9248 (N_9248,N_4168,N_66);
or U9249 (N_9249,N_3336,N_1064);
xnor U9250 (N_9250,N_1623,N_1285);
or U9251 (N_9251,N_4382,N_4374);
xor U9252 (N_9252,N_2331,N_1390);
nand U9253 (N_9253,N_573,N_2156);
nor U9254 (N_9254,N_40,N_4182);
xnor U9255 (N_9255,N_2235,N_1557);
or U9256 (N_9256,N_859,N_2989);
nor U9257 (N_9257,N_3909,N_3926);
and U9258 (N_9258,N_1545,N_2424);
nand U9259 (N_9259,N_3294,N_4297);
and U9260 (N_9260,N_295,N_4795);
nand U9261 (N_9261,N_1727,N_413);
or U9262 (N_9262,N_2717,N_2920);
and U9263 (N_9263,N_4302,N_294);
or U9264 (N_9264,N_3052,N_2140);
nor U9265 (N_9265,N_420,N_429);
nand U9266 (N_9266,N_4648,N_4350);
nor U9267 (N_9267,N_2939,N_3304);
xnor U9268 (N_9268,N_2883,N_2959);
nand U9269 (N_9269,N_3067,N_3221);
nor U9270 (N_9270,N_2860,N_1214);
xnor U9271 (N_9271,N_3611,N_1994);
nor U9272 (N_9272,N_1587,N_4005);
xnor U9273 (N_9273,N_1316,N_3390);
xnor U9274 (N_9274,N_353,N_3734);
nor U9275 (N_9275,N_793,N_2910);
nand U9276 (N_9276,N_3174,N_3164);
nand U9277 (N_9277,N_4945,N_1981);
xnor U9278 (N_9278,N_2654,N_4331);
or U9279 (N_9279,N_109,N_1700);
or U9280 (N_9280,N_4257,N_403);
and U9281 (N_9281,N_4090,N_2288);
xor U9282 (N_9282,N_3982,N_3152);
nand U9283 (N_9283,N_3493,N_3691);
or U9284 (N_9284,N_4260,N_3571);
or U9285 (N_9285,N_3312,N_2568);
nand U9286 (N_9286,N_2660,N_4265);
nand U9287 (N_9287,N_24,N_3927);
nor U9288 (N_9288,N_4423,N_4705);
nor U9289 (N_9289,N_1665,N_2493);
and U9290 (N_9290,N_3122,N_3625);
nand U9291 (N_9291,N_2174,N_761);
and U9292 (N_9292,N_814,N_1908);
nor U9293 (N_9293,N_4281,N_2152);
and U9294 (N_9294,N_1656,N_3438);
xor U9295 (N_9295,N_3204,N_630);
or U9296 (N_9296,N_4954,N_2784);
xor U9297 (N_9297,N_1591,N_2678);
nand U9298 (N_9298,N_2984,N_1200);
and U9299 (N_9299,N_1720,N_3666);
xor U9300 (N_9300,N_1578,N_2886);
or U9301 (N_9301,N_1003,N_1770);
and U9302 (N_9302,N_797,N_3354);
xor U9303 (N_9303,N_3292,N_915);
nand U9304 (N_9304,N_1842,N_3681);
nor U9305 (N_9305,N_1775,N_4732);
nor U9306 (N_9306,N_4670,N_2655);
and U9307 (N_9307,N_4419,N_2011);
or U9308 (N_9308,N_253,N_81);
nor U9309 (N_9309,N_2281,N_392);
or U9310 (N_9310,N_1004,N_2350);
or U9311 (N_9311,N_3106,N_2627);
or U9312 (N_9312,N_1007,N_4080);
xor U9313 (N_9313,N_2740,N_4426);
xnor U9314 (N_9314,N_1926,N_41);
or U9315 (N_9315,N_4769,N_3092);
xnor U9316 (N_9316,N_4264,N_2160);
nor U9317 (N_9317,N_3360,N_2774);
nor U9318 (N_9318,N_497,N_2822);
or U9319 (N_9319,N_4637,N_1886);
nand U9320 (N_9320,N_108,N_4797);
xnor U9321 (N_9321,N_2353,N_3676);
xor U9322 (N_9322,N_883,N_3650);
nor U9323 (N_9323,N_2411,N_3230);
and U9324 (N_9324,N_2743,N_4241);
xor U9325 (N_9325,N_330,N_806);
xor U9326 (N_9326,N_3186,N_1168);
nor U9327 (N_9327,N_3664,N_3563);
and U9328 (N_9328,N_3985,N_1288);
xnor U9329 (N_9329,N_202,N_1240);
nor U9330 (N_9330,N_4684,N_2727);
nand U9331 (N_9331,N_677,N_3244);
and U9332 (N_9332,N_2348,N_3612);
nor U9333 (N_9333,N_4417,N_2546);
nor U9334 (N_9334,N_2308,N_3417);
xnor U9335 (N_9335,N_1758,N_543);
nor U9336 (N_9336,N_4810,N_3622);
or U9337 (N_9337,N_3095,N_4025);
or U9338 (N_9338,N_4806,N_2764);
xor U9339 (N_9339,N_1239,N_1423);
nand U9340 (N_9340,N_4205,N_4767);
nor U9341 (N_9341,N_4167,N_3203);
xor U9342 (N_9342,N_1016,N_4621);
xor U9343 (N_9343,N_4668,N_3760);
nand U9344 (N_9344,N_804,N_3872);
or U9345 (N_9345,N_614,N_1510);
xnor U9346 (N_9346,N_1922,N_3684);
nand U9347 (N_9347,N_1281,N_4925);
nand U9348 (N_9348,N_3554,N_1398);
xor U9349 (N_9349,N_236,N_1091);
xnor U9350 (N_9350,N_1718,N_2080);
and U9351 (N_9351,N_2208,N_4720);
nor U9352 (N_9352,N_4058,N_4364);
xnor U9353 (N_9353,N_3850,N_4611);
xnor U9354 (N_9354,N_1984,N_2198);
and U9355 (N_9355,N_2082,N_1896);
nor U9356 (N_9356,N_2928,N_2110);
nand U9357 (N_9357,N_1717,N_15);
nand U9358 (N_9358,N_4541,N_4228);
nand U9359 (N_9359,N_2964,N_2614);
nand U9360 (N_9360,N_247,N_4418);
nor U9361 (N_9361,N_2587,N_1270);
nor U9362 (N_9362,N_4140,N_3427);
and U9363 (N_9363,N_75,N_452);
nor U9364 (N_9364,N_2426,N_1887);
xnor U9365 (N_9365,N_1915,N_4236);
nor U9366 (N_9366,N_706,N_835);
or U9367 (N_9367,N_1976,N_287);
xor U9368 (N_9368,N_3226,N_1741);
xor U9369 (N_9369,N_2948,N_566);
xor U9370 (N_9370,N_804,N_762);
xor U9371 (N_9371,N_1639,N_3160);
xnor U9372 (N_9372,N_4693,N_119);
nor U9373 (N_9373,N_701,N_2146);
or U9374 (N_9374,N_4665,N_3096);
or U9375 (N_9375,N_2925,N_4787);
and U9376 (N_9376,N_227,N_2716);
xor U9377 (N_9377,N_663,N_1599);
nor U9378 (N_9378,N_3781,N_3638);
nand U9379 (N_9379,N_1743,N_4578);
xnor U9380 (N_9380,N_1040,N_2611);
and U9381 (N_9381,N_4489,N_2289);
xor U9382 (N_9382,N_1645,N_1039);
nand U9383 (N_9383,N_4638,N_4142);
nor U9384 (N_9384,N_1174,N_253);
nor U9385 (N_9385,N_1370,N_3446);
and U9386 (N_9386,N_1131,N_2569);
nand U9387 (N_9387,N_3056,N_3409);
xnor U9388 (N_9388,N_20,N_109);
nand U9389 (N_9389,N_3487,N_1504);
nor U9390 (N_9390,N_3093,N_4683);
nand U9391 (N_9391,N_4355,N_4558);
nand U9392 (N_9392,N_1760,N_968);
nand U9393 (N_9393,N_4976,N_3745);
xor U9394 (N_9394,N_1565,N_731);
nand U9395 (N_9395,N_3883,N_75);
or U9396 (N_9396,N_4071,N_0);
nand U9397 (N_9397,N_2304,N_1638);
xor U9398 (N_9398,N_1095,N_1232);
nand U9399 (N_9399,N_4255,N_39);
nand U9400 (N_9400,N_1902,N_1458);
nor U9401 (N_9401,N_3596,N_2559);
xnor U9402 (N_9402,N_4461,N_810);
xor U9403 (N_9403,N_3662,N_3278);
and U9404 (N_9404,N_3397,N_2180);
nand U9405 (N_9405,N_2711,N_1536);
nor U9406 (N_9406,N_94,N_2472);
and U9407 (N_9407,N_2250,N_2630);
nand U9408 (N_9408,N_4302,N_2853);
xnor U9409 (N_9409,N_4982,N_2654);
or U9410 (N_9410,N_1741,N_1275);
nand U9411 (N_9411,N_4268,N_520);
nor U9412 (N_9412,N_4833,N_2428);
nor U9413 (N_9413,N_2104,N_873);
nor U9414 (N_9414,N_3736,N_3213);
xnor U9415 (N_9415,N_102,N_4378);
or U9416 (N_9416,N_2650,N_8);
nor U9417 (N_9417,N_839,N_525);
and U9418 (N_9418,N_2818,N_2501);
xor U9419 (N_9419,N_3519,N_563);
nor U9420 (N_9420,N_3425,N_4574);
and U9421 (N_9421,N_2123,N_3830);
or U9422 (N_9422,N_1100,N_4805);
and U9423 (N_9423,N_1085,N_3926);
xor U9424 (N_9424,N_4994,N_3599);
nand U9425 (N_9425,N_1302,N_2879);
and U9426 (N_9426,N_1048,N_2500);
xnor U9427 (N_9427,N_3360,N_4253);
or U9428 (N_9428,N_1609,N_2783);
nor U9429 (N_9429,N_2750,N_3763);
and U9430 (N_9430,N_901,N_4581);
or U9431 (N_9431,N_1488,N_1251);
nor U9432 (N_9432,N_3577,N_2328);
and U9433 (N_9433,N_1087,N_3986);
nand U9434 (N_9434,N_81,N_4880);
nand U9435 (N_9435,N_4716,N_2366);
nor U9436 (N_9436,N_2201,N_693);
nor U9437 (N_9437,N_363,N_359);
nor U9438 (N_9438,N_4974,N_3137);
xor U9439 (N_9439,N_1217,N_1267);
xor U9440 (N_9440,N_1718,N_4708);
xnor U9441 (N_9441,N_4022,N_2903);
nand U9442 (N_9442,N_815,N_2660);
or U9443 (N_9443,N_4872,N_4699);
or U9444 (N_9444,N_3400,N_276);
nand U9445 (N_9445,N_2228,N_1667);
and U9446 (N_9446,N_1679,N_1914);
nor U9447 (N_9447,N_4438,N_4241);
nand U9448 (N_9448,N_2465,N_4287);
xnor U9449 (N_9449,N_3406,N_4429);
or U9450 (N_9450,N_3747,N_3496);
and U9451 (N_9451,N_1216,N_2444);
xnor U9452 (N_9452,N_2311,N_2245);
nor U9453 (N_9453,N_2641,N_4900);
or U9454 (N_9454,N_3708,N_4398);
nor U9455 (N_9455,N_4922,N_3576);
or U9456 (N_9456,N_1871,N_2088);
nor U9457 (N_9457,N_1835,N_351);
nand U9458 (N_9458,N_113,N_3266);
xnor U9459 (N_9459,N_2521,N_3667);
or U9460 (N_9460,N_900,N_1277);
nand U9461 (N_9461,N_4836,N_1362);
xnor U9462 (N_9462,N_4491,N_1496);
xor U9463 (N_9463,N_2152,N_3126);
xor U9464 (N_9464,N_4663,N_2625);
nor U9465 (N_9465,N_2391,N_4271);
and U9466 (N_9466,N_1929,N_873);
nor U9467 (N_9467,N_3063,N_2691);
xor U9468 (N_9468,N_1781,N_455);
nand U9469 (N_9469,N_800,N_4188);
nand U9470 (N_9470,N_3075,N_4035);
nand U9471 (N_9471,N_195,N_1860);
xnor U9472 (N_9472,N_4190,N_3058);
nand U9473 (N_9473,N_4821,N_2331);
and U9474 (N_9474,N_499,N_237);
nor U9475 (N_9475,N_2595,N_1661);
xnor U9476 (N_9476,N_4930,N_3008);
and U9477 (N_9477,N_4331,N_4097);
nor U9478 (N_9478,N_3844,N_4676);
nand U9479 (N_9479,N_2961,N_4507);
and U9480 (N_9480,N_3332,N_40);
or U9481 (N_9481,N_589,N_4278);
nor U9482 (N_9482,N_1667,N_2001);
xnor U9483 (N_9483,N_850,N_3519);
nor U9484 (N_9484,N_1332,N_4145);
nor U9485 (N_9485,N_2096,N_2542);
nor U9486 (N_9486,N_3390,N_297);
or U9487 (N_9487,N_3307,N_2911);
xnor U9488 (N_9488,N_3046,N_3768);
nor U9489 (N_9489,N_1112,N_3899);
nand U9490 (N_9490,N_1065,N_1428);
and U9491 (N_9491,N_538,N_2181);
or U9492 (N_9492,N_2078,N_3618);
nand U9493 (N_9493,N_1667,N_1121);
nor U9494 (N_9494,N_3752,N_919);
or U9495 (N_9495,N_2309,N_4083);
nand U9496 (N_9496,N_1401,N_4085);
and U9497 (N_9497,N_1163,N_4980);
nand U9498 (N_9498,N_4524,N_2334);
or U9499 (N_9499,N_4628,N_2170);
xnor U9500 (N_9500,N_2266,N_3360);
or U9501 (N_9501,N_3411,N_4410);
or U9502 (N_9502,N_4689,N_3458);
xnor U9503 (N_9503,N_1944,N_265);
or U9504 (N_9504,N_2373,N_2401);
nand U9505 (N_9505,N_338,N_2584);
xor U9506 (N_9506,N_586,N_949);
xor U9507 (N_9507,N_3274,N_2278);
or U9508 (N_9508,N_4039,N_4988);
nand U9509 (N_9509,N_2721,N_4473);
or U9510 (N_9510,N_4239,N_494);
xnor U9511 (N_9511,N_369,N_2973);
and U9512 (N_9512,N_1414,N_2954);
xor U9513 (N_9513,N_3852,N_4788);
and U9514 (N_9514,N_2392,N_1706);
xor U9515 (N_9515,N_3615,N_2866);
nand U9516 (N_9516,N_591,N_399);
nor U9517 (N_9517,N_3047,N_2071);
nand U9518 (N_9518,N_3304,N_1764);
or U9519 (N_9519,N_355,N_1950);
and U9520 (N_9520,N_3390,N_4553);
or U9521 (N_9521,N_4271,N_2890);
and U9522 (N_9522,N_441,N_1603);
nand U9523 (N_9523,N_2653,N_529);
nand U9524 (N_9524,N_2028,N_408);
nor U9525 (N_9525,N_2502,N_594);
xor U9526 (N_9526,N_4376,N_426);
xor U9527 (N_9527,N_4837,N_380);
nor U9528 (N_9528,N_2095,N_364);
or U9529 (N_9529,N_1811,N_2370);
and U9530 (N_9530,N_4488,N_2203);
and U9531 (N_9531,N_2684,N_1035);
nand U9532 (N_9532,N_2802,N_1381);
xnor U9533 (N_9533,N_2052,N_1267);
nor U9534 (N_9534,N_1193,N_166);
or U9535 (N_9535,N_426,N_4946);
or U9536 (N_9536,N_4783,N_4999);
xor U9537 (N_9537,N_4138,N_3772);
or U9538 (N_9538,N_1626,N_4968);
xnor U9539 (N_9539,N_2210,N_1555);
and U9540 (N_9540,N_3698,N_2320);
nand U9541 (N_9541,N_3726,N_1181);
nor U9542 (N_9542,N_3547,N_4047);
and U9543 (N_9543,N_3935,N_4482);
nand U9544 (N_9544,N_3028,N_559);
xnor U9545 (N_9545,N_3261,N_4702);
and U9546 (N_9546,N_172,N_3258);
nand U9547 (N_9547,N_1206,N_2055);
and U9548 (N_9548,N_4429,N_2769);
xnor U9549 (N_9549,N_234,N_2803);
or U9550 (N_9550,N_3261,N_2291);
nand U9551 (N_9551,N_1078,N_465);
nand U9552 (N_9552,N_1696,N_1512);
nand U9553 (N_9553,N_2089,N_2990);
nor U9554 (N_9554,N_2330,N_274);
nand U9555 (N_9555,N_2636,N_3274);
nand U9556 (N_9556,N_1699,N_837);
nor U9557 (N_9557,N_2110,N_4205);
xor U9558 (N_9558,N_1946,N_3549);
or U9559 (N_9559,N_3717,N_1513);
xnor U9560 (N_9560,N_2163,N_1753);
and U9561 (N_9561,N_3596,N_3857);
nor U9562 (N_9562,N_3029,N_1064);
or U9563 (N_9563,N_3183,N_2141);
or U9564 (N_9564,N_620,N_616);
nor U9565 (N_9565,N_3179,N_4677);
nor U9566 (N_9566,N_268,N_4165);
and U9567 (N_9567,N_2236,N_3423);
nor U9568 (N_9568,N_4728,N_4488);
or U9569 (N_9569,N_256,N_510);
nor U9570 (N_9570,N_4930,N_205);
and U9571 (N_9571,N_1071,N_4775);
nor U9572 (N_9572,N_4148,N_2831);
xor U9573 (N_9573,N_935,N_841);
and U9574 (N_9574,N_1820,N_1558);
nand U9575 (N_9575,N_220,N_1790);
nor U9576 (N_9576,N_340,N_3865);
nor U9577 (N_9577,N_230,N_4933);
nor U9578 (N_9578,N_4786,N_2094);
and U9579 (N_9579,N_1586,N_2709);
nand U9580 (N_9580,N_2686,N_2784);
nor U9581 (N_9581,N_639,N_4770);
xnor U9582 (N_9582,N_4584,N_4681);
nor U9583 (N_9583,N_2561,N_3420);
nand U9584 (N_9584,N_4589,N_761);
and U9585 (N_9585,N_2677,N_4806);
xnor U9586 (N_9586,N_3982,N_2842);
nor U9587 (N_9587,N_4706,N_4578);
and U9588 (N_9588,N_4190,N_4873);
nand U9589 (N_9589,N_185,N_3191);
and U9590 (N_9590,N_419,N_3216);
and U9591 (N_9591,N_1179,N_2824);
and U9592 (N_9592,N_4416,N_629);
or U9593 (N_9593,N_1625,N_363);
nor U9594 (N_9594,N_2756,N_4791);
and U9595 (N_9595,N_3887,N_2683);
xnor U9596 (N_9596,N_2915,N_683);
xnor U9597 (N_9597,N_2355,N_3822);
xor U9598 (N_9598,N_4958,N_2673);
nand U9599 (N_9599,N_2283,N_4246);
nor U9600 (N_9600,N_2144,N_4325);
xor U9601 (N_9601,N_3434,N_2145);
xnor U9602 (N_9602,N_745,N_3514);
nand U9603 (N_9603,N_4624,N_2268);
or U9604 (N_9604,N_1077,N_277);
nand U9605 (N_9605,N_2371,N_3248);
nand U9606 (N_9606,N_4962,N_1705);
xnor U9607 (N_9607,N_1342,N_2839);
and U9608 (N_9608,N_3240,N_2151);
nor U9609 (N_9609,N_3484,N_1671);
and U9610 (N_9610,N_74,N_32);
nand U9611 (N_9611,N_4547,N_3870);
nand U9612 (N_9612,N_9,N_1684);
xnor U9613 (N_9613,N_809,N_1540);
xor U9614 (N_9614,N_713,N_650);
xor U9615 (N_9615,N_2620,N_4186);
or U9616 (N_9616,N_2068,N_956);
xor U9617 (N_9617,N_1426,N_800);
nor U9618 (N_9618,N_4643,N_3771);
nor U9619 (N_9619,N_3914,N_4251);
xor U9620 (N_9620,N_4469,N_1739);
nand U9621 (N_9621,N_1331,N_1831);
nor U9622 (N_9622,N_206,N_3029);
xnor U9623 (N_9623,N_1946,N_690);
nor U9624 (N_9624,N_4330,N_328);
or U9625 (N_9625,N_4473,N_1585);
nand U9626 (N_9626,N_3192,N_1549);
and U9627 (N_9627,N_539,N_545);
nor U9628 (N_9628,N_1368,N_4849);
xnor U9629 (N_9629,N_14,N_1403);
or U9630 (N_9630,N_4136,N_4681);
and U9631 (N_9631,N_4275,N_4337);
and U9632 (N_9632,N_2479,N_2926);
nand U9633 (N_9633,N_3646,N_4156);
or U9634 (N_9634,N_1214,N_3322);
xor U9635 (N_9635,N_1750,N_555);
and U9636 (N_9636,N_4023,N_3802);
xnor U9637 (N_9637,N_1829,N_3131);
nor U9638 (N_9638,N_544,N_2850);
xnor U9639 (N_9639,N_4317,N_4360);
or U9640 (N_9640,N_2017,N_2315);
or U9641 (N_9641,N_4507,N_1189);
or U9642 (N_9642,N_4341,N_2331);
and U9643 (N_9643,N_3287,N_72);
or U9644 (N_9644,N_3112,N_4011);
nor U9645 (N_9645,N_2188,N_71);
and U9646 (N_9646,N_335,N_2573);
and U9647 (N_9647,N_1215,N_1231);
or U9648 (N_9648,N_2555,N_3244);
nor U9649 (N_9649,N_4180,N_2630);
nand U9650 (N_9650,N_2566,N_769);
nand U9651 (N_9651,N_1648,N_2910);
or U9652 (N_9652,N_1590,N_4504);
nor U9653 (N_9653,N_4656,N_4989);
and U9654 (N_9654,N_3046,N_2780);
or U9655 (N_9655,N_76,N_1806);
or U9656 (N_9656,N_2267,N_1342);
nor U9657 (N_9657,N_224,N_3926);
nand U9658 (N_9658,N_2010,N_1804);
nor U9659 (N_9659,N_639,N_1533);
nand U9660 (N_9660,N_4156,N_549);
or U9661 (N_9661,N_1739,N_2856);
or U9662 (N_9662,N_3208,N_4201);
and U9663 (N_9663,N_3542,N_4061);
and U9664 (N_9664,N_32,N_1100);
and U9665 (N_9665,N_618,N_3866);
and U9666 (N_9666,N_1838,N_1862);
nor U9667 (N_9667,N_1853,N_1952);
xnor U9668 (N_9668,N_738,N_3054);
and U9669 (N_9669,N_4900,N_188);
and U9670 (N_9670,N_713,N_1107);
xnor U9671 (N_9671,N_3949,N_1720);
and U9672 (N_9672,N_1494,N_3847);
nor U9673 (N_9673,N_4815,N_3024);
and U9674 (N_9674,N_600,N_624);
nand U9675 (N_9675,N_1181,N_4707);
xor U9676 (N_9676,N_1945,N_3780);
xnor U9677 (N_9677,N_1188,N_3907);
nand U9678 (N_9678,N_4081,N_4838);
xor U9679 (N_9679,N_2832,N_2249);
xor U9680 (N_9680,N_3601,N_454);
xnor U9681 (N_9681,N_1683,N_2237);
or U9682 (N_9682,N_546,N_1586);
nor U9683 (N_9683,N_4406,N_2893);
and U9684 (N_9684,N_57,N_1448);
and U9685 (N_9685,N_3593,N_3316);
and U9686 (N_9686,N_52,N_938);
xnor U9687 (N_9687,N_662,N_3257);
nand U9688 (N_9688,N_476,N_2302);
and U9689 (N_9689,N_2284,N_4016);
and U9690 (N_9690,N_3335,N_872);
xor U9691 (N_9691,N_4637,N_512);
nand U9692 (N_9692,N_4820,N_4453);
nand U9693 (N_9693,N_4338,N_1286);
and U9694 (N_9694,N_401,N_1578);
xnor U9695 (N_9695,N_4535,N_2104);
nand U9696 (N_9696,N_4828,N_1312);
xnor U9697 (N_9697,N_1261,N_909);
nand U9698 (N_9698,N_1899,N_4821);
xnor U9699 (N_9699,N_1987,N_3796);
or U9700 (N_9700,N_3646,N_4686);
and U9701 (N_9701,N_2947,N_1693);
or U9702 (N_9702,N_2862,N_813);
and U9703 (N_9703,N_646,N_2586);
and U9704 (N_9704,N_1400,N_3472);
and U9705 (N_9705,N_3057,N_2777);
and U9706 (N_9706,N_3062,N_4713);
or U9707 (N_9707,N_2479,N_4992);
xor U9708 (N_9708,N_4498,N_1744);
xnor U9709 (N_9709,N_1600,N_4834);
xor U9710 (N_9710,N_3263,N_4085);
nand U9711 (N_9711,N_3429,N_180);
and U9712 (N_9712,N_4843,N_1179);
nor U9713 (N_9713,N_4060,N_2275);
nand U9714 (N_9714,N_2756,N_1721);
or U9715 (N_9715,N_1262,N_1059);
or U9716 (N_9716,N_2983,N_4107);
and U9717 (N_9717,N_163,N_167);
nor U9718 (N_9718,N_2714,N_4058);
nand U9719 (N_9719,N_2156,N_823);
xor U9720 (N_9720,N_4086,N_1328);
nor U9721 (N_9721,N_908,N_999);
nand U9722 (N_9722,N_4046,N_3381);
nand U9723 (N_9723,N_2525,N_3548);
nand U9724 (N_9724,N_4659,N_4430);
or U9725 (N_9725,N_2038,N_2848);
or U9726 (N_9726,N_3463,N_88);
and U9727 (N_9727,N_1080,N_4604);
and U9728 (N_9728,N_2635,N_709);
nor U9729 (N_9729,N_3650,N_3620);
xor U9730 (N_9730,N_4659,N_4840);
xor U9731 (N_9731,N_1032,N_1355);
nor U9732 (N_9732,N_195,N_2922);
or U9733 (N_9733,N_2264,N_3490);
or U9734 (N_9734,N_3974,N_166);
nor U9735 (N_9735,N_4772,N_2512);
xnor U9736 (N_9736,N_2612,N_4641);
and U9737 (N_9737,N_1024,N_249);
or U9738 (N_9738,N_2384,N_4636);
and U9739 (N_9739,N_3232,N_3532);
xnor U9740 (N_9740,N_956,N_2762);
nor U9741 (N_9741,N_1907,N_2459);
and U9742 (N_9742,N_58,N_2932);
or U9743 (N_9743,N_3199,N_4663);
and U9744 (N_9744,N_4641,N_1098);
xnor U9745 (N_9745,N_3389,N_1094);
and U9746 (N_9746,N_903,N_169);
nor U9747 (N_9747,N_1357,N_3076);
xor U9748 (N_9748,N_2869,N_1640);
nor U9749 (N_9749,N_2722,N_3066);
xor U9750 (N_9750,N_2222,N_489);
and U9751 (N_9751,N_2256,N_800);
nand U9752 (N_9752,N_1896,N_159);
or U9753 (N_9753,N_4662,N_3442);
or U9754 (N_9754,N_4444,N_3241);
nand U9755 (N_9755,N_9,N_4982);
nor U9756 (N_9756,N_2529,N_678);
nand U9757 (N_9757,N_1951,N_445);
xor U9758 (N_9758,N_1130,N_399);
xnor U9759 (N_9759,N_4903,N_988);
xnor U9760 (N_9760,N_3124,N_2638);
nor U9761 (N_9761,N_2012,N_4102);
nand U9762 (N_9762,N_473,N_2655);
or U9763 (N_9763,N_317,N_2171);
nor U9764 (N_9764,N_2009,N_4066);
xnor U9765 (N_9765,N_433,N_734);
nor U9766 (N_9766,N_837,N_1831);
or U9767 (N_9767,N_1,N_2396);
xor U9768 (N_9768,N_1335,N_1132);
nand U9769 (N_9769,N_3716,N_4898);
or U9770 (N_9770,N_27,N_3160);
nand U9771 (N_9771,N_3040,N_1209);
nand U9772 (N_9772,N_3298,N_4261);
nor U9773 (N_9773,N_2796,N_2961);
xor U9774 (N_9774,N_308,N_4064);
or U9775 (N_9775,N_4204,N_4213);
xor U9776 (N_9776,N_2863,N_3073);
or U9777 (N_9777,N_1965,N_2598);
or U9778 (N_9778,N_2851,N_3958);
nor U9779 (N_9779,N_976,N_1412);
nand U9780 (N_9780,N_52,N_4411);
xnor U9781 (N_9781,N_2262,N_1981);
nand U9782 (N_9782,N_3943,N_4292);
and U9783 (N_9783,N_685,N_1843);
nor U9784 (N_9784,N_975,N_3518);
or U9785 (N_9785,N_4441,N_2535);
or U9786 (N_9786,N_4836,N_1083);
xnor U9787 (N_9787,N_3029,N_932);
and U9788 (N_9788,N_2697,N_4181);
or U9789 (N_9789,N_3504,N_3023);
and U9790 (N_9790,N_3993,N_3527);
nand U9791 (N_9791,N_1910,N_4361);
nor U9792 (N_9792,N_2802,N_3339);
and U9793 (N_9793,N_2989,N_3579);
and U9794 (N_9794,N_4804,N_1503);
and U9795 (N_9795,N_4071,N_3187);
xor U9796 (N_9796,N_3253,N_1800);
nor U9797 (N_9797,N_2229,N_2839);
nor U9798 (N_9798,N_2309,N_2381);
nor U9799 (N_9799,N_3049,N_2985);
or U9800 (N_9800,N_389,N_130);
nand U9801 (N_9801,N_2287,N_2904);
nand U9802 (N_9802,N_3649,N_3348);
nor U9803 (N_9803,N_3128,N_372);
xnor U9804 (N_9804,N_1488,N_2005);
or U9805 (N_9805,N_818,N_2076);
nand U9806 (N_9806,N_2718,N_4675);
xor U9807 (N_9807,N_963,N_252);
nor U9808 (N_9808,N_4913,N_4201);
and U9809 (N_9809,N_4096,N_3529);
xor U9810 (N_9810,N_3267,N_49);
nor U9811 (N_9811,N_1942,N_1106);
and U9812 (N_9812,N_1919,N_3729);
xnor U9813 (N_9813,N_4267,N_4407);
or U9814 (N_9814,N_3029,N_4134);
nor U9815 (N_9815,N_1683,N_3131);
xnor U9816 (N_9816,N_2666,N_4272);
or U9817 (N_9817,N_4438,N_3416);
nor U9818 (N_9818,N_3229,N_4678);
or U9819 (N_9819,N_1268,N_324);
xnor U9820 (N_9820,N_3261,N_2095);
nand U9821 (N_9821,N_4472,N_3299);
or U9822 (N_9822,N_4189,N_1489);
nand U9823 (N_9823,N_3904,N_4236);
nand U9824 (N_9824,N_4814,N_178);
nand U9825 (N_9825,N_1841,N_4924);
xor U9826 (N_9826,N_1747,N_3994);
or U9827 (N_9827,N_3282,N_591);
or U9828 (N_9828,N_3198,N_2088);
xor U9829 (N_9829,N_1967,N_4175);
nand U9830 (N_9830,N_3428,N_1263);
and U9831 (N_9831,N_2182,N_3957);
and U9832 (N_9832,N_1242,N_4617);
nor U9833 (N_9833,N_3663,N_1007);
and U9834 (N_9834,N_4372,N_4431);
xor U9835 (N_9835,N_3172,N_763);
nand U9836 (N_9836,N_787,N_790);
or U9837 (N_9837,N_2425,N_81);
xnor U9838 (N_9838,N_3400,N_237);
nor U9839 (N_9839,N_3758,N_3460);
nand U9840 (N_9840,N_517,N_2704);
or U9841 (N_9841,N_4819,N_1482);
and U9842 (N_9842,N_4364,N_4117);
or U9843 (N_9843,N_3641,N_58);
nor U9844 (N_9844,N_3071,N_699);
nand U9845 (N_9845,N_2420,N_3418);
and U9846 (N_9846,N_2442,N_1094);
nor U9847 (N_9847,N_1771,N_104);
or U9848 (N_9848,N_4907,N_1165);
and U9849 (N_9849,N_1545,N_1483);
or U9850 (N_9850,N_3677,N_4292);
nand U9851 (N_9851,N_2302,N_4807);
nor U9852 (N_9852,N_766,N_2470);
or U9853 (N_9853,N_4082,N_3236);
or U9854 (N_9854,N_3782,N_662);
or U9855 (N_9855,N_3509,N_733);
or U9856 (N_9856,N_388,N_1814);
nor U9857 (N_9857,N_4257,N_2864);
nand U9858 (N_9858,N_4679,N_4822);
nand U9859 (N_9859,N_1288,N_1279);
nand U9860 (N_9860,N_2582,N_4794);
nor U9861 (N_9861,N_3943,N_2035);
nor U9862 (N_9862,N_4650,N_4543);
nand U9863 (N_9863,N_1328,N_3955);
and U9864 (N_9864,N_944,N_4693);
xnor U9865 (N_9865,N_3934,N_4353);
nand U9866 (N_9866,N_36,N_1340);
xnor U9867 (N_9867,N_855,N_708);
xor U9868 (N_9868,N_1059,N_3833);
nor U9869 (N_9869,N_2529,N_3947);
nand U9870 (N_9870,N_730,N_4250);
and U9871 (N_9871,N_572,N_4136);
xor U9872 (N_9872,N_3930,N_4415);
or U9873 (N_9873,N_2959,N_4639);
and U9874 (N_9874,N_2106,N_2674);
or U9875 (N_9875,N_4725,N_254);
xor U9876 (N_9876,N_2780,N_1057);
xor U9877 (N_9877,N_4588,N_3232);
or U9878 (N_9878,N_4478,N_4916);
xor U9879 (N_9879,N_556,N_2987);
and U9880 (N_9880,N_208,N_4690);
nor U9881 (N_9881,N_1946,N_4655);
and U9882 (N_9882,N_4709,N_2518);
nand U9883 (N_9883,N_2540,N_4647);
xor U9884 (N_9884,N_1791,N_269);
nand U9885 (N_9885,N_3321,N_872);
and U9886 (N_9886,N_2374,N_1283);
nand U9887 (N_9887,N_2772,N_2291);
nor U9888 (N_9888,N_2878,N_1603);
xor U9889 (N_9889,N_4455,N_3922);
nand U9890 (N_9890,N_252,N_1732);
nor U9891 (N_9891,N_777,N_3163);
nand U9892 (N_9892,N_1584,N_122);
and U9893 (N_9893,N_2853,N_4301);
nor U9894 (N_9894,N_464,N_2024);
and U9895 (N_9895,N_2282,N_2436);
nor U9896 (N_9896,N_1161,N_960);
nor U9897 (N_9897,N_2110,N_2806);
or U9898 (N_9898,N_363,N_4802);
and U9899 (N_9899,N_1887,N_525);
or U9900 (N_9900,N_3818,N_2796);
nand U9901 (N_9901,N_1036,N_1290);
nor U9902 (N_9902,N_3433,N_2756);
nand U9903 (N_9903,N_4338,N_3543);
or U9904 (N_9904,N_2666,N_717);
nand U9905 (N_9905,N_342,N_3811);
xor U9906 (N_9906,N_4018,N_39);
nor U9907 (N_9907,N_1723,N_1350);
nor U9908 (N_9908,N_2957,N_1999);
nor U9909 (N_9909,N_4134,N_3826);
nor U9910 (N_9910,N_2264,N_2922);
nor U9911 (N_9911,N_149,N_4589);
and U9912 (N_9912,N_3962,N_2510);
xnor U9913 (N_9913,N_535,N_3343);
and U9914 (N_9914,N_2111,N_1058);
and U9915 (N_9915,N_380,N_311);
and U9916 (N_9916,N_1388,N_1809);
or U9917 (N_9917,N_1572,N_4167);
xor U9918 (N_9918,N_895,N_4199);
or U9919 (N_9919,N_1482,N_1845);
xnor U9920 (N_9920,N_2918,N_1772);
nand U9921 (N_9921,N_322,N_3185);
nand U9922 (N_9922,N_3774,N_2388);
and U9923 (N_9923,N_4222,N_3502);
or U9924 (N_9924,N_8,N_2045);
or U9925 (N_9925,N_3959,N_2216);
or U9926 (N_9926,N_803,N_3523);
or U9927 (N_9927,N_1094,N_2375);
or U9928 (N_9928,N_4090,N_56);
xnor U9929 (N_9929,N_1099,N_1726);
or U9930 (N_9930,N_1799,N_71);
and U9931 (N_9931,N_1664,N_2390);
nand U9932 (N_9932,N_3883,N_568);
nor U9933 (N_9933,N_1696,N_2387);
xnor U9934 (N_9934,N_2029,N_3416);
nand U9935 (N_9935,N_2134,N_4034);
and U9936 (N_9936,N_2461,N_646);
nor U9937 (N_9937,N_291,N_1958);
xnor U9938 (N_9938,N_1150,N_210);
xor U9939 (N_9939,N_2551,N_1661);
xor U9940 (N_9940,N_4721,N_3994);
nor U9941 (N_9941,N_3658,N_3421);
or U9942 (N_9942,N_3991,N_2257);
and U9943 (N_9943,N_3847,N_487);
or U9944 (N_9944,N_275,N_3276);
or U9945 (N_9945,N_4464,N_2724);
and U9946 (N_9946,N_4058,N_3335);
and U9947 (N_9947,N_3805,N_2581);
nor U9948 (N_9948,N_3668,N_1840);
xnor U9949 (N_9949,N_158,N_2137);
nand U9950 (N_9950,N_831,N_417);
nor U9951 (N_9951,N_4187,N_2851);
xnor U9952 (N_9952,N_4371,N_131);
and U9953 (N_9953,N_4571,N_4080);
xnor U9954 (N_9954,N_4826,N_3568);
and U9955 (N_9955,N_3861,N_4564);
nor U9956 (N_9956,N_1708,N_3628);
nand U9957 (N_9957,N_2983,N_739);
or U9958 (N_9958,N_3190,N_219);
nand U9959 (N_9959,N_4969,N_1297);
nor U9960 (N_9960,N_1714,N_1562);
or U9961 (N_9961,N_1686,N_2703);
xnor U9962 (N_9962,N_1958,N_344);
or U9963 (N_9963,N_981,N_2889);
or U9964 (N_9964,N_1464,N_780);
nor U9965 (N_9965,N_1413,N_1923);
nor U9966 (N_9966,N_3690,N_2845);
nor U9967 (N_9967,N_310,N_4387);
xnor U9968 (N_9968,N_2729,N_554);
nand U9969 (N_9969,N_3196,N_1463);
nand U9970 (N_9970,N_1605,N_4181);
xor U9971 (N_9971,N_2522,N_2137);
and U9972 (N_9972,N_728,N_1667);
nor U9973 (N_9973,N_100,N_3199);
xnor U9974 (N_9974,N_462,N_4795);
or U9975 (N_9975,N_66,N_1511);
xnor U9976 (N_9976,N_4697,N_3615);
or U9977 (N_9977,N_2698,N_3888);
nand U9978 (N_9978,N_4360,N_2133);
xor U9979 (N_9979,N_1058,N_1513);
and U9980 (N_9980,N_369,N_160);
nor U9981 (N_9981,N_1936,N_3085);
or U9982 (N_9982,N_3298,N_4523);
xor U9983 (N_9983,N_1699,N_2202);
and U9984 (N_9984,N_918,N_39);
and U9985 (N_9985,N_3845,N_2906);
or U9986 (N_9986,N_2287,N_1004);
xnor U9987 (N_9987,N_1756,N_2740);
and U9988 (N_9988,N_174,N_2013);
or U9989 (N_9989,N_3158,N_3028);
nand U9990 (N_9990,N_2835,N_4379);
xor U9991 (N_9991,N_4452,N_1286);
nor U9992 (N_9992,N_1013,N_3179);
nor U9993 (N_9993,N_1211,N_2907);
xnor U9994 (N_9994,N_3957,N_3952);
nand U9995 (N_9995,N_2085,N_1241);
xor U9996 (N_9996,N_2097,N_3707);
nor U9997 (N_9997,N_4116,N_2433);
nor U9998 (N_9998,N_2730,N_2259);
and U9999 (N_9999,N_1728,N_2619);
nand U10000 (N_10000,N_7099,N_7338);
or U10001 (N_10001,N_7213,N_5022);
nand U10002 (N_10002,N_9131,N_8894);
and U10003 (N_10003,N_5369,N_9043);
nor U10004 (N_10004,N_6774,N_8384);
nand U10005 (N_10005,N_8893,N_9986);
and U10006 (N_10006,N_9057,N_9313);
or U10007 (N_10007,N_7634,N_8828);
xnor U10008 (N_10008,N_5165,N_6694);
and U10009 (N_10009,N_7810,N_5595);
nand U10010 (N_10010,N_7719,N_6157);
xor U10011 (N_10011,N_6371,N_5336);
nor U10012 (N_10012,N_9568,N_9252);
and U10013 (N_10013,N_8511,N_9185);
and U10014 (N_10014,N_9961,N_6740);
or U10015 (N_10015,N_6907,N_8514);
nor U10016 (N_10016,N_8379,N_5224);
and U10017 (N_10017,N_9555,N_8190);
or U10018 (N_10018,N_7987,N_5434);
xnor U10019 (N_10019,N_5605,N_6129);
or U10020 (N_10020,N_5966,N_6957);
or U10021 (N_10021,N_6817,N_5351);
nand U10022 (N_10022,N_9166,N_8691);
nand U10023 (N_10023,N_9471,N_9953);
and U10024 (N_10024,N_7764,N_5887);
and U10025 (N_10025,N_5046,N_7212);
xnor U10026 (N_10026,N_7761,N_6646);
xor U10027 (N_10027,N_5185,N_7113);
xor U10028 (N_10028,N_5058,N_9734);
nor U10029 (N_10029,N_7836,N_6836);
nor U10030 (N_10030,N_8347,N_7564);
and U10031 (N_10031,N_9881,N_5973);
nor U10032 (N_10032,N_9498,N_5540);
nand U10033 (N_10033,N_5702,N_7499);
xnor U10034 (N_10034,N_6331,N_8901);
or U10035 (N_10035,N_8789,N_7921);
nand U10036 (N_10036,N_5982,N_8058);
and U10037 (N_10037,N_9743,N_8534);
nor U10038 (N_10038,N_9490,N_8790);
xnor U10039 (N_10039,N_6118,N_6744);
xor U10040 (N_10040,N_8985,N_9692);
xnor U10041 (N_10041,N_5546,N_8301);
xnor U10042 (N_10042,N_9807,N_7732);
or U10043 (N_10043,N_6108,N_5190);
or U10044 (N_10044,N_7097,N_6903);
and U10045 (N_10045,N_6031,N_9606);
nor U10046 (N_10046,N_9048,N_8442);
and U10047 (N_10047,N_8427,N_7453);
and U10048 (N_10048,N_7833,N_7854);
or U10049 (N_10049,N_9010,N_9376);
and U10050 (N_10050,N_6120,N_7523);
and U10051 (N_10051,N_8770,N_6585);
xor U10052 (N_10052,N_5263,N_7762);
or U10053 (N_10053,N_8975,N_5220);
or U10054 (N_10054,N_9759,N_7901);
and U10055 (N_10055,N_6521,N_5312);
or U10056 (N_10056,N_5355,N_5164);
nor U10057 (N_10057,N_5929,N_6075);
or U10058 (N_10058,N_8703,N_8783);
xor U10059 (N_10059,N_8211,N_5675);
xnor U10060 (N_10060,N_7163,N_7891);
nand U10061 (N_10061,N_8880,N_9538);
and U10062 (N_10062,N_6698,N_6516);
or U10063 (N_10063,N_8295,N_6720);
nand U10064 (N_10064,N_7411,N_6218);
or U10065 (N_10065,N_7277,N_9429);
and U10066 (N_10066,N_7627,N_5236);
and U10067 (N_10067,N_5709,N_7646);
nand U10068 (N_10068,N_5961,N_9639);
nand U10069 (N_10069,N_6579,N_6524);
xor U10070 (N_10070,N_6601,N_7573);
or U10071 (N_10071,N_8484,N_6767);
nand U10072 (N_10072,N_8808,N_8272);
nor U10073 (N_10073,N_7154,N_8537);
and U10074 (N_10074,N_7856,N_7100);
and U10075 (N_10075,N_9314,N_8191);
or U10076 (N_10076,N_9911,N_5097);
nor U10077 (N_10077,N_5377,N_8735);
xnor U10078 (N_10078,N_7580,N_7758);
nand U10079 (N_10079,N_7557,N_9387);
xnor U10080 (N_10080,N_5813,N_8164);
xnor U10081 (N_10081,N_9181,N_8357);
or U10082 (N_10082,N_7045,N_6448);
xnor U10083 (N_10083,N_5326,N_9199);
and U10084 (N_10084,N_6576,N_5379);
nand U10085 (N_10085,N_7023,N_7363);
xnor U10086 (N_10086,N_9742,N_6475);
and U10087 (N_10087,N_9629,N_7668);
nor U10088 (N_10088,N_5138,N_7805);
xnor U10089 (N_10089,N_9381,N_9090);
and U10090 (N_10090,N_7400,N_5948);
and U10091 (N_10091,N_6865,N_8026);
nor U10092 (N_10092,N_7979,N_7597);
nand U10093 (N_10093,N_7519,N_6064);
or U10094 (N_10094,N_5755,N_6630);
xnor U10095 (N_10095,N_7455,N_8268);
and U10096 (N_10096,N_6933,N_8928);
and U10097 (N_10097,N_5510,N_9589);
nor U10098 (N_10098,N_9765,N_8418);
and U10099 (N_10099,N_5261,N_5426);
xor U10100 (N_10100,N_7983,N_9627);
or U10101 (N_10101,N_7418,N_8128);
nor U10102 (N_10102,N_7806,N_9413);
nand U10103 (N_10103,N_5584,N_6117);
xor U10104 (N_10104,N_7847,N_5036);
xnor U10105 (N_10105,N_7948,N_5012);
nor U10106 (N_10106,N_7509,N_5057);
xnor U10107 (N_10107,N_5989,N_7579);
xnor U10108 (N_10108,N_9192,N_7943);
nand U10109 (N_10109,N_8512,N_9642);
nand U10110 (N_10110,N_6388,N_9912);
and U10111 (N_10111,N_7117,N_6258);
xor U10112 (N_10112,N_9885,N_5944);
or U10113 (N_10113,N_8391,N_6586);
nand U10114 (N_10114,N_8800,N_6358);
nand U10115 (N_10115,N_5829,N_8791);
and U10116 (N_10116,N_7750,N_8728);
nor U10117 (N_10117,N_6423,N_7393);
nand U10118 (N_10118,N_7966,N_7310);
nand U10119 (N_10119,N_7636,N_6239);
or U10120 (N_10120,N_8948,N_9258);
nor U10121 (N_10121,N_5218,N_6590);
or U10122 (N_10122,N_6793,N_9619);
xor U10123 (N_10123,N_7725,N_6806);
xor U10124 (N_10124,N_9528,N_8621);
nand U10125 (N_10125,N_5625,N_7803);
and U10126 (N_10126,N_6783,N_7716);
xnor U10127 (N_10127,N_5958,N_7133);
nor U10128 (N_10128,N_7532,N_7216);
and U10129 (N_10129,N_8792,N_9355);
or U10130 (N_10130,N_9943,N_8570);
or U10131 (N_10131,N_6544,N_7791);
or U10132 (N_10132,N_6187,N_5331);
and U10133 (N_10133,N_6024,N_8297);
or U10134 (N_10134,N_8571,N_6899);
xor U10135 (N_10135,N_7221,N_9557);
or U10136 (N_10136,N_5309,N_5700);
and U10137 (N_10137,N_7250,N_9263);
or U10138 (N_10138,N_7409,N_9366);
nor U10139 (N_10139,N_6619,N_6476);
or U10140 (N_10140,N_5200,N_6846);
nor U10141 (N_10141,N_7735,N_5025);
and U10142 (N_10142,N_9651,N_6926);
xor U10143 (N_10143,N_5452,N_9180);
xor U10144 (N_10144,N_7884,N_7047);
xnor U10145 (N_10145,N_8669,N_8102);
xor U10146 (N_10146,N_6508,N_6425);
nor U10147 (N_10147,N_5541,N_9794);
nand U10148 (N_10148,N_7318,N_5542);
or U10149 (N_10149,N_6844,N_7570);
nand U10150 (N_10150,N_8978,N_6878);
xor U10151 (N_10151,N_5802,N_8101);
nor U10152 (N_10152,N_7687,N_7688);
xnor U10153 (N_10153,N_7392,N_9100);
xnor U10154 (N_10154,N_5677,N_9145);
xor U10155 (N_10155,N_8374,N_6324);
xor U10156 (N_10156,N_6299,N_7026);
or U10157 (N_10157,N_9107,N_7878);
nand U10158 (N_10158,N_9507,N_7641);
nand U10159 (N_10159,N_7441,N_6278);
xor U10160 (N_10160,N_5945,N_9595);
nand U10161 (N_10161,N_5979,N_9855);
xor U10162 (N_10162,N_6677,N_7741);
and U10163 (N_10163,N_7281,N_8806);
or U10164 (N_10164,N_5711,N_8244);
or U10165 (N_10165,N_6528,N_8865);
and U10166 (N_10166,N_7477,N_9927);
or U10167 (N_10167,N_9310,N_6773);
nand U10168 (N_10168,N_6682,N_9160);
or U10169 (N_10169,N_6302,N_7322);
nor U10170 (N_10170,N_7932,N_8736);
or U10171 (N_10171,N_9663,N_6447);
nand U10172 (N_10172,N_5791,N_6203);
xor U10173 (N_10173,N_7558,N_7146);
and U10174 (N_10174,N_5681,N_6693);
nor U10175 (N_10175,N_9929,N_6623);
xnor U10176 (N_10176,N_6000,N_7490);
xnor U10177 (N_10177,N_5300,N_9847);
and U10178 (N_10178,N_6385,N_5226);
or U10179 (N_10179,N_9036,N_9977);
nor U10180 (N_10180,N_6639,N_7300);
nor U10181 (N_10181,N_5091,N_6155);
nand U10182 (N_10182,N_8997,N_7141);
xor U10183 (N_10183,N_8335,N_5960);
and U10184 (N_10184,N_6548,N_9624);
and U10185 (N_10185,N_5494,N_7914);
or U10186 (N_10186,N_8771,N_9753);
or U10187 (N_10187,N_8499,N_5021);
or U10188 (N_10188,N_7357,N_5810);
nor U10189 (N_10189,N_9229,N_7612);
nand U10190 (N_10190,N_8710,N_8944);
or U10191 (N_10191,N_6925,N_8955);
or U10192 (N_10192,N_6483,N_8200);
nand U10193 (N_10193,N_9841,N_7463);
nand U10194 (N_10194,N_5382,N_6479);
xor U10195 (N_10195,N_8554,N_9712);
nor U10196 (N_10196,N_9359,N_9604);
nand U10197 (N_10197,N_6819,N_6849);
nor U10198 (N_10198,N_5969,N_9935);
and U10199 (N_10199,N_5832,N_8830);
and U10200 (N_10200,N_5668,N_7662);
xor U10201 (N_10201,N_7497,N_6684);
nor U10202 (N_10202,N_6478,N_7187);
and U10203 (N_10203,N_7984,N_5478);
and U10204 (N_10204,N_8594,N_8535);
nand U10205 (N_10205,N_9364,N_8553);
xor U10206 (N_10206,N_7958,N_8708);
xnor U10207 (N_10207,N_5198,N_5536);
xnor U10208 (N_10208,N_6100,N_5234);
xor U10209 (N_10209,N_5061,N_6622);
xor U10210 (N_10210,N_9669,N_8763);
nand U10211 (N_10211,N_5713,N_6496);
nor U10212 (N_10212,N_5282,N_8358);
nand U10213 (N_10213,N_8748,N_8834);
or U10214 (N_10214,N_6618,N_9632);
nand U10215 (N_10215,N_6431,N_6626);
nor U10216 (N_10216,N_5499,N_9078);
nand U10217 (N_10217,N_7412,N_6067);
and U10218 (N_10218,N_7759,N_7886);
and U10219 (N_10219,N_8049,N_9979);
nor U10220 (N_10220,N_7107,N_6053);
nand U10221 (N_10221,N_9170,N_8714);
and U10222 (N_10222,N_5622,N_5667);
nand U10223 (N_10223,N_9288,N_7071);
nor U10224 (N_10224,N_5910,N_8139);
xnor U10225 (N_10225,N_6073,N_9427);
nand U10226 (N_10226,N_6871,N_5741);
or U10227 (N_10227,N_7399,N_6914);
xnor U10228 (N_10228,N_5586,N_6341);
or U10229 (N_10229,N_8724,N_9227);
nand U10230 (N_10230,N_8014,N_9725);
nor U10231 (N_10231,N_6964,N_7653);
nand U10232 (N_10232,N_9957,N_6551);
or U10233 (N_10233,N_9491,N_9484);
xor U10234 (N_10234,N_5123,N_8394);
nand U10235 (N_10235,N_9660,N_9793);
and U10236 (N_10236,N_8019,N_9330);
xnor U10237 (N_10237,N_9201,N_7429);
or U10238 (N_10238,N_9674,N_7583);
nand U10239 (N_10239,N_5160,N_8930);
nor U10240 (N_10240,N_8879,N_7291);
and U10241 (N_10241,N_6344,N_7718);
or U10242 (N_10242,N_9095,N_5275);
or U10243 (N_10243,N_8671,N_9294);
nor U10244 (N_10244,N_5335,N_7252);
nand U10245 (N_10245,N_6082,N_9138);
nor U10246 (N_10246,N_6301,N_9579);
or U10247 (N_10247,N_8994,N_6246);
and U10248 (N_10248,N_8832,N_7031);
nor U10249 (N_10249,N_7695,N_5816);
xor U10250 (N_10250,N_6690,N_5323);
nor U10251 (N_10251,N_6180,N_6657);
nor U10252 (N_10252,N_5620,N_6389);
and U10253 (N_10253,N_7960,N_6975);
xnor U10254 (N_10254,N_6598,N_6578);
nor U10255 (N_10255,N_9705,N_8424);
xnor U10256 (N_10256,N_9840,N_7872);
nand U10257 (N_10257,N_7443,N_9634);
or U10258 (N_10258,N_6285,N_5628);
nor U10259 (N_10259,N_5408,N_7950);
or U10260 (N_10260,N_8551,N_8317);
nand U10261 (N_10261,N_7027,N_7843);
nand U10262 (N_10262,N_5767,N_9880);
nand U10263 (N_10263,N_9316,N_9800);
and U10264 (N_10264,N_5936,N_6864);
or U10265 (N_10265,N_5116,N_5462);
and U10266 (N_10266,N_5397,N_5512);
nand U10267 (N_10267,N_6281,N_5135);
and U10268 (N_10268,N_7711,N_6854);
xnor U10269 (N_10269,N_9854,N_6300);
xor U10270 (N_10270,N_8324,N_8812);
nor U10271 (N_10271,N_8827,N_6788);
xor U10272 (N_10272,N_6858,N_6036);
xor U10273 (N_10273,N_5154,N_9803);
or U10274 (N_10274,N_6127,N_9871);
or U10275 (N_10275,N_7421,N_8527);
xor U10276 (N_10276,N_8677,N_8895);
or U10277 (N_10277,N_6104,N_5330);
nand U10278 (N_10278,N_9221,N_9578);
nand U10279 (N_10279,N_8543,N_7427);
and U10280 (N_10280,N_9018,N_5492);
and U10281 (N_10281,N_7637,N_7489);
nand U10282 (N_10282,N_5465,N_6821);
and U10283 (N_10283,N_6007,N_7140);
nor U10284 (N_10284,N_9340,N_8114);
and U10285 (N_10285,N_9923,N_6125);
nand U10286 (N_10286,N_6613,N_8127);
nand U10287 (N_10287,N_9818,N_5819);
or U10288 (N_10288,N_8521,N_9388);
or U10289 (N_10289,N_9984,N_9142);
nand U10290 (N_10290,N_5780,N_8867);
xnor U10291 (N_10291,N_5597,N_9951);
or U10292 (N_10292,N_9037,N_6928);
xnor U10293 (N_10293,N_6947,N_6786);
nand U10294 (N_10294,N_7424,N_5642);
nand U10295 (N_10295,N_6028,N_7743);
or U10296 (N_10296,N_6137,N_7237);
nand U10297 (N_10297,N_6881,N_6374);
xor U10298 (N_10298,N_6497,N_6756);
nor U10299 (N_10299,N_9990,N_9396);
nor U10300 (N_10300,N_7957,N_9715);
and U10301 (N_10301,N_9703,N_9457);
nor U10302 (N_10302,N_8953,N_7470);
and U10303 (N_10303,N_9781,N_6839);
xor U10304 (N_10304,N_5208,N_6348);
or U10305 (N_10305,N_9958,N_8775);
nor U10306 (N_10306,N_8129,N_9339);
xor U10307 (N_10307,N_5483,N_7143);
xor U10308 (N_10308,N_7933,N_8130);
or U10309 (N_10309,N_9292,N_5578);
nor U10310 (N_10310,N_6828,N_5750);
and U10311 (N_10311,N_7828,N_9102);
xor U10312 (N_10312,N_9699,N_5604);
and U10313 (N_10313,N_8426,N_5360);
and U10314 (N_10314,N_7265,N_5946);
or U10315 (N_10315,N_5029,N_5735);
xnor U10316 (N_10316,N_8638,N_6018);
nand U10317 (N_10317,N_8480,N_7209);
and U10318 (N_10318,N_7576,N_7912);
xnor U10319 (N_10319,N_7638,N_7474);
nand U10320 (N_10320,N_9477,N_8900);
xor U10321 (N_10321,N_5556,N_7348);
nor U10322 (N_10322,N_9426,N_8608);
nor U10323 (N_10323,N_6996,N_7486);
and U10324 (N_10324,N_9442,N_8449);
nand U10325 (N_10325,N_5757,N_6621);
nor U10326 (N_10326,N_9972,N_7178);
nand U10327 (N_10327,N_8366,N_9909);
xnor U10328 (N_10328,N_5919,N_7610);
xnor U10329 (N_10329,N_7088,N_6002);
xor U10330 (N_10330,N_5993,N_7425);
or U10331 (N_10331,N_7385,N_7572);
xor U10332 (N_10332,N_9744,N_5939);
and U10333 (N_10333,N_8675,N_6445);
nand U10334 (N_10334,N_7793,N_9779);
xor U10335 (N_10335,N_9539,N_8633);
and U10336 (N_10336,N_8959,N_9474);
nand U10337 (N_10337,N_7368,N_7076);
or U10338 (N_10338,N_9347,N_8623);
or U10339 (N_10339,N_5392,N_7752);
or U10340 (N_10340,N_6591,N_6874);
and U10341 (N_10341,N_7458,N_6495);
xor U10342 (N_10342,N_6319,N_6805);
nand U10343 (N_10343,N_7606,N_7065);
or U10344 (N_10344,N_5161,N_7297);
or U10345 (N_10345,N_6294,N_8483);
and U10346 (N_10346,N_5056,N_9256);
nor U10347 (N_10347,N_7101,N_9400);
and U10348 (N_10348,N_9092,N_6199);
nand U10349 (N_10349,N_5108,N_8151);
nand U10350 (N_10350,N_9144,N_9875);
and U10351 (N_10351,N_5761,N_5143);
xor U10352 (N_10352,N_6843,N_7740);
or U10353 (N_10353,N_6503,N_5346);
nand U10354 (N_10354,N_7595,N_9924);
or U10355 (N_10355,N_6046,N_5828);
nor U10356 (N_10356,N_5406,N_9769);
or U10357 (N_10357,N_8022,N_8653);
xnor U10358 (N_10358,N_8686,N_6109);
xnor U10359 (N_10359,N_7650,N_8194);
or U10360 (N_10360,N_6257,N_9513);
or U10361 (N_10361,N_5039,N_9159);
nor U10362 (N_10362,N_8363,N_9419);
and U10363 (N_10363,N_5296,N_6310);
and U10364 (N_10364,N_6215,N_8839);
nor U10365 (N_10365,N_9571,N_7457);
xnor U10366 (N_10366,N_8174,N_6494);
and U10367 (N_10367,N_9675,N_7785);
xor U10368 (N_10368,N_8343,N_5402);
nand U10369 (N_10369,N_8096,N_7705);
or U10370 (N_10370,N_5603,N_7386);
nand U10371 (N_10371,N_8933,N_5322);
nor U10372 (N_10372,N_8060,N_5691);
or U10373 (N_10373,N_8001,N_6340);
nor U10374 (N_10374,N_8250,N_6200);
and U10375 (N_10375,N_9008,N_9780);
nand U10376 (N_10376,N_5202,N_7186);
or U10377 (N_10377,N_7751,N_6372);
nor U10378 (N_10378,N_6818,N_6008);
nand U10379 (N_10379,N_6972,N_8607);
and U10380 (N_10380,N_7858,N_9939);
and U10381 (N_10381,N_7316,N_6277);
nor U10382 (N_10382,N_7450,N_8273);
nand U10383 (N_10383,N_8729,N_5067);
xnor U10384 (N_10384,N_8977,N_7218);
or U10385 (N_10385,N_7816,N_9547);
nand U10386 (N_10386,N_7929,N_7563);
nand U10387 (N_10387,N_5196,N_7551);
xnor U10388 (N_10388,N_6406,N_8012);
nor U10389 (N_10389,N_7547,N_9284);
nor U10390 (N_10390,N_7295,N_7736);
and U10391 (N_10391,N_7371,N_5228);
xor U10392 (N_10392,N_5368,N_8110);
or U10393 (N_10393,N_8257,N_5089);
xor U10394 (N_10394,N_6399,N_7536);
and U10395 (N_10395,N_8654,N_7378);
nor U10396 (N_10396,N_7164,N_5192);
nor U10397 (N_10397,N_6955,N_8218);
and U10398 (N_10398,N_6671,N_6550);
nand U10399 (N_10399,N_7849,N_8848);
nand U10400 (N_10400,N_9895,N_8302);
nor U10401 (N_10401,N_6059,N_8940);
or U10402 (N_10402,N_6848,N_5136);
nor U10403 (N_10403,N_7661,N_7655);
nor U10404 (N_10404,N_8986,N_6553);
nand U10405 (N_10405,N_5823,N_5571);
nand U10406 (N_10406,N_9168,N_9823);
or U10407 (N_10407,N_5696,N_9422);
xor U10408 (N_10408,N_8443,N_7428);
xor U10409 (N_10409,N_8903,N_7203);
and U10410 (N_10410,N_7248,N_5239);
nand U10411 (N_10411,N_9319,N_9024);
and U10412 (N_10412,N_6438,N_6173);
nor U10413 (N_10413,N_6205,N_6672);
nand U10414 (N_10414,N_9563,N_8744);
nand U10415 (N_10415,N_6889,N_6823);
xor U10416 (N_10416,N_9545,N_6969);
or U10417 (N_10417,N_6570,N_9352);
and U10418 (N_10418,N_6739,N_7120);
and U10419 (N_10419,N_5343,N_6396);
nand U10420 (N_10420,N_7207,N_5815);
xor U10421 (N_10421,N_5518,N_9820);
and U10422 (N_10422,N_5291,N_9161);
xor U10423 (N_10423,N_9281,N_9852);
nor U10424 (N_10424,N_6620,N_7728);
nand U10425 (N_10425,N_5428,N_9942);
nor U10426 (N_10426,N_8841,N_6432);
and U10427 (N_10427,N_5646,N_7435);
nand U10428 (N_10428,N_7152,N_7276);
xnor U10429 (N_10429,N_9460,N_8531);
nand U10430 (N_10430,N_5693,N_5888);
nor U10431 (N_10431,N_5078,N_5252);
or U10432 (N_10432,N_6454,N_7122);
and U10433 (N_10433,N_5028,N_7440);
xor U10434 (N_10434,N_9424,N_9446);
and U10435 (N_10435,N_5787,N_8312);
or U10436 (N_10436,N_9534,N_5447);
nor U10437 (N_10437,N_9623,N_7928);
nand U10438 (N_10438,N_6317,N_5390);
nand U10439 (N_10439,N_7312,N_6184);
nor U10440 (N_10440,N_7342,N_6984);
nand U10441 (N_10441,N_9752,N_7776);
or U10442 (N_10442,N_7404,N_6559);
nor U10443 (N_10443,N_5384,N_5784);
nand U10444 (N_10444,N_7516,N_9197);
nor U10445 (N_10445,N_9384,N_6163);
or U10446 (N_10446,N_6139,N_6212);
and U10447 (N_10447,N_5125,N_8912);
xor U10448 (N_10448,N_8741,N_7666);
or U10449 (N_10449,N_7787,N_5177);
and U10450 (N_10450,N_9104,N_8068);
nor U10451 (N_10451,N_8353,N_7430);
nor U10452 (N_10452,N_6932,N_8138);
nor U10453 (N_10453,N_6997,N_9717);
and U10454 (N_10454,N_5126,N_7083);
xor U10455 (N_10455,N_8971,N_5055);
and U10456 (N_10456,N_9709,N_7370);
or U10457 (N_10457,N_7451,N_5371);
xor U10458 (N_10458,N_5880,N_8784);
nor U10459 (N_10459,N_5068,N_6297);
xor U10460 (N_10460,N_6336,N_8469);
xnor U10461 (N_10461,N_9030,N_7993);
xnor U10462 (N_10462,N_9874,N_5773);
or U10463 (N_10463,N_8630,N_8267);
and U10464 (N_10464,N_9701,N_5931);
nor U10465 (N_10465,N_6021,N_6295);
and U10466 (N_10466,N_9337,N_9262);
nor U10467 (N_10467,N_8329,N_5474);
and U10468 (N_10468,N_6992,N_6575);
and U10469 (N_10469,N_9960,N_9832);
nand U10470 (N_10470,N_8592,N_7041);
xor U10471 (N_10471,N_7330,N_6275);
xor U10472 (N_10472,N_5339,N_6781);
nor U10473 (N_10473,N_7234,N_7746);
nor U10474 (N_10474,N_6851,N_5023);
or U10475 (N_10475,N_5487,N_6020);
nand U10476 (N_10476,N_7364,N_6261);
nand U10477 (N_10477,N_8029,N_6769);
or U10478 (N_10478,N_8204,N_9069);
nor U10479 (N_10479,N_5159,N_8451);
xnor U10480 (N_10480,N_5533,N_8316);
xor U10481 (N_10481,N_5516,N_9916);
xnor U10482 (N_10482,N_9115,N_5444);
or U10483 (N_10483,N_5588,N_6242);
nor U10484 (N_10484,N_9375,N_8846);
or U10485 (N_10485,N_9487,N_6323);
or U10486 (N_10486,N_7714,N_5304);
nand U10487 (N_10487,N_6599,N_8210);
nor U10488 (N_10488,N_5890,N_5648);
nand U10489 (N_10489,N_8196,N_7320);
xnor U10490 (N_10490,N_8146,N_6255);
or U10491 (N_10491,N_9383,N_7329);
nand U10492 (N_10492,N_9906,N_7643);
or U10493 (N_10493,N_6262,N_8546);
nand U10494 (N_10494,N_7080,N_7414);
nand U10495 (N_10495,N_7383,N_7199);
xor U10496 (N_10496,N_6446,N_5180);
nor U10497 (N_10497,N_9249,N_8497);
nand U10498 (N_10498,N_9282,N_7842);
or U10499 (N_10499,N_8702,N_9931);
xor U10500 (N_10500,N_5685,N_5650);
nand U10501 (N_10501,N_6128,N_6052);
xnor U10502 (N_10502,N_6654,N_7147);
xor U10503 (N_10503,N_6350,N_9804);
or U10504 (N_10504,N_7883,N_8380);
xnor U10505 (N_10505,N_5488,N_5651);
nor U10506 (N_10506,N_7520,N_5844);
nand U10507 (N_10507,N_8387,N_7201);
and U10508 (N_10508,N_5457,N_6349);
nor U10509 (N_10509,N_8208,N_7394);
nand U10510 (N_10510,N_5598,N_7894);
or U10511 (N_10511,N_5289,N_6329);
xor U10512 (N_10512,N_7998,N_5801);
nand U10513 (N_10513,N_9338,N_7305);
nor U10514 (N_10514,N_9033,N_6343);
or U10515 (N_10515,N_8436,N_7992);
nand U10516 (N_10516,N_6896,N_7157);
nor U10517 (N_10517,N_7920,N_6791);
xor U10518 (N_10518,N_7206,N_7376);
and U10519 (N_10519,N_5800,N_7593);
xnor U10520 (N_10520,N_7881,N_6229);
or U10521 (N_10521,N_9679,N_8408);
xnor U10522 (N_10522,N_5834,N_5900);
xnor U10523 (N_10523,N_8486,N_6443);
xnor U10524 (N_10524,N_7888,N_5140);
xor U10525 (N_10525,N_7697,N_8159);
xor U10526 (N_10526,N_6605,N_7156);
and U10527 (N_10527,N_7895,N_8574);
nor U10528 (N_10528,N_7500,N_5174);
or U10529 (N_10529,N_5972,N_6920);
nor U10530 (N_10530,N_6051,N_6063);
and U10531 (N_10531,N_7682,N_6900);
xor U10532 (N_10532,N_5042,N_7644);
xnor U10533 (N_10533,N_7652,N_9582);
xor U10534 (N_10534,N_8361,N_8352);
xor U10535 (N_10535,N_9049,N_8938);
xnor U10536 (N_10536,N_6243,N_5701);
or U10537 (N_10537,N_5520,N_5376);
and U10538 (N_10538,N_7259,N_9905);
and U10539 (N_10539,N_7515,N_7261);
nand U10540 (N_10540,N_7321,N_9122);
or U10541 (N_10541,N_5420,N_8406);
and U10542 (N_10542,N_6142,N_7674);
xnor U10543 (N_10543,N_6703,N_8287);
or U10544 (N_10544,N_9700,N_5258);
and U10545 (N_10545,N_9593,N_8787);
nand U10546 (N_10546,N_5082,N_9401);
xnor U10547 (N_10547,N_9889,N_6967);
xnor U10548 (N_10548,N_9328,N_9118);
nor U10549 (N_10549,N_9599,N_6629);
and U10550 (N_10550,N_6826,N_8993);
or U10551 (N_10551,N_5708,N_8091);
nor U10552 (N_10552,N_9265,N_6678);
nand U10553 (N_10553,N_8690,N_9940);
nand U10554 (N_10554,N_9902,N_6596);
nor U10555 (N_10555,N_5134,N_8399);
nor U10556 (N_10556,N_8382,N_6434);
xor U10557 (N_10557,N_9654,N_5484);
nor U10558 (N_10558,N_7108,N_6870);
and U10559 (N_10559,N_6332,N_5652);
nor U10560 (N_10560,N_6581,N_5153);
nand U10561 (N_10561,N_8254,N_6572);
xnor U10562 (N_10562,N_7043,N_7049);
nand U10563 (N_10563,N_8502,N_9272);
xnor U10564 (N_10564,N_8713,N_6689);
and U10565 (N_10565,N_7915,N_5502);
xor U10566 (N_10566,N_8261,N_8305);
and U10567 (N_10567,N_6604,N_6418);
nand U10568 (N_10568,N_5493,N_6283);
nor U10569 (N_10569,N_7623,N_6238);
xnor U10570 (N_10570,N_5285,N_8863);
or U10571 (N_10571,N_7035,N_8627);
nand U10572 (N_10572,N_5468,N_7040);
nor U10573 (N_10573,N_8400,N_7491);
nand U10574 (N_10574,N_5596,N_7562);
xor U10575 (N_10575,N_7339,N_6845);
and U10576 (N_10576,N_7072,N_5785);
or U10577 (N_10577,N_8233,N_6792);
nand U10578 (N_10578,N_7734,N_9811);
nor U10579 (N_10579,N_6561,N_6269);
xnor U10580 (N_10580,N_6259,N_9345);
nand U10581 (N_10581,N_8336,N_6722);
nand U10582 (N_10582,N_9919,N_7530);
or U10583 (N_10583,N_9097,N_7158);
nand U10584 (N_10584,N_9859,N_5987);
xor U10585 (N_10585,N_8518,N_8025);
xnor U10586 (N_10586,N_5010,N_5230);
nor U10587 (N_10587,N_7304,N_7826);
nor U10588 (N_10588,N_6426,N_5666);
nand U10589 (N_10589,N_8581,N_5740);
nand U10590 (N_10590,N_7887,N_5414);
xnor U10591 (N_10591,N_9494,N_5537);
xnor U10592 (N_10592,N_5265,N_8507);
or U10593 (N_10593,N_6663,N_8754);
nor U10594 (N_10594,N_8921,N_9128);
and U10595 (N_10595,N_8354,N_7105);
nand U10596 (N_10596,N_6417,N_8999);
or U10597 (N_10597,N_6135,N_9127);
nand U10598 (N_10598,N_6251,N_9285);
nor U10599 (N_10599,N_8673,N_8919);
xor U10600 (N_10600,N_8651,N_9303);
nor U10601 (N_10601,N_9341,N_6867);
nand U10602 (N_10602,N_7538,N_6614);
and U10603 (N_10603,N_5366,N_6363);
nor U10604 (N_10604,N_6264,N_7372);
nand U10605 (N_10605,N_6178,N_5908);
nand U10606 (N_10606,N_9827,N_9501);
or U10607 (N_10607,N_9938,N_7931);
nor U10608 (N_10608,N_6961,N_6760);
or U10609 (N_10609,N_7846,N_9226);
xnor U10610 (N_10610,N_9948,N_9783);
nand U10611 (N_10611,N_5047,N_5992);
xnor U10612 (N_10612,N_9837,N_5325);
xor U10613 (N_10613,N_5051,N_7387);
or U10614 (N_10614,N_8455,N_9395);
xor U10615 (N_10615,N_6347,N_8116);
or U10616 (N_10616,N_9708,N_8960);
nand U10617 (N_10617,N_5521,N_8003);
and U10618 (N_10618,N_6342,N_7771);
and U10619 (N_10619,N_9215,N_5026);
nand U10620 (N_10620,N_6412,N_8052);
nor U10621 (N_10621,N_5233,N_9857);
or U10622 (N_10622,N_9011,N_8038);
nand U10623 (N_10623,N_8871,N_6138);
or U10624 (N_10624,N_6315,N_6022);
and U10625 (N_10625,N_9596,N_6768);
and U10626 (N_10626,N_7438,N_7664);
nand U10627 (N_10627,N_7433,N_8359);
xor U10628 (N_10628,N_7543,N_6824);
xnor U10629 (N_10629,N_8145,N_9760);
nand U10630 (N_10630,N_6025,N_5508);
and U10631 (N_10631,N_8652,N_8011);
and U10632 (N_10632,N_7258,N_9397);
and U10633 (N_10633,N_6633,N_7266);
and U10634 (N_10634,N_9451,N_5805);
xor U10635 (N_10635,N_8346,N_8550);
nor U10636 (N_10636,N_7225,N_8524);
xnor U10637 (N_10637,N_6183,N_8464);
nand U10638 (N_10638,N_9843,N_6640);
or U10639 (N_10639,N_9059,N_6536);
nor U10640 (N_10640,N_6395,N_7654);
nor U10641 (N_10641,N_6987,N_9653);
xnor U10642 (N_10642,N_9936,N_9182);
xor U10643 (N_10643,N_7723,N_8006);
and U10644 (N_10644,N_7838,N_7864);
or U10645 (N_10645,N_6529,N_8614);
and U10646 (N_10646,N_7374,N_5762);
nor U10647 (N_10647,N_6898,N_9791);
nand U10648 (N_10648,N_9416,N_8926);
and U10649 (N_10649,N_6355,N_8536);
nor U10650 (N_10650,N_9649,N_6884);
nand U10651 (N_10651,N_8516,N_6723);
nand U10652 (N_10652,N_7899,N_8881);
nor U10653 (N_10653,N_9560,N_7116);
nor U10654 (N_10654,N_9019,N_7945);
and U10655 (N_10655,N_6832,N_8568);
or U10656 (N_10656,N_6436,N_8279);
xor U10657 (N_10657,N_9731,N_6866);
nand U10658 (N_10658,N_8197,N_8509);
nand U10659 (N_10659,N_6413,N_6291);
nor U10660 (N_10660,N_6979,N_6091);
nor U10661 (N_10661,N_6804,N_6699);
nor U10662 (N_10662,N_5002,N_5418);
nand U10663 (N_10663,N_9559,N_5223);
xor U10664 (N_10664,N_5614,N_5922);
xor U10665 (N_10665,N_5370,N_8080);
and U10666 (N_10666,N_5245,N_7037);
nand U10667 (N_10667,N_8106,N_8746);
and U10668 (N_10668,N_9354,N_5114);
or U10669 (N_10669,N_6507,N_9088);
nand U10670 (N_10670,N_7681,N_7229);
nand U10671 (N_10671,N_5974,N_8171);
nand U10672 (N_10672,N_8781,N_6398);
or U10673 (N_10673,N_6519,N_6597);
nand U10674 (N_10674,N_8477,N_7459);
or U10675 (N_10675,N_7969,N_9235);
or U10676 (N_10676,N_8582,N_8296);
or U10677 (N_10677,N_7510,N_8017);
nor U10678 (N_10678,N_6842,N_6513);
nor U10679 (N_10679,N_5187,N_8162);
xnor U10680 (N_10680,N_5712,N_8332);
and U10681 (N_10681,N_8811,N_9436);
or U10682 (N_10682,N_9955,N_7568);
and U10683 (N_10683,N_8717,N_8872);
nand U10684 (N_10684,N_7622,N_8243);
or U10685 (N_10685,N_7264,N_5102);
nand U10686 (N_10686,N_9710,N_8041);
nand U10687 (N_10687,N_7939,N_7090);
xnor U10688 (N_10688,N_9207,N_6681);
xnor U10689 (N_10689,N_9497,N_6069);
nor U10690 (N_10690,N_7254,N_9299);
or U10691 (N_10691,N_9601,N_5415);
or U10692 (N_10692,N_6256,N_6411);
nor U10693 (N_10693,N_5117,N_7460);
nand U10694 (N_10694,N_6841,N_5416);
or U10695 (N_10695,N_7050,N_5354);
or U10696 (N_10696,N_7786,N_6304);
nor U10697 (N_10697,N_6154,N_5237);
and U10698 (N_10698,N_5806,N_9452);
or U10699 (N_10699,N_8056,N_9480);
nand U10700 (N_10700,N_9810,N_7645);
nor U10701 (N_10701,N_9719,N_9728);
nand U10702 (N_10702,N_8457,N_7524);
xor U10703 (N_10703,N_6812,N_6111);
nor U10704 (N_10704,N_9861,N_6404);
nand U10705 (N_10705,N_5727,N_8161);
nor U10706 (N_10706,N_7533,N_5615);
xor U10707 (N_10707,N_7823,N_8050);
nand U10708 (N_10708,N_5580,N_9266);
nor U10709 (N_10709,N_8961,N_8591);
or U10710 (N_10710,N_7260,N_8737);
xor U10711 (N_10711,N_8866,N_5710);
and U10712 (N_10712,N_6840,N_6352);
nand U10713 (N_10713,N_9581,N_9683);
xnor U10714 (N_10714,N_6778,N_7684);
and U10715 (N_10715,N_6938,N_8131);
nor U10716 (N_10716,N_9365,N_7468);
nor U10717 (N_10717,N_8722,N_7150);
or U10718 (N_10718,N_7292,N_5456);
xor U10719 (N_10719,N_8949,N_8241);
nand U10720 (N_10720,N_7985,N_9468);
nand U10721 (N_10721,N_8917,N_7640);
or U10722 (N_10722,N_9952,N_6166);
nor U10723 (N_10723,N_8918,N_9063);
or U10724 (N_10724,N_8108,N_9407);
nand U10725 (N_10725,N_6643,N_9334);
and U10726 (N_10726,N_6181,N_6208);
or U10727 (N_10727,N_5895,N_9763);
and U10728 (N_10728,N_9598,N_7119);
xor U10729 (N_10729,N_6017,N_7446);
and U10730 (N_10730,N_8631,N_9311);
and U10731 (N_10731,N_8923,N_8456);
nand U10732 (N_10732,N_7663,N_6713);
or U10733 (N_10733,N_6160,N_8586);
and U10734 (N_10734,N_5315,N_6897);
or U10735 (N_10735,N_8890,N_7056);
or U10736 (N_10736,N_8280,N_6087);
xor U10737 (N_10737,N_5594,N_6511);
nand U10738 (N_10738,N_5074,N_9223);
or U10739 (N_10739,N_6980,N_6060);
and U10740 (N_10740,N_5599,N_7792);
or U10741 (N_10741,N_9937,N_8804);
nand U10742 (N_10742,N_6292,N_8247);
or U10743 (N_10743,N_9084,N_6473);
xor U10744 (N_10744,N_9724,N_5865);
nand U10745 (N_10745,N_6588,N_7124);
or U10746 (N_10746,N_6225,N_9682);
or U10747 (N_10747,N_7036,N_8344);
and U10748 (N_10748,N_8206,N_7988);
nand U10749 (N_10749,N_5647,N_7136);
xnor U10750 (N_10750,N_7789,N_9594);
or U10751 (N_10751,N_6666,N_6041);
and U10752 (N_10752,N_9917,N_6400);
and U10753 (N_10753,N_7841,N_7042);
or U10754 (N_10754,N_5139,N_8320);
and U10755 (N_10755,N_8618,N_5133);
nand U10756 (N_10756,N_7565,N_5501);
nand U10757 (N_10757,N_9346,N_6172);
and U10758 (N_10758,N_9934,N_9757);
or U10759 (N_10759,N_7021,N_8141);
or U10760 (N_10760,N_8298,N_8409);
and U10761 (N_10761,N_5127,N_8904);
nand U10762 (N_10762,N_9625,N_5294);
nor U10763 (N_10763,N_6466,N_9371);
nor U10764 (N_10764,N_9722,N_6244);
and U10765 (N_10765,N_9195,N_7253);
nor U10766 (N_10766,N_5694,N_8860);
nor U10767 (N_10767,N_7845,N_9826);
nand U10768 (N_10768,N_5387,N_6962);
or U10769 (N_10769,N_7760,N_6776);
and U10770 (N_10770,N_9716,N_5684);
xnor U10771 (N_10771,N_6130,N_9850);
nand U10772 (N_10772,N_8788,N_7419);
and U10773 (N_10773,N_8077,N_8485);
and U10774 (N_10774,N_7809,N_9255);
nand U10775 (N_10775,N_5424,N_8356);
xnor U10776 (N_10776,N_6763,N_5576);
and U10777 (N_10777,N_7680,N_5409);
nor U10778 (N_10778,N_9411,N_8648);
and U10779 (N_10779,N_5404,N_5758);
nor U10780 (N_10780,N_8560,N_9739);
and U10781 (N_10781,N_6534,N_5024);
nand U10782 (N_10782,N_8984,N_9171);
nand U10783 (N_10783,N_9296,N_7626);
nor U10784 (N_10784,N_6488,N_8567);
nor U10785 (N_10785,N_6730,N_8795);
and U10786 (N_10786,N_6949,N_8444);
nand U10787 (N_10787,N_8668,N_9041);
nand U10788 (N_10788,N_6484,N_9532);
nor U10789 (N_10789,N_7362,N_9778);
nor U10790 (N_10790,N_6945,N_9344);
xor U10791 (N_10791,N_6742,N_8692);
xnor U10792 (N_10792,N_5871,N_6356);
nand U10793 (N_10793,N_9521,N_7507);
nor U10794 (N_10794,N_6141,N_5303);
and U10795 (N_10795,N_7332,N_8371);
or U10796 (N_10796,N_9863,N_8888);
and U10797 (N_10797,N_9989,N_5121);
or U10798 (N_10798,N_8433,N_9662);
xor U10799 (N_10799,N_7202,N_5188);
nand U10800 (N_10800,N_9430,N_7968);
xor U10801 (N_10801,N_8508,N_9495);
and U10802 (N_10802,N_9925,N_9026);
or U10803 (N_10803,N_5720,N_7768);
or U10804 (N_10804,N_9481,N_7704);
or U10805 (N_10805,N_9833,N_6422);
nor U10806 (N_10806,N_6209,N_5031);
nor U10807 (N_10807,N_9470,N_9997);
or U10808 (N_10808,N_5147,N_5380);
nand U10809 (N_10809,N_6015,N_6748);
nor U10810 (N_10810,N_8051,N_7618);
and U10811 (N_10811,N_8235,N_6393);
and U10812 (N_10812,N_6869,N_6383);
xnor U10813 (N_10813,N_9814,N_9154);
xnor U10814 (N_10814,N_7267,N_7569);
nor U10815 (N_10815,N_7594,N_9825);
xnor U10816 (N_10816,N_6929,N_5340);
or U10817 (N_10817,N_5737,N_8153);
nand U10818 (N_10818,N_6862,N_7749);
xor U10819 (N_10819,N_5915,N_8002);
nand U10820 (N_10820,N_5181,N_6661);
nor U10821 (N_10821,N_6729,N_6440);
or U10822 (N_10822,N_5803,N_6764);
and U10823 (N_10823,N_9790,N_7379);
nand U10824 (N_10824,N_6942,N_7567);
and U10825 (N_10825,N_8231,N_8160);
or U10826 (N_10826,N_9218,N_7584);
nor U10827 (N_10827,N_8698,N_7817);
nor U10828 (N_10828,N_5095,N_6977);
or U10829 (N_10829,N_8681,N_6761);
nand U10830 (N_10830,N_7600,N_6068);
xor U10831 (N_10831,N_7639,N_5917);
nand U10832 (N_10832,N_8750,N_5877);
xor U10833 (N_10833,N_9458,N_8598);
nor U10834 (N_10834,N_8142,N_9295);
or U10835 (N_10835,N_5814,N_6611);
nand U10836 (N_10836,N_6882,N_5334);
nand U10837 (N_10837,N_6078,N_5035);
or U10838 (N_10838,N_8558,N_7947);
xnor U10839 (N_10839,N_7631,N_8613);
xnor U10840 (N_10840,N_8385,N_8005);
nor U10841 (N_10841,N_5600,N_5454);
nand U10842 (N_10842,N_7916,N_5267);
nor U10843 (N_10843,N_9830,N_5683);
and U10844 (N_10844,N_5792,N_5724);
nor U10845 (N_10845,N_5847,N_9461);
and U10846 (N_10846,N_6110,N_5726);
or U10847 (N_10847,N_6481,N_7487);
nand U10848 (N_10848,N_7128,N_6707);
and U10849 (N_10849,N_9136,N_5498);
or U10850 (N_10850,N_7997,N_7602);
xnor U10851 (N_10851,N_8246,N_5697);
nor U10852 (N_10852,N_8958,N_5295);
xnor U10853 (N_10853,N_6088,N_8459);
xor U10854 (N_10854,N_7578,N_6433);
or U10855 (N_10855,N_7198,N_7492);
nand U10856 (N_10856,N_9044,N_6922);
nand U10857 (N_10857,N_7114,N_9969);
nor U10858 (N_10858,N_8124,N_5951);
xnor U10859 (N_10859,N_7829,N_6293);
xor U10860 (N_10860,N_6056,N_7647);
or U10861 (N_10861,N_5216,N_8020);
xnor U10862 (N_10862,N_5372,N_9524);
or U10863 (N_10863,N_6048,N_9317);
or U10864 (N_10864,N_9082,N_8411);
and U10865 (N_10865,N_8381,N_6974);
xor U10866 (N_10866,N_5995,N_7946);
nor U10867 (N_10867,N_7676,N_9094);
and U10868 (N_10868,N_5768,N_6627);
xnor U10869 (N_10869,N_6676,N_7135);
or U10870 (N_10870,N_7951,N_5643);
and U10871 (N_10871,N_9329,N_8605);
or U10872 (N_10872,N_6971,N_8873);
nand U10873 (N_10873,N_7867,N_8637);
nor U10874 (N_10874,N_8532,N_7422);
nor U10875 (N_10875,N_9378,N_5551);
nor U10876 (N_10876,N_7195,N_5149);
and U10877 (N_10877,N_5207,N_7375);
and U10878 (N_10878,N_7763,N_5171);
or U10879 (N_10879,N_9023,N_9809);
nand U10880 (N_10880,N_7483,N_8883);
and U10881 (N_10881,N_9636,N_5563);
or U10882 (N_10882,N_5754,N_5013);
nand U10883 (N_10883,N_6600,N_5011);
nor U10884 (N_10884,N_7098,N_5231);
nand U10885 (N_10885,N_7361,N_8037);
nor U10886 (N_10886,N_8562,N_9637);
nand U10887 (N_10887,N_5473,N_9110);
nand U10888 (N_10888,N_7690,N_6263);
or U10889 (N_10889,N_9664,N_8747);
or U10890 (N_10890,N_7351,N_8886);
nor U10891 (N_10891,N_5215,N_8115);
nand U10892 (N_10892,N_8099,N_8033);
or U10893 (N_10893,N_5778,N_6080);
xor U10894 (N_10894,N_9746,N_9659);
nand U10895 (N_10895,N_8528,N_6515);
nor U10896 (N_10896,N_5019,N_8490);
nand U10897 (N_10897,N_8487,N_8435);
xnor U10898 (N_10898,N_7247,N_9867);
xnor U10899 (N_10899,N_9806,N_8851);
and U10900 (N_10900,N_9587,N_7068);
and U10901 (N_10901,N_6005,N_8857);
nor U10902 (N_10902,N_5901,N_8650);
xor U10903 (N_10903,N_5676,N_6050);
xnor U10904 (N_10904,N_8263,N_6379);
xor U10905 (N_10905,N_5670,N_5736);
or U10906 (N_10906,N_6248,N_8237);
nand U10907 (N_10907,N_9405,N_9479);
and U10908 (N_10908,N_6790,N_5978);
or U10909 (N_10909,N_8810,N_7813);
xor U10910 (N_10910,N_5004,N_5725);
and U10911 (N_10911,N_6337,N_5278);
nand U10912 (N_10912,N_8664,N_8719);
nor U10913 (N_10913,N_7189,N_5348);
and U10914 (N_10914,N_5490,N_5932);
nor U10915 (N_10915,N_9516,N_8018);
nand U10916 (N_10916,N_9193,N_9987);
nand U10917 (N_10917,N_8939,N_7005);
and U10918 (N_10918,N_5213,N_8201);
or U10919 (N_10919,N_6562,N_9277);
nor U10920 (N_10920,N_8688,N_9504);
nand U10921 (N_10921,N_5318,N_9995);
or U10922 (N_10922,N_8794,N_7087);
nor U10923 (N_10923,N_7293,N_9891);
and U10924 (N_10924,N_7811,N_5554);
and U10925 (N_10925,N_9020,N_5417);
and U10926 (N_10926,N_6233,N_6963);
nor U10927 (N_10927,N_6345,N_7502);
nor U10928 (N_10928,N_8898,N_6738);
and U10929 (N_10929,N_7000,N_5703);
and U10930 (N_10930,N_8695,N_7781);
xnor U10931 (N_10931,N_7301,N_9202);
and U10932 (N_10932,N_6517,N_5286);
xor U10933 (N_10933,N_5636,N_5385);
nor U10934 (N_10934,N_7089,N_6023);
xnor U10935 (N_10935,N_8821,N_7729);
and U10936 (N_10936,N_8465,N_6107);
nor U10937 (N_10937,N_6968,N_8544);
nand U10938 (N_10938,N_9543,N_7066);
nor U10939 (N_10939,N_8707,N_7648);
nor U10940 (N_10940,N_6094,N_5519);
xnor U10941 (N_10941,N_8226,N_9126);
or U10942 (N_10942,N_9541,N_6775);
nand U10943 (N_10943,N_8331,N_8629);
nand U10944 (N_10944,N_5319,N_7844);
nor U10945 (N_10945,N_7624,N_5730);
nor U10946 (N_10946,N_7073,N_7183);
or U10947 (N_10947,N_6658,N_9004);
and U10948 (N_10948,N_8557,N_6835);
or U10949 (N_10949,N_9775,N_9439);
nor U10950 (N_10950,N_5751,N_6565);
or U10951 (N_10951,N_6182,N_8803);
nand U10952 (N_10952,N_8522,N_9234);
and U10953 (N_10953,N_8739,N_6958);
or U10954 (N_10954,N_9707,N_9549);
and U10955 (N_10955,N_8285,N_6033);
nand U10956 (N_10956,N_6186,N_7131);
nand U10957 (N_10957,N_5203,N_5015);
xor U10958 (N_10958,N_8039,N_5680);
and U10959 (N_10959,N_6989,N_7609);
nor U10960 (N_10960,N_8414,N_6480);
xnor U10961 (N_10961,N_6563,N_7629);
and U10962 (N_10962,N_5491,N_5328);
or U10963 (N_10963,N_9173,N_5898);
or U10964 (N_10964,N_6230,N_8609);
xnor U10965 (N_10965,N_8437,N_7512);
nand U10966 (N_10966,N_9113,N_9655);
xor U10967 (N_10967,N_7619,N_7397);
and U10968 (N_10968,N_7866,N_9244);
or U10969 (N_10969,N_8583,N_9762);
nand U10970 (N_10970,N_7757,N_7169);
nor U10971 (N_10971,N_5933,N_8705);
nand U10972 (N_10972,N_6545,N_7903);
xnor U10973 (N_10973,N_9431,N_5256);
nand U10974 (N_10974,N_5113,N_7820);
and U10975 (N_10975,N_5870,N_9815);
xor U10976 (N_10976,N_9836,N_8170);
nand U10977 (N_10977,N_5217,N_7380);
xor U10978 (N_10978,N_7715,N_6512);
nand U10979 (N_10979,N_7280,N_7571);
nand U10980 (N_10980,N_7333,N_8333);
or U10981 (N_10981,N_9304,N_9824);
xnor U10982 (N_10982,N_6011,N_7611);
and U10983 (N_10983,N_6361,N_6606);
or U10984 (N_10984,N_6547,N_5451);
nor U10985 (N_10985,N_6102,N_9671);
nand U10986 (N_10986,N_5530,N_6628);
and U10987 (N_10987,N_7539,N_5431);
nor U10988 (N_10988,N_7358,N_8079);
nor U10989 (N_10989,N_6490,N_6453);
xnor U10990 (N_10990,N_6795,N_9022);
or U10991 (N_10991,N_8645,N_9914);
and U10992 (N_10992,N_8420,N_7415);
and U10993 (N_10993,N_7355,N_5441);
nor U10994 (N_10994,N_8133,N_6759);
and U10995 (N_10995,N_7522,N_5259);
and U10996 (N_10996,N_5349,N_8661);
nand U10997 (N_10997,N_8094,N_6280);
nor U10998 (N_10998,N_9737,N_5503);
or U10999 (N_10999,N_9290,N_9155);
or U11000 (N_11000,N_9245,N_5955);
xnor U11001 (N_11001,N_9661,N_8966);
nand U11002 (N_11002,N_8962,N_5069);
xnor U11003 (N_11003,N_7104,N_5201);
nand U11004 (N_11004,N_7109,N_7581);
or U11005 (N_11005,N_5826,N_9975);
nand U11006 (N_11006,N_5308,N_8488);
xor U11007 (N_11007,N_6014,N_9351);
and U11008 (N_11008,N_6065,N_6308);
xnor U11009 (N_11009,N_8992,N_6114);
and U11010 (N_11010,N_7256,N_8264);
and U11011 (N_11011,N_6799,N_7959);
or U11012 (N_11012,N_6538,N_7656);
and U11013 (N_11013,N_7182,N_9846);
and U11014 (N_11014,N_5071,N_8517);
xnor U11015 (N_11015,N_6273,N_8797);
or U11016 (N_11016,N_6772,N_6918);
or U11017 (N_11017,N_5505,N_8310);
and U11018 (N_11018,N_5893,N_5671);
xnor U11019 (N_11019,N_8165,N_7024);
nor U11020 (N_11020,N_9738,N_9733);
nand U11021 (N_11021,N_9964,N_9251);
xor U11022 (N_11022,N_8943,N_9297);
nor U11023 (N_11023,N_9101,N_9998);
xnor U11024 (N_11024,N_9119,N_9379);
nand U11025 (N_11025,N_7726,N_7337);
and U11026 (N_11026,N_5882,N_7591);
or U11027 (N_11027,N_7590,N_9702);
and U11028 (N_11028,N_6384,N_6577);
nand U11029 (N_11029,N_8956,N_5050);
and U11030 (N_11030,N_8896,N_7048);
or U11031 (N_11031,N_6333,N_5122);
xnor U11032 (N_11032,N_9212,N_6027);
nand U11033 (N_11033,N_7461,N_8375);
nand U11034 (N_11034,N_6266,N_8727);
or U11035 (N_11035,N_7155,N_6857);
nand U11036 (N_11036,N_5141,N_7798);
nand U11037 (N_11037,N_7287,N_8085);
or U11038 (N_11038,N_9967,N_7765);
nand U11039 (N_11039,N_9112,N_6032);
and U11040 (N_11040,N_6410,N_8816);
or U11041 (N_11041,N_7669,N_5897);
or U11042 (N_11042,N_7880,N_8925);
or U11043 (N_11043,N_5843,N_9456);
xor U11044 (N_11044,N_9465,N_5257);
nand U11045 (N_11045,N_7307,N_5475);
xor U11046 (N_11046,N_7142,N_9741);
nand U11047 (N_11047,N_5830,N_7925);
nor U11048 (N_11048,N_7127,N_9921);
xnor U11049 (N_11049,N_5427,N_9856);
nor U11050 (N_11050,N_9302,N_8258);
or U11051 (N_11051,N_6461,N_5894);
nand U11052 (N_11052,N_9129,N_9574);
nand U11053 (N_11053,N_5283,N_9009);
xor U11054 (N_11054,N_5049,N_8207);
or U11055 (N_11055,N_9335,N_9079);
and U11056 (N_11056,N_6901,N_9821);
xnor U11057 (N_11057,N_7922,N_6822);
or U11058 (N_11058,N_9766,N_5769);
nand U11059 (N_11059,N_7941,N_9877);
nand U11060 (N_11060,N_8338,N_9150);
nor U11061 (N_11061,N_6725,N_8225);
or U11062 (N_11062,N_7956,N_9271);
and U11063 (N_11063,N_5509,N_7085);
and U11064 (N_11064,N_6625,N_7621);
nand U11065 (N_11065,N_5616,N_7496);
or U11066 (N_11066,N_5629,N_5442);
nor U11067 (N_11067,N_7166,N_7814);
and U11068 (N_11068,N_8445,N_5206);
and U11069 (N_11069,N_6346,N_8450);
nand U11070 (N_11070,N_5137,N_7955);
nor U11071 (N_11071,N_9070,N_8230);
nor U11072 (N_11072,N_5495,N_7092);
nor U11073 (N_11073,N_6539,N_7737);
xor U11074 (N_11074,N_7044,N_6449);
nor U11075 (N_11075,N_8205,N_5538);
xnor U11076 (N_11076,N_9838,N_6816);
nand U11077 (N_11077,N_5212,N_9175);
or U11078 (N_11078,N_5221,N_8227);
nand U11079 (N_11079,N_6201,N_9399);
nand U11080 (N_11080,N_7445,N_6126);
xnor U11081 (N_11081,N_5460,N_8852);
xor U11082 (N_11082,N_8734,N_9415);
or U11083 (N_11083,N_6149,N_7633);
or U11084 (N_11084,N_5144,N_9332);
and U11085 (N_11085,N_8600,N_5774);
xnor U11086 (N_11086,N_8876,N_9608);
or U11087 (N_11087,N_5060,N_6168);
nor U11088 (N_11088,N_9051,N_5449);
xor U11089 (N_11089,N_7575,N_7420);
or U11090 (N_11090,N_7720,N_9350);
xnor U11091 (N_11091,N_5555,N_5688);
xor U11092 (N_11092,N_7153,N_6644);
or U11093 (N_11093,N_9805,N_8307);
nor U11094 (N_11094,N_8423,N_7032);
nor U11095 (N_11095,N_9508,N_5436);
xnor U11096 (N_11096,N_7685,N_6680);
xnor U11097 (N_11097,N_7635,N_7898);
xor U11098 (N_11098,N_6733,N_7560);
nand U11099 (N_11099,N_8251,N_8579);
or U11100 (N_11100,N_8242,N_6589);
nor U11101 (N_11101,N_8136,N_7262);
xnor U11102 (N_11102,N_7465,N_8533);
xnor U11103 (N_11103,N_6095,N_7288);
nand U11104 (N_11104,N_8172,N_7309);
and U11105 (N_11105,N_7008,N_9086);
xor U11106 (N_11106,N_6282,N_8983);
xor U11107 (N_11107,N_6852,N_9901);
and U11108 (N_11108,N_9729,N_8685);
and U11109 (N_11109,N_6717,N_7906);
or U11110 (N_11110,N_6668,N_8620);
or U11111 (N_11111,N_8213,N_9777);
nand U11112 (N_11112,N_6030,N_7184);
and U11113 (N_11113,N_8377,N_9576);
and U11114 (N_11114,N_7228,N_5515);
or U11115 (N_11115,N_6134,N_5214);
xor U11116 (N_11116,N_5746,N_9174);
nand U11117 (N_11117,N_8689,N_8548);
nand U11118 (N_11118,N_9455,N_6701);
and U11119 (N_11119,N_5853,N_7148);
nor U11120 (N_11120,N_5527,N_8054);
nand U11121 (N_11121,N_9828,N_8432);
nor U11122 (N_11122,N_5763,N_7853);
and U11123 (N_11123,N_7642,N_8275);
or U11124 (N_11124,N_8539,N_8271);
and U11125 (N_11125,N_9527,N_9795);
nand U11126 (N_11126,N_9754,N_8897);
xnor U11127 (N_11127,N_8615,N_7381);
and U11128 (N_11128,N_8044,N_9076);
nor U11129 (N_11129,N_7517,N_9887);
nand U11130 (N_11130,N_5885,N_9247);
or U11131 (N_11131,N_5999,N_8040);
and U11132 (N_11132,N_6530,N_8425);
and U11133 (N_11133,N_8089,N_5940);
or U11134 (N_11134,N_9801,N_7665);
or U11135 (N_11135,N_7278,N_8882);
xor U11136 (N_11136,N_9188,N_8337);
nor U11137 (N_11137,N_5965,N_9349);
and U11138 (N_11138,N_6766,N_9552);
xor U11139 (N_11139,N_8665,N_9691);
xor U11140 (N_11140,N_8809,N_7598);
xnor U11141 (N_11141,N_6460,N_5962);
or U11142 (N_11142,N_5110,N_7238);
or U11143 (N_11143,N_7129,N_6416);
and U11144 (N_11144,N_8023,N_8318);
or U11145 (N_11145,N_5321,N_9485);
nand U11146 (N_11146,N_9280,N_5131);
nand U11147 (N_11147,N_6421,N_9514);
xnor U11148 (N_11148,N_7529,N_9512);
and U11149 (N_11149,N_7191,N_8772);
and U11150 (N_11150,N_7054,N_7241);
xnor U11151 (N_11151,N_5169,N_5255);
or U11152 (N_11152,N_9536,N_7038);
nand U11153 (N_11153,N_8762,N_5038);
xor U11154 (N_11154,N_9853,N_8090);
nor U11155 (N_11155,N_6192,N_6636);
and U11156 (N_11156,N_7011,N_8199);
xnor U11157 (N_11157,N_7077,N_5242);
nand U11158 (N_11158,N_9164,N_5471);
or U11159 (N_11159,N_8048,N_8454);
nand U11160 (N_11160,N_7353,N_5375);
or U11161 (N_11161,N_7018,N_7033);
nor U11162 (N_11162,N_6930,N_6617);
and U11163 (N_11163,N_7482,N_9264);
or U11164 (N_11164,N_5653,N_8221);
and U11165 (N_11165,N_6662,N_5391);
nand U11166 (N_11166,N_5970,N_6779);
nor U11167 (N_11167,N_8369,N_9231);
nor U11168 (N_11168,N_6210,N_9808);
nand U11169 (N_11169,N_6714,N_8416);
nand U11170 (N_11170,N_8072,N_5570);
nand U11171 (N_11171,N_5400,N_6504);
nor U11172 (N_11172,N_5352,N_8742);
or U11173 (N_11173,N_6656,N_6850);
nor U11174 (N_11174,N_7692,N_8120);
nor U11175 (N_11175,N_9488,N_5916);
nand U11176 (N_11176,N_7395,N_8697);
and U11177 (N_11177,N_8283,N_8282);
and U11178 (N_11178,N_8348,N_7194);
nand U11179 (N_11179,N_5253,N_7269);
nand U11180 (N_11180,N_8679,N_5535);
nand U11181 (N_11181,N_5638,N_5511);
nor U11182 (N_11182,N_5017,N_9301);
or U11183 (N_11183,N_8849,N_8855);
or U11184 (N_11184,N_5222,N_7555);
or U11185 (N_11185,N_7745,N_5225);
xnor U11186 (N_11186,N_5356,N_9237);
and U11187 (N_11187,N_6058,N_8957);
nand U11188 (N_11188,N_5184,N_7797);
nand U11189 (N_11189,N_7767,N_7188);
nor U11190 (N_11190,N_6966,N_6593);
nor U11191 (N_11191,N_9611,N_8458);
xnor U11192 (N_11192,N_7020,N_6594);
nor U11193 (N_11193,N_9677,N_9890);
and U11194 (N_11194,N_9609,N_5876);
nor U11195 (N_11195,N_9767,N_8767);
and U11196 (N_11196,N_7480,N_6810);
and U11197 (N_11197,N_8008,N_5799);
nand U11198 (N_11198,N_8157,N_6197);
xnor U11199 (N_11199,N_6514,N_7756);
or U11200 (N_11200,N_7981,N_5860);
or U11201 (N_11201,N_7110,N_5790);
nand U11202 (N_11202,N_7210,N_7965);
xnor U11203 (N_11203,N_6670,N_9016);
or U11204 (N_11204,N_5130,N_9817);
xnor U11205 (N_11205,N_6382,N_9648);
xor U11206 (N_11206,N_5663,N_8202);
xnor U11207 (N_11207,N_7678,N_8046);
or U11208 (N_11208,N_9822,N_6526);
nand U11209 (N_11209,N_6868,N_7323);
and U11210 (N_11210,N_7649,N_9915);
xnor U11211 (N_11211,N_9950,N_6664);
or U11212 (N_11212,N_9798,N_8482);
or U11213 (N_11213,N_8004,N_7738);
or U11214 (N_11214,N_9075,N_6831);
nor U11215 (N_11215,N_9434,N_5301);
nor U11216 (N_11216,N_6133,N_5260);
nor U11217 (N_11217,N_6367,N_6815);
and U11218 (N_11218,N_8972,N_8389);
nor U11219 (N_11219,N_5118,N_7437);
nor U11220 (N_11220,N_5789,N_9322);
and U11221 (N_11221,N_5094,N_7022);
xor U11222 (N_11222,N_9466,N_6121);
nor U11223 (N_11223,N_6207,N_8780);
and U11224 (N_11224,N_5313,N_5388);
and U11225 (N_11225,N_5607,N_8470);
xnor U11226 (N_11226,N_9447,N_5332);
nor U11227 (N_11227,N_7462,N_7257);
and U11228 (N_11228,N_7605,N_5904);
xnor U11229 (N_11229,N_9133,N_6250);
and U11230 (N_11230,N_5875,N_6334);
or U11231 (N_11231,N_6359,N_5561);
nand U11232 (N_11232,N_7439,N_5627);
nand U11233 (N_11233,N_9377,N_5807);
nor U11234 (N_11234,N_9540,N_9505);
nand U11235 (N_11235,N_8290,N_6362);
or U11236 (N_11236,N_5399,N_9693);
and U11237 (N_11237,N_8034,N_6540);
or U11238 (N_11238,N_5085,N_8155);
xor U11239 (N_11239,N_5066,N_8475);
nand U11240 (N_11240,N_5040,N_5514);
nand U11241 (N_11241,N_7535,N_7926);
or U11242 (N_11242,N_9257,N_9414);
nand U11243 (N_11243,N_5623,N_9186);
nor U11244 (N_11244,N_8779,N_8922);
nor U11245 (N_11245,N_8850,N_9668);
and U11246 (N_11246,N_9949,N_5818);
and U11247 (N_11247,N_8663,N_5363);
nand U11248 (N_11248,N_5766,N_8240);
and U11249 (N_11249,N_9721,N_5795);
and U11250 (N_11250,N_5549,N_7670);
nand U11251 (N_11251,N_5151,N_8186);
xor U11252 (N_11252,N_9570,N_5007);
xnor U11253 (N_11253,N_7336,N_7174);
xnor U11254 (N_11254,N_6981,N_6234);
and U11255 (N_11255,N_8216,N_5985);
xnor U11256 (N_11256,N_9876,N_5000);
nand U11257 (N_11257,N_7545,N_8228);
or U11258 (N_11258,N_5158,N_5080);
and U11259 (N_11259,N_6700,N_9156);
and U11260 (N_11260,N_9443,N_9402);
or U11261 (N_11261,N_9926,N_9353);
nand U11262 (N_11262,N_8150,N_6754);
nor U11263 (N_11263,N_6592,N_7927);
nand U11264 (N_11264,N_7689,N_8217);
and U11265 (N_11265,N_6351,N_7471);
and U11266 (N_11266,N_7493,N_6814);
nor U11267 (N_11267,N_9398,N_7343);
nand U11268 (N_11268,N_9872,N_5695);
nor U11269 (N_11269,N_6045,N_7871);
xnor U11270 (N_11270,N_5883,N_7405);
nor U11271 (N_11271,N_8364,N_9382);
nand U11272 (N_11272,N_6189,N_6247);
nand U11273 (N_11273,N_5907,N_5299);
nor U11274 (N_11274,N_6441,N_6276);
nand U11275 (N_11275,N_9928,N_6704);
or U11276 (N_11276,N_8678,N_9813);
nor U11277 (N_11277,N_6152,N_9014);
nand U11278 (N_11278,N_5659,N_8936);
nor U11279 (N_11279,N_5862,N_7279);
and U11280 (N_11280,N_8982,N_9962);
xnor U11281 (N_11281,N_6198,N_8326);
xor U11282 (N_11282,N_9670,N_9620);
and U11283 (N_11283,N_9061,N_8974);
xnor U11284 (N_11284,N_5073,N_6659);
xnor U11285 (N_11285,N_9954,N_8109);
or U11286 (N_11286,N_7952,N_8061);
and U11287 (N_11287,N_8178,N_8765);
and U11288 (N_11288,N_9342,N_5827);
xnor U11289 (N_11289,N_6734,N_6691);
or U11290 (N_11290,N_6115,N_6265);
xnor U11291 (N_11291,N_9445,N_6279);
and U11292 (N_11292,N_8229,N_8604);
and U11293 (N_11293,N_7890,N_6062);
or U11294 (N_11294,N_9006,N_8910);
or U11295 (N_11295,N_5101,N_6378);
and U11296 (N_11296,N_5575,N_5528);
nand U11297 (N_11297,N_6077,N_8253);
or U11298 (N_11298,N_6765,N_5896);
and U11299 (N_11299,N_6893,N_7973);
xor U11300 (N_11300,N_9530,N_9183);
or U11301 (N_11301,N_7138,N_9130);
xor U11302 (N_11302,N_8676,N_6408);
nor U11303 (N_11303,N_5195,N_5170);
or U11304 (N_11304,N_7311,N_9565);
xnor U11305 (N_11305,N_5854,N_7837);
xor U11306 (N_11306,N_7053,N_9904);
nor U11307 (N_11307,N_5178,N_7334);
or U11308 (N_11308,N_7231,N_9641);
nor U11309 (N_11309,N_5324,N_5994);
nand U11310 (N_11310,N_5631,N_9312);
nand U11311 (N_11311,N_6687,N_6191);
or U11312 (N_11312,N_7010,N_5284);
and U11313 (N_11313,N_5497,N_6119);
and U11314 (N_11314,N_9091,N_6309);
nand U11315 (N_11315,N_8503,N_6313);
or U11316 (N_11316,N_6407,N_9784);
xnor U11317 (N_11317,N_5395,N_5606);
xnor U11318 (N_11318,N_8148,N_8989);
nand U11319 (N_11319,N_9327,N_9918);
nor U11320 (N_11320,N_9034,N_8838);
nand U11321 (N_11321,N_7444,N_6727);
or U11322 (N_11322,N_6649,N_5477);
nor U11323 (N_11323,N_6631,N_9315);
xnor U11324 (N_11324,N_5959,N_5840);
nand U11325 (N_11325,N_5087,N_9772);
nor U11326 (N_11326,N_5448,N_6338);
or U11327 (N_11327,N_6771,N_8603);
xnor U11328 (N_11328,N_5043,N_5821);
and U11329 (N_11329,N_9616,N_8107);
xor U11330 (N_11330,N_8215,N_8438);
nand U11331 (N_11331,N_9065,N_9203);
nor U11332 (N_11332,N_9971,N_8446);
xor U11333 (N_11333,N_6369,N_8440);
and U11334 (N_11334,N_6289,N_7126);
nor U11335 (N_11335,N_6464,N_9058);
nor U11336 (N_11336,N_5928,N_6960);
xnor U11337 (N_11337,N_6003,N_5771);
or U11338 (N_11338,N_8826,N_9441);
and U11339 (N_11339,N_8768,N_5981);
or U11340 (N_11340,N_7900,N_8501);
xnor U11341 (N_11341,N_5088,N_6745);
or U11342 (N_11342,N_7808,N_6685);
nand U11343 (N_11343,N_8097,N_5569);
xor U11344 (N_11344,N_6004,N_9900);
or U11345 (N_11345,N_8564,N_5866);
nor U11346 (N_11346,N_8473,N_6435);
and U11347 (N_11347,N_7586,N_9910);
or U11348 (N_11348,N_8667,N_6098);
and U11349 (N_11349,N_7025,N_5119);
nor U11350 (N_11350,N_9137,N_6546);
and U11351 (N_11351,N_8193,N_9116);
nor U11352 (N_11352,N_6327,N_9569);
and U11353 (N_11353,N_9209,N_9740);
and U11354 (N_11354,N_5742,N_5619);
or U11355 (N_11355,N_9732,N_5500);
or U11356 (N_11356,N_7577,N_5016);
and U11357 (N_11357,N_8341,N_6943);
nand U11358 (N_11358,N_5439,N_5592);
nand U11359 (N_11359,N_9357,N_5037);
nor U11360 (N_11360,N_6245,N_6485);
or U11361 (N_11361,N_5189,N_7236);
xnor U11362 (N_11362,N_6206,N_7106);
and U11363 (N_11363,N_9704,N_9553);
xor U11364 (N_11364,N_5558,N_9028);
nor U11365 (N_11365,N_9370,N_9356);
nand U11366 (N_11366,N_6039,N_8047);
nor U11367 (N_11367,N_6885,N_5034);
nor U11368 (N_11368,N_8773,N_6489);
nor U11369 (N_11369,N_5156,N_9678);
and U11370 (N_11370,N_6632,N_8774);
nand U11371 (N_11371,N_7103,N_8415);
or U11372 (N_11372,N_5914,N_8585);
nor U11373 (N_11373,N_9308,N_5086);
or U11374 (N_11374,N_5243,N_8030);
nor U11375 (N_11375,N_7075,N_8981);
xnor U11376 (N_11376,N_7683,N_6807);
nor U11377 (N_11377,N_6165,N_6148);
xnor U11378 (N_11378,N_8493,N_8071);
and U11379 (N_11379,N_8149,N_8552);
nand U11380 (N_11380,N_8419,N_7475);
nor U11381 (N_11381,N_5532,N_5027);
nand U11382 (N_11382,N_9067,N_7093);
nand U11383 (N_11383,N_5472,N_7904);
nand U11384 (N_11384,N_5093,N_8311);
nand U11385 (N_11385,N_8672,N_9253);
nand U11386 (N_11386,N_5655,N_5199);
xor U11387 (N_11387,N_7175,N_7476);
nor U11388 (N_11388,N_5639,N_7830);
nand U11389 (N_11389,N_9469,N_5227);
and U11390 (N_11390,N_7877,N_9566);
nand U11391 (N_11391,N_7975,N_9564);
nor U11392 (N_11392,N_9776,N_6803);
nor U11393 (N_11393,N_8647,N_8840);
nor U11394 (N_11394,N_7840,N_9638);
xnor U11395 (N_11395,N_8606,N_6794);
xnor U11396 (N_11396,N_7620,N_8463);
xnor U11397 (N_11397,N_8612,N_7677);
nor U11398 (N_11398,N_7002,N_6641);
nor U11399 (N_11399,N_5852,N_6518);
nand U11400 (N_11400,N_6735,N_6861);
xnor U11401 (N_11401,N_8682,N_7999);
and U11402 (N_11402,N_8820,N_5718);
and U11403 (N_11403,N_6492,N_5062);
nand U11404 (N_11404,N_6161,N_5634);
and U11405 (N_11405,N_7971,N_5338);
and U11406 (N_11406,N_5838,N_6419);
nand U11407 (N_11407,N_9796,N_5878);
nor U11408 (N_11408,N_7319,N_8700);
nor U11409 (N_11409,N_5583,N_7913);
nor U11410 (N_11410,N_5272,N_6886);
nor U11411 (N_11411,N_7964,N_9007);
xor U11412 (N_11412,N_5523,N_8350);
and U11413 (N_11413,N_8776,N_5817);
and U11414 (N_11414,N_6944,N_7942);
nand U11415 (N_11415,N_5846,N_6079);
or U11416 (N_11416,N_8813,N_5645);
and U11417 (N_11417,N_9764,N_8980);
nor U11418 (N_11418,N_8801,N_9015);
or U11419 (N_11419,N_5783,N_7873);
or U11420 (N_11420,N_9268,N_7812);
nand U11421 (N_11421,N_9882,N_7693);
nand U11422 (N_11422,N_7860,N_5884);
or U11423 (N_11423,N_9274,N_5811);
and U11424 (N_11424,N_9771,N_5176);
or U11425 (N_11425,N_5689,N_6159);
or U11426 (N_11426,N_8082,N_7501);
and U11427 (N_11427,N_5341,N_6811);
xnor U11428 (N_11428,N_8368,N_6386);
nand U11429 (N_11429,N_5824,N_8626);
or U11430 (N_11430,N_7707,N_8417);
xnor U11431 (N_11431,N_8814,N_5954);
and U11432 (N_11432,N_7897,N_7391);
or U11433 (N_11433,N_9886,N_8907);
and U11434 (N_11434,N_6872,N_5926);
nand U11435 (N_11435,N_8911,N_8059);
nor U11436 (N_11436,N_7286,N_6482);
nor U11437 (N_11437,N_5593,N_9748);
and U11438 (N_11438,N_6252,N_8758);
or U11439 (N_11439,N_6555,N_6465);
nor U11440 (N_11440,N_8963,N_7986);
and U11441 (N_11441,N_6424,N_7667);
nand U11442 (N_11442,N_7713,N_5661);
or U11443 (N_11443,N_8074,N_8909);
nor U11444 (N_11444,N_5874,N_9038);
or U11445 (N_11445,N_6364,N_7962);
xor U11446 (N_11446,N_9333,N_7795);
nand U11447 (N_11447,N_9829,N_7859);
and U11448 (N_11448,N_5585,N_9162);
nand U11449 (N_11449,N_5937,N_5975);
nor U11450 (N_11450,N_6837,N_7373);
or U11451 (N_11451,N_8987,N_6451);
nor U11452 (N_11452,N_6220,N_7019);
nand U11453 (N_11453,N_5264,N_6474);
and U11454 (N_11454,N_7546,N_5986);
nor U11455 (N_11455,N_9930,N_5314);
nor U11456 (N_11456,N_6813,N_5271);
or U11457 (N_11457,N_6456,N_5729);
nor U11458 (N_11458,N_7778,N_6762);
xnor U11459 (N_11459,N_6890,N_7346);
xor U11460 (N_11460,N_5759,N_5544);
or U11461 (N_11461,N_5238,N_5486);
and U11462 (N_11462,N_5633,N_5531);
nor U11463 (N_11463,N_9472,N_5009);
nand U11464 (N_11464,N_6368,N_7488);
and U11465 (N_11465,N_8701,N_6876);
nand U11466 (N_11466,N_8088,N_6912);
nor U11467 (N_11467,N_5132,N_8284);
nor U11468 (N_11468,N_7972,N_9172);
and U11469 (N_11469,N_9141,N_5732);
or U11470 (N_11470,N_6743,N_8843);
nand U11471 (N_11471,N_8439,N_5429);
or U11472 (N_11472,N_9276,N_8073);
nor U11473 (N_11473,N_8256,N_7834);
xor U11474 (N_11474,N_5344,N_9718);
and U11475 (N_11475,N_9425,N_5298);
xor U11476 (N_11476,N_9493,N_8970);
and U11477 (N_11477,N_9306,N_8365);
or U11478 (N_11478,N_9684,N_6099);
and U11479 (N_11479,N_9433,N_8624);
nand U11480 (N_11480,N_9454,N_5794);
nor U11481 (N_11481,N_7818,N_9042);
nor U11482 (N_11482,N_9947,N_5268);
nor U11483 (N_11483,N_9321,N_5573);
or U11484 (N_11484,N_8718,N_9657);
xor U11485 (N_11485,N_6875,N_8565);
or U11486 (N_11486,N_8396,N_9073);
nor U11487 (N_11487,N_7341,N_5033);
or U11488 (N_11488,N_5240,N_8222);
or U11489 (N_11489,N_5211,N_7396);
nand U11490 (N_11490,N_7923,N_6612);
nand U11491 (N_11491,N_9363,N_9689);
xor U11492 (N_11492,N_6923,N_6660);
nand U11493 (N_11493,N_7616,N_7325);
nor U11494 (N_11494,N_5772,N_6655);
xnor U11495 (N_11495,N_8819,N_8602);
or U11496 (N_11496,N_8035,N_8288);
or U11497 (N_11497,N_9993,N_6505);
or U11498 (N_11498,N_8319,N_6272);
xor U11499 (N_11499,N_5856,N_9982);
nor U11500 (N_11500,N_7940,N_6736);
nor U11501 (N_11501,N_5836,N_8064);
nor U11502 (N_11502,N_5105,N_5744);
or U11503 (N_11503,N_7004,N_6950);
xnor U11504 (N_11504,N_5466,N_8740);
and U11505 (N_11505,N_6146,N_6533);
and U11506 (N_11506,N_5699,N_7874);
nor U11507 (N_11507,N_7566,N_6525);
or U11508 (N_11508,N_6268,N_9575);
nand U11509 (N_11509,N_6983,N_9420);
and U11510 (N_11510,N_5839,N_8942);
nand U11511 (N_11511,N_5728,N_9688);
xor U11512 (N_11512,N_6397,N_9500);
and U11513 (N_11513,N_7995,N_7554);
nand U11514 (N_11514,N_5411,N_9066);
xnor U11515 (N_11515,N_7733,N_7479);
nand U11516 (N_11516,N_9694,N_6228);
or U11517 (N_11517,N_6043,N_7603);
nand U11518 (N_11518,N_5849,N_8092);
xnor U11519 (N_11519,N_7352,N_8125);
nand U11520 (N_11520,N_7485,N_7513);
xor U11521 (N_11521,N_7944,N_6954);
and U11522 (N_11522,N_5980,N_9751);
or U11523 (N_11523,N_6829,N_7615);
xor U11524 (N_11524,N_5241,N_6798);
nor U11525 (N_11525,N_8169,N_5587);
nor U11526 (N_11526,N_6204,N_7058);
and U11527 (N_11527,N_5096,N_7275);
nor U11528 (N_11528,N_6132,N_7151);
nand U11529 (N_11529,N_9697,N_8260);
and U11530 (N_11530,N_6888,N_8761);
and U11531 (N_11531,N_7744,N_9064);
nand U11532 (N_11532,N_5705,N_7980);
or U11533 (N_11533,N_8723,N_9279);
nand U11534 (N_11534,N_9473,N_7879);
or U11535 (N_11535,N_8467,N_8899);
nand U11536 (N_11536,N_7908,N_7531);
xnor U11537 (N_11537,N_6231,N_9147);
xnor U11538 (N_11538,N_9851,N_6477);
or U11539 (N_11539,N_6236,N_5539);
and U11540 (N_11540,N_9367,N_7125);
nor U11541 (N_11541,N_8214,N_5244);
and U11542 (N_11542,N_9054,N_7772);
or U11543 (N_11543,N_9358,N_5459);
xor U11544 (N_11544,N_9017,N_7220);
or U11545 (N_11545,N_9860,N_8759);
nor U11546 (N_11546,N_7698,N_5777);
xnor U11547 (N_11547,N_6749,N_8122);
nor U11548 (N_11548,N_6373,N_8870);
or U11549 (N_11549,N_9590,N_6405);
xnor U11550 (N_11550,N_6937,N_8466);
or U11551 (N_11551,N_5453,N_7748);
nand U11552 (N_11552,N_6800,N_7977);
and U11553 (N_11553,N_6906,N_5293);
nand U11554 (N_11554,N_5529,N_8616);
nor U11555 (N_11555,N_7657,N_5835);
or U11556 (N_11556,N_8504,N_9774);
nand U11557 (N_11557,N_5383,N_8478);
and U11558 (N_11558,N_6715,N_6084);
nand U11559 (N_11559,N_7967,N_6401);
or U11560 (N_11560,N_5998,N_5889);
nor U11561 (N_11561,N_6175,N_6635);
and U11562 (N_11562,N_7824,N_9978);
nand U11563 (N_11563,N_5179,N_8495);
xnor U11564 (N_11564,N_9149,N_6894);
nand U11565 (N_11565,N_5438,N_8549);
or U11566 (N_11566,N_8135,N_8403);
or U11567 (N_11567,N_6787,N_8167);
nand U11568 (N_11568,N_8836,N_9673);
or U11569 (N_11569,N_9747,N_6223);
nand U11570 (N_11570,N_7782,N_9348);
nand U11571 (N_11571,N_7062,N_8434);
or U11572 (N_11572,N_7863,N_5124);
xor U11573 (N_11573,N_8156,N_7671);
xnor U11574 (N_11574,N_5581,N_6956);
or U11575 (N_11575,N_7494,N_5574);
nand U11576 (N_11576,N_6113,N_5470);
xor U11577 (N_11577,N_5562,N_5347);
or U11578 (N_11578,N_8709,N_6339);
nor U11579 (N_11579,N_9117,N_5006);
xnor U11580 (N_11580,N_7284,N_6891);
or U11581 (N_11581,N_8891,N_6927);
and U11582 (N_11582,N_7534,N_8769);
and U11583 (N_11583,N_5063,N_8249);
xor U11584 (N_11584,N_8009,N_9232);
and U11585 (N_11585,N_9558,N_5273);
nand U11586 (N_11586,N_5820,N_8931);
or U11587 (N_11587,N_6366,N_6782);
xnor U11588 (N_11588,N_9002,N_7514);
nand U11589 (N_11589,N_6746,N_5458);
or U11590 (N_11590,N_9444,N_6040);
nor U11591 (N_11591,N_6224,N_8144);
nor U11592 (N_11592,N_9561,N_5734);
xnor U11593 (N_11593,N_7176,N_8715);
or U11594 (N_11594,N_8027,N_7354);
or U11595 (N_11595,N_6491,N_7398);
nor U11596 (N_11596,N_6566,N_9792);
or U11597 (N_11597,N_9585,N_9320);
nor U11598 (N_11598,N_7658,N_7007);
xor U11599 (N_11599,N_5350,N_9027);
xnor U11600 (N_11600,N_6158,N_7014);
nor U11601 (N_11601,N_5522,N_8412);
nor U11602 (N_11602,N_9106,N_9453);
nand U11603 (N_11603,N_7607,N_5873);
nand U11604 (N_11604,N_9556,N_8786);
and U11605 (N_11605,N_6859,N_8721);
xor U11606 (N_11606,N_9602,N_6307);
and U11607 (N_11607,N_6542,N_9412);
or U11608 (N_11608,N_7982,N_5378);
nand U11609 (N_11609,N_5274,N_5567);
xor U11610 (N_11610,N_8525,N_7403);
nand U11611 (N_11611,N_8515,N_7431);
and U11612 (N_11612,N_9959,N_5869);
and U11613 (N_11613,N_8118,N_9167);
or U11614 (N_11614,N_6156,N_8304);
nand U11615 (N_11615,N_7390,N_9610);
or U11616 (N_11616,N_9768,N_8644);
nand U11617 (N_11617,N_5186,N_6103);
nand U11618 (N_11618,N_6042,N_5635);
nor U11619 (N_11619,N_6044,N_6924);
and U11620 (N_11620,N_5861,N_6164);
nand U11621 (N_11621,N_9148,N_5476);
nor U11622 (N_11622,N_7953,N_8578);
xnor U11623 (N_11623,N_5317,N_7200);
and U11624 (N_11624,N_7774,N_8158);
nand U11625 (N_11625,N_6669,N_7162);
or U11626 (N_11626,N_9224,N_5545);
and U11627 (N_11627,N_6931,N_6190);
and U11628 (N_11628,N_8687,N_7770);
nand U11629 (N_11629,N_7067,N_5892);
or U11630 (N_11630,N_6122,N_8360);
xnor U11631 (N_11631,N_9908,N_9687);
and U11632 (N_11632,N_5398,N_6202);
xnor U11633 (N_11633,N_9184,N_8147);
xnor U11634 (N_11634,N_8075,N_7139);
xnor U11635 (N_11635,N_5739,N_7601);
nand U11636 (N_11636,N_9099,N_6780);
xnor U11637 (N_11637,N_9385,N_5867);
xnor U11638 (N_11638,N_6751,N_8979);
nand U11639 (N_11639,N_9621,N_6560);
nor U11640 (N_11640,N_6902,N_7215);
nor U11641 (N_11641,N_6615,N_9695);
nand U11642 (N_11642,N_8494,N_9893);
xor U11643 (N_11643,N_8745,N_9526);
nand U11644 (N_11644,N_8383,N_7063);
or U11645 (N_11645,N_5796,N_7889);
nor U11646 (N_11646,N_9869,N_6237);
or U11647 (N_11647,N_5445,N_5090);
nor U11648 (N_11648,N_8386,N_8757);
and U11649 (N_11649,N_5367,N_5327);
xnor U11650 (N_11650,N_7679,N_9421);
or U11651 (N_11651,N_9205,N_6090);
xnor U11652 (N_11652,N_6522,N_9134);
xnor U11653 (N_11653,N_9839,N_9211);
xor U11654 (N_11654,N_5579,N_6072);
or U11655 (N_11655,N_9369,N_9289);
xor U11656 (N_11656,N_6608,N_6123);
nand U11657 (N_11657,N_7039,N_9206);
nor U11658 (N_11658,N_5641,N_9782);
nand U11659 (N_11659,N_9981,N_9482);
nand U11660 (N_11660,N_9849,N_9755);
nand U11661 (N_11661,N_9770,N_5841);
nand U11662 (N_11662,N_6226,N_5446);
xnor U11663 (N_11663,N_7233,N_5964);
xor U11664 (N_11664,N_7862,N_5747);
and U11665 (N_11665,N_9177,N_8590);
and U11666 (N_11666,N_5756,N_5851);
nor U11667 (N_11667,N_6106,N_8063);
and U11668 (N_11668,N_5485,N_8589);
and U11669 (N_11669,N_9685,N_8314);
or U11670 (N_11670,N_8293,N_7825);
nor U11671 (N_11671,N_9228,N_9124);
nand U11672 (N_11672,N_6784,N_6330);
and U11673 (N_11673,N_9991,N_6809);
nor U11674 (N_11674,N_9614,N_9730);
or U11675 (N_11675,N_7314,N_7608);
or U11676 (N_11676,N_7498,N_6501);
xor U11677 (N_11677,N_8069,N_6353);
xnor U11678 (N_11678,N_9246,N_7717);
and U11679 (N_11679,N_7302,N_9176);
and U11680 (N_11680,N_9467,N_5906);
xor U11681 (N_11681,N_6016,N_8932);
xor U11682 (N_11682,N_5565,N_7585);
and U11683 (N_11683,N_7875,N_9021);
nor U11684 (N_11684,N_8505,N_9278);
and U11685 (N_11685,N_5142,N_7699);
nand U11686 (N_11686,N_7831,N_5941);
xnor U11687 (N_11687,N_5950,N_8658);
xnor U11688 (N_11688,N_6086,N_8696);
or U11689 (N_11689,N_9056,N_7541);
nand U11690 (N_11690,N_6240,N_9326);
or U11691 (N_11691,N_9799,N_9053);
xnor U11692 (N_11692,N_6674,N_9690);
nor U11693 (N_11693,N_8111,N_7246);
nor U11694 (N_11694,N_7788,N_7739);
nor U11695 (N_11695,N_8429,N_7937);
and U11696 (N_11696,N_5808,N_5764);
or U11697 (N_11697,N_8100,N_6549);
nand U11698 (N_11698,N_6089,N_7227);
xnor U11699 (N_11699,N_7994,N_6569);
nor U11700 (N_11700,N_8500,N_9163);
or U11701 (N_11701,N_5333,N_9372);
and U11702 (N_11702,N_5048,N_7224);
or U11703 (N_11703,N_8636,N_8642);
or U11704 (N_11704,N_9392,N_5968);
nand U11705 (N_11705,N_5722,N_7804);
and U11706 (N_11706,N_5128,N_6993);
xor U11707 (N_11707,N_6541,N_6318);
xnor U11708 (N_11708,N_8991,N_7423);
nor U11709 (N_11709,N_8777,N_8410);
or U11710 (N_11710,N_6602,N_7436);
xor U11711 (N_11711,N_7408,N_7028);
or U11712 (N_11712,N_8935,N_9945);
nor U11713 (N_11713,N_6527,N_8325);
nor U11714 (N_11714,N_9259,N_6370);
nand U11715 (N_11715,N_8853,N_9213);
or U11716 (N_11716,N_5996,N_6357);
and U11717 (N_11717,N_8413,N_5084);
and U11718 (N_11718,N_6711,N_7559);
or U11719 (N_11719,N_5419,N_5290);
nor U11720 (N_11720,N_5568,N_8778);
nor U11721 (N_11721,N_9250,N_5292);
nor U11722 (N_11722,N_8113,N_6394);
or U11723 (N_11723,N_8447,N_7340);
xor U11724 (N_11724,N_6070,N_8431);
and U11725 (N_11725,N_8576,N_8441);
nor U11726 (N_11726,N_8649,N_8632);
nor U11727 (N_11727,N_5362,N_8601);
and U11728 (N_11728,N_6936,N_5864);
nor U11729 (N_11729,N_8062,N_9045);
nand U11730 (N_11730,N_9985,N_8000);
nor U11731 (N_11731,N_8937,N_5752);
nand U11732 (N_11732,N_8292,N_6188);
and U11733 (N_11733,N_6595,N_5163);
nand U11734 (N_11734,N_6651,N_9248);
or U11735 (N_11735,N_6140,N_7095);
and U11736 (N_11736,N_8245,N_6976);
or U11737 (N_11737,N_6998,N_5822);
nor U11738 (N_11738,N_7777,N_8738);
or U11739 (N_11739,N_6564,N_9318);
nor U11740 (N_11740,N_9374,N_7160);
or U11741 (N_11741,N_8181,N_9503);
and U11742 (N_11742,N_5467,N_5534);
nor U11743 (N_11743,N_7504,N_8238);
or U11744 (N_11744,N_9298,N_8028);
nand U11745 (N_11745,N_9047,N_5672);
and U11746 (N_11746,N_9121,N_8117);
or U11747 (N_11747,N_7659,N_5552);
nor U11748 (N_11748,N_7773,N_9275);
nor U11749 (N_11749,N_5717,N_8328);
or U11750 (N_11750,N_5967,N_8641);
and U11751 (N_11751,N_9676,N_8998);
nor U11752 (N_11752,N_9214,N_9720);
nor U11753 (N_11753,N_6314,N_5566);
nor U11754 (N_11754,N_7478,N_9542);
nor U11755 (N_11755,N_8266,N_8968);
xor U11756 (N_11756,N_7290,N_6335);
nand U11757 (N_11757,N_8802,N_6650);
or U11758 (N_11758,N_9864,N_8224);
xor U11759 (N_11759,N_6731,N_8584);
nand U11760 (N_11760,N_8580,N_6892);
xor U11761 (N_11761,N_6354,N_9440);
or U11762 (N_11762,N_7588,N_8862);
nand U11763 (N_11763,N_8660,N_8760);
or U11764 (N_11764,N_9153,N_6910);
xnor U11765 (N_11765,N_7503,N_8373);
nand U11766 (N_11766,N_8878,N_8752);
and U11767 (N_11767,N_5674,N_5682);
xnor U11768 (N_11768,N_7766,N_6101);
nand U11769 (N_11769,N_8842,N_6306);
or U11770 (N_11770,N_7240,N_9956);
nand U11771 (N_11771,N_8462,N_9152);
nor U11772 (N_11772,N_7754,N_8322);
xor U11773 (N_11773,N_6375,N_8468);
nand U11774 (N_11774,N_9907,N_7384);
nor U11775 (N_11775,N_5649,N_5788);
and U11776 (N_11776,N_7177,N_5482);
nand U11777 (N_11777,N_5437,N_7294);
nand U11778 (N_11778,N_5957,N_9511);
nand U11779 (N_11779,N_7328,N_9380);
or U11780 (N_11780,N_6948,N_6653);
and U11781 (N_11781,N_6287,N_8868);
nand U11782 (N_11782,N_6176,N_9432);
nand U11783 (N_11783,N_6402,N_7244);
or U11784 (N_11784,N_8276,N_9287);
xnor U11785 (N_11785,N_8262,N_8952);
nor U11786 (N_11786,N_6986,N_8662);
or U11787 (N_11787,N_7700,N_7057);
xor U11788 (N_11788,N_8858,N_6777);
and U11789 (N_11789,N_6470,N_7839);
and U11790 (N_11790,N_6170,N_9980);
xnor U11791 (N_11791,N_5760,N_9533);
or U11792 (N_11792,N_8969,N_5393);
nand U11793 (N_11793,N_6797,N_5345);
nand U11794 (N_11794,N_9068,N_9029);
or U11795 (N_11795,N_5765,N_5613);
nand U11796 (N_11796,N_7473,N_6409);
or U11797 (N_11797,N_7919,N_6708);
or U11798 (N_11798,N_8313,N_9583);
and U11799 (N_11799,N_8720,N_7780);
nand U11800 (N_11800,N_9403,N_8805);
nand U11801 (N_11801,N_6185,N_5107);
nand U11802 (N_11802,N_9970,N_5266);
and U11803 (N_11803,N_7978,N_5450);
xor U11804 (N_11804,N_6403,N_9586);
or U11805 (N_11805,N_5320,N_6609);
nor U11806 (N_11806,N_7852,N_5716);
or U11807 (N_11807,N_6458,N_8861);
nand U11808 (N_11808,N_5997,N_8597);
and U11809 (N_11809,N_8239,N_8659);
and U11810 (N_11810,N_7709,N_9787);
xor U11811 (N_11811,N_7268,N_7167);
or U11812 (N_11812,N_9647,N_9615);
and U11813 (N_11813,N_7905,N_5601);
or U11814 (N_11814,N_5364,N_7285);
nand U11815 (N_11815,N_8055,N_7911);
xnor U11816 (N_11816,N_6116,N_6747);
nand U11817 (N_11817,N_5842,N_9242);
or U11818 (N_11818,N_9081,N_8185);
and U11819 (N_11819,N_9309,N_7870);
xor U11820 (N_11820,N_7850,N_7059);
or U11821 (N_11821,N_8340,N_9105);
xor U11822 (N_11822,N_7556,N_7550);
nand U11823 (N_11823,N_8946,N_5248);
nand U11824 (N_11824,N_7344,N_7800);
nand U11825 (N_11825,N_8947,N_8134);
xnor U11826 (N_11826,N_8951,N_9756);
xor U11827 (N_11827,N_5183,N_7892);
nor U11828 (N_11828,N_8007,N_6284);
nand U11829 (N_11829,N_7970,N_8405);
and U11830 (N_11830,N_8976,N_5690);
or U11831 (N_11831,N_7472,N_9788);
or U11832 (N_11832,N_8854,N_8782);
and U11833 (N_11833,N_9658,N_8013);
nand U11834 (N_11834,N_5065,N_6387);
or U11835 (N_11835,N_5032,N_8825);
or U11836 (N_11836,N_7861,N_5423);
nor U11837 (N_11837,N_7508,N_5020);
xor U11838 (N_11838,N_5543,N_6012);
or U11839 (N_11839,N_7625,N_9394);
and U11840 (N_11840,N_5776,N_7434);
and U11841 (N_11841,N_5443,N_8908);
nor U11842 (N_11842,N_7335,N_8057);
xnor U11843 (N_11843,N_8699,N_6940);
or U11844 (N_11844,N_9135,N_5270);
xnor U11845 (N_11845,N_7755,N_7180);
nor U11846 (N_11846,N_9613,N_8281);
or U11847 (N_11847,N_5891,N_6904);
nor U11848 (N_11848,N_6978,N_6953);
xor U11849 (N_11849,N_9217,N_7614);
nor U11850 (N_11850,N_9665,N_9178);
and U11851 (N_11851,N_9644,N_8015);
xnor U11852 (N_11852,N_9331,N_8392);
xnor U11853 (N_11853,N_8530,N_6909);
xor U11854 (N_11854,N_9974,N_6096);
nor U11855 (N_11855,N_9267,N_8683);
xnor U11856 (N_11856,N_5129,N_7542);
xnor U11857 (N_11857,N_9537,N_8885);
and U11858 (N_11858,N_5109,N_7303);
xnor U11859 (N_11859,N_5976,N_6194);
or U11860 (N_11860,N_9031,N_8749);
xnor U11861 (N_11861,N_5194,N_6444);
or U11862 (N_11862,N_6179,N_9963);
nand U11863 (N_11863,N_9208,N_9233);
or U11864 (N_11864,N_5316,N_7855);
and U11865 (N_11865,N_8277,N_7179);
and U11866 (N_11866,N_8887,N_7365);
nand U11867 (N_11867,N_9646,N_9976);
or U11868 (N_11868,N_6193,N_7909);
nand U11869 (N_11869,N_5277,N_5657);
or U11870 (N_11870,N_7413,N_6946);
xnor U11871 (N_11871,N_5394,N_5786);
xor U11872 (N_11872,N_9125,N_6026);
nand U11873 (N_11873,N_5076,N_9220);
nand U11874 (N_11874,N_9667,N_5098);
xor U11875 (N_11875,N_9554,N_9899);
nand U11876 (N_11876,N_5337,N_7938);
xnor U11877 (N_11877,N_8884,N_5513);
nor U11878 (N_11878,N_7144,N_7086);
or U11879 (N_11879,N_6195,N_9200);
and U11880 (N_11880,N_8093,N_5001);
xnor U11881 (N_11881,N_7217,N_9216);
xor U11882 (N_11882,N_9584,N_5389);
and U11883 (N_11883,N_8081,N_6414);
nand U11884 (N_11884,N_8704,N_8327);
and U11885 (N_11885,N_9476,N_8220);
or U11886 (N_11886,N_7359,N_5079);
xor U11887 (N_11887,N_7052,N_8785);
or U11888 (N_11888,N_5182,N_7271);
or U11889 (N_11889,N_6752,N_5193);
nor U11890 (N_11890,N_6741,N_9103);
nand U11891 (N_11891,N_9139,N_6177);
or U11892 (N_11892,N_7094,N_8452);
and U11893 (N_11893,N_6716,N_7651);
xnor U11894 (N_11894,N_6217,N_9039);
or U11895 (N_11895,N_9093,N_5410);
and U11896 (N_11896,N_7675,N_9588);
and U11897 (N_11897,N_9735,N_8192);
and U11898 (N_11898,N_6216,N_8523);
nor U11899 (N_11899,N_5173,N_5553);
nand U11900 (N_11900,N_9373,N_6877);
xor U11901 (N_11901,N_5723,N_5678);
and U11902 (N_11902,N_5731,N_9812);
and U11903 (N_11903,N_5602,N_8934);
and U11904 (N_11904,N_9390,N_5698);
xnor U11905 (N_11905,N_9410,N_9510);
and U11906 (N_11906,N_5956,N_9114);
and U11907 (N_11907,N_6750,N_7449);
and U11908 (N_11908,N_6568,N_7055);
xnor U11909 (N_11909,N_5311,N_9550);
nor U11910 (N_11910,N_7299,N_9922);
and U11911 (N_11911,N_5353,N_5374);
xor U11912 (N_11912,N_7009,N_5191);
or U11913 (N_11913,N_9666,N_8756);
nor U11914 (N_11914,N_8555,N_6468);
xor U11915 (N_11915,N_9518,N_9071);
or U11916 (N_11916,N_9096,N_7401);
or U11917 (N_11917,N_6437,N_5934);
nor U11918 (N_11918,N_7949,N_8693);
or U11919 (N_11919,N_9238,N_6227);
nor U11920 (N_11920,N_9123,N_5881);
nor U11921 (N_11921,N_8542,N_7190);
nor U11922 (N_11922,N_8187,N_8547);
and U11923 (N_11923,N_7315,N_8104);
nor U11924 (N_11924,N_8859,N_8189);
and U11925 (N_11925,N_6785,N_5507);
or U11926 (N_11926,N_7481,N_9577);
or U11927 (N_11927,N_6880,N_8822);
xnor U11928 (N_11928,N_6493,N_8345);
or U11929 (N_11929,N_5302,N_5548);
and U11930 (N_11930,N_5361,N_8563);
nand U11931 (N_11931,N_5611,N_6219);
nor U11932 (N_11932,N_9062,N_9723);
xor U11933 (N_11933,N_9531,N_6211);
xor U11934 (N_11934,N_8823,N_8234);
and U11935 (N_11935,N_9750,N_5210);
or U11936 (N_11936,N_6951,N_5938);
and U11937 (N_11937,N_8753,N_6274);
nor U11938 (N_11938,N_8036,N_7832);
nor U11939 (N_11939,N_6035,N_6390);
or U11940 (N_11940,N_5111,N_9831);
and U11941 (N_11941,N_6833,N_9140);
nor U11942 (N_11942,N_9269,N_9966);
nor U11943 (N_11943,N_9055,N_6939);
nand U11944 (N_11944,N_9243,N_6074);
xnor U11945 (N_11945,N_5952,N_6144);
nor U11946 (N_11946,N_5770,N_9165);
and U11947 (N_11947,N_8617,N_5637);
and U11948 (N_11948,N_7081,N_8684);
nor U11949 (N_11949,N_9423,N_9143);
nor U11950 (N_11950,N_8315,N_6169);
nand U11951 (N_11951,N_5572,N_6487);
nor U11952 (N_11952,N_8203,N_9600);
nand U11953 (N_11953,N_8010,N_9409);
or U11954 (N_11954,N_7298,N_9797);
xor U11955 (N_11955,N_8905,N_9992);
nand U11956 (N_11956,N_7382,N_5525);
or U11957 (N_11957,N_8913,N_6667);
or U11958 (N_11958,N_6532,N_6995);
xor U11959 (N_11959,N_6696,N_9509);
nand U11960 (N_11960,N_9239,N_9343);
xnor U11961 (N_11961,N_6624,N_9968);
nand U11962 (N_11962,N_8397,N_9046);
or U11963 (N_11963,N_8053,N_5632);
or U11964 (N_11964,N_7230,N_9194);
xnor U11965 (N_11965,N_7193,N_8674);
nor U11966 (N_11966,N_6510,N_9761);
nor U11967 (N_11967,N_7185,N_5150);
xnor U11968 (N_11968,N_6472,N_8393);
or U11969 (N_11969,N_7417,N_9300);
nor U11970 (N_11970,N_9633,N_5254);
and U11971 (N_11971,N_8286,N_8941);
or U11972 (N_11972,N_7822,N_8489);
xor U11973 (N_11973,N_9802,N_5609);
nor U11974 (N_11974,N_6066,N_7821);
xor U11975 (N_11975,N_8545,N_6573);
xor U11976 (N_11976,N_7902,N_5879);
nor U11977 (N_11977,N_8807,N_9612);
and U11978 (N_11978,N_9631,N_5083);
nand U11979 (N_11979,N_8198,N_9187);
nor U11980 (N_11980,N_8067,N_7544);
nor U11981 (N_11981,N_7790,N_6753);
nor U11982 (N_11982,N_8666,N_5658);
nand U11983 (N_11983,N_5249,N_7416);
xor U11984 (N_11984,N_7801,N_8209);
or U11985 (N_11985,N_5644,N_6990);
or U11986 (N_11986,N_9158,N_8177);
xnor U11987 (N_11987,N_9463,N_8291);
nor U11988 (N_11988,N_9551,N_7694);
or U11989 (N_11989,N_6392,N_7521);
or U11990 (N_11990,N_6320,N_8378);
nand U11991 (N_11991,N_5175,N_9210);
nor U11992 (N_11992,N_5115,N_7282);
or U11993 (N_11993,N_5988,N_5664);
or U11994 (N_11994,N_9080,N_6267);
nor U11995 (N_11995,N_8407,N_5924);
nor U11996 (N_11996,N_5617,N_6883);
nand U11997 (N_11997,N_5251,N_7882);
or U11998 (N_11998,N_9592,N_8967);
nor U11999 (N_11999,N_9449,N_7961);
or U12000 (N_12000,N_7060,N_5219);
or U12001 (N_12001,N_7165,N_7722);
xor U12002 (N_12002,N_8330,N_7226);
nand U12003 (N_12003,N_6887,N_9622);
or U12004 (N_12004,N_8712,N_9464);
nor U12005 (N_12005,N_5005,N_8182);
xnor U12006 (N_12006,N_9222,N_8078);
xnor U12007 (N_12007,N_5749,N_9529);
nor U12008 (N_12008,N_8016,N_7017);
and U12009 (N_12009,N_6558,N_7410);
and U12010 (N_12010,N_7006,N_8526);
or U12011 (N_12011,N_9617,N_9428);
xor U12012 (N_12012,N_5455,N_8732);
nand U12013 (N_12013,N_9913,N_6019);
nand U12014 (N_12014,N_9108,N_5721);
xnor U12015 (N_12015,N_9973,N_9535);
or U12016 (N_12016,N_9072,N_6686);
and U12017 (N_12017,N_5863,N_7495);
nand U12018 (N_12018,N_8847,N_6584);
nand U12019 (N_12019,N_5977,N_6006);
nor U12020 (N_12020,N_8180,N_6825);
nor U12021 (N_12021,N_8175,N_5719);
or U12022 (N_12022,N_9894,N_5280);
or U12023 (N_12023,N_5469,N_6537);
nor U12024 (N_12024,N_8070,N_6520);
nand U12025 (N_12025,N_5166,N_8706);
or U12026 (N_12026,N_6915,N_9437);
xnor U12027 (N_12027,N_6847,N_5381);
nand U12028 (N_12028,N_5425,N_8596);
and U12029 (N_12029,N_5903,N_6970);
or U12030 (N_12030,N_8112,N_9842);
nand U12031 (N_12031,N_8634,N_7255);
and U12032 (N_12032,N_9361,N_8929);
or U12033 (N_12033,N_7628,N_8076);
xnor U12034 (N_12034,N_6298,N_7245);
nand U12035 (N_12035,N_8152,N_6830);
or U12036 (N_12036,N_5481,N_8619);
nand U12037 (N_12037,N_7506,N_8404);
and U12038 (N_12038,N_6162,N_5112);
or U12039 (N_12039,N_9883,N_5984);
nand U12040 (N_12040,N_7673,N_5120);
xnor U12041 (N_12041,N_8733,N_5557);
nor U12042 (N_12042,N_9523,N_5407);
xnor U12043 (N_12043,N_5923,N_8481);
nand U12044 (N_12044,N_6083,N_6683);
or U12045 (N_12045,N_6311,N_9005);
nor U12046 (N_12046,N_8755,N_5745);
nand U12047 (N_12047,N_6934,N_5433);
or U12048 (N_12048,N_6254,N_7592);
or U12049 (N_12049,N_6556,N_7360);
nand U12050 (N_12050,N_6092,N_9994);
or U12051 (N_12051,N_8965,N_6913);
nand U12052 (N_12052,N_9000,N_8764);
nand U12053 (N_12053,N_8188,N_9844);
or U12054 (N_12054,N_8349,N_9305);
xor U12055 (N_12055,N_7121,N_6459);
xor U12056 (N_12056,N_8538,N_9706);
nand U12057 (N_12057,N_8042,N_6919);
and U12058 (N_12058,N_6692,N_7604);
nor U12059 (N_12059,N_7930,N_8575);
nor U12060 (N_12060,N_6895,N_7936);
and U12061 (N_12061,N_6574,N_7197);
xnor U12062 (N_12062,N_9941,N_9230);
and U12063 (N_12063,N_7289,N_7799);
xor U12064 (N_12064,N_5365,N_7051);
or U12065 (N_12065,N_5612,N_6724);
or U12066 (N_12066,N_7907,N_7196);
and U12067 (N_12067,N_6959,N_6174);
or U12068 (N_12068,N_6429,N_5812);
nor U12069 (N_12069,N_6013,N_8043);
nand U12070 (N_12070,N_5044,N_7130);
or U12071 (N_12071,N_6873,N_7070);
or U12072 (N_12072,N_6582,N_5692);
nand U12073 (N_12073,N_5911,N_7326);
xnor U12074 (N_12074,N_8173,N_9572);
nor U12075 (N_12075,N_7448,N_6855);
nand U12076 (N_12076,N_8259,N_8829);
or U12077 (N_12077,N_5912,N_5205);
nand U12078 (N_12078,N_8587,N_6143);
nor U12079 (N_12079,N_8864,N_6719);
nor U12080 (N_12080,N_7242,N_9098);
xnor U12081 (N_12081,N_6853,N_6732);
nor U12082 (N_12082,N_6634,N_8300);
nor U12083 (N_12083,N_8388,N_7672);
nand U12084 (N_12084,N_7168,N_7079);
xor U12085 (N_12085,N_7172,N_5902);
xnor U12086 (N_12086,N_7349,N_5868);
nor U12087 (N_12087,N_6271,N_5262);
nand U12088 (N_12088,N_9003,N_7549);
nor U12089 (N_12089,N_7134,N_5358);
or U12090 (N_12090,N_7454,N_6552);
nand U12091 (N_12091,N_8799,N_7691);
xor U12092 (N_12092,N_8278,N_8796);
nand U12093 (N_12093,N_7013,N_6652);
and U12094 (N_12094,N_8945,N_8103);
nand U12095 (N_12095,N_7708,N_8856);
and U12096 (N_12096,N_9681,N_9645);
nor U12097 (N_12097,N_9448,N_7367);
and U12098 (N_12098,N_5656,N_7137);
nor U12099 (N_12099,N_9858,N_7123);
nand U12100 (N_12100,N_8725,N_8646);
nand U12101 (N_12101,N_8421,N_8460);
xor U12102 (N_12102,N_6463,N_9696);
nor U12103 (N_12103,N_5053,N_8265);
xnor U12104 (N_12104,N_5162,N_9489);
nand U12105 (N_12105,N_8513,N_7012);
xor U12106 (N_12106,N_7747,N_5991);
or U12107 (N_12107,N_6726,N_5971);
and U12108 (N_12108,N_8168,N_7452);
nand U12109 (N_12109,N_8471,N_9459);
nand U12110 (N_12110,N_8476,N_5235);
nor U12111 (N_12111,N_5288,N_5920);
or U12112 (N_12112,N_8566,N_5075);
or U12113 (N_12113,N_6502,N_7769);
and U12114 (N_12114,N_7934,N_6112);
xnor U12115 (N_12115,N_6001,N_9548);
nand U12116 (N_12116,N_9225,N_6580);
or U12117 (N_12117,N_7511,N_7388);
xor U12118 (N_12118,N_5106,N_6391);
nand U12119 (N_12119,N_8541,N_7484);
nor U12120 (N_12120,N_6105,N_6994);
or U12121 (N_12121,N_6150,N_9496);
nand U12122 (N_12122,N_5797,N_7989);
and U12123 (N_12123,N_6469,N_7331);
xnor U12124 (N_12124,N_7064,N_6009);
or U12125 (N_12125,N_8066,N_7171);
nand U12126 (N_12126,N_9404,N_7518);
or U12127 (N_12127,N_8430,N_8355);
and U12128 (N_12128,N_9435,N_6718);
and U12129 (N_12129,N_8132,N_6097);
nor U12130 (N_12130,N_7345,N_5148);
nand U12131 (N_12131,N_9786,N_5092);
nand U12132 (N_12132,N_9618,N_7091);
and U12133 (N_12133,N_8342,N_8163);
nor U12134 (N_12134,N_6770,N_8496);
nor U12135 (N_12135,N_6758,N_5793);
and U12136 (N_12136,N_6312,N_8395);
nor U12137 (N_12137,N_9591,N_9562);
nor U12138 (N_12138,N_5640,N_5909);
nor U12139 (N_12139,N_7918,N_9758);
or U12140 (N_12140,N_5825,N_8299);
or U12141 (N_12141,N_8334,N_5782);
and U12142 (N_12142,N_6253,N_8448);
nor U12143 (N_12143,N_6071,N_5850);
and U12144 (N_12144,N_5845,N_5479);
or U12145 (N_12145,N_5152,N_9475);
nand U12146 (N_12146,N_8098,N_8176);
nor U12147 (N_12147,N_9146,N_8367);
nor U12148 (N_12148,N_5305,N_8223);
or U12149 (N_12149,N_5401,N_6856);
and U12150 (N_12150,N_7084,N_5168);
nand U12151 (N_12151,N_5276,N_5733);
nor U12152 (N_12152,N_6991,N_7308);
nor U12153 (N_12153,N_7974,N_7991);
and U12154 (N_12154,N_7274,N_8321);
nor U12155 (N_12155,N_6705,N_5686);
nand U12156 (N_12156,N_8398,N_5953);
and U12157 (N_12157,N_5781,N_5526);
nor U12158 (N_12158,N_6531,N_9862);
nor U12159 (N_12159,N_5610,N_5704);
or U12160 (N_12160,N_6973,N_7851);
or U12161 (N_12161,N_8372,N_7819);
xnor U12162 (N_12162,N_8021,N_9157);
xor U12163 (N_12163,N_9074,N_5624);
nand U12164 (N_12164,N_7827,N_6467);
and U12165 (N_12165,N_7306,N_5517);
xnor U12166 (N_12166,N_9462,N_8086);
and U12167 (N_12167,N_6911,N_8655);
or U12168 (N_12168,N_9672,N_7389);
or U12169 (N_12169,N_6322,N_7350);
nand U12170 (N_12170,N_7115,N_6695);
xnor U12171 (N_12171,N_9025,N_5918);
xnor U12172 (N_12172,N_7802,N_9189);
and U12173 (N_12173,N_5269,N_9519);
and U12174 (N_12174,N_5386,N_6796);
xor U12175 (N_12175,N_5145,N_9580);
nor U12176 (N_12176,N_5560,N_7935);
and U12177 (N_12177,N_7917,N_6952);
or U12178 (N_12178,N_5591,N_9879);
nand U12179 (N_12179,N_8323,N_8996);
or U12180 (N_12180,N_7742,N_6710);
nand U12181 (N_12181,N_5524,N_6860);
and U12182 (N_12182,N_5621,N_7046);
or U12183 (N_12183,N_6702,N_6834);
or U12184 (N_12184,N_6325,N_5310);
or U12185 (N_12185,N_7442,N_8031);
nand U12186 (N_12186,N_9052,N_7132);
or U12187 (N_12187,N_7074,N_8506);
nor U12188 (N_12188,N_9261,N_7016);
nor U12189 (N_12189,N_7204,N_8274);
or U12190 (N_12190,N_5246,N_9727);
or U12191 (N_12191,N_7096,N_6296);
or U12192 (N_12192,N_5209,N_7313);
and U12193 (N_12193,N_7061,N_6241);
or U12194 (N_12194,N_6365,N_8119);
nor U12195 (N_12195,N_8520,N_6153);
nor U12196 (N_12196,N_9368,N_8519);
or U12197 (N_12197,N_7526,N_6081);
xor U12198 (N_12198,N_8556,N_9241);
and U12199 (N_12199,N_7954,N_6908);
nor U12200 (N_12200,N_8628,N_5279);
xor U12201 (N_12201,N_8339,N_9362);
nand U12202 (N_12202,N_6038,N_8143);
nand U12203 (N_12203,N_7865,N_8422);
and U12204 (N_12204,N_5229,N_9903);
nor U12205 (N_12205,N_5008,N_6147);
nand U12206 (N_12206,N_6982,N_7243);
nand U12207 (N_12207,N_7467,N_9486);
or U12208 (N_12208,N_9169,N_8569);
nand U12209 (N_12209,N_9870,N_7251);
nand U12210 (N_12210,N_8877,N_6603);
nand U12211 (N_12211,N_5100,N_9878);
nor U12212 (N_12212,N_8491,N_7102);
xnor U12213 (N_12213,N_5405,N_7296);
xnor U12214 (N_12214,N_9273,N_5899);
nand U12215 (N_12215,N_5155,N_6637);
nand U12216 (N_12216,N_7596,N_6728);
xnor U12217 (N_12217,N_5547,N_5589);
or U12218 (N_12218,N_6642,N_7015);
nand U12219 (N_12219,N_9270,N_5003);
nand U12220 (N_12220,N_9643,N_6665);
or U12221 (N_12221,N_8179,N_5913);
and U12222 (N_12222,N_6290,N_9040);
xnor U12223 (N_12223,N_5430,N_5753);
or U12224 (N_12224,N_8625,N_8835);
xor U12225 (N_12225,N_9785,N_5848);
xnor U12226 (N_12226,N_6679,N_7283);
and U12227 (N_12227,N_9884,N_7910);
nor U12228 (N_12228,N_8390,N_9866);
and U12229 (N_12229,N_7239,N_9630);
xnor U12230 (N_12230,N_6567,N_9087);
and U12231 (N_12231,N_7552,N_6286);
nor U12232 (N_12232,N_8798,N_8916);
nor U12233 (N_12233,N_6270,N_6688);
nand U12234 (N_12234,N_5070,N_6430);
or U12235 (N_12235,N_6376,N_9417);
xor U12236 (N_12236,N_5359,N_6055);
xnor U12237 (N_12237,N_6462,N_6863);
or U12238 (N_12238,N_9898,N_6450);
nand U12239 (N_12239,N_6571,N_8083);
and U12240 (N_12240,N_9254,N_8376);
xor U12241 (N_12241,N_9408,N_7069);
or U12242 (N_12242,N_9711,N_6801);
and U12243 (N_12243,N_5014,N_8219);
xnor U12244 (N_12244,N_9603,N_5925);
xnor U12245 (N_12245,N_8726,N_7528);
xnor U12246 (N_12246,N_6638,N_8593);
xnor U12247 (N_12247,N_7848,N_7553);
nor U12248 (N_12248,N_7402,N_6136);
nand U12249 (N_12249,N_6076,N_9517);
or U12250 (N_12250,N_8529,N_8474);
and U12251 (N_12251,N_8351,N_9865);
and U12252 (N_12252,N_7145,N_5577);
or U12253 (N_12253,N_6085,N_8610);
and U12254 (N_12254,N_8294,N_5480);
xor U12255 (N_12255,N_5064,N_5798);
and U12256 (N_12256,N_6706,N_9083);
and U12257 (N_12257,N_6820,N_6917);
xnor U12258 (N_12258,N_7896,N_7222);
nor U12259 (N_12259,N_5804,N_6037);
xor U12260 (N_12260,N_8308,N_9132);
or U12261 (N_12261,N_5329,N_5963);
or U12262 (N_12262,N_8032,N_5935);
and U12263 (N_12263,N_6420,N_9845);
nor U12264 (N_12264,N_5564,N_5104);
nor U12265 (N_12265,N_5687,N_9544);
or U12266 (N_12266,N_5018,N_5660);
and U12267 (N_12267,N_8140,N_8844);
or U12268 (N_12268,N_7924,N_6827);
nor U12269 (N_12269,N_6757,N_9035);
and U12270 (N_12270,N_8255,N_5905);
xor U12271 (N_12271,N_5232,N_5943);
xor U12272 (N_12272,N_5947,N_8498);
or U12273 (N_12273,N_6999,N_5059);
nor U12274 (N_12274,N_9567,N_7963);
xor U12275 (N_12275,N_8577,N_8954);
xnor U12276 (N_12276,N_5831,N_6061);
or U12277 (N_12277,N_9946,N_7223);
and U12278 (N_12278,N_7587,N_6305);
or U12279 (N_12279,N_9714,N_8766);
nand U12280 (N_12280,N_7613,N_6543);
xor U12281 (N_12281,N_5157,N_6935);
or U12282 (N_12282,N_8212,N_9492);
nand U12283 (N_12283,N_5281,N_5504);
and U12284 (N_12284,N_5738,N_8635);
or U12285 (N_12285,N_9520,N_7505);
nor U12286 (N_12286,N_7730,N_5930);
and U12287 (N_12287,N_6499,N_7327);
nand U12288 (N_12288,N_8306,N_7001);
nor U12289 (N_12289,N_7869,N_5582);
xor U12290 (N_12290,N_6057,N_7078);
and U12291 (N_12291,N_7525,N_9713);
and U12292 (N_12292,N_7034,N_7366);
nand U12293 (N_12293,N_6802,N_6712);
and U12294 (N_12294,N_7701,N_8716);
xnor U12295 (N_12295,N_9789,N_9933);
and U12296 (N_12296,N_9386,N_8561);
nand U12297 (N_12297,N_9988,N_8902);
nor U12298 (N_12298,N_9522,N_6196);
and U12299 (N_12299,N_7779,N_7235);
or U12300 (N_12300,N_6457,N_8643);
or U12301 (N_12301,N_5297,N_8479);
nand U12302 (N_12302,N_8269,N_9060);
or U12303 (N_12303,N_9336,N_6535);
or U12304 (N_12304,N_8831,N_8914);
and U12305 (N_12305,N_7996,N_6047);
nand U12306 (N_12306,N_6151,N_8588);
xnor U12307 (N_12307,N_5857,N_9597);
and U12308 (N_12308,N_5030,N_6721);
nor U12309 (N_12309,N_5949,N_9418);
xor U12310 (N_12310,N_8973,N_7784);
nand U12311 (N_12311,N_6921,N_5373);
nand U12312 (N_12312,N_8402,N_9483);
and U12313 (N_12313,N_6442,N_8845);
and U12314 (N_12314,N_7112,N_7161);
nand U12315 (N_12315,N_6249,N_7347);
xor U12316 (N_12316,N_5247,N_9190);
nand U12317 (N_12317,N_6213,N_9816);
nand U12318 (N_12318,N_5983,N_6321);
or U12319 (N_12319,N_7232,N_6965);
nand U12320 (N_12320,N_9323,N_7030);
and U12321 (N_12321,N_8818,N_8874);
and U12322 (N_12322,N_8950,N_6452);
and U12323 (N_12323,N_7407,N_7876);
nand U12324 (N_12324,N_7630,N_9111);
nand U12325 (N_12325,N_8195,N_5052);
nand U12326 (N_12326,N_9965,N_5357);
and U12327 (N_12327,N_6583,N_9686);
or U12328 (N_12328,N_8599,N_7149);
xnor U12329 (N_12329,N_7317,N_9515);
or U12330 (N_12330,N_7270,N_9835);
or U12331 (N_12331,N_6049,N_5559);
nand U12332 (N_12332,N_8540,N_8024);
nand U12333 (N_12333,N_9179,N_5673);
xnor U12334 (N_12334,N_7783,N_6985);
xnor U12335 (N_12335,N_6607,N_6709);
and U12336 (N_12336,N_9450,N_6167);
or U12337 (N_12337,N_8990,N_8869);
and U12338 (N_12338,N_7537,N_5250);
nand U12339 (N_12339,N_8657,N_5306);
or U12340 (N_12340,N_6380,N_6616);
and U12341 (N_12341,N_9191,N_7192);
xnor U12342 (N_12342,N_9896,N_7589);
xor U12343 (N_12343,N_7796,N_8303);
or U12344 (N_12344,N_7527,N_7447);
nand U12345 (N_12345,N_8236,N_9286);
nand U12346 (N_12346,N_6054,N_7753);
or U12347 (N_12347,N_9325,N_5630);
nand U12348 (N_12348,N_9013,N_6554);
xor U12349 (N_12349,N_8639,N_5775);
nor U12350 (N_12350,N_8731,N_9650);
nor U12351 (N_12351,N_7170,N_8694);
nand U12352 (N_12352,N_9680,N_9546);
xnor U12353 (N_12353,N_6941,N_7249);
or U12354 (N_12354,N_9920,N_9204);
nand U12355 (N_12355,N_9012,N_7219);
and U12356 (N_12356,N_6506,N_9773);
nand U12357 (N_12357,N_6235,N_9085);
nor U12358 (N_12358,N_7835,N_6288);
nor U12359 (N_12359,N_6523,N_8084);
and U12360 (N_12360,N_9283,N_7731);
xor U12361 (N_12361,N_5081,N_9260);
and U12362 (N_12362,N_5859,N_8711);
nor U12363 (N_12363,N_7857,N_9652);
and U12364 (N_12364,N_9656,N_9324);
nor U12365 (N_12365,N_5461,N_9726);
and U12366 (N_12366,N_6326,N_9291);
nor U12367 (N_12367,N_8510,N_5707);
xnor U12368 (N_12368,N_9607,N_6439);
nand U12369 (N_12369,N_7003,N_5167);
or U12370 (N_12370,N_5412,N_8095);
xor U12371 (N_12371,N_9819,N_9848);
and U12372 (N_12372,N_8817,N_8461);
or U12373 (N_12373,N_9120,N_8252);
and U12374 (N_12374,N_9999,N_5858);
and U12375 (N_12375,N_8837,N_7118);
or U12376 (N_12376,N_5886,N_9001);
nor U12377 (N_12377,N_8889,N_7456);
nor U12378 (N_12378,N_7702,N_5669);
nand U12379 (N_12379,N_5855,N_5679);
or U12380 (N_12380,N_7432,N_9240);
or U12381 (N_12381,N_8751,N_9888);
xnor U12382 (N_12382,N_7356,N_5396);
or U12383 (N_12383,N_9151,N_6360);
and U12384 (N_12384,N_6093,N_5103);
xor U12385 (N_12385,N_8362,N_6034);
nor U12386 (N_12386,N_6303,N_5714);
nand U12387 (N_12387,N_6789,N_7976);
and U12388 (N_12388,N_5942,N_6377);
nand U12389 (N_12389,N_5662,N_6610);
nor U12390 (N_12390,N_6381,N_5204);
nand U12391 (N_12391,N_7426,N_6428);
or U12392 (N_12392,N_5779,N_7599);
nand U12393 (N_12393,N_6647,N_9219);
xor U12394 (N_12394,N_8640,N_9499);
nand U12395 (N_12395,N_6260,N_7990);
xnor U12396 (N_12396,N_5197,N_8270);
nand U12397 (N_12397,N_5172,N_6221);
nor U12398 (N_12398,N_6145,N_7893);
or U12399 (N_12399,N_5608,N_9032);
nand U12400 (N_12400,N_7469,N_6455);
nor U12401 (N_12401,N_6471,N_6316);
and U12402 (N_12402,N_5748,N_8309);
nor U12403 (N_12403,N_6232,N_9236);
nor U12404 (N_12404,N_5654,N_8370);
xnor U12405 (N_12405,N_8428,N_9628);
or U12406 (N_12406,N_7377,N_5342);
and U12407 (N_12407,N_9635,N_7807);
or U12408 (N_12408,N_9745,N_7712);
nand U12409 (N_12409,N_5489,N_7406);
and U12410 (N_12410,N_5146,N_7703);
xnor U12411 (N_12411,N_6755,N_7868);
or U12412 (N_12412,N_5665,N_6838);
or U12413 (N_12413,N_5432,N_8559);
nor U12414 (N_12414,N_7686,N_9749);
or U12415 (N_12415,N_8289,N_9307);
nor U12416 (N_12416,N_8573,N_7696);
xor U12417 (N_12417,N_7574,N_6587);
and U12418 (N_12418,N_8126,N_8670);
or U12419 (N_12419,N_6222,N_6415);
or U12420 (N_12420,N_7324,N_9196);
xor U12421 (N_12421,N_8680,N_8492);
xor U12422 (N_12422,N_8793,N_9506);
nor U12423 (N_12423,N_5464,N_6131);
nor U12424 (N_12424,N_5618,N_8875);
nand U12425 (N_12425,N_7159,N_5872);
and U12426 (N_12426,N_7724,N_5626);
nand U12427 (N_12427,N_8920,N_9897);
or U12428 (N_12428,N_8045,N_6737);
and U12429 (N_12429,N_9626,N_6010);
and U12430 (N_12430,N_6648,N_7885);
xor U12431 (N_12431,N_5045,N_8572);
nor U12432 (N_12432,N_5403,N_5743);
nor U12433 (N_12433,N_8815,N_9389);
xor U12434 (N_12434,N_7815,N_5550);
nor U12435 (N_12435,N_6808,N_7111);
or U12436 (N_12436,N_5072,N_7082);
nor U12437 (N_12437,N_5506,N_7029);
nand U12438 (N_12438,N_7369,N_7660);
nor U12439 (N_12439,N_5413,N_6697);
and U12440 (N_12440,N_9996,N_5463);
and U12441 (N_12441,N_6171,N_5809);
nand U12442 (N_12442,N_9393,N_5590);
and U12443 (N_12443,N_9089,N_8184);
and U12444 (N_12444,N_7721,N_9573);
and U12445 (N_12445,N_9868,N_8824);
and U12446 (N_12446,N_5927,N_9698);
nand U12447 (N_12447,N_6988,N_9502);
nand U12448 (N_12448,N_9640,N_9932);
xnor U12449 (N_12449,N_8906,N_9605);
nor U12450 (N_12450,N_8622,N_7263);
nand U12451 (N_12451,N_8065,N_8248);
nand U12452 (N_12452,N_7208,N_9873);
nand U12453 (N_12453,N_5715,N_6498);
and U12454 (N_12454,N_5440,N_5921);
or U12455 (N_12455,N_6486,N_7466);
nand U12456 (N_12456,N_8472,N_7710);
nor U12457 (N_12457,N_6645,N_7775);
and U12458 (N_12458,N_8401,N_8121);
or U12459 (N_12459,N_5990,N_7561);
xnor U12460 (N_12460,N_8995,N_9391);
nand U12461 (N_12461,N_8166,N_7794);
nand U12462 (N_12462,N_9944,N_8915);
xnor U12463 (N_12463,N_7632,N_7617);
or U12464 (N_12464,N_6557,N_9478);
or U12465 (N_12465,N_5837,N_6500);
and U12466 (N_12466,N_6214,N_8105);
xnor U12467 (N_12467,N_5054,N_5041);
or U12468 (N_12468,N_7173,N_7582);
xnor U12469 (N_12469,N_5496,N_8988);
and U12470 (N_12470,N_8924,N_6673);
and U12471 (N_12471,N_9360,N_9109);
and U12472 (N_12472,N_6509,N_9050);
nand U12473 (N_12473,N_6879,N_9834);
nand U12474 (N_12474,N_7214,N_8595);
or U12475 (N_12475,N_8892,N_8927);
or U12476 (N_12476,N_8611,N_7727);
and U12477 (N_12477,N_6675,N_8730);
nor U12478 (N_12478,N_5099,N_5706);
nand U12479 (N_12479,N_7273,N_7272);
or U12480 (N_12480,N_6916,N_6905);
nor U12481 (N_12481,N_8833,N_8232);
xor U12482 (N_12482,N_5307,N_9198);
nand U12483 (N_12483,N_8183,N_7540);
and U12484 (N_12484,N_7464,N_8453);
and U12485 (N_12485,N_5435,N_5077);
or U12486 (N_12486,N_6427,N_9077);
xor U12487 (N_12487,N_7706,N_8154);
nor U12488 (N_12488,N_7205,N_6029);
nor U12489 (N_12489,N_8964,N_7548);
nand U12490 (N_12490,N_9892,N_6124);
xor U12491 (N_12491,N_9525,N_5422);
xor U12492 (N_12492,N_5421,N_9293);
nand U12493 (N_12493,N_6328,N_9983);
nor U12494 (N_12494,N_7181,N_9438);
or U12495 (N_12495,N_8656,N_8087);
nand U12496 (N_12496,N_9736,N_8123);
and U12497 (N_12497,N_8743,N_9406);
and U12498 (N_12498,N_7211,N_8137);
or U12499 (N_12499,N_5833,N_5287);
xnor U12500 (N_12500,N_6756,N_9872);
and U12501 (N_12501,N_9039,N_5815);
and U12502 (N_12502,N_6086,N_6560);
xnor U12503 (N_12503,N_9915,N_6086);
nor U12504 (N_12504,N_8773,N_7212);
nand U12505 (N_12505,N_6691,N_9480);
or U12506 (N_12506,N_7613,N_7256);
or U12507 (N_12507,N_5998,N_6593);
nor U12508 (N_12508,N_6980,N_6510);
nor U12509 (N_12509,N_5325,N_9498);
and U12510 (N_12510,N_9733,N_9053);
and U12511 (N_12511,N_6851,N_8214);
or U12512 (N_12512,N_7804,N_6631);
or U12513 (N_12513,N_8781,N_9466);
or U12514 (N_12514,N_8088,N_9348);
nor U12515 (N_12515,N_9566,N_9520);
xnor U12516 (N_12516,N_5832,N_6219);
nand U12517 (N_12517,N_9257,N_9785);
nand U12518 (N_12518,N_9711,N_5296);
or U12519 (N_12519,N_8036,N_9024);
and U12520 (N_12520,N_9232,N_7510);
or U12521 (N_12521,N_8366,N_7359);
nor U12522 (N_12522,N_8960,N_5201);
xnor U12523 (N_12523,N_6466,N_8227);
nor U12524 (N_12524,N_6285,N_5534);
or U12525 (N_12525,N_9458,N_6985);
and U12526 (N_12526,N_9858,N_6891);
nand U12527 (N_12527,N_7318,N_7117);
xnor U12528 (N_12528,N_7889,N_9956);
xnor U12529 (N_12529,N_6933,N_7489);
and U12530 (N_12530,N_7261,N_8437);
nor U12531 (N_12531,N_6216,N_5639);
xor U12532 (N_12532,N_5697,N_7752);
or U12533 (N_12533,N_6764,N_8325);
and U12534 (N_12534,N_5481,N_9137);
and U12535 (N_12535,N_7885,N_5587);
and U12536 (N_12536,N_5417,N_5429);
nor U12537 (N_12537,N_8974,N_5922);
nor U12538 (N_12538,N_6212,N_6318);
xor U12539 (N_12539,N_8489,N_9053);
nand U12540 (N_12540,N_8362,N_8011);
nor U12541 (N_12541,N_9060,N_7335);
xor U12542 (N_12542,N_6338,N_8522);
or U12543 (N_12543,N_8818,N_5787);
nor U12544 (N_12544,N_8902,N_5893);
nor U12545 (N_12545,N_9386,N_5438);
nand U12546 (N_12546,N_7496,N_9243);
and U12547 (N_12547,N_7136,N_8319);
and U12548 (N_12548,N_6822,N_5253);
nor U12549 (N_12549,N_5125,N_5940);
or U12550 (N_12550,N_9680,N_6164);
and U12551 (N_12551,N_5563,N_6545);
and U12552 (N_12552,N_5486,N_6901);
xor U12553 (N_12553,N_8314,N_9504);
nand U12554 (N_12554,N_7584,N_5999);
and U12555 (N_12555,N_9715,N_7410);
nand U12556 (N_12556,N_6169,N_8146);
nand U12557 (N_12557,N_7052,N_5999);
nor U12558 (N_12558,N_5888,N_8260);
xor U12559 (N_12559,N_6588,N_5499);
xor U12560 (N_12560,N_9749,N_7211);
xor U12561 (N_12561,N_7946,N_9670);
or U12562 (N_12562,N_5058,N_7722);
nand U12563 (N_12563,N_9230,N_8156);
nand U12564 (N_12564,N_9190,N_7015);
or U12565 (N_12565,N_8376,N_5212);
nor U12566 (N_12566,N_6532,N_8904);
and U12567 (N_12567,N_6655,N_9409);
xor U12568 (N_12568,N_5507,N_6254);
nand U12569 (N_12569,N_9863,N_7803);
or U12570 (N_12570,N_9320,N_5394);
xor U12571 (N_12571,N_8887,N_5388);
xor U12572 (N_12572,N_9485,N_8805);
xnor U12573 (N_12573,N_7461,N_8788);
nor U12574 (N_12574,N_7414,N_6065);
or U12575 (N_12575,N_5165,N_5542);
xor U12576 (N_12576,N_8112,N_8372);
nand U12577 (N_12577,N_7509,N_5895);
or U12578 (N_12578,N_5580,N_6408);
and U12579 (N_12579,N_9965,N_8540);
and U12580 (N_12580,N_7859,N_5810);
xor U12581 (N_12581,N_6281,N_6902);
nor U12582 (N_12582,N_5564,N_5750);
and U12583 (N_12583,N_9479,N_8335);
xnor U12584 (N_12584,N_8667,N_9890);
xnor U12585 (N_12585,N_6778,N_6887);
or U12586 (N_12586,N_9579,N_7290);
nor U12587 (N_12587,N_7706,N_8258);
or U12588 (N_12588,N_6140,N_6283);
nor U12589 (N_12589,N_7369,N_9310);
nand U12590 (N_12590,N_8367,N_7240);
or U12591 (N_12591,N_6753,N_5937);
nor U12592 (N_12592,N_5591,N_8856);
and U12593 (N_12593,N_5340,N_6977);
nor U12594 (N_12594,N_5573,N_7271);
nand U12595 (N_12595,N_9148,N_7601);
xor U12596 (N_12596,N_7149,N_5881);
nand U12597 (N_12597,N_7013,N_8131);
or U12598 (N_12598,N_6386,N_9413);
nor U12599 (N_12599,N_7575,N_8576);
nand U12600 (N_12600,N_9203,N_7078);
and U12601 (N_12601,N_8810,N_5057);
and U12602 (N_12602,N_7072,N_7065);
or U12603 (N_12603,N_6672,N_6297);
xor U12604 (N_12604,N_5106,N_5637);
xor U12605 (N_12605,N_5472,N_5630);
and U12606 (N_12606,N_9900,N_6675);
or U12607 (N_12607,N_5486,N_6277);
nand U12608 (N_12608,N_6424,N_6247);
xnor U12609 (N_12609,N_8936,N_8034);
nand U12610 (N_12610,N_6537,N_5117);
nand U12611 (N_12611,N_9656,N_8173);
and U12612 (N_12612,N_7283,N_5500);
nor U12613 (N_12613,N_7281,N_6890);
and U12614 (N_12614,N_8898,N_9880);
nand U12615 (N_12615,N_8666,N_9215);
or U12616 (N_12616,N_8392,N_6145);
xnor U12617 (N_12617,N_9283,N_8303);
nand U12618 (N_12618,N_7383,N_8770);
nor U12619 (N_12619,N_8714,N_6961);
nand U12620 (N_12620,N_5520,N_6581);
or U12621 (N_12621,N_9477,N_6878);
nand U12622 (N_12622,N_6310,N_6236);
or U12623 (N_12623,N_7278,N_8437);
nor U12624 (N_12624,N_6327,N_7765);
and U12625 (N_12625,N_6510,N_8818);
or U12626 (N_12626,N_7679,N_9242);
xor U12627 (N_12627,N_5508,N_7707);
xor U12628 (N_12628,N_6072,N_5975);
or U12629 (N_12629,N_8877,N_5614);
nand U12630 (N_12630,N_7854,N_9536);
or U12631 (N_12631,N_9843,N_9828);
nand U12632 (N_12632,N_7262,N_7137);
and U12633 (N_12633,N_7518,N_6057);
nand U12634 (N_12634,N_7333,N_7622);
or U12635 (N_12635,N_5155,N_6104);
nand U12636 (N_12636,N_7899,N_8589);
or U12637 (N_12637,N_6435,N_5278);
nor U12638 (N_12638,N_5113,N_6064);
xor U12639 (N_12639,N_6835,N_9404);
nand U12640 (N_12640,N_9703,N_6080);
and U12641 (N_12641,N_5590,N_9322);
and U12642 (N_12642,N_9247,N_7575);
and U12643 (N_12643,N_7173,N_6738);
or U12644 (N_12644,N_6439,N_5122);
nor U12645 (N_12645,N_8989,N_8443);
nand U12646 (N_12646,N_5763,N_6325);
nor U12647 (N_12647,N_6984,N_6234);
nor U12648 (N_12648,N_7295,N_5524);
nand U12649 (N_12649,N_7092,N_8726);
or U12650 (N_12650,N_6788,N_8963);
or U12651 (N_12651,N_9195,N_7580);
nor U12652 (N_12652,N_9137,N_6176);
nor U12653 (N_12653,N_5882,N_6499);
nand U12654 (N_12654,N_9296,N_5667);
xnor U12655 (N_12655,N_9359,N_9242);
xnor U12656 (N_12656,N_8411,N_5262);
xnor U12657 (N_12657,N_9566,N_6560);
nand U12658 (N_12658,N_5506,N_9164);
xor U12659 (N_12659,N_8857,N_6689);
and U12660 (N_12660,N_7582,N_6681);
nor U12661 (N_12661,N_5519,N_7850);
or U12662 (N_12662,N_5177,N_6554);
nand U12663 (N_12663,N_9929,N_9263);
xnor U12664 (N_12664,N_8066,N_6172);
xor U12665 (N_12665,N_8779,N_6262);
or U12666 (N_12666,N_5768,N_7151);
xnor U12667 (N_12667,N_5118,N_9511);
and U12668 (N_12668,N_9211,N_7176);
nand U12669 (N_12669,N_8046,N_7040);
nand U12670 (N_12670,N_9371,N_5708);
nand U12671 (N_12671,N_5798,N_7688);
nand U12672 (N_12672,N_9093,N_6889);
nand U12673 (N_12673,N_7775,N_8446);
or U12674 (N_12674,N_6589,N_5779);
and U12675 (N_12675,N_6354,N_5394);
nand U12676 (N_12676,N_9093,N_8477);
and U12677 (N_12677,N_6387,N_8556);
nand U12678 (N_12678,N_6044,N_8201);
xnor U12679 (N_12679,N_5048,N_7955);
or U12680 (N_12680,N_5061,N_8918);
nor U12681 (N_12681,N_9348,N_7769);
nor U12682 (N_12682,N_8315,N_5105);
or U12683 (N_12683,N_6997,N_5566);
nor U12684 (N_12684,N_6583,N_9574);
nor U12685 (N_12685,N_9603,N_9102);
xnor U12686 (N_12686,N_6283,N_7602);
nand U12687 (N_12687,N_8723,N_8643);
xor U12688 (N_12688,N_9682,N_8241);
or U12689 (N_12689,N_8342,N_5584);
and U12690 (N_12690,N_7263,N_7381);
nand U12691 (N_12691,N_7470,N_8757);
or U12692 (N_12692,N_7134,N_8347);
and U12693 (N_12693,N_5564,N_5738);
or U12694 (N_12694,N_6391,N_6057);
and U12695 (N_12695,N_6596,N_7411);
nand U12696 (N_12696,N_5230,N_9509);
xor U12697 (N_12697,N_8791,N_8189);
nand U12698 (N_12698,N_9556,N_7799);
and U12699 (N_12699,N_8496,N_6393);
and U12700 (N_12700,N_6642,N_9956);
and U12701 (N_12701,N_6981,N_5654);
nand U12702 (N_12702,N_9569,N_5832);
nor U12703 (N_12703,N_9461,N_7898);
nand U12704 (N_12704,N_5314,N_5970);
nand U12705 (N_12705,N_5243,N_5770);
or U12706 (N_12706,N_9156,N_9247);
xnor U12707 (N_12707,N_9384,N_9791);
xor U12708 (N_12708,N_6358,N_9750);
xor U12709 (N_12709,N_5590,N_9088);
or U12710 (N_12710,N_6628,N_7199);
nand U12711 (N_12711,N_9112,N_5975);
and U12712 (N_12712,N_9441,N_5489);
or U12713 (N_12713,N_7109,N_7100);
or U12714 (N_12714,N_5595,N_5631);
nor U12715 (N_12715,N_5383,N_5954);
or U12716 (N_12716,N_5569,N_9806);
nand U12717 (N_12717,N_7806,N_9382);
and U12718 (N_12718,N_8606,N_8320);
and U12719 (N_12719,N_7924,N_9222);
or U12720 (N_12720,N_5088,N_7566);
or U12721 (N_12721,N_8135,N_5402);
or U12722 (N_12722,N_6670,N_7509);
and U12723 (N_12723,N_9810,N_9142);
and U12724 (N_12724,N_5762,N_5337);
or U12725 (N_12725,N_9138,N_8091);
or U12726 (N_12726,N_8036,N_6285);
and U12727 (N_12727,N_7061,N_6499);
xnor U12728 (N_12728,N_8035,N_9072);
nand U12729 (N_12729,N_8017,N_5449);
or U12730 (N_12730,N_8264,N_9454);
nor U12731 (N_12731,N_5498,N_5078);
nand U12732 (N_12732,N_6999,N_6318);
and U12733 (N_12733,N_9318,N_6778);
nand U12734 (N_12734,N_9155,N_8431);
xor U12735 (N_12735,N_6115,N_7716);
nor U12736 (N_12736,N_9847,N_9700);
and U12737 (N_12737,N_6415,N_8917);
xnor U12738 (N_12738,N_5383,N_8551);
and U12739 (N_12739,N_6966,N_9436);
nand U12740 (N_12740,N_5295,N_6076);
and U12741 (N_12741,N_8450,N_6428);
nand U12742 (N_12742,N_9170,N_7095);
nand U12743 (N_12743,N_8372,N_5954);
or U12744 (N_12744,N_8063,N_8823);
xor U12745 (N_12745,N_6807,N_7495);
or U12746 (N_12746,N_7361,N_7254);
xnor U12747 (N_12747,N_6435,N_7230);
xor U12748 (N_12748,N_9165,N_7158);
nand U12749 (N_12749,N_7155,N_9841);
nor U12750 (N_12750,N_7096,N_6757);
and U12751 (N_12751,N_5142,N_6503);
or U12752 (N_12752,N_6739,N_7082);
or U12753 (N_12753,N_7403,N_7796);
nor U12754 (N_12754,N_8386,N_5363);
and U12755 (N_12755,N_7030,N_8208);
nand U12756 (N_12756,N_9823,N_6594);
and U12757 (N_12757,N_7039,N_9353);
xnor U12758 (N_12758,N_7139,N_7560);
and U12759 (N_12759,N_6055,N_9504);
or U12760 (N_12760,N_6188,N_7228);
and U12761 (N_12761,N_9084,N_9520);
nand U12762 (N_12762,N_9545,N_6098);
nand U12763 (N_12763,N_8579,N_7355);
nor U12764 (N_12764,N_9802,N_6654);
xor U12765 (N_12765,N_5772,N_9776);
and U12766 (N_12766,N_8724,N_9582);
nand U12767 (N_12767,N_9683,N_5364);
xnor U12768 (N_12768,N_5009,N_9881);
and U12769 (N_12769,N_7906,N_7823);
or U12770 (N_12770,N_7685,N_6523);
and U12771 (N_12771,N_8890,N_8281);
xor U12772 (N_12772,N_5911,N_6321);
and U12773 (N_12773,N_9276,N_9264);
nand U12774 (N_12774,N_6055,N_9767);
and U12775 (N_12775,N_5495,N_6265);
nand U12776 (N_12776,N_5294,N_5502);
xor U12777 (N_12777,N_5066,N_9551);
nor U12778 (N_12778,N_7861,N_5339);
xnor U12779 (N_12779,N_8993,N_8717);
xnor U12780 (N_12780,N_5357,N_6729);
or U12781 (N_12781,N_5003,N_6635);
or U12782 (N_12782,N_9370,N_7227);
or U12783 (N_12783,N_9592,N_7552);
nand U12784 (N_12784,N_9024,N_6304);
or U12785 (N_12785,N_7240,N_5037);
xnor U12786 (N_12786,N_6270,N_8182);
nand U12787 (N_12787,N_9177,N_6186);
nand U12788 (N_12788,N_7560,N_8865);
and U12789 (N_12789,N_6823,N_9173);
and U12790 (N_12790,N_8969,N_6179);
nand U12791 (N_12791,N_6020,N_9174);
or U12792 (N_12792,N_5695,N_5510);
xnor U12793 (N_12793,N_7785,N_8632);
and U12794 (N_12794,N_5714,N_9580);
or U12795 (N_12795,N_7954,N_6871);
nor U12796 (N_12796,N_8372,N_9205);
xnor U12797 (N_12797,N_6629,N_5818);
and U12798 (N_12798,N_9944,N_8762);
nand U12799 (N_12799,N_7473,N_8972);
xor U12800 (N_12800,N_5669,N_7878);
or U12801 (N_12801,N_5953,N_5920);
nor U12802 (N_12802,N_8091,N_9742);
or U12803 (N_12803,N_7120,N_9852);
xnor U12804 (N_12804,N_9308,N_8744);
nor U12805 (N_12805,N_8292,N_8562);
or U12806 (N_12806,N_9834,N_8044);
xnor U12807 (N_12807,N_9880,N_5481);
nor U12808 (N_12808,N_9166,N_8800);
nor U12809 (N_12809,N_6706,N_8744);
and U12810 (N_12810,N_9018,N_5862);
xnor U12811 (N_12811,N_9581,N_8960);
xor U12812 (N_12812,N_9910,N_7862);
and U12813 (N_12813,N_7119,N_9049);
nand U12814 (N_12814,N_6895,N_5604);
nand U12815 (N_12815,N_8420,N_6453);
nor U12816 (N_12816,N_9383,N_8175);
nor U12817 (N_12817,N_7501,N_9887);
and U12818 (N_12818,N_9941,N_6843);
xor U12819 (N_12819,N_7302,N_5167);
or U12820 (N_12820,N_5003,N_7934);
and U12821 (N_12821,N_6884,N_8559);
nand U12822 (N_12822,N_5354,N_6016);
and U12823 (N_12823,N_6474,N_6437);
nor U12824 (N_12824,N_9717,N_9097);
nor U12825 (N_12825,N_9414,N_7426);
nand U12826 (N_12826,N_5267,N_6048);
nor U12827 (N_12827,N_6274,N_9578);
nor U12828 (N_12828,N_7131,N_9347);
nand U12829 (N_12829,N_5301,N_5510);
xnor U12830 (N_12830,N_8266,N_7628);
or U12831 (N_12831,N_8596,N_8605);
or U12832 (N_12832,N_7108,N_9794);
nor U12833 (N_12833,N_7883,N_5805);
nand U12834 (N_12834,N_7973,N_8200);
or U12835 (N_12835,N_7085,N_8260);
xnor U12836 (N_12836,N_7141,N_7991);
xnor U12837 (N_12837,N_6304,N_6340);
nand U12838 (N_12838,N_9408,N_5101);
nand U12839 (N_12839,N_6387,N_7799);
nor U12840 (N_12840,N_6819,N_6489);
nand U12841 (N_12841,N_5057,N_9337);
nor U12842 (N_12842,N_5901,N_9882);
and U12843 (N_12843,N_5444,N_8302);
xor U12844 (N_12844,N_8784,N_8906);
nor U12845 (N_12845,N_9684,N_5874);
and U12846 (N_12846,N_8255,N_5637);
or U12847 (N_12847,N_7283,N_5733);
or U12848 (N_12848,N_5561,N_6312);
and U12849 (N_12849,N_9390,N_9051);
or U12850 (N_12850,N_8654,N_6978);
xor U12851 (N_12851,N_7142,N_5750);
nor U12852 (N_12852,N_9027,N_6544);
nor U12853 (N_12853,N_7180,N_6020);
and U12854 (N_12854,N_6671,N_6658);
xor U12855 (N_12855,N_8752,N_8108);
or U12856 (N_12856,N_5656,N_7168);
xnor U12857 (N_12857,N_5807,N_8640);
and U12858 (N_12858,N_8630,N_7783);
xnor U12859 (N_12859,N_8444,N_7910);
or U12860 (N_12860,N_9975,N_5364);
xnor U12861 (N_12861,N_9643,N_8958);
xor U12862 (N_12862,N_9046,N_7215);
nand U12863 (N_12863,N_9937,N_5844);
or U12864 (N_12864,N_9701,N_8523);
nor U12865 (N_12865,N_8071,N_7688);
nand U12866 (N_12866,N_9616,N_5614);
nor U12867 (N_12867,N_6984,N_5556);
nor U12868 (N_12868,N_6759,N_9119);
and U12869 (N_12869,N_5332,N_8585);
nand U12870 (N_12870,N_7622,N_6491);
xor U12871 (N_12871,N_6847,N_7565);
nand U12872 (N_12872,N_9383,N_9373);
xnor U12873 (N_12873,N_6133,N_8009);
xor U12874 (N_12874,N_8410,N_7872);
nor U12875 (N_12875,N_5857,N_8994);
nor U12876 (N_12876,N_5554,N_9677);
xor U12877 (N_12877,N_5100,N_5245);
nor U12878 (N_12878,N_8879,N_7556);
nand U12879 (N_12879,N_8875,N_6341);
or U12880 (N_12880,N_6548,N_7068);
nand U12881 (N_12881,N_6084,N_5728);
and U12882 (N_12882,N_5384,N_5676);
or U12883 (N_12883,N_8262,N_7364);
nand U12884 (N_12884,N_6522,N_9007);
and U12885 (N_12885,N_7288,N_5593);
xnor U12886 (N_12886,N_5666,N_6333);
and U12887 (N_12887,N_5700,N_9230);
or U12888 (N_12888,N_6982,N_6992);
nand U12889 (N_12889,N_9538,N_9803);
or U12890 (N_12890,N_8222,N_8791);
and U12891 (N_12891,N_8748,N_9978);
or U12892 (N_12892,N_6849,N_9441);
or U12893 (N_12893,N_7301,N_7855);
and U12894 (N_12894,N_9247,N_8118);
nor U12895 (N_12895,N_9685,N_8643);
nor U12896 (N_12896,N_9831,N_8364);
or U12897 (N_12897,N_9964,N_9268);
or U12898 (N_12898,N_8126,N_9850);
xnor U12899 (N_12899,N_5272,N_9951);
nand U12900 (N_12900,N_6782,N_7877);
or U12901 (N_12901,N_6544,N_6042);
and U12902 (N_12902,N_9498,N_7478);
xnor U12903 (N_12903,N_8761,N_9301);
and U12904 (N_12904,N_9877,N_7498);
nand U12905 (N_12905,N_7999,N_6994);
xnor U12906 (N_12906,N_8099,N_8886);
and U12907 (N_12907,N_5259,N_6556);
or U12908 (N_12908,N_8351,N_8617);
nand U12909 (N_12909,N_6305,N_8443);
xor U12910 (N_12910,N_6055,N_6340);
xor U12911 (N_12911,N_6568,N_5955);
nor U12912 (N_12912,N_8317,N_5362);
nor U12913 (N_12913,N_6001,N_8324);
xor U12914 (N_12914,N_9118,N_5324);
and U12915 (N_12915,N_9085,N_8945);
nand U12916 (N_12916,N_7861,N_8986);
and U12917 (N_12917,N_6168,N_7258);
nor U12918 (N_12918,N_9252,N_5819);
nand U12919 (N_12919,N_5615,N_8499);
nor U12920 (N_12920,N_9658,N_9696);
or U12921 (N_12921,N_6703,N_6035);
or U12922 (N_12922,N_8297,N_5484);
nor U12923 (N_12923,N_7222,N_9777);
xnor U12924 (N_12924,N_5919,N_6903);
xnor U12925 (N_12925,N_8712,N_7891);
nand U12926 (N_12926,N_7567,N_9463);
nor U12927 (N_12927,N_8263,N_6700);
and U12928 (N_12928,N_6379,N_6516);
nand U12929 (N_12929,N_6105,N_9918);
nand U12930 (N_12930,N_7448,N_7712);
xor U12931 (N_12931,N_7116,N_8141);
nor U12932 (N_12932,N_8407,N_8505);
or U12933 (N_12933,N_6409,N_5125);
nor U12934 (N_12934,N_6484,N_7628);
or U12935 (N_12935,N_7151,N_7553);
xor U12936 (N_12936,N_6013,N_8882);
and U12937 (N_12937,N_9749,N_6668);
xor U12938 (N_12938,N_6739,N_8668);
or U12939 (N_12939,N_9638,N_8503);
nor U12940 (N_12940,N_8044,N_7370);
nand U12941 (N_12941,N_5040,N_5378);
xor U12942 (N_12942,N_9743,N_7980);
and U12943 (N_12943,N_6067,N_5527);
and U12944 (N_12944,N_6370,N_7023);
xor U12945 (N_12945,N_9858,N_6331);
and U12946 (N_12946,N_6304,N_7682);
nor U12947 (N_12947,N_5515,N_7669);
nor U12948 (N_12948,N_7949,N_6315);
nand U12949 (N_12949,N_5025,N_6454);
xor U12950 (N_12950,N_7055,N_6923);
or U12951 (N_12951,N_5311,N_6133);
nor U12952 (N_12952,N_9475,N_5088);
xnor U12953 (N_12953,N_5460,N_6537);
nor U12954 (N_12954,N_6216,N_7913);
xor U12955 (N_12955,N_6097,N_9711);
xnor U12956 (N_12956,N_7394,N_6288);
xor U12957 (N_12957,N_9729,N_6128);
xor U12958 (N_12958,N_8317,N_7328);
nor U12959 (N_12959,N_7626,N_6913);
nor U12960 (N_12960,N_9924,N_6997);
and U12961 (N_12961,N_6363,N_6341);
or U12962 (N_12962,N_9392,N_8107);
nand U12963 (N_12963,N_8391,N_6890);
or U12964 (N_12964,N_5050,N_8434);
xnor U12965 (N_12965,N_9183,N_8700);
and U12966 (N_12966,N_6857,N_8182);
nand U12967 (N_12967,N_7861,N_5863);
xor U12968 (N_12968,N_5866,N_8022);
or U12969 (N_12969,N_8315,N_9158);
nand U12970 (N_12970,N_5379,N_9131);
nand U12971 (N_12971,N_7791,N_5062);
nor U12972 (N_12972,N_5800,N_9282);
xor U12973 (N_12973,N_6566,N_6036);
nand U12974 (N_12974,N_5504,N_7065);
or U12975 (N_12975,N_6459,N_9442);
nor U12976 (N_12976,N_5903,N_9712);
and U12977 (N_12977,N_6715,N_8361);
nor U12978 (N_12978,N_5699,N_7191);
xnor U12979 (N_12979,N_5216,N_8199);
xnor U12980 (N_12980,N_8866,N_5283);
nor U12981 (N_12981,N_7577,N_6704);
nand U12982 (N_12982,N_6418,N_6899);
xnor U12983 (N_12983,N_6770,N_8949);
nor U12984 (N_12984,N_8803,N_5294);
xnor U12985 (N_12985,N_6517,N_9165);
or U12986 (N_12986,N_8429,N_9624);
nand U12987 (N_12987,N_7121,N_8990);
nand U12988 (N_12988,N_5576,N_8980);
or U12989 (N_12989,N_5075,N_6331);
nand U12990 (N_12990,N_8090,N_9197);
or U12991 (N_12991,N_9297,N_5483);
nor U12992 (N_12992,N_8681,N_7214);
or U12993 (N_12993,N_9798,N_7362);
xor U12994 (N_12994,N_5036,N_8702);
or U12995 (N_12995,N_7030,N_6775);
nor U12996 (N_12996,N_8743,N_9651);
nand U12997 (N_12997,N_7251,N_9725);
and U12998 (N_12998,N_7141,N_8815);
nor U12999 (N_12999,N_5239,N_9713);
xor U13000 (N_13000,N_9028,N_9842);
and U13001 (N_13001,N_9931,N_6829);
nor U13002 (N_13002,N_9321,N_8864);
nand U13003 (N_13003,N_6411,N_6533);
nand U13004 (N_13004,N_8517,N_5018);
and U13005 (N_13005,N_9357,N_6525);
nand U13006 (N_13006,N_5331,N_7829);
xor U13007 (N_13007,N_9729,N_7367);
nor U13008 (N_13008,N_7074,N_5714);
nand U13009 (N_13009,N_6404,N_5611);
or U13010 (N_13010,N_8822,N_7165);
xor U13011 (N_13011,N_8916,N_5426);
and U13012 (N_13012,N_6494,N_5107);
or U13013 (N_13013,N_5713,N_6860);
or U13014 (N_13014,N_9684,N_8914);
or U13015 (N_13015,N_6412,N_9831);
or U13016 (N_13016,N_9478,N_9523);
nor U13017 (N_13017,N_9821,N_5253);
and U13018 (N_13018,N_7749,N_5726);
or U13019 (N_13019,N_5976,N_9793);
xor U13020 (N_13020,N_8347,N_5672);
or U13021 (N_13021,N_7303,N_6222);
nand U13022 (N_13022,N_6448,N_8573);
and U13023 (N_13023,N_7477,N_6703);
or U13024 (N_13024,N_8734,N_5108);
and U13025 (N_13025,N_9295,N_6992);
xnor U13026 (N_13026,N_6332,N_7524);
xor U13027 (N_13027,N_8743,N_8885);
and U13028 (N_13028,N_9564,N_5706);
or U13029 (N_13029,N_7947,N_8529);
or U13030 (N_13030,N_9599,N_5059);
nor U13031 (N_13031,N_5844,N_7358);
and U13032 (N_13032,N_5837,N_9421);
or U13033 (N_13033,N_8277,N_5744);
and U13034 (N_13034,N_7104,N_5856);
nor U13035 (N_13035,N_5470,N_6765);
xor U13036 (N_13036,N_7246,N_8095);
nor U13037 (N_13037,N_7953,N_8282);
nand U13038 (N_13038,N_5500,N_6280);
nand U13039 (N_13039,N_8247,N_8090);
or U13040 (N_13040,N_7547,N_7282);
and U13041 (N_13041,N_9230,N_7921);
xnor U13042 (N_13042,N_6049,N_6273);
xnor U13043 (N_13043,N_6014,N_9831);
or U13044 (N_13044,N_6949,N_6556);
nor U13045 (N_13045,N_7328,N_5492);
and U13046 (N_13046,N_6631,N_6092);
or U13047 (N_13047,N_5100,N_9218);
or U13048 (N_13048,N_8989,N_7287);
nand U13049 (N_13049,N_7586,N_7665);
and U13050 (N_13050,N_5901,N_7550);
or U13051 (N_13051,N_5439,N_5098);
xor U13052 (N_13052,N_8030,N_6955);
or U13053 (N_13053,N_5769,N_8944);
nor U13054 (N_13054,N_9587,N_8125);
nor U13055 (N_13055,N_5614,N_8099);
xnor U13056 (N_13056,N_6540,N_5217);
xor U13057 (N_13057,N_9574,N_8844);
xnor U13058 (N_13058,N_7382,N_9380);
nor U13059 (N_13059,N_5244,N_5499);
and U13060 (N_13060,N_5551,N_5557);
xnor U13061 (N_13061,N_7469,N_7589);
nand U13062 (N_13062,N_7817,N_8009);
nand U13063 (N_13063,N_6186,N_5300);
nor U13064 (N_13064,N_5450,N_5956);
and U13065 (N_13065,N_6982,N_5699);
or U13066 (N_13066,N_9234,N_9862);
or U13067 (N_13067,N_8001,N_9960);
and U13068 (N_13068,N_5020,N_6157);
and U13069 (N_13069,N_5240,N_7120);
nand U13070 (N_13070,N_9939,N_6657);
and U13071 (N_13071,N_8574,N_6871);
or U13072 (N_13072,N_6725,N_5700);
or U13073 (N_13073,N_8632,N_9265);
or U13074 (N_13074,N_5161,N_7382);
and U13075 (N_13075,N_7602,N_7913);
xnor U13076 (N_13076,N_9461,N_9740);
nor U13077 (N_13077,N_5015,N_7839);
nor U13078 (N_13078,N_7882,N_8679);
or U13079 (N_13079,N_5942,N_6135);
nand U13080 (N_13080,N_5367,N_7615);
or U13081 (N_13081,N_9077,N_6402);
nand U13082 (N_13082,N_5175,N_7427);
nand U13083 (N_13083,N_9587,N_9987);
and U13084 (N_13084,N_5350,N_5016);
nand U13085 (N_13085,N_5743,N_5130);
nor U13086 (N_13086,N_6917,N_5568);
and U13087 (N_13087,N_5045,N_9504);
nor U13088 (N_13088,N_5273,N_5439);
nor U13089 (N_13089,N_5364,N_6841);
xor U13090 (N_13090,N_6650,N_5601);
nand U13091 (N_13091,N_5704,N_5973);
nand U13092 (N_13092,N_5458,N_8799);
xor U13093 (N_13093,N_9735,N_9297);
and U13094 (N_13094,N_8264,N_6107);
nand U13095 (N_13095,N_8627,N_8977);
nand U13096 (N_13096,N_6182,N_9177);
and U13097 (N_13097,N_5819,N_5206);
xor U13098 (N_13098,N_9597,N_9676);
nor U13099 (N_13099,N_8741,N_6658);
or U13100 (N_13100,N_9186,N_6350);
xnor U13101 (N_13101,N_7305,N_8946);
nand U13102 (N_13102,N_7537,N_6429);
nand U13103 (N_13103,N_5421,N_8635);
or U13104 (N_13104,N_6009,N_9346);
and U13105 (N_13105,N_5849,N_7523);
nor U13106 (N_13106,N_8404,N_5570);
nand U13107 (N_13107,N_8536,N_5189);
nand U13108 (N_13108,N_6145,N_6032);
nand U13109 (N_13109,N_7753,N_8891);
xor U13110 (N_13110,N_7356,N_6002);
and U13111 (N_13111,N_8503,N_8805);
nand U13112 (N_13112,N_5101,N_8010);
nand U13113 (N_13113,N_9382,N_8188);
nand U13114 (N_13114,N_6671,N_6984);
and U13115 (N_13115,N_9645,N_8781);
xor U13116 (N_13116,N_7966,N_9655);
nand U13117 (N_13117,N_6433,N_5764);
and U13118 (N_13118,N_9184,N_6787);
and U13119 (N_13119,N_6277,N_5271);
and U13120 (N_13120,N_8740,N_8452);
and U13121 (N_13121,N_7461,N_5398);
and U13122 (N_13122,N_6185,N_6550);
xor U13123 (N_13123,N_5699,N_6432);
nor U13124 (N_13124,N_6290,N_7697);
and U13125 (N_13125,N_7725,N_5192);
and U13126 (N_13126,N_5576,N_8032);
nor U13127 (N_13127,N_8460,N_5549);
and U13128 (N_13128,N_7384,N_5613);
or U13129 (N_13129,N_9948,N_5793);
nand U13130 (N_13130,N_7175,N_7120);
nor U13131 (N_13131,N_6801,N_6523);
xnor U13132 (N_13132,N_9393,N_5469);
nand U13133 (N_13133,N_7276,N_8797);
or U13134 (N_13134,N_8750,N_5449);
nor U13135 (N_13135,N_9649,N_6166);
nand U13136 (N_13136,N_8372,N_7647);
or U13137 (N_13137,N_8848,N_7530);
and U13138 (N_13138,N_9967,N_8481);
nand U13139 (N_13139,N_6202,N_5718);
nand U13140 (N_13140,N_9965,N_6531);
xnor U13141 (N_13141,N_8509,N_9973);
xnor U13142 (N_13142,N_7928,N_6572);
or U13143 (N_13143,N_7842,N_8224);
nand U13144 (N_13144,N_7667,N_8133);
xor U13145 (N_13145,N_5540,N_7824);
nor U13146 (N_13146,N_6566,N_8418);
and U13147 (N_13147,N_9832,N_5721);
nand U13148 (N_13148,N_5779,N_8814);
nor U13149 (N_13149,N_7723,N_9238);
and U13150 (N_13150,N_8582,N_9452);
and U13151 (N_13151,N_7334,N_7369);
nand U13152 (N_13152,N_5869,N_9367);
nand U13153 (N_13153,N_8625,N_8546);
xnor U13154 (N_13154,N_8520,N_8594);
xor U13155 (N_13155,N_7832,N_8544);
nand U13156 (N_13156,N_6074,N_9341);
nor U13157 (N_13157,N_9550,N_7246);
nor U13158 (N_13158,N_9422,N_9123);
or U13159 (N_13159,N_9803,N_5597);
nand U13160 (N_13160,N_7675,N_7078);
or U13161 (N_13161,N_5746,N_8827);
nor U13162 (N_13162,N_9832,N_8204);
and U13163 (N_13163,N_7584,N_8731);
xor U13164 (N_13164,N_7018,N_9889);
nor U13165 (N_13165,N_9936,N_9703);
or U13166 (N_13166,N_7419,N_5779);
nor U13167 (N_13167,N_8985,N_5394);
or U13168 (N_13168,N_9809,N_8001);
and U13169 (N_13169,N_7286,N_7422);
nor U13170 (N_13170,N_7593,N_8042);
nor U13171 (N_13171,N_8173,N_7943);
nor U13172 (N_13172,N_9996,N_9266);
nand U13173 (N_13173,N_7503,N_7826);
and U13174 (N_13174,N_9317,N_9757);
and U13175 (N_13175,N_9157,N_6483);
xnor U13176 (N_13176,N_9858,N_9310);
nor U13177 (N_13177,N_8944,N_9582);
nand U13178 (N_13178,N_5726,N_6663);
or U13179 (N_13179,N_9513,N_8673);
or U13180 (N_13180,N_9822,N_8280);
nand U13181 (N_13181,N_8499,N_7353);
nor U13182 (N_13182,N_7185,N_5414);
nor U13183 (N_13183,N_9598,N_5369);
nand U13184 (N_13184,N_8990,N_6308);
nor U13185 (N_13185,N_6514,N_6576);
nand U13186 (N_13186,N_9861,N_9576);
xor U13187 (N_13187,N_8502,N_8374);
nand U13188 (N_13188,N_7242,N_5296);
nand U13189 (N_13189,N_6024,N_8075);
or U13190 (N_13190,N_7697,N_8661);
nor U13191 (N_13191,N_7096,N_5561);
or U13192 (N_13192,N_6837,N_6600);
and U13193 (N_13193,N_7897,N_9152);
nor U13194 (N_13194,N_7087,N_8426);
and U13195 (N_13195,N_8616,N_7615);
and U13196 (N_13196,N_6768,N_8351);
and U13197 (N_13197,N_9533,N_5985);
xor U13198 (N_13198,N_9343,N_8468);
and U13199 (N_13199,N_7738,N_5028);
xor U13200 (N_13200,N_6379,N_6746);
xnor U13201 (N_13201,N_5481,N_7655);
and U13202 (N_13202,N_6524,N_7270);
xor U13203 (N_13203,N_7837,N_9227);
nor U13204 (N_13204,N_7744,N_9635);
nor U13205 (N_13205,N_6708,N_8515);
or U13206 (N_13206,N_7558,N_5873);
nor U13207 (N_13207,N_9726,N_8284);
nor U13208 (N_13208,N_8645,N_5453);
and U13209 (N_13209,N_5146,N_5104);
and U13210 (N_13210,N_9058,N_8602);
or U13211 (N_13211,N_7050,N_7904);
or U13212 (N_13212,N_7067,N_8515);
xnor U13213 (N_13213,N_8017,N_8140);
nand U13214 (N_13214,N_9405,N_5035);
nand U13215 (N_13215,N_7520,N_5188);
xor U13216 (N_13216,N_6436,N_6297);
nand U13217 (N_13217,N_6792,N_8637);
nor U13218 (N_13218,N_5983,N_9574);
and U13219 (N_13219,N_9772,N_9315);
xor U13220 (N_13220,N_9856,N_7818);
nand U13221 (N_13221,N_6138,N_5846);
xor U13222 (N_13222,N_6974,N_7114);
nor U13223 (N_13223,N_6307,N_8947);
nand U13224 (N_13224,N_5399,N_8891);
xnor U13225 (N_13225,N_6820,N_8328);
nand U13226 (N_13226,N_8992,N_8755);
nor U13227 (N_13227,N_5421,N_9006);
or U13228 (N_13228,N_8449,N_7971);
and U13229 (N_13229,N_7644,N_9242);
nor U13230 (N_13230,N_6908,N_8064);
nand U13231 (N_13231,N_7374,N_5053);
and U13232 (N_13232,N_7253,N_9220);
xnor U13233 (N_13233,N_6941,N_8422);
or U13234 (N_13234,N_6142,N_6456);
and U13235 (N_13235,N_5780,N_6431);
xor U13236 (N_13236,N_7624,N_8946);
or U13237 (N_13237,N_6427,N_7488);
and U13238 (N_13238,N_6049,N_6587);
xor U13239 (N_13239,N_8703,N_5368);
nor U13240 (N_13240,N_7691,N_5125);
nor U13241 (N_13241,N_9598,N_8005);
nand U13242 (N_13242,N_6184,N_9604);
nand U13243 (N_13243,N_6461,N_5400);
nand U13244 (N_13244,N_5391,N_9047);
nor U13245 (N_13245,N_6037,N_6093);
nor U13246 (N_13246,N_6853,N_9501);
nand U13247 (N_13247,N_5366,N_6545);
and U13248 (N_13248,N_8868,N_6718);
and U13249 (N_13249,N_9211,N_5438);
nand U13250 (N_13250,N_5299,N_7501);
or U13251 (N_13251,N_7678,N_8995);
nand U13252 (N_13252,N_8650,N_6252);
and U13253 (N_13253,N_9625,N_9568);
and U13254 (N_13254,N_5768,N_7181);
nand U13255 (N_13255,N_7490,N_9068);
nand U13256 (N_13256,N_6658,N_6069);
xor U13257 (N_13257,N_7043,N_6031);
nor U13258 (N_13258,N_7487,N_8473);
nor U13259 (N_13259,N_5855,N_9641);
nor U13260 (N_13260,N_7941,N_8749);
or U13261 (N_13261,N_7980,N_5581);
nor U13262 (N_13262,N_6233,N_8909);
and U13263 (N_13263,N_8924,N_9499);
or U13264 (N_13264,N_7528,N_9073);
nor U13265 (N_13265,N_7572,N_9620);
nand U13266 (N_13266,N_8416,N_7443);
nor U13267 (N_13267,N_8784,N_5611);
or U13268 (N_13268,N_6193,N_8808);
xnor U13269 (N_13269,N_8729,N_7192);
nor U13270 (N_13270,N_7458,N_6363);
or U13271 (N_13271,N_5372,N_8072);
xnor U13272 (N_13272,N_9090,N_8248);
nand U13273 (N_13273,N_8211,N_6198);
nor U13274 (N_13274,N_9290,N_5125);
and U13275 (N_13275,N_8039,N_7804);
and U13276 (N_13276,N_9065,N_6194);
or U13277 (N_13277,N_7832,N_6005);
xnor U13278 (N_13278,N_8824,N_5419);
or U13279 (N_13279,N_5873,N_7923);
or U13280 (N_13280,N_9788,N_9672);
nor U13281 (N_13281,N_9296,N_6763);
xnor U13282 (N_13282,N_9936,N_6013);
or U13283 (N_13283,N_9580,N_8370);
nor U13284 (N_13284,N_8087,N_7008);
nand U13285 (N_13285,N_5704,N_5005);
and U13286 (N_13286,N_9381,N_8507);
or U13287 (N_13287,N_7554,N_5529);
nor U13288 (N_13288,N_5430,N_8998);
nand U13289 (N_13289,N_6154,N_9240);
and U13290 (N_13290,N_5788,N_6040);
nor U13291 (N_13291,N_7689,N_8496);
nand U13292 (N_13292,N_5637,N_6386);
or U13293 (N_13293,N_5228,N_5165);
nand U13294 (N_13294,N_6018,N_9002);
and U13295 (N_13295,N_9470,N_7938);
nand U13296 (N_13296,N_9673,N_9777);
nor U13297 (N_13297,N_9101,N_8679);
nor U13298 (N_13298,N_5248,N_9659);
or U13299 (N_13299,N_7461,N_6015);
xnor U13300 (N_13300,N_7257,N_5622);
or U13301 (N_13301,N_8868,N_8000);
nor U13302 (N_13302,N_7043,N_5630);
and U13303 (N_13303,N_6309,N_8255);
nand U13304 (N_13304,N_6130,N_7267);
or U13305 (N_13305,N_7099,N_5321);
xnor U13306 (N_13306,N_6295,N_5302);
and U13307 (N_13307,N_5008,N_9778);
or U13308 (N_13308,N_7283,N_5435);
nand U13309 (N_13309,N_5006,N_6077);
nor U13310 (N_13310,N_6136,N_5636);
nor U13311 (N_13311,N_8112,N_8754);
and U13312 (N_13312,N_9527,N_7575);
nor U13313 (N_13313,N_9853,N_8569);
or U13314 (N_13314,N_5422,N_6235);
nor U13315 (N_13315,N_6726,N_6952);
and U13316 (N_13316,N_5235,N_6549);
xnor U13317 (N_13317,N_6801,N_8469);
nand U13318 (N_13318,N_5580,N_5816);
or U13319 (N_13319,N_6040,N_8680);
nor U13320 (N_13320,N_8143,N_6855);
xnor U13321 (N_13321,N_8933,N_6048);
nor U13322 (N_13322,N_6960,N_9327);
nand U13323 (N_13323,N_8173,N_8788);
nor U13324 (N_13324,N_7179,N_7652);
and U13325 (N_13325,N_8039,N_8473);
and U13326 (N_13326,N_6736,N_5269);
nor U13327 (N_13327,N_5102,N_7830);
and U13328 (N_13328,N_7776,N_9661);
xor U13329 (N_13329,N_8241,N_6916);
and U13330 (N_13330,N_5463,N_6269);
nand U13331 (N_13331,N_5428,N_5757);
and U13332 (N_13332,N_9157,N_6357);
xnor U13333 (N_13333,N_6390,N_8095);
nand U13334 (N_13334,N_8120,N_6813);
and U13335 (N_13335,N_5042,N_5013);
and U13336 (N_13336,N_6832,N_5372);
or U13337 (N_13337,N_5836,N_5077);
xnor U13338 (N_13338,N_7192,N_8340);
xnor U13339 (N_13339,N_6957,N_6136);
or U13340 (N_13340,N_8820,N_9768);
xnor U13341 (N_13341,N_8009,N_6531);
nor U13342 (N_13342,N_8003,N_5067);
and U13343 (N_13343,N_8578,N_7602);
or U13344 (N_13344,N_7729,N_6539);
or U13345 (N_13345,N_9916,N_6600);
nand U13346 (N_13346,N_5840,N_8259);
and U13347 (N_13347,N_6159,N_6223);
nor U13348 (N_13348,N_6781,N_9996);
nor U13349 (N_13349,N_5764,N_5024);
nand U13350 (N_13350,N_8103,N_7955);
and U13351 (N_13351,N_7262,N_5173);
nor U13352 (N_13352,N_9583,N_5114);
xor U13353 (N_13353,N_5334,N_7627);
and U13354 (N_13354,N_8949,N_6843);
nor U13355 (N_13355,N_9375,N_9621);
and U13356 (N_13356,N_6784,N_7581);
nor U13357 (N_13357,N_6389,N_7683);
xnor U13358 (N_13358,N_6241,N_7596);
nand U13359 (N_13359,N_9016,N_5458);
or U13360 (N_13360,N_7760,N_9929);
and U13361 (N_13361,N_5581,N_8793);
or U13362 (N_13362,N_9516,N_5204);
or U13363 (N_13363,N_6339,N_7849);
or U13364 (N_13364,N_7372,N_7367);
nand U13365 (N_13365,N_5454,N_7706);
xor U13366 (N_13366,N_8014,N_6239);
or U13367 (N_13367,N_6393,N_6594);
and U13368 (N_13368,N_6231,N_7994);
and U13369 (N_13369,N_6522,N_9147);
nand U13370 (N_13370,N_8153,N_5663);
nand U13371 (N_13371,N_8810,N_5086);
and U13372 (N_13372,N_7563,N_7654);
nor U13373 (N_13373,N_7690,N_7404);
xnor U13374 (N_13374,N_9364,N_8056);
or U13375 (N_13375,N_6221,N_7036);
and U13376 (N_13376,N_6680,N_8918);
xor U13377 (N_13377,N_8603,N_6400);
nor U13378 (N_13378,N_8342,N_6784);
xor U13379 (N_13379,N_5273,N_8220);
nor U13380 (N_13380,N_7163,N_5389);
nand U13381 (N_13381,N_7654,N_9452);
or U13382 (N_13382,N_7220,N_6458);
or U13383 (N_13383,N_7648,N_5740);
or U13384 (N_13384,N_6408,N_7054);
or U13385 (N_13385,N_6255,N_6259);
xnor U13386 (N_13386,N_8352,N_7150);
and U13387 (N_13387,N_6118,N_9913);
or U13388 (N_13388,N_5687,N_5037);
xor U13389 (N_13389,N_6112,N_5497);
nand U13390 (N_13390,N_5480,N_8582);
or U13391 (N_13391,N_7515,N_5151);
and U13392 (N_13392,N_9799,N_7169);
and U13393 (N_13393,N_6006,N_5740);
nand U13394 (N_13394,N_6977,N_6189);
xnor U13395 (N_13395,N_7727,N_5960);
or U13396 (N_13396,N_9323,N_8279);
xor U13397 (N_13397,N_5697,N_5408);
or U13398 (N_13398,N_9883,N_9865);
nor U13399 (N_13399,N_8001,N_5372);
nand U13400 (N_13400,N_8187,N_5201);
and U13401 (N_13401,N_5654,N_5406);
xor U13402 (N_13402,N_7024,N_6658);
nor U13403 (N_13403,N_6264,N_9564);
nand U13404 (N_13404,N_9023,N_9996);
or U13405 (N_13405,N_7289,N_8226);
or U13406 (N_13406,N_6606,N_8414);
or U13407 (N_13407,N_7515,N_7308);
nor U13408 (N_13408,N_8282,N_7070);
nand U13409 (N_13409,N_8972,N_5444);
or U13410 (N_13410,N_9288,N_7749);
and U13411 (N_13411,N_8297,N_5194);
nand U13412 (N_13412,N_7959,N_5664);
nand U13413 (N_13413,N_5338,N_7173);
and U13414 (N_13414,N_8769,N_8380);
or U13415 (N_13415,N_9567,N_6218);
xnor U13416 (N_13416,N_7406,N_6960);
nand U13417 (N_13417,N_8132,N_6239);
nor U13418 (N_13418,N_7853,N_7636);
or U13419 (N_13419,N_8866,N_5067);
xor U13420 (N_13420,N_5004,N_9636);
xnor U13421 (N_13421,N_5079,N_9646);
or U13422 (N_13422,N_6090,N_6796);
xor U13423 (N_13423,N_7019,N_9308);
or U13424 (N_13424,N_8756,N_8175);
nor U13425 (N_13425,N_7827,N_6472);
xor U13426 (N_13426,N_7619,N_5289);
nand U13427 (N_13427,N_8223,N_8010);
and U13428 (N_13428,N_8443,N_5252);
xor U13429 (N_13429,N_6833,N_9816);
xnor U13430 (N_13430,N_6754,N_9485);
nand U13431 (N_13431,N_8584,N_5336);
xor U13432 (N_13432,N_7388,N_8689);
and U13433 (N_13433,N_9871,N_8525);
or U13434 (N_13434,N_6080,N_5151);
xor U13435 (N_13435,N_7754,N_8796);
xnor U13436 (N_13436,N_5136,N_6782);
nor U13437 (N_13437,N_7607,N_7522);
and U13438 (N_13438,N_7533,N_9758);
or U13439 (N_13439,N_7991,N_6203);
and U13440 (N_13440,N_5806,N_8695);
nand U13441 (N_13441,N_5603,N_7985);
xor U13442 (N_13442,N_8135,N_5503);
or U13443 (N_13443,N_6685,N_7585);
nand U13444 (N_13444,N_9631,N_6692);
nor U13445 (N_13445,N_7350,N_9816);
nand U13446 (N_13446,N_7307,N_9375);
nor U13447 (N_13447,N_5270,N_5855);
or U13448 (N_13448,N_7414,N_7716);
and U13449 (N_13449,N_7480,N_6019);
xnor U13450 (N_13450,N_5403,N_6742);
xnor U13451 (N_13451,N_9058,N_6990);
xnor U13452 (N_13452,N_7294,N_8119);
and U13453 (N_13453,N_8730,N_5663);
nand U13454 (N_13454,N_6165,N_7055);
and U13455 (N_13455,N_9772,N_9110);
or U13456 (N_13456,N_6782,N_8609);
nor U13457 (N_13457,N_9704,N_8824);
and U13458 (N_13458,N_7351,N_9016);
or U13459 (N_13459,N_5470,N_9899);
or U13460 (N_13460,N_7275,N_6547);
and U13461 (N_13461,N_8074,N_5796);
xnor U13462 (N_13462,N_5032,N_9828);
and U13463 (N_13463,N_5615,N_9259);
xor U13464 (N_13464,N_6617,N_8419);
xor U13465 (N_13465,N_9206,N_9693);
nand U13466 (N_13466,N_7087,N_6596);
nand U13467 (N_13467,N_6933,N_8255);
nand U13468 (N_13468,N_8492,N_7541);
or U13469 (N_13469,N_7661,N_7539);
xor U13470 (N_13470,N_7839,N_5781);
xor U13471 (N_13471,N_8723,N_5021);
and U13472 (N_13472,N_9332,N_6232);
nor U13473 (N_13473,N_9300,N_8212);
and U13474 (N_13474,N_5843,N_9505);
nand U13475 (N_13475,N_6626,N_8142);
xor U13476 (N_13476,N_7870,N_9562);
nor U13477 (N_13477,N_9090,N_9365);
nor U13478 (N_13478,N_9701,N_7787);
nand U13479 (N_13479,N_9764,N_5339);
nor U13480 (N_13480,N_8161,N_9620);
or U13481 (N_13481,N_9586,N_8232);
nor U13482 (N_13482,N_7132,N_6353);
xnor U13483 (N_13483,N_6266,N_7688);
and U13484 (N_13484,N_5336,N_7191);
nand U13485 (N_13485,N_6909,N_8129);
and U13486 (N_13486,N_5741,N_6224);
nor U13487 (N_13487,N_7270,N_8707);
or U13488 (N_13488,N_5503,N_6701);
and U13489 (N_13489,N_7856,N_8970);
nand U13490 (N_13490,N_8541,N_8569);
and U13491 (N_13491,N_5443,N_8734);
or U13492 (N_13492,N_6527,N_9761);
nor U13493 (N_13493,N_6160,N_8715);
and U13494 (N_13494,N_5991,N_8701);
nand U13495 (N_13495,N_5308,N_5365);
and U13496 (N_13496,N_6192,N_6221);
and U13497 (N_13497,N_9689,N_6837);
nor U13498 (N_13498,N_6577,N_6952);
nor U13499 (N_13499,N_7596,N_9290);
and U13500 (N_13500,N_6813,N_9492);
and U13501 (N_13501,N_5103,N_8824);
nand U13502 (N_13502,N_8110,N_5919);
and U13503 (N_13503,N_5822,N_9886);
or U13504 (N_13504,N_5025,N_9781);
or U13505 (N_13505,N_8905,N_5018);
or U13506 (N_13506,N_7655,N_7521);
and U13507 (N_13507,N_5154,N_5615);
xor U13508 (N_13508,N_9377,N_5296);
or U13509 (N_13509,N_6644,N_7668);
xor U13510 (N_13510,N_7664,N_5631);
or U13511 (N_13511,N_8322,N_8170);
or U13512 (N_13512,N_6986,N_7747);
or U13513 (N_13513,N_6785,N_6958);
nand U13514 (N_13514,N_8743,N_7297);
and U13515 (N_13515,N_9190,N_6055);
and U13516 (N_13516,N_7546,N_8111);
or U13517 (N_13517,N_6854,N_5611);
or U13518 (N_13518,N_8961,N_6945);
or U13519 (N_13519,N_8679,N_7840);
or U13520 (N_13520,N_7863,N_8092);
nand U13521 (N_13521,N_8815,N_9694);
and U13522 (N_13522,N_7477,N_9449);
or U13523 (N_13523,N_8719,N_9147);
and U13524 (N_13524,N_6173,N_8637);
xor U13525 (N_13525,N_6578,N_6266);
xnor U13526 (N_13526,N_9744,N_5421);
nand U13527 (N_13527,N_7747,N_8444);
nand U13528 (N_13528,N_8084,N_6427);
and U13529 (N_13529,N_8085,N_5286);
nor U13530 (N_13530,N_7622,N_6489);
xnor U13531 (N_13531,N_9295,N_5437);
nand U13532 (N_13532,N_8524,N_9645);
nand U13533 (N_13533,N_8349,N_7741);
nand U13534 (N_13534,N_9860,N_7160);
nand U13535 (N_13535,N_6064,N_8192);
nand U13536 (N_13536,N_7857,N_8833);
nor U13537 (N_13537,N_9936,N_5915);
xor U13538 (N_13538,N_9602,N_5302);
xor U13539 (N_13539,N_8556,N_5922);
or U13540 (N_13540,N_6311,N_8654);
nand U13541 (N_13541,N_7232,N_8095);
nor U13542 (N_13542,N_8098,N_9607);
and U13543 (N_13543,N_5771,N_9346);
and U13544 (N_13544,N_8664,N_8713);
nor U13545 (N_13545,N_6045,N_6560);
and U13546 (N_13546,N_8330,N_8264);
and U13547 (N_13547,N_6110,N_5863);
and U13548 (N_13548,N_6592,N_6474);
xor U13549 (N_13549,N_5532,N_6510);
nand U13550 (N_13550,N_9489,N_8089);
or U13551 (N_13551,N_8270,N_7599);
nand U13552 (N_13552,N_5944,N_5582);
nor U13553 (N_13553,N_9378,N_8639);
nand U13554 (N_13554,N_9711,N_5174);
xor U13555 (N_13555,N_8474,N_6861);
nand U13556 (N_13556,N_9555,N_9520);
nor U13557 (N_13557,N_6620,N_5385);
and U13558 (N_13558,N_9685,N_7920);
nor U13559 (N_13559,N_6733,N_8511);
or U13560 (N_13560,N_6365,N_7182);
nor U13561 (N_13561,N_7711,N_6911);
xnor U13562 (N_13562,N_8014,N_8767);
or U13563 (N_13563,N_6797,N_6470);
nand U13564 (N_13564,N_9802,N_9913);
nor U13565 (N_13565,N_8519,N_5157);
nor U13566 (N_13566,N_5637,N_8213);
xor U13567 (N_13567,N_6598,N_9246);
nor U13568 (N_13568,N_6861,N_5258);
nor U13569 (N_13569,N_5669,N_8761);
or U13570 (N_13570,N_6047,N_5915);
nand U13571 (N_13571,N_8568,N_7676);
xnor U13572 (N_13572,N_5998,N_6907);
xor U13573 (N_13573,N_5139,N_8697);
or U13574 (N_13574,N_9063,N_8975);
or U13575 (N_13575,N_7699,N_6830);
or U13576 (N_13576,N_5174,N_6700);
xor U13577 (N_13577,N_6693,N_5907);
xnor U13578 (N_13578,N_8384,N_9647);
nor U13579 (N_13579,N_6785,N_9372);
nor U13580 (N_13580,N_8738,N_7627);
xnor U13581 (N_13581,N_9610,N_6636);
nor U13582 (N_13582,N_7703,N_5210);
or U13583 (N_13583,N_8231,N_9878);
nand U13584 (N_13584,N_9842,N_8533);
xnor U13585 (N_13585,N_8882,N_8545);
nand U13586 (N_13586,N_6164,N_9432);
and U13587 (N_13587,N_8905,N_7349);
and U13588 (N_13588,N_8393,N_9614);
or U13589 (N_13589,N_6002,N_5833);
nand U13590 (N_13590,N_7458,N_8596);
and U13591 (N_13591,N_8849,N_6985);
nand U13592 (N_13592,N_7050,N_8914);
nand U13593 (N_13593,N_8408,N_7299);
nor U13594 (N_13594,N_8984,N_6123);
or U13595 (N_13595,N_7924,N_5320);
or U13596 (N_13596,N_6706,N_7901);
and U13597 (N_13597,N_6888,N_5435);
nand U13598 (N_13598,N_5703,N_7807);
nand U13599 (N_13599,N_8827,N_5387);
and U13600 (N_13600,N_8534,N_5182);
nor U13601 (N_13601,N_6196,N_6823);
nand U13602 (N_13602,N_9742,N_9655);
xnor U13603 (N_13603,N_6033,N_7276);
and U13604 (N_13604,N_7476,N_6570);
xor U13605 (N_13605,N_9146,N_8016);
or U13606 (N_13606,N_5882,N_8048);
and U13607 (N_13607,N_9008,N_6051);
nand U13608 (N_13608,N_7859,N_8025);
and U13609 (N_13609,N_5688,N_8313);
nand U13610 (N_13610,N_6015,N_6285);
xnor U13611 (N_13611,N_7011,N_6058);
and U13612 (N_13612,N_7454,N_7994);
nor U13613 (N_13613,N_5310,N_5577);
nand U13614 (N_13614,N_7340,N_7460);
and U13615 (N_13615,N_5779,N_7541);
and U13616 (N_13616,N_8457,N_8438);
or U13617 (N_13617,N_9155,N_7895);
nand U13618 (N_13618,N_8737,N_9191);
and U13619 (N_13619,N_9280,N_7939);
nand U13620 (N_13620,N_6738,N_8793);
nor U13621 (N_13621,N_9260,N_9447);
nand U13622 (N_13622,N_7812,N_7527);
or U13623 (N_13623,N_6262,N_5937);
nand U13624 (N_13624,N_8748,N_8623);
and U13625 (N_13625,N_7827,N_6399);
nand U13626 (N_13626,N_5536,N_5699);
nand U13627 (N_13627,N_5084,N_9285);
and U13628 (N_13628,N_6304,N_7544);
or U13629 (N_13629,N_5763,N_7616);
nor U13630 (N_13630,N_9296,N_9317);
and U13631 (N_13631,N_5874,N_9508);
or U13632 (N_13632,N_6517,N_7527);
or U13633 (N_13633,N_8870,N_5585);
xor U13634 (N_13634,N_8227,N_7069);
and U13635 (N_13635,N_7857,N_7732);
nand U13636 (N_13636,N_8111,N_9695);
nand U13637 (N_13637,N_6299,N_5371);
nand U13638 (N_13638,N_7091,N_5953);
nor U13639 (N_13639,N_5690,N_6181);
or U13640 (N_13640,N_9584,N_6808);
xnor U13641 (N_13641,N_5071,N_5901);
and U13642 (N_13642,N_5649,N_7518);
nand U13643 (N_13643,N_8828,N_7438);
xor U13644 (N_13644,N_8716,N_9165);
nor U13645 (N_13645,N_8051,N_9897);
and U13646 (N_13646,N_6422,N_8727);
or U13647 (N_13647,N_6680,N_7583);
and U13648 (N_13648,N_9187,N_5064);
nor U13649 (N_13649,N_9941,N_9309);
and U13650 (N_13650,N_6017,N_7781);
or U13651 (N_13651,N_9446,N_6996);
nand U13652 (N_13652,N_7281,N_6962);
nor U13653 (N_13653,N_5189,N_8278);
and U13654 (N_13654,N_8772,N_6049);
nor U13655 (N_13655,N_9417,N_9680);
xor U13656 (N_13656,N_7846,N_8910);
nor U13657 (N_13657,N_5234,N_7028);
or U13658 (N_13658,N_9492,N_5922);
or U13659 (N_13659,N_7331,N_6312);
nand U13660 (N_13660,N_8570,N_5476);
nand U13661 (N_13661,N_9028,N_7470);
xor U13662 (N_13662,N_5108,N_6107);
nand U13663 (N_13663,N_9003,N_8875);
and U13664 (N_13664,N_5497,N_9008);
nand U13665 (N_13665,N_7287,N_5301);
or U13666 (N_13666,N_6242,N_5809);
and U13667 (N_13667,N_6696,N_8023);
nand U13668 (N_13668,N_7247,N_6975);
xor U13669 (N_13669,N_7453,N_5826);
nand U13670 (N_13670,N_5623,N_7771);
nand U13671 (N_13671,N_5853,N_5033);
nor U13672 (N_13672,N_7220,N_7070);
or U13673 (N_13673,N_7474,N_5556);
nor U13674 (N_13674,N_6631,N_6403);
or U13675 (N_13675,N_8107,N_6290);
and U13676 (N_13676,N_7634,N_9883);
nand U13677 (N_13677,N_7960,N_7597);
xor U13678 (N_13678,N_9306,N_7142);
nor U13679 (N_13679,N_9483,N_5562);
nand U13680 (N_13680,N_7348,N_7727);
and U13681 (N_13681,N_5424,N_7982);
and U13682 (N_13682,N_8224,N_6348);
nor U13683 (N_13683,N_9991,N_7266);
nor U13684 (N_13684,N_5178,N_5443);
xor U13685 (N_13685,N_9700,N_8250);
or U13686 (N_13686,N_5145,N_5980);
nand U13687 (N_13687,N_9722,N_6112);
nand U13688 (N_13688,N_8202,N_5150);
nand U13689 (N_13689,N_9528,N_7755);
or U13690 (N_13690,N_7228,N_7100);
nor U13691 (N_13691,N_6748,N_5290);
nor U13692 (N_13692,N_7355,N_8084);
nand U13693 (N_13693,N_5618,N_8981);
and U13694 (N_13694,N_9809,N_5757);
nor U13695 (N_13695,N_8844,N_9678);
xnor U13696 (N_13696,N_5887,N_9872);
nor U13697 (N_13697,N_5227,N_6366);
xor U13698 (N_13698,N_9670,N_9478);
or U13699 (N_13699,N_7988,N_6104);
or U13700 (N_13700,N_7397,N_5090);
nand U13701 (N_13701,N_8493,N_9286);
nor U13702 (N_13702,N_9573,N_8136);
or U13703 (N_13703,N_8383,N_5990);
and U13704 (N_13704,N_7122,N_9887);
nor U13705 (N_13705,N_5276,N_9519);
or U13706 (N_13706,N_6400,N_8435);
xor U13707 (N_13707,N_7079,N_7122);
nor U13708 (N_13708,N_9698,N_9791);
and U13709 (N_13709,N_7777,N_5589);
or U13710 (N_13710,N_9248,N_5474);
nand U13711 (N_13711,N_5470,N_8721);
xnor U13712 (N_13712,N_6730,N_9034);
nor U13713 (N_13713,N_7703,N_7644);
nand U13714 (N_13714,N_7372,N_5838);
nand U13715 (N_13715,N_5903,N_9542);
or U13716 (N_13716,N_7274,N_6856);
xor U13717 (N_13717,N_8478,N_5465);
or U13718 (N_13718,N_7478,N_5165);
nand U13719 (N_13719,N_6153,N_7638);
and U13720 (N_13720,N_5242,N_9867);
and U13721 (N_13721,N_5159,N_6570);
or U13722 (N_13722,N_7189,N_9907);
and U13723 (N_13723,N_9115,N_9419);
or U13724 (N_13724,N_9349,N_8260);
xor U13725 (N_13725,N_6507,N_8161);
or U13726 (N_13726,N_5771,N_5160);
nand U13727 (N_13727,N_9579,N_7811);
or U13728 (N_13728,N_7587,N_9798);
nor U13729 (N_13729,N_5930,N_5713);
and U13730 (N_13730,N_6690,N_7196);
nand U13731 (N_13731,N_9888,N_9831);
nor U13732 (N_13732,N_5236,N_7711);
nand U13733 (N_13733,N_6588,N_8933);
nand U13734 (N_13734,N_7268,N_8055);
xor U13735 (N_13735,N_9811,N_5378);
and U13736 (N_13736,N_5104,N_5315);
xor U13737 (N_13737,N_8445,N_6893);
xnor U13738 (N_13738,N_9401,N_8908);
nand U13739 (N_13739,N_6747,N_7196);
nand U13740 (N_13740,N_5589,N_8907);
and U13741 (N_13741,N_8346,N_6619);
and U13742 (N_13742,N_5333,N_8038);
nor U13743 (N_13743,N_7957,N_5539);
and U13744 (N_13744,N_5856,N_9230);
or U13745 (N_13745,N_5371,N_9966);
nand U13746 (N_13746,N_7667,N_8641);
and U13747 (N_13747,N_9431,N_6568);
nand U13748 (N_13748,N_5384,N_9290);
or U13749 (N_13749,N_7061,N_7820);
and U13750 (N_13750,N_7818,N_9404);
xnor U13751 (N_13751,N_6007,N_5445);
nand U13752 (N_13752,N_7259,N_6595);
xnor U13753 (N_13753,N_5959,N_6339);
or U13754 (N_13754,N_7632,N_9567);
xor U13755 (N_13755,N_6480,N_9186);
or U13756 (N_13756,N_8271,N_7979);
nand U13757 (N_13757,N_9146,N_7345);
nor U13758 (N_13758,N_9469,N_8688);
or U13759 (N_13759,N_9155,N_9539);
xnor U13760 (N_13760,N_6303,N_6845);
nor U13761 (N_13761,N_8246,N_8447);
and U13762 (N_13762,N_5642,N_6407);
and U13763 (N_13763,N_9354,N_8690);
nor U13764 (N_13764,N_8346,N_5884);
nand U13765 (N_13765,N_8814,N_8474);
nor U13766 (N_13766,N_6839,N_6567);
and U13767 (N_13767,N_6137,N_9901);
xnor U13768 (N_13768,N_5241,N_6800);
or U13769 (N_13769,N_5426,N_7845);
and U13770 (N_13770,N_7669,N_5574);
nand U13771 (N_13771,N_9894,N_7098);
nand U13772 (N_13772,N_8321,N_9964);
nand U13773 (N_13773,N_5020,N_7201);
and U13774 (N_13774,N_7794,N_6985);
nor U13775 (N_13775,N_5686,N_8805);
nor U13776 (N_13776,N_9585,N_9481);
nor U13777 (N_13777,N_7048,N_8439);
and U13778 (N_13778,N_8974,N_5086);
and U13779 (N_13779,N_9016,N_5685);
or U13780 (N_13780,N_8013,N_7063);
nand U13781 (N_13781,N_9578,N_5176);
or U13782 (N_13782,N_9600,N_6848);
or U13783 (N_13783,N_7081,N_5574);
nand U13784 (N_13784,N_8368,N_9448);
nand U13785 (N_13785,N_6788,N_5812);
or U13786 (N_13786,N_7382,N_8833);
and U13787 (N_13787,N_8639,N_5731);
and U13788 (N_13788,N_8219,N_9747);
xor U13789 (N_13789,N_7454,N_5703);
nand U13790 (N_13790,N_7977,N_8191);
and U13791 (N_13791,N_8690,N_9407);
nand U13792 (N_13792,N_9303,N_7814);
and U13793 (N_13793,N_5955,N_9750);
xnor U13794 (N_13794,N_7994,N_5983);
nor U13795 (N_13795,N_5236,N_6304);
or U13796 (N_13796,N_6402,N_6231);
and U13797 (N_13797,N_5771,N_9256);
or U13798 (N_13798,N_8593,N_5757);
and U13799 (N_13799,N_6400,N_6755);
xnor U13800 (N_13800,N_9243,N_8651);
or U13801 (N_13801,N_6820,N_5947);
nand U13802 (N_13802,N_9137,N_9951);
and U13803 (N_13803,N_8688,N_5795);
nand U13804 (N_13804,N_5030,N_8995);
nor U13805 (N_13805,N_9907,N_5060);
and U13806 (N_13806,N_5282,N_8704);
nand U13807 (N_13807,N_5006,N_8591);
xor U13808 (N_13808,N_9026,N_9722);
nor U13809 (N_13809,N_5537,N_5458);
nand U13810 (N_13810,N_8709,N_5348);
and U13811 (N_13811,N_6798,N_5178);
or U13812 (N_13812,N_6341,N_6230);
xor U13813 (N_13813,N_9936,N_8312);
nand U13814 (N_13814,N_8653,N_8382);
xnor U13815 (N_13815,N_7910,N_5503);
xor U13816 (N_13816,N_6778,N_7722);
or U13817 (N_13817,N_8363,N_7279);
nor U13818 (N_13818,N_7745,N_5447);
or U13819 (N_13819,N_9186,N_7908);
and U13820 (N_13820,N_6310,N_7908);
xor U13821 (N_13821,N_8644,N_9851);
nor U13822 (N_13822,N_8775,N_6737);
nand U13823 (N_13823,N_5387,N_6702);
nand U13824 (N_13824,N_7647,N_9328);
and U13825 (N_13825,N_8994,N_7547);
and U13826 (N_13826,N_7419,N_5068);
and U13827 (N_13827,N_5533,N_9799);
xnor U13828 (N_13828,N_8602,N_8987);
nor U13829 (N_13829,N_8321,N_6577);
and U13830 (N_13830,N_6641,N_8297);
and U13831 (N_13831,N_6941,N_9676);
or U13832 (N_13832,N_7896,N_5501);
and U13833 (N_13833,N_5626,N_6606);
nand U13834 (N_13834,N_9407,N_5593);
nand U13835 (N_13835,N_5984,N_5836);
nand U13836 (N_13836,N_8760,N_5581);
xnor U13837 (N_13837,N_7023,N_6443);
or U13838 (N_13838,N_8813,N_5830);
nand U13839 (N_13839,N_9308,N_9916);
nand U13840 (N_13840,N_7332,N_9406);
nand U13841 (N_13841,N_9033,N_6928);
or U13842 (N_13842,N_6854,N_7224);
xor U13843 (N_13843,N_9683,N_5052);
or U13844 (N_13844,N_7494,N_9780);
xor U13845 (N_13845,N_6503,N_5245);
nand U13846 (N_13846,N_6190,N_9887);
and U13847 (N_13847,N_9999,N_6262);
xor U13848 (N_13848,N_9018,N_6815);
or U13849 (N_13849,N_7067,N_6073);
nor U13850 (N_13850,N_6486,N_8944);
nand U13851 (N_13851,N_6595,N_8849);
xor U13852 (N_13852,N_9823,N_7065);
and U13853 (N_13853,N_8868,N_7630);
nand U13854 (N_13854,N_6756,N_9864);
nand U13855 (N_13855,N_5173,N_5639);
or U13856 (N_13856,N_7700,N_7440);
and U13857 (N_13857,N_5898,N_7761);
nor U13858 (N_13858,N_8799,N_5172);
and U13859 (N_13859,N_8325,N_8801);
nor U13860 (N_13860,N_8896,N_6511);
or U13861 (N_13861,N_7553,N_5330);
xor U13862 (N_13862,N_9490,N_7799);
nor U13863 (N_13863,N_9942,N_8724);
nor U13864 (N_13864,N_9724,N_9696);
xnor U13865 (N_13865,N_8814,N_5629);
nand U13866 (N_13866,N_7751,N_5055);
nor U13867 (N_13867,N_8289,N_9898);
and U13868 (N_13868,N_6138,N_8241);
and U13869 (N_13869,N_5009,N_7138);
xnor U13870 (N_13870,N_7156,N_8156);
nand U13871 (N_13871,N_6495,N_6689);
nor U13872 (N_13872,N_6978,N_8472);
or U13873 (N_13873,N_8317,N_7220);
or U13874 (N_13874,N_5617,N_5689);
xnor U13875 (N_13875,N_6342,N_8546);
or U13876 (N_13876,N_9601,N_6816);
and U13877 (N_13877,N_8450,N_6820);
nand U13878 (N_13878,N_8024,N_7605);
xor U13879 (N_13879,N_9261,N_6746);
xor U13880 (N_13880,N_6508,N_7936);
or U13881 (N_13881,N_7298,N_8082);
nand U13882 (N_13882,N_6309,N_5781);
xnor U13883 (N_13883,N_6987,N_6358);
or U13884 (N_13884,N_7932,N_7469);
and U13885 (N_13885,N_7161,N_5625);
or U13886 (N_13886,N_9302,N_6877);
xnor U13887 (N_13887,N_8627,N_9800);
nor U13888 (N_13888,N_6254,N_8709);
or U13889 (N_13889,N_8234,N_5266);
nand U13890 (N_13890,N_6160,N_6145);
nor U13891 (N_13891,N_8209,N_7869);
nor U13892 (N_13892,N_7063,N_8645);
nor U13893 (N_13893,N_6128,N_6783);
nand U13894 (N_13894,N_5032,N_5241);
nand U13895 (N_13895,N_8405,N_8770);
and U13896 (N_13896,N_8442,N_7376);
xnor U13897 (N_13897,N_6337,N_6859);
or U13898 (N_13898,N_9093,N_7808);
nor U13899 (N_13899,N_8960,N_5862);
nor U13900 (N_13900,N_5074,N_8995);
nor U13901 (N_13901,N_7490,N_9058);
xor U13902 (N_13902,N_7296,N_9727);
or U13903 (N_13903,N_9247,N_9408);
nand U13904 (N_13904,N_6158,N_6525);
and U13905 (N_13905,N_9957,N_6138);
nor U13906 (N_13906,N_8071,N_8483);
xor U13907 (N_13907,N_5350,N_7611);
nand U13908 (N_13908,N_6576,N_6811);
xnor U13909 (N_13909,N_8053,N_5843);
or U13910 (N_13910,N_9052,N_5719);
xor U13911 (N_13911,N_9399,N_9989);
or U13912 (N_13912,N_8164,N_5886);
or U13913 (N_13913,N_5171,N_8275);
nor U13914 (N_13914,N_9370,N_6736);
nor U13915 (N_13915,N_9010,N_7006);
xnor U13916 (N_13916,N_5672,N_8476);
nor U13917 (N_13917,N_8125,N_9310);
nand U13918 (N_13918,N_8392,N_5341);
nor U13919 (N_13919,N_9467,N_6226);
nor U13920 (N_13920,N_9121,N_5322);
and U13921 (N_13921,N_8838,N_5461);
or U13922 (N_13922,N_7075,N_5507);
xnor U13923 (N_13923,N_9681,N_8620);
nand U13924 (N_13924,N_8438,N_9379);
nor U13925 (N_13925,N_8579,N_6425);
xnor U13926 (N_13926,N_6913,N_9664);
and U13927 (N_13927,N_6026,N_9912);
nand U13928 (N_13928,N_5629,N_8059);
and U13929 (N_13929,N_7182,N_7936);
and U13930 (N_13930,N_7373,N_5649);
nor U13931 (N_13931,N_5368,N_8727);
nor U13932 (N_13932,N_5448,N_8911);
or U13933 (N_13933,N_5633,N_8111);
or U13934 (N_13934,N_9423,N_9789);
nand U13935 (N_13935,N_7050,N_5744);
or U13936 (N_13936,N_6198,N_6545);
xnor U13937 (N_13937,N_7252,N_8589);
nand U13938 (N_13938,N_9868,N_7321);
nor U13939 (N_13939,N_7526,N_6810);
or U13940 (N_13940,N_8024,N_9600);
or U13941 (N_13941,N_7543,N_9437);
and U13942 (N_13942,N_9955,N_7722);
and U13943 (N_13943,N_6609,N_9084);
and U13944 (N_13944,N_7914,N_9725);
xnor U13945 (N_13945,N_9462,N_8309);
and U13946 (N_13946,N_5769,N_8670);
nor U13947 (N_13947,N_7072,N_9220);
nand U13948 (N_13948,N_7162,N_9745);
xnor U13949 (N_13949,N_5775,N_9811);
nand U13950 (N_13950,N_8007,N_7591);
and U13951 (N_13951,N_7410,N_9713);
or U13952 (N_13952,N_6822,N_9181);
nand U13953 (N_13953,N_7147,N_5580);
xor U13954 (N_13954,N_7559,N_6988);
nand U13955 (N_13955,N_8343,N_5936);
nor U13956 (N_13956,N_8847,N_8725);
and U13957 (N_13957,N_7316,N_5561);
or U13958 (N_13958,N_5423,N_9097);
xor U13959 (N_13959,N_8161,N_8630);
nand U13960 (N_13960,N_7261,N_6233);
nor U13961 (N_13961,N_9129,N_5897);
or U13962 (N_13962,N_7761,N_5434);
nor U13963 (N_13963,N_6951,N_6950);
nand U13964 (N_13964,N_6844,N_8257);
nand U13965 (N_13965,N_6941,N_5422);
nor U13966 (N_13966,N_7724,N_8092);
nand U13967 (N_13967,N_6453,N_9259);
xnor U13968 (N_13968,N_5886,N_5958);
and U13969 (N_13969,N_6684,N_7474);
nand U13970 (N_13970,N_8188,N_8264);
xor U13971 (N_13971,N_8527,N_9059);
nor U13972 (N_13972,N_8926,N_8245);
xnor U13973 (N_13973,N_5683,N_5807);
nand U13974 (N_13974,N_5087,N_7965);
xor U13975 (N_13975,N_6843,N_7020);
or U13976 (N_13976,N_6314,N_8192);
nand U13977 (N_13977,N_5181,N_7230);
or U13978 (N_13978,N_7695,N_5974);
nand U13979 (N_13979,N_7918,N_7479);
and U13980 (N_13980,N_6629,N_5529);
nand U13981 (N_13981,N_8905,N_7189);
nand U13982 (N_13982,N_8935,N_7608);
and U13983 (N_13983,N_8715,N_9894);
or U13984 (N_13984,N_5808,N_7949);
and U13985 (N_13985,N_6660,N_8208);
and U13986 (N_13986,N_6909,N_7034);
xnor U13987 (N_13987,N_7682,N_9552);
xnor U13988 (N_13988,N_9056,N_5253);
and U13989 (N_13989,N_8924,N_9086);
or U13990 (N_13990,N_7661,N_9130);
nor U13991 (N_13991,N_7499,N_8341);
or U13992 (N_13992,N_9316,N_9351);
and U13993 (N_13993,N_5055,N_5818);
or U13994 (N_13994,N_5393,N_9811);
xnor U13995 (N_13995,N_9357,N_6700);
nor U13996 (N_13996,N_6972,N_8094);
and U13997 (N_13997,N_7691,N_7892);
and U13998 (N_13998,N_7977,N_8329);
xor U13999 (N_13999,N_8235,N_5812);
nand U14000 (N_14000,N_6552,N_9430);
and U14001 (N_14001,N_8625,N_6274);
xnor U14002 (N_14002,N_8789,N_6882);
nand U14003 (N_14003,N_8728,N_5092);
or U14004 (N_14004,N_8435,N_6439);
xnor U14005 (N_14005,N_9383,N_9655);
xor U14006 (N_14006,N_9025,N_7568);
nand U14007 (N_14007,N_7799,N_5772);
nand U14008 (N_14008,N_7341,N_7117);
or U14009 (N_14009,N_5770,N_9013);
and U14010 (N_14010,N_7811,N_9060);
nand U14011 (N_14011,N_8777,N_9665);
xnor U14012 (N_14012,N_8977,N_6410);
nand U14013 (N_14013,N_8083,N_9962);
nand U14014 (N_14014,N_9893,N_7404);
and U14015 (N_14015,N_8731,N_7993);
nand U14016 (N_14016,N_7971,N_9941);
nand U14017 (N_14017,N_7697,N_5084);
xnor U14018 (N_14018,N_5370,N_9632);
or U14019 (N_14019,N_7949,N_8950);
xnor U14020 (N_14020,N_5276,N_5864);
and U14021 (N_14021,N_9929,N_6455);
nor U14022 (N_14022,N_5453,N_7369);
xor U14023 (N_14023,N_8233,N_8358);
nor U14024 (N_14024,N_7814,N_8867);
xnor U14025 (N_14025,N_6593,N_7475);
xor U14026 (N_14026,N_5095,N_9775);
nor U14027 (N_14027,N_5605,N_9364);
and U14028 (N_14028,N_7193,N_7242);
nor U14029 (N_14029,N_5129,N_6887);
xnor U14030 (N_14030,N_8989,N_8553);
xor U14031 (N_14031,N_8887,N_7576);
nand U14032 (N_14032,N_8869,N_8255);
and U14033 (N_14033,N_9603,N_5019);
and U14034 (N_14034,N_8254,N_7197);
and U14035 (N_14035,N_9073,N_9236);
or U14036 (N_14036,N_7068,N_8130);
nor U14037 (N_14037,N_7495,N_7517);
and U14038 (N_14038,N_6652,N_8614);
nand U14039 (N_14039,N_9387,N_5666);
nand U14040 (N_14040,N_6929,N_8642);
xor U14041 (N_14041,N_5122,N_7738);
xor U14042 (N_14042,N_7783,N_9758);
and U14043 (N_14043,N_7810,N_6556);
xor U14044 (N_14044,N_6132,N_7642);
nand U14045 (N_14045,N_7534,N_9860);
xor U14046 (N_14046,N_8340,N_5977);
and U14047 (N_14047,N_5522,N_6433);
or U14048 (N_14048,N_6506,N_5121);
and U14049 (N_14049,N_9057,N_8092);
or U14050 (N_14050,N_6966,N_7275);
nand U14051 (N_14051,N_6963,N_6894);
nor U14052 (N_14052,N_8977,N_8485);
nor U14053 (N_14053,N_5885,N_9029);
nor U14054 (N_14054,N_7853,N_8622);
xnor U14055 (N_14055,N_9932,N_5999);
xnor U14056 (N_14056,N_7519,N_5742);
nand U14057 (N_14057,N_8361,N_9722);
nand U14058 (N_14058,N_5845,N_8050);
xnor U14059 (N_14059,N_7096,N_6233);
or U14060 (N_14060,N_9578,N_7589);
and U14061 (N_14061,N_6358,N_9673);
nand U14062 (N_14062,N_8456,N_7892);
and U14063 (N_14063,N_9723,N_6378);
xor U14064 (N_14064,N_7811,N_7645);
nor U14065 (N_14065,N_8764,N_8188);
and U14066 (N_14066,N_5360,N_9133);
xnor U14067 (N_14067,N_9225,N_7593);
and U14068 (N_14068,N_7397,N_5277);
nor U14069 (N_14069,N_7887,N_8626);
nand U14070 (N_14070,N_9237,N_7533);
and U14071 (N_14071,N_9872,N_9318);
and U14072 (N_14072,N_7998,N_7591);
and U14073 (N_14073,N_7938,N_6316);
and U14074 (N_14074,N_7241,N_6268);
nor U14075 (N_14075,N_9098,N_9910);
nand U14076 (N_14076,N_5674,N_8821);
xnor U14077 (N_14077,N_8652,N_5494);
or U14078 (N_14078,N_6571,N_5174);
nand U14079 (N_14079,N_8602,N_5442);
or U14080 (N_14080,N_6222,N_9593);
xnor U14081 (N_14081,N_9667,N_7652);
xor U14082 (N_14082,N_9203,N_5776);
nand U14083 (N_14083,N_6834,N_5794);
or U14084 (N_14084,N_6076,N_9735);
xnor U14085 (N_14085,N_6591,N_9148);
xnor U14086 (N_14086,N_5693,N_9303);
and U14087 (N_14087,N_9142,N_5720);
and U14088 (N_14088,N_5226,N_5977);
and U14089 (N_14089,N_6668,N_6628);
xnor U14090 (N_14090,N_9449,N_9071);
or U14091 (N_14091,N_6991,N_7610);
nor U14092 (N_14092,N_7460,N_5290);
or U14093 (N_14093,N_6219,N_5983);
and U14094 (N_14094,N_7641,N_6284);
and U14095 (N_14095,N_7150,N_7318);
and U14096 (N_14096,N_5610,N_8930);
or U14097 (N_14097,N_9476,N_5812);
nor U14098 (N_14098,N_8758,N_9294);
or U14099 (N_14099,N_7648,N_5498);
nor U14100 (N_14100,N_9591,N_5604);
or U14101 (N_14101,N_7567,N_6566);
or U14102 (N_14102,N_6278,N_5892);
nand U14103 (N_14103,N_7424,N_5149);
and U14104 (N_14104,N_9150,N_7227);
nor U14105 (N_14105,N_7011,N_5798);
nand U14106 (N_14106,N_5081,N_7490);
xor U14107 (N_14107,N_7742,N_9884);
xnor U14108 (N_14108,N_6683,N_5610);
nand U14109 (N_14109,N_7587,N_9680);
nor U14110 (N_14110,N_6567,N_6068);
nand U14111 (N_14111,N_5935,N_5228);
and U14112 (N_14112,N_6669,N_9601);
nand U14113 (N_14113,N_5463,N_7866);
or U14114 (N_14114,N_8130,N_6617);
and U14115 (N_14115,N_9501,N_9982);
and U14116 (N_14116,N_8685,N_9414);
xnor U14117 (N_14117,N_6428,N_6332);
nor U14118 (N_14118,N_9771,N_6853);
nand U14119 (N_14119,N_5967,N_8204);
or U14120 (N_14120,N_5566,N_5784);
nand U14121 (N_14121,N_9984,N_9344);
and U14122 (N_14122,N_6475,N_8244);
and U14123 (N_14123,N_7493,N_7074);
xor U14124 (N_14124,N_8613,N_8423);
or U14125 (N_14125,N_7092,N_5289);
or U14126 (N_14126,N_6021,N_9384);
xor U14127 (N_14127,N_6924,N_5966);
or U14128 (N_14128,N_5643,N_8840);
or U14129 (N_14129,N_7825,N_5847);
or U14130 (N_14130,N_8358,N_5074);
xnor U14131 (N_14131,N_7503,N_5550);
xor U14132 (N_14132,N_5603,N_9995);
nand U14133 (N_14133,N_8597,N_6252);
xnor U14134 (N_14134,N_6669,N_9172);
or U14135 (N_14135,N_8975,N_9112);
nor U14136 (N_14136,N_8762,N_7504);
nor U14137 (N_14137,N_8371,N_9179);
and U14138 (N_14138,N_5799,N_6064);
and U14139 (N_14139,N_7470,N_9743);
or U14140 (N_14140,N_8812,N_5004);
and U14141 (N_14141,N_9601,N_7075);
nand U14142 (N_14142,N_5772,N_6711);
and U14143 (N_14143,N_5378,N_9399);
or U14144 (N_14144,N_9955,N_5109);
nand U14145 (N_14145,N_6089,N_7241);
or U14146 (N_14146,N_7583,N_7264);
xnor U14147 (N_14147,N_9012,N_5016);
nor U14148 (N_14148,N_8572,N_8412);
nand U14149 (N_14149,N_5448,N_9510);
nand U14150 (N_14150,N_7461,N_7608);
nand U14151 (N_14151,N_8190,N_7687);
or U14152 (N_14152,N_7151,N_9551);
xnor U14153 (N_14153,N_6538,N_7427);
nand U14154 (N_14154,N_8336,N_8168);
or U14155 (N_14155,N_7182,N_9472);
nand U14156 (N_14156,N_7820,N_8752);
nor U14157 (N_14157,N_6339,N_7744);
xnor U14158 (N_14158,N_9309,N_8173);
nand U14159 (N_14159,N_5128,N_7208);
nand U14160 (N_14160,N_7649,N_7266);
nor U14161 (N_14161,N_5120,N_7947);
nor U14162 (N_14162,N_6568,N_7215);
xnor U14163 (N_14163,N_6727,N_5638);
nand U14164 (N_14164,N_8523,N_7697);
xor U14165 (N_14165,N_6112,N_5463);
nand U14166 (N_14166,N_6156,N_6837);
nand U14167 (N_14167,N_7149,N_6784);
or U14168 (N_14168,N_6827,N_7696);
or U14169 (N_14169,N_6965,N_6167);
xnor U14170 (N_14170,N_9134,N_6957);
and U14171 (N_14171,N_9662,N_7039);
or U14172 (N_14172,N_8192,N_9594);
xnor U14173 (N_14173,N_5645,N_8125);
nor U14174 (N_14174,N_7742,N_9328);
nand U14175 (N_14175,N_9119,N_6529);
or U14176 (N_14176,N_7342,N_5161);
nor U14177 (N_14177,N_6444,N_8954);
nand U14178 (N_14178,N_6642,N_7089);
and U14179 (N_14179,N_6979,N_5683);
nand U14180 (N_14180,N_8777,N_8714);
and U14181 (N_14181,N_8224,N_7547);
and U14182 (N_14182,N_5298,N_7397);
nor U14183 (N_14183,N_8083,N_9844);
xor U14184 (N_14184,N_8014,N_9119);
or U14185 (N_14185,N_8608,N_8505);
nand U14186 (N_14186,N_8275,N_8899);
xnor U14187 (N_14187,N_8721,N_5773);
or U14188 (N_14188,N_7810,N_9410);
nor U14189 (N_14189,N_9270,N_9364);
and U14190 (N_14190,N_8731,N_9940);
xor U14191 (N_14191,N_8776,N_7017);
xor U14192 (N_14192,N_7127,N_5719);
nand U14193 (N_14193,N_6107,N_9327);
and U14194 (N_14194,N_6091,N_8227);
nor U14195 (N_14195,N_7298,N_7340);
nor U14196 (N_14196,N_5901,N_9211);
xnor U14197 (N_14197,N_7217,N_7986);
xor U14198 (N_14198,N_7966,N_8581);
nand U14199 (N_14199,N_6327,N_7752);
nand U14200 (N_14200,N_6233,N_8540);
or U14201 (N_14201,N_6613,N_6804);
nand U14202 (N_14202,N_7343,N_6033);
or U14203 (N_14203,N_6434,N_9207);
nor U14204 (N_14204,N_6728,N_9034);
xor U14205 (N_14205,N_5836,N_6816);
or U14206 (N_14206,N_7686,N_8391);
nand U14207 (N_14207,N_6805,N_6808);
and U14208 (N_14208,N_6957,N_7513);
nor U14209 (N_14209,N_8375,N_7215);
xnor U14210 (N_14210,N_8919,N_5095);
and U14211 (N_14211,N_5891,N_6387);
xor U14212 (N_14212,N_7095,N_7216);
and U14213 (N_14213,N_8534,N_7442);
nand U14214 (N_14214,N_9219,N_9373);
xnor U14215 (N_14215,N_8873,N_6857);
and U14216 (N_14216,N_8507,N_8285);
nand U14217 (N_14217,N_5183,N_9894);
xnor U14218 (N_14218,N_5189,N_9438);
nor U14219 (N_14219,N_5464,N_6909);
xnor U14220 (N_14220,N_6514,N_7015);
nor U14221 (N_14221,N_8630,N_5262);
xnor U14222 (N_14222,N_5723,N_9328);
xnor U14223 (N_14223,N_7043,N_8877);
or U14224 (N_14224,N_5924,N_6301);
xor U14225 (N_14225,N_7328,N_8461);
and U14226 (N_14226,N_8954,N_5150);
or U14227 (N_14227,N_8645,N_8529);
or U14228 (N_14228,N_8153,N_6112);
and U14229 (N_14229,N_7718,N_5284);
or U14230 (N_14230,N_9177,N_7028);
and U14231 (N_14231,N_7685,N_7920);
xnor U14232 (N_14232,N_9275,N_8666);
xnor U14233 (N_14233,N_9969,N_8813);
nor U14234 (N_14234,N_7152,N_7834);
xnor U14235 (N_14235,N_5783,N_9561);
xor U14236 (N_14236,N_8828,N_5805);
nand U14237 (N_14237,N_7431,N_7574);
nand U14238 (N_14238,N_7530,N_7785);
nor U14239 (N_14239,N_8488,N_8220);
or U14240 (N_14240,N_5692,N_5227);
nand U14241 (N_14241,N_8931,N_6632);
nand U14242 (N_14242,N_6043,N_7795);
nand U14243 (N_14243,N_5313,N_9829);
and U14244 (N_14244,N_6394,N_9819);
or U14245 (N_14245,N_7618,N_7534);
nand U14246 (N_14246,N_7171,N_5520);
nand U14247 (N_14247,N_9316,N_7420);
or U14248 (N_14248,N_6533,N_7135);
xor U14249 (N_14249,N_9306,N_6974);
nand U14250 (N_14250,N_6404,N_9478);
xnor U14251 (N_14251,N_6302,N_5403);
nor U14252 (N_14252,N_9623,N_5798);
nand U14253 (N_14253,N_5854,N_9101);
or U14254 (N_14254,N_8036,N_8051);
nor U14255 (N_14255,N_8374,N_6927);
or U14256 (N_14256,N_6071,N_8602);
nor U14257 (N_14257,N_9286,N_9769);
nor U14258 (N_14258,N_9220,N_5423);
xor U14259 (N_14259,N_5047,N_8541);
xnor U14260 (N_14260,N_5218,N_7708);
and U14261 (N_14261,N_6020,N_5250);
nand U14262 (N_14262,N_6372,N_9461);
and U14263 (N_14263,N_5568,N_9713);
or U14264 (N_14264,N_8950,N_5221);
nor U14265 (N_14265,N_5752,N_7248);
xnor U14266 (N_14266,N_9288,N_8480);
xor U14267 (N_14267,N_9597,N_6062);
or U14268 (N_14268,N_5495,N_6915);
xor U14269 (N_14269,N_8905,N_9485);
nor U14270 (N_14270,N_7906,N_5952);
xor U14271 (N_14271,N_9550,N_8150);
nand U14272 (N_14272,N_7202,N_8597);
xnor U14273 (N_14273,N_7103,N_6776);
nand U14274 (N_14274,N_5394,N_6045);
xor U14275 (N_14275,N_7356,N_9474);
nor U14276 (N_14276,N_6083,N_9178);
and U14277 (N_14277,N_5471,N_6052);
xor U14278 (N_14278,N_5567,N_6883);
nand U14279 (N_14279,N_5179,N_5758);
nand U14280 (N_14280,N_8271,N_8839);
xor U14281 (N_14281,N_8445,N_5708);
nor U14282 (N_14282,N_5040,N_7652);
and U14283 (N_14283,N_8069,N_9975);
and U14284 (N_14284,N_7815,N_5764);
nor U14285 (N_14285,N_9485,N_6499);
or U14286 (N_14286,N_9687,N_8876);
or U14287 (N_14287,N_7710,N_7640);
and U14288 (N_14288,N_7214,N_8557);
nand U14289 (N_14289,N_6000,N_6874);
nand U14290 (N_14290,N_6476,N_8023);
and U14291 (N_14291,N_9881,N_6373);
xor U14292 (N_14292,N_6427,N_6845);
xor U14293 (N_14293,N_7708,N_7270);
nor U14294 (N_14294,N_7296,N_5017);
xor U14295 (N_14295,N_9056,N_9884);
nand U14296 (N_14296,N_7680,N_8066);
nor U14297 (N_14297,N_8460,N_6451);
and U14298 (N_14298,N_9390,N_8182);
nand U14299 (N_14299,N_5656,N_5413);
and U14300 (N_14300,N_5614,N_9224);
nand U14301 (N_14301,N_8298,N_6672);
or U14302 (N_14302,N_8774,N_5701);
xnor U14303 (N_14303,N_6220,N_5307);
and U14304 (N_14304,N_6609,N_9076);
xnor U14305 (N_14305,N_7624,N_7977);
nand U14306 (N_14306,N_7291,N_8102);
nand U14307 (N_14307,N_8274,N_9413);
nand U14308 (N_14308,N_7376,N_6101);
or U14309 (N_14309,N_9576,N_8272);
nand U14310 (N_14310,N_9430,N_7395);
nand U14311 (N_14311,N_6648,N_8806);
nor U14312 (N_14312,N_8384,N_7634);
xor U14313 (N_14313,N_6527,N_5544);
or U14314 (N_14314,N_8387,N_6285);
and U14315 (N_14315,N_5618,N_8285);
and U14316 (N_14316,N_8206,N_8318);
nand U14317 (N_14317,N_6466,N_9608);
nand U14318 (N_14318,N_7110,N_7255);
xor U14319 (N_14319,N_9942,N_8117);
nand U14320 (N_14320,N_6778,N_5895);
nor U14321 (N_14321,N_8732,N_7701);
nor U14322 (N_14322,N_5719,N_8687);
nor U14323 (N_14323,N_6711,N_8296);
nor U14324 (N_14324,N_6544,N_8844);
and U14325 (N_14325,N_8962,N_7534);
nor U14326 (N_14326,N_6801,N_9814);
xor U14327 (N_14327,N_6674,N_5556);
or U14328 (N_14328,N_5957,N_7995);
and U14329 (N_14329,N_6122,N_6360);
xor U14330 (N_14330,N_5179,N_6746);
or U14331 (N_14331,N_9357,N_9156);
and U14332 (N_14332,N_5238,N_9452);
and U14333 (N_14333,N_6335,N_6886);
nand U14334 (N_14334,N_5243,N_6450);
nor U14335 (N_14335,N_7504,N_8683);
xor U14336 (N_14336,N_9442,N_7869);
or U14337 (N_14337,N_6548,N_7443);
and U14338 (N_14338,N_7842,N_5634);
and U14339 (N_14339,N_7626,N_7732);
nand U14340 (N_14340,N_5750,N_8551);
and U14341 (N_14341,N_7113,N_8065);
xor U14342 (N_14342,N_9191,N_6205);
xnor U14343 (N_14343,N_9118,N_7324);
and U14344 (N_14344,N_6804,N_6275);
and U14345 (N_14345,N_5170,N_7143);
or U14346 (N_14346,N_5195,N_5267);
nor U14347 (N_14347,N_6990,N_7083);
nor U14348 (N_14348,N_5424,N_7313);
nand U14349 (N_14349,N_7202,N_5957);
and U14350 (N_14350,N_7634,N_6553);
nor U14351 (N_14351,N_8667,N_6332);
nor U14352 (N_14352,N_9893,N_7301);
and U14353 (N_14353,N_6207,N_6631);
and U14354 (N_14354,N_6992,N_5866);
nor U14355 (N_14355,N_7031,N_9494);
and U14356 (N_14356,N_8471,N_6749);
nand U14357 (N_14357,N_8606,N_7427);
and U14358 (N_14358,N_5314,N_9793);
xor U14359 (N_14359,N_9067,N_6813);
xor U14360 (N_14360,N_9836,N_5761);
nor U14361 (N_14361,N_9584,N_6052);
nand U14362 (N_14362,N_8241,N_5731);
nor U14363 (N_14363,N_6742,N_9483);
or U14364 (N_14364,N_7546,N_7395);
nand U14365 (N_14365,N_9475,N_7571);
xnor U14366 (N_14366,N_6984,N_8196);
xor U14367 (N_14367,N_6190,N_6767);
nor U14368 (N_14368,N_8284,N_9128);
nor U14369 (N_14369,N_8684,N_6683);
nor U14370 (N_14370,N_6781,N_6790);
nor U14371 (N_14371,N_7984,N_7619);
nor U14372 (N_14372,N_7328,N_8312);
or U14373 (N_14373,N_8350,N_9941);
or U14374 (N_14374,N_9188,N_6583);
xnor U14375 (N_14375,N_7811,N_8019);
nand U14376 (N_14376,N_8565,N_9950);
or U14377 (N_14377,N_9289,N_7882);
nor U14378 (N_14378,N_8159,N_6200);
or U14379 (N_14379,N_9518,N_9224);
and U14380 (N_14380,N_8316,N_7140);
and U14381 (N_14381,N_9241,N_7360);
nor U14382 (N_14382,N_7524,N_8996);
nand U14383 (N_14383,N_5415,N_6085);
or U14384 (N_14384,N_6459,N_5910);
nand U14385 (N_14385,N_9621,N_9108);
nor U14386 (N_14386,N_8269,N_6612);
and U14387 (N_14387,N_5255,N_8873);
xnor U14388 (N_14388,N_9352,N_7308);
or U14389 (N_14389,N_7540,N_6259);
or U14390 (N_14390,N_5780,N_8044);
nor U14391 (N_14391,N_5012,N_5077);
and U14392 (N_14392,N_6201,N_9217);
xnor U14393 (N_14393,N_8585,N_5776);
xnor U14394 (N_14394,N_9247,N_5142);
nor U14395 (N_14395,N_7502,N_9940);
nor U14396 (N_14396,N_5457,N_7585);
nand U14397 (N_14397,N_9110,N_8519);
and U14398 (N_14398,N_9499,N_7549);
nor U14399 (N_14399,N_8172,N_8705);
nor U14400 (N_14400,N_8922,N_7015);
xor U14401 (N_14401,N_9272,N_8121);
nor U14402 (N_14402,N_8436,N_5158);
nor U14403 (N_14403,N_7911,N_8912);
or U14404 (N_14404,N_8879,N_9810);
or U14405 (N_14405,N_6611,N_7207);
and U14406 (N_14406,N_9167,N_7491);
or U14407 (N_14407,N_6145,N_7128);
nor U14408 (N_14408,N_7590,N_8812);
and U14409 (N_14409,N_5581,N_8153);
xor U14410 (N_14410,N_8564,N_6184);
or U14411 (N_14411,N_8438,N_9304);
or U14412 (N_14412,N_8246,N_5013);
and U14413 (N_14413,N_8797,N_6234);
or U14414 (N_14414,N_7035,N_6985);
or U14415 (N_14415,N_7343,N_8228);
or U14416 (N_14416,N_8810,N_7857);
xor U14417 (N_14417,N_8161,N_6185);
nand U14418 (N_14418,N_6404,N_9953);
and U14419 (N_14419,N_8062,N_7077);
and U14420 (N_14420,N_8166,N_5909);
nand U14421 (N_14421,N_6246,N_8347);
or U14422 (N_14422,N_9373,N_7319);
and U14423 (N_14423,N_7211,N_5515);
nand U14424 (N_14424,N_6342,N_8460);
or U14425 (N_14425,N_7418,N_8693);
nand U14426 (N_14426,N_8060,N_5259);
nand U14427 (N_14427,N_9951,N_7670);
or U14428 (N_14428,N_7480,N_7320);
nand U14429 (N_14429,N_8061,N_9728);
nand U14430 (N_14430,N_8701,N_9922);
or U14431 (N_14431,N_7943,N_9955);
nor U14432 (N_14432,N_9280,N_8467);
xor U14433 (N_14433,N_7908,N_9756);
xnor U14434 (N_14434,N_9971,N_7337);
and U14435 (N_14435,N_9217,N_9544);
nor U14436 (N_14436,N_9097,N_5395);
xor U14437 (N_14437,N_6358,N_6911);
xnor U14438 (N_14438,N_9734,N_6234);
and U14439 (N_14439,N_6916,N_5421);
nor U14440 (N_14440,N_8678,N_6186);
and U14441 (N_14441,N_5580,N_6453);
or U14442 (N_14442,N_7712,N_5539);
nand U14443 (N_14443,N_9928,N_7630);
xnor U14444 (N_14444,N_7021,N_9961);
nand U14445 (N_14445,N_8984,N_7448);
xor U14446 (N_14446,N_5508,N_9977);
or U14447 (N_14447,N_8224,N_6430);
nand U14448 (N_14448,N_7990,N_7387);
nor U14449 (N_14449,N_5285,N_6619);
nor U14450 (N_14450,N_9169,N_7187);
and U14451 (N_14451,N_5754,N_8696);
or U14452 (N_14452,N_5494,N_8727);
or U14453 (N_14453,N_5964,N_5050);
and U14454 (N_14454,N_7657,N_5349);
or U14455 (N_14455,N_6605,N_5849);
nor U14456 (N_14456,N_5189,N_7731);
nor U14457 (N_14457,N_6445,N_5099);
nand U14458 (N_14458,N_9170,N_8661);
xor U14459 (N_14459,N_7672,N_9637);
and U14460 (N_14460,N_5639,N_6722);
and U14461 (N_14461,N_9353,N_5806);
nor U14462 (N_14462,N_8679,N_5941);
nand U14463 (N_14463,N_5600,N_8055);
xnor U14464 (N_14464,N_7672,N_8490);
xnor U14465 (N_14465,N_9773,N_8855);
or U14466 (N_14466,N_6502,N_6119);
and U14467 (N_14467,N_7272,N_5248);
nand U14468 (N_14468,N_5432,N_5956);
and U14469 (N_14469,N_9905,N_7329);
or U14470 (N_14470,N_7289,N_9100);
and U14471 (N_14471,N_8557,N_7107);
nand U14472 (N_14472,N_8184,N_9364);
nor U14473 (N_14473,N_5957,N_5033);
or U14474 (N_14474,N_5436,N_8437);
nand U14475 (N_14475,N_8809,N_8717);
xnor U14476 (N_14476,N_5525,N_8241);
xor U14477 (N_14477,N_7392,N_8722);
nand U14478 (N_14478,N_5341,N_7796);
or U14479 (N_14479,N_8090,N_8522);
and U14480 (N_14480,N_9650,N_9208);
or U14481 (N_14481,N_8460,N_6560);
and U14482 (N_14482,N_5421,N_7465);
nor U14483 (N_14483,N_8131,N_9025);
nor U14484 (N_14484,N_8973,N_6335);
nand U14485 (N_14485,N_7840,N_8123);
xnor U14486 (N_14486,N_7847,N_8465);
nand U14487 (N_14487,N_7326,N_5589);
and U14488 (N_14488,N_5803,N_9798);
nor U14489 (N_14489,N_6287,N_7859);
or U14490 (N_14490,N_8234,N_7375);
nand U14491 (N_14491,N_7002,N_8812);
xor U14492 (N_14492,N_7643,N_8971);
or U14493 (N_14493,N_7013,N_8995);
nor U14494 (N_14494,N_7081,N_6601);
xnor U14495 (N_14495,N_6342,N_6516);
nor U14496 (N_14496,N_8690,N_9762);
nor U14497 (N_14497,N_6492,N_6165);
xnor U14498 (N_14498,N_6651,N_8382);
nand U14499 (N_14499,N_7562,N_7566);
nor U14500 (N_14500,N_8911,N_6543);
nand U14501 (N_14501,N_9016,N_9255);
nand U14502 (N_14502,N_8570,N_7006);
or U14503 (N_14503,N_7772,N_7657);
or U14504 (N_14504,N_9745,N_8369);
nand U14505 (N_14505,N_5179,N_5403);
and U14506 (N_14506,N_7383,N_8324);
nor U14507 (N_14507,N_6737,N_8100);
xor U14508 (N_14508,N_6153,N_5120);
nand U14509 (N_14509,N_7256,N_5366);
and U14510 (N_14510,N_5993,N_7452);
nand U14511 (N_14511,N_9246,N_8511);
or U14512 (N_14512,N_7466,N_8858);
nor U14513 (N_14513,N_6562,N_9238);
xor U14514 (N_14514,N_9847,N_5927);
xnor U14515 (N_14515,N_9841,N_9822);
and U14516 (N_14516,N_6545,N_8881);
xnor U14517 (N_14517,N_9018,N_8555);
xnor U14518 (N_14518,N_8679,N_8019);
nor U14519 (N_14519,N_6840,N_7460);
or U14520 (N_14520,N_8918,N_5875);
and U14521 (N_14521,N_6246,N_5792);
or U14522 (N_14522,N_8469,N_5570);
nand U14523 (N_14523,N_7788,N_9785);
nor U14524 (N_14524,N_6060,N_6563);
xor U14525 (N_14525,N_5069,N_5006);
or U14526 (N_14526,N_5570,N_5982);
nand U14527 (N_14527,N_6047,N_6292);
xor U14528 (N_14528,N_7176,N_6094);
nand U14529 (N_14529,N_7185,N_5896);
nand U14530 (N_14530,N_5075,N_6629);
and U14531 (N_14531,N_9669,N_7777);
nor U14532 (N_14532,N_5513,N_9127);
and U14533 (N_14533,N_6784,N_5469);
or U14534 (N_14534,N_5197,N_5576);
and U14535 (N_14535,N_9071,N_9153);
nor U14536 (N_14536,N_8110,N_6604);
nand U14537 (N_14537,N_8669,N_9795);
nand U14538 (N_14538,N_9875,N_9893);
nor U14539 (N_14539,N_5663,N_8692);
nor U14540 (N_14540,N_5767,N_5619);
nor U14541 (N_14541,N_6050,N_7770);
xnor U14542 (N_14542,N_6367,N_7959);
nor U14543 (N_14543,N_9338,N_6352);
or U14544 (N_14544,N_5019,N_6345);
nor U14545 (N_14545,N_5100,N_7811);
nand U14546 (N_14546,N_8378,N_9757);
and U14547 (N_14547,N_7905,N_8101);
nor U14548 (N_14548,N_8083,N_9401);
or U14549 (N_14549,N_7940,N_5354);
xor U14550 (N_14550,N_5613,N_5299);
nand U14551 (N_14551,N_7943,N_6763);
nor U14552 (N_14552,N_6958,N_7153);
nand U14553 (N_14553,N_8132,N_8265);
xor U14554 (N_14554,N_6221,N_9116);
nand U14555 (N_14555,N_8644,N_5043);
nor U14556 (N_14556,N_6019,N_5294);
and U14557 (N_14557,N_8544,N_9626);
nor U14558 (N_14558,N_6691,N_8248);
and U14559 (N_14559,N_5729,N_8743);
or U14560 (N_14560,N_7066,N_5330);
and U14561 (N_14561,N_8224,N_8322);
nor U14562 (N_14562,N_5758,N_5664);
xnor U14563 (N_14563,N_9233,N_7949);
xnor U14564 (N_14564,N_6388,N_9012);
xor U14565 (N_14565,N_8524,N_6197);
or U14566 (N_14566,N_9602,N_8907);
nor U14567 (N_14567,N_9862,N_9517);
nand U14568 (N_14568,N_9159,N_9214);
nor U14569 (N_14569,N_7447,N_6744);
xor U14570 (N_14570,N_6367,N_9450);
nand U14571 (N_14571,N_6604,N_6616);
nor U14572 (N_14572,N_5477,N_6460);
nand U14573 (N_14573,N_9899,N_6939);
xnor U14574 (N_14574,N_6654,N_8369);
and U14575 (N_14575,N_6808,N_6937);
and U14576 (N_14576,N_9964,N_7543);
nand U14577 (N_14577,N_7106,N_9699);
and U14578 (N_14578,N_8571,N_8725);
xor U14579 (N_14579,N_5770,N_7454);
nor U14580 (N_14580,N_6252,N_6666);
nor U14581 (N_14581,N_7454,N_5431);
and U14582 (N_14582,N_9542,N_7166);
xnor U14583 (N_14583,N_7507,N_6333);
or U14584 (N_14584,N_7588,N_9213);
and U14585 (N_14585,N_6514,N_5258);
xor U14586 (N_14586,N_7981,N_6548);
or U14587 (N_14587,N_6408,N_6919);
and U14588 (N_14588,N_7305,N_5569);
or U14589 (N_14589,N_9149,N_5911);
and U14590 (N_14590,N_7985,N_7048);
xnor U14591 (N_14591,N_6896,N_8981);
or U14592 (N_14592,N_8209,N_5400);
nand U14593 (N_14593,N_6235,N_6923);
nand U14594 (N_14594,N_6620,N_5884);
or U14595 (N_14595,N_5425,N_9503);
and U14596 (N_14596,N_9941,N_7731);
and U14597 (N_14597,N_8326,N_6492);
nor U14598 (N_14598,N_9786,N_5851);
xor U14599 (N_14599,N_6252,N_5188);
xor U14600 (N_14600,N_7173,N_9909);
nand U14601 (N_14601,N_7252,N_5560);
xor U14602 (N_14602,N_8403,N_6891);
xnor U14603 (N_14603,N_8654,N_6235);
xor U14604 (N_14604,N_6443,N_6474);
nand U14605 (N_14605,N_8667,N_5920);
nand U14606 (N_14606,N_8124,N_5116);
xnor U14607 (N_14607,N_9983,N_8379);
or U14608 (N_14608,N_7201,N_9555);
nand U14609 (N_14609,N_9956,N_6489);
and U14610 (N_14610,N_8075,N_5188);
nand U14611 (N_14611,N_9924,N_9776);
nand U14612 (N_14612,N_5219,N_8628);
xnor U14613 (N_14613,N_7193,N_7973);
nor U14614 (N_14614,N_8562,N_5696);
xnor U14615 (N_14615,N_7865,N_5372);
xor U14616 (N_14616,N_6583,N_7181);
xnor U14617 (N_14617,N_5612,N_8135);
nand U14618 (N_14618,N_8471,N_8000);
or U14619 (N_14619,N_6911,N_8450);
nand U14620 (N_14620,N_7592,N_9663);
xnor U14621 (N_14621,N_8455,N_6858);
nor U14622 (N_14622,N_6776,N_5097);
nor U14623 (N_14623,N_6503,N_9677);
xor U14624 (N_14624,N_7334,N_5126);
and U14625 (N_14625,N_9597,N_8460);
nor U14626 (N_14626,N_6856,N_7542);
or U14627 (N_14627,N_7866,N_5579);
nor U14628 (N_14628,N_7992,N_9587);
xnor U14629 (N_14629,N_7587,N_8858);
or U14630 (N_14630,N_6919,N_8651);
and U14631 (N_14631,N_9499,N_8273);
nor U14632 (N_14632,N_6524,N_5460);
and U14633 (N_14633,N_7822,N_6972);
or U14634 (N_14634,N_9289,N_7643);
nor U14635 (N_14635,N_9731,N_8560);
nand U14636 (N_14636,N_9877,N_6111);
xnor U14637 (N_14637,N_6154,N_7213);
xnor U14638 (N_14638,N_9915,N_8353);
nor U14639 (N_14639,N_8539,N_8708);
nor U14640 (N_14640,N_7989,N_6332);
or U14641 (N_14641,N_6858,N_9479);
or U14642 (N_14642,N_9122,N_6573);
nand U14643 (N_14643,N_5697,N_9287);
xnor U14644 (N_14644,N_8432,N_5722);
nor U14645 (N_14645,N_8555,N_9029);
and U14646 (N_14646,N_8132,N_9802);
xnor U14647 (N_14647,N_6003,N_8057);
xor U14648 (N_14648,N_5261,N_8805);
nor U14649 (N_14649,N_8576,N_9574);
or U14650 (N_14650,N_9007,N_6684);
nand U14651 (N_14651,N_7411,N_8950);
nor U14652 (N_14652,N_6635,N_6761);
or U14653 (N_14653,N_7462,N_9565);
nor U14654 (N_14654,N_6667,N_8622);
or U14655 (N_14655,N_6669,N_6397);
and U14656 (N_14656,N_5095,N_6728);
nand U14657 (N_14657,N_7084,N_8769);
nand U14658 (N_14658,N_5514,N_9616);
or U14659 (N_14659,N_6256,N_6306);
and U14660 (N_14660,N_9675,N_6072);
and U14661 (N_14661,N_8383,N_8053);
nor U14662 (N_14662,N_8871,N_9433);
and U14663 (N_14663,N_7544,N_5034);
nand U14664 (N_14664,N_9825,N_7185);
and U14665 (N_14665,N_5675,N_5559);
or U14666 (N_14666,N_9952,N_7277);
nor U14667 (N_14667,N_6348,N_5415);
and U14668 (N_14668,N_5776,N_6349);
and U14669 (N_14669,N_5589,N_5102);
nor U14670 (N_14670,N_7054,N_9767);
nor U14671 (N_14671,N_9331,N_5606);
xor U14672 (N_14672,N_9258,N_6966);
and U14673 (N_14673,N_6658,N_9862);
nand U14674 (N_14674,N_5437,N_5104);
nor U14675 (N_14675,N_9373,N_8175);
nor U14676 (N_14676,N_8574,N_7393);
and U14677 (N_14677,N_7200,N_6308);
or U14678 (N_14678,N_9499,N_6698);
xnor U14679 (N_14679,N_6853,N_7828);
nor U14680 (N_14680,N_6403,N_6593);
nand U14681 (N_14681,N_7755,N_8921);
xor U14682 (N_14682,N_7559,N_6332);
nand U14683 (N_14683,N_8257,N_8926);
nor U14684 (N_14684,N_7133,N_6787);
nand U14685 (N_14685,N_6305,N_8617);
or U14686 (N_14686,N_7216,N_8816);
nand U14687 (N_14687,N_7612,N_9047);
nand U14688 (N_14688,N_7054,N_8772);
nand U14689 (N_14689,N_8170,N_7723);
nand U14690 (N_14690,N_7615,N_7287);
and U14691 (N_14691,N_8770,N_5056);
xor U14692 (N_14692,N_8781,N_5660);
nand U14693 (N_14693,N_9517,N_5788);
or U14694 (N_14694,N_7733,N_9551);
xor U14695 (N_14695,N_9747,N_5718);
or U14696 (N_14696,N_5687,N_6425);
nor U14697 (N_14697,N_7494,N_9275);
and U14698 (N_14698,N_9435,N_5356);
or U14699 (N_14699,N_5219,N_9666);
xor U14700 (N_14700,N_5940,N_6539);
and U14701 (N_14701,N_6570,N_7078);
and U14702 (N_14702,N_6049,N_7995);
nand U14703 (N_14703,N_5433,N_5457);
xnor U14704 (N_14704,N_7547,N_7782);
or U14705 (N_14705,N_5119,N_7363);
xor U14706 (N_14706,N_8505,N_6816);
or U14707 (N_14707,N_8945,N_6693);
xnor U14708 (N_14708,N_9345,N_9330);
xor U14709 (N_14709,N_6185,N_6687);
nor U14710 (N_14710,N_5373,N_6267);
nand U14711 (N_14711,N_6602,N_6926);
or U14712 (N_14712,N_5436,N_5355);
xor U14713 (N_14713,N_7041,N_8132);
xnor U14714 (N_14714,N_7956,N_7998);
nand U14715 (N_14715,N_5729,N_7187);
and U14716 (N_14716,N_9640,N_5696);
and U14717 (N_14717,N_8082,N_6421);
nor U14718 (N_14718,N_6918,N_9384);
nor U14719 (N_14719,N_9280,N_5386);
nor U14720 (N_14720,N_8934,N_6758);
or U14721 (N_14721,N_8426,N_5178);
and U14722 (N_14722,N_6950,N_6473);
xor U14723 (N_14723,N_8010,N_6811);
or U14724 (N_14724,N_6566,N_6863);
or U14725 (N_14725,N_5316,N_6435);
nor U14726 (N_14726,N_5585,N_8182);
nand U14727 (N_14727,N_5175,N_7237);
or U14728 (N_14728,N_9345,N_9130);
and U14729 (N_14729,N_9174,N_5283);
nor U14730 (N_14730,N_5955,N_5627);
xor U14731 (N_14731,N_6989,N_7606);
xor U14732 (N_14732,N_7429,N_8620);
xor U14733 (N_14733,N_6703,N_7316);
and U14734 (N_14734,N_8267,N_8281);
xor U14735 (N_14735,N_5198,N_6564);
nor U14736 (N_14736,N_6708,N_5590);
or U14737 (N_14737,N_9880,N_6415);
nor U14738 (N_14738,N_9967,N_8241);
and U14739 (N_14739,N_7987,N_5648);
nor U14740 (N_14740,N_7397,N_7598);
xor U14741 (N_14741,N_8024,N_8081);
and U14742 (N_14742,N_8408,N_5254);
xnor U14743 (N_14743,N_7324,N_6086);
xor U14744 (N_14744,N_9571,N_6348);
xnor U14745 (N_14745,N_5672,N_7224);
xnor U14746 (N_14746,N_6355,N_8187);
or U14747 (N_14747,N_6627,N_7440);
nor U14748 (N_14748,N_5768,N_8719);
nor U14749 (N_14749,N_5422,N_7790);
nor U14750 (N_14750,N_8513,N_5223);
xor U14751 (N_14751,N_9874,N_8088);
nor U14752 (N_14752,N_5572,N_8367);
or U14753 (N_14753,N_7742,N_7103);
nor U14754 (N_14754,N_8059,N_5507);
xnor U14755 (N_14755,N_8284,N_7486);
nor U14756 (N_14756,N_5327,N_7282);
nand U14757 (N_14757,N_9015,N_9972);
nand U14758 (N_14758,N_7443,N_7728);
nand U14759 (N_14759,N_7102,N_7522);
and U14760 (N_14760,N_5336,N_6583);
xor U14761 (N_14761,N_7205,N_5451);
xnor U14762 (N_14762,N_8407,N_7203);
or U14763 (N_14763,N_5855,N_5107);
and U14764 (N_14764,N_6130,N_8357);
or U14765 (N_14765,N_5603,N_5182);
or U14766 (N_14766,N_5560,N_7486);
and U14767 (N_14767,N_6889,N_5557);
or U14768 (N_14768,N_6412,N_5905);
xnor U14769 (N_14769,N_5974,N_9191);
xnor U14770 (N_14770,N_6464,N_5320);
or U14771 (N_14771,N_7504,N_8684);
xor U14772 (N_14772,N_6075,N_9101);
xnor U14773 (N_14773,N_5874,N_5486);
xnor U14774 (N_14774,N_9745,N_6624);
nand U14775 (N_14775,N_6493,N_7275);
nor U14776 (N_14776,N_7583,N_9338);
and U14777 (N_14777,N_8649,N_9762);
xnor U14778 (N_14778,N_5459,N_8054);
xor U14779 (N_14779,N_9685,N_8211);
and U14780 (N_14780,N_9015,N_7962);
or U14781 (N_14781,N_5850,N_7918);
or U14782 (N_14782,N_5820,N_5244);
or U14783 (N_14783,N_9079,N_6067);
nor U14784 (N_14784,N_5559,N_5047);
and U14785 (N_14785,N_6705,N_5601);
and U14786 (N_14786,N_9280,N_5779);
and U14787 (N_14787,N_7901,N_9820);
xnor U14788 (N_14788,N_5199,N_9090);
nand U14789 (N_14789,N_6241,N_9515);
nand U14790 (N_14790,N_5885,N_7419);
xnor U14791 (N_14791,N_7933,N_6544);
or U14792 (N_14792,N_8812,N_7293);
or U14793 (N_14793,N_7358,N_8674);
and U14794 (N_14794,N_5908,N_6150);
and U14795 (N_14795,N_8929,N_7665);
or U14796 (N_14796,N_6807,N_8315);
or U14797 (N_14797,N_6600,N_5925);
and U14798 (N_14798,N_9699,N_9604);
nand U14799 (N_14799,N_8624,N_9635);
or U14800 (N_14800,N_8403,N_9048);
nand U14801 (N_14801,N_8957,N_9019);
xor U14802 (N_14802,N_7816,N_9359);
xnor U14803 (N_14803,N_6885,N_6697);
nand U14804 (N_14804,N_7653,N_7963);
xnor U14805 (N_14805,N_8050,N_5498);
nor U14806 (N_14806,N_9558,N_9639);
nand U14807 (N_14807,N_7847,N_9599);
nor U14808 (N_14808,N_5645,N_7922);
and U14809 (N_14809,N_7013,N_6162);
nand U14810 (N_14810,N_8803,N_5631);
nand U14811 (N_14811,N_7659,N_7592);
nand U14812 (N_14812,N_6891,N_6220);
nor U14813 (N_14813,N_5431,N_5053);
xor U14814 (N_14814,N_9012,N_6566);
or U14815 (N_14815,N_6666,N_6047);
xnor U14816 (N_14816,N_8312,N_7058);
xor U14817 (N_14817,N_5024,N_7845);
nor U14818 (N_14818,N_8357,N_6204);
or U14819 (N_14819,N_9408,N_5093);
xor U14820 (N_14820,N_9311,N_7556);
nor U14821 (N_14821,N_6823,N_9562);
nand U14822 (N_14822,N_7585,N_5880);
nor U14823 (N_14823,N_6458,N_8649);
nor U14824 (N_14824,N_5875,N_8794);
or U14825 (N_14825,N_5126,N_5152);
or U14826 (N_14826,N_9672,N_6316);
nand U14827 (N_14827,N_7270,N_8693);
nor U14828 (N_14828,N_5675,N_9174);
nor U14829 (N_14829,N_6031,N_9528);
xnor U14830 (N_14830,N_8786,N_7288);
nand U14831 (N_14831,N_9822,N_7292);
nand U14832 (N_14832,N_9600,N_9131);
or U14833 (N_14833,N_8950,N_7414);
or U14834 (N_14834,N_7427,N_9232);
nand U14835 (N_14835,N_8236,N_8686);
nand U14836 (N_14836,N_9155,N_9073);
xnor U14837 (N_14837,N_7993,N_5697);
nor U14838 (N_14838,N_9606,N_8762);
nand U14839 (N_14839,N_8530,N_9113);
or U14840 (N_14840,N_8913,N_7199);
or U14841 (N_14841,N_8335,N_5199);
xor U14842 (N_14842,N_8361,N_7924);
nor U14843 (N_14843,N_6826,N_5628);
nor U14844 (N_14844,N_7682,N_9753);
nor U14845 (N_14845,N_7363,N_6925);
nor U14846 (N_14846,N_6427,N_6403);
nand U14847 (N_14847,N_7020,N_8894);
or U14848 (N_14848,N_6057,N_5129);
or U14849 (N_14849,N_7116,N_7256);
xor U14850 (N_14850,N_8548,N_6085);
or U14851 (N_14851,N_5567,N_6476);
and U14852 (N_14852,N_5188,N_5523);
nand U14853 (N_14853,N_6330,N_5268);
xnor U14854 (N_14854,N_8976,N_9015);
nor U14855 (N_14855,N_8558,N_7599);
and U14856 (N_14856,N_9420,N_5154);
xnor U14857 (N_14857,N_9143,N_9247);
and U14858 (N_14858,N_6296,N_6835);
xor U14859 (N_14859,N_5553,N_8927);
xor U14860 (N_14860,N_9183,N_9886);
nor U14861 (N_14861,N_8212,N_6281);
xor U14862 (N_14862,N_8846,N_6443);
or U14863 (N_14863,N_9942,N_5697);
or U14864 (N_14864,N_9687,N_5635);
or U14865 (N_14865,N_7995,N_7984);
nor U14866 (N_14866,N_5923,N_6559);
and U14867 (N_14867,N_7797,N_7649);
and U14868 (N_14868,N_8402,N_7849);
xnor U14869 (N_14869,N_9378,N_5616);
xor U14870 (N_14870,N_8107,N_7199);
nand U14871 (N_14871,N_5763,N_9885);
or U14872 (N_14872,N_6793,N_6837);
xor U14873 (N_14873,N_7216,N_6412);
nand U14874 (N_14874,N_5476,N_5042);
and U14875 (N_14875,N_5473,N_7179);
or U14876 (N_14876,N_9027,N_7840);
and U14877 (N_14877,N_8872,N_9555);
and U14878 (N_14878,N_8180,N_9317);
or U14879 (N_14879,N_8322,N_6146);
nor U14880 (N_14880,N_7926,N_9136);
nor U14881 (N_14881,N_7100,N_6282);
and U14882 (N_14882,N_7079,N_7177);
or U14883 (N_14883,N_9365,N_8575);
nand U14884 (N_14884,N_6108,N_9276);
nand U14885 (N_14885,N_5997,N_7214);
and U14886 (N_14886,N_8693,N_8996);
nor U14887 (N_14887,N_9400,N_5300);
xnor U14888 (N_14888,N_5260,N_8035);
and U14889 (N_14889,N_5810,N_7828);
nand U14890 (N_14890,N_7944,N_7340);
or U14891 (N_14891,N_5304,N_6124);
xor U14892 (N_14892,N_6110,N_6580);
xor U14893 (N_14893,N_9932,N_7219);
xor U14894 (N_14894,N_5684,N_9760);
xnor U14895 (N_14895,N_9113,N_9472);
nor U14896 (N_14896,N_7680,N_8651);
xor U14897 (N_14897,N_8949,N_7911);
nor U14898 (N_14898,N_7418,N_8274);
or U14899 (N_14899,N_8865,N_6289);
nand U14900 (N_14900,N_6999,N_7039);
nor U14901 (N_14901,N_6568,N_7237);
xnor U14902 (N_14902,N_6863,N_9675);
or U14903 (N_14903,N_8091,N_8953);
nor U14904 (N_14904,N_6035,N_9918);
nand U14905 (N_14905,N_6206,N_8672);
nor U14906 (N_14906,N_7156,N_8291);
xor U14907 (N_14907,N_7859,N_6851);
nand U14908 (N_14908,N_6705,N_9605);
nand U14909 (N_14909,N_9220,N_5103);
xnor U14910 (N_14910,N_7581,N_7419);
or U14911 (N_14911,N_5870,N_7739);
nor U14912 (N_14912,N_7252,N_5889);
and U14913 (N_14913,N_5836,N_8612);
or U14914 (N_14914,N_9486,N_7986);
nor U14915 (N_14915,N_7627,N_8039);
xor U14916 (N_14916,N_7007,N_9469);
nor U14917 (N_14917,N_6618,N_5997);
or U14918 (N_14918,N_9678,N_6135);
or U14919 (N_14919,N_9782,N_8896);
xor U14920 (N_14920,N_9121,N_8326);
and U14921 (N_14921,N_8785,N_7850);
xnor U14922 (N_14922,N_6696,N_5745);
or U14923 (N_14923,N_7281,N_6253);
nor U14924 (N_14924,N_5672,N_5492);
xor U14925 (N_14925,N_7289,N_6306);
or U14926 (N_14926,N_9587,N_5610);
or U14927 (N_14927,N_6083,N_8505);
and U14928 (N_14928,N_5417,N_7727);
nand U14929 (N_14929,N_9762,N_9634);
and U14930 (N_14930,N_6796,N_6857);
xor U14931 (N_14931,N_8331,N_5395);
or U14932 (N_14932,N_6756,N_7448);
or U14933 (N_14933,N_8504,N_6087);
or U14934 (N_14934,N_7423,N_9546);
and U14935 (N_14935,N_8891,N_9791);
xnor U14936 (N_14936,N_8532,N_6963);
nand U14937 (N_14937,N_5834,N_7350);
xor U14938 (N_14938,N_9593,N_8914);
or U14939 (N_14939,N_8746,N_6720);
nand U14940 (N_14940,N_5201,N_8188);
nand U14941 (N_14941,N_5500,N_8182);
nand U14942 (N_14942,N_7193,N_9244);
nand U14943 (N_14943,N_9082,N_5561);
nor U14944 (N_14944,N_9872,N_8772);
and U14945 (N_14945,N_7667,N_5699);
nor U14946 (N_14946,N_9070,N_6057);
or U14947 (N_14947,N_9066,N_8838);
nor U14948 (N_14948,N_7304,N_5306);
and U14949 (N_14949,N_8391,N_5951);
or U14950 (N_14950,N_7098,N_7052);
xnor U14951 (N_14951,N_8178,N_9359);
xor U14952 (N_14952,N_5106,N_6028);
or U14953 (N_14953,N_7500,N_9682);
nor U14954 (N_14954,N_8010,N_9008);
nor U14955 (N_14955,N_8127,N_9123);
and U14956 (N_14956,N_5594,N_9837);
nor U14957 (N_14957,N_7233,N_7530);
or U14958 (N_14958,N_7546,N_8566);
and U14959 (N_14959,N_8381,N_9239);
nor U14960 (N_14960,N_9932,N_9957);
or U14961 (N_14961,N_8818,N_6729);
nor U14962 (N_14962,N_5940,N_7478);
and U14963 (N_14963,N_6898,N_7735);
or U14964 (N_14964,N_6608,N_8804);
or U14965 (N_14965,N_9268,N_5906);
and U14966 (N_14966,N_5565,N_8238);
nand U14967 (N_14967,N_6833,N_8464);
nor U14968 (N_14968,N_7610,N_6432);
xnor U14969 (N_14969,N_8645,N_9306);
nor U14970 (N_14970,N_9539,N_8892);
and U14971 (N_14971,N_6100,N_7806);
nand U14972 (N_14972,N_8170,N_5222);
nand U14973 (N_14973,N_7835,N_5944);
nor U14974 (N_14974,N_7107,N_8611);
xor U14975 (N_14975,N_6381,N_6355);
xnor U14976 (N_14976,N_8036,N_7487);
nand U14977 (N_14977,N_6566,N_6358);
or U14978 (N_14978,N_7238,N_5750);
nand U14979 (N_14979,N_8179,N_8429);
xor U14980 (N_14980,N_6680,N_5032);
nor U14981 (N_14981,N_9355,N_8512);
and U14982 (N_14982,N_9161,N_8047);
or U14983 (N_14983,N_9628,N_9407);
and U14984 (N_14984,N_8390,N_6124);
xnor U14985 (N_14985,N_8923,N_8809);
nor U14986 (N_14986,N_5772,N_9113);
and U14987 (N_14987,N_5188,N_5722);
and U14988 (N_14988,N_6469,N_6875);
nand U14989 (N_14989,N_6820,N_7582);
and U14990 (N_14990,N_8632,N_7138);
nand U14991 (N_14991,N_8991,N_9101);
nand U14992 (N_14992,N_9860,N_6804);
and U14993 (N_14993,N_9572,N_9644);
or U14994 (N_14994,N_7426,N_8690);
or U14995 (N_14995,N_9294,N_5259);
xor U14996 (N_14996,N_6987,N_6970);
xor U14997 (N_14997,N_5085,N_5799);
xor U14998 (N_14998,N_9674,N_5570);
and U14999 (N_14999,N_6268,N_6191);
and U15000 (N_15000,N_10502,N_13350);
and U15001 (N_15001,N_10433,N_10994);
xnor U15002 (N_15002,N_10827,N_13337);
or U15003 (N_15003,N_14340,N_12674);
and U15004 (N_15004,N_13671,N_11114);
nor U15005 (N_15005,N_11362,N_11562);
xnor U15006 (N_15006,N_14830,N_10438);
xnor U15007 (N_15007,N_13156,N_12590);
xor U15008 (N_15008,N_12748,N_13652);
xor U15009 (N_15009,N_13631,N_14226);
nand U15010 (N_15010,N_13401,N_11402);
and U15011 (N_15011,N_10245,N_11128);
or U15012 (N_15012,N_14642,N_12872);
nand U15013 (N_15013,N_10058,N_12751);
nor U15014 (N_15014,N_13324,N_14635);
or U15015 (N_15015,N_14441,N_13625);
or U15016 (N_15016,N_12167,N_11747);
or U15017 (N_15017,N_11609,N_11111);
and U15018 (N_15018,N_12449,N_13693);
and U15019 (N_15019,N_10603,N_10895);
xnor U15020 (N_15020,N_12883,N_10369);
xor U15021 (N_15021,N_10723,N_10393);
and U15022 (N_15022,N_13835,N_14159);
or U15023 (N_15023,N_10992,N_14557);
and U15024 (N_15024,N_12684,N_11031);
or U15025 (N_15025,N_14383,N_14227);
or U15026 (N_15026,N_14810,N_14558);
xor U15027 (N_15027,N_10932,N_13511);
and U15028 (N_15028,N_12757,N_11168);
or U15029 (N_15029,N_10066,N_13753);
xor U15030 (N_15030,N_12252,N_10922);
nor U15031 (N_15031,N_11729,N_12814);
nand U15032 (N_15032,N_10456,N_10589);
and U15033 (N_15033,N_12375,N_14670);
xor U15034 (N_15034,N_11869,N_13115);
xnor U15035 (N_15035,N_14724,N_13894);
xor U15036 (N_15036,N_13119,N_12950);
nand U15037 (N_15037,N_11406,N_14435);
nor U15038 (N_15038,N_13045,N_13615);
or U15039 (N_15039,N_11877,N_11893);
xor U15040 (N_15040,N_12810,N_14440);
nand U15041 (N_15041,N_14154,N_10725);
nor U15042 (N_15042,N_13692,N_10270);
nand U15043 (N_15043,N_14399,N_10694);
and U15044 (N_15044,N_14068,N_14965);
and U15045 (N_15045,N_12229,N_12924);
xor U15046 (N_15046,N_11834,N_11004);
nor U15047 (N_15047,N_11595,N_12691);
xnor U15048 (N_15048,N_10790,N_12463);
nor U15049 (N_15049,N_11918,N_12288);
or U15050 (N_15050,N_10791,N_10681);
or U15051 (N_15051,N_12609,N_13140);
xor U15052 (N_15052,N_13378,N_10033);
or U15053 (N_15053,N_13367,N_13272);
xor U15054 (N_15054,N_10864,N_10943);
nand U15055 (N_15055,N_13138,N_10746);
and U15056 (N_15056,N_14752,N_14938);
or U15057 (N_15057,N_11571,N_14732);
or U15058 (N_15058,N_10722,N_10689);
nor U15059 (N_15059,N_14939,N_12307);
nor U15060 (N_15060,N_11758,N_12969);
and U15061 (N_15061,N_12854,N_14375);
nor U15062 (N_15062,N_14048,N_13175);
and U15063 (N_15063,N_12379,N_12442);
or U15064 (N_15064,N_12276,N_10670);
nand U15065 (N_15065,N_12516,N_11070);
and U15066 (N_15066,N_11140,N_14082);
xnor U15067 (N_15067,N_11134,N_12006);
nor U15068 (N_15068,N_12890,N_13764);
nor U15069 (N_15069,N_14478,N_10903);
nand U15070 (N_15070,N_12411,N_10545);
xor U15071 (N_15071,N_11984,N_10053);
xnor U15072 (N_15072,N_12472,N_11813);
xnor U15073 (N_15073,N_11645,N_14660);
and U15074 (N_15074,N_14023,N_13650);
nand U15075 (N_15075,N_13078,N_13912);
and U15076 (N_15076,N_10985,N_12283);
nor U15077 (N_15077,N_11244,N_11184);
nand U15078 (N_15078,N_14964,N_13204);
xor U15079 (N_15079,N_10902,N_12504);
and U15080 (N_15080,N_13900,N_12237);
or U15081 (N_15081,N_10726,N_14090);
xnor U15082 (N_15082,N_10044,N_10884);
or U15083 (N_15083,N_10473,N_13387);
and U15084 (N_15084,N_10976,N_11042);
or U15085 (N_15085,N_11584,N_13022);
or U15086 (N_15086,N_14827,N_14006);
and U15087 (N_15087,N_14518,N_12700);
nor U15088 (N_15088,N_11471,N_11724);
and U15089 (N_15089,N_14208,N_13634);
and U15090 (N_15090,N_11920,N_12423);
and U15091 (N_15091,N_11195,N_13209);
and U15092 (N_15092,N_10754,N_11662);
nor U15093 (N_15093,N_13215,N_14760);
or U15094 (N_15094,N_14743,N_13741);
nor U15095 (N_15095,N_10811,N_10182);
nand U15096 (N_15096,N_12913,N_12736);
nor U15097 (N_15097,N_12014,N_10751);
and U15098 (N_15098,N_13677,N_13609);
and U15099 (N_15099,N_13114,N_14057);
nand U15100 (N_15100,N_10516,N_10996);
nor U15101 (N_15101,N_12117,N_14326);
or U15102 (N_15102,N_13702,N_10036);
xor U15103 (N_15103,N_12210,N_13549);
and U15104 (N_15104,N_12944,N_10767);
and U15105 (N_15105,N_14607,N_13039);
nor U15106 (N_15106,N_13815,N_10301);
and U15107 (N_15107,N_10259,N_13133);
and U15108 (N_15108,N_13909,N_14354);
xnor U15109 (N_15109,N_12614,N_11702);
and U15110 (N_15110,N_14843,N_12498);
and U15111 (N_15111,N_14776,N_14346);
or U15112 (N_15112,N_14749,N_11993);
xnor U15113 (N_15113,N_11247,N_10410);
and U15114 (N_15114,N_10623,N_10257);
and U15115 (N_15115,N_14894,N_12205);
or U15116 (N_15116,N_14608,N_10345);
nor U15117 (N_15117,N_12137,N_10839);
nor U15118 (N_15118,N_12085,N_10304);
xor U15119 (N_15119,N_14523,N_12079);
xor U15120 (N_15120,N_13176,N_10511);
nor U15121 (N_15121,N_10376,N_12104);
nand U15122 (N_15122,N_11684,N_11650);
and U15123 (N_15123,N_12999,N_11257);
and U15124 (N_15124,N_10163,N_11916);
nor U15125 (N_15125,N_10834,N_10889);
and U15126 (N_15126,N_13059,N_14519);
xnor U15127 (N_15127,N_13755,N_10606);
and U15128 (N_15128,N_13129,N_10750);
nand U15129 (N_15129,N_11826,N_14682);
nor U15130 (N_15130,N_14838,N_12032);
nand U15131 (N_15131,N_12733,N_10558);
and U15132 (N_15132,N_13493,N_10665);
xnor U15133 (N_15133,N_14224,N_14053);
nor U15134 (N_15134,N_13206,N_14485);
and U15135 (N_15135,N_13787,N_12653);
nand U15136 (N_15136,N_11763,N_14066);
xor U15137 (N_15137,N_13203,N_13111);
xor U15138 (N_15138,N_14344,N_12677);
nand U15139 (N_15139,N_12529,N_14751);
xor U15140 (N_15140,N_11485,N_14305);
or U15141 (N_15141,N_12439,N_10367);
or U15142 (N_15142,N_11632,N_14113);
nand U15143 (N_15143,N_11078,N_10200);
nor U15144 (N_15144,N_14954,N_12535);
xnor U15145 (N_15145,N_14417,N_12289);
nor U15146 (N_15146,N_11517,N_12774);
or U15147 (N_15147,N_13485,N_13807);
or U15148 (N_15148,N_11976,N_13273);
xnor U15149 (N_15149,N_12465,N_10557);
and U15150 (N_15150,N_12941,N_11617);
and U15151 (N_15151,N_13211,N_12040);
or U15152 (N_15152,N_11428,N_10318);
xor U15153 (N_15153,N_11383,N_11855);
nor U15154 (N_15154,N_13369,N_10408);
and U15155 (N_15155,N_14299,N_10204);
xor U15156 (N_15156,N_11413,N_10073);
and U15157 (N_15157,N_12355,N_13905);
nor U15158 (N_15158,N_12042,N_10832);
and U15159 (N_15159,N_10439,N_12448);
or U15160 (N_15160,N_10296,N_12022);
and U15161 (N_15161,N_10309,N_12324);
xnor U15162 (N_15162,N_14033,N_13380);
or U15163 (N_15163,N_10003,N_10009);
or U15164 (N_15164,N_10535,N_12271);
or U15165 (N_15165,N_10607,N_14505);
or U15166 (N_15166,N_12063,N_11147);
and U15167 (N_15167,N_10045,N_10714);
nand U15168 (N_15168,N_13656,N_14579);
nor U15169 (N_15169,N_10372,N_12335);
xor U15170 (N_15170,N_13540,N_11012);
nand U15171 (N_15171,N_13551,N_11232);
xor U15172 (N_15172,N_10274,N_14825);
nor U15173 (N_15173,N_14698,N_10674);
and U15174 (N_15174,N_12018,N_14144);
nand U15175 (N_15175,N_11896,N_14168);
nor U15176 (N_15176,N_13995,N_10704);
and U15177 (N_15177,N_12038,N_11935);
and U15178 (N_15178,N_14194,N_10284);
or U15179 (N_15179,N_13978,N_10398);
nand U15180 (N_15180,N_10043,N_14389);
and U15181 (N_15181,N_14055,N_14906);
xnor U15182 (N_15182,N_12513,N_14611);
or U15183 (N_15183,N_10685,N_11167);
or U15184 (N_15184,N_13112,N_14193);
and U15185 (N_15185,N_12719,N_11782);
nor U15186 (N_15186,N_10119,N_13240);
or U15187 (N_15187,N_12139,N_14216);
nor U15188 (N_15188,N_10786,N_12203);
or U15189 (N_15189,N_11882,N_10350);
or U15190 (N_15190,N_14653,N_14811);
and U15191 (N_15191,N_12783,N_11902);
or U15192 (N_15192,N_12727,N_12239);
nand U15193 (N_15193,N_10952,N_10621);
or U15194 (N_15194,N_10476,N_13033);
xnor U15195 (N_15195,N_10961,N_14912);
nor U15196 (N_15196,N_10165,N_10818);
nand U15197 (N_15197,N_13734,N_11020);
xnor U15198 (N_15198,N_10243,N_10303);
nor U15199 (N_15199,N_13896,N_14177);
nand U15200 (N_15200,N_14323,N_14260);
nand U15201 (N_15201,N_13405,N_10383);
or U15202 (N_15202,N_12746,N_14133);
nand U15203 (N_15203,N_12300,N_11898);
nor U15204 (N_15204,N_13824,N_11526);
and U15205 (N_15205,N_14669,N_11041);
or U15206 (N_15206,N_13883,N_11365);
and U15207 (N_15207,N_10890,N_14275);
nand U15208 (N_15208,N_12604,N_13015);
nand U15209 (N_15209,N_13368,N_10297);
or U15210 (N_15210,N_11460,N_14138);
nor U15211 (N_15211,N_13803,N_10211);
and U15212 (N_15212,N_10155,N_14387);
or U15213 (N_15213,N_13359,N_13305);
xor U15214 (N_15214,N_13520,N_12739);
xnor U15215 (N_15215,N_11330,N_11243);
xor U15216 (N_15216,N_10249,N_12019);
xor U15217 (N_15217,N_13960,N_12780);
nand U15218 (N_15218,N_10615,N_12051);
and U15219 (N_15219,N_10339,N_10300);
xnor U15220 (N_15220,N_12563,N_12671);
xor U15221 (N_15221,N_14726,N_13688);
xnor U15222 (N_15222,N_12346,N_11603);
xnor U15223 (N_15223,N_12470,N_13619);
nor U15224 (N_15224,N_14393,N_12192);
nand U15225 (N_15225,N_12928,N_10935);
and U15226 (N_15226,N_10748,N_14991);
nand U15227 (N_15227,N_12392,N_10507);
or U15228 (N_15228,N_14277,N_12220);
nor U15229 (N_15229,N_11141,N_10595);
or U15230 (N_15230,N_12143,N_10328);
and U15231 (N_15231,N_12997,N_12860);
or U15232 (N_15232,N_14334,N_10065);
and U15233 (N_15233,N_12973,N_12793);
xnor U15234 (N_15234,N_10776,N_13184);
or U15235 (N_15235,N_10133,N_10466);
xnor U15236 (N_15236,N_10288,N_14846);
nor U15237 (N_15237,N_14714,N_13366);
nand U15238 (N_15238,N_11072,N_14818);
nand U15239 (N_15239,N_14034,N_14832);
nand U15240 (N_15240,N_12459,N_10930);
or U15241 (N_15241,N_12919,N_13210);
and U15242 (N_15242,N_12618,N_14099);
xor U15243 (N_15243,N_10015,N_14378);
xnor U15244 (N_15244,N_13729,N_11319);
nor U15245 (N_15245,N_12873,N_14444);
or U15246 (N_15246,N_11313,N_11207);
nand U15247 (N_15247,N_14515,N_13443);
xnor U15248 (N_15248,N_10458,N_14243);
or U15249 (N_15249,N_11862,N_11710);
nand U15250 (N_15250,N_12643,N_12017);
xnor U15251 (N_15251,N_12937,N_10272);
or U15252 (N_15252,N_12495,N_13792);
nand U15253 (N_15253,N_12194,N_12331);
xnor U15254 (N_15254,N_13416,N_11727);
and U15255 (N_15255,N_12053,N_14329);
or U15256 (N_15256,N_10882,N_11488);
xnor U15257 (N_15257,N_13576,N_10465);
nor U15258 (N_15258,N_13126,N_14000);
xnor U15259 (N_15259,N_10397,N_11371);
nand U15260 (N_15260,N_12790,N_12650);
nand U15261 (N_15261,N_12743,N_14974);
nand U15262 (N_15262,N_13881,N_11624);
xnor U15263 (N_15263,N_11473,N_14943);
and U15264 (N_15264,N_11891,N_14336);
or U15265 (N_15265,N_12845,N_14876);
xor U15266 (N_15266,N_12875,N_14641);
and U15267 (N_15267,N_11796,N_14308);
nand U15268 (N_15268,N_10757,N_11556);
xnor U15269 (N_15269,N_12371,N_10377);
or U15270 (N_15270,N_12593,N_14929);
nor U15271 (N_15271,N_11574,N_11146);
xor U15272 (N_15272,N_13424,N_13944);
nor U15273 (N_15273,N_13445,N_10821);
nor U15274 (N_15274,N_12382,N_14552);
xor U15275 (N_15275,N_13591,N_13635);
xor U15276 (N_15276,N_13128,N_14459);
and U15277 (N_15277,N_11079,N_12804);
nor U15278 (N_15278,N_13708,N_10753);
or U15279 (N_15279,N_13021,N_14274);
nor U15280 (N_15280,N_13185,N_13202);
and U15281 (N_15281,N_11331,N_11676);
nor U15282 (N_15282,N_14950,N_14796);
nor U15283 (N_15283,N_14266,N_11956);
or U15284 (N_15284,N_14145,N_10205);
nor U15285 (N_15285,N_13774,N_11176);
and U15286 (N_15286,N_14903,N_13229);
nand U15287 (N_15287,N_12044,N_10368);
nand U15288 (N_15288,N_10203,N_10760);
and U15289 (N_15289,N_14699,N_12909);
nor U15290 (N_15290,N_14426,N_10178);
nand U15291 (N_15291,N_12791,N_14486);
nand U15292 (N_15292,N_11316,N_12138);
or U15293 (N_15293,N_10349,N_11550);
nand U15294 (N_15294,N_10954,N_12679);
and U15295 (N_15295,N_11756,N_13618);
or U15296 (N_15296,N_13054,N_14317);
nor U15297 (N_15297,N_14960,N_10072);
nor U15298 (N_15298,N_14195,N_12939);
or U15299 (N_15299,N_14215,N_10405);
nand U15300 (N_15300,N_13189,N_11116);
nand U15301 (N_15301,N_13053,N_10820);
nor U15302 (N_15302,N_11503,N_11281);
or U15303 (N_15303,N_13519,N_13796);
and U15304 (N_15304,N_14210,N_14065);
nand U15305 (N_15305,N_10384,N_13010);
or U15306 (N_15306,N_12446,N_14001);
nor U15307 (N_15307,N_13194,N_14504);
nor U15308 (N_15308,N_10306,N_12620);
nor U15309 (N_15309,N_11117,N_10088);
and U15310 (N_15310,N_14596,N_10712);
xor U15311 (N_15311,N_12586,N_11478);
and U15312 (N_15312,N_12067,N_12078);
nor U15313 (N_15313,N_13178,N_10641);
nor U15314 (N_15314,N_14905,N_14119);
xor U15315 (N_15315,N_12430,N_12594);
nand U15316 (N_15316,N_13550,N_10179);
or U15317 (N_15317,N_12011,N_12437);
and U15318 (N_15318,N_13349,N_11443);
nor U15319 (N_15319,N_10892,N_14135);
xor U15320 (N_15320,N_13085,N_14118);
nor U15321 (N_15321,N_14438,N_12365);
nor U15322 (N_15322,N_11021,N_10069);
and U15323 (N_15323,N_10220,N_13426);
nor U15324 (N_15324,N_14487,N_14924);
and U15325 (N_15325,N_13235,N_12405);
xor U15326 (N_15326,N_14716,N_13145);
nor U15327 (N_15327,N_12369,N_12977);
xnor U15328 (N_15328,N_12359,N_13725);
xor U15329 (N_15329,N_14044,N_12092);
or U15330 (N_15330,N_11329,N_12427);
nor U15331 (N_15331,N_13707,N_11071);
or U15332 (N_15332,N_12047,N_13208);
nand U15333 (N_15333,N_10140,N_13398);
and U15334 (N_15334,N_12701,N_12926);
nand U15335 (N_15335,N_13122,N_14311);
or U15336 (N_15336,N_14396,N_13422);
nor U15337 (N_15337,N_11044,N_13850);
nor U15338 (N_15338,N_12234,N_10057);
xor U15339 (N_15339,N_11604,N_11265);
nor U15340 (N_15340,N_14946,N_12110);
nor U15341 (N_15341,N_13105,N_11465);
xnor U15342 (N_15342,N_12056,N_12169);
and U15343 (N_15343,N_10455,N_12059);
or U15344 (N_15344,N_11880,N_14802);
nor U15345 (N_15345,N_11267,N_14182);
or U15346 (N_15346,N_14548,N_10565);
xor U15347 (N_15347,N_12720,N_10646);
nand U15348 (N_15348,N_12407,N_14136);
nand U15349 (N_15349,N_14790,N_11721);
nand U15350 (N_15350,N_13641,N_10861);
and U15351 (N_15351,N_10653,N_12779);
xor U15352 (N_15352,N_14879,N_10187);
and U15353 (N_15353,N_12471,N_10267);
or U15354 (N_15354,N_12799,N_14294);
xnor U15355 (N_15355,N_14728,N_14453);
nand U15356 (N_15356,N_11082,N_14298);
nor U15357 (N_15357,N_11714,N_12238);
or U15358 (N_15358,N_14956,N_12180);
nand U15359 (N_15359,N_14497,N_11932);
or U15360 (N_15360,N_14106,N_13512);
nand U15361 (N_15361,N_10871,N_11785);
and U15362 (N_15362,N_10823,N_10109);
nand U15363 (N_15363,N_11236,N_14436);
xnor U15364 (N_15364,N_10115,N_11717);
and U15365 (N_15365,N_14831,N_11974);
xor U15366 (N_15366,N_13680,N_12281);
nor U15367 (N_15367,N_12605,N_13452);
xor U15368 (N_15368,N_13507,N_13775);
and U15369 (N_15369,N_11551,N_12897);
xnor U15370 (N_15370,N_14447,N_14073);
and U15371 (N_15371,N_13567,N_10276);
xnor U15372 (N_15372,N_10809,N_12415);
nand U15373 (N_15373,N_14615,N_10000);
nor U15374 (N_15374,N_13454,N_11618);
xor U15375 (N_15375,N_12633,N_13274);
or U15376 (N_15376,N_12390,N_10807);
nand U15377 (N_15377,N_14165,N_14704);
or U15378 (N_15378,N_10008,N_13417);
nand U15379 (N_15379,N_11969,N_10797);
xnor U15380 (N_15380,N_10112,N_12333);
nor U15381 (N_15381,N_11892,N_10246);
nand U15382 (N_15382,N_13862,N_13546);
and U15383 (N_15383,N_10358,N_10352);
or U15384 (N_15384,N_14061,N_12921);
nor U15385 (N_15385,N_13303,N_10283);
xnor U15386 (N_15386,N_10958,N_10873);
nand U15387 (N_15387,N_14403,N_12468);
and U15388 (N_15388,N_12023,N_13298);
and U15389 (N_15389,N_10857,N_10979);
or U15390 (N_15390,N_13199,N_11288);
nor U15391 (N_15391,N_12957,N_14619);
nor U15392 (N_15392,N_11991,N_11800);
and U15393 (N_15393,N_13221,N_11028);
nor U15394 (N_15394,N_14640,N_14139);
nor U15395 (N_15395,N_14588,N_12069);
nand U15396 (N_15396,N_10196,N_13795);
nor U15397 (N_15397,N_14744,N_13327);
xnor U15398 (N_15398,N_11143,N_10080);
nand U15399 (N_15399,N_12822,N_10153);
and U15400 (N_15400,N_10830,N_13365);
and U15401 (N_15401,N_10527,N_14576);
or U15402 (N_15402,N_10879,N_12843);
nor U15403 (N_15403,N_11376,N_10174);
xnor U15404 (N_15404,N_12091,N_11469);
nand U15405 (N_15405,N_14002,N_14780);
and U15406 (N_15406,N_14499,N_14148);
nand U15407 (N_15407,N_10425,N_13694);
nand U15408 (N_15408,N_14856,N_12140);
and U15409 (N_15409,N_10340,N_13379);
and U15410 (N_15410,N_12106,N_11711);
nor U15411 (N_15411,N_13790,N_12596);
nor U15412 (N_15412,N_14069,N_12721);
nand U15413 (N_15413,N_13034,N_12217);
and U15414 (N_15414,N_13411,N_13435);
and U15415 (N_15415,N_12482,N_12813);
or U15416 (N_15416,N_14854,N_12664);
or U15417 (N_15417,N_11718,N_12298);
nand U15418 (N_15418,N_14872,N_14857);
and U15419 (N_15419,N_12157,N_12545);
or U15420 (N_15420,N_13318,N_11080);
and U15421 (N_15421,N_11516,N_11568);
or U15422 (N_15422,N_10039,N_12826);
and U15423 (N_15423,N_11001,N_11417);
nand U15424 (N_15424,N_14004,N_13330);
xnor U15425 (N_15425,N_12877,N_14821);
and U15426 (N_15426,N_14968,N_12703);
nor U15427 (N_15427,N_10856,N_14031);
nand U15428 (N_15428,N_12174,N_14997);
nor U15429 (N_15429,N_10012,N_12555);
or U15430 (N_15430,N_13354,N_11672);
or U15431 (N_15431,N_10237,N_11981);
xor U15432 (N_15432,N_11347,N_10103);
nand U15433 (N_15433,N_12863,N_10035);
nand U15434 (N_15434,N_14680,N_11621);
nand U15435 (N_15435,N_12986,N_12706);
and U15436 (N_15436,N_12064,N_13752);
xor U15437 (N_15437,N_11546,N_10662);
xnor U15438 (N_15438,N_11597,N_13780);
or U15439 (N_15439,N_12981,N_12848);
nor U15440 (N_15440,N_12539,N_13713);
nand U15441 (N_15441,N_14464,N_11532);
and U15442 (N_15442,N_14644,N_13396);
nor U15443 (N_15443,N_13395,N_12917);
nor U15444 (N_15444,N_10354,N_13453);
nand U15445 (N_15445,N_10128,N_14042);
and U15446 (N_15446,N_10142,N_10462);
nand U15447 (N_15447,N_11849,N_10987);
nor U15448 (N_15448,N_13664,N_11848);
nand U15449 (N_15449,N_11045,N_11298);
and U15450 (N_15450,N_11129,N_10635);
nand U15451 (N_15451,N_10238,N_13169);
xor U15452 (N_15452,N_13413,N_13997);
nand U15453 (N_15453,N_14643,N_14922);
or U15454 (N_15454,N_14650,N_14676);
nand U15455 (N_15455,N_14245,N_11846);
and U15456 (N_15456,N_12233,N_11404);
or U15457 (N_15457,N_14463,N_11278);
nor U15458 (N_15458,N_13344,N_10449);
or U15459 (N_15459,N_10337,N_14592);
xnor U15460 (N_15460,N_10002,N_11456);
and U15461 (N_15461,N_12606,N_12345);
nor U15462 (N_15462,N_13012,N_12998);
or U15463 (N_15463,N_13648,N_12306);
xnor U15464 (N_15464,N_14989,N_13726);
or U15465 (N_15465,N_13351,N_10404);
or U15466 (N_15466,N_10239,N_11507);
and U15467 (N_15467,N_14541,N_12797);
or U15468 (N_15468,N_11335,N_11219);
and U15469 (N_15469,N_13630,N_11457);
and U15470 (N_15470,N_10501,N_11198);
xnor U15471 (N_15471,N_12885,N_12553);
nand U15472 (N_15472,N_13977,N_11054);
xor U15473 (N_15473,N_12569,N_14324);
nand U15474 (N_15474,N_13825,N_11753);
xnor U15475 (N_15475,N_12168,N_14862);
and U15476 (N_15476,N_14705,N_13687);
and U15477 (N_15477,N_14049,N_12805);
xor U15478 (N_15478,N_11132,N_12114);
xnor U15479 (N_15479,N_13312,N_11124);
nand U15480 (N_15480,N_13139,N_10763);
nor U15481 (N_15481,N_10280,N_12214);
nand U15482 (N_15482,N_10394,N_10251);
xnor U15483 (N_15483,N_11238,N_11358);
or U15484 (N_15484,N_14470,N_10840);
nand U15485 (N_15485,N_11157,N_11450);
and U15486 (N_15486,N_13762,N_14240);
xnor U15487 (N_15487,N_12968,N_13296);
and U15488 (N_15488,N_14767,N_11351);
or U15489 (N_15489,N_13794,N_14223);
nor U15490 (N_15490,N_14142,N_14390);
xnor U15491 (N_15491,N_13653,N_10855);
or U15492 (N_15492,N_13098,N_12216);
nor U15493 (N_15493,N_11751,N_11486);
xor U15494 (N_15494,N_14820,N_12292);
xor U15495 (N_15495,N_10552,N_11937);
nand U15496 (N_15496,N_14875,N_14225);
nor U15497 (N_15497,N_10441,N_11424);
nor U15498 (N_15498,N_14778,N_13243);
and U15499 (N_15499,N_14409,N_10286);
and U15500 (N_15500,N_12408,N_12878);
xor U15501 (N_15501,N_13218,N_14775);
or U15502 (N_15502,N_12978,N_13992);
nand U15503 (N_15503,N_14202,N_10341);
xnor U15504 (N_15504,N_12982,N_13160);
nand U15505 (N_15505,N_10324,N_10866);
nor U15506 (N_15506,N_10459,N_14238);
and U15507 (N_15507,N_11350,N_12934);
xnor U15508 (N_15508,N_14022,N_13593);
xnor U15509 (N_15509,N_10982,N_12501);
xnor U15510 (N_15510,N_10546,N_11502);
xnor U15511 (N_15511,N_12828,N_13481);
xnor U15512 (N_15512,N_14629,N_11085);
xor U15513 (N_15513,N_14721,N_11646);
or U15514 (N_15514,N_13621,N_13584);
xnor U15515 (N_15515,N_11734,N_12071);
xnor U15516 (N_15516,N_10244,N_11757);
nor U15517 (N_15517,N_10530,N_11011);
and U15518 (N_15518,N_12574,N_11366);
nand U15519 (N_15519,N_13101,N_10815);
and U15520 (N_15520,N_13295,N_12947);
or U15521 (N_15521,N_13751,N_14581);
or U15522 (N_15522,N_14567,N_11576);
xor U15523 (N_15523,N_11459,N_12565);
xor U15524 (N_15524,N_13757,N_13885);
nand U15525 (N_15525,N_11377,N_11035);
and U15526 (N_15526,N_14534,N_13321);
or U15527 (N_15527,N_13892,N_11878);
nor U15528 (N_15528,N_13225,N_11825);
xor U15529 (N_15529,N_14014,N_10877);
nand U15530 (N_15530,N_11814,N_10627);
xor U15531 (N_15531,N_14708,N_14196);
xor U15532 (N_15532,N_10566,N_10347);
or U15533 (N_15533,N_10362,N_13756);
or U15534 (N_15534,N_10361,N_13724);
nor U15535 (N_15535,N_12418,N_12290);
or U15536 (N_15536,N_13293,N_12515);
or U15537 (N_15537,N_11802,N_10988);
or U15538 (N_15538,N_10293,N_11370);
nand U15539 (N_15539,N_14539,N_13533);
nor U15540 (N_15540,N_10129,N_13980);
nor U15541 (N_15541,N_10937,N_11569);
nand U15542 (N_15542,N_12128,N_11156);
xnor U15543 (N_15543,N_11125,N_13237);
nand U15544 (N_15544,N_10567,N_12160);
nor U15545 (N_15545,N_13938,N_12838);
or U15546 (N_15546,N_12726,N_14799);
or U15547 (N_15547,N_10156,N_13107);
nor U15548 (N_15548,N_12849,N_11346);
xnor U15549 (N_15549,N_14170,N_11374);
or U15550 (N_15550,N_11705,N_13425);
nor U15551 (N_15551,N_11017,N_10878);
nor U15552 (N_15552,N_14722,N_14500);
and U15553 (N_15553,N_14738,N_14803);
nor U15554 (N_15554,N_13587,N_13700);
xnor U15555 (N_15555,N_12915,N_13962);
nand U15556 (N_15556,N_10225,N_14127);
xnor U15557 (N_15557,N_12587,N_14916);
nor U15558 (N_15558,N_14442,N_11636);
xnor U15559 (N_15559,N_11911,N_13331);
xor U15560 (N_15560,N_14306,N_13709);
nand U15561 (N_15561,N_14586,N_13510);
or U15562 (N_15562,N_11241,N_10747);
or U15563 (N_15563,N_13501,N_12268);
xor U15564 (N_15564,N_13370,N_10998);
or U15565 (N_15565,N_10396,N_11679);
xor U15566 (N_15566,N_10030,N_13152);
nor U15567 (N_15567,N_11689,N_14754);
nand U15568 (N_15568,N_13504,N_14176);
nor U15569 (N_15569,N_10770,N_10395);
nand U15570 (N_15570,N_11699,N_14162);
nand U15571 (N_15571,N_10317,N_13627);
nor U15572 (N_15572,N_10680,N_11590);
xor U15573 (N_15573,N_11613,N_12540);
and U15574 (N_15574,N_12918,N_10049);
nor U15575 (N_15575,N_12476,N_11175);
and U15576 (N_15576,N_14385,N_13539);
and U15577 (N_15577,N_12894,N_13649);
and U15578 (N_15578,N_13838,N_11749);
and U15579 (N_15579,N_14483,N_13127);
or U15580 (N_15580,N_14062,N_10814);
nand U15581 (N_15581,N_13744,N_11263);
nand U15582 (N_15582,N_10305,N_14087);
nand U15583 (N_15583,N_11222,N_13784);
and U15584 (N_15584,N_12551,N_10067);
or U15585 (N_15585,N_11737,N_11399);
or U15586 (N_15586,N_14423,N_14679);
nor U15587 (N_15587,N_14358,N_11707);
nand U15588 (N_15588,N_13827,N_12480);
xnor U15589 (N_15589,N_12963,N_14788);
xor U15590 (N_15590,N_12571,N_11180);
nor U15591 (N_15591,N_10229,N_10240);
nor U15592 (N_15592,N_10143,N_14612);
and U15593 (N_15593,N_11823,N_12589);
nand U15594 (N_15594,N_14647,N_13891);
or U15595 (N_15595,N_14807,N_14840);
nor U15596 (N_15596,N_12638,N_14445);
xor U15597 (N_15597,N_11353,N_10083);
nor U15598 (N_15598,N_13719,N_12466);
xnor U15599 (N_15599,N_12729,N_10228);
or U15600 (N_15600,N_12055,N_12108);
or U15601 (N_15601,N_10087,N_12562);
nor U15602 (N_15602,N_14864,N_11492);
nand U15603 (N_15603,N_13582,N_11629);
and U15604 (N_15604,N_12827,N_12158);
nor U15605 (N_15605,N_14590,N_11306);
nand U15606 (N_15606,N_11775,N_13389);
xnor U15607 (N_15607,N_14511,N_12487);
nand U15608 (N_15608,N_13926,N_11959);
xnor U15609 (N_15609,N_11029,N_10478);
xnor U15610 (N_15610,N_10656,N_13356);
xor U15611 (N_15611,N_12990,N_14718);
or U15612 (N_15612,N_10338,N_14921);
nand U15613 (N_15613,N_12243,N_10254);
and U15614 (N_15614,N_10215,N_10901);
or U15615 (N_15615,N_14747,N_13890);
xnor U15616 (N_15616,N_13937,N_10938);
nand U15617 (N_15617,N_12955,N_12146);
xnor U15618 (N_15618,N_12887,N_12457);
nand U15619 (N_15619,N_14187,N_13856);
or U15620 (N_15620,N_12505,N_12475);
and U15621 (N_15621,N_14010,N_13491);
or U15622 (N_15622,N_11716,N_12364);
nand U15623 (N_15623,N_14429,N_10264);
xor U15624 (N_15624,N_14510,N_11754);
nand U15625 (N_15625,N_10480,N_14132);
or U15626 (N_15626,N_14254,N_12906);
xnor U15627 (N_15627,N_11586,N_13313);
nor U15628 (N_15628,N_14600,N_13721);
nor U15629 (N_15629,N_14488,N_10782);
and U15630 (N_15630,N_11250,N_13831);
or U15631 (N_15631,N_12512,N_13782);
nor U15632 (N_15632,N_14571,N_10374);
xnor U15633 (N_15633,N_11811,N_10197);
and U15634 (N_15634,N_13182,N_11284);
and U15635 (N_15635,N_12253,N_13505);
or U15636 (N_15636,N_10571,N_11889);
or U15637 (N_15637,N_13684,N_10150);
nor U15638 (N_15638,N_13248,N_14525);
xnor U15639 (N_15639,N_14116,N_14517);
or U15640 (N_15640,N_14784,N_11339);
xnor U15641 (N_15641,N_14836,N_11401);
or U15642 (N_15642,N_10071,N_14457);
and U15643 (N_15643,N_11549,N_11675);
xor U15644 (N_15644,N_14040,N_12549);
nor U15645 (N_15645,N_13953,N_12485);
nand U15646 (N_15646,N_12202,N_10166);
nand U15647 (N_15647,N_14878,N_10108);
nor U15648 (N_15648,N_10365,N_14562);
or U15649 (N_15649,N_11873,N_13468);
nor U15650 (N_15650,N_11127,N_14494);
nand U15651 (N_15651,N_14758,N_11870);
nand U15652 (N_15652,N_14804,N_10848);
and U15653 (N_15653,N_11519,N_10638);
or U15654 (N_15654,N_13834,N_10587);
nand U15655 (N_15655,N_13355,N_13830);
nand U15656 (N_15656,N_12244,N_13842);
nand U15657 (N_15657,N_12230,N_10787);
xor U15658 (N_15658,N_10184,N_14130);
or U15659 (N_15659,N_11121,N_13474);
nor U15660 (N_15660,N_12450,N_11148);
nand U15661 (N_15661,N_12199,N_13144);
nand U15662 (N_15662,N_11697,N_14434);
nor U15663 (N_15663,N_11227,N_10562);
xor U15664 (N_15664,N_14121,N_12734);
nor U15665 (N_15665,N_11731,N_11229);
nand U15666 (N_15666,N_11518,N_13959);
nor U15667 (N_15667,N_13746,N_12511);
or U15668 (N_15668,N_13456,N_10801);
xor U15669 (N_15669,N_12107,N_11384);
nand U15670 (N_15670,N_12387,N_11230);
nor U15671 (N_15671,N_12082,N_10308);
nand U15672 (N_15672,N_12548,N_10876);
nor U15673 (N_15673,N_12547,N_10634);
and U15674 (N_15674,N_13222,N_11499);
and U15675 (N_15675,N_11678,N_12984);
nor U15676 (N_15676,N_12975,N_14931);
xnor U15677 (N_15677,N_11952,N_10648);
nand U15678 (N_15678,N_13277,N_14076);
and U15679 (N_15679,N_11933,N_14634);
xnor U15680 (N_15680,N_14105,N_10250);
nand U15681 (N_15681,N_12759,N_13857);
nor U15682 (N_15682,N_14757,N_13785);
or U15683 (N_15683,N_12744,N_11260);
nand U15684 (N_15684,N_13095,N_12223);
nand U15685 (N_15685,N_12133,N_10134);
nor U15686 (N_15686,N_14771,N_10843);
nor U15687 (N_15687,N_13437,N_14080);
xor U15688 (N_15688,N_14030,N_13712);
xor U15689 (N_15689,N_12386,N_11554);
nor U15690 (N_15690,N_12747,N_10946);
xor U15691 (N_15691,N_10631,N_14404);
and U15692 (N_15692,N_12231,N_10241);
xor U15693 (N_15693,N_14287,N_11965);
and U15694 (N_15694,N_13142,N_10464);
and U15695 (N_15695,N_14772,N_13736);
xnor U15696 (N_15696,N_14092,N_12367);
nor U15697 (N_15697,N_11565,N_11939);
xnor U15698 (N_15698,N_10554,N_10391);
nand U15699 (N_15699,N_13074,N_12745);
xor U15700 (N_15700,N_11564,N_10001);
or U15701 (N_15701,N_11744,N_12640);
xor U15702 (N_15702,N_12096,N_12583);
xor U15703 (N_15703,N_14462,N_12543);
nor U15704 (N_15704,N_10208,N_12186);
nand U15705 (N_15705,N_12348,N_12440);
nor U15706 (N_15706,N_13297,N_13728);
nor U15707 (N_15707,N_10331,N_12401);
xnor U15708 (N_15708,N_10661,N_11842);
nor U15709 (N_15709,N_11039,N_14219);
xnor U15710 (N_15710,N_14628,N_12994);
xor U15711 (N_15711,N_13058,N_11867);
and U15712 (N_15712,N_13906,N_10936);
xor U15713 (N_15713,N_14668,N_12458);
and U15714 (N_15714,N_14431,N_13000);
nor U15715 (N_15715,N_12844,N_11214);
nand U15716 (N_15716,N_12777,N_14867);
or U15717 (N_15717,N_12851,N_11592);
nor U15718 (N_15718,N_11123,N_14887);
nand U15719 (N_15719,N_14995,N_12478);
nor U15720 (N_15720,N_10392,N_10375);
nor U15721 (N_15721,N_12372,N_14295);
or U15722 (N_15722,N_10925,N_11671);
nor U15723 (N_15723,N_11599,N_11327);
or U15724 (N_15724,N_14468,N_14316);
nand U15725 (N_15725,N_10772,N_10960);
nand U15726 (N_15726,N_13286,N_14214);
nor U15727 (N_15727,N_14941,N_12221);
and U15728 (N_15728,N_13594,N_12380);
nor U15729 (N_15729,N_12956,N_14885);
and U15730 (N_15730,N_14573,N_10173);
xnor U15731 (N_15731,N_11352,N_12097);
nand U15732 (N_15732,N_13662,N_14252);
or U15733 (N_15733,N_13245,N_11542);
and U15734 (N_15734,N_14161,N_14267);
and U15735 (N_15735,N_14928,N_10461);
and U15736 (N_15736,N_13023,N_10944);
nand U15737 (N_15737,N_14866,N_12122);
xnor U15738 (N_15738,N_14310,N_10584);
and U15739 (N_15739,N_12525,N_10513);
or U15740 (N_15740,N_10381,N_12902);
nor U15741 (N_15741,N_14149,N_14098);
xnor U15742 (N_15742,N_14394,N_10819);
nor U15743 (N_15743,N_13050,N_10736);
nor U15744 (N_15744,N_14550,N_14814);
and U15745 (N_15745,N_14764,N_13872);
xor U15746 (N_15746,N_12796,N_12383);
nor U15747 (N_15747,N_11396,N_10643);
nand U15748 (N_15748,N_11448,N_13002);
nor U15749 (N_15749,N_12648,N_13920);
and U15750 (N_15750,N_11144,N_11953);
or U15751 (N_15751,N_11628,N_10011);
or U15752 (N_15752,N_14249,N_13984);
and U15753 (N_15753,N_12899,N_12996);
or U15754 (N_15754,N_11611,N_12240);
xnor U15755 (N_15755,N_12989,N_13574);
nor U15756 (N_15756,N_10500,N_12980);
nor U15757 (N_15757,N_10533,N_12004);
or U15758 (N_15758,N_11474,N_10553);
and U15759 (N_15759,N_11701,N_13147);
or U15760 (N_15760,N_10435,N_13542);
nor U15761 (N_15761,N_13320,N_13974);
nor U15762 (N_15762,N_10062,N_14942);
or U15763 (N_15763,N_11226,N_10741);
and U15764 (N_15764,N_13340,N_14703);
xnor U15765 (N_15765,N_14236,N_13093);
nor U15766 (N_15766,N_14111,N_12285);
or U15767 (N_15767,N_12497,N_14985);
or U15768 (N_15768,N_11868,N_11234);
or U15769 (N_15769,N_14029,N_13250);
and U15770 (N_15770,N_13394,N_10055);
nor U15771 (N_15771,N_11381,N_14564);
or U15772 (N_15772,N_10403,N_11282);
nand U15773 (N_15773,N_10497,N_11348);
or U15774 (N_15774,N_12301,N_10260);
or U15775 (N_15775,N_13490,N_12841);
nand U15776 (N_15776,N_11799,N_11997);
nand U15777 (N_15777,N_14707,N_14904);
or U15778 (N_15778,N_12600,N_14582);
and U15779 (N_15779,N_10282,N_10835);
or U15780 (N_15780,N_10170,N_10457);
xnor U15781 (N_15781,N_10123,N_14839);
nand U15782 (N_15782,N_11760,N_12147);
or U15783 (N_15783,N_13839,N_11103);
nor U15784 (N_15784,N_13388,N_13057);
or U15785 (N_15785,N_11067,N_14246);
nor U15786 (N_15786,N_13092,N_13352);
or U15787 (N_15787,N_11588,N_11706);
xor U15788 (N_15788,N_12403,N_14524);
nand U15789 (N_15789,N_11687,N_13457);
xor U15790 (N_15790,N_10774,N_12646);
nand U15791 (N_15791,N_12248,N_11808);
nand U15792 (N_15792,N_13307,N_10953);
or U15793 (N_15793,N_10942,N_14819);
nand U15794 (N_15794,N_10614,N_14675);
nor U15795 (N_15795,N_11836,N_12710);
or U15796 (N_15796,N_10056,N_10484);
and U15797 (N_15797,N_11722,N_10453);
nor U15798 (N_15798,N_12629,N_10572);
and U15799 (N_15799,N_13106,N_14253);
or U15800 (N_15800,N_14734,N_12690);
nand U15801 (N_15801,N_10612,N_10909);
nor U15802 (N_15802,N_13716,N_13345);
or U15803 (N_15803,N_12767,N_14250);
xnor U15804 (N_15804,N_11324,N_13465);
nor U15805 (N_15805,N_10190,N_13314);
xor U15806 (N_15806,N_13283,N_10788);
nand U15807 (N_15807,N_13954,N_14597);
and U15808 (N_15808,N_13889,N_14452);
xor U15809 (N_15809,N_13528,N_11924);
and U15810 (N_15810,N_12645,N_12388);
and U15811 (N_15811,N_12073,N_11179);
xnor U15812 (N_15812,N_12770,N_11224);
and U15813 (N_15813,N_10730,N_13943);
or U15814 (N_15814,N_11663,N_14183);
and U15815 (N_15815,N_11508,N_10269);
xnor U15816 (N_15816,N_11762,N_10256);
and U15817 (N_15817,N_14451,N_13503);
or U15818 (N_15818,N_11791,N_14833);
or U15819 (N_15819,N_10136,N_11667);
nor U15820 (N_15820,N_13628,N_10262);
nand U15821 (N_15821,N_12182,N_10907);
or U15822 (N_15822,N_12842,N_13444);
nor U15823 (N_15823,N_14798,N_14684);
nand U15824 (N_15824,N_12730,N_12426);
nor U15825 (N_15825,N_10407,N_13779);
xnor U15826 (N_15826,N_12507,N_11971);
and U15827 (N_15827,N_10939,N_12867);
or U15828 (N_15828,N_14327,N_11895);
xor U15829 (N_15829,N_11988,N_11563);
nand U15830 (N_15830,N_10816,N_14472);
nand U15831 (N_15831,N_12870,N_10735);
or U15832 (N_15832,N_10602,N_11016);
nand U15833 (N_15833,N_13999,N_12630);
nand U15834 (N_15834,N_12607,N_12315);
nand U15835 (N_15835,N_11528,N_14918);
nor U15836 (N_15836,N_12198,N_12050);
and U15837 (N_15837,N_13590,N_11567);
and U15838 (N_15838,N_10771,N_13941);
nor U15839 (N_15839,N_12735,N_13645);
or U15840 (N_15840,N_13073,N_12871);
xnor U15841 (N_15841,N_11187,N_11733);
nand U15842 (N_15842,N_14218,N_13604);
nor U15843 (N_15843,N_13212,N_14067);
nand U15844 (N_15844,N_13083,N_14792);
or U15845 (N_15845,N_14212,N_14008);
xor U15846 (N_15846,N_14056,N_11246);
xor U15847 (N_15847,N_11913,N_13806);
nand U15848 (N_15848,N_14793,N_10997);
or U15849 (N_15849,N_13675,N_13915);
nand U15850 (N_15850,N_14540,N_11197);
or U15851 (N_15851,N_10232,N_14570);
nor U15852 (N_15852,N_12181,N_10637);
nand U15853 (N_15853,N_11531,N_11695);
or U15854 (N_15854,N_12013,N_10990);
and U15855 (N_15855,N_14364,N_13099);
xnor U15856 (N_15856,N_13403,N_11462);
or U15857 (N_15857,N_14551,N_14400);
or U15858 (N_15858,N_11126,N_13028);
and U15859 (N_15859,N_10632,N_10451);
xor U15860 (N_15860,N_12812,N_13482);
or U15861 (N_15861,N_14658,N_14870);
nor U15862 (N_15862,N_10382,N_13506);
nand U15863 (N_15863,N_12868,N_13372);
and U15864 (N_15864,N_11375,N_12820);
nand U15865 (N_15865,N_14662,N_14109);
xor U15866 (N_15866,N_11333,N_14314);
or U15867 (N_15867,N_12687,N_14038);
nand U15868 (N_15868,N_13983,N_14824);
nand U15869 (N_15869,N_14028,N_13768);
xnor U15870 (N_15870,N_13769,N_10379);
xor U15871 (N_15871,N_13441,N_12111);
or U15872 (N_15872,N_13685,N_12326);
or U15873 (N_15873,N_10590,N_14186);
and U15874 (N_15874,N_14659,N_13778);
xor U15875 (N_15875,N_11906,N_11289);
nor U15876 (N_15876,N_12792,N_10102);
and U15877 (N_15877,N_10869,N_12250);
or U15878 (N_15878,N_13930,N_12264);
or U15879 (N_15879,N_12960,N_10863);
and U15880 (N_15880,N_12030,N_14986);
nand U15881 (N_15881,N_14263,N_11816);
or U15882 (N_15882,N_14933,N_13601);
xor U15883 (N_15883,N_13617,N_10910);
xnor U15884 (N_15884,N_11680,N_11093);
xor U15885 (N_15885,N_12958,N_11302);
and U15886 (N_15886,N_10755,N_11925);
nor U15887 (N_15887,N_14781,N_13442);
xnor U15888 (N_15888,N_14609,N_14203);
nor U15889 (N_15889,N_10444,N_12705);
xor U15890 (N_15890,N_14533,N_13942);
nor U15891 (N_15891,N_14353,N_12644);
nand U15892 (N_15892,N_12094,N_11277);
xor U15893 (N_15893,N_13672,N_11165);
nand U15894 (N_15894,N_10418,N_11287);
nand U15895 (N_15895,N_10221,N_12215);
xor U15896 (N_15896,N_13090,N_13793);
xnor U15897 (N_15897,N_12105,N_10217);
or U15898 (N_15898,N_11641,N_13907);
nand U15899 (N_15899,N_13407,N_10042);
or U15900 (N_15900,N_10806,N_12966);
and U15901 (N_15901,N_13742,N_12876);
nand U15902 (N_15902,N_11538,N_14632);
xor U15903 (N_15903,N_14256,N_11455);
and U15904 (N_15904,N_12654,N_11199);
or U15905 (N_15905,N_11967,N_14897);
nor U15906 (N_15906,N_10758,N_11086);
and U15907 (N_15907,N_14054,N_13259);
xor U15908 (N_15908,N_14012,N_11496);
or U15909 (N_15909,N_14766,N_10107);
nand U15910 (N_15910,N_11866,N_12658);
nand U15911 (N_15911,N_10991,N_13771);
nand U15912 (N_15912,N_14542,N_11831);
or U15913 (N_15913,N_11098,N_13154);
nor U15914 (N_15914,N_11090,N_13919);
nand U15915 (N_15915,N_12016,N_10739);
or U15916 (N_15916,N_14123,N_11092);
xor U15917 (N_15917,N_11378,N_11583);
xor U15918 (N_15918,N_11635,N_12099);
nand U15919 (N_15919,N_14015,N_14156);
nor U15920 (N_15920,N_14374,N_14826);
nand U15921 (N_15921,N_11024,N_13945);
or U15922 (N_15922,N_11387,N_11688);
or U15923 (N_15923,N_12119,N_13922);
nor U15924 (N_15924,N_14032,N_13660);
nor U15925 (N_15925,N_12080,N_10534);
and U15926 (N_15926,N_14770,N_10506);
or U15927 (N_15927,N_12584,N_11515);
or U15928 (N_15928,N_11158,N_13291);
or U15929 (N_15929,N_12327,N_10499);
nor U15930 (N_15930,N_13228,N_14179);
xor U15931 (N_15931,N_14321,N_11328);
and U15932 (N_15932,N_12731,N_13921);
nor U15933 (N_15933,N_13265,N_13451);
xnor U15934 (N_15934,N_14858,N_13747);
or U15935 (N_15935,N_11790,N_13161);
nand U15936 (N_15936,N_14496,N_10016);
and U15937 (N_15937,N_11480,N_11212);
or U15938 (N_15938,N_12723,N_11467);
or U15939 (N_15939,N_13864,N_13385);
nand U15940 (N_15940,N_13661,N_10113);
and U15941 (N_15941,N_10579,N_11622);
xor U15942 (N_15942,N_10768,N_13665);
xor U15943 (N_15943,N_13766,N_12431);
nand U15944 (N_15944,N_14126,N_10868);
xnor U15945 (N_15945,N_13262,N_11852);
nor U15946 (N_15946,N_14815,N_10914);
xnor U15947 (N_15947,N_10277,N_11767);
xnor U15948 (N_15948,N_13480,N_10813);
or U15949 (N_15949,N_12136,N_13633);
or U15950 (N_15950,N_10683,N_10964);
nor U15951 (N_15951,N_13530,N_11573);
nand U15952 (N_15952,N_14454,N_11630);
nor U15953 (N_15953,N_10471,N_12862);
or U15954 (N_15954,N_14695,N_13866);
nor U15955 (N_15955,N_13571,N_14391);
and U15956 (N_15956,N_11600,N_11326);
and U15957 (N_15957,N_12683,N_10738);
nor U15958 (N_15958,N_13874,N_11188);
or U15959 (N_15959,N_12046,N_13108);
nand U15960 (N_15960,N_10891,N_14529);
nand U15961 (N_15961,N_14951,N_10414);
xnor U15962 (N_15962,N_13924,N_14425);
or U15963 (N_15963,N_14401,N_11720);
nand U15964 (N_15964,N_10149,N_10655);
nand U15965 (N_15965,N_13730,N_12962);
nor U15966 (N_15966,N_11343,N_13535);
xnor U15967 (N_15967,N_12336,N_10716);
nor U15968 (N_15968,N_14809,N_11610);
or U15969 (N_15969,N_14146,N_10978);
nand U15970 (N_15970,N_13516,N_14777);
and U15971 (N_15971,N_14197,N_10486);
nor U15972 (N_15972,N_10503,N_11412);
and U15973 (N_15973,N_12279,N_12761);
and U15974 (N_15974,N_12803,N_13258);
nor U15975 (N_15975,N_14151,N_13767);
xnor U15976 (N_15976,N_14880,N_14143);
xnor U15977 (N_15977,N_14657,N_11320);
or U15978 (N_15978,N_11627,N_11838);
or U15979 (N_15979,N_13289,N_12628);
and U15980 (N_15980,N_12712,N_12286);
or U15981 (N_15981,N_12582,N_10494);
nor U15982 (N_15982,N_12001,N_13438);
nor U15983 (N_15983,N_11256,N_11213);
or U15984 (N_15984,N_13255,N_14547);
xor U15985 (N_15985,N_10137,N_12178);
and U15986 (N_15986,N_12932,N_13300);
and U15987 (N_15987,N_10667,N_12741);
nand U15988 (N_15988,N_14513,N_14907);
or U15989 (N_15989,N_10447,N_11897);
and U15990 (N_15990,N_13132,N_10348);
nor U15991 (N_15991,N_11345,N_14617);
and U15992 (N_15992,N_14291,N_11944);
nand U15993 (N_15993,N_12889,N_13181);
xor U15994 (N_15994,N_13412,N_11361);
xnor U15995 (N_15995,N_14959,N_13879);
nand U15996 (N_15996,N_12669,N_12208);
nor U15997 (N_15997,N_13466,N_10980);
and U15998 (N_15998,N_10152,N_11173);
or U15999 (N_15999,N_11703,N_14180);
nand U16000 (N_16000,N_10721,N_13809);
or U16001 (N_16001,N_10972,N_11803);
and U16002 (N_16002,N_14174,N_11704);
and U16003 (N_16003,N_13553,N_14890);
or U16004 (N_16004,N_10852,N_10707);
nor U16005 (N_16005,N_13137,N_11088);
xnor U16006 (N_16006,N_13932,N_10508);
and U16007 (N_16007,N_13068,N_11101);
nor U16008 (N_16008,N_10146,N_11014);
xnor U16009 (N_16009,N_14373,N_11102);
nor U16010 (N_16010,N_13014,N_12952);
xnor U16011 (N_16011,N_12323,N_11652);
xor U16012 (N_16012,N_13056,N_10364);
nand U16013 (N_16013,N_11391,N_10279);
nor U16014 (N_16014,N_12191,N_12124);
nand U16015 (N_16015,N_13036,N_10966);
nor U16016 (N_16016,N_10131,N_12591);
nand U16017 (N_16017,N_11612,N_14681);
and U16018 (N_16018,N_11447,N_10523);
nand U16019 (N_16019,N_12451,N_12358);
xor U16020 (N_16020,N_14655,N_10519);
xnor U16021 (N_16021,N_10912,N_10619);
nand U16022 (N_16022,N_11850,N_12778);
xnor U16023 (N_16023,N_11040,N_11859);
or U16024 (N_16024,N_12473,N_14339);
nor U16025 (N_16025,N_12914,N_14688);
nand U16026 (N_16026,N_12681,N_14633);
xor U16027 (N_16027,N_11741,N_13802);
nor U16028 (N_16028,N_12623,N_11725);
nor U16029 (N_16029,N_13903,N_13979);
or U16030 (N_16030,N_11992,N_10518);
nand U16031 (N_16031,N_12577,N_12162);
and U16032 (N_16032,N_11970,N_13311);
nor U16033 (N_16033,N_11510,N_10047);
and U16034 (N_16034,N_10693,N_11183);
and U16035 (N_16035,N_14666,N_14901);
nand U16036 (N_16036,N_12344,N_14412);
or U16037 (N_16037,N_12524,N_12992);
nand U16038 (N_16038,N_14561,N_11363);
nor U16039 (N_16039,N_14258,N_10028);
nand U16040 (N_16040,N_12673,N_14140);
nand U16041 (N_16041,N_14091,N_13823);
nand U16042 (N_16042,N_14637,N_13738);
nand U16043 (N_16043,N_11372,N_13699);
nor U16044 (N_16044,N_14262,N_11639);
xor U16045 (N_16045,N_11013,N_11581);
xor U16046 (N_16046,N_12794,N_12764);
nor U16047 (N_16047,N_10216,N_10517);
nor U16048 (N_16048,N_10636,N_13976);
nor U16049 (N_16049,N_14678,N_11489);
xnor U16050 (N_16050,N_10054,N_11009);
and U16051 (N_16051,N_11781,N_13884);
xnor U16052 (N_16052,N_11962,N_10540);
nor U16053 (N_16053,N_12699,N_14071);
and U16054 (N_16054,N_10265,N_14602);
nand U16055 (N_16055,N_10018,N_12795);
nor U16056 (N_16056,N_11620,N_14247);
and U16057 (N_16057,N_13723,N_13357);
or U16058 (N_16058,N_14131,N_10483);
or U16059 (N_16059,N_13801,N_10366);
nand U16060 (N_16060,N_14779,N_14475);
or U16061 (N_16061,N_10542,N_11801);
nand U16062 (N_16062,N_11659,N_13691);
nor U16063 (N_16063,N_14458,N_11658);
and U16064 (N_16064,N_13326,N_12696);
and U16065 (N_16065,N_10548,N_14677);
and U16066 (N_16066,N_11369,N_14328);
xnor U16067 (N_16067,N_13711,N_13536);
nor U16068 (N_16068,N_14433,N_14914);
nor U16069 (N_16069,N_10191,N_13348);
nand U16070 (N_16070,N_11694,N_13573);
and U16071 (N_16071,N_14025,N_11888);
and U16072 (N_16072,N_12927,N_11110);
and U16073 (N_16073,N_11050,N_10431);
nor U16074 (N_16074,N_13153,N_11779);
xor U16075 (N_16075,N_10333,N_11740);
nand U16076 (N_16076,N_11596,N_10188);
and U16077 (N_16077,N_13096,N_10906);
nor U16078 (N_16078,N_14521,N_14153);
xor U16079 (N_16079,N_10106,N_14969);
nor U16080 (N_16080,N_14893,N_14998);
or U16081 (N_16081,N_12948,N_11661);
nand U16082 (N_16082,N_12912,N_12429);
and U16083 (N_16083,N_11708,N_12940);
xnor U16084 (N_16084,N_11557,N_11765);
xor U16085 (N_16085,N_11525,N_13902);
and U16086 (N_16086,N_12561,N_14495);
nor U16087 (N_16087,N_14967,N_14302);
and U16088 (N_16088,N_11209,N_10756);
and U16089 (N_16089,N_13271,N_13005);
nor U16090 (N_16090,N_12882,N_10373);
or U16091 (N_16091,N_10695,N_13875);
or U16092 (N_16092,N_13180,N_14763);
xor U16093 (N_16093,N_13841,N_13239);
xnor U16094 (N_16094,N_11177,N_10611);
xor U16095 (N_16095,N_12891,N_12489);
xnor U16096 (N_16096,N_11651,N_14584);
nand U16097 (N_16097,N_14762,N_13048);
or U16098 (N_16098,N_10538,N_14844);
xor U16099 (N_16099,N_13432,N_11033);
xnor U16100 (N_16100,N_13955,N_10195);
xnor U16101 (N_16101,N_13242,N_11691);
and U16102 (N_16102,N_14211,N_12130);
nand U16103 (N_16103,N_12148,N_12144);
nand U16104 (N_16104,N_14282,N_10313);
nor U16105 (N_16105,N_11936,N_14522);
nand U16106 (N_16106,N_11410,N_11360);
and U16107 (N_16107,N_12247,N_13509);
or U16108 (N_16108,N_14095,N_13025);
nor U16109 (N_16109,N_11615,N_12752);
xor U16110 (N_16110,N_13760,N_13667);
nand U16111 (N_16111,N_12760,N_10355);
nand U16112 (N_16112,N_14384,N_12299);
xor U16113 (N_16113,N_11470,N_14284);
nor U16114 (N_16114,N_13616,N_12716);
and U16115 (N_16115,N_12066,N_11860);
and U16116 (N_16116,N_14898,N_12093);
xnor U16117 (N_16117,N_12021,N_13174);
nand U16118 (N_16118,N_12008,N_11797);
and U16119 (N_16119,N_14083,N_13973);
xnor U16120 (N_16120,N_14992,N_12965);
xnor U16121 (N_16121,N_11342,N_13611);
xnor U16122 (N_16122,N_13064,N_10475);
xor U16123 (N_16123,N_13384,N_13637);
xor U16124 (N_16124,N_12376,N_13009);
nand U16125 (N_16125,N_11750,N_12542);
nand U16126 (N_16126,N_13612,N_14925);
and U16127 (N_16127,N_11393,N_11769);
nor U16128 (N_16128,N_10900,N_14993);
and U16129 (N_16129,N_12277,N_13047);
or U16130 (N_16130,N_13749,N_12617);
xor U16131 (N_16131,N_14027,N_11318);
nor U16132 (N_16132,N_13136,N_14817);
nand U16133 (N_16133,N_12781,N_12702);
or U16134 (N_16134,N_14013,N_14566);
nand U16135 (N_16135,N_12452,N_13044);
nor U16136 (N_16136,N_14791,N_14631);
nand U16137 (N_16137,N_13958,N_11746);
nand U16138 (N_16138,N_12821,N_11007);
xnor U16139 (N_16139,N_13390,N_11931);
or U16140 (N_16140,N_12165,N_13103);
or U16141 (N_16141,N_14686,N_14514);
xor U16142 (N_16142,N_11297,N_12598);
or U16143 (N_16143,N_11792,N_11440);
nand U16144 (N_16144,N_14392,N_12857);
xor U16145 (N_16145,N_12776,N_14812);
nand U16146 (N_16146,N_14852,N_12931);
nor U16147 (N_16147,N_13897,N_13759);
nand U16148 (N_16148,N_10325,N_12213);
and U16149 (N_16149,N_14307,N_11301);
and U16150 (N_16150,N_13299,N_14554);
and U16151 (N_16151,N_14737,N_12161);
or U16152 (N_16152,N_13964,N_14293);
nand U16153 (N_16153,N_11458,N_13450);
nor U16154 (N_16154,N_10298,N_11258);
nand U16155 (N_16155,N_11879,N_12422);
xor U16156 (N_16156,N_10981,N_12295);
nor U16157 (N_16157,N_13788,N_10803);
or U16158 (N_16158,N_13579,N_14768);
or U16159 (N_16159,N_11577,N_13475);
xnor U16160 (N_16160,N_10514,N_10401);
or U16161 (N_16161,N_12808,N_11666);
nor U16162 (N_16162,N_12464,N_10915);
xnor U16163 (N_16163,N_13067,N_11973);
nand U16164 (N_16164,N_10201,N_12424);
nor U16165 (N_16165,N_14665,N_11248);
nor U16166 (N_16166,N_13052,N_12432);
or U16167 (N_16167,N_11926,N_12152);
xor U16168 (N_16168,N_10094,N_11139);
xor U16169 (N_16169,N_11354,N_11190);
nor U16170 (N_16170,N_13971,N_14430);
nand U16171 (N_16171,N_13434,N_14041);
nor U16172 (N_16172,N_10784,N_13580);
nand U16173 (N_16173,N_11425,N_10380);
and U16174 (N_16174,N_12121,N_10493);
nand U16175 (N_16175,N_11591,N_13562);
and U16176 (N_16176,N_10620,N_12395);
or U16177 (N_16177,N_13494,N_14234);
or U16178 (N_16178,N_10193,N_11713);
xnor U16179 (N_16179,N_10273,N_12142);
nand U16180 (N_16180,N_10490,N_10872);
or U16181 (N_16181,N_11649,N_11990);
nand U16182 (N_16182,N_14480,N_12678);
nand U16183 (N_16183,N_10967,N_14627);
xor U16184 (N_16184,N_14842,N_14322);
xor U16185 (N_16185,N_12737,N_11774);
xnor U16186 (N_16186,N_10027,N_13391);
nand U16187 (N_16187,N_10111,N_12579);
nand U16188 (N_16188,N_11048,N_11109);
or U16189 (N_16189,N_14437,N_10696);
or U16190 (N_16190,N_12077,N_13529);
xnor U16191 (N_16191,N_11081,N_12166);
nor U16192 (N_16192,N_12806,N_13463);
xnor U16193 (N_16193,N_12786,N_14624);
xnor U16194 (N_16194,N_13565,N_11783);
nor U16195 (N_16195,N_10581,N_13223);
or U16196 (N_16196,N_13893,N_12062);
xor U16197 (N_16197,N_11804,N_12740);
xor U16198 (N_16198,N_12722,N_12763);
nand U16199 (N_16199,N_11191,N_12400);
nand U16200 (N_16200,N_14977,N_11872);
and U16201 (N_16201,N_11657,N_14278);
or U16202 (N_16202,N_10520,N_14248);
and U16203 (N_16203,N_11415,N_12313);
nand U16204 (N_16204,N_13278,N_12532);
or U16205 (N_16205,N_10599,N_14636);
nand U16206 (N_16206,N_14072,N_14449);
or U16207 (N_16207,N_11322,N_12045);
and U16208 (N_16208,N_10737,N_12869);
nor U16209 (N_16209,N_11540,N_12033);
nand U16210 (N_16210,N_11023,N_14691);
or U16211 (N_16211,N_13323,N_12758);
and U16212 (N_16212,N_11270,N_12413);
nor U16213 (N_16213,N_11237,N_11057);
or U16214 (N_16214,N_11451,N_11770);
and U16215 (N_16215,N_13798,N_13492);
nand U16216 (N_16216,N_10529,N_10789);
and U16217 (N_16217,N_11827,N_13910);
or U16218 (N_16218,N_11601,N_11883);
and U16219 (N_16219,N_14088,N_12211);
or U16220 (N_16220,N_13201,N_14325);
xnor U16221 (N_16221,N_10639,N_13217);
nand U16222 (N_16222,N_13765,N_14537);
nor U16223 (N_16223,N_13043,N_13247);
and U16224 (N_16224,N_13346,N_13901);
nor U16225 (N_16225,N_12352,N_11522);
or U16226 (N_16226,N_10858,N_14007);
nor U16227 (N_16227,N_14594,N_10091);
xnor U16228 (N_16228,N_11951,N_11152);
xnor U16229 (N_16229,N_13342,N_13219);
nor U16230 (N_16230,N_14232,N_14018);
and U16231 (N_16231,N_11185,N_13588);
and U16232 (N_16232,N_11547,N_13703);
nand U16233 (N_16233,N_13031,N_11521);
and U16234 (N_16234,N_12865,N_10918);
xnor U16235 (N_16235,N_14037,N_11940);
and U16236 (N_16236,N_14125,N_13393);
or U16237 (N_16237,N_12893,N_11171);
nand U16238 (N_16238,N_12809,N_11500);
and U16239 (N_16239,N_13007,N_11491);
xnor U16240 (N_16240,N_10117,N_11084);
nor U16241 (N_16241,N_11299,N_12043);
and U16242 (N_16242,N_12789,N_11264);
or U16243 (N_16243,N_11530,N_10311);
and U16244 (N_16244,N_12892,N_13965);
and U16245 (N_16245,N_10715,N_13957);
nand U16246 (N_16246,N_11164,N_12619);
nor U16247 (N_16247,N_10319,N_12823);
and U16248 (N_16248,N_13063,N_10616);
and U16249 (N_16249,N_13789,N_13880);
nand U16250 (N_16250,N_13041,N_13682);
nand U16251 (N_16251,N_10468,N_14604);
or U16252 (N_16252,N_11545,N_13249);
nor U16253 (N_16253,N_12559,N_10007);
and U16254 (N_16254,N_13689,N_12325);
xor U16255 (N_16255,N_13695,N_13069);
xnor U16256 (N_16256,N_11625,N_10528);
and U16257 (N_16257,N_10329,N_10886);
and U16258 (N_16258,N_13363,N_11431);
nor U16259 (N_16259,N_12782,N_10336);
nor U16260 (N_16260,N_12098,N_13353);
and U16261 (N_16261,N_12573,N_12188);
xor U16262 (N_16262,N_12496,N_12567);
xor U16263 (N_16263,N_10762,N_14172);
nor U16264 (N_16264,N_14410,N_14687);
nand U16265 (N_16265,N_13179,N_14381);
and U16266 (N_16266,N_11523,N_11166);
and U16267 (N_16267,N_12935,N_13508);
nand U16268 (N_16268,N_10020,N_13216);
nand U16269 (N_16269,N_13018,N_12322);
or U16270 (N_16270,N_14181,N_14415);
or U16271 (N_16271,N_14837,N_13079);
nor U16272 (N_16272,N_10085,N_14097);
or U16273 (N_16273,N_12245,N_13280);
nor U16274 (N_16274,N_13994,N_11172);
and U16275 (N_16275,N_11995,N_13720);
nor U16276 (N_16276,N_13526,N_10100);
nor U16277 (N_16277,N_12852,N_12929);
nand U16278 (N_16278,N_11477,N_14755);
nor U16279 (N_16279,N_12036,N_13317);
and U16280 (N_16280,N_10626,N_14280);
xor U16281 (N_16281,N_13737,N_14963);
nor U16282 (N_16282,N_13309,N_11514);
or U16283 (N_16283,N_14823,N_13523);
xnor U16284 (N_16284,N_12200,N_11421);
or U16285 (N_16285,N_14063,N_10829);
and U16286 (N_16286,N_12120,N_14580);
and U16287 (N_16287,N_11921,N_14654);
nor U16288 (N_16288,N_10547,N_14935);
or U16289 (N_16289,N_14477,N_10874);
or U16290 (N_16290,N_11422,N_12749);
and U16291 (N_16291,N_13935,N_10779);
nor U16292 (N_16292,N_12988,N_10625);
nor U16293 (N_16293,N_12132,N_13524);
nor U16294 (N_16294,N_12444,N_13038);
and U16295 (N_16295,N_12766,N_12837);
nand U16296 (N_16296,N_14712,N_14889);
or U16297 (N_16297,N_11154,N_14395);
or U16298 (N_16298,N_11664,N_14782);
and U16299 (N_16299,N_14808,N_10063);
nor U16300 (N_16300,N_12488,N_10841);
or U16301 (N_16301,N_10064,N_11314);
nand U16302 (N_16302,N_14101,N_11784);
nor U16303 (N_16303,N_13555,N_12154);
nor U16304 (N_16304,N_11325,N_10052);
nand U16305 (N_16305,N_14797,N_12509);
nor U16306 (N_16306,N_14482,N_14512);
xor U16307 (N_16307,N_12839,N_14990);
nor U16308 (N_16308,N_14865,N_14932);
xnor U16309 (N_16309,N_13968,N_13406);
or U16310 (N_16310,N_10568,N_10026);
nor U16311 (N_16311,N_14466,N_10622);
nor U16312 (N_16312,N_11829,N_11960);
nand U16313 (N_16313,N_13776,N_13557);
and U16314 (N_16314,N_14369,N_12204);
and U16315 (N_16315,N_12049,N_10686);
or U16316 (N_16316,N_13735,N_13446);
xnor U16317 (N_16317,N_11653,N_11809);
and U16318 (N_16318,N_10749,N_10539);
nand U16319 (N_16319,N_10780,N_14122);
and U16320 (N_16320,N_11427,N_13654);
and U16321 (N_16321,N_10186,N_12101);
and U16322 (N_16322,N_12209,N_11812);
or U16323 (N_16323,N_13545,N_10314);
xor U16324 (N_16324,N_13404,N_12499);
nor U16325 (N_16325,N_12552,N_10479);
nor U16326 (N_16326,N_12544,N_10983);
nand U16327 (N_16327,N_12310,N_12257);
and U16328 (N_16328,N_10732,N_12788);
xnor U16329 (N_16329,N_10209,N_12193);
xor U16330 (N_16330,N_10161,N_13308);
and U16331 (N_16331,N_10962,N_10831);
nand U16332 (N_16332,N_14024,N_10263);
nand U16333 (N_16333,N_10921,N_14332);
nand U16334 (N_16334,N_11696,N_12874);
and U16335 (N_16335,N_13544,N_13024);
or U16336 (N_16336,N_10743,N_13822);
and U16337 (N_16337,N_10316,N_10101);
and U16338 (N_16338,N_10923,N_12141);
nor U16339 (N_16339,N_13560,N_14128);
or U16340 (N_16340,N_10989,N_14958);
xnor U16341 (N_16341,N_10198,N_10929);
or U16342 (N_16342,N_14296,N_14003);
or U16343 (N_16343,N_10443,N_12126);
and U16344 (N_16344,N_13614,N_12688);
xor U16345 (N_16345,N_14577,N_11133);
xor U16346 (N_16346,N_13256,N_10629);
or U16347 (N_16347,N_14841,N_12724);
nand U16348 (N_16348,N_11052,N_10031);
or U16349 (N_16349,N_10713,N_12317);
nand U16350 (N_16350,N_14503,N_13328);
xor U16351 (N_16351,N_13626,N_12212);
xnor U16352 (N_16352,N_12267,N_12293);
xnor U16353 (N_16353,N_10860,N_13745);
and U16354 (N_16354,N_10154,N_14911);
xnor U16355 (N_16355,N_13414,N_12771);
or U16356 (N_16356,N_10048,N_12732);
xor U16357 (N_16357,N_14583,N_13836);
nand U16358 (N_16358,N_13559,N_14835);
and U16359 (N_16359,N_12454,N_12836);
nand U16360 (N_16360,N_12846,N_13763);
or U16361 (N_16361,N_10114,N_11272);
xor U16362 (N_16362,N_14987,N_10908);
or U16363 (N_16363,N_12557,N_11060);
and U16364 (N_16364,N_11305,N_12404);
or U16365 (N_16365,N_14376,N_10956);
nor U16366 (N_16366,N_10668,N_12641);
or U16367 (N_16367,N_13008,N_13409);
xor U16368 (N_16368,N_14086,N_12076);
nor U16369 (N_16369,N_11064,N_13042);
xnor U16370 (N_16370,N_14971,N_11311);
nand U16371 (N_16371,N_11607,N_13686);
nand U16372 (N_16372,N_13362,N_14360);
nand U16373 (N_16373,N_14058,N_13914);
and U16374 (N_16374,N_11647,N_14598);
nand U16375 (N_16375,N_12296,N_11739);
or U16376 (N_16376,N_11323,N_12249);
nor U16377 (N_16377,N_14421,N_13819);
or U16378 (N_16378,N_11553,N_14418);
or U16379 (N_16379,N_11454,N_11690);
or U16380 (N_16380,N_11527,N_12768);
nor U16381 (N_16381,N_10728,N_13499);
and U16382 (N_16382,N_14685,N_12282);
nor U16383 (N_16383,N_12546,N_11794);
and U16384 (N_16384,N_11835,N_11631);
xnor U16385 (N_16385,N_14077,N_11056);
nor U16386 (N_16386,N_12177,N_10825);
or U16387 (N_16387,N_14506,N_13301);
and U16388 (N_16388,N_13123,N_10084);
or U16389 (N_16389,N_11856,N_14241);
nand U16390 (N_16390,N_12636,N_10521);
nor U16391 (N_16391,N_13118,N_13399);
nor U16392 (N_16392,N_12005,N_10802);
or U16393 (N_16393,N_11534,N_13996);
nor U16394 (N_16394,N_12456,N_10255);
or U16395 (N_16395,N_13155,N_12065);
and U16396 (N_16396,N_13636,N_10999);
and U16397 (N_16397,N_10068,N_10650);
nand U16398 (N_16398,N_10618,N_14753);
xnor U16399 (N_16399,N_13548,N_11186);
nor U16400 (N_16400,N_13644,N_12682);
nor U16401 (N_16401,N_11235,N_13592);
xnor U16402 (N_16402,N_12224,N_10281);
nand U16403 (N_16403,N_12637,N_14761);
and U16404 (N_16404,N_13904,N_10420);
nand U16405 (N_16405,N_12460,N_13563);
nor U16406 (N_16406,N_12599,N_11580);
xor U16407 (N_16407,N_10321,N_13800);
xor U16408 (N_16408,N_13055,N_10388);
and U16409 (N_16409,N_11810,N_14574);
and U16410 (N_16410,N_12183,N_11901);
nor U16411 (N_16411,N_10740,N_14147);
xnor U16412 (N_16412,N_14930,N_12007);
or U16413 (N_16413,N_14289,N_13513);
nor U16414 (N_16414,N_10343,N_10824);
or U16415 (N_16415,N_14114,N_12340);
and U16416 (N_16416,N_12414,N_13568);
or U16417 (N_16417,N_11642,N_12354);
and U16418 (N_16418,N_11681,N_10893);
nor U16419 (N_16419,N_13867,N_11795);
xor U16420 (N_16420,N_14304,N_14966);
xor U16421 (N_16421,N_14994,N_10292);
xor U16422 (N_16422,N_13683,N_11206);
and U16423 (N_16423,N_10927,N_12807);
nand U16424 (N_16424,N_13448,N_12254);
nor U16425 (N_16425,N_13287,N_14649);
or U16426 (N_16426,N_10817,N_14701);
and U16427 (N_16427,N_11449,N_13855);
and U16428 (N_16428,N_10213,N_14021);
nand U16429 (N_16429,N_11105,N_12608);
or U16430 (N_16430,N_13869,N_13537);
and U16431 (N_16431,N_13075,N_14926);
nand U16432 (N_16432,N_14117,N_13382);
and U16433 (N_16433,N_12566,N_13143);
nor U16434 (N_16434,N_10158,N_11076);
nor U16435 (N_16435,N_13887,N_10498);
xnor U16436 (N_16436,N_11979,N_14805);
nand U16437 (N_16437,N_13674,N_11548);
xor U16438 (N_16438,N_14089,N_13061);
xor U16439 (N_16439,N_14093,N_13758);
or U16440 (N_16440,N_13319,N_13761);
nand U16441 (N_16441,N_14816,N_11181);
or U16442 (N_16442,N_12337,N_13418);
and U16443 (N_16443,N_10076,N_13214);
nand U16444 (N_16444,N_12455,N_14947);
nor U16445 (N_16445,N_13197,N_14335);
and U16446 (N_16446,N_12201,N_12985);
nand U16447 (N_16447,N_12942,N_14661);
and U16448 (N_16448,N_12127,N_10504);
nand U16449 (N_16449,N_10531,N_13917);
nand U16450 (N_16450,N_14970,N_10442);
nor U16451 (N_16451,N_11392,N_14908);
or U16452 (N_16452,N_12672,N_10230);
xnor U16453 (N_16453,N_12389,N_14264);
nand U16454 (N_16454,N_13525,N_13543);
or U16455 (N_16455,N_10120,N_10294);
nand U16456 (N_16456,N_11269,N_13589);
or U16457 (N_16457,N_14787,N_13213);
nor U16458 (N_16458,N_14813,N_13514);
or U16459 (N_16459,N_13120,N_12171);
or U16460 (N_16460,N_13420,N_12905);
or U16461 (N_16461,N_13988,N_12189);
xnor U16462 (N_16462,N_11887,N_13013);
and U16463 (N_16463,N_14368,N_14261);
and U16464 (N_16464,N_14011,N_10600);
nand U16465 (N_16465,N_10147,N_10593);
nor U16466 (N_16466,N_12087,N_11341);
and U16467 (N_16467,N_12908,N_14439);
nor U16468 (N_16468,N_14544,N_14155);
nor U16469 (N_16469,N_13080,N_11634);
or U16470 (N_16470,N_10096,N_14829);
or U16471 (N_16471,N_11983,N_14896);
xnor U16472 (N_16472,N_11948,N_13517);
nand U16473 (N_16473,N_10842,N_14736);
nor U16474 (N_16474,N_14386,N_13261);
or U16475 (N_16475,N_14422,N_12341);
nor U16476 (N_16476,N_11777,N_11018);
xnor U16477 (N_16477,N_12462,N_11999);
nand U16478 (N_16478,N_11481,N_10719);
and U16479 (N_16479,N_11200,N_14806);
or U16480 (N_16480,N_12493,N_10454);
or U16481 (N_16481,N_12438,N_12187);
xor U16482 (N_16482,N_14616,N_10389);
nand U16483 (N_16483,N_14221,N_10731);
nand U16484 (N_16484,N_14999,N_13975);
xnor U16485 (N_16485,N_11472,N_11068);
nand U16486 (N_16486,N_13035,N_12859);
and U16487 (N_16487,N_10710,N_14367);
and U16488 (N_16488,N_11598,N_10700);
nand U16489 (N_16489,N_14349,N_13566);
xor U16490 (N_16490,N_12519,N_12398);
xor U16491 (N_16491,N_11065,N_11512);
nor U16492 (N_16492,N_13062,N_14005);
and U16493 (N_16493,N_14882,N_13315);
or U16494 (N_16494,N_12350,N_10975);
xnor U16495 (N_16495,N_12084,N_11097);
and U16496 (N_16496,N_14190,N_14152);
nor U16497 (N_16497,N_14319,N_13581);
nand U16498 (N_16498,N_13923,N_11682);
or U16499 (N_16499,N_11755,N_11915);
or U16500 (N_16500,N_10573,N_14070);
or U16501 (N_16501,N_14892,N_13072);
nor U16502 (N_16502,N_11107,N_14257);
or U16503 (N_16503,N_13704,N_13849);
xor U16504 (N_16504,N_14697,N_11941);
xor U16505 (N_16505,N_12537,N_12366);
and U16506 (N_16506,N_13227,N_11464);
or U16507 (N_16507,N_10409,N_12588);
and U16508 (N_16508,N_14270,N_11698);
xnor U16509 (N_16509,N_13459,N_14886);
nor U16510 (N_16510,N_13376,N_12694);
or U16511 (N_16511,N_11069,N_10752);
and U16512 (N_16512,N_11290,N_10974);
or U16513 (N_16513,N_10799,N_13911);
nand U16514 (N_16514,N_10310,N_12920);
or U16515 (N_16515,N_12241,N_12125);
nand U16516 (N_16516,N_13084,N_13863);
xor U16517 (N_16517,N_10253,N_14330);
and U16518 (N_16518,N_12560,N_13610);
xnor U16519 (N_16519,N_13731,N_10334);
or U16520 (N_16520,N_11619,N_11986);
nor U16521 (N_16521,N_12274,N_14745);
xor U16522 (N_16522,N_11876,N_12585);
nand U16523 (N_16523,N_13164,N_13421);
nand U16524 (N_16524,N_13449,N_13386);
nand U16525 (N_16525,N_10037,N_10588);
nor U16526 (N_16526,N_12159,N_11429);
nor U16527 (N_16527,N_11038,N_14493);
or U16528 (N_16528,N_12302,N_12632);
nor U16529 (N_16529,N_10701,N_14331);
nand U16530 (N_16530,N_12070,N_11294);
or U16531 (N_16531,N_11321,N_13276);
nor U16532 (N_16532,N_10729,N_10227);
nor U16533 (N_16533,N_10853,N_11494);
or U16534 (N_16534,N_14110,N_12259);
nand U16535 (N_16535,N_11821,N_11605);
or U16536 (N_16536,N_10580,N_12635);
and U16537 (N_16537,N_13845,N_11759);
nand U16538 (N_16538,N_11245,N_12113);
nor U16539 (N_16539,N_12351,N_11334);
nand U16540 (N_16540,N_13032,N_14471);
nor U16541 (N_16541,N_11034,N_13647);
xnor U16542 (N_16542,N_14456,N_11058);
or U16543 (N_16543,N_12625,N_14377);
and U16544 (N_16544,N_13461,N_13339);
or U16545 (N_16545,N_13715,N_10759);
nor U16546 (N_16546,N_14303,N_14213);
nor U16547 (N_16547,N_10171,N_11077);
nor U16548 (N_16548,N_13663,N_11405);
xnor U16549 (N_16549,N_10234,N_14874);
and U16550 (N_16550,N_10424,N_11159);
nand U16551 (N_16551,N_14899,N_14774);
and U16552 (N_16552,N_14595,N_14085);
nor U16553 (N_16553,N_12811,N_11433);
nand U16554 (N_16554,N_13004,N_11890);
and U16555 (N_16555,N_14124,N_12242);
xor U16556 (N_16556,N_12953,N_14988);
or U16557 (N_16557,N_10385,N_14730);
nand U16558 (N_16558,N_11400,N_10440);
xnor U16559 (N_16559,N_10804,N_10660);
xnor U16560 (N_16560,N_14884,N_11726);
xor U16561 (N_16561,N_11438,N_14568);
nand U16562 (N_16562,N_12481,N_10812);
nand U16563 (N_16563,N_13681,N_12834);
or U16564 (N_16564,N_14955,N_10005);
nand U16565 (N_16565,N_11466,N_10450);
nand U16566 (N_16566,N_14313,N_14184);
nor U16567 (N_16567,N_12680,N_10617);
or U16568 (N_16568,N_13773,N_13172);
xnor U16569 (N_16569,N_11894,N_13282);
or U16570 (N_16570,N_13336,N_13440);
nand U16571 (N_16571,N_11637,N_13292);
nand U16572 (N_16572,N_10630,N_14465);
or U16573 (N_16573,N_13158,N_13882);
nor U16574 (N_16574,N_10720,N_13624);
nand U16575 (N_16575,N_11752,N_12474);
xnor U16576 (N_16576,N_11149,N_12003);
xnor U16577 (N_16577,N_13832,N_12184);
and U16578 (N_16578,N_14913,N_11616);
nand U16579 (N_16579,N_14427,N_13531);
nand U16580 (N_16580,N_11259,N_13739);
or U16581 (N_16581,N_10793,N_13060);
nand U16582 (N_16582,N_11379,N_13607);
nand U16583 (N_16583,N_14414,N_12207);
nand U16584 (N_16584,N_14881,N_11942);
nor U16585 (N_16585,N_12833,N_11655);
nor U16586 (N_16586,N_12294,N_13876);
xor U16587 (N_16587,N_12568,N_14443);
and U16588 (N_16588,N_10095,N_12251);
nand U16589 (N_16589,N_13019,N_13149);
nor U16590 (N_16590,N_12888,N_12129);
nor U16591 (N_16591,N_11394,N_12541);
xor U16592 (N_16592,N_14244,N_10092);
nand U16593 (N_16593,N_11309,N_11182);
xnor U16594 (N_16594,N_11793,N_12765);
or U16595 (N_16595,N_11441,N_12227);
or U16596 (N_16596,N_13518,N_14674);
xor U16597 (N_16597,N_11497,N_14508);
nand U16598 (N_16598,N_10082,N_10427);
nor U16599 (N_16599,N_12949,N_11231);
and U16600 (N_16600,N_14446,N_11950);
xor U16601 (N_16601,N_12373,N_14272);
or U16602 (N_16602,N_11211,N_12024);
or U16603 (N_16603,N_13469,N_13498);
xnor U16604 (N_16604,N_11833,N_14715);
xor U16605 (N_16605,N_12409,N_14268);
nor U16606 (N_16606,N_12936,N_11388);
xor U16607 (N_16607,N_13497,N_14795);
or U16608 (N_16608,N_13981,N_12491);
nor U16609 (N_16609,N_11262,N_10359);
or U16610 (N_16610,N_13471,N_10977);
nor U16611 (N_16611,N_12520,N_13808);
xnor U16612 (N_16612,N_13853,N_10727);
or U16613 (N_16613,N_14713,N_10970);
and U16614 (N_16614,N_13026,N_10127);
nand U16615 (N_16615,N_12558,N_13840);
or U16616 (N_16616,N_14199,N_12176);
or U16617 (N_16617,N_10399,N_14052);
nor U16618 (N_16618,N_12081,N_14948);
or U16619 (N_16619,N_12634,N_12343);
xor U16620 (N_16620,N_10859,N_12621);
xor U16621 (N_16621,N_13748,N_12602);
or U16622 (N_16622,N_10132,N_10219);
and U16623 (N_16623,N_11349,N_11291);
xnor U16624 (N_16624,N_14605,N_13110);
nor U16625 (N_16625,N_10652,N_13124);
nor U16626 (N_16626,N_10029,N_11006);
and U16627 (N_16627,N_14692,N_10148);
nand U16628 (N_16628,N_10965,N_11420);
or U16629 (N_16629,N_14405,N_13325);
nand U16630 (N_16630,N_11865,N_10469);
nand U16631 (N_16631,N_14312,N_12530);
nand U16632 (N_16632,N_11955,N_14448);
nor U16633 (N_16633,N_14983,N_11909);
or U16634 (N_16634,N_12801,N_10070);
nor U16635 (N_16635,N_10116,N_14276);
or U16636 (N_16636,N_14285,N_14163);
or U16637 (N_16637,N_12420,N_10826);
and U16638 (N_16638,N_14046,N_11844);
nand U16639 (N_16639,N_13086,N_10598);
and U16640 (N_16640,N_12399,N_13322);
nor U16641 (N_16641,N_11668,N_14585);
nand U16642 (N_16642,N_10708,N_10613);
nand U16643 (N_16643,N_10560,N_12959);
nand U16644 (N_16644,N_13088,N_12311);
and U16645 (N_16645,N_12048,N_10223);
nor U16646 (N_16646,N_13577,N_11730);
nand U16647 (N_16647,N_13569,N_12447);
nand U16648 (N_16648,N_11037,N_11633);
nor U16649 (N_16649,N_11253,N_13241);
nor U16650 (N_16650,N_13310,N_10951);
nand U16651 (N_16651,N_13844,N_14207);
xor U16652 (N_16652,N_13783,N_12775);
or U16653 (N_16653,N_12425,N_11162);
or U16654 (N_16654,N_11957,N_14980);
nor U16655 (N_16655,N_14923,N_14337);
and U16656 (N_16656,N_14538,N_11251);
and U16657 (N_16657,N_10950,N_13733);
nor U16658 (N_16658,N_14150,N_11505);
and U16659 (N_16659,N_11160,N_14690);
or U16660 (N_16660,N_11426,N_10657);
nand U16661 (N_16661,N_11837,N_12831);
xnor U16662 (N_16662,N_13374,N_10684);
and U16663 (N_16663,N_14228,N_11196);
xor U16664 (N_16664,N_10097,N_12009);
or U16665 (N_16665,N_14020,N_14075);
nor U16666 (N_16666,N_14379,N_11218);
and U16667 (N_16667,N_13332,N_14402);
or U16668 (N_16668,N_12134,N_11122);
xor U16669 (N_16669,N_12269,N_10032);
nor U16670 (N_16670,N_11886,N_10586);
or U16671 (N_16671,N_11900,N_11626);
nand U16672 (N_16672,N_11046,N_14084);
nor U16673 (N_16673,N_11027,N_11150);
xnor U16674 (N_16674,N_11773,N_12601);
xnor U16675 (N_16675,N_13812,N_11963);
xor U16676 (N_16676,N_10993,N_13679);
xor U16677 (N_16677,N_11764,N_12278);
or U16678 (N_16678,N_12698,N_12670);
or U16679 (N_16679,N_13361,N_10664);
nand U16680 (N_16680,N_11602,N_11089);
or U16681 (N_16681,N_13848,N_13198);
nor U16682 (N_16682,N_12967,N_12858);
and U16683 (N_16683,N_12676,N_11660);
or U16684 (N_16684,N_12697,N_10761);
nor U16685 (N_16685,N_14663,N_14078);
and U16686 (N_16686,N_12273,N_11798);
nand U16687 (N_16687,N_13231,N_12964);
or U16688 (N_16688,N_10118,N_14348);
nor U16689 (N_16689,N_13392,N_11304);
nand U16690 (N_16690,N_13837,N_10640);
nor U16691 (N_16691,N_10025,N_10104);
xor U16692 (N_16692,N_11312,N_12695);
or U16693 (N_16693,N_12469,N_12647);
xor U16694 (N_16694,N_13030,N_10411);
or U16695 (N_16695,N_11169,N_14733);
nand U16696 (N_16696,N_10472,N_10537);
nor U16697 (N_16697,N_12356,N_12015);
xor U16698 (N_16698,N_10647,N_10505);
and U16699 (N_16699,N_13089,N_11025);
xnor U16700 (N_16700,N_10955,N_13329);
nand U16701 (N_16701,N_13159,N_11778);
nand U16702 (N_16702,N_10061,N_14419);
or U16703 (N_16703,N_11135,N_10577);
and U16704 (N_16704,N_14290,N_14587);
and U16705 (N_16705,N_10854,N_10181);
and U16706 (N_16706,N_11280,N_12338);
and U16707 (N_16707,N_12039,N_13166);
and U16708 (N_16708,N_13916,N_14492);
nand U16709 (N_16709,N_14909,N_10549);
nor U16710 (N_16710,N_12416,N_10833);
nand U16711 (N_16711,N_14834,N_13608);
or U16712 (N_16712,N_11529,N_13640);
and U16713 (N_16713,N_13121,N_11049);
nor U16714 (N_16714,N_14861,N_14689);
or U16715 (N_16715,N_11487,N_12443);
xor U16716 (N_16716,N_13931,N_12370);
and U16717 (N_16717,N_10551,N_13541);
or U16718 (N_16718,N_12612,N_10287);
xor U16719 (N_16719,N_14167,N_11719);
and U16720 (N_16720,N_13597,N_11654);
nor U16721 (N_16721,N_12164,N_12898);
nand U16722 (N_16722,N_11819,N_12156);
xor U16723 (N_16723,N_10489,N_12109);
or U16724 (N_16724,N_13473,N_13602);
nor U16725 (N_16725,N_10164,N_10452);
and U16726 (N_16726,N_11344,N_10969);
nand U16727 (N_16727,N_10445,N_14350);
nor U16728 (N_16728,N_12075,N_13521);
and U16729 (N_16729,N_10671,N_14871);
nor U16730 (N_16730,N_14982,N_10406);
nand U16731 (N_16731,N_10093,N_14209);
nor U16732 (N_16732,N_11220,N_12433);
or U16733 (N_16733,N_10845,N_12490);
and U16734 (N_16734,N_10928,N_14507);
or U16735 (N_16735,N_12334,N_14900);
or U16736 (N_16736,N_10675,N_10838);
xor U16737 (N_16737,N_11818,N_11715);
or U16738 (N_16738,N_12626,N_13097);
or U16739 (N_16739,N_11841,N_10959);
nand U16740 (N_16740,N_14560,N_12419);
nor U16741 (N_16741,N_11203,N_14555);
xor U16742 (N_16742,N_13146,N_12708);
xor U16743 (N_16743,N_10322,N_12534);
xnor U16744 (N_16744,N_14694,N_12514);
and U16745 (N_16745,N_14621,N_13447);
and U16746 (N_16746,N_13294,N_10933);
xnor U16747 (N_16747,N_12010,N_12769);
nand U16748 (N_16748,N_11386,N_14079);
nand U16749 (N_16749,N_10488,N_14388);
nor U16750 (N_16750,N_13486,N_12406);
nand U16751 (N_16751,N_10416,N_13415);
and U16752 (N_16752,N_12291,N_11985);
nand U16753 (N_16753,N_14520,N_10995);
nand U16754 (N_16754,N_14949,N_10014);
or U16755 (N_16755,N_12639,N_13236);
or U16756 (N_16756,N_11905,N_11771);
or U16757 (N_16757,N_11131,N_13410);
xor U16758 (N_16758,N_13436,N_13646);
or U16759 (N_16759,N_13797,N_13552);
xnor U16760 (N_16760,N_11987,N_10214);
nor U16761 (N_16761,N_10268,N_11938);
and U16762 (N_16762,N_10285,N_12258);
and U16763 (N_16763,N_12523,N_12508);
and U16764 (N_16764,N_13642,N_13183);
and U16765 (N_16765,N_13859,N_10346);
or U16766 (N_16766,N_12576,N_14850);
nor U16767 (N_16767,N_11061,N_12903);
or U16768 (N_16768,N_10022,N_13304);
and U16769 (N_16769,N_14927,N_13263);
and U16770 (N_16770,N_14318,N_13659);
xnor U16771 (N_16771,N_12100,N_11772);
nand U16772 (N_16772,N_13770,N_13400);
nor U16773 (N_16773,N_11539,N_14639);
xnor U16774 (N_16774,N_14137,N_10202);
xnor U16775 (N_16775,N_13843,N_10126);
nand U16776 (N_16776,N_13116,N_10744);
nand U16777 (N_16777,N_11385,N_13586);
xor U16778 (N_16778,N_10963,N_13316);
or U16779 (N_16779,N_10040,N_10446);
and U16780 (N_16780,N_12377,N_12506);
and U16781 (N_16781,N_11208,N_11145);
nor U16782 (N_16782,N_11130,N_13267);
xnor U16783 (N_16783,N_11115,N_11776);
xnor U16784 (N_16784,N_14606,N_13186);
nand U16785 (N_16785,N_10672,N_10415);
and U16786 (N_16786,N_14398,N_11083);
and U16787 (N_16787,N_12265,N_11582);
xnor U16788 (N_16788,N_11216,N_13467);
and U16789 (N_16789,N_12825,N_11215);
xnor U16790 (N_16790,N_13087,N_14357);
nand U16791 (N_16791,N_12616,N_11927);
xor U16792 (N_16792,N_10851,N_14102);
and U16793 (N_16793,N_13956,N_11533);
or U16794 (N_16794,N_13335,N_13264);
nor U16795 (N_16795,N_12510,N_13639);
nor U16796 (N_16796,N_12012,N_13538);
nand U16797 (N_16797,N_11570,N_11559);
xnor U16798 (N_16798,N_13065,N_10525);
nand U16799 (N_16799,N_14978,N_14543);
nand U16800 (N_16800,N_11585,N_13460);
and U16801 (N_16801,N_10805,N_12742);
and U16802 (N_16802,N_13561,N_13596);
xor U16803 (N_16803,N_12262,N_10004);
xor U16804 (N_16804,N_13260,N_10176);
and U16805 (N_16805,N_11692,N_14406);
or U16806 (N_16806,N_12528,N_11461);
or U16807 (N_16807,N_11677,N_14622);
nor U16808 (N_16808,N_10984,N_14696);
and U16809 (N_16809,N_13858,N_11240);
nand U16810 (N_16810,N_13714,N_10236);
nand U16811 (N_16811,N_11806,N_11047);
xor U16812 (N_16812,N_13358,N_11008);
or U16813 (N_16813,N_12412,N_12225);
xnor U16814 (N_16814,N_11934,N_12175);
and U16815 (N_16815,N_13613,N_10850);
nor U16816 (N_16816,N_13377,N_12961);
or U16817 (N_16817,N_13428,N_11832);
xnor U16818 (N_16818,N_14944,N_14545);
xnor U16819 (N_16819,N_14064,N_11511);
nor U16820 (N_16820,N_11051,N_14259);
nand U16821 (N_16821,N_12627,N_10110);
and U16822 (N_16822,N_13908,N_11665);
nand U16823 (N_16823,N_12613,N_10585);
nor U16824 (N_16824,N_11780,N_11279);
or U16825 (N_16825,N_13570,N_10777);
nor U16826 (N_16826,N_12725,N_12824);
or U16827 (N_16827,N_12853,N_11643);
and U16828 (N_16828,N_14822,N_13865);
and U16829 (N_16829,N_14671,N_14359);
nor U16830 (N_16830,N_12342,N_11587);
or U16831 (N_16831,N_11606,N_10904);
nand U16832 (N_16832,N_11483,N_14934);
nor U16833 (N_16833,N_13343,N_12861);
xnor U16834 (N_16834,N_14188,N_11919);
and U16835 (N_16835,N_12718,N_13001);
and U16836 (N_16836,N_10034,N_11445);
or U16837 (N_16837,N_14345,N_12993);
nor U16838 (N_16838,N_12320,N_12925);
nor U16839 (N_16839,N_13193,N_14589);
xor U16840 (N_16840,N_10423,N_11223);
nor U16841 (N_16841,N_11432,N_14891);
nand U16842 (N_16842,N_13925,N_13347);
nand U16843 (N_16843,N_12219,N_11498);
nor U16844 (N_16844,N_11390,N_10888);
xnor U16845 (N_16845,N_14801,N_13049);
or U16846 (N_16846,N_11340,N_14710);
xnor U16847 (N_16847,N_12058,N_10421);
and U16848 (N_16848,N_14281,N_13833);
or U16849 (N_16849,N_14420,N_10583);
nor U16850 (N_16850,N_10733,N_14652);
or U16851 (N_16851,N_13082,N_11015);
and U16852 (N_16852,N_10682,N_11839);
or U16853 (N_16853,N_12753,N_14646);
xor U16854 (N_16854,N_10973,N_13595);
nand U16855 (N_16855,N_12486,N_11815);
xnor U16856 (N_16856,N_14157,N_12235);
nor U16857 (N_16857,N_10160,N_14411);
nand U16858 (N_16858,N_10931,N_12363);
and U16859 (N_16859,N_14432,N_14700);
xnor U16860 (N_16860,N_10896,N_13727);
nor U16861 (N_16861,N_13854,N_11736);
xor U16862 (N_16862,N_10496,N_14860);
nor U16863 (N_16863,N_10582,N_12266);
nor U16864 (N_16864,N_14474,N_13846);
nand U16865 (N_16865,N_14273,N_11910);
nor U16866 (N_16866,N_10881,N_13017);
nand U16867 (N_16867,N_12232,N_13643);
nand U16868 (N_16868,N_14397,N_13016);
nand U16869 (N_16869,N_10601,N_13196);
and U16870 (N_16870,N_12652,N_11536);
and U16871 (N_16871,N_11861,N_10159);
xnor U16872 (N_16872,N_11463,N_14851);
or U16873 (N_16873,N_12115,N_10766);
and U16874 (N_16874,N_13658,N_14108);
or U16875 (N_16875,N_12123,N_11178);
nor U16876 (N_16876,N_13927,N_12663);
nand U16877 (N_16877,N_11853,N_10510);
xor U16878 (N_16878,N_14171,N_10649);
nand U16879 (N_16879,N_12610,N_14491);
xnor U16880 (N_16880,N_11436,N_10041);
nand U16881 (N_16881,N_12256,N_14026);
and U16882 (N_16882,N_11274,N_11112);
xor U16883 (N_16883,N_13269,N_10428);
nand U16884 (N_16884,N_10578,N_11958);
or U16885 (N_16885,N_14169,N_13572);
or U16886 (N_16886,N_12536,N_10162);
nand U16887 (N_16887,N_10609,N_13982);
and U16888 (N_16888,N_13117,N_11656);
and U16889 (N_16889,N_11903,N_10885);
and U16890 (N_16890,N_11066,N_12597);
xor U16891 (N_16891,N_13990,N_10792);
xor U16892 (N_16892,N_12661,N_10669);
and U16893 (N_16893,N_10765,N_10718);
xnor U16894 (N_16894,N_12910,N_14725);
nor U16895 (N_16895,N_11120,N_10226);
nor U16896 (N_16896,N_11036,N_11153);
xor U16897 (N_16897,N_14638,N_11273);
xnor U16898 (N_16898,N_13165,N_12798);
or U16899 (N_16899,N_14626,N_12879);
xnor U16900 (N_16900,N_12381,N_10555);
and U16901 (N_16901,N_10524,N_14413);
nand U16902 (N_16902,N_10413,N_11395);
or U16903 (N_16903,N_12665,N_13195);
xnor U16904 (N_16904,N_12900,N_10323);
and U16905 (N_16905,N_11010,N_11828);
nand U16906 (N_16906,N_10275,N_11106);
nand U16907 (N_16907,N_12991,N_13104);
nor U16908 (N_16908,N_14484,N_13556);
and U16909 (N_16909,N_13998,N_11544);
nor U16910 (N_16910,N_10883,N_13632);
and U16911 (N_16911,N_13168,N_13816);
nand U16912 (N_16912,N_10785,N_13948);
or U16913 (N_16913,N_14920,N_13829);
nor U16914 (N_16914,N_12052,N_13046);
and U16915 (N_16915,N_14206,N_14288);
nor U16916 (N_16916,N_12850,N_10894);
or U16917 (N_16917,N_14455,N_11310);
nor U16918 (N_16918,N_10561,N_12880);
or U16919 (N_16919,N_12580,N_11968);
nand U16920 (N_16920,N_13781,N_12938);
or U16921 (N_16921,N_12773,N_12972);
nand U16922 (N_16922,N_10941,N_11874);
xnor U16923 (N_16923,N_13020,N_12847);
or U16924 (N_16924,N_11000,N_13458);
xor U16925 (N_16925,N_14672,N_14320);
nand U16926 (N_16926,N_10124,N_10130);
nor U16927 (N_16927,N_12556,N_11638);
nand U16928 (N_16928,N_10610,N_11857);
nor U16929 (N_16929,N_13371,N_12197);
nor U16930 (N_16930,N_11686,N_13439);
nor U16931 (N_16931,N_11572,N_10312);
nand U16932 (N_16932,N_10090,N_14045);
xor U16933 (N_16933,N_11275,N_12819);
and U16934 (N_16934,N_13464,N_11104);
xor U16935 (N_16935,N_13238,N_14910);
xnor U16936 (N_16936,N_14112,N_13657);
xnor U16937 (N_16937,N_11738,N_13606);
xnor U16938 (N_16938,N_12305,N_12494);
nor U16939 (N_16939,N_11266,N_14370);
xor U16940 (N_16940,N_11555,N_10098);
or U16941 (N_16941,N_11444,N_13246);
xnor U16942 (N_16942,N_12185,N_11520);
nand U16943 (N_16943,N_11912,N_11271);
nor U16944 (N_16944,N_11964,N_12060);
and U16945 (N_16945,N_11367,N_14855);
xnor U16946 (N_16946,N_13871,N_10430);
and U16947 (N_16947,N_11881,N_11484);
or U16948 (N_16948,N_14711,N_13698);
nor U16949 (N_16949,N_10172,N_10745);
nor U16950 (N_16950,N_12086,N_12284);
xnor U16951 (N_16951,N_13192,N_11748);
and U16952 (N_16952,N_10307,N_10724);
nand U16953 (N_16953,N_14863,N_10541);
xor U16954 (N_16954,N_11674,N_13777);
or U16955 (N_16955,N_10327,N_12954);
nand U16956 (N_16956,N_10828,N_10013);
nor U16957 (N_16957,N_13888,N_12660);
and U16958 (N_16958,N_10673,N_10808);
xnor U16959 (N_16959,N_11332,N_12656);
nor U16960 (N_16960,N_11452,N_13820);
nand U16961 (N_16961,N_13585,N_13952);
nand U16962 (N_16962,N_10386,N_10105);
nor U16963 (N_16963,N_10291,N_11099);
nand U16964 (N_16964,N_13027,N_14727);
nand U16965 (N_16965,N_14019,N_10569);
or U16966 (N_16966,N_10949,N_14341);
nor U16967 (N_16967,N_14853,N_10717);
nor U16968 (N_16968,N_11095,N_11561);
nand U16969 (N_16969,N_14372,N_10773);
nand U16970 (N_16970,N_13268,N_13934);
nor U16971 (N_16971,N_11490,N_11501);
nand U16972 (N_16972,N_13224,N_10764);
nor U16973 (N_16973,N_14731,N_12484);
xnor U16974 (N_16974,N_13554,N_14269);
and U16975 (N_16975,N_12830,N_14363);
nand U16976 (N_16976,N_11252,N_13488);
nand U16977 (N_16977,N_13966,N_14229);
or U16978 (N_16978,N_11904,N_10658);
and U16979 (N_16979,N_10278,N_10604);
nand U16980 (N_16980,N_12907,N_10290);
and U16981 (N_16981,N_10060,N_11308);
nor U16982 (N_16982,N_11096,N_11249);
or U16983 (N_16983,N_12309,N_12421);
nor U16984 (N_16984,N_11614,N_10509);
and U16985 (N_16985,N_11063,N_14198);
nand U16986 (N_16986,N_14120,N_14189);
and U16987 (N_16987,N_11541,N_14756);
or U16988 (N_16988,N_12153,N_10482);
nor U16989 (N_16989,N_12103,N_13134);
nand U16990 (N_16990,N_11817,N_12384);
and U16991 (N_16991,N_12397,N_10659);
nand U16992 (N_16992,N_10371,N_14656);
nand U16993 (N_16993,N_10271,N_10837);
nor U16994 (N_16994,N_12163,N_14526);
xor U16995 (N_16995,N_14546,N_13599);
and U16996 (N_16996,N_14362,N_14532);
nor U16997 (N_16997,N_10218,N_12349);
nand U16998 (N_16998,N_10436,N_10688);
and U16999 (N_16999,N_14975,N_10138);
nor U17000 (N_17000,N_12195,N_10387);
or U17001 (N_17001,N_13989,N_12312);
nand U17002 (N_17002,N_10676,N_10899);
or U17003 (N_17003,N_10363,N_10532);
xor U17004 (N_17004,N_14572,N_14984);
and U17005 (N_17005,N_11558,N_10426);
xor U17006 (N_17006,N_10677,N_13402);
nand U17007 (N_17007,N_13961,N_13939);
nor U17008 (N_17008,N_10905,N_10870);
or U17009 (N_17009,N_12657,N_10687);
nor U17010 (N_17010,N_10019,N_13131);
nor U17011 (N_17011,N_10467,N_11100);
nor U17012 (N_17012,N_12328,N_14047);
nand U17013 (N_17013,N_12715,N_10957);
xnor U17014 (N_17014,N_11994,N_11292);
nor U17015 (N_17015,N_12668,N_13220);
nand U17016 (N_17016,N_10515,N_13091);
or U17017 (N_17017,N_10550,N_11685);
nor U17018 (N_17018,N_11506,N_12666);
xnor U17019 (N_17019,N_13419,N_12581);
nor U17020 (N_17020,N_13575,N_10017);
nand U17021 (N_17021,N_14039,N_12642);
nor U17022 (N_17022,N_14309,N_12945);
nor U17023 (N_17023,N_14673,N_13037);
or U17024 (N_17024,N_14888,N_11998);
nand U17025 (N_17025,N_14859,N_10575);
nor U17026 (N_17026,N_11380,N_10477);
and U17027 (N_17027,N_12521,N_13547);
xnor U17028 (N_17028,N_13479,N_11972);
nand U17029 (N_17029,N_12533,N_12260);
or U17030 (N_17030,N_11189,N_10169);
or U17031 (N_17031,N_11822,N_10206);
and U17032 (N_17032,N_13710,N_11355);
or U17033 (N_17033,N_13969,N_13826);
nor U17034 (N_17034,N_11728,N_13993);
nand U17035 (N_17035,N_14917,N_11296);
nor U17036 (N_17036,N_13470,N_13171);
nor U17037 (N_17037,N_12150,N_13290);
nand U17038 (N_17038,N_13071,N_13130);
nor U17039 (N_17039,N_13847,N_14104);
nand U17040 (N_17040,N_11608,N_10326);
nand U17041 (N_17041,N_13804,N_10594);
xor U17042 (N_17042,N_10847,N_14074);
nand U17043 (N_17043,N_13430,N_12374);
xnor U17044 (N_17044,N_14769,N_11151);
xor U17045 (N_17045,N_10320,N_11476);
or U17046 (N_17046,N_11943,N_13814);
xor U17047 (N_17047,N_10046,N_11091);
and U17048 (N_17048,N_13423,N_11192);
nand U17049 (N_17049,N_12396,N_14201);
nand U17050 (N_17050,N_12930,N_11359);
or U17051 (N_17051,N_14043,N_12353);
nor U17052 (N_17052,N_10180,N_11768);
or U17053 (N_17053,N_13200,N_10261);
xor U17054 (N_17054,N_10222,N_12713);
or U17055 (N_17055,N_10351,N_14164);
nor U17056 (N_17056,N_14160,N_11966);
nand U17057 (N_17057,N_14648,N_10947);
and U17058 (N_17058,N_10412,N_13638);
nor U17059 (N_17059,N_12261,N_10536);
xnor U17060 (N_17060,N_10920,N_12173);
nor U17061 (N_17061,N_12118,N_13936);
xor U17062 (N_17062,N_13040,N_11669);
or U17063 (N_17063,N_12206,N_10862);
and U17064 (N_17064,N_14501,N_13852);
or U17065 (N_17065,N_11840,N_10705);
and U17066 (N_17066,N_12031,N_13113);
nor U17067 (N_17067,N_14235,N_10926);
nor U17068 (N_17068,N_12483,N_12402);
and U17069 (N_17069,N_13288,N_14741);
nand U17070 (N_17070,N_12360,N_13861);
nor U17071 (N_17071,N_14717,N_11201);
or U17072 (N_17072,N_14740,N_13705);
xnor U17073 (N_17073,N_12467,N_10141);
xor U17074 (N_17074,N_14848,N_14603);
and U17075 (N_17075,N_13690,N_11648);
or U17076 (N_17076,N_14178,N_12755);
xor U17077 (N_17077,N_12864,N_12068);
and U17078 (N_17078,N_12172,N_13254);
nand U17079 (N_17079,N_13483,N_14599);
nand U17080 (N_17080,N_13963,N_11094);
nand U17081 (N_17081,N_11854,N_10121);
xnor U17082 (N_17082,N_11947,N_12570);
and U17083 (N_17083,N_10645,N_10678);
nor U17084 (N_17084,N_12922,N_10175);
or U17085 (N_17085,N_13029,N_10706);
nor U17086 (N_17086,N_14620,N_12611);
or U17087 (N_17087,N_14973,N_10079);
nor U17088 (N_17088,N_11059,N_14103);
or U17089 (N_17089,N_11403,N_13818);
nor U17090 (N_17090,N_12693,N_12622);
or U17091 (N_17091,N_13477,N_12394);
xor U17092 (N_17092,N_14563,N_11210);
and U17093 (N_17093,N_12028,N_11242);
nor U17094 (N_17094,N_14315,N_13851);
or U17095 (N_17095,N_13102,N_10916);
xnor U17096 (N_17096,N_10709,N_10697);
nor U17097 (N_17097,N_12750,N_12951);
or U17098 (N_17098,N_11142,N_12946);
or U17099 (N_17099,N_12866,N_10099);
and U17100 (N_17100,N_11745,N_10711);
nand U17101 (N_17101,N_12116,N_13207);
or U17102 (N_17102,N_12155,N_12531);
nor U17103 (N_17103,N_12500,N_12391);
or U17104 (N_17104,N_10919,N_11255);
or U17105 (N_17105,N_11949,N_14301);
nand U17106 (N_17106,N_12029,N_12002);
and U17107 (N_17107,N_11700,N_12976);
nand U17108 (N_17108,N_13397,N_10419);
or U17109 (N_17109,N_13151,N_11005);
xor U17110 (N_17110,N_11138,N_13226);
xnor U17111 (N_17111,N_11373,N_10078);
xor U17112 (N_17112,N_11414,N_10224);
nor U17113 (N_17113,N_12685,N_13177);
nand U17114 (N_17114,N_14516,N_14481);
and U17115 (N_17115,N_14271,N_10775);
and U17116 (N_17116,N_11254,N_10051);
nand U17117 (N_17117,N_14936,N_14883);
xnor U17118 (N_17118,N_11961,N_12089);
or U17119 (N_17119,N_11261,N_13673);
nand U17120 (N_17120,N_10794,N_12881);
or U17121 (N_17121,N_11914,N_11766);
xnor U17122 (N_17122,N_10898,N_13929);
nor U17123 (N_17123,N_14051,N_10522);
nand U17124 (N_17124,N_14173,N_12330);
xor U17125 (N_17125,N_10434,N_10781);
nor U17126 (N_17126,N_13583,N_14498);
nor U17127 (N_17127,N_13873,N_12943);
xor U17128 (N_17128,N_12983,N_13558);
xnor U17129 (N_17129,N_13266,N_10266);
nand U17130 (N_17130,N_13813,N_12856);
and U17131 (N_17131,N_12901,N_14601);
xnor U17132 (N_17132,N_11315,N_11233);
or U17133 (N_17133,N_11788,N_11761);
and U17134 (N_17134,N_12686,N_12971);
and U17135 (N_17135,N_13070,N_11398);
and U17136 (N_17136,N_12000,N_10021);
and U17137 (N_17137,N_10247,N_10390);
nand U17138 (N_17138,N_13167,N_13375);
nor U17139 (N_17139,N_11975,N_12436);
or U17140 (N_17140,N_10470,N_12517);
xnor U17141 (N_17141,N_10703,N_14528);
nand U17142 (N_17142,N_14017,N_14961);
and U17143 (N_17143,N_12667,N_12575);
nand U17144 (N_17144,N_10402,N_14706);
nor U17145 (N_17145,N_10940,N_10563);
nand U17146 (N_17146,N_11239,N_11434);
and U17147 (N_17147,N_11043,N_14937);
and U17148 (N_17148,N_13669,N_14343);
nor U17149 (N_17149,N_13148,N_14785);
xor U17150 (N_17150,N_10783,N_11743);
and U17151 (N_17151,N_12445,N_14972);
nand U17152 (N_17152,N_14723,N_11858);
xnor U17153 (N_17153,N_12970,N_14338);
nor U17154 (N_17154,N_13895,N_13364);
xor U17155 (N_17155,N_14407,N_12784);
nor U17156 (N_17156,N_11475,N_13429);
or U17157 (N_17157,N_12649,N_10633);
nand U17158 (N_17158,N_11204,N_14371);
or U17159 (N_17159,N_11118,N_10332);
xnor U17160 (N_17160,N_14789,N_13868);
or U17161 (N_17161,N_11593,N_12378);
nand U17162 (N_17162,N_10663,N_13605);
nor U17163 (N_17163,N_12704,N_10086);
xor U17164 (N_17164,N_14773,N_13534);
or U17165 (N_17165,N_13281,N_14509);
or U17166 (N_17166,N_13676,N_13629);
nand U17167 (N_17167,N_11566,N_14709);
nor U17168 (N_17168,N_14100,N_12357);
nor U17169 (N_17169,N_14915,N_13408);
nor U17170 (N_17170,N_11578,N_14962);
and U17171 (N_17171,N_12603,N_12308);
and U17172 (N_17172,N_14895,N_14735);
or U17173 (N_17173,N_14009,N_14347);
xnor U17174 (N_17174,N_11442,N_10836);
and U17175 (N_17175,N_11356,N_13696);
or U17176 (N_17176,N_12287,N_11789);
or U17177 (N_17177,N_10125,N_13076);
xor U17178 (N_17178,N_11644,N_13821);
and U17179 (N_17179,N_10559,N_14094);
nor U17180 (N_17180,N_11225,N_10880);
and U17181 (N_17181,N_10233,N_11640);
or U17182 (N_17182,N_13373,N_14428);
and U17183 (N_17183,N_14489,N_13947);
nand U17184 (N_17184,N_12911,N_13564);
and U17185 (N_17185,N_14683,N_13141);
or U17186 (N_17186,N_13173,N_11884);
nand U17187 (N_17187,N_12886,N_12572);
nand U17188 (N_17188,N_11113,N_11830);
or U17189 (N_17189,N_12020,N_10157);
nor U17190 (N_17190,N_12417,N_10591);
nand U17191 (N_17191,N_14382,N_12347);
nand U17192 (N_17192,N_13603,N_13496);
or U17193 (N_17193,N_11276,N_10370);
nor U17194 (N_17194,N_13455,N_11217);
nor U17195 (N_17195,N_13985,N_14300);
nor U17196 (N_17196,N_14578,N_11732);
nor U17197 (N_17197,N_14556,N_11589);
nor U17198 (N_17198,N_12709,N_13933);
and U17199 (N_17199,N_13810,N_13502);
nor U17200 (N_17200,N_12368,N_11293);
xor U17201 (N_17201,N_13285,N_10865);
and U17202 (N_17202,N_11228,N_12835);
xnor U17203 (N_17203,N_11338,N_13986);
and U17204 (N_17204,N_14096,N_14719);
and U17205 (N_17205,N_14531,N_12659);
and U17206 (N_17206,N_14565,N_11283);
nor U17207 (N_17207,N_10597,N_10654);
and U17208 (N_17208,N_12527,N_13191);
nor U17209 (N_17209,N_11357,N_10945);
or U17210 (N_17210,N_13234,N_10258);
and U17211 (N_17211,N_13100,N_11437);
or U17212 (N_17212,N_10526,N_11382);
or U17213 (N_17213,N_11824,N_14297);
and U17214 (N_17214,N_14115,N_12329);
xnor U17215 (N_17215,N_10135,N_14530);
or U17216 (N_17216,N_14016,N_14591);
or U17217 (N_17217,N_14460,N_13515);
nand U17218 (N_17218,N_10252,N_10081);
nand U17219 (N_17219,N_12090,N_11923);
or U17220 (N_17220,N_14365,N_14869);
and U17221 (N_17221,N_13279,N_13527);
nor U17222 (N_17222,N_13791,N_12135);
and U17223 (N_17223,N_11899,N_11397);
nand U17224 (N_17224,N_11055,N_13532);
xnor U17225 (N_17225,N_14623,N_12035);
nor U17226 (N_17226,N_13991,N_13135);
nand U17227 (N_17227,N_13655,N_11087);
or U17228 (N_17228,N_10360,N_10330);
or U17229 (N_17229,N_13427,N_10344);
nand U17230 (N_17230,N_10849,N_10010);
and U17231 (N_17231,N_10342,N_12410);
and U17232 (N_17232,N_14873,N_10592);
xnor U17233 (N_17233,N_12304,N_12061);
nor U17234 (N_17234,N_13949,N_14292);
or U17235 (N_17235,N_14618,N_12280);
nand U17236 (N_17236,N_11418,N_13077);
nand U17237 (N_17237,N_12662,N_11435);
nor U17238 (N_17238,N_13125,N_14490);
or U17239 (N_17239,N_14952,N_12318);
nand U17240 (N_17240,N_11408,N_10248);
and U17241 (N_17241,N_10690,N_10075);
xor U17242 (N_17242,N_12995,N_11430);
nor U17243 (N_17243,N_12787,N_14251);
nand U17244 (N_17244,N_10844,N_13860);
nand U17245 (N_17245,N_12027,N_12631);
nor U17246 (N_17246,N_14352,N_13928);
or U17247 (N_17247,N_12624,N_10194);
nor U17248 (N_17248,N_12041,N_11003);
xnor U17249 (N_17249,N_13051,N_14416);
and U17250 (N_17250,N_11980,N_10778);
or U17251 (N_17251,N_12829,N_12314);
or U17252 (N_17252,N_11851,N_14783);
and U17253 (N_17253,N_10167,N_13170);
and U17254 (N_17254,N_11885,N_12088);
xnor U17255 (N_17255,N_12707,N_10570);
xor U17256 (N_17256,N_12170,N_13651);
or U17257 (N_17257,N_10934,N_11307);
nand U17258 (N_17258,N_13886,N_12054);
or U17259 (N_17259,N_13522,N_14750);
xor U17260 (N_17260,N_14239,N_10050);
xor U17261 (N_17261,N_13743,N_13972);
nand U17262 (N_17262,N_11336,N_10074);
and U17263 (N_17263,N_10168,N_10335);
or U17264 (N_17264,N_14059,N_14286);
nor U17265 (N_17265,N_12772,N_12228);
and U17266 (N_17266,N_13302,N_14366);
xnor U17267 (N_17267,N_10692,N_10207);
and U17268 (N_17268,N_13257,N_14527);
nor U17269 (N_17269,N_10556,N_11845);
or U17270 (N_17270,N_10487,N_13478);
nand U17271 (N_17271,N_13489,N_10491);
or U17272 (N_17272,N_11221,N_13163);
xor U17273 (N_17273,N_12785,N_10769);
or U17274 (N_17274,N_11928,N_11155);
and U17275 (N_17275,N_14220,N_10189);
xnor U17276 (N_17276,N_11174,N_12503);
and U17277 (N_17277,N_13786,N_12554);
or U17278 (N_17278,N_14200,N_12818);
xnor U17279 (N_17279,N_10356,N_14036);
xnor U17280 (N_17280,N_14981,N_11560);
or U17281 (N_17281,N_11368,N_12297);
nand U17282 (N_17282,N_12754,N_12026);
nand U17283 (N_17283,N_12595,N_11108);
and U17284 (N_17284,N_12095,N_13162);
nor U17285 (N_17285,N_10492,N_12428);
xor U17286 (N_17286,N_13251,N_10495);
or U17287 (N_17287,N_14050,N_11074);
and U17288 (N_17288,N_12149,N_11693);
and U17289 (N_17289,N_12933,N_12896);
nand U17290 (N_17290,N_13718,N_10122);
xnor U17291 (N_17291,N_13701,N_13006);
and U17292 (N_17292,N_12025,N_11579);
or U17293 (N_17293,N_11285,N_13244);
nand U17294 (N_17294,N_14476,N_11053);
or U17295 (N_17295,N_13495,N_12979);
or U17296 (N_17296,N_13487,N_13697);
or U17297 (N_17297,N_12840,N_13670);
and U17298 (N_17298,N_13431,N_10024);
nor U17299 (N_17299,N_11446,N_11495);
nand U17300 (N_17300,N_12074,N_10986);
nor U17301 (N_17301,N_14081,N_11295);
nand U17302 (N_17302,N_11439,N_14035);
nand U17303 (N_17303,N_11989,N_14794);
xor U17304 (N_17304,N_14473,N_11594);
xnor U17305 (N_17305,N_14467,N_13306);
xnor U17306 (N_17306,N_13946,N_12538);
and U17307 (N_17307,N_10867,N_12987);
nor U17308 (N_17308,N_14424,N_14729);
nand U17309 (N_17309,N_10800,N_12236);
nand U17310 (N_17310,N_10315,N_13205);
nand U17311 (N_17311,N_11205,N_10485);
nand U17312 (N_17312,N_11493,N_12385);
nor U17313 (N_17313,N_12131,N_10212);
and U17314 (N_17314,N_11032,N_11864);
xor U17315 (N_17315,N_11922,N_14380);
nor U17316 (N_17316,N_14233,N_10199);
nor U17317 (N_17317,N_13187,N_12800);
and U17318 (N_17318,N_11202,N_14746);
nor U17319 (N_17319,N_10077,N_12255);
and U17320 (N_17320,N_13811,N_12522);
nor U17321 (N_17321,N_13230,N_12756);
nand U17322 (N_17322,N_12112,N_14175);
nor U17323 (N_17323,N_11787,N_11303);
nand U17324 (N_17324,N_13472,N_14919);
or U17325 (N_17325,N_10796,N_12855);
and U17326 (N_17326,N_14630,N_14469);
or U17327 (N_17327,N_10596,N_11945);
nand U17328 (N_17328,N_11843,N_12711);
nand U17329 (N_17329,N_14356,N_11364);
or U17330 (N_17330,N_11161,N_10432);
nand U17331 (N_17331,N_11419,N_10185);
or U17332 (N_17332,N_13109,N_10608);
nor U17333 (N_17333,N_12738,N_11847);
and U17334 (N_17334,N_10512,N_13232);
nand U17335 (N_17335,N_12361,N_13066);
or U17336 (N_17336,N_11954,N_13750);
or U17337 (N_17337,N_13717,N_14158);
nor U17338 (N_17338,N_13360,N_13188);
xor U17339 (N_17339,N_11137,N_14945);
and U17340 (N_17340,N_14279,N_11479);
or U17341 (N_17341,N_12578,N_12689);
or U17342 (N_17342,N_14355,N_13950);
or U17343 (N_17343,N_11552,N_14786);
or U17344 (N_17344,N_12816,N_11871);
or U17345 (N_17345,N_12275,N_10295);
and U17346 (N_17346,N_12615,N_11062);
xnor U17347 (N_17347,N_13383,N_13252);
or U17348 (N_17348,N_14192,N_14702);
or U17349 (N_17349,N_13333,N_11683);
and U17350 (N_17350,N_13270,N_10400);
or U17351 (N_17351,N_12270,N_13805);
or U17352 (N_17352,N_10242,N_11712);
nand U17353 (N_17353,N_14283,N_10679);
xor U17354 (N_17354,N_13623,N_10357);
xnor U17355 (N_17355,N_12034,N_13598);
xor U17356 (N_17356,N_11453,N_12179);
nand U17357 (N_17357,N_13870,N_10544);
xor U17358 (N_17358,N_11193,N_11709);
or U17359 (N_17359,N_12651,N_13967);
or U17360 (N_17360,N_13578,N_11170);
nand U17361 (N_17361,N_10822,N_12884);
or U17362 (N_17362,N_12802,N_10642);
and U17363 (N_17363,N_13011,N_13732);
xnor U17364 (N_17364,N_14141,N_11537);
and U17365 (N_17365,N_11996,N_11535);
nand U17366 (N_17366,N_11509,N_11423);
and U17367 (N_17367,N_13275,N_10177);
or U17368 (N_17368,N_12728,N_14479);
and U17369 (N_17369,N_14759,N_11337);
nor U17370 (N_17370,N_11742,N_11389);
or U17371 (N_17371,N_10576,N_12393);
nor U17372 (N_17372,N_14800,N_12895);
nand U17373 (N_17373,N_11875,N_14996);
or U17374 (N_17374,N_14667,N_11820);
nor U17375 (N_17375,N_14361,N_14351);
nor U17376 (N_17376,N_12518,N_14569);
xnor U17377 (N_17377,N_11468,N_12072);
nand U17378 (N_17378,N_13799,N_10644);
or U17379 (N_17379,N_11019,N_10437);
or U17380 (N_17380,N_13828,N_10948);
and U17381 (N_17381,N_14845,N_14976);
xnor U17382 (N_17382,N_11946,N_14902);
nand U17383 (N_17383,N_10913,N_14651);
nand U17384 (N_17384,N_14230,N_11673);
nand U17385 (N_17385,N_10231,N_12339);
and U17386 (N_17386,N_12272,N_11411);
nor U17387 (N_17387,N_10474,N_13918);
or U17388 (N_17388,N_10183,N_13600);
or U17389 (N_17389,N_11907,N_11268);
and U17390 (N_17390,N_10038,N_14408);
nand U17391 (N_17391,N_14536,N_14828);
nand U17392 (N_17392,N_12904,N_10605);
or U17393 (N_17393,N_13817,N_13913);
xnor U17394 (N_17394,N_10698,N_11030);
xor U17395 (N_17395,N_13284,N_10289);
nor U17396 (N_17396,N_14645,N_10151);
or U17397 (N_17397,N_10702,N_14553);
nor U17398 (N_17398,N_11930,N_11073);
or U17399 (N_17399,N_11978,N_13898);
or U17400 (N_17400,N_12762,N_10810);
and U17401 (N_17401,N_14265,N_12717);
and U17402 (N_17402,N_10235,N_11026);
nand U17403 (N_17403,N_12692,N_11575);
or U17404 (N_17404,N_11194,N_10145);
nor U17405 (N_17405,N_13233,N_12246);
nor U17406 (N_17406,N_10887,N_10666);
and U17407 (N_17407,N_11524,N_10139);
nand U17408 (N_17408,N_13500,N_11119);
or U17409 (N_17409,N_11513,N_14575);
nor U17410 (N_17410,N_12923,N_14957);
nor U17411 (N_17411,N_12083,N_14847);
or U17412 (N_17412,N_12263,N_14742);
and U17413 (N_17413,N_12222,N_14979);
xnor U17414 (N_17414,N_10422,N_10460);
xnor U17415 (N_17415,N_11908,N_10302);
nor U17416 (N_17416,N_10448,N_10846);
and U17417 (N_17417,N_14166,N_13877);
and U17418 (N_17418,N_11735,N_10059);
xnor U17419 (N_17419,N_12196,N_13334);
nor U17420 (N_17420,N_13150,N_10897);
nand U17421 (N_17421,N_14222,N_13970);
and U17422 (N_17422,N_13003,N_10089);
and U17423 (N_17423,N_14191,N_13878);
xor U17424 (N_17424,N_12102,N_10429);
xnor U17425 (N_17425,N_13462,N_14342);
or U17426 (N_17426,N_11929,N_12037);
xnor U17427 (N_17427,N_10742,N_10911);
nand U17428 (N_17428,N_13622,N_10968);
xnor U17429 (N_17429,N_12057,N_10299);
nor U17430 (N_17430,N_12714,N_13722);
nor U17431 (N_17431,N_10795,N_12502);
xnor U17432 (N_17432,N_12319,N_12492);
and U17433 (N_17433,N_13740,N_13666);
nor U17434 (N_17434,N_13157,N_14614);
xnor U17435 (N_17435,N_14625,N_14549);
xnor U17436 (N_17436,N_13706,N_10798);
and U17437 (N_17437,N_11786,N_14720);
nor U17438 (N_17438,N_14765,N_11163);
nand U17439 (N_17439,N_13899,N_10023);
or U17440 (N_17440,N_10192,N_13668);
and U17441 (N_17441,N_14242,N_11136);
or U17442 (N_17442,N_12916,N_13433);
or U17443 (N_17443,N_14060,N_14231);
or U17444 (N_17444,N_14739,N_13484);
and U17445 (N_17445,N_14204,N_10481);
nand U17446 (N_17446,N_11482,N_13381);
and U17447 (N_17447,N_13094,N_11917);
and U17448 (N_17448,N_12362,N_14877);
or U17449 (N_17449,N_14610,N_12435);
or U17450 (N_17450,N_11407,N_11002);
nand U17451 (N_17451,N_14461,N_12592);
or U17452 (N_17452,N_10353,N_10378);
nand U17453 (N_17453,N_14953,N_11075);
nor U17454 (N_17454,N_10210,N_13081);
and U17455 (N_17455,N_14849,N_12332);
nand U17456 (N_17456,N_14664,N_11543);
nor U17457 (N_17457,N_11863,N_11623);
xnor U17458 (N_17458,N_12316,N_10564);
and U17459 (N_17459,N_13620,N_13754);
and U17460 (N_17460,N_10543,N_11022);
nand U17461 (N_17461,N_12526,N_10463);
or U17462 (N_17462,N_14593,N_12303);
nor U17463 (N_17463,N_13940,N_14559);
nor U17464 (N_17464,N_14868,N_14940);
nor U17465 (N_17465,N_12817,N_13987);
or U17466 (N_17466,N_13190,N_13338);
nor U17467 (N_17467,N_14255,N_13772);
xnor U17468 (N_17468,N_12321,N_11317);
and U17469 (N_17469,N_14748,N_10924);
nand U17470 (N_17470,N_12226,N_13951);
or U17471 (N_17471,N_12815,N_12974);
or U17472 (N_17472,N_10917,N_14237);
nor U17473 (N_17473,N_11807,N_12145);
nand U17474 (N_17474,N_12550,N_11300);
and U17475 (N_17475,N_12564,N_12151);
or U17476 (N_17476,N_12655,N_10971);
and U17477 (N_17477,N_10574,N_14129);
or U17478 (N_17478,N_12434,N_10006);
xor U17479 (N_17479,N_12441,N_11982);
and U17480 (N_17480,N_12477,N_14450);
nand U17481 (N_17481,N_14205,N_10734);
and U17482 (N_17482,N_13476,N_12479);
xor U17483 (N_17483,N_11409,N_14134);
nor U17484 (N_17484,N_14613,N_11670);
nand U17485 (N_17485,N_14693,N_12832);
or U17486 (N_17486,N_11416,N_12218);
nand U17487 (N_17487,N_14502,N_14185);
xor U17488 (N_17488,N_13253,N_14333);
nor U17489 (N_17489,N_14217,N_10651);
xor U17490 (N_17490,N_14107,N_10628);
and U17491 (N_17491,N_12675,N_10144);
nor U17492 (N_17492,N_14535,N_10624);
nand U17493 (N_17493,N_13678,N_11286);
and U17494 (N_17494,N_11805,N_10691);
xnor U17495 (N_17495,N_13341,N_11977);
xor U17496 (N_17496,N_10699,N_12461);
nor U17497 (N_17497,N_10417,N_11504);
nand U17498 (N_17498,N_12453,N_10875);
and U17499 (N_17499,N_11723,N_12190);
or U17500 (N_17500,N_13207,N_13540);
nor U17501 (N_17501,N_11161,N_14269);
or U17502 (N_17502,N_14901,N_13431);
or U17503 (N_17503,N_10137,N_13179);
or U17504 (N_17504,N_12307,N_11804);
or U17505 (N_17505,N_13838,N_14371);
nand U17506 (N_17506,N_13471,N_14983);
nand U17507 (N_17507,N_12954,N_12203);
and U17508 (N_17508,N_13531,N_10226);
xor U17509 (N_17509,N_10427,N_12758);
nor U17510 (N_17510,N_10734,N_11673);
nand U17511 (N_17511,N_12180,N_12112);
and U17512 (N_17512,N_14882,N_12261);
and U17513 (N_17513,N_10313,N_10889);
and U17514 (N_17514,N_13913,N_14445);
xor U17515 (N_17515,N_13537,N_12688);
nand U17516 (N_17516,N_14522,N_12202);
or U17517 (N_17517,N_14485,N_11247);
xor U17518 (N_17518,N_10726,N_14089);
and U17519 (N_17519,N_10201,N_10567);
nor U17520 (N_17520,N_12267,N_10489);
xor U17521 (N_17521,N_14116,N_13212);
nand U17522 (N_17522,N_14762,N_13662);
nand U17523 (N_17523,N_10962,N_13018);
or U17524 (N_17524,N_12884,N_11016);
xor U17525 (N_17525,N_13637,N_14665);
xor U17526 (N_17526,N_12934,N_10938);
nand U17527 (N_17527,N_13289,N_14550);
xor U17528 (N_17528,N_14688,N_12750);
nand U17529 (N_17529,N_12007,N_10790);
xor U17530 (N_17530,N_10194,N_12913);
or U17531 (N_17531,N_11251,N_11921);
xor U17532 (N_17532,N_10951,N_13569);
or U17533 (N_17533,N_13100,N_10282);
nor U17534 (N_17534,N_11915,N_13301);
or U17535 (N_17535,N_12377,N_10784);
nand U17536 (N_17536,N_11821,N_14503);
and U17537 (N_17537,N_11235,N_12279);
or U17538 (N_17538,N_12731,N_10334);
and U17539 (N_17539,N_12205,N_12742);
nand U17540 (N_17540,N_10987,N_14274);
xor U17541 (N_17541,N_13060,N_14617);
nor U17542 (N_17542,N_11107,N_12823);
and U17543 (N_17543,N_10552,N_14113);
nor U17544 (N_17544,N_13044,N_14806);
or U17545 (N_17545,N_14752,N_11117);
xor U17546 (N_17546,N_13991,N_14081);
and U17547 (N_17547,N_11898,N_14210);
xnor U17548 (N_17548,N_13519,N_13948);
or U17549 (N_17549,N_14853,N_10274);
nand U17550 (N_17550,N_12821,N_12591);
or U17551 (N_17551,N_14785,N_10762);
or U17552 (N_17552,N_12470,N_14353);
nand U17553 (N_17553,N_13067,N_14230);
nand U17554 (N_17554,N_14956,N_11502);
xor U17555 (N_17555,N_14337,N_12917);
nor U17556 (N_17556,N_12494,N_11160);
nor U17557 (N_17557,N_10356,N_13709);
nand U17558 (N_17558,N_12157,N_11015);
nor U17559 (N_17559,N_13999,N_13898);
or U17560 (N_17560,N_11156,N_13436);
or U17561 (N_17561,N_11134,N_10352);
nand U17562 (N_17562,N_12925,N_13156);
or U17563 (N_17563,N_12936,N_14409);
nand U17564 (N_17564,N_10520,N_10673);
xor U17565 (N_17565,N_10878,N_11839);
nor U17566 (N_17566,N_13552,N_11555);
xnor U17567 (N_17567,N_11501,N_10238);
or U17568 (N_17568,N_14681,N_10552);
and U17569 (N_17569,N_13179,N_11134);
and U17570 (N_17570,N_13388,N_12902);
nand U17571 (N_17571,N_13204,N_10939);
nor U17572 (N_17572,N_12994,N_13474);
nor U17573 (N_17573,N_11308,N_12012);
nor U17574 (N_17574,N_10207,N_11685);
and U17575 (N_17575,N_14988,N_14689);
and U17576 (N_17576,N_13712,N_11948);
xnor U17577 (N_17577,N_10294,N_12244);
nand U17578 (N_17578,N_11384,N_12325);
nor U17579 (N_17579,N_14606,N_12039);
and U17580 (N_17580,N_14834,N_14780);
and U17581 (N_17581,N_11391,N_12430);
and U17582 (N_17582,N_12976,N_11048);
nor U17583 (N_17583,N_13286,N_14656);
nand U17584 (N_17584,N_14678,N_11527);
xor U17585 (N_17585,N_11459,N_14874);
nor U17586 (N_17586,N_14441,N_10554);
nand U17587 (N_17587,N_14613,N_11733);
nand U17588 (N_17588,N_12349,N_14842);
or U17589 (N_17589,N_13142,N_10543);
and U17590 (N_17590,N_11612,N_12391);
xnor U17591 (N_17591,N_14494,N_14879);
xnor U17592 (N_17592,N_14280,N_12591);
nor U17593 (N_17593,N_14544,N_14235);
xor U17594 (N_17594,N_13507,N_10490);
and U17595 (N_17595,N_14578,N_12170);
nor U17596 (N_17596,N_13310,N_11335);
xnor U17597 (N_17597,N_14490,N_11878);
or U17598 (N_17598,N_14445,N_14251);
nor U17599 (N_17599,N_12603,N_13774);
and U17600 (N_17600,N_14639,N_10086);
nand U17601 (N_17601,N_12234,N_11270);
nor U17602 (N_17602,N_14857,N_10715);
nor U17603 (N_17603,N_11300,N_13051);
and U17604 (N_17604,N_13358,N_14730);
and U17605 (N_17605,N_10505,N_14993);
nand U17606 (N_17606,N_11852,N_13277);
nand U17607 (N_17607,N_13257,N_14112);
nor U17608 (N_17608,N_11167,N_10586);
xor U17609 (N_17609,N_13834,N_11931);
and U17610 (N_17610,N_14632,N_13471);
or U17611 (N_17611,N_13186,N_14119);
nand U17612 (N_17612,N_14743,N_14339);
nand U17613 (N_17613,N_11622,N_14500);
xor U17614 (N_17614,N_12074,N_12159);
nor U17615 (N_17615,N_13157,N_11815);
xnor U17616 (N_17616,N_11732,N_10874);
xnor U17617 (N_17617,N_12430,N_13135);
nand U17618 (N_17618,N_13260,N_13395);
nand U17619 (N_17619,N_10691,N_10005);
nand U17620 (N_17620,N_11043,N_10387);
nand U17621 (N_17621,N_10460,N_14784);
nand U17622 (N_17622,N_14290,N_10480);
xor U17623 (N_17623,N_10622,N_10127);
xor U17624 (N_17624,N_11991,N_14882);
or U17625 (N_17625,N_10579,N_13899);
or U17626 (N_17626,N_11209,N_14892);
nand U17627 (N_17627,N_14026,N_13003);
and U17628 (N_17628,N_14911,N_14655);
or U17629 (N_17629,N_14548,N_10210);
or U17630 (N_17630,N_12454,N_11868);
and U17631 (N_17631,N_11487,N_12791);
or U17632 (N_17632,N_10053,N_14120);
nand U17633 (N_17633,N_11887,N_11961);
and U17634 (N_17634,N_13256,N_13321);
or U17635 (N_17635,N_10537,N_11858);
nor U17636 (N_17636,N_10839,N_14643);
nand U17637 (N_17637,N_11993,N_14138);
and U17638 (N_17638,N_13858,N_13073);
xnor U17639 (N_17639,N_13644,N_13180);
nor U17640 (N_17640,N_14743,N_14522);
and U17641 (N_17641,N_14904,N_11866);
nor U17642 (N_17642,N_12785,N_13064);
nor U17643 (N_17643,N_14312,N_10438);
or U17644 (N_17644,N_10420,N_14254);
xnor U17645 (N_17645,N_10387,N_14195);
nor U17646 (N_17646,N_13914,N_14915);
and U17647 (N_17647,N_12405,N_13106);
nor U17648 (N_17648,N_14007,N_13145);
nand U17649 (N_17649,N_10299,N_14402);
xnor U17650 (N_17650,N_11299,N_13512);
nand U17651 (N_17651,N_12338,N_11567);
or U17652 (N_17652,N_14618,N_12103);
and U17653 (N_17653,N_14685,N_12081);
nand U17654 (N_17654,N_11739,N_10258);
and U17655 (N_17655,N_11416,N_14960);
xor U17656 (N_17656,N_12903,N_13898);
or U17657 (N_17657,N_14281,N_12276);
and U17658 (N_17658,N_13671,N_14450);
xor U17659 (N_17659,N_11916,N_11938);
nand U17660 (N_17660,N_11752,N_14249);
nand U17661 (N_17661,N_10968,N_12278);
nor U17662 (N_17662,N_10360,N_11896);
nor U17663 (N_17663,N_12623,N_11274);
xor U17664 (N_17664,N_14255,N_14776);
xor U17665 (N_17665,N_11164,N_10138);
or U17666 (N_17666,N_14047,N_11179);
xor U17667 (N_17667,N_14485,N_12297);
xor U17668 (N_17668,N_13459,N_12166);
nand U17669 (N_17669,N_11725,N_13064);
and U17670 (N_17670,N_13335,N_10046);
and U17671 (N_17671,N_14089,N_11858);
nor U17672 (N_17672,N_14932,N_13100);
and U17673 (N_17673,N_10594,N_13383);
xor U17674 (N_17674,N_11017,N_13435);
and U17675 (N_17675,N_14632,N_13610);
nor U17676 (N_17676,N_12691,N_10720);
nor U17677 (N_17677,N_12845,N_14662);
and U17678 (N_17678,N_12140,N_12906);
nand U17679 (N_17679,N_14881,N_12514);
or U17680 (N_17680,N_12037,N_10329);
xnor U17681 (N_17681,N_12060,N_11956);
nand U17682 (N_17682,N_12767,N_10379);
xnor U17683 (N_17683,N_14086,N_13200);
nand U17684 (N_17684,N_14159,N_13911);
nand U17685 (N_17685,N_11230,N_14357);
nor U17686 (N_17686,N_12739,N_12129);
nor U17687 (N_17687,N_10642,N_13407);
and U17688 (N_17688,N_10237,N_11709);
and U17689 (N_17689,N_10790,N_14953);
and U17690 (N_17690,N_11419,N_13747);
xnor U17691 (N_17691,N_10082,N_13992);
or U17692 (N_17692,N_13092,N_12668);
or U17693 (N_17693,N_13000,N_10917);
nand U17694 (N_17694,N_10572,N_13283);
xnor U17695 (N_17695,N_13422,N_10328);
and U17696 (N_17696,N_13510,N_12309);
nand U17697 (N_17697,N_12733,N_13030);
or U17698 (N_17698,N_14209,N_11562);
nand U17699 (N_17699,N_14841,N_12751);
nand U17700 (N_17700,N_12248,N_14781);
and U17701 (N_17701,N_12848,N_12000);
nand U17702 (N_17702,N_11235,N_14565);
nor U17703 (N_17703,N_13731,N_12502);
nand U17704 (N_17704,N_10860,N_13166);
or U17705 (N_17705,N_12917,N_14024);
nand U17706 (N_17706,N_10390,N_10702);
and U17707 (N_17707,N_11345,N_10817);
and U17708 (N_17708,N_13583,N_10561);
xor U17709 (N_17709,N_12796,N_13720);
xnor U17710 (N_17710,N_13948,N_14168);
xor U17711 (N_17711,N_13684,N_12344);
nor U17712 (N_17712,N_11906,N_11172);
xnor U17713 (N_17713,N_13460,N_13729);
nor U17714 (N_17714,N_12450,N_13542);
nor U17715 (N_17715,N_11506,N_12857);
nor U17716 (N_17716,N_14991,N_12548);
or U17717 (N_17717,N_14848,N_13907);
nor U17718 (N_17718,N_10776,N_11807);
nor U17719 (N_17719,N_12999,N_12761);
xnor U17720 (N_17720,N_13389,N_13012);
nand U17721 (N_17721,N_11843,N_13765);
or U17722 (N_17722,N_14164,N_12408);
nand U17723 (N_17723,N_11015,N_13145);
and U17724 (N_17724,N_14103,N_14657);
nand U17725 (N_17725,N_12881,N_13717);
and U17726 (N_17726,N_13005,N_14361);
and U17727 (N_17727,N_13995,N_14712);
xnor U17728 (N_17728,N_14714,N_10393);
and U17729 (N_17729,N_14349,N_14638);
nand U17730 (N_17730,N_13358,N_14355);
nand U17731 (N_17731,N_12585,N_12888);
nor U17732 (N_17732,N_11291,N_11562);
nor U17733 (N_17733,N_13058,N_12814);
nand U17734 (N_17734,N_12282,N_13761);
nand U17735 (N_17735,N_13950,N_10558);
nor U17736 (N_17736,N_14291,N_12748);
nor U17737 (N_17737,N_10012,N_12934);
nand U17738 (N_17738,N_12383,N_12423);
or U17739 (N_17739,N_14188,N_12516);
or U17740 (N_17740,N_14305,N_12088);
nor U17741 (N_17741,N_11003,N_11265);
xor U17742 (N_17742,N_13148,N_12584);
xor U17743 (N_17743,N_13673,N_14437);
nand U17744 (N_17744,N_11022,N_10755);
and U17745 (N_17745,N_14178,N_12252);
xnor U17746 (N_17746,N_14906,N_10148);
nand U17747 (N_17747,N_14216,N_10496);
or U17748 (N_17748,N_10291,N_12604);
and U17749 (N_17749,N_10751,N_10877);
nor U17750 (N_17750,N_13772,N_12211);
and U17751 (N_17751,N_11515,N_14790);
nor U17752 (N_17752,N_13747,N_13138);
nand U17753 (N_17753,N_11610,N_13906);
and U17754 (N_17754,N_10622,N_12428);
xnor U17755 (N_17755,N_10515,N_11603);
or U17756 (N_17756,N_12879,N_13096);
or U17757 (N_17757,N_10864,N_13508);
nand U17758 (N_17758,N_14196,N_14108);
xnor U17759 (N_17759,N_12821,N_10367);
xnor U17760 (N_17760,N_13836,N_11348);
and U17761 (N_17761,N_11245,N_14875);
nor U17762 (N_17762,N_12070,N_10182);
xor U17763 (N_17763,N_11160,N_10034);
xnor U17764 (N_17764,N_12040,N_10357);
nand U17765 (N_17765,N_14365,N_12345);
xnor U17766 (N_17766,N_11399,N_14785);
and U17767 (N_17767,N_10618,N_14253);
and U17768 (N_17768,N_11609,N_14207);
nand U17769 (N_17769,N_12169,N_12136);
nand U17770 (N_17770,N_13944,N_10032);
and U17771 (N_17771,N_12810,N_10974);
xnor U17772 (N_17772,N_12864,N_10296);
xor U17773 (N_17773,N_10346,N_13938);
xnor U17774 (N_17774,N_10154,N_11018);
nand U17775 (N_17775,N_13492,N_14826);
nand U17776 (N_17776,N_14134,N_13515);
nor U17777 (N_17777,N_14852,N_14091);
or U17778 (N_17778,N_10326,N_11163);
xnor U17779 (N_17779,N_10273,N_12051);
nand U17780 (N_17780,N_10697,N_14027);
xnor U17781 (N_17781,N_13286,N_12065);
nand U17782 (N_17782,N_13603,N_11371);
and U17783 (N_17783,N_11637,N_10493);
nand U17784 (N_17784,N_13514,N_11703);
nand U17785 (N_17785,N_10733,N_13813);
xor U17786 (N_17786,N_14680,N_14589);
or U17787 (N_17787,N_14334,N_10110);
and U17788 (N_17788,N_11464,N_12305);
and U17789 (N_17789,N_12873,N_10106);
xor U17790 (N_17790,N_11860,N_10038);
nand U17791 (N_17791,N_14488,N_10357);
and U17792 (N_17792,N_12984,N_12631);
nand U17793 (N_17793,N_14867,N_13505);
or U17794 (N_17794,N_11074,N_12713);
xor U17795 (N_17795,N_14318,N_11257);
and U17796 (N_17796,N_10154,N_13487);
or U17797 (N_17797,N_11243,N_13086);
or U17798 (N_17798,N_14535,N_10201);
and U17799 (N_17799,N_13045,N_11790);
xor U17800 (N_17800,N_11692,N_12646);
xnor U17801 (N_17801,N_13261,N_14347);
nor U17802 (N_17802,N_13863,N_12594);
and U17803 (N_17803,N_14190,N_12563);
nor U17804 (N_17804,N_12226,N_12048);
nor U17805 (N_17805,N_11631,N_14601);
xnor U17806 (N_17806,N_14989,N_14227);
and U17807 (N_17807,N_11082,N_10024);
or U17808 (N_17808,N_11467,N_12250);
or U17809 (N_17809,N_14908,N_12265);
and U17810 (N_17810,N_12145,N_11131);
or U17811 (N_17811,N_13285,N_13808);
xor U17812 (N_17812,N_10193,N_13347);
or U17813 (N_17813,N_13665,N_12724);
nor U17814 (N_17814,N_13780,N_14741);
or U17815 (N_17815,N_14239,N_13356);
and U17816 (N_17816,N_14721,N_13421);
xnor U17817 (N_17817,N_11565,N_12242);
or U17818 (N_17818,N_14035,N_13022);
nand U17819 (N_17819,N_12327,N_14374);
and U17820 (N_17820,N_13129,N_11261);
nor U17821 (N_17821,N_14729,N_12949);
nand U17822 (N_17822,N_13757,N_12949);
nand U17823 (N_17823,N_14040,N_10396);
nor U17824 (N_17824,N_13701,N_12020);
nand U17825 (N_17825,N_10342,N_14759);
and U17826 (N_17826,N_12617,N_11509);
nand U17827 (N_17827,N_13382,N_10686);
xnor U17828 (N_17828,N_11979,N_10101);
nand U17829 (N_17829,N_10416,N_13931);
or U17830 (N_17830,N_14615,N_11982);
nand U17831 (N_17831,N_11211,N_14098);
or U17832 (N_17832,N_13929,N_14734);
or U17833 (N_17833,N_12449,N_14066);
xnor U17834 (N_17834,N_14304,N_10792);
and U17835 (N_17835,N_10451,N_14908);
or U17836 (N_17836,N_10366,N_11462);
and U17837 (N_17837,N_10601,N_14105);
nand U17838 (N_17838,N_12969,N_12960);
nand U17839 (N_17839,N_12674,N_13777);
nand U17840 (N_17840,N_10982,N_10140);
and U17841 (N_17841,N_14498,N_12281);
nand U17842 (N_17842,N_13874,N_11734);
and U17843 (N_17843,N_14812,N_14926);
and U17844 (N_17844,N_12785,N_14487);
and U17845 (N_17845,N_13669,N_13357);
or U17846 (N_17846,N_14181,N_14304);
xnor U17847 (N_17847,N_12159,N_14788);
and U17848 (N_17848,N_12714,N_12646);
and U17849 (N_17849,N_14398,N_12665);
xnor U17850 (N_17850,N_13228,N_12815);
or U17851 (N_17851,N_10250,N_12900);
xnor U17852 (N_17852,N_10030,N_11983);
or U17853 (N_17853,N_14109,N_11833);
or U17854 (N_17854,N_13634,N_11259);
and U17855 (N_17855,N_13861,N_12063);
or U17856 (N_17856,N_10558,N_10578);
nand U17857 (N_17857,N_10272,N_11036);
or U17858 (N_17858,N_12624,N_11765);
or U17859 (N_17859,N_14130,N_10060);
and U17860 (N_17860,N_13276,N_14769);
xor U17861 (N_17861,N_11409,N_14759);
nor U17862 (N_17862,N_13419,N_14096);
and U17863 (N_17863,N_13113,N_10081);
or U17864 (N_17864,N_14345,N_12685);
nor U17865 (N_17865,N_11913,N_13815);
and U17866 (N_17866,N_10215,N_11348);
and U17867 (N_17867,N_12905,N_11413);
or U17868 (N_17868,N_13028,N_13306);
nand U17869 (N_17869,N_12377,N_13514);
xor U17870 (N_17870,N_11825,N_10999);
or U17871 (N_17871,N_13631,N_12885);
nand U17872 (N_17872,N_13111,N_13048);
xor U17873 (N_17873,N_12929,N_10603);
nor U17874 (N_17874,N_14962,N_12708);
nor U17875 (N_17875,N_12177,N_14722);
nand U17876 (N_17876,N_10192,N_14086);
or U17877 (N_17877,N_10858,N_14570);
and U17878 (N_17878,N_11348,N_12100);
or U17879 (N_17879,N_12925,N_12701);
xor U17880 (N_17880,N_10890,N_11314);
xnor U17881 (N_17881,N_10580,N_11564);
nor U17882 (N_17882,N_13040,N_14736);
xor U17883 (N_17883,N_11558,N_12899);
and U17884 (N_17884,N_14946,N_10459);
or U17885 (N_17885,N_10316,N_12383);
nor U17886 (N_17886,N_13431,N_12383);
or U17887 (N_17887,N_11337,N_11818);
or U17888 (N_17888,N_14217,N_10179);
and U17889 (N_17889,N_10576,N_12416);
nand U17890 (N_17890,N_13127,N_10421);
nand U17891 (N_17891,N_14630,N_12239);
or U17892 (N_17892,N_11497,N_14332);
xor U17893 (N_17893,N_13889,N_12755);
nor U17894 (N_17894,N_14189,N_10727);
or U17895 (N_17895,N_11303,N_12095);
xnor U17896 (N_17896,N_14766,N_10775);
xnor U17897 (N_17897,N_11861,N_10757);
xor U17898 (N_17898,N_13871,N_13127);
and U17899 (N_17899,N_13318,N_13221);
or U17900 (N_17900,N_12828,N_10154);
and U17901 (N_17901,N_10419,N_13405);
and U17902 (N_17902,N_14618,N_10239);
nor U17903 (N_17903,N_12168,N_10321);
nand U17904 (N_17904,N_10467,N_12701);
or U17905 (N_17905,N_13256,N_10481);
and U17906 (N_17906,N_14674,N_12524);
nand U17907 (N_17907,N_13316,N_13514);
or U17908 (N_17908,N_14263,N_14556);
or U17909 (N_17909,N_12309,N_11601);
or U17910 (N_17910,N_14865,N_13011);
nand U17911 (N_17911,N_11712,N_14574);
nand U17912 (N_17912,N_10601,N_13403);
nor U17913 (N_17913,N_12070,N_10160);
nand U17914 (N_17914,N_10418,N_12598);
and U17915 (N_17915,N_13819,N_13964);
nand U17916 (N_17916,N_14931,N_12632);
nand U17917 (N_17917,N_14005,N_11431);
xnor U17918 (N_17918,N_11060,N_14226);
and U17919 (N_17919,N_10588,N_14213);
xor U17920 (N_17920,N_13148,N_11275);
nand U17921 (N_17921,N_11247,N_10677);
nand U17922 (N_17922,N_11736,N_11431);
and U17923 (N_17923,N_12952,N_10929);
nor U17924 (N_17924,N_14479,N_10295);
nand U17925 (N_17925,N_11852,N_13105);
and U17926 (N_17926,N_13056,N_10746);
xnor U17927 (N_17927,N_10900,N_11939);
xor U17928 (N_17928,N_14531,N_14241);
and U17929 (N_17929,N_10306,N_12349);
or U17930 (N_17930,N_12008,N_14786);
or U17931 (N_17931,N_12765,N_11912);
xnor U17932 (N_17932,N_11276,N_11497);
xor U17933 (N_17933,N_14302,N_10907);
and U17934 (N_17934,N_12949,N_10430);
or U17935 (N_17935,N_10537,N_13592);
nand U17936 (N_17936,N_14099,N_10459);
nand U17937 (N_17937,N_12922,N_14916);
and U17938 (N_17938,N_14381,N_12776);
xor U17939 (N_17939,N_14653,N_12595);
nor U17940 (N_17940,N_12459,N_14926);
nand U17941 (N_17941,N_10374,N_12341);
nor U17942 (N_17942,N_14284,N_13050);
xnor U17943 (N_17943,N_13586,N_14025);
nor U17944 (N_17944,N_14429,N_12767);
nand U17945 (N_17945,N_11790,N_14668);
and U17946 (N_17946,N_11333,N_14315);
nor U17947 (N_17947,N_10862,N_13839);
xnor U17948 (N_17948,N_10831,N_14999);
nand U17949 (N_17949,N_14753,N_10739);
xnor U17950 (N_17950,N_11110,N_12962);
and U17951 (N_17951,N_11146,N_13884);
xnor U17952 (N_17952,N_10357,N_12376);
and U17953 (N_17953,N_12723,N_10148);
nor U17954 (N_17954,N_12783,N_13019);
nor U17955 (N_17955,N_12055,N_14077);
xnor U17956 (N_17956,N_11151,N_10495);
nor U17957 (N_17957,N_11259,N_10875);
xor U17958 (N_17958,N_14718,N_11579);
nor U17959 (N_17959,N_12078,N_13995);
nand U17960 (N_17960,N_14934,N_11914);
and U17961 (N_17961,N_13024,N_13095);
nand U17962 (N_17962,N_13055,N_10644);
or U17963 (N_17963,N_10070,N_10273);
or U17964 (N_17964,N_13018,N_11038);
and U17965 (N_17965,N_10163,N_13892);
xor U17966 (N_17966,N_10919,N_13927);
xor U17967 (N_17967,N_10325,N_14603);
or U17968 (N_17968,N_14005,N_11921);
or U17969 (N_17969,N_11867,N_13364);
or U17970 (N_17970,N_10119,N_14052);
or U17971 (N_17971,N_12039,N_12483);
and U17972 (N_17972,N_14632,N_14780);
nor U17973 (N_17973,N_10384,N_10230);
nand U17974 (N_17974,N_12923,N_13425);
nand U17975 (N_17975,N_12446,N_12909);
and U17976 (N_17976,N_14643,N_11298);
xor U17977 (N_17977,N_13964,N_12567);
nor U17978 (N_17978,N_13460,N_10701);
or U17979 (N_17979,N_10932,N_13214);
nor U17980 (N_17980,N_12936,N_11813);
and U17981 (N_17981,N_14498,N_12086);
xor U17982 (N_17982,N_12481,N_12772);
or U17983 (N_17983,N_13814,N_13607);
nand U17984 (N_17984,N_10036,N_13093);
or U17985 (N_17985,N_13905,N_12154);
and U17986 (N_17986,N_10608,N_11683);
and U17987 (N_17987,N_10239,N_10283);
xor U17988 (N_17988,N_13767,N_13501);
xor U17989 (N_17989,N_10224,N_10136);
nor U17990 (N_17990,N_11376,N_10702);
nand U17991 (N_17991,N_14669,N_13588);
nand U17992 (N_17992,N_12391,N_12147);
xor U17993 (N_17993,N_11597,N_14744);
nor U17994 (N_17994,N_10228,N_10277);
nand U17995 (N_17995,N_12341,N_11157);
nor U17996 (N_17996,N_13138,N_10734);
or U17997 (N_17997,N_10655,N_10073);
nand U17998 (N_17998,N_12429,N_13003);
nor U17999 (N_17999,N_10617,N_11167);
or U18000 (N_18000,N_14298,N_12216);
or U18001 (N_18001,N_12805,N_11660);
nand U18002 (N_18002,N_13931,N_11903);
and U18003 (N_18003,N_11597,N_14090);
xnor U18004 (N_18004,N_13447,N_12959);
and U18005 (N_18005,N_11850,N_12279);
and U18006 (N_18006,N_12247,N_11412);
or U18007 (N_18007,N_10589,N_14493);
nor U18008 (N_18008,N_12408,N_10082);
nand U18009 (N_18009,N_11743,N_14528);
nor U18010 (N_18010,N_13618,N_11919);
and U18011 (N_18011,N_13328,N_10678);
nor U18012 (N_18012,N_12424,N_13491);
nor U18013 (N_18013,N_13044,N_14189);
nand U18014 (N_18014,N_10809,N_12077);
nor U18015 (N_18015,N_13086,N_10063);
nand U18016 (N_18016,N_10936,N_12053);
or U18017 (N_18017,N_13932,N_14871);
and U18018 (N_18018,N_11809,N_14330);
xor U18019 (N_18019,N_14830,N_14190);
xnor U18020 (N_18020,N_13900,N_14499);
xnor U18021 (N_18021,N_14757,N_10172);
xnor U18022 (N_18022,N_14376,N_10223);
or U18023 (N_18023,N_12724,N_11469);
and U18024 (N_18024,N_14104,N_12888);
nand U18025 (N_18025,N_11855,N_13301);
and U18026 (N_18026,N_14981,N_12672);
xor U18027 (N_18027,N_13702,N_10820);
or U18028 (N_18028,N_12640,N_13819);
nand U18029 (N_18029,N_14657,N_13784);
xor U18030 (N_18030,N_10989,N_14675);
or U18031 (N_18031,N_14191,N_13700);
or U18032 (N_18032,N_12160,N_11851);
nand U18033 (N_18033,N_12859,N_13528);
and U18034 (N_18034,N_12538,N_14502);
nand U18035 (N_18035,N_10312,N_10252);
or U18036 (N_18036,N_11401,N_14263);
nor U18037 (N_18037,N_14574,N_10878);
nand U18038 (N_18038,N_11468,N_10156);
nand U18039 (N_18039,N_11089,N_10827);
or U18040 (N_18040,N_10753,N_10820);
and U18041 (N_18041,N_10219,N_11959);
nor U18042 (N_18042,N_13030,N_12224);
nand U18043 (N_18043,N_12282,N_13970);
xnor U18044 (N_18044,N_10414,N_12260);
or U18045 (N_18045,N_14918,N_11450);
or U18046 (N_18046,N_10286,N_11301);
xnor U18047 (N_18047,N_11009,N_14550);
and U18048 (N_18048,N_12556,N_10883);
and U18049 (N_18049,N_10512,N_11922);
nand U18050 (N_18050,N_13331,N_13000);
or U18051 (N_18051,N_11564,N_10647);
and U18052 (N_18052,N_12090,N_10960);
nand U18053 (N_18053,N_12356,N_12835);
or U18054 (N_18054,N_12606,N_10878);
nand U18055 (N_18055,N_13516,N_12653);
nor U18056 (N_18056,N_10870,N_12313);
or U18057 (N_18057,N_12231,N_11796);
or U18058 (N_18058,N_12014,N_10719);
nor U18059 (N_18059,N_12178,N_13253);
xnor U18060 (N_18060,N_11494,N_13836);
xor U18061 (N_18061,N_11515,N_14038);
nor U18062 (N_18062,N_12105,N_10609);
nand U18063 (N_18063,N_12250,N_12962);
nand U18064 (N_18064,N_14759,N_13092);
xnor U18065 (N_18065,N_11538,N_11702);
nor U18066 (N_18066,N_12596,N_13207);
nand U18067 (N_18067,N_10500,N_12951);
or U18068 (N_18068,N_11093,N_11985);
nor U18069 (N_18069,N_11370,N_14749);
xnor U18070 (N_18070,N_12954,N_10584);
or U18071 (N_18071,N_10943,N_12111);
or U18072 (N_18072,N_13012,N_13923);
xnor U18073 (N_18073,N_14989,N_12154);
nand U18074 (N_18074,N_13437,N_13593);
nand U18075 (N_18075,N_14114,N_14325);
xnor U18076 (N_18076,N_13493,N_10089);
xor U18077 (N_18077,N_10776,N_13652);
or U18078 (N_18078,N_11704,N_12400);
nor U18079 (N_18079,N_13056,N_14971);
or U18080 (N_18080,N_12098,N_12595);
nor U18081 (N_18081,N_12007,N_10804);
and U18082 (N_18082,N_13968,N_10251);
xnor U18083 (N_18083,N_13160,N_12921);
nor U18084 (N_18084,N_10361,N_13866);
nand U18085 (N_18085,N_10683,N_11116);
xor U18086 (N_18086,N_12650,N_11575);
nor U18087 (N_18087,N_14827,N_14756);
or U18088 (N_18088,N_13379,N_12301);
nor U18089 (N_18089,N_13777,N_10618);
nor U18090 (N_18090,N_11924,N_14499);
or U18091 (N_18091,N_11585,N_12382);
nand U18092 (N_18092,N_13628,N_13539);
or U18093 (N_18093,N_13790,N_12405);
xnor U18094 (N_18094,N_11880,N_11537);
and U18095 (N_18095,N_10308,N_10673);
or U18096 (N_18096,N_10399,N_13939);
nor U18097 (N_18097,N_14678,N_14329);
nor U18098 (N_18098,N_12648,N_13076);
or U18099 (N_18099,N_14401,N_13106);
xnor U18100 (N_18100,N_14238,N_13329);
and U18101 (N_18101,N_12553,N_11448);
or U18102 (N_18102,N_12519,N_12820);
nor U18103 (N_18103,N_12199,N_10374);
and U18104 (N_18104,N_13567,N_12408);
and U18105 (N_18105,N_13580,N_10132);
and U18106 (N_18106,N_12441,N_13094);
nor U18107 (N_18107,N_11512,N_13648);
nor U18108 (N_18108,N_12459,N_13567);
and U18109 (N_18109,N_12631,N_13656);
and U18110 (N_18110,N_10155,N_10640);
nor U18111 (N_18111,N_12017,N_14623);
nor U18112 (N_18112,N_13570,N_14840);
nor U18113 (N_18113,N_13101,N_13891);
xor U18114 (N_18114,N_11681,N_13823);
and U18115 (N_18115,N_14642,N_13167);
or U18116 (N_18116,N_12787,N_14297);
nand U18117 (N_18117,N_12785,N_14213);
nor U18118 (N_18118,N_13974,N_12994);
nand U18119 (N_18119,N_13569,N_12585);
nor U18120 (N_18120,N_12579,N_13072);
and U18121 (N_18121,N_10823,N_13803);
or U18122 (N_18122,N_11984,N_14113);
and U18123 (N_18123,N_11353,N_12062);
and U18124 (N_18124,N_13152,N_11138);
and U18125 (N_18125,N_14119,N_11253);
nand U18126 (N_18126,N_10993,N_14166);
or U18127 (N_18127,N_14269,N_11446);
xnor U18128 (N_18128,N_11076,N_12831);
and U18129 (N_18129,N_14488,N_14613);
or U18130 (N_18130,N_13101,N_10695);
nor U18131 (N_18131,N_12526,N_13304);
xnor U18132 (N_18132,N_14763,N_11465);
xnor U18133 (N_18133,N_11864,N_13202);
nor U18134 (N_18134,N_12513,N_10526);
and U18135 (N_18135,N_12661,N_13847);
nand U18136 (N_18136,N_11033,N_11341);
or U18137 (N_18137,N_14739,N_11794);
and U18138 (N_18138,N_12712,N_12352);
nor U18139 (N_18139,N_11701,N_14520);
and U18140 (N_18140,N_12236,N_14653);
nor U18141 (N_18141,N_10604,N_11425);
nor U18142 (N_18142,N_12887,N_12467);
or U18143 (N_18143,N_10427,N_13723);
nand U18144 (N_18144,N_14081,N_14353);
and U18145 (N_18145,N_14617,N_10859);
and U18146 (N_18146,N_13487,N_14279);
xor U18147 (N_18147,N_14855,N_14002);
nand U18148 (N_18148,N_12556,N_12035);
or U18149 (N_18149,N_11655,N_13271);
or U18150 (N_18150,N_11022,N_10147);
nand U18151 (N_18151,N_14929,N_11324);
or U18152 (N_18152,N_10019,N_13986);
nand U18153 (N_18153,N_13021,N_13330);
xor U18154 (N_18154,N_13150,N_10415);
nand U18155 (N_18155,N_14660,N_12790);
xor U18156 (N_18156,N_11492,N_10589);
and U18157 (N_18157,N_13286,N_11527);
or U18158 (N_18158,N_11503,N_11220);
nand U18159 (N_18159,N_11861,N_14610);
xnor U18160 (N_18160,N_14345,N_10595);
nor U18161 (N_18161,N_12029,N_12872);
nand U18162 (N_18162,N_13962,N_11356);
or U18163 (N_18163,N_11841,N_14082);
nand U18164 (N_18164,N_10360,N_13757);
or U18165 (N_18165,N_10921,N_10528);
nor U18166 (N_18166,N_13723,N_14258);
nor U18167 (N_18167,N_12141,N_14869);
and U18168 (N_18168,N_10415,N_10236);
or U18169 (N_18169,N_10294,N_13479);
and U18170 (N_18170,N_11669,N_11619);
nand U18171 (N_18171,N_13685,N_12911);
xor U18172 (N_18172,N_12275,N_12473);
and U18173 (N_18173,N_12033,N_12389);
and U18174 (N_18174,N_10586,N_10829);
and U18175 (N_18175,N_10852,N_14346);
or U18176 (N_18176,N_14801,N_12057);
xor U18177 (N_18177,N_10238,N_11766);
and U18178 (N_18178,N_10587,N_13493);
nor U18179 (N_18179,N_14148,N_14223);
or U18180 (N_18180,N_11847,N_12091);
and U18181 (N_18181,N_12455,N_13566);
or U18182 (N_18182,N_10344,N_14486);
xnor U18183 (N_18183,N_11774,N_13734);
nor U18184 (N_18184,N_14900,N_14693);
or U18185 (N_18185,N_12419,N_11959);
nor U18186 (N_18186,N_14169,N_13578);
xnor U18187 (N_18187,N_11588,N_13239);
or U18188 (N_18188,N_11588,N_11142);
nand U18189 (N_18189,N_11523,N_13375);
or U18190 (N_18190,N_12928,N_10824);
nand U18191 (N_18191,N_12085,N_12838);
nand U18192 (N_18192,N_14793,N_12835);
xnor U18193 (N_18193,N_10015,N_11669);
nand U18194 (N_18194,N_13926,N_14170);
nand U18195 (N_18195,N_12436,N_11647);
nand U18196 (N_18196,N_13381,N_13694);
nor U18197 (N_18197,N_13111,N_10668);
nand U18198 (N_18198,N_13995,N_10531);
nand U18199 (N_18199,N_13369,N_12467);
nor U18200 (N_18200,N_11577,N_10824);
nand U18201 (N_18201,N_12570,N_12940);
xnor U18202 (N_18202,N_11962,N_11906);
and U18203 (N_18203,N_12265,N_13073);
nand U18204 (N_18204,N_11663,N_10784);
or U18205 (N_18205,N_13914,N_10236);
xnor U18206 (N_18206,N_14700,N_14292);
xnor U18207 (N_18207,N_11894,N_14221);
and U18208 (N_18208,N_14755,N_11185);
nand U18209 (N_18209,N_12206,N_10340);
and U18210 (N_18210,N_11385,N_12787);
xor U18211 (N_18211,N_14345,N_10250);
and U18212 (N_18212,N_14668,N_14610);
or U18213 (N_18213,N_13789,N_13326);
nor U18214 (N_18214,N_14478,N_10350);
nor U18215 (N_18215,N_11014,N_12222);
or U18216 (N_18216,N_11916,N_13976);
xor U18217 (N_18217,N_10253,N_13195);
xor U18218 (N_18218,N_13043,N_14802);
xor U18219 (N_18219,N_11213,N_11714);
xor U18220 (N_18220,N_10672,N_14695);
nand U18221 (N_18221,N_10489,N_13969);
or U18222 (N_18222,N_10178,N_14031);
and U18223 (N_18223,N_13219,N_11673);
and U18224 (N_18224,N_14085,N_11886);
and U18225 (N_18225,N_13467,N_13948);
nor U18226 (N_18226,N_12557,N_12996);
xnor U18227 (N_18227,N_12942,N_10061);
nor U18228 (N_18228,N_13769,N_11344);
nor U18229 (N_18229,N_14506,N_13742);
xnor U18230 (N_18230,N_11511,N_14557);
nand U18231 (N_18231,N_12597,N_10368);
or U18232 (N_18232,N_14076,N_14053);
or U18233 (N_18233,N_10670,N_13756);
nand U18234 (N_18234,N_12632,N_14553);
nand U18235 (N_18235,N_11022,N_10031);
nand U18236 (N_18236,N_12437,N_12116);
nor U18237 (N_18237,N_10401,N_13063);
nor U18238 (N_18238,N_10967,N_14381);
xor U18239 (N_18239,N_14599,N_12609);
nor U18240 (N_18240,N_13797,N_11102);
nand U18241 (N_18241,N_12095,N_12049);
nand U18242 (N_18242,N_13700,N_10848);
xor U18243 (N_18243,N_14083,N_13878);
xor U18244 (N_18244,N_14932,N_11717);
nor U18245 (N_18245,N_14435,N_13009);
and U18246 (N_18246,N_14267,N_12482);
and U18247 (N_18247,N_12263,N_14926);
and U18248 (N_18248,N_11643,N_13280);
nor U18249 (N_18249,N_13996,N_13382);
nand U18250 (N_18250,N_10677,N_12742);
nor U18251 (N_18251,N_13665,N_11624);
and U18252 (N_18252,N_10446,N_14476);
xnor U18253 (N_18253,N_13068,N_14879);
or U18254 (N_18254,N_10465,N_10978);
or U18255 (N_18255,N_11938,N_14744);
nor U18256 (N_18256,N_10922,N_10624);
nor U18257 (N_18257,N_14458,N_11615);
xnor U18258 (N_18258,N_14351,N_14051);
nand U18259 (N_18259,N_13742,N_11626);
nor U18260 (N_18260,N_13010,N_13742);
nor U18261 (N_18261,N_11011,N_14925);
nor U18262 (N_18262,N_12231,N_11885);
nand U18263 (N_18263,N_11801,N_14973);
nor U18264 (N_18264,N_14537,N_10282);
or U18265 (N_18265,N_13757,N_11134);
nor U18266 (N_18266,N_14882,N_10557);
or U18267 (N_18267,N_13088,N_11966);
nor U18268 (N_18268,N_11980,N_13215);
nand U18269 (N_18269,N_11953,N_10327);
and U18270 (N_18270,N_10305,N_11182);
or U18271 (N_18271,N_14664,N_13780);
or U18272 (N_18272,N_10052,N_14582);
and U18273 (N_18273,N_10715,N_11354);
or U18274 (N_18274,N_12019,N_11783);
or U18275 (N_18275,N_13011,N_10285);
or U18276 (N_18276,N_10568,N_10958);
and U18277 (N_18277,N_13597,N_11087);
or U18278 (N_18278,N_10773,N_10570);
and U18279 (N_18279,N_10302,N_13396);
nand U18280 (N_18280,N_12062,N_11780);
or U18281 (N_18281,N_11717,N_14565);
nor U18282 (N_18282,N_11503,N_12515);
and U18283 (N_18283,N_13957,N_12623);
or U18284 (N_18284,N_14787,N_11284);
nand U18285 (N_18285,N_11608,N_12726);
nand U18286 (N_18286,N_10998,N_13524);
xor U18287 (N_18287,N_10277,N_14992);
and U18288 (N_18288,N_10131,N_10631);
xnor U18289 (N_18289,N_12201,N_13846);
and U18290 (N_18290,N_14370,N_10097);
nand U18291 (N_18291,N_12948,N_11990);
or U18292 (N_18292,N_12491,N_12702);
or U18293 (N_18293,N_14448,N_10018);
or U18294 (N_18294,N_12016,N_10890);
xnor U18295 (N_18295,N_12162,N_11489);
xor U18296 (N_18296,N_10430,N_14441);
xor U18297 (N_18297,N_10062,N_12363);
nand U18298 (N_18298,N_11054,N_10994);
nor U18299 (N_18299,N_11171,N_13035);
nor U18300 (N_18300,N_12032,N_14223);
and U18301 (N_18301,N_11869,N_13033);
or U18302 (N_18302,N_14065,N_10309);
xor U18303 (N_18303,N_14711,N_10203);
nor U18304 (N_18304,N_12761,N_10094);
nand U18305 (N_18305,N_11077,N_11247);
and U18306 (N_18306,N_10335,N_11968);
or U18307 (N_18307,N_13632,N_12918);
and U18308 (N_18308,N_11351,N_14221);
xnor U18309 (N_18309,N_14531,N_14902);
and U18310 (N_18310,N_14346,N_14245);
xor U18311 (N_18311,N_10287,N_11046);
or U18312 (N_18312,N_11221,N_14757);
or U18313 (N_18313,N_14495,N_11121);
and U18314 (N_18314,N_11352,N_13641);
nor U18315 (N_18315,N_13386,N_12072);
or U18316 (N_18316,N_12857,N_12052);
or U18317 (N_18317,N_12526,N_13606);
or U18318 (N_18318,N_14021,N_11284);
nor U18319 (N_18319,N_11496,N_14794);
or U18320 (N_18320,N_10559,N_12595);
and U18321 (N_18321,N_14527,N_14628);
or U18322 (N_18322,N_11487,N_13853);
nand U18323 (N_18323,N_10979,N_13203);
xnor U18324 (N_18324,N_12032,N_10929);
and U18325 (N_18325,N_11971,N_11151);
or U18326 (N_18326,N_10745,N_11343);
xnor U18327 (N_18327,N_14855,N_14661);
nand U18328 (N_18328,N_14530,N_13751);
nand U18329 (N_18329,N_12653,N_12580);
xnor U18330 (N_18330,N_11852,N_10143);
xnor U18331 (N_18331,N_10758,N_10439);
or U18332 (N_18332,N_13905,N_11557);
nor U18333 (N_18333,N_11663,N_11210);
or U18334 (N_18334,N_12133,N_11504);
or U18335 (N_18335,N_10914,N_12360);
or U18336 (N_18336,N_14183,N_13999);
nand U18337 (N_18337,N_10078,N_13939);
or U18338 (N_18338,N_14351,N_12896);
nand U18339 (N_18339,N_14266,N_12509);
xor U18340 (N_18340,N_11209,N_10761);
and U18341 (N_18341,N_11872,N_13754);
nor U18342 (N_18342,N_11660,N_10479);
and U18343 (N_18343,N_10911,N_11239);
xor U18344 (N_18344,N_11148,N_13919);
nand U18345 (N_18345,N_12587,N_12223);
xnor U18346 (N_18346,N_14136,N_12090);
nor U18347 (N_18347,N_14179,N_12221);
xnor U18348 (N_18348,N_12879,N_14601);
and U18349 (N_18349,N_12306,N_14981);
or U18350 (N_18350,N_14419,N_11483);
or U18351 (N_18351,N_11231,N_14117);
nor U18352 (N_18352,N_11020,N_12246);
xor U18353 (N_18353,N_13692,N_12688);
xnor U18354 (N_18354,N_11148,N_11447);
or U18355 (N_18355,N_13887,N_10274);
xnor U18356 (N_18356,N_14821,N_12944);
xor U18357 (N_18357,N_12541,N_10460);
and U18358 (N_18358,N_12415,N_12672);
and U18359 (N_18359,N_13946,N_11230);
and U18360 (N_18360,N_12178,N_13073);
nand U18361 (N_18361,N_14793,N_13499);
and U18362 (N_18362,N_14113,N_14806);
xor U18363 (N_18363,N_13038,N_11483);
and U18364 (N_18364,N_11648,N_10759);
nand U18365 (N_18365,N_11290,N_10006);
nand U18366 (N_18366,N_13803,N_11116);
or U18367 (N_18367,N_11202,N_10624);
nor U18368 (N_18368,N_10794,N_14943);
xnor U18369 (N_18369,N_10749,N_12490);
or U18370 (N_18370,N_13527,N_10685);
xnor U18371 (N_18371,N_13557,N_13483);
and U18372 (N_18372,N_11330,N_14233);
nand U18373 (N_18373,N_10487,N_11293);
or U18374 (N_18374,N_14509,N_14614);
nand U18375 (N_18375,N_11715,N_14500);
and U18376 (N_18376,N_11493,N_11119);
nor U18377 (N_18377,N_10467,N_14820);
or U18378 (N_18378,N_13134,N_13132);
xnor U18379 (N_18379,N_13041,N_14719);
nand U18380 (N_18380,N_13179,N_11342);
or U18381 (N_18381,N_12614,N_12192);
and U18382 (N_18382,N_14252,N_10511);
nor U18383 (N_18383,N_12363,N_12056);
nor U18384 (N_18384,N_12692,N_14413);
xnor U18385 (N_18385,N_13157,N_13957);
or U18386 (N_18386,N_10272,N_12699);
or U18387 (N_18387,N_12039,N_14858);
or U18388 (N_18388,N_12970,N_10754);
and U18389 (N_18389,N_13263,N_11781);
nand U18390 (N_18390,N_10955,N_12229);
nor U18391 (N_18391,N_14893,N_11658);
nor U18392 (N_18392,N_12930,N_12873);
and U18393 (N_18393,N_14427,N_14571);
xor U18394 (N_18394,N_11724,N_10119);
nor U18395 (N_18395,N_11260,N_13882);
xnor U18396 (N_18396,N_12655,N_12455);
and U18397 (N_18397,N_11106,N_14400);
nor U18398 (N_18398,N_14606,N_13193);
xnor U18399 (N_18399,N_13950,N_13410);
and U18400 (N_18400,N_12573,N_11250);
nor U18401 (N_18401,N_12238,N_12461);
nand U18402 (N_18402,N_10622,N_13284);
or U18403 (N_18403,N_10230,N_13543);
nand U18404 (N_18404,N_14594,N_11882);
or U18405 (N_18405,N_13878,N_11215);
nor U18406 (N_18406,N_14536,N_12203);
xor U18407 (N_18407,N_11776,N_14550);
and U18408 (N_18408,N_12467,N_13301);
nor U18409 (N_18409,N_10951,N_12166);
and U18410 (N_18410,N_13896,N_14985);
nand U18411 (N_18411,N_14413,N_12826);
nor U18412 (N_18412,N_14629,N_11974);
or U18413 (N_18413,N_12506,N_14463);
nor U18414 (N_18414,N_11199,N_12619);
xor U18415 (N_18415,N_13903,N_12056);
xnor U18416 (N_18416,N_11034,N_14401);
nand U18417 (N_18417,N_10436,N_12334);
nand U18418 (N_18418,N_13190,N_13975);
xnor U18419 (N_18419,N_13287,N_10721);
and U18420 (N_18420,N_12078,N_11341);
xor U18421 (N_18421,N_11416,N_11715);
and U18422 (N_18422,N_13803,N_13607);
nand U18423 (N_18423,N_13870,N_12217);
nand U18424 (N_18424,N_10958,N_12251);
and U18425 (N_18425,N_14913,N_12124);
xor U18426 (N_18426,N_10219,N_11276);
and U18427 (N_18427,N_11753,N_13766);
nor U18428 (N_18428,N_13470,N_13600);
xor U18429 (N_18429,N_11932,N_10135);
or U18430 (N_18430,N_13899,N_11188);
xor U18431 (N_18431,N_10064,N_12788);
or U18432 (N_18432,N_13737,N_12030);
nor U18433 (N_18433,N_13662,N_14355);
xor U18434 (N_18434,N_14173,N_13976);
and U18435 (N_18435,N_13989,N_11607);
xnor U18436 (N_18436,N_11361,N_11321);
xor U18437 (N_18437,N_14084,N_10083);
xnor U18438 (N_18438,N_13739,N_14878);
nand U18439 (N_18439,N_13302,N_10379);
nor U18440 (N_18440,N_11098,N_12784);
nand U18441 (N_18441,N_13770,N_10889);
or U18442 (N_18442,N_12070,N_14846);
or U18443 (N_18443,N_12756,N_14942);
or U18444 (N_18444,N_12684,N_10191);
xnor U18445 (N_18445,N_11300,N_13706);
or U18446 (N_18446,N_10279,N_14412);
nand U18447 (N_18447,N_12416,N_10084);
nor U18448 (N_18448,N_14617,N_11003);
nor U18449 (N_18449,N_11008,N_10636);
xor U18450 (N_18450,N_14345,N_14242);
and U18451 (N_18451,N_11630,N_14160);
nand U18452 (N_18452,N_10142,N_11582);
and U18453 (N_18453,N_13697,N_10574);
xnor U18454 (N_18454,N_14532,N_10420);
nor U18455 (N_18455,N_13134,N_12386);
nor U18456 (N_18456,N_11273,N_11138);
and U18457 (N_18457,N_11969,N_11741);
nor U18458 (N_18458,N_11980,N_12132);
or U18459 (N_18459,N_11576,N_13862);
nor U18460 (N_18460,N_12789,N_13713);
nand U18461 (N_18461,N_12373,N_13383);
xor U18462 (N_18462,N_12849,N_12619);
xor U18463 (N_18463,N_11521,N_11064);
nor U18464 (N_18464,N_12984,N_14293);
xor U18465 (N_18465,N_12785,N_12708);
xor U18466 (N_18466,N_13093,N_11551);
or U18467 (N_18467,N_12281,N_13180);
or U18468 (N_18468,N_14302,N_11254);
nand U18469 (N_18469,N_10107,N_11140);
nand U18470 (N_18470,N_12431,N_12712);
xnor U18471 (N_18471,N_10624,N_10711);
or U18472 (N_18472,N_11825,N_13237);
or U18473 (N_18473,N_11052,N_11821);
and U18474 (N_18474,N_10733,N_11899);
nand U18475 (N_18475,N_12008,N_13393);
and U18476 (N_18476,N_11027,N_10961);
nor U18477 (N_18477,N_12682,N_13487);
xnor U18478 (N_18478,N_10477,N_13768);
xnor U18479 (N_18479,N_14945,N_14131);
and U18480 (N_18480,N_12447,N_13625);
nor U18481 (N_18481,N_14866,N_13019);
nand U18482 (N_18482,N_14487,N_13471);
and U18483 (N_18483,N_12112,N_10742);
xor U18484 (N_18484,N_13433,N_11703);
xor U18485 (N_18485,N_14869,N_10681);
nand U18486 (N_18486,N_10856,N_12299);
and U18487 (N_18487,N_13947,N_14209);
or U18488 (N_18488,N_13545,N_12701);
or U18489 (N_18489,N_14235,N_10809);
and U18490 (N_18490,N_11723,N_11528);
xor U18491 (N_18491,N_11036,N_12601);
nand U18492 (N_18492,N_10666,N_10601);
and U18493 (N_18493,N_11747,N_14011);
xor U18494 (N_18494,N_10388,N_11377);
xor U18495 (N_18495,N_10407,N_13318);
xor U18496 (N_18496,N_14007,N_13739);
or U18497 (N_18497,N_13157,N_11125);
nand U18498 (N_18498,N_13880,N_13321);
xor U18499 (N_18499,N_14609,N_14168);
nand U18500 (N_18500,N_12340,N_12501);
nand U18501 (N_18501,N_10957,N_12055);
xnor U18502 (N_18502,N_11624,N_14202);
nand U18503 (N_18503,N_13276,N_13805);
or U18504 (N_18504,N_14276,N_11096);
or U18505 (N_18505,N_12970,N_10376);
nor U18506 (N_18506,N_10926,N_11578);
xor U18507 (N_18507,N_12458,N_13188);
and U18508 (N_18508,N_11666,N_13397);
nor U18509 (N_18509,N_14539,N_13461);
xor U18510 (N_18510,N_11934,N_14829);
and U18511 (N_18511,N_11446,N_12135);
nand U18512 (N_18512,N_13396,N_13616);
or U18513 (N_18513,N_11601,N_10220);
and U18514 (N_18514,N_11000,N_12953);
nand U18515 (N_18515,N_12606,N_12675);
or U18516 (N_18516,N_10890,N_11959);
or U18517 (N_18517,N_13255,N_10813);
or U18518 (N_18518,N_14607,N_10216);
and U18519 (N_18519,N_12973,N_14225);
xnor U18520 (N_18520,N_13939,N_10626);
or U18521 (N_18521,N_12037,N_13116);
nor U18522 (N_18522,N_14835,N_12568);
nand U18523 (N_18523,N_12894,N_10303);
and U18524 (N_18524,N_13916,N_14211);
and U18525 (N_18525,N_11471,N_13779);
nand U18526 (N_18526,N_14176,N_12527);
and U18527 (N_18527,N_10072,N_14817);
or U18528 (N_18528,N_12200,N_12941);
nor U18529 (N_18529,N_11045,N_13187);
or U18530 (N_18530,N_11668,N_10812);
xnor U18531 (N_18531,N_10345,N_14257);
and U18532 (N_18532,N_13433,N_13542);
and U18533 (N_18533,N_10319,N_13103);
or U18534 (N_18534,N_13762,N_13201);
nor U18535 (N_18535,N_12374,N_13336);
nand U18536 (N_18536,N_10564,N_14760);
or U18537 (N_18537,N_12741,N_11750);
xor U18538 (N_18538,N_10868,N_14768);
nor U18539 (N_18539,N_14435,N_10677);
or U18540 (N_18540,N_12127,N_12632);
or U18541 (N_18541,N_13376,N_11194);
nor U18542 (N_18542,N_13123,N_13900);
or U18543 (N_18543,N_13187,N_11878);
xnor U18544 (N_18544,N_12399,N_11687);
xor U18545 (N_18545,N_14851,N_12680);
xnor U18546 (N_18546,N_12714,N_14357);
and U18547 (N_18547,N_14517,N_11152);
and U18548 (N_18548,N_14460,N_10576);
nand U18549 (N_18549,N_10073,N_12615);
or U18550 (N_18550,N_13547,N_13561);
nor U18551 (N_18551,N_12015,N_13063);
nand U18552 (N_18552,N_10538,N_13246);
or U18553 (N_18553,N_14863,N_11707);
xor U18554 (N_18554,N_12801,N_11225);
nor U18555 (N_18555,N_14587,N_12909);
nand U18556 (N_18556,N_12552,N_10900);
nor U18557 (N_18557,N_11831,N_13238);
and U18558 (N_18558,N_11336,N_12586);
nor U18559 (N_18559,N_13666,N_14867);
xnor U18560 (N_18560,N_11706,N_10240);
xor U18561 (N_18561,N_14077,N_10192);
or U18562 (N_18562,N_13617,N_10593);
nor U18563 (N_18563,N_13593,N_11557);
xnor U18564 (N_18564,N_12963,N_11269);
and U18565 (N_18565,N_11726,N_13736);
xor U18566 (N_18566,N_14863,N_13125);
and U18567 (N_18567,N_14952,N_13404);
nor U18568 (N_18568,N_13300,N_10559);
nand U18569 (N_18569,N_14133,N_13697);
and U18570 (N_18570,N_13212,N_14412);
and U18571 (N_18571,N_10129,N_11471);
nor U18572 (N_18572,N_10070,N_11577);
xnor U18573 (N_18573,N_13856,N_10460);
nor U18574 (N_18574,N_11973,N_12385);
xor U18575 (N_18575,N_11259,N_10918);
xor U18576 (N_18576,N_14345,N_10820);
xor U18577 (N_18577,N_10983,N_11324);
xnor U18578 (N_18578,N_11959,N_12074);
and U18579 (N_18579,N_12167,N_10611);
nor U18580 (N_18580,N_12061,N_10284);
nor U18581 (N_18581,N_11637,N_13993);
and U18582 (N_18582,N_13402,N_10445);
nor U18583 (N_18583,N_10402,N_12483);
nor U18584 (N_18584,N_10080,N_12746);
xor U18585 (N_18585,N_10254,N_10626);
nand U18586 (N_18586,N_13855,N_14593);
nor U18587 (N_18587,N_11099,N_13647);
nor U18588 (N_18588,N_13773,N_12477);
or U18589 (N_18589,N_12009,N_11459);
nand U18590 (N_18590,N_13284,N_10084);
nor U18591 (N_18591,N_10965,N_13706);
or U18592 (N_18592,N_14510,N_12480);
and U18593 (N_18593,N_12225,N_11393);
nand U18594 (N_18594,N_11342,N_11480);
xnor U18595 (N_18595,N_12450,N_10013);
or U18596 (N_18596,N_11458,N_10569);
nor U18597 (N_18597,N_11456,N_11666);
and U18598 (N_18598,N_14310,N_14242);
xnor U18599 (N_18599,N_13446,N_14750);
xor U18600 (N_18600,N_13930,N_12971);
and U18601 (N_18601,N_14478,N_13027);
nand U18602 (N_18602,N_11872,N_11632);
nand U18603 (N_18603,N_13146,N_13007);
nor U18604 (N_18604,N_11261,N_14074);
nand U18605 (N_18605,N_14910,N_13128);
or U18606 (N_18606,N_11926,N_10859);
and U18607 (N_18607,N_12809,N_14698);
xnor U18608 (N_18608,N_13958,N_14903);
and U18609 (N_18609,N_12954,N_11944);
nor U18610 (N_18610,N_13730,N_10998);
or U18611 (N_18611,N_13654,N_14508);
and U18612 (N_18612,N_12573,N_11391);
xor U18613 (N_18613,N_12084,N_14213);
nor U18614 (N_18614,N_12449,N_14927);
xnor U18615 (N_18615,N_14107,N_13004);
and U18616 (N_18616,N_14080,N_13280);
nor U18617 (N_18617,N_10888,N_10373);
nand U18618 (N_18618,N_10602,N_14548);
and U18619 (N_18619,N_13138,N_12072);
or U18620 (N_18620,N_10518,N_11004);
and U18621 (N_18621,N_10520,N_10984);
and U18622 (N_18622,N_10330,N_14348);
and U18623 (N_18623,N_10654,N_12099);
nand U18624 (N_18624,N_12119,N_11322);
nand U18625 (N_18625,N_10591,N_13930);
nor U18626 (N_18626,N_13264,N_12878);
xnor U18627 (N_18627,N_13927,N_12875);
nor U18628 (N_18628,N_13765,N_12785);
xor U18629 (N_18629,N_10939,N_10838);
and U18630 (N_18630,N_14534,N_12221);
nor U18631 (N_18631,N_10296,N_11108);
xnor U18632 (N_18632,N_10810,N_11099);
xor U18633 (N_18633,N_11245,N_13000);
or U18634 (N_18634,N_11611,N_13928);
nor U18635 (N_18635,N_12289,N_14653);
nand U18636 (N_18636,N_14022,N_10328);
nand U18637 (N_18637,N_13290,N_14628);
nor U18638 (N_18638,N_11058,N_10181);
nor U18639 (N_18639,N_13888,N_12160);
xor U18640 (N_18640,N_10359,N_13702);
nand U18641 (N_18641,N_12687,N_14792);
and U18642 (N_18642,N_13246,N_10932);
nor U18643 (N_18643,N_10503,N_11020);
nand U18644 (N_18644,N_13973,N_11739);
and U18645 (N_18645,N_14442,N_12133);
nand U18646 (N_18646,N_11757,N_14719);
xor U18647 (N_18647,N_11697,N_13077);
xnor U18648 (N_18648,N_13927,N_14753);
nor U18649 (N_18649,N_10399,N_12511);
nor U18650 (N_18650,N_14181,N_14864);
xnor U18651 (N_18651,N_10131,N_12466);
or U18652 (N_18652,N_11809,N_10845);
or U18653 (N_18653,N_11573,N_12434);
or U18654 (N_18654,N_14589,N_13979);
xnor U18655 (N_18655,N_10034,N_14434);
or U18656 (N_18656,N_11995,N_12112);
nor U18657 (N_18657,N_13947,N_10904);
nand U18658 (N_18658,N_12771,N_13248);
nor U18659 (N_18659,N_12156,N_13005);
nor U18660 (N_18660,N_12843,N_12892);
or U18661 (N_18661,N_10562,N_14134);
xnor U18662 (N_18662,N_12018,N_12156);
nand U18663 (N_18663,N_10533,N_11481);
nand U18664 (N_18664,N_14967,N_14634);
xnor U18665 (N_18665,N_14409,N_10869);
xor U18666 (N_18666,N_14648,N_11582);
or U18667 (N_18667,N_13394,N_11240);
or U18668 (N_18668,N_12767,N_14961);
or U18669 (N_18669,N_11991,N_13215);
nand U18670 (N_18670,N_12226,N_14057);
and U18671 (N_18671,N_14999,N_14655);
nand U18672 (N_18672,N_14380,N_13711);
or U18673 (N_18673,N_11264,N_14282);
and U18674 (N_18674,N_14045,N_12470);
xor U18675 (N_18675,N_14707,N_12844);
and U18676 (N_18676,N_11810,N_13042);
or U18677 (N_18677,N_13829,N_13170);
nand U18678 (N_18678,N_11081,N_10669);
xor U18679 (N_18679,N_11253,N_10943);
or U18680 (N_18680,N_12124,N_12621);
and U18681 (N_18681,N_13863,N_12083);
or U18682 (N_18682,N_11776,N_14527);
xor U18683 (N_18683,N_14021,N_13827);
and U18684 (N_18684,N_14005,N_13823);
xor U18685 (N_18685,N_13750,N_11445);
nand U18686 (N_18686,N_14090,N_11925);
and U18687 (N_18687,N_13031,N_14773);
nand U18688 (N_18688,N_11151,N_14634);
xor U18689 (N_18689,N_13853,N_10552);
nor U18690 (N_18690,N_13196,N_13427);
and U18691 (N_18691,N_10644,N_10802);
or U18692 (N_18692,N_14584,N_11058);
xnor U18693 (N_18693,N_10540,N_13657);
or U18694 (N_18694,N_13647,N_10160);
nand U18695 (N_18695,N_13757,N_13329);
nor U18696 (N_18696,N_14834,N_11801);
xnor U18697 (N_18697,N_12993,N_13958);
nor U18698 (N_18698,N_12311,N_12176);
and U18699 (N_18699,N_12332,N_14212);
xnor U18700 (N_18700,N_11931,N_10788);
nand U18701 (N_18701,N_10454,N_14977);
and U18702 (N_18702,N_13192,N_13800);
xnor U18703 (N_18703,N_11215,N_13679);
nand U18704 (N_18704,N_14468,N_13537);
and U18705 (N_18705,N_14247,N_14043);
nand U18706 (N_18706,N_12809,N_14399);
nor U18707 (N_18707,N_14814,N_11011);
xor U18708 (N_18708,N_13053,N_10510);
and U18709 (N_18709,N_12057,N_14526);
nand U18710 (N_18710,N_12258,N_12110);
nor U18711 (N_18711,N_11547,N_13298);
nor U18712 (N_18712,N_11697,N_10265);
xnor U18713 (N_18713,N_13401,N_12928);
or U18714 (N_18714,N_13174,N_13772);
or U18715 (N_18715,N_13215,N_10837);
xor U18716 (N_18716,N_13693,N_14383);
nand U18717 (N_18717,N_11235,N_13088);
nand U18718 (N_18718,N_10715,N_12676);
or U18719 (N_18719,N_10915,N_12910);
xnor U18720 (N_18720,N_12236,N_14351);
and U18721 (N_18721,N_10512,N_12894);
nor U18722 (N_18722,N_10290,N_12493);
and U18723 (N_18723,N_12708,N_10706);
xnor U18724 (N_18724,N_10015,N_13747);
xnor U18725 (N_18725,N_12401,N_13088);
nand U18726 (N_18726,N_11477,N_14158);
or U18727 (N_18727,N_12060,N_10470);
and U18728 (N_18728,N_14140,N_13097);
nor U18729 (N_18729,N_10889,N_13330);
nand U18730 (N_18730,N_10707,N_11718);
xor U18731 (N_18731,N_14476,N_12541);
xor U18732 (N_18732,N_11898,N_12111);
or U18733 (N_18733,N_14176,N_13647);
nand U18734 (N_18734,N_10730,N_11724);
nor U18735 (N_18735,N_11433,N_12126);
or U18736 (N_18736,N_11350,N_14181);
nand U18737 (N_18737,N_10147,N_12437);
nor U18738 (N_18738,N_10181,N_14176);
and U18739 (N_18739,N_12565,N_11755);
xnor U18740 (N_18740,N_14421,N_10801);
nor U18741 (N_18741,N_10167,N_13051);
nor U18742 (N_18742,N_14485,N_10150);
and U18743 (N_18743,N_14897,N_14392);
and U18744 (N_18744,N_12550,N_13205);
nor U18745 (N_18745,N_10845,N_13543);
xor U18746 (N_18746,N_11962,N_10973);
and U18747 (N_18747,N_11768,N_12390);
nor U18748 (N_18748,N_12307,N_14704);
or U18749 (N_18749,N_11936,N_12519);
xor U18750 (N_18750,N_13470,N_14578);
or U18751 (N_18751,N_12047,N_14429);
and U18752 (N_18752,N_12264,N_12965);
xnor U18753 (N_18753,N_10463,N_12053);
nand U18754 (N_18754,N_12581,N_11129);
xnor U18755 (N_18755,N_13919,N_14442);
or U18756 (N_18756,N_10576,N_14398);
and U18757 (N_18757,N_10657,N_14266);
xnor U18758 (N_18758,N_11145,N_11537);
nor U18759 (N_18759,N_11573,N_13384);
nor U18760 (N_18760,N_14521,N_11061);
nor U18761 (N_18761,N_13573,N_10760);
xnor U18762 (N_18762,N_10746,N_13315);
nand U18763 (N_18763,N_11104,N_13057);
xnor U18764 (N_18764,N_14994,N_10747);
nand U18765 (N_18765,N_14638,N_11517);
nand U18766 (N_18766,N_11049,N_13429);
nand U18767 (N_18767,N_13659,N_11697);
xor U18768 (N_18768,N_13234,N_10164);
xor U18769 (N_18769,N_11154,N_11429);
nand U18770 (N_18770,N_10187,N_13246);
xnor U18771 (N_18771,N_10628,N_11695);
nand U18772 (N_18772,N_14984,N_14003);
or U18773 (N_18773,N_13967,N_12368);
nand U18774 (N_18774,N_14035,N_10802);
xor U18775 (N_18775,N_13039,N_11679);
nor U18776 (N_18776,N_13126,N_10631);
nor U18777 (N_18777,N_12263,N_11651);
xor U18778 (N_18778,N_12288,N_13928);
nor U18779 (N_18779,N_10563,N_14393);
nor U18780 (N_18780,N_11082,N_11564);
or U18781 (N_18781,N_13901,N_10623);
or U18782 (N_18782,N_13546,N_11666);
xor U18783 (N_18783,N_10770,N_12227);
or U18784 (N_18784,N_14792,N_11894);
or U18785 (N_18785,N_14853,N_10998);
nand U18786 (N_18786,N_10597,N_10129);
or U18787 (N_18787,N_10191,N_10994);
and U18788 (N_18788,N_12965,N_10709);
nor U18789 (N_18789,N_13508,N_14325);
nand U18790 (N_18790,N_13466,N_10126);
and U18791 (N_18791,N_13200,N_12877);
nor U18792 (N_18792,N_11482,N_12688);
xnor U18793 (N_18793,N_12128,N_12901);
and U18794 (N_18794,N_12266,N_10261);
nand U18795 (N_18795,N_12064,N_13820);
or U18796 (N_18796,N_13699,N_10030);
nor U18797 (N_18797,N_10051,N_14923);
nand U18798 (N_18798,N_11709,N_11570);
nand U18799 (N_18799,N_10225,N_10929);
and U18800 (N_18800,N_14644,N_12037);
nor U18801 (N_18801,N_12523,N_14077);
or U18802 (N_18802,N_10621,N_12623);
xor U18803 (N_18803,N_10155,N_13905);
and U18804 (N_18804,N_12807,N_10770);
and U18805 (N_18805,N_10482,N_13186);
and U18806 (N_18806,N_14151,N_11001);
or U18807 (N_18807,N_12032,N_10049);
or U18808 (N_18808,N_11659,N_10570);
and U18809 (N_18809,N_14248,N_12295);
nand U18810 (N_18810,N_11066,N_14325);
nor U18811 (N_18811,N_13269,N_13855);
nand U18812 (N_18812,N_10141,N_11203);
nand U18813 (N_18813,N_13049,N_13187);
or U18814 (N_18814,N_11331,N_11942);
and U18815 (N_18815,N_14690,N_11635);
nor U18816 (N_18816,N_11287,N_12975);
or U18817 (N_18817,N_14544,N_13735);
xor U18818 (N_18818,N_12044,N_11064);
and U18819 (N_18819,N_10740,N_10546);
xor U18820 (N_18820,N_10328,N_12906);
nor U18821 (N_18821,N_11207,N_10016);
xnor U18822 (N_18822,N_11348,N_13518);
or U18823 (N_18823,N_10622,N_12481);
and U18824 (N_18824,N_14365,N_14787);
xnor U18825 (N_18825,N_13736,N_13878);
and U18826 (N_18826,N_11323,N_14290);
and U18827 (N_18827,N_12429,N_14270);
or U18828 (N_18828,N_10672,N_10851);
xor U18829 (N_18829,N_14440,N_10168);
nor U18830 (N_18830,N_10251,N_11048);
or U18831 (N_18831,N_13772,N_13865);
nor U18832 (N_18832,N_12704,N_11617);
and U18833 (N_18833,N_10719,N_11000);
and U18834 (N_18834,N_10186,N_12436);
nand U18835 (N_18835,N_10166,N_12345);
or U18836 (N_18836,N_11344,N_12462);
nand U18837 (N_18837,N_12811,N_11725);
nor U18838 (N_18838,N_13172,N_12537);
nand U18839 (N_18839,N_11596,N_13647);
nand U18840 (N_18840,N_14131,N_10716);
or U18841 (N_18841,N_11125,N_12181);
nor U18842 (N_18842,N_14961,N_11298);
nand U18843 (N_18843,N_10840,N_10850);
xor U18844 (N_18844,N_13472,N_10166);
xor U18845 (N_18845,N_14198,N_11378);
or U18846 (N_18846,N_11618,N_13779);
and U18847 (N_18847,N_12097,N_13084);
xnor U18848 (N_18848,N_13917,N_10862);
or U18849 (N_18849,N_10772,N_10178);
nor U18850 (N_18850,N_12445,N_14016);
nor U18851 (N_18851,N_13923,N_12259);
or U18852 (N_18852,N_11834,N_13857);
nand U18853 (N_18853,N_14882,N_12884);
nand U18854 (N_18854,N_11184,N_14734);
nand U18855 (N_18855,N_10704,N_10378);
nand U18856 (N_18856,N_12616,N_11606);
and U18857 (N_18857,N_10044,N_11578);
xor U18858 (N_18858,N_12875,N_13494);
or U18859 (N_18859,N_11413,N_13587);
nor U18860 (N_18860,N_14841,N_11211);
and U18861 (N_18861,N_13463,N_11417);
xor U18862 (N_18862,N_12537,N_14593);
nand U18863 (N_18863,N_12988,N_11409);
nor U18864 (N_18864,N_13577,N_12407);
nor U18865 (N_18865,N_12714,N_10321);
nand U18866 (N_18866,N_11281,N_10208);
or U18867 (N_18867,N_12309,N_14914);
and U18868 (N_18868,N_14120,N_14577);
nor U18869 (N_18869,N_14954,N_11157);
and U18870 (N_18870,N_10921,N_14510);
or U18871 (N_18871,N_13869,N_12185);
nand U18872 (N_18872,N_11159,N_14810);
nor U18873 (N_18873,N_12158,N_11427);
xor U18874 (N_18874,N_10147,N_14662);
nand U18875 (N_18875,N_11072,N_14113);
nor U18876 (N_18876,N_14370,N_10043);
or U18877 (N_18877,N_12491,N_13441);
nor U18878 (N_18878,N_11748,N_14195);
or U18879 (N_18879,N_10307,N_10444);
nand U18880 (N_18880,N_12817,N_14522);
and U18881 (N_18881,N_10784,N_10918);
xor U18882 (N_18882,N_10447,N_10059);
xor U18883 (N_18883,N_12890,N_10149);
nor U18884 (N_18884,N_14193,N_11120);
xor U18885 (N_18885,N_11581,N_14758);
nor U18886 (N_18886,N_13313,N_13844);
nand U18887 (N_18887,N_13368,N_13692);
or U18888 (N_18888,N_11603,N_10947);
xor U18889 (N_18889,N_11845,N_13552);
or U18890 (N_18890,N_10038,N_13701);
or U18891 (N_18891,N_12729,N_13980);
nand U18892 (N_18892,N_13263,N_14380);
nor U18893 (N_18893,N_12112,N_12485);
and U18894 (N_18894,N_14754,N_13914);
xnor U18895 (N_18895,N_12990,N_10314);
or U18896 (N_18896,N_10488,N_14696);
and U18897 (N_18897,N_13170,N_11471);
nor U18898 (N_18898,N_13171,N_10577);
and U18899 (N_18899,N_13206,N_12622);
nor U18900 (N_18900,N_14460,N_12507);
and U18901 (N_18901,N_12010,N_11699);
or U18902 (N_18902,N_11338,N_12307);
or U18903 (N_18903,N_13792,N_12482);
nand U18904 (N_18904,N_11720,N_11333);
xor U18905 (N_18905,N_12938,N_11480);
xnor U18906 (N_18906,N_14941,N_14966);
and U18907 (N_18907,N_11634,N_12694);
and U18908 (N_18908,N_12651,N_14325);
nand U18909 (N_18909,N_14447,N_11426);
and U18910 (N_18910,N_13315,N_13895);
or U18911 (N_18911,N_13665,N_11277);
or U18912 (N_18912,N_12607,N_12251);
xnor U18913 (N_18913,N_11496,N_12402);
and U18914 (N_18914,N_11399,N_12665);
xnor U18915 (N_18915,N_13993,N_10827);
nand U18916 (N_18916,N_11635,N_13673);
and U18917 (N_18917,N_12288,N_10361);
and U18918 (N_18918,N_12517,N_12329);
or U18919 (N_18919,N_14782,N_13892);
and U18920 (N_18920,N_14430,N_11301);
xnor U18921 (N_18921,N_10336,N_14645);
nand U18922 (N_18922,N_11448,N_10981);
xor U18923 (N_18923,N_13537,N_14893);
xor U18924 (N_18924,N_12874,N_12904);
or U18925 (N_18925,N_14679,N_12050);
and U18926 (N_18926,N_11936,N_14251);
and U18927 (N_18927,N_12297,N_13656);
and U18928 (N_18928,N_10238,N_13454);
nand U18929 (N_18929,N_14432,N_12842);
nor U18930 (N_18930,N_14944,N_10462);
nand U18931 (N_18931,N_11648,N_10453);
xor U18932 (N_18932,N_14456,N_12714);
nor U18933 (N_18933,N_12129,N_10996);
nand U18934 (N_18934,N_11573,N_10483);
nand U18935 (N_18935,N_13700,N_10796);
xor U18936 (N_18936,N_14989,N_12173);
nand U18937 (N_18937,N_14927,N_12814);
nor U18938 (N_18938,N_11881,N_12110);
xor U18939 (N_18939,N_13173,N_13315);
nor U18940 (N_18940,N_14818,N_12986);
or U18941 (N_18941,N_14606,N_13695);
and U18942 (N_18942,N_11063,N_10642);
nor U18943 (N_18943,N_13608,N_11515);
xnor U18944 (N_18944,N_11423,N_14433);
or U18945 (N_18945,N_14151,N_11508);
nand U18946 (N_18946,N_14630,N_12164);
xnor U18947 (N_18947,N_14942,N_11108);
and U18948 (N_18948,N_13381,N_12932);
or U18949 (N_18949,N_12301,N_11284);
nand U18950 (N_18950,N_11219,N_10957);
nand U18951 (N_18951,N_14624,N_13920);
nand U18952 (N_18952,N_11596,N_10369);
nor U18953 (N_18953,N_13945,N_10236);
or U18954 (N_18954,N_11389,N_11814);
nor U18955 (N_18955,N_10559,N_11935);
nand U18956 (N_18956,N_10072,N_10660);
and U18957 (N_18957,N_11765,N_14077);
xnor U18958 (N_18958,N_10545,N_11046);
nor U18959 (N_18959,N_12366,N_12580);
and U18960 (N_18960,N_12612,N_11912);
nand U18961 (N_18961,N_12905,N_10565);
nand U18962 (N_18962,N_13986,N_11898);
nand U18963 (N_18963,N_14272,N_10272);
nand U18964 (N_18964,N_12983,N_14059);
and U18965 (N_18965,N_11866,N_14306);
xnor U18966 (N_18966,N_11632,N_12169);
xor U18967 (N_18967,N_14411,N_14560);
or U18968 (N_18968,N_12652,N_10481);
and U18969 (N_18969,N_12706,N_14919);
or U18970 (N_18970,N_11304,N_10123);
and U18971 (N_18971,N_12473,N_11578);
or U18972 (N_18972,N_11396,N_13930);
or U18973 (N_18973,N_11948,N_10924);
or U18974 (N_18974,N_12507,N_10951);
xor U18975 (N_18975,N_13262,N_13478);
nand U18976 (N_18976,N_11390,N_10007);
or U18977 (N_18977,N_10124,N_14665);
xor U18978 (N_18978,N_13022,N_11206);
and U18979 (N_18979,N_12193,N_11747);
or U18980 (N_18980,N_11627,N_11828);
xnor U18981 (N_18981,N_13613,N_12080);
or U18982 (N_18982,N_12197,N_14732);
nand U18983 (N_18983,N_14247,N_13899);
and U18984 (N_18984,N_12886,N_13751);
and U18985 (N_18985,N_14482,N_11444);
xor U18986 (N_18986,N_12189,N_14529);
nand U18987 (N_18987,N_14845,N_10854);
nor U18988 (N_18988,N_11711,N_10504);
nand U18989 (N_18989,N_12842,N_11007);
nor U18990 (N_18990,N_10561,N_12048);
and U18991 (N_18991,N_10583,N_13016);
nand U18992 (N_18992,N_14416,N_11332);
nor U18993 (N_18993,N_12293,N_12884);
xor U18994 (N_18994,N_11021,N_13277);
nand U18995 (N_18995,N_11530,N_14933);
or U18996 (N_18996,N_13075,N_11620);
or U18997 (N_18997,N_11279,N_13127);
nor U18998 (N_18998,N_11392,N_10675);
nand U18999 (N_18999,N_10154,N_11584);
nor U19000 (N_19000,N_11852,N_13192);
or U19001 (N_19001,N_13802,N_11978);
and U19002 (N_19002,N_13502,N_11717);
or U19003 (N_19003,N_12498,N_10844);
nand U19004 (N_19004,N_11880,N_12499);
nand U19005 (N_19005,N_10384,N_13032);
and U19006 (N_19006,N_10898,N_12911);
nand U19007 (N_19007,N_11774,N_10179);
nor U19008 (N_19008,N_11108,N_12824);
xnor U19009 (N_19009,N_10704,N_13237);
or U19010 (N_19010,N_12692,N_12153);
or U19011 (N_19011,N_12317,N_12294);
nor U19012 (N_19012,N_13866,N_14463);
or U19013 (N_19013,N_12835,N_10386);
or U19014 (N_19014,N_11327,N_10134);
nand U19015 (N_19015,N_11283,N_10821);
and U19016 (N_19016,N_14484,N_11787);
and U19017 (N_19017,N_12765,N_13587);
xor U19018 (N_19018,N_13571,N_10788);
nand U19019 (N_19019,N_14317,N_13594);
xnor U19020 (N_19020,N_14602,N_13308);
nor U19021 (N_19021,N_13985,N_13647);
xor U19022 (N_19022,N_11320,N_12698);
nand U19023 (N_19023,N_14206,N_14117);
and U19024 (N_19024,N_11010,N_11391);
nand U19025 (N_19025,N_10437,N_11993);
nand U19026 (N_19026,N_14692,N_10613);
nor U19027 (N_19027,N_11630,N_14571);
nor U19028 (N_19028,N_12486,N_10944);
xor U19029 (N_19029,N_10217,N_10381);
or U19030 (N_19030,N_11348,N_11811);
or U19031 (N_19031,N_14952,N_10906);
or U19032 (N_19032,N_12456,N_13352);
or U19033 (N_19033,N_14456,N_10298);
and U19034 (N_19034,N_14073,N_13861);
nor U19035 (N_19035,N_13413,N_13084);
or U19036 (N_19036,N_12124,N_12165);
nor U19037 (N_19037,N_14663,N_12999);
nand U19038 (N_19038,N_13155,N_12659);
nand U19039 (N_19039,N_11337,N_11551);
xor U19040 (N_19040,N_14678,N_11647);
nor U19041 (N_19041,N_12473,N_13052);
nor U19042 (N_19042,N_12228,N_12464);
nand U19043 (N_19043,N_14716,N_10041);
nor U19044 (N_19044,N_11976,N_11513);
and U19045 (N_19045,N_12368,N_14743);
xor U19046 (N_19046,N_12062,N_14525);
or U19047 (N_19047,N_11081,N_12394);
nand U19048 (N_19048,N_11088,N_14087);
xor U19049 (N_19049,N_12862,N_12774);
nor U19050 (N_19050,N_13621,N_12757);
nor U19051 (N_19051,N_14841,N_14901);
nand U19052 (N_19052,N_11962,N_13289);
or U19053 (N_19053,N_11750,N_12864);
and U19054 (N_19054,N_14040,N_12963);
and U19055 (N_19055,N_10138,N_11700);
or U19056 (N_19056,N_10474,N_10035);
xor U19057 (N_19057,N_13650,N_11782);
or U19058 (N_19058,N_10654,N_12839);
xor U19059 (N_19059,N_12371,N_10254);
or U19060 (N_19060,N_11512,N_13901);
or U19061 (N_19061,N_11527,N_14100);
and U19062 (N_19062,N_10542,N_13518);
nand U19063 (N_19063,N_11386,N_11832);
or U19064 (N_19064,N_14780,N_11908);
or U19065 (N_19065,N_11293,N_12914);
nand U19066 (N_19066,N_11552,N_14762);
and U19067 (N_19067,N_14493,N_13968);
and U19068 (N_19068,N_12394,N_12123);
and U19069 (N_19069,N_11098,N_11489);
xor U19070 (N_19070,N_12022,N_14777);
xor U19071 (N_19071,N_13903,N_13098);
and U19072 (N_19072,N_14972,N_11193);
and U19073 (N_19073,N_14490,N_11550);
nor U19074 (N_19074,N_12714,N_12808);
nor U19075 (N_19075,N_14070,N_11300);
and U19076 (N_19076,N_10873,N_13869);
nor U19077 (N_19077,N_14579,N_10702);
nor U19078 (N_19078,N_13459,N_12809);
or U19079 (N_19079,N_14774,N_10775);
nand U19080 (N_19080,N_14814,N_14701);
or U19081 (N_19081,N_11759,N_11441);
and U19082 (N_19082,N_12872,N_13223);
or U19083 (N_19083,N_11368,N_10791);
nand U19084 (N_19084,N_11064,N_11206);
nor U19085 (N_19085,N_13978,N_12292);
or U19086 (N_19086,N_14522,N_10309);
nor U19087 (N_19087,N_14967,N_11751);
or U19088 (N_19088,N_14695,N_13546);
xnor U19089 (N_19089,N_10319,N_11646);
and U19090 (N_19090,N_11392,N_12365);
xor U19091 (N_19091,N_14756,N_10142);
and U19092 (N_19092,N_13049,N_10183);
or U19093 (N_19093,N_11210,N_13582);
xnor U19094 (N_19094,N_14746,N_13082);
nor U19095 (N_19095,N_10256,N_12272);
xnor U19096 (N_19096,N_13951,N_12136);
and U19097 (N_19097,N_10081,N_11868);
xnor U19098 (N_19098,N_12249,N_13084);
and U19099 (N_19099,N_14393,N_12865);
nor U19100 (N_19100,N_13738,N_10343);
and U19101 (N_19101,N_12173,N_13101);
xor U19102 (N_19102,N_13271,N_14218);
and U19103 (N_19103,N_14875,N_10785);
nand U19104 (N_19104,N_13952,N_10898);
or U19105 (N_19105,N_12946,N_13447);
nand U19106 (N_19106,N_13613,N_11496);
or U19107 (N_19107,N_11444,N_14529);
nand U19108 (N_19108,N_14728,N_11008);
nor U19109 (N_19109,N_11433,N_11292);
xnor U19110 (N_19110,N_11984,N_14291);
or U19111 (N_19111,N_12074,N_14797);
nand U19112 (N_19112,N_13634,N_12460);
nor U19113 (N_19113,N_10284,N_13026);
xor U19114 (N_19114,N_14104,N_11280);
nand U19115 (N_19115,N_10947,N_11584);
xnor U19116 (N_19116,N_11487,N_10273);
xnor U19117 (N_19117,N_10608,N_10465);
or U19118 (N_19118,N_12016,N_10277);
nand U19119 (N_19119,N_13698,N_10614);
or U19120 (N_19120,N_11813,N_14139);
nand U19121 (N_19121,N_11269,N_14868);
xor U19122 (N_19122,N_13774,N_12665);
xnor U19123 (N_19123,N_13240,N_11646);
nand U19124 (N_19124,N_11409,N_14556);
or U19125 (N_19125,N_10625,N_11615);
or U19126 (N_19126,N_10761,N_14589);
nand U19127 (N_19127,N_11975,N_12821);
and U19128 (N_19128,N_14704,N_12972);
nand U19129 (N_19129,N_10667,N_11124);
nor U19130 (N_19130,N_14625,N_12018);
and U19131 (N_19131,N_12610,N_12995);
or U19132 (N_19132,N_13767,N_10458);
nor U19133 (N_19133,N_12257,N_11416);
and U19134 (N_19134,N_12668,N_11710);
xor U19135 (N_19135,N_14481,N_12353);
nor U19136 (N_19136,N_13730,N_11071);
and U19137 (N_19137,N_11417,N_14873);
or U19138 (N_19138,N_11937,N_14851);
nand U19139 (N_19139,N_13603,N_13156);
and U19140 (N_19140,N_10694,N_12041);
xor U19141 (N_19141,N_11701,N_12377);
nor U19142 (N_19142,N_11340,N_10639);
nand U19143 (N_19143,N_12077,N_10226);
and U19144 (N_19144,N_12449,N_12715);
nor U19145 (N_19145,N_12761,N_14259);
xnor U19146 (N_19146,N_12402,N_12341);
nor U19147 (N_19147,N_14537,N_11917);
or U19148 (N_19148,N_11153,N_11618);
and U19149 (N_19149,N_13660,N_11055);
or U19150 (N_19150,N_14647,N_12463);
nor U19151 (N_19151,N_12735,N_12131);
nor U19152 (N_19152,N_11920,N_12320);
nor U19153 (N_19153,N_13029,N_12536);
nand U19154 (N_19154,N_10257,N_11351);
nand U19155 (N_19155,N_13105,N_11062);
nand U19156 (N_19156,N_12777,N_11227);
xor U19157 (N_19157,N_11882,N_13333);
and U19158 (N_19158,N_14625,N_12805);
or U19159 (N_19159,N_11662,N_11341);
nand U19160 (N_19160,N_11626,N_12076);
xnor U19161 (N_19161,N_12939,N_14668);
nand U19162 (N_19162,N_11953,N_14756);
or U19163 (N_19163,N_13003,N_13488);
xor U19164 (N_19164,N_12541,N_11480);
or U19165 (N_19165,N_14776,N_13319);
xnor U19166 (N_19166,N_11469,N_11647);
or U19167 (N_19167,N_13605,N_10981);
xor U19168 (N_19168,N_12346,N_14644);
and U19169 (N_19169,N_10443,N_13324);
and U19170 (N_19170,N_10721,N_10436);
xnor U19171 (N_19171,N_13572,N_10852);
nand U19172 (N_19172,N_11464,N_10144);
xnor U19173 (N_19173,N_14858,N_10646);
nor U19174 (N_19174,N_14053,N_11799);
xnor U19175 (N_19175,N_11004,N_13203);
and U19176 (N_19176,N_10623,N_13980);
and U19177 (N_19177,N_14002,N_13984);
or U19178 (N_19178,N_12567,N_13542);
nor U19179 (N_19179,N_10083,N_13471);
or U19180 (N_19180,N_12790,N_10370);
nor U19181 (N_19181,N_10530,N_13950);
and U19182 (N_19182,N_10016,N_14840);
nand U19183 (N_19183,N_10334,N_13618);
nor U19184 (N_19184,N_14817,N_10551);
or U19185 (N_19185,N_14348,N_11192);
xnor U19186 (N_19186,N_11121,N_13553);
nand U19187 (N_19187,N_12961,N_11863);
and U19188 (N_19188,N_12855,N_14464);
nand U19189 (N_19189,N_14399,N_13828);
or U19190 (N_19190,N_10482,N_13206);
xor U19191 (N_19191,N_14048,N_13348);
nor U19192 (N_19192,N_14732,N_11098);
xor U19193 (N_19193,N_12750,N_12142);
and U19194 (N_19194,N_11337,N_10408);
nor U19195 (N_19195,N_10298,N_13591);
and U19196 (N_19196,N_14591,N_14803);
xnor U19197 (N_19197,N_10226,N_13159);
and U19198 (N_19198,N_12633,N_12870);
nand U19199 (N_19199,N_14004,N_10539);
nand U19200 (N_19200,N_13823,N_12717);
and U19201 (N_19201,N_13171,N_14335);
and U19202 (N_19202,N_14044,N_12756);
nand U19203 (N_19203,N_12768,N_14233);
and U19204 (N_19204,N_13374,N_10203);
nor U19205 (N_19205,N_11315,N_11394);
nand U19206 (N_19206,N_11588,N_10333);
or U19207 (N_19207,N_12704,N_12307);
nand U19208 (N_19208,N_12754,N_12182);
nor U19209 (N_19209,N_12536,N_10445);
nand U19210 (N_19210,N_12451,N_11700);
and U19211 (N_19211,N_14441,N_11488);
nand U19212 (N_19212,N_13103,N_12777);
nand U19213 (N_19213,N_14172,N_10295);
nand U19214 (N_19214,N_13752,N_12044);
xnor U19215 (N_19215,N_12329,N_12060);
xnor U19216 (N_19216,N_14409,N_11101);
or U19217 (N_19217,N_12379,N_14654);
or U19218 (N_19218,N_10790,N_11824);
nor U19219 (N_19219,N_10123,N_12240);
and U19220 (N_19220,N_12603,N_10109);
and U19221 (N_19221,N_14240,N_12992);
nor U19222 (N_19222,N_12791,N_11803);
or U19223 (N_19223,N_13823,N_10933);
nand U19224 (N_19224,N_10857,N_13016);
nor U19225 (N_19225,N_14647,N_14300);
or U19226 (N_19226,N_14583,N_13265);
nand U19227 (N_19227,N_11814,N_14670);
and U19228 (N_19228,N_11555,N_10101);
or U19229 (N_19229,N_12388,N_12305);
nand U19230 (N_19230,N_13535,N_13427);
nor U19231 (N_19231,N_11422,N_14012);
xor U19232 (N_19232,N_11866,N_12724);
and U19233 (N_19233,N_10527,N_14338);
nand U19234 (N_19234,N_13099,N_14575);
nand U19235 (N_19235,N_10445,N_14136);
xnor U19236 (N_19236,N_10983,N_13318);
and U19237 (N_19237,N_11684,N_12634);
nor U19238 (N_19238,N_10174,N_12705);
or U19239 (N_19239,N_11840,N_14660);
nand U19240 (N_19240,N_10589,N_14481);
nor U19241 (N_19241,N_12490,N_11929);
nor U19242 (N_19242,N_12922,N_11848);
xnor U19243 (N_19243,N_14996,N_11076);
and U19244 (N_19244,N_10601,N_14721);
or U19245 (N_19245,N_12970,N_11788);
nor U19246 (N_19246,N_12666,N_11771);
xnor U19247 (N_19247,N_10738,N_13183);
or U19248 (N_19248,N_11934,N_12126);
or U19249 (N_19249,N_13270,N_10520);
xor U19250 (N_19250,N_12123,N_11037);
xor U19251 (N_19251,N_12197,N_10824);
nor U19252 (N_19252,N_14866,N_12570);
xor U19253 (N_19253,N_11864,N_10138);
and U19254 (N_19254,N_11680,N_12379);
or U19255 (N_19255,N_10663,N_12494);
xor U19256 (N_19256,N_14085,N_13760);
nand U19257 (N_19257,N_13220,N_11830);
or U19258 (N_19258,N_14911,N_13411);
xnor U19259 (N_19259,N_14871,N_12582);
or U19260 (N_19260,N_11217,N_13447);
nand U19261 (N_19261,N_11295,N_11683);
xnor U19262 (N_19262,N_12711,N_12937);
nand U19263 (N_19263,N_13309,N_12145);
xnor U19264 (N_19264,N_11905,N_13466);
nor U19265 (N_19265,N_12107,N_11845);
nand U19266 (N_19266,N_13835,N_11731);
xor U19267 (N_19267,N_14541,N_13546);
xor U19268 (N_19268,N_10273,N_11282);
nand U19269 (N_19269,N_12033,N_14320);
nand U19270 (N_19270,N_12092,N_13563);
nor U19271 (N_19271,N_14619,N_13935);
xnor U19272 (N_19272,N_12128,N_11010);
and U19273 (N_19273,N_11290,N_13416);
xnor U19274 (N_19274,N_14469,N_13550);
xnor U19275 (N_19275,N_10994,N_14640);
xnor U19276 (N_19276,N_13105,N_10687);
xnor U19277 (N_19277,N_10235,N_11644);
or U19278 (N_19278,N_13974,N_10824);
and U19279 (N_19279,N_11639,N_11365);
nand U19280 (N_19280,N_13866,N_11197);
nor U19281 (N_19281,N_14402,N_13280);
nand U19282 (N_19282,N_10155,N_11374);
nor U19283 (N_19283,N_14979,N_13520);
or U19284 (N_19284,N_12424,N_14011);
and U19285 (N_19285,N_10098,N_11148);
nand U19286 (N_19286,N_14567,N_12879);
and U19287 (N_19287,N_13119,N_13294);
nor U19288 (N_19288,N_10222,N_10311);
nor U19289 (N_19289,N_12081,N_10888);
nand U19290 (N_19290,N_14116,N_14259);
xor U19291 (N_19291,N_13440,N_13566);
or U19292 (N_19292,N_13272,N_12173);
and U19293 (N_19293,N_10830,N_10571);
or U19294 (N_19294,N_13336,N_13384);
nand U19295 (N_19295,N_12806,N_11196);
xor U19296 (N_19296,N_12388,N_13949);
xor U19297 (N_19297,N_12315,N_12698);
nand U19298 (N_19298,N_10397,N_10779);
xnor U19299 (N_19299,N_10281,N_12706);
or U19300 (N_19300,N_11536,N_10025);
or U19301 (N_19301,N_14249,N_11545);
nor U19302 (N_19302,N_11820,N_14775);
or U19303 (N_19303,N_10991,N_11855);
or U19304 (N_19304,N_14395,N_13216);
and U19305 (N_19305,N_10318,N_12143);
nor U19306 (N_19306,N_13747,N_13166);
xnor U19307 (N_19307,N_14445,N_11883);
nor U19308 (N_19308,N_10716,N_12904);
nand U19309 (N_19309,N_13585,N_14316);
and U19310 (N_19310,N_13574,N_12874);
nor U19311 (N_19311,N_10175,N_11189);
nand U19312 (N_19312,N_10346,N_14287);
or U19313 (N_19313,N_10629,N_13492);
xor U19314 (N_19314,N_12133,N_14597);
nor U19315 (N_19315,N_11465,N_12038);
or U19316 (N_19316,N_13605,N_12371);
xnor U19317 (N_19317,N_10616,N_14355);
nor U19318 (N_19318,N_10789,N_11000);
nor U19319 (N_19319,N_10162,N_12015);
nand U19320 (N_19320,N_10318,N_13974);
and U19321 (N_19321,N_13851,N_10323);
xor U19322 (N_19322,N_10589,N_12632);
nand U19323 (N_19323,N_13880,N_11464);
xnor U19324 (N_19324,N_10102,N_10112);
and U19325 (N_19325,N_13879,N_13836);
nand U19326 (N_19326,N_14109,N_11831);
and U19327 (N_19327,N_13946,N_10649);
and U19328 (N_19328,N_13703,N_11626);
nand U19329 (N_19329,N_11337,N_11244);
xnor U19330 (N_19330,N_13508,N_13927);
nor U19331 (N_19331,N_13760,N_12422);
xnor U19332 (N_19332,N_12592,N_13317);
nand U19333 (N_19333,N_14332,N_12888);
or U19334 (N_19334,N_13306,N_13886);
nor U19335 (N_19335,N_14458,N_13174);
nand U19336 (N_19336,N_10942,N_10785);
nand U19337 (N_19337,N_11282,N_12453);
nand U19338 (N_19338,N_10655,N_12216);
xnor U19339 (N_19339,N_14837,N_10434);
and U19340 (N_19340,N_10581,N_11412);
and U19341 (N_19341,N_13736,N_13230);
or U19342 (N_19342,N_14828,N_12827);
nor U19343 (N_19343,N_12818,N_10293);
or U19344 (N_19344,N_13340,N_13335);
xnor U19345 (N_19345,N_11074,N_12547);
or U19346 (N_19346,N_12064,N_11808);
nor U19347 (N_19347,N_13185,N_11019);
nand U19348 (N_19348,N_14583,N_13497);
xor U19349 (N_19349,N_13422,N_14321);
xnor U19350 (N_19350,N_10867,N_14968);
xor U19351 (N_19351,N_13154,N_12821);
xnor U19352 (N_19352,N_10358,N_11303);
nand U19353 (N_19353,N_13005,N_14128);
nor U19354 (N_19354,N_13225,N_14057);
or U19355 (N_19355,N_10302,N_10613);
xor U19356 (N_19356,N_11510,N_14852);
or U19357 (N_19357,N_12824,N_14320);
xor U19358 (N_19358,N_13012,N_12213);
and U19359 (N_19359,N_10188,N_14228);
and U19360 (N_19360,N_12387,N_14000);
and U19361 (N_19361,N_12830,N_14484);
nand U19362 (N_19362,N_10080,N_12657);
xnor U19363 (N_19363,N_11864,N_10911);
xor U19364 (N_19364,N_10299,N_12103);
xnor U19365 (N_19365,N_12691,N_13977);
and U19366 (N_19366,N_12868,N_11043);
and U19367 (N_19367,N_14971,N_12239);
and U19368 (N_19368,N_14667,N_13277);
nor U19369 (N_19369,N_12769,N_14553);
or U19370 (N_19370,N_13585,N_10554);
nor U19371 (N_19371,N_12195,N_13612);
xor U19372 (N_19372,N_12410,N_13844);
nand U19373 (N_19373,N_14844,N_10836);
xnor U19374 (N_19374,N_10774,N_11841);
and U19375 (N_19375,N_13649,N_13845);
nor U19376 (N_19376,N_14775,N_11699);
and U19377 (N_19377,N_13882,N_12264);
xnor U19378 (N_19378,N_10997,N_13051);
nor U19379 (N_19379,N_14504,N_10554);
or U19380 (N_19380,N_11685,N_11932);
or U19381 (N_19381,N_13990,N_13090);
nand U19382 (N_19382,N_10758,N_12493);
xor U19383 (N_19383,N_13836,N_10204);
xor U19384 (N_19384,N_11852,N_10986);
nand U19385 (N_19385,N_11808,N_13572);
and U19386 (N_19386,N_10751,N_10963);
and U19387 (N_19387,N_14381,N_12322);
nand U19388 (N_19388,N_12777,N_12639);
or U19389 (N_19389,N_10035,N_11848);
nand U19390 (N_19390,N_11802,N_14836);
nand U19391 (N_19391,N_12360,N_13244);
and U19392 (N_19392,N_12198,N_13111);
or U19393 (N_19393,N_13612,N_13470);
xnor U19394 (N_19394,N_10942,N_14133);
nor U19395 (N_19395,N_11714,N_10804);
xnor U19396 (N_19396,N_13624,N_12525);
or U19397 (N_19397,N_12602,N_10063);
and U19398 (N_19398,N_10894,N_10782);
nor U19399 (N_19399,N_10030,N_10851);
or U19400 (N_19400,N_11583,N_14276);
nand U19401 (N_19401,N_14109,N_11942);
nand U19402 (N_19402,N_11916,N_14252);
or U19403 (N_19403,N_13284,N_13954);
xor U19404 (N_19404,N_12394,N_12293);
nand U19405 (N_19405,N_12302,N_11940);
or U19406 (N_19406,N_11738,N_12424);
xnor U19407 (N_19407,N_10223,N_14165);
xor U19408 (N_19408,N_14307,N_13350);
xor U19409 (N_19409,N_13665,N_11444);
xor U19410 (N_19410,N_12145,N_14345);
nor U19411 (N_19411,N_10915,N_13056);
or U19412 (N_19412,N_13209,N_11377);
nor U19413 (N_19413,N_13475,N_13305);
or U19414 (N_19414,N_10111,N_12540);
nand U19415 (N_19415,N_12216,N_11187);
nor U19416 (N_19416,N_10830,N_11759);
and U19417 (N_19417,N_13890,N_11388);
nor U19418 (N_19418,N_12984,N_12206);
and U19419 (N_19419,N_14804,N_11934);
nor U19420 (N_19420,N_14188,N_11008);
nor U19421 (N_19421,N_11230,N_11983);
xor U19422 (N_19422,N_12684,N_14822);
or U19423 (N_19423,N_10988,N_11141);
nor U19424 (N_19424,N_14838,N_12930);
nor U19425 (N_19425,N_10522,N_13634);
nand U19426 (N_19426,N_13590,N_12278);
xor U19427 (N_19427,N_10672,N_14129);
or U19428 (N_19428,N_11300,N_11327);
nor U19429 (N_19429,N_12705,N_10146);
nor U19430 (N_19430,N_11589,N_11392);
and U19431 (N_19431,N_14475,N_11736);
and U19432 (N_19432,N_14988,N_10727);
nand U19433 (N_19433,N_10086,N_10231);
xnor U19434 (N_19434,N_12793,N_13712);
and U19435 (N_19435,N_13055,N_11499);
xnor U19436 (N_19436,N_13709,N_11033);
and U19437 (N_19437,N_11194,N_11907);
nor U19438 (N_19438,N_12311,N_13856);
nor U19439 (N_19439,N_14794,N_13055);
xnor U19440 (N_19440,N_10168,N_13404);
nor U19441 (N_19441,N_12544,N_14372);
or U19442 (N_19442,N_12868,N_13692);
nor U19443 (N_19443,N_10920,N_13695);
or U19444 (N_19444,N_13033,N_13200);
nand U19445 (N_19445,N_14324,N_14250);
xnor U19446 (N_19446,N_12335,N_14917);
xor U19447 (N_19447,N_10404,N_14746);
xor U19448 (N_19448,N_13503,N_12561);
xnor U19449 (N_19449,N_12867,N_13216);
nor U19450 (N_19450,N_14060,N_10249);
nand U19451 (N_19451,N_11090,N_11753);
xor U19452 (N_19452,N_10807,N_14437);
xnor U19453 (N_19453,N_14399,N_12708);
and U19454 (N_19454,N_10349,N_11838);
nand U19455 (N_19455,N_12501,N_11832);
nor U19456 (N_19456,N_12347,N_14077);
nor U19457 (N_19457,N_12813,N_10212);
nand U19458 (N_19458,N_11590,N_12831);
nand U19459 (N_19459,N_11809,N_10233);
nor U19460 (N_19460,N_14719,N_13722);
or U19461 (N_19461,N_10545,N_14743);
nand U19462 (N_19462,N_11607,N_12242);
xor U19463 (N_19463,N_12012,N_12651);
nand U19464 (N_19464,N_12132,N_13051);
nand U19465 (N_19465,N_10456,N_12683);
xnor U19466 (N_19466,N_12552,N_11538);
and U19467 (N_19467,N_14531,N_14342);
xor U19468 (N_19468,N_12969,N_13485);
or U19469 (N_19469,N_11249,N_12899);
or U19470 (N_19470,N_10867,N_13744);
and U19471 (N_19471,N_13031,N_10832);
and U19472 (N_19472,N_12527,N_13568);
or U19473 (N_19473,N_13483,N_12899);
nor U19474 (N_19474,N_14435,N_14135);
nand U19475 (N_19475,N_13969,N_11136);
xnor U19476 (N_19476,N_10981,N_10992);
or U19477 (N_19477,N_11885,N_14361);
nand U19478 (N_19478,N_14374,N_12461);
nand U19479 (N_19479,N_12763,N_11710);
nor U19480 (N_19480,N_13280,N_12041);
or U19481 (N_19481,N_13963,N_10946);
or U19482 (N_19482,N_14800,N_13413);
nor U19483 (N_19483,N_14836,N_11456);
xor U19484 (N_19484,N_14753,N_11795);
xor U19485 (N_19485,N_12630,N_12599);
nor U19486 (N_19486,N_10898,N_12172);
and U19487 (N_19487,N_14771,N_10400);
nand U19488 (N_19488,N_13073,N_10970);
nor U19489 (N_19489,N_13905,N_11092);
and U19490 (N_19490,N_11984,N_11055);
or U19491 (N_19491,N_11280,N_14807);
xnor U19492 (N_19492,N_13228,N_11660);
nor U19493 (N_19493,N_14735,N_11757);
xnor U19494 (N_19494,N_13275,N_14854);
xor U19495 (N_19495,N_11533,N_10942);
nand U19496 (N_19496,N_13267,N_12706);
or U19497 (N_19497,N_13980,N_12727);
nor U19498 (N_19498,N_14532,N_13424);
or U19499 (N_19499,N_13537,N_13458);
or U19500 (N_19500,N_11320,N_12530);
xor U19501 (N_19501,N_14709,N_11057);
and U19502 (N_19502,N_10591,N_11804);
and U19503 (N_19503,N_10611,N_13959);
or U19504 (N_19504,N_12306,N_12002);
and U19505 (N_19505,N_10660,N_10460);
nand U19506 (N_19506,N_14993,N_12591);
xor U19507 (N_19507,N_14886,N_12298);
and U19508 (N_19508,N_11654,N_14308);
xor U19509 (N_19509,N_13425,N_10252);
nand U19510 (N_19510,N_13951,N_12006);
and U19511 (N_19511,N_10950,N_10699);
xor U19512 (N_19512,N_10323,N_13523);
nand U19513 (N_19513,N_11612,N_13613);
and U19514 (N_19514,N_11314,N_14347);
nor U19515 (N_19515,N_13337,N_13879);
or U19516 (N_19516,N_11486,N_13288);
and U19517 (N_19517,N_12212,N_13720);
nor U19518 (N_19518,N_12439,N_12545);
nand U19519 (N_19519,N_13039,N_12882);
nor U19520 (N_19520,N_12655,N_13763);
nand U19521 (N_19521,N_12812,N_10806);
xnor U19522 (N_19522,N_13263,N_11234);
and U19523 (N_19523,N_13779,N_13806);
nor U19524 (N_19524,N_10733,N_14692);
and U19525 (N_19525,N_10967,N_13828);
nand U19526 (N_19526,N_14455,N_14217);
xnor U19527 (N_19527,N_13382,N_12748);
nand U19528 (N_19528,N_11173,N_12022);
or U19529 (N_19529,N_13842,N_12060);
and U19530 (N_19530,N_14104,N_12231);
or U19531 (N_19531,N_11915,N_11427);
nor U19532 (N_19532,N_12027,N_11969);
nand U19533 (N_19533,N_11536,N_11408);
nand U19534 (N_19534,N_14342,N_13219);
xor U19535 (N_19535,N_13969,N_11313);
or U19536 (N_19536,N_12494,N_12697);
nand U19537 (N_19537,N_13898,N_11095);
or U19538 (N_19538,N_13740,N_14777);
nand U19539 (N_19539,N_14137,N_12643);
xor U19540 (N_19540,N_10885,N_13359);
nor U19541 (N_19541,N_12650,N_10432);
xor U19542 (N_19542,N_13165,N_12228);
and U19543 (N_19543,N_10971,N_12432);
and U19544 (N_19544,N_12183,N_10711);
and U19545 (N_19545,N_13330,N_13270);
nor U19546 (N_19546,N_12401,N_11478);
or U19547 (N_19547,N_14271,N_10115);
xnor U19548 (N_19548,N_12164,N_13666);
xnor U19549 (N_19549,N_13769,N_11371);
nand U19550 (N_19550,N_14612,N_10690);
nand U19551 (N_19551,N_14611,N_12196);
nand U19552 (N_19552,N_12024,N_11050);
nor U19553 (N_19553,N_10088,N_11509);
nand U19554 (N_19554,N_11986,N_10765);
nand U19555 (N_19555,N_13538,N_12685);
nand U19556 (N_19556,N_13543,N_11437);
nand U19557 (N_19557,N_13749,N_10728);
and U19558 (N_19558,N_13173,N_13269);
nor U19559 (N_19559,N_10135,N_14121);
or U19560 (N_19560,N_14444,N_10759);
xnor U19561 (N_19561,N_13322,N_11343);
nand U19562 (N_19562,N_14231,N_13121);
and U19563 (N_19563,N_12987,N_10100);
or U19564 (N_19564,N_12415,N_13003);
or U19565 (N_19565,N_12112,N_14415);
nand U19566 (N_19566,N_10976,N_13045);
nand U19567 (N_19567,N_10634,N_10221);
and U19568 (N_19568,N_10377,N_14045);
nor U19569 (N_19569,N_14645,N_10183);
and U19570 (N_19570,N_12213,N_12445);
xor U19571 (N_19571,N_11363,N_14873);
or U19572 (N_19572,N_11377,N_14666);
and U19573 (N_19573,N_12865,N_14289);
or U19574 (N_19574,N_12780,N_11181);
nor U19575 (N_19575,N_12033,N_10695);
and U19576 (N_19576,N_14960,N_12254);
nor U19577 (N_19577,N_10054,N_11811);
xnor U19578 (N_19578,N_11707,N_14391);
or U19579 (N_19579,N_13616,N_11973);
and U19580 (N_19580,N_11511,N_12258);
nor U19581 (N_19581,N_12421,N_14049);
or U19582 (N_19582,N_13408,N_14682);
xor U19583 (N_19583,N_10446,N_12674);
nand U19584 (N_19584,N_13360,N_12528);
nor U19585 (N_19585,N_10561,N_14482);
nand U19586 (N_19586,N_10090,N_11153);
nand U19587 (N_19587,N_12094,N_10229);
nand U19588 (N_19588,N_14032,N_14204);
xnor U19589 (N_19589,N_14872,N_12600);
or U19590 (N_19590,N_10039,N_14739);
nor U19591 (N_19591,N_12292,N_13534);
nand U19592 (N_19592,N_14143,N_12969);
xnor U19593 (N_19593,N_12805,N_12467);
nand U19594 (N_19594,N_13157,N_14546);
xnor U19595 (N_19595,N_12558,N_12170);
nand U19596 (N_19596,N_12356,N_10706);
and U19597 (N_19597,N_14428,N_11194);
nand U19598 (N_19598,N_14085,N_10515);
xnor U19599 (N_19599,N_14005,N_14632);
nor U19600 (N_19600,N_14108,N_14701);
xor U19601 (N_19601,N_13158,N_11273);
or U19602 (N_19602,N_10339,N_11781);
nor U19603 (N_19603,N_12446,N_12821);
and U19604 (N_19604,N_10485,N_14210);
or U19605 (N_19605,N_13025,N_14189);
and U19606 (N_19606,N_14205,N_14880);
and U19607 (N_19607,N_10457,N_12836);
or U19608 (N_19608,N_13317,N_10882);
or U19609 (N_19609,N_11829,N_14789);
and U19610 (N_19610,N_10827,N_10463);
xor U19611 (N_19611,N_12202,N_13375);
xnor U19612 (N_19612,N_10550,N_10488);
or U19613 (N_19613,N_11226,N_12228);
nand U19614 (N_19614,N_14207,N_11285);
and U19615 (N_19615,N_13356,N_13812);
xnor U19616 (N_19616,N_11097,N_12482);
and U19617 (N_19617,N_12139,N_14781);
nand U19618 (N_19618,N_10172,N_13629);
or U19619 (N_19619,N_14414,N_12904);
and U19620 (N_19620,N_10831,N_12443);
xor U19621 (N_19621,N_14863,N_10631);
xor U19622 (N_19622,N_11468,N_14414);
nor U19623 (N_19623,N_11698,N_13224);
nor U19624 (N_19624,N_13786,N_14691);
or U19625 (N_19625,N_14071,N_10689);
nand U19626 (N_19626,N_14829,N_10644);
and U19627 (N_19627,N_11190,N_11029);
xor U19628 (N_19628,N_11197,N_12143);
or U19629 (N_19629,N_13503,N_14402);
nand U19630 (N_19630,N_11886,N_11068);
and U19631 (N_19631,N_12265,N_11323);
or U19632 (N_19632,N_13510,N_11834);
nor U19633 (N_19633,N_13162,N_10130);
nor U19634 (N_19634,N_13769,N_12493);
and U19635 (N_19635,N_12244,N_13879);
nor U19636 (N_19636,N_10313,N_10477);
nor U19637 (N_19637,N_13281,N_10204);
nor U19638 (N_19638,N_14295,N_10049);
xor U19639 (N_19639,N_11912,N_11421);
xor U19640 (N_19640,N_11339,N_11701);
and U19641 (N_19641,N_13318,N_10768);
nor U19642 (N_19642,N_13704,N_14894);
nor U19643 (N_19643,N_14056,N_10175);
and U19644 (N_19644,N_13910,N_10771);
and U19645 (N_19645,N_12461,N_12512);
nor U19646 (N_19646,N_13365,N_13852);
nor U19647 (N_19647,N_11522,N_11739);
xnor U19648 (N_19648,N_14910,N_11378);
or U19649 (N_19649,N_12902,N_10152);
and U19650 (N_19650,N_13546,N_14379);
or U19651 (N_19651,N_14398,N_12056);
nor U19652 (N_19652,N_11926,N_11686);
nand U19653 (N_19653,N_10998,N_11822);
or U19654 (N_19654,N_13011,N_12344);
xor U19655 (N_19655,N_13211,N_14000);
nor U19656 (N_19656,N_11659,N_12316);
nand U19657 (N_19657,N_13107,N_14812);
xnor U19658 (N_19658,N_11801,N_14223);
xor U19659 (N_19659,N_14821,N_13403);
or U19660 (N_19660,N_12443,N_14770);
xnor U19661 (N_19661,N_13879,N_13134);
nor U19662 (N_19662,N_13946,N_11307);
nor U19663 (N_19663,N_11127,N_13590);
or U19664 (N_19664,N_12986,N_11775);
xor U19665 (N_19665,N_10972,N_13523);
nor U19666 (N_19666,N_13442,N_14406);
xnor U19667 (N_19667,N_14544,N_10450);
xor U19668 (N_19668,N_10394,N_12694);
nand U19669 (N_19669,N_13044,N_11820);
and U19670 (N_19670,N_12970,N_14941);
or U19671 (N_19671,N_14438,N_14453);
or U19672 (N_19672,N_14493,N_14712);
and U19673 (N_19673,N_13400,N_14188);
and U19674 (N_19674,N_12715,N_11312);
nor U19675 (N_19675,N_14203,N_11679);
nand U19676 (N_19676,N_14999,N_12984);
xnor U19677 (N_19677,N_14820,N_11143);
or U19678 (N_19678,N_13258,N_11533);
and U19679 (N_19679,N_10381,N_12714);
or U19680 (N_19680,N_11079,N_14061);
nor U19681 (N_19681,N_14319,N_10343);
xor U19682 (N_19682,N_12197,N_14974);
and U19683 (N_19683,N_13722,N_14501);
nand U19684 (N_19684,N_13889,N_11218);
nand U19685 (N_19685,N_10327,N_14899);
xnor U19686 (N_19686,N_11274,N_11717);
or U19687 (N_19687,N_11909,N_13303);
nand U19688 (N_19688,N_12612,N_10238);
nand U19689 (N_19689,N_12789,N_14304);
and U19690 (N_19690,N_11864,N_10531);
xor U19691 (N_19691,N_13165,N_14744);
xnor U19692 (N_19692,N_12673,N_13223);
and U19693 (N_19693,N_11026,N_12906);
xnor U19694 (N_19694,N_11827,N_11468);
nand U19695 (N_19695,N_12922,N_10414);
nand U19696 (N_19696,N_13369,N_14625);
nand U19697 (N_19697,N_11349,N_14010);
xor U19698 (N_19698,N_10330,N_12490);
nand U19699 (N_19699,N_13872,N_12721);
xnor U19700 (N_19700,N_11846,N_11557);
or U19701 (N_19701,N_12262,N_10159);
nand U19702 (N_19702,N_14171,N_12788);
or U19703 (N_19703,N_10760,N_11814);
xor U19704 (N_19704,N_12695,N_14636);
and U19705 (N_19705,N_10784,N_11160);
and U19706 (N_19706,N_11755,N_13600);
and U19707 (N_19707,N_13300,N_14805);
nor U19708 (N_19708,N_12181,N_14471);
or U19709 (N_19709,N_12955,N_11815);
xor U19710 (N_19710,N_14100,N_14851);
nand U19711 (N_19711,N_13599,N_10315);
nand U19712 (N_19712,N_12503,N_14270);
nor U19713 (N_19713,N_13925,N_10192);
or U19714 (N_19714,N_14086,N_11613);
xnor U19715 (N_19715,N_11186,N_14551);
nor U19716 (N_19716,N_11716,N_12097);
nor U19717 (N_19717,N_10954,N_10322);
nand U19718 (N_19718,N_13049,N_12403);
and U19719 (N_19719,N_13043,N_13511);
nand U19720 (N_19720,N_14506,N_11919);
xnor U19721 (N_19721,N_13525,N_12659);
and U19722 (N_19722,N_11968,N_14734);
and U19723 (N_19723,N_14403,N_11885);
xor U19724 (N_19724,N_14712,N_13087);
xnor U19725 (N_19725,N_14764,N_12212);
nor U19726 (N_19726,N_13227,N_14386);
or U19727 (N_19727,N_14861,N_12197);
nor U19728 (N_19728,N_13247,N_14874);
or U19729 (N_19729,N_12700,N_12669);
or U19730 (N_19730,N_10852,N_13270);
or U19731 (N_19731,N_14356,N_14661);
xnor U19732 (N_19732,N_12468,N_14320);
and U19733 (N_19733,N_10723,N_11063);
nor U19734 (N_19734,N_10335,N_10809);
nor U19735 (N_19735,N_11795,N_13608);
or U19736 (N_19736,N_12725,N_12179);
and U19737 (N_19737,N_10834,N_14983);
or U19738 (N_19738,N_13497,N_10535);
nor U19739 (N_19739,N_12202,N_11434);
xor U19740 (N_19740,N_13217,N_12114);
xnor U19741 (N_19741,N_10249,N_11911);
nand U19742 (N_19742,N_10985,N_13578);
and U19743 (N_19743,N_12659,N_13969);
nand U19744 (N_19744,N_14496,N_13545);
xnor U19745 (N_19745,N_14498,N_12296);
nand U19746 (N_19746,N_14103,N_11148);
nand U19747 (N_19747,N_10041,N_13780);
nor U19748 (N_19748,N_12899,N_10588);
xnor U19749 (N_19749,N_14212,N_12523);
and U19750 (N_19750,N_14949,N_14140);
nor U19751 (N_19751,N_13478,N_11366);
xnor U19752 (N_19752,N_11355,N_12314);
xnor U19753 (N_19753,N_14502,N_14020);
or U19754 (N_19754,N_12484,N_11215);
and U19755 (N_19755,N_12988,N_12127);
nor U19756 (N_19756,N_11992,N_12971);
xnor U19757 (N_19757,N_14105,N_14349);
or U19758 (N_19758,N_12321,N_11120);
and U19759 (N_19759,N_12035,N_14655);
and U19760 (N_19760,N_10982,N_10943);
nand U19761 (N_19761,N_10633,N_13366);
nor U19762 (N_19762,N_11022,N_14537);
and U19763 (N_19763,N_14770,N_14548);
nand U19764 (N_19764,N_10707,N_14646);
and U19765 (N_19765,N_12222,N_14877);
nand U19766 (N_19766,N_11179,N_14370);
nor U19767 (N_19767,N_11312,N_11474);
nor U19768 (N_19768,N_14310,N_13398);
nand U19769 (N_19769,N_14962,N_13209);
nor U19770 (N_19770,N_13919,N_11865);
xnor U19771 (N_19771,N_10971,N_10374);
and U19772 (N_19772,N_10649,N_11571);
and U19773 (N_19773,N_12299,N_11534);
xor U19774 (N_19774,N_14090,N_12749);
xor U19775 (N_19775,N_13498,N_13878);
and U19776 (N_19776,N_11999,N_10450);
nand U19777 (N_19777,N_14031,N_12726);
and U19778 (N_19778,N_10980,N_13998);
or U19779 (N_19779,N_12281,N_11852);
nand U19780 (N_19780,N_10789,N_13207);
or U19781 (N_19781,N_12549,N_14978);
nor U19782 (N_19782,N_11703,N_12977);
nand U19783 (N_19783,N_13923,N_14726);
nor U19784 (N_19784,N_13981,N_12663);
xnor U19785 (N_19785,N_13757,N_11696);
or U19786 (N_19786,N_12026,N_10028);
nor U19787 (N_19787,N_14651,N_14729);
xor U19788 (N_19788,N_12761,N_11308);
or U19789 (N_19789,N_11286,N_14233);
or U19790 (N_19790,N_10835,N_14947);
nor U19791 (N_19791,N_12177,N_11167);
or U19792 (N_19792,N_12057,N_13150);
xor U19793 (N_19793,N_10070,N_12192);
or U19794 (N_19794,N_11582,N_10817);
and U19795 (N_19795,N_10079,N_10662);
xnor U19796 (N_19796,N_14458,N_12584);
or U19797 (N_19797,N_14956,N_13500);
nor U19798 (N_19798,N_13180,N_12488);
xor U19799 (N_19799,N_13025,N_13290);
nor U19800 (N_19800,N_11335,N_13037);
and U19801 (N_19801,N_12593,N_14738);
and U19802 (N_19802,N_14563,N_13899);
or U19803 (N_19803,N_11802,N_11429);
and U19804 (N_19804,N_14313,N_12849);
nand U19805 (N_19805,N_11170,N_10063);
or U19806 (N_19806,N_14617,N_10395);
xor U19807 (N_19807,N_12607,N_12835);
xnor U19808 (N_19808,N_13920,N_12390);
nor U19809 (N_19809,N_10470,N_12280);
nand U19810 (N_19810,N_14659,N_12708);
and U19811 (N_19811,N_12243,N_13876);
nand U19812 (N_19812,N_13086,N_11599);
nand U19813 (N_19813,N_14899,N_12587);
or U19814 (N_19814,N_13095,N_12514);
xnor U19815 (N_19815,N_13838,N_10617);
and U19816 (N_19816,N_14728,N_13451);
and U19817 (N_19817,N_11406,N_11929);
nand U19818 (N_19818,N_10583,N_14691);
xnor U19819 (N_19819,N_12529,N_11625);
and U19820 (N_19820,N_10034,N_11821);
nand U19821 (N_19821,N_13446,N_14036);
nor U19822 (N_19822,N_12577,N_14473);
or U19823 (N_19823,N_10556,N_11768);
nand U19824 (N_19824,N_12433,N_12424);
or U19825 (N_19825,N_11200,N_11904);
nand U19826 (N_19826,N_11108,N_13307);
or U19827 (N_19827,N_12744,N_11999);
nand U19828 (N_19828,N_14863,N_11275);
or U19829 (N_19829,N_13829,N_11101);
and U19830 (N_19830,N_13379,N_13344);
nand U19831 (N_19831,N_10592,N_12435);
nand U19832 (N_19832,N_14128,N_13955);
nor U19833 (N_19833,N_11979,N_11976);
nor U19834 (N_19834,N_12071,N_13580);
nor U19835 (N_19835,N_14847,N_14515);
xor U19836 (N_19836,N_10079,N_10327);
nor U19837 (N_19837,N_11562,N_12115);
nand U19838 (N_19838,N_10563,N_13093);
or U19839 (N_19839,N_10030,N_12094);
or U19840 (N_19840,N_12025,N_14035);
or U19841 (N_19841,N_11313,N_11654);
or U19842 (N_19842,N_13011,N_10027);
nor U19843 (N_19843,N_14546,N_12252);
nand U19844 (N_19844,N_11926,N_12554);
nor U19845 (N_19845,N_10895,N_13859);
nand U19846 (N_19846,N_11587,N_11443);
nor U19847 (N_19847,N_14992,N_11419);
or U19848 (N_19848,N_14522,N_11791);
or U19849 (N_19849,N_12931,N_11576);
xor U19850 (N_19850,N_10807,N_13810);
nand U19851 (N_19851,N_13931,N_14955);
xor U19852 (N_19852,N_11531,N_10776);
nor U19853 (N_19853,N_14546,N_10197);
nand U19854 (N_19854,N_13021,N_13941);
xor U19855 (N_19855,N_13990,N_11549);
nand U19856 (N_19856,N_10848,N_12794);
xnor U19857 (N_19857,N_10368,N_14641);
xnor U19858 (N_19858,N_12927,N_11195);
or U19859 (N_19859,N_14458,N_14516);
nor U19860 (N_19860,N_12373,N_11139);
xor U19861 (N_19861,N_14572,N_13134);
xor U19862 (N_19862,N_10565,N_11096);
nor U19863 (N_19863,N_10797,N_12147);
nand U19864 (N_19864,N_10486,N_14247);
or U19865 (N_19865,N_10403,N_11037);
and U19866 (N_19866,N_11857,N_11538);
or U19867 (N_19867,N_13792,N_10818);
nor U19868 (N_19868,N_12869,N_13963);
and U19869 (N_19869,N_13709,N_10761);
and U19870 (N_19870,N_10397,N_10432);
and U19871 (N_19871,N_14859,N_10118);
or U19872 (N_19872,N_10543,N_14529);
nand U19873 (N_19873,N_10277,N_12359);
xor U19874 (N_19874,N_14487,N_13259);
nor U19875 (N_19875,N_12084,N_12179);
or U19876 (N_19876,N_14304,N_12377);
nor U19877 (N_19877,N_10855,N_11208);
nand U19878 (N_19878,N_11643,N_11287);
xor U19879 (N_19879,N_11301,N_12098);
nand U19880 (N_19880,N_14036,N_12507);
nand U19881 (N_19881,N_13957,N_12218);
xnor U19882 (N_19882,N_12619,N_11582);
xor U19883 (N_19883,N_12054,N_13508);
nor U19884 (N_19884,N_12208,N_14975);
or U19885 (N_19885,N_12814,N_14928);
or U19886 (N_19886,N_10687,N_12344);
nand U19887 (N_19887,N_10208,N_13453);
nand U19888 (N_19888,N_10614,N_11447);
nor U19889 (N_19889,N_11931,N_14828);
xnor U19890 (N_19890,N_11559,N_11248);
and U19891 (N_19891,N_12696,N_11545);
nor U19892 (N_19892,N_11012,N_11267);
and U19893 (N_19893,N_14155,N_13157);
or U19894 (N_19894,N_10457,N_14657);
nand U19895 (N_19895,N_14930,N_10093);
xnor U19896 (N_19896,N_10476,N_12968);
and U19897 (N_19897,N_13395,N_13833);
nand U19898 (N_19898,N_11772,N_11025);
nor U19899 (N_19899,N_12011,N_13006);
or U19900 (N_19900,N_11632,N_11343);
and U19901 (N_19901,N_13940,N_12737);
xnor U19902 (N_19902,N_13244,N_10597);
nor U19903 (N_19903,N_10423,N_14106);
nor U19904 (N_19904,N_11618,N_11009);
xor U19905 (N_19905,N_10362,N_13532);
xnor U19906 (N_19906,N_14404,N_13623);
xnor U19907 (N_19907,N_13698,N_14844);
nand U19908 (N_19908,N_11424,N_11311);
or U19909 (N_19909,N_14483,N_11055);
nor U19910 (N_19910,N_14401,N_13009);
and U19911 (N_19911,N_11764,N_14452);
and U19912 (N_19912,N_14201,N_12092);
nand U19913 (N_19913,N_14266,N_10124);
nand U19914 (N_19914,N_12849,N_10901);
or U19915 (N_19915,N_14967,N_11540);
nand U19916 (N_19916,N_13092,N_10618);
nor U19917 (N_19917,N_12957,N_14663);
xnor U19918 (N_19918,N_13219,N_12189);
and U19919 (N_19919,N_12986,N_10263);
or U19920 (N_19920,N_12836,N_11656);
nand U19921 (N_19921,N_12341,N_14110);
or U19922 (N_19922,N_10781,N_13955);
xnor U19923 (N_19923,N_14249,N_14161);
nand U19924 (N_19924,N_10513,N_14927);
nand U19925 (N_19925,N_13564,N_10773);
or U19926 (N_19926,N_10793,N_14144);
xor U19927 (N_19927,N_12981,N_11893);
nor U19928 (N_19928,N_10323,N_11784);
nor U19929 (N_19929,N_11462,N_10944);
and U19930 (N_19930,N_10630,N_13148);
and U19931 (N_19931,N_12179,N_13721);
nand U19932 (N_19932,N_14891,N_13151);
nand U19933 (N_19933,N_13834,N_14928);
xor U19934 (N_19934,N_11612,N_11138);
and U19935 (N_19935,N_12781,N_13137);
or U19936 (N_19936,N_10671,N_14669);
xnor U19937 (N_19937,N_14928,N_13587);
nand U19938 (N_19938,N_12285,N_14278);
or U19939 (N_19939,N_12513,N_10980);
xnor U19940 (N_19940,N_14188,N_10139);
xor U19941 (N_19941,N_10939,N_10182);
xor U19942 (N_19942,N_10683,N_13714);
xor U19943 (N_19943,N_10919,N_13026);
nor U19944 (N_19944,N_13393,N_13139);
or U19945 (N_19945,N_14182,N_13697);
xnor U19946 (N_19946,N_13959,N_11289);
or U19947 (N_19947,N_11818,N_14953);
and U19948 (N_19948,N_10903,N_13161);
xor U19949 (N_19949,N_11187,N_12672);
or U19950 (N_19950,N_10204,N_14840);
xnor U19951 (N_19951,N_14484,N_12244);
and U19952 (N_19952,N_12897,N_12762);
nand U19953 (N_19953,N_12121,N_12371);
nand U19954 (N_19954,N_14652,N_13398);
nand U19955 (N_19955,N_10776,N_10444);
nand U19956 (N_19956,N_10596,N_12902);
or U19957 (N_19957,N_12991,N_12074);
or U19958 (N_19958,N_12010,N_11651);
nand U19959 (N_19959,N_11104,N_14565);
and U19960 (N_19960,N_13446,N_10704);
or U19961 (N_19961,N_12495,N_13773);
or U19962 (N_19962,N_12965,N_14557);
nand U19963 (N_19963,N_11049,N_11159);
nor U19964 (N_19964,N_12769,N_10582);
and U19965 (N_19965,N_12726,N_14590);
or U19966 (N_19966,N_11752,N_11207);
nand U19967 (N_19967,N_12757,N_11040);
nor U19968 (N_19968,N_13618,N_13718);
or U19969 (N_19969,N_11706,N_14245);
and U19970 (N_19970,N_10725,N_13715);
xnor U19971 (N_19971,N_11052,N_13568);
xnor U19972 (N_19972,N_12557,N_11187);
nand U19973 (N_19973,N_11272,N_13199);
nand U19974 (N_19974,N_11158,N_14746);
nand U19975 (N_19975,N_14252,N_11102);
and U19976 (N_19976,N_14132,N_11826);
nor U19977 (N_19977,N_12933,N_10354);
nand U19978 (N_19978,N_14738,N_11913);
or U19979 (N_19979,N_13664,N_10330);
nand U19980 (N_19980,N_12895,N_14308);
xor U19981 (N_19981,N_14078,N_12312);
and U19982 (N_19982,N_11808,N_13792);
and U19983 (N_19983,N_12878,N_10975);
nand U19984 (N_19984,N_13084,N_14313);
or U19985 (N_19985,N_11278,N_13990);
or U19986 (N_19986,N_12074,N_14690);
and U19987 (N_19987,N_10775,N_10581);
or U19988 (N_19988,N_13842,N_10983);
nand U19989 (N_19989,N_13347,N_13894);
nor U19990 (N_19990,N_11161,N_14189);
or U19991 (N_19991,N_11798,N_14023);
nand U19992 (N_19992,N_12864,N_12052);
nor U19993 (N_19993,N_14525,N_10174);
nor U19994 (N_19994,N_12752,N_13378);
and U19995 (N_19995,N_13760,N_11378);
nor U19996 (N_19996,N_14433,N_13169);
or U19997 (N_19997,N_13459,N_13677);
nor U19998 (N_19998,N_13596,N_10217);
nor U19999 (N_19999,N_14760,N_14986);
nand UO_0 (O_0,N_16944,N_15999);
and UO_1 (O_1,N_17649,N_17383);
xnor UO_2 (O_2,N_19946,N_18070);
or UO_3 (O_3,N_16796,N_19057);
nand UO_4 (O_4,N_18064,N_17174);
or UO_5 (O_5,N_16902,N_15607);
or UO_6 (O_6,N_19265,N_15772);
nand UO_7 (O_7,N_16424,N_18924);
nand UO_8 (O_8,N_17090,N_16004);
and UO_9 (O_9,N_18975,N_16867);
and UO_10 (O_10,N_17559,N_16248);
nor UO_11 (O_11,N_16865,N_15466);
nor UO_12 (O_12,N_17165,N_18711);
xnor UO_13 (O_13,N_15762,N_16486);
xor UO_14 (O_14,N_18909,N_16606);
nand UO_15 (O_15,N_15023,N_15227);
nor UO_16 (O_16,N_15906,N_16889);
and UO_17 (O_17,N_15964,N_16336);
nand UO_18 (O_18,N_15660,N_18578);
or UO_19 (O_19,N_17733,N_17319);
nor UO_20 (O_20,N_17023,N_16392);
or UO_21 (O_21,N_15550,N_19628);
nand UO_22 (O_22,N_17399,N_17230);
or UO_23 (O_23,N_16899,N_17601);
nor UO_24 (O_24,N_17200,N_16370);
or UO_25 (O_25,N_18891,N_15666);
or UO_26 (O_26,N_15232,N_19240);
or UO_27 (O_27,N_17953,N_18503);
nor UO_28 (O_28,N_18979,N_18886);
or UO_29 (O_29,N_18019,N_16096);
nor UO_30 (O_30,N_19899,N_19267);
xor UO_31 (O_31,N_19724,N_16909);
xor UO_32 (O_32,N_19187,N_17515);
and UO_33 (O_33,N_15858,N_16303);
nor UO_34 (O_34,N_18466,N_16629);
nor UO_35 (O_35,N_16518,N_15729);
xnor UO_36 (O_36,N_16761,N_19823);
nor UO_37 (O_37,N_17665,N_16066);
or UO_38 (O_38,N_18295,N_16536);
or UO_39 (O_39,N_19526,N_17007);
nand UO_40 (O_40,N_19186,N_17751);
nand UO_41 (O_41,N_15676,N_17414);
nand UO_42 (O_42,N_19742,N_16449);
or UO_43 (O_43,N_16516,N_19533);
xnor UO_44 (O_44,N_15400,N_17377);
nand UO_45 (O_45,N_17458,N_19014);
and UO_46 (O_46,N_16210,N_16841);
and UO_47 (O_47,N_17641,N_17854);
xnor UO_48 (O_48,N_15256,N_18446);
and UO_49 (O_49,N_17940,N_17056);
or UO_50 (O_50,N_18003,N_18903);
xor UO_51 (O_51,N_16553,N_19335);
nand UO_52 (O_52,N_16159,N_15047);
nand UO_53 (O_53,N_18098,N_15138);
xor UO_54 (O_54,N_16979,N_16595);
and UO_55 (O_55,N_16640,N_15013);
or UO_56 (O_56,N_19867,N_17771);
xor UO_57 (O_57,N_17283,N_17690);
and UO_58 (O_58,N_15016,N_18919);
nor UO_59 (O_59,N_16737,N_16344);
and UO_60 (O_60,N_18196,N_17606);
nor UO_61 (O_61,N_19914,N_15057);
nor UO_62 (O_62,N_16877,N_15587);
nand UO_63 (O_63,N_19484,N_19405);
nand UO_64 (O_64,N_19120,N_19391);
and UO_65 (O_65,N_16133,N_18881);
xor UO_66 (O_66,N_16713,N_18202);
xor UO_67 (O_67,N_17125,N_15565);
or UO_68 (O_68,N_18255,N_15625);
nor UO_69 (O_69,N_19771,N_15902);
and UO_70 (O_70,N_19140,N_17578);
nand UO_71 (O_71,N_15284,N_19833);
or UO_72 (O_72,N_17322,N_17583);
xnor UO_73 (O_73,N_17931,N_16590);
nand UO_74 (O_74,N_17916,N_19220);
or UO_75 (O_75,N_19446,N_17813);
or UO_76 (O_76,N_17190,N_16472);
or UO_77 (O_77,N_18766,N_15879);
nand UO_78 (O_78,N_19569,N_18786);
nor UO_79 (O_79,N_17505,N_16884);
or UO_80 (O_80,N_15490,N_16932);
xor UO_81 (O_81,N_18483,N_17946);
xnor UO_82 (O_82,N_17514,N_18710);
nand UO_83 (O_83,N_16772,N_19314);
nor UO_84 (O_84,N_15793,N_18474);
and UO_85 (O_85,N_15020,N_19884);
nor UO_86 (O_86,N_19115,N_16119);
xnor UO_87 (O_87,N_16235,N_15350);
or UO_88 (O_88,N_19069,N_18228);
xnor UO_89 (O_89,N_18203,N_19308);
nand UO_90 (O_90,N_19002,N_19476);
xor UO_91 (O_91,N_17517,N_15730);
nand UO_92 (O_92,N_15201,N_17543);
xor UO_93 (O_93,N_18637,N_18490);
nand UO_94 (O_94,N_15408,N_19514);
nor UO_95 (O_95,N_17356,N_18308);
nor UO_96 (O_96,N_15344,N_15129);
and UO_97 (O_97,N_16810,N_16948);
or UO_98 (O_98,N_18966,N_19895);
or UO_99 (O_99,N_17851,N_18081);
nor UO_100 (O_100,N_19355,N_17353);
nand UO_101 (O_101,N_18819,N_15100);
and UO_102 (O_102,N_18524,N_19725);
nor UO_103 (O_103,N_18007,N_19189);
or UO_104 (O_104,N_16842,N_18166);
xnor UO_105 (O_105,N_17636,N_16854);
nor UO_106 (O_106,N_18132,N_19126);
nor UO_107 (O_107,N_19481,N_19862);
or UO_108 (O_108,N_18762,N_16749);
and UO_109 (O_109,N_15656,N_16880);
and UO_110 (O_110,N_19516,N_15334);
xor UO_111 (O_111,N_18247,N_15875);
nor UO_112 (O_112,N_17484,N_18596);
xnor UO_113 (O_113,N_18194,N_17588);
nor UO_114 (O_114,N_16738,N_19709);
or UO_115 (O_115,N_16950,N_15121);
xor UO_116 (O_116,N_19550,N_18883);
xor UO_117 (O_117,N_18626,N_16381);
xor UO_118 (O_118,N_18587,N_19045);
nand UO_119 (O_119,N_16489,N_18276);
nor UO_120 (O_120,N_17693,N_18516);
nand UO_121 (O_121,N_17951,N_18195);
xor UO_122 (O_122,N_17538,N_19434);
nand UO_123 (O_123,N_15886,N_19989);
xnor UO_124 (O_124,N_15120,N_18404);
nor UO_125 (O_125,N_15795,N_16929);
nand UO_126 (O_126,N_18436,N_19772);
or UO_127 (O_127,N_16132,N_15953);
or UO_128 (O_128,N_15220,N_15473);
nand UO_129 (O_129,N_19842,N_16218);
xor UO_130 (O_130,N_15367,N_16304);
nor UO_131 (O_131,N_18902,N_19567);
nor UO_132 (O_132,N_19806,N_15544);
and UO_133 (O_133,N_19848,N_17914);
xor UO_134 (O_134,N_16460,N_18629);
nor UO_135 (O_135,N_16388,N_17460);
and UO_136 (O_136,N_15911,N_16898);
or UO_137 (O_137,N_18890,N_19111);
nand UO_138 (O_138,N_19036,N_15123);
or UO_139 (O_139,N_18409,N_17391);
nand UO_140 (O_140,N_15713,N_18319);
or UO_141 (O_141,N_18406,N_19900);
or UO_142 (O_142,N_19441,N_17386);
nor UO_143 (O_143,N_16627,N_18821);
nor UO_144 (O_144,N_17078,N_18770);
nor UO_145 (O_145,N_18817,N_17720);
nand UO_146 (O_146,N_18021,N_18478);
and UO_147 (O_147,N_17626,N_18367);
nand UO_148 (O_148,N_16168,N_16419);
or UO_149 (O_149,N_17985,N_18192);
nand UO_150 (O_150,N_19046,N_15492);
and UO_151 (O_151,N_17909,N_18048);
nand UO_152 (O_152,N_17066,N_19143);
nor UO_153 (O_153,N_19557,N_16915);
or UO_154 (O_154,N_17186,N_19455);
or UO_155 (O_155,N_17969,N_16679);
or UO_156 (O_156,N_15766,N_17518);
or UO_157 (O_157,N_16125,N_17416);
nor UO_158 (O_158,N_16745,N_17836);
nor UO_159 (O_159,N_18805,N_18914);
xnor UO_160 (O_160,N_17135,N_16414);
or UO_161 (O_161,N_17777,N_18469);
or UO_162 (O_162,N_17536,N_16395);
nand UO_163 (O_163,N_18664,N_17662);
nand UO_164 (O_164,N_15166,N_15005);
xor UO_165 (O_165,N_15074,N_17509);
or UO_166 (O_166,N_17139,N_19438);
nor UO_167 (O_167,N_19788,N_19775);
nand UO_168 (O_168,N_16289,N_16998);
xor UO_169 (O_169,N_16971,N_18097);
or UO_170 (O_170,N_19356,N_15157);
or UO_171 (O_171,N_19810,N_15050);
nor UO_172 (O_172,N_17858,N_16873);
or UO_173 (O_173,N_15931,N_16314);
and UO_174 (O_174,N_18125,N_17779);
nor UO_175 (O_175,N_16162,N_16150);
xor UO_176 (O_176,N_16102,N_15663);
xnor UO_177 (O_177,N_19590,N_19875);
and UO_178 (O_178,N_18075,N_16957);
nand UO_179 (O_179,N_16740,N_15867);
and UO_180 (O_180,N_16729,N_15131);
or UO_181 (O_181,N_15611,N_17154);
xor UO_182 (O_182,N_18504,N_17264);
or UO_183 (O_183,N_16712,N_17256);
and UO_184 (O_184,N_15692,N_15465);
nor UO_185 (O_185,N_19419,N_17823);
and UO_186 (O_186,N_15298,N_19483);
nor UO_187 (O_187,N_15234,N_15533);
and UO_188 (O_188,N_19085,N_19197);
nor UO_189 (O_189,N_19161,N_19676);
and UO_190 (O_190,N_19912,N_16819);
xor UO_191 (O_191,N_15240,N_17705);
nand UO_192 (O_192,N_15045,N_16940);
xnor UO_193 (O_193,N_15064,N_15345);
xor UO_194 (O_194,N_17421,N_19926);
and UO_195 (O_195,N_15303,N_18254);
nand UO_196 (O_196,N_15147,N_15900);
nor UO_197 (O_197,N_18912,N_16912);
or UO_198 (O_198,N_17191,N_17840);
and UO_199 (O_199,N_17932,N_17899);
nor UO_200 (O_200,N_19089,N_18784);
xor UO_201 (O_201,N_17491,N_19889);
xor UO_202 (O_202,N_19565,N_19431);
nor UO_203 (O_203,N_15788,N_19191);
and UO_204 (O_204,N_18213,N_16888);
nand UO_205 (O_205,N_18672,N_15545);
xor UO_206 (O_206,N_18355,N_15778);
xnor UO_207 (O_207,N_15436,N_19216);
xor UO_208 (O_208,N_16617,N_18414);
nand UO_209 (O_209,N_19644,N_16562);
or UO_210 (O_210,N_17954,N_15258);
and UO_211 (O_211,N_19805,N_15073);
nor UO_212 (O_212,N_19773,N_18403);
xor UO_213 (O_213,N_18759,N_17841);
or UO_214 (O_214,N_19188,N_17017);
nand UO_215 (O_215,N_18282,N_16667);
nand UO_216 (O_216,N_18984,N_16665);
nand UO_217 (O_217,N_19378,N_17292);
or UO_218 (O_218,N_18158,N_17281);
nand UO_219 (O_219,N_18811,N_18065);
xor UO_220 (O_220,N_15719,N_17702);
xnor UO_221 (O_221,N_16184,N_17326);
xor UO_222 (O_222,N_19148,N_19545);
nand UO_223 (O_223,N_15280,N_15851);
nand UO_224 (O_224,N_16148,N_16837);
and UO_225 (O_225,N_16934,N_16101);
xor UO_226 (O_226,N_16324,N_15110);
xor UO_227 (O_227,N_19517,N_15049);
xnor UO_228 (O_228,N_19118,N_16636);
and UO_229 (O_229,N_19741,N_16782);
xnor UO_230 (O_230,N_16069,N_16992);
and UO_231 (O_231,N_16196,N_15387);
and UO_232 (O_232,N_16339,N_19876);
nor UO_233 (O_233,N_19341,N_15595);
nor UO_234 (O_234,N_16579,N_17555);
nor UO_235 (O_235,N_18602,N_19655);
nand UO_236 (O_236,N_17815,N_16718);
or UO_237 (O_237,N_17520,N_16759);
xnor UO_238 (O_238,N_16177,N_19090);
and UO_239 (O_239,N_17005,N_15554);
and UO_240 (O_240,N_19698,N_15101);
xnor UO_241 (O_241,N_15153,N_15773);
and UO_242 (O_242,N_17506,N_19262);
and UO_243 (O_243,N_19025,N_15892);
nand UO_244 (O_244,N_17558,N_17318);
nor UO_245 (O_245,N_18391,N_16300);
and UO_246 (O_246,N_17409,N_19092);
xor UO_247 (O_247,N_17730,N_15756);
nor UO_248 (O_248,N_16316,N_17067);
or UO_249 (O_249,N_19368,N_16987);
or UO_250 (O_250,N_17596,N_18031);
or UO_251 (O_251,N_17622,N_16400);
xor UO_252 (O_252,N_15839,N_19803);
or UO_253 (O_253,N_16268,N_15286);
or UO_254 (O_254,N_15021,N_15551);
and UO_255 (O_255,N_16391,N_16361);
or UO_256 (O_256,N_16373,N_16770);
xnor UO_257 (O_257,N_17568,N_18684);
xnor UO_258 (O_258,N_18143,N_18157);
xnor UO_259 (O_259,N_17585,N_18865);
xor UO_260 (O_260,N_15525,N_17146);
nor UO_261 (O_261,N_15965,N_19997);
nand UO_262 (O_262,N_16876,N_19540);
and UO_263 (O_263,N_16193,N_17224);
and UO_264 (O_264,N_19019,N_18178);
xnor UO_265 (O_265,N_18101,N_17285);
nand UO_266 (O_266,N_15685,N_15883);
or UO_267 (O_267,N_19583,N_16242);
xor UO_268 (O_268,N_16448,N_16188);
or UO_269 (O_269,N_18253,N_19711);
nand UO_270 (O_270,N_19326,N_17493);
xnor UO_271 (O_271,N_17642,N_18802);
nand UO_272 (O_272,N_17324,N_19001);
or UO_273 (O_273,N_16806,N_16180);
nor UO_274 (O_274,N_16223,N_19690);
xor UO_275 (O_275,N_19662,N_16163);
and UO_276 (O_276,N_17406,N_15094);
xnor UO_277 (O_277,N_18991,N_17167);
nand UO_278 (O_278,N_15877,N_15861);
nand UO_279 (O_279,N_18614,N_15508);
or UO_280 (O_280,N_15113,N_16386);
and UO_281 (O_281,N_17994,N_16698);
nand UO_282 (O_282,N_15461,N_15152);
and UO_283 (O_283,N_16769,N_16099);
nand UO_284 (O_284,N_15959,N_16885);
and UO_285 (O_285,N_17850,N_19641);
nand UO_286 (O_286,N_15469,N_17692);
and UO_287 (O_287,N_15184,N_19653);
nor UO_288 (O_288,N_15882,N_17437);
nand UO_289 (O_289,N_18686,N_19897);
nor UO_290 (O_290,N_18080,N_17158);
or UO_291 (O_291,N_15535,N_19928);
nand UO_292 (O_292,N_18564,N_18956);
xnor UO_293 (O_293,N_16130,N_18520);
nand UO_294 (O_294,N_18592,N_16609);
and UO_295 (O_295,N_19903,N_17420);
and UO_296 (O_296,N_19617,N_17431);
and UO_297 (O_297,N_17508,N_15828);
nor UO_298 (O_298,N_15962,N_19620);
xnor UO_299 (O_299,N_15249,N_16530);
xor UO_300 (O_300,N_16656,N_16312);
or UO_301 (O_301,N_16702,N_18808);
xor UO_302 (O_302,N_19196,N_15395);
nor UO_303 (O_303,N_19064,N_18868);
nor UO_304 (O_304,N_15104,N_15415);
nor UO_305 (O_305,N_18576,N_18959);
or UO_306 (O_306,N_18094,N_17894);
nand UO_307 (O_307,N_18451,N_18087);
nand UO_308 (O_308,N_17166,N_17624);
xor UO_309 (O_309,N_19223,N_16387);
nand UO_310 (O_310,N_18559,N_15869);
or UO_311 (O_311,N_15680,N_17474);
or UO_312 (O_312,N_17922,N_16097);
nand UO_313 (O_313,N_19295,N_19443);
nand UO_314 (O_314,N_18339,N_16956);
xor UO_315 (O_315,N_19638,N_17463);
nand UO_316 (O_316,N_18565,N_15504);
nor UO_317 (O_317,N_16278,N_15615);
nor UO_318 (O_318,N_19561,N_19871);
nand UO_319 (O_319,N_16155,N_16550);
nor UO_320 (O_320,N_17625,N_18974);
and UO_321 (O_321,N_16081,N_16493);
nor UO_322 (O_322,N_19944,N_16285);
nand UO_323 (O_323,N_17749,N_17072);
or UO_324 (O_324,N_17092,N_15293);
and UO_325 (O_325,N_19865,N_16980);
xnor UO_326 (O_326,N_16653,N_17832);
or UO_327 (O_327,N_16778,N_16129);
nor UO_328 (O_328,N_16820,N_17127);
or UO_329 (O_329,N_15938,N_19408);
and UO_330 (O_330,N_18977,N_17401);
and UO_331 (O_331,N_15035,N_15758);
xor UO_332 (O_332,N_18329,N_16247);
nand UO_333 (O_333,N_18286,N_18941);
nor UO_334 (O_334,N_17239,N_16900);
nor UO_335 (O_335,N_18230,N_15951);
and UO_336 (O_336,N_16657,N_18111);
or UO_337 (O_337,N_15079,N_16996);
xor UO_338 (O_338,N_19398,N_17222);
nor UO_339 (O_339,N_17796,N_18826);
and UO_340 (O_340,N_17184,N_19168);
nor UO_341 (O_341,N_17615,N_17159);
xnor UO_342 (O_342,N_18476,N_18754);
nand UO_343 (O_343,N_15389,N_17883);
nor UO_344 (O_344,N_19736,N_17580);
nand UO_345 (O_345,N_18427,N_16243);
or UO_346 (O_346,N_15827,N_17701);
xnor UO_347 (O_347,N_15777,N_15488);
nor UO_348 (O_348,N_17422,N_17889);
xor UO_349 (O_349,N_15106,N_19785);
nor UO_350 (O_350,N_15144,N_15026);
and UO_351 (O_351,N_18036,N_18069);
or UO_352 (O_352,N_16661,N_17773);
or UO_353 (O_353,N_18349,N_19246);
and UO_354 (O_354,N_19327,N_18803);
xnor UO_355 (O_355,N_15610,N_18088);
nand UO_356 (O_356,N_15829,N_15042);
nand UO_357 (O_357,N_15752,N_17896);
or UO_358 (O_358,N_18740,N_15011);
xor UO_359 (O_359,N_18357,N_17470);
and UO_360 (O_360,N_17545,N_15384);
nand UO_361 (O_361,N_19983,N_18508);
nor UO_362 (O_362,N_19682,N_19253);
or UO_363 (O_363,N_18972,N_17074);
xor UO_364 (O_364,N_17328,N_19898);
nand UO_365 (O_365,N_15336,N_17130);
xnor UO_366 (O_366,N_18314,N_19630);
and UO_367 (O_367,N_17358,N_15580);
nor UO_368 (O_368,N_17959,N_19645);
nor UO_369 (O_369,N_18463,N_18638);
nor UO_370 (O_370,N_17251,N_15063);
nand UO_371 (O_371,N_16141,N_15321);
nor UO_372 (O_372,N_17361,N_17941);
or UO_373 (O_373,N_18313,N_15404);
and UO_374 (O_374,N_16746,N_17404);
xnor UO_375 (O_375,N_18677,N_18795);
and UO_376 (O_376,N_19131,N_15746);
and UO_377 (O_377,N_19496,N_17289);
and UO_378 (O_378,N_18591,N_17863);
xor UO_379 (O_379,N_17982,N_18407);
or UO_380 (O_380,N_17069,N_16574);
nand UO_381 (O_381,N_18497,N_15994);
or UO_382 (O_382,N_16359,N_18814);
nor UO_383 (O_383,N_17085,N_18015);
xor UO_384 (O_384,N_18144,N_19538);
xor UO_385 (O_385,N_18692,N_19468);
nor UO_386 (O_386,N_15443,N_16869);
nand UO_387 (O_387,N_17974,N_15439);
nand UO_388 (O_388,N_15522,N_18009);
xor UO_389 (O_389,N_18259,N_16585);
xnor UO_390 (O_390,N_17402,N_15142);
nor UO_391 (O_391,N_15645,N_18574);
or UO_392 (O_392,N_15216,N_18491);
nand UO_393 (O_393,N_19905,N_18535);
or UO_394 (O_394,N_18550,N_15192);
or UO_395 (O_395,N_18226,N_16350);
nor UO_396 (O_396,N_18204,N_15688);
and UO_397 (O_397,N_17478,N_16024);
nand UO_398 (O_398,N_16542,N_19844);
nor UO_399 (O_399,N_17288,N_18187);
or UO_400 (O_400,N_16468,N_17465);
nor UO_401 (O_401,N_17270,N_16306);
nand UO_402 (O_402,N_18791,N_15163);
xnor UO_403 (O_403,N_19534,N_17774);
xnor UO_404 (O_404,N_19859,N_16402);
nor UO_405 (O_405,N_18525,N_15181);
or UO_406 (O_406,N_17025,N_16100);
and UO_407 (O_407,N_18774,N_19554);
and UO_408 (O_408,N_17189,N_15718);
and UO_409 (O_409,N_18417,N_17030);
xor UO_410 (O_410,N_18742,N_19563);
or UO_411 (O_411,N_18617,N_15686);
xnor UO_412 (O_412,N_15483,N_16255);
xor UO_413 (O_413,N_17581,N_16134);
or UO_414 (O_414,N_17084,N_15654);
nand UO_415 (O_415,N_19358,N_17181);
nand UO_416 (O_416,N_19809,N_17263);
xnor UO_417 (O_417,N_15934,N_19519);
or UO_418 (O_418,N_19461,N_17816);
xnor UO_419 (O_419,N_16645,N_18618);
or UO_420 (O_420,N_15391,N_19420);
nand UO_421 (O_421,N_17698,N_17249);
nand UO_422 (O_422,N_17440,N_19937);
or UO_423 (O_423,N_19656,N_18248);
or UO_424 (O_424,N_19510,N_18221);
nor UO_425 (O_425,N_17253,N_15392);
nor UO_426 (O_426,N_15175,N_17717);
and UO_427 (O_427,N_15428,N_17111);
or UO_428 (O_428,N_15797,N_19680);
nand UO_429 (O_429,N_19421,N_16685);
xnor UO_430 (O_430,N_18370,N_19023);
or UO_431 (O_431,N_15449,N_17104);
or UO_432 (O_432,N_19225,N_16525);
or UO_433 (O_433,N_17845,N_18948);
nor UO_434 (O_434,N_18269,N_18756);
nand UO_435 (O_435,N_18796,N_18785);
or UO_436 (O_436,N_19782,N_19179);
xor UO_437 (O_437,N_19750,N_17619);
or UO_438 (O_438,N_19920,N_17312);
nor UO_439 (O_439,N_18631,N_16890);
xnor UO_440 (O_440,N_16117,N_19570);
and UO_441 (O_441,N_18452,N_19024);
and UO_442 (O_442,N_18289,N_17811);
xor UO_443 (O_443,N_18034,N_17878);
nor UO_444 (O_444,N_17640,N_16994);
or UO_445 (O_445,N_15173,N_17812);
or UO_446 (O_446,N_19674,N_19702);
nor UO_447 (O_447,N_17419,N_15834);
nor UO_448 (O_448,N_17041,N_17029);
or UO_449 (O_449,N_19864,N_17043);
xor UO_450 (O_450,N_16744,N_18706);
nand UO_451 (O_451,N_18245,N_19054);
nor UO_452 (O_452,N_16354,N_19342);
xor UO_453 (O_453,N_19917,N_18641);
and UO_454 (O_454,N_18378,N_17728);
and UO_455 (O_455,N_19047,N_15600);
and UO_456 (O_456,N_17193,N_16821);
and UO_457 (O_457,N_18229,N_17477);
or UO_458 (O_458,N_15307,N_18183);
nand UO_459 (O_459,N_19406,N_16385);
nor UO_460 (O_460,N_18887,N_16379);
or UO_461 (O_461,N_15559,N_19137);
or UO_462 (O_462,N_17233,N_16591);
nand UO_463 (O_463,N_17810,N_17218);
nand UO_464 (O_464,N_15993,N_16474);
xor UO_465 (O_465,N_16683,N_18857);
nor UO_466 (O_466,N_17036,N_16431);
nand UO_467 (O_467,N_17516,N_16908);
and UO_468 (O_468,N_17427,N_19537);
and UO_469 (O_469,N_18600,N_17929);
and UO_470 (O_470,N_15689,N_19058);
nand UO_471 (O_471,N_16347,N_17337);
or UO_472 (O_472,N_16990,N_18863);
and UO_473 (O_473,N_17497,N_17485);
nand UO_474 (O_474,N_15316,N_18346);
nor UO_475 (O_475,N_15859,N_17781);
or UO_476 (O_476,N_16538,N_17088);
and UO_477 (O_477,N_19088,N_18904);
nor UO_478 (O_478,N_16958,N_17028);
nor UO_479 (O_479,N_17550,N_17411);
or UO_480 (O_480,N_17140,N_19780);
xor UO_481 (O_481,N_15915,N_17524);
nor UO_482 (O_482,N_19093,N_16642);
nand UO_483 (O_483,N_16846,N_19022);
or UO_484 (O_484,N_18438,N_15921);
and UO_485 (O_485,N_19735,N_19953);
nand UO_486 (O_486,N_18652,N_17480);
nand UO_487 (O_487,N_18944,N_16153);
nor UO_488 (O_488,N_17594,N_16140);
nand UO_489 (O_489,N_18413,N_16721);
nor UO_490 (O_490,N_18200,N_18170);
or UO_491 (O_491,N_16845,N_15233);
or UO_492 (O_492,N_15223,N_16641);
nand UO_493 (O_493,N_17081,N_18586);
and UO_494 (O_494,N_18274,N_18921);
and UO_495 (O_495,N_16149,N_15831);
xor UO_496 (O_496,N_16090,N_15908);
and UO_497 (O_497,N_18743,N_16480);
nand UO_498 (O_498,N_19360,N_15382);
xor UO_499 (O_499,N_18655,N_15204);
nand UO_500 (O_500,N_19269,N_17540);
nor UO_501 (O_501,N_15048,N_19904);
nor UO_502 (O_502,N_19606,N_16157);
and UO_503 (O_503,N_18102,N_16710);
nor UO_504 (O_504,N_19011,N_19751);
nor UO_505 (O_505,N_17449,N_18606);
nand UO_506 (O_506,N_16521,N_17790);
or UO_507 (O_507,N_17937,N_18444);
and UO_508 (O_508,N_18371,N_19247);
nand UO_509 (O_509,N_16105,N_15310);
nand UO_510 (O_510,N_17826,N_19227);
and UO_511 (O_511,N_18117,N_18934);
nor UO_512 (O_512,N_17955,N_17210);
nor UO_513 (O_513,N_18970,N_18067);
nand UO_514 (O_514,N_16547,N_19930);
nor UO_515 (O_515,N_15720,N_17003);
nor UO_516 (O_516,N_16704,N_18842);
or UO_517 (O_517,N_18118,N_17639);
nor UO_518 (O_518,N_15226,N_18053);
or UO_519 (O_519,N_19721,N_15261);
nand UO_520 (O_520,N_16205,N_15178);
and UO_521 (O_521,N_17780,N_19171);
and UO_522 (O_522,N_18643,N_15036);
nand UO_523 (O_523,N_19999,N_18176);
nor UO_524 (O_524,N_16762,N_19273);
xnor UO_525 (O_525,N_15529,N_18401);
or UO_526 (O_526,N_16785,N_16112);
nand UO_527 (O_527,N_19598,N_17302);
and UO_528 (O_528,N_19470,N_15741);
or UO_529 (O_529,N_19511,N_15275);
xnor UO_530 (O_530,N_15717,N_17742);
and UO_531 (O_531,N_18880,N_19457);
and UO_532 (O_532,N_16798,N_17576);
or UO_533 (O_533,N_19575,N_17128);
xor UO_534 (O_534,N_16263,N_17907);
xor UO_535 (O_535,N_18581,N_17521);
nand UO_536 (O_536,N_17424,N_15653);
xnor UO_537 (O_537,N_18733,N_17142);
or UO_538 (O_538,N_16111,N_18698);
nand UO_539 (O_539,N_17898,N_15972);
nand UO_540 (O_540,N_15700,N_17874);
or UO_541 (O_541,N_16213,N_19053);
xor UO_542 (O_542,N_19901,N_16577);
nand UO_543 (O_543,N_15760,N_15354);
xor UO_544 (O_544,N_15297,N_15608);
nor UO_545 (O_545,N_15547,N_17468);
and UO_546 (O_546,N_17152,N_19843);
xnor UO_547 (O_547,N_17689,N_18555);
or UO_548 (O_548,N_19718,N_16041);
nand UO_549 (O_549,N_19489,N_19757);
nand UO_550 (O_550,N_17155,N_19693);
and UO_551 (O_551,N_19166,N_19228);
and UO_552 (O_552,N_18411,N_17494);
xnor UO_553 (O_553,N_18046,N_19594);
xnor UO_554 (O_554,N_16116,N_19943);
nor UO_555 (O_555,N_16531,N_18116);
and UO_556 (O_556,N_18639,N_18584);
xor UO_557 (O_557,N_18376,N_18268);
and UO_558 (O_558,N_15989,N_17204);
xnor UO_559 (O_559,N_16559,N_15599);
nand UO_560 (O_560,N_15523,N_16028);
nand UO_561 (O_561,N_18512,N_15218);
nand UO_562 (O_562,N_18461,N_15602);
nor UO_563 (O_563,N_19350,N_19633);
nor UO_564 (O_564,N_16127,N_18416);
xor UO_565 (O_565,N_19153,N_15088);
or UO_566 (O_566,N_19888,N_19384);
nand UO_567 (O_567,N_19527,N_19243);
nor UO_568 (O_568,N_19941,N_16974);
and UO_569 (O_569,N_19242,N_19659);
or UO_570 (O_570,N_15821,N_19287);
and UO_571 (O_571,N_19248,N_16437);
nor UO_572 (O_572,N_18205,N_19480);
nand UO_573 (O_573,N_18457,N_19529);
or UO_574 (O_574,N_18372,N_19499);
nor UO_575 (O_575,N_16494,N_15573);
and UO_576 (O_576,N_16254,N_15749);
nand UO_577 (O_577,N_19060,N_15271);
and UO_578 (O_578,N_17561,N_18611);
nand UO_579 (O_579,N_17169,N_16930);
and UO_580 (O_580,N_17651,N_15670);
nand UO_581 (O_581,N_17280,N_18043);
and UO_582 (O_582,N_17163,N_17978);
xor UO_583 (O_583,N_17379,N_18062);
and UO_584 (O_584,N_16768,N_18073);
and UO_585 (O_585,N_17714,N_15920);
xnor UO_586 (O_586,N_18800,N_17064);
nor UO_587 (O_587,N_16274,N_15576);
nor UO_588 (O_588,N_18761,N_17661);
and UO_589 (O_589,N_15311,N_16808);
or UO_590 (O_590,N_16561,N_16755);
xnor UO_591 (O_591,N_17993,N_16327);
and UO_592 (O_592,N_17392,N_19648);
and UO_593 (O_593,N_19947,N_16620);
or UO_594 (O_594,N_16410,N_16673);
xor UO_595 (O_595,N_18347,N_15407);
and UO_596 (O_596,N_15860,N_19739);
and UO_597 (O_597,N_18682,N_16995);
and UO_598 (O_598,N_18971,N_17102);
nor UO_599 (O_599,N_17235,N_17713);
and UO_600 (O_600,N_18235,N_17400);
or UO_601 (O_601,N_19144,N_19439);
nand UO_602 (O_602,N_17217,N_17196);
nor UO_603 (O_603,N_16797,N_19547);
nand UO_604 (O_604,N_15910,N_17984);
nor UO_605 (O_605,N_15198,N_15030);
or UO_606 (O_606,N_17327,N_18764);
nor UO_607 (O_607,N_19918,N_18901);
or UO_608 (O_608,N_19017,N_18730);
and UO_609 (O_609,N_19146,N_19832);
nand UO_610 (O_610,N_17997,N_16891);
or UO_611 (O_611,N_17935,N_18322);
xor UO_612 (O_612,N_18471,N_18310);
or UO_613 (O_613,N_18128,N_18693);
nor UO_614 (O_614,N_19173,N_17229);
and UO_615 (O_615,N_19464,N_18331);
and UO_616 (O_616,N_16094,N_19365);
xnor UO_617 (O_617,N_19256,N_15784);
nor UO_618 (O_618,N_19654,N_16910);
nor UO_619 (O_619,N_16522,N_19056);
xnor UO_620 (O_620,N_17925,N_19042);
xnor UO_621 (O_621,N_15446,N_19968);
and UO_622 (O_622,N_16363,N_18123);
xor UO_623 (O_623,N_17972,N_19581);
xnor UO_624 (O_624,N_16011,N_18623);
xor UO_625 (O_625,N_19156,N_19874);
xnor UO_626 (O_626,N_17394,N_18445);
or UO_627 (O_627,N_18769,N_18396);
or UO_628 (O_628,N_17187,N_16857);
nand UO_629 (O_629,N_15257,N_17047);
nor UO_630 (O_630,N_18177,N_15146);
nor UO_631 (O_631,N_17246,N_17620);
nand UO_632 (O_632,N_17346,N_16396);
xnor UO_633 (O_633,N_18237,N_19134);
or UO_634 (O_634,N_15538,N_18537);
nand UO_635 (O_635,N_16364,N_19445);
nand UO_636 (O_636,N_19579,N_18701);
and UO_637 (O_637,N_15474,N_18056);
or UO_638 (O_638,N_18323,N_17123);
or UO_639 (O_639,N_19004,N_15695);
xnor UO_640 (O_640,N_16824,N_15108);
and UO_641 (O_641,N_15497,N_18100);
and UO_642 (O_642,N_18316,N_16047);
and UO_643 (O_643,N_17244,N_18344);
xnor UO_644 (O_644,N_17808,N_15913);
nand UO_645 (O_645,N_17310,N_18035);
and UO_646 (O_646,N_17799,N_15505);
nor UO_647 (O_647,N_15534,N_16734);
xor UO_648 (O_648,N_15854,N_17022);
nor UO_649 (O_649,N_17892,N_17048);
nand UO_650 (O_650,N_17975,N_19774);
or UO_651 (O_651,N_15374,N_19755);
nor UO_652 (O_652,N_19417,N_16195);
nand UO_653 (O_653,N_19040,N_16715);
nor UO_654 (O_654,N_16811,N_17008);
nor UO_655 (O_655,N_17838,N_16850);
and UO_656 (O_656,N_19963,N_17179);
nand UO_657 (O_657,N_18460,N_15300);
or UO_658 (O_658,N_18251,N_18820);
nor UO_659 (O_659,N_17110,N_15633);
or UO_660 (O_660,N_18683,N_18138);
xor UO_661 (O_661,N_16126,N_16475);
or UO_662 (O_662,N_19770,N_15781);
nor UO_663 (O_663,N_15805,N_15812);
or UO_664 (O_664,N_16378,N_19440);
xor UO_665 (O_665,N_15242,N_15744);
nor UO_666 (O_666,N_17475,N_15751);
xnor UO_667 (O_667,N_19430,N_17254);
nand UO_668 (O_668,N_19133,N_16812);
nand UO_669 (O_669,N_19392,N_17259);
nand UO_670 (O_670,N_17214,N_19613);
or UO_671 (O_671,N_19410,N_18473);
xor UO_672 (O_672,N_19415,N_17643);
nand UO_673 (O_673,N_19710,N_19942);
or UO_674 (O_674,N_16167,N_16628);
nor UO_675 (O_675,N_17557,N_18889);
nand UO_676 (O_676,N_15032,N_18831);
nor UO_677 (O_677,N_15228,N_18663);
xor UO_678 (O_678,N_18258,N_18109);
xor UO_679 (O_679,N_19348,N_19856);
nand UO_680 (O_680,N_19629,N_19652);
nor UO_681 (O_681,N_15025,N_18499);
or UO_682 (O_682,N_15299,N_16211);
nand UO_683 (O_683,N_16332,N_16032);
nor UO_684 (O_684,N_18467,N_19883);
and UO_685 (O_685,N_15808,N_17413);
or UO_686 (O_686,N_17671,N_18619);
nand UO_687 (O_687,N_16064,N_18536);
and UO_688 (O_688,N_15487,N_18728);
xor UO_689 (O_689,N_19595,N_19500);
nor UO_690 (O_690,N_18214,N_19727);
xnor UO_691 (O_691,N_15506,N_17862);
nor UO_692 (O_692,N_17716,N_15949);
or UO_693 (O_693,N_16688,N_18078);
nand UO_694 (O_694,N_15331,N_17407);
or UO_695 (O_695,N_18448,N_17706);
xnor UO_696 (O_696,N_16413,N_15673);
xnor UO_697 (O_697,N_15456,N_18940);
and UO_698 (O_698,N_17112,N_17355);
or UO_699 (O_699,N_15434,N_15804);
and UO_700 (O_700,N_16085,N_15421);
xor UO_701 (O_701,N_18968,N_16997);
xnor UO_702 (O_702,N_19010,N_16537);
nand UO_703 (O_703,N_18060,N_15935);
and UO_704 (O_704,N_18152,N_15151);
and UO_705 (O_705,N_15897,N_15753);
xnor UO_706 (O_706,N_15698,N_16010);
or UO_707 (O_707,N_19677,N_18219);
nor UO_708 (O_708,N_17425,N_18992);
xnor UO_709 (O_709,N_19967,N_19082);
or UO_710 (O_710,N_19190,N_16103);
nor UO_711 (O_711,N_19008,N_18494);
or UO_712 (O_712,N_19665,N_17635);
and UO_713 (O_713,N_17454,N_15557);
or UO_714 (O_714,N_18562,N_17888);
xnor UO_715 (O_715,N_16551,N_18949);
nor UO_716 (O_716,N_18825,N_15838);
and UO_717 (O_717,N_16831,N_16446);
nand UO_718 (O_718,N_17527,N_16800);
or UO_719 (O_719,N_16731,N_18266);
and UO_720 (O_720,N_17430,N_15546);
nor UO_721 (O_721,N_15058,N_16924);
xnor UO_722 (O_722,N_15619,N_18822);
or UO_723 (O_723,N_16652,N_18767);
nor UO_724 (O_724,N_16786,N_19080);
nor UO_725 (O_725,N_15349,N_17272);
nand UO_726 (O_726,N_19518,N_17040);
and UO_727 (O_727,N_15195,N_19119);
or UO_728 (O_728,N_19478,N_15393);
nor UO_729 (O_729,N_15780,N_15306);
and UO_730 (O_730,N_16926,N_19063);
nand UO_731 (O_731,N_17247,N_19294);
nor UO_732 (O_732,N_19395,N_15641);
nor UO_733 (O_733,N_15319,N_17829);
and UO_734 (O_734,N_19670,N_16204);
nor UO_735 (O_735,N_19873,N_17153);
nand UO_736 (O_736,N_19103,N_16593);
and UO_737 (O_737,N_16978,N_17080);
xnor UO_738 (O_738,N_17569,N_19385);
nor UO_739 (O_739,N_15176,N_18801);
xnor UO_740 (O_740,N_15420,N_16695);
or UO_741 (O_741,N_16430,N_15197);
xnor UO_742 (O_742,N_16697,N_17293);
nand UO_743 (O_743,N_15651,N_16835);
xnor UO_744 (O_744,N_19451,N_18418);
nor UO_745 (O_745,N_16404,N_19170);
and UO_746 (O_746,N_19456,N_17418);
xnor UO_747 (O_747,N_18644,N_15136);
or UO_748 (O_748,N_16478,N_17171);
nand UO_749 (O_749,N_18841,N_19473);
and UO_750 (O_750,N_16804,N_17991);
nor UO_751 (O_751,N_18963,N_16907);
or UO_752 (O_752,N_15621,N_18810);
xor UO_753 (O_753,N_18885,N_18998);
nor UO_754 (O_754,N_18813,N_19099);
xor UO_755 (O_755,N_18379,N_19882);
and UO_756 (O_756,N_19700,N_15982);
xor UO_757 (O_757,N_19094,N_15085);
and UO_758 (O_758,N_15842,N_18160);
nor UO_759 (O_759,N_15706,N_16788);
nand UO_760 (O_760,N_15833,N_19834);
or UO_761 (O_761,N_19282,N_17274);
xnor UO_762 (O_762,N_16981,N_17176);
or UO_763 (O_763,N_18783,N_16533);
nor UO_764 (O_764,N_19009,N_16662);
or UO_765 (O_765,N_15914,N_17282);
and UO_766 (O_766,N_15253,N_15000);
nand UO_767 (O_767,N_18747,N_19779);
or UO_768 (O_768,N_16625,N_15418);
xnor UO_769 (O_769,N_19673,N_18239);
nor UO_770 (O_770,N_19167,N_19651);
and UO_771 (O_771,N_18561,N_16110);
and UO_772 (O_772,N_18571,N_16461);
or UO_773 (O_773,N_19769,N_17161);
nor UO_774 (O_774,N_15442,N_15937);
xor UO_775 (O_775,N_17262,N_15657);
or UO_776 (O_776,N_16427,N_16190);
and UO_777 (O_777,N_18270,N_15411);
nand UO_778 (O_778,N_18315,N_15454);
nand UO_779 (O_779,N_15588,N_18543);
and UO_780 (O_780,N_15664,N_19891);
nor UO_781 (O_781,N_19236,N_18753);
or UO_782 (O_782,N_18724,N_18439);
or UO_783 (O_783,N_17782,N_16859);
nor UO_784 (O_784,N_18025,N_19340);
or UO_785 (O_785,N_15478,N_15904);
xnor UO_786 (O_786,N_15230,N_15884);
nand UO_787 (O_787,N_17768,N_18580);
nor UO_788 (O_788,N_18627,N_16941);
and UO_789 (O_789,N_15918,N_16014);
and UO_790 (O_790,N_19345,N_19396);
nor UO_791 (O_791,N_15145,N_15618);
nand UO_792 (O_792,N_15432,N_15422);
or UO_793 (O_793,N_16145,N_16281);
or UO_794 (O_794,N_16725,N_18656);
nor UO_795 (O_795,N_19343,N_15863);
xor UO_796 (O_796,N_18425,N_17119);
or UO_797 (O_797,N_16690,N_17800);
xnor UO_798 (O_798,N_18326,N_19381);
xnor UO_799 (O_799,N_19536,N_18135);
and UO_800 (O_800,N_18377,N_16977);
nor UO_801 (O_801,N_15274,N_15090);
xnor UO_802 (O_802,N_17467,N_15806);
and UO_803 (O_803,N_16421,N_16042);
and UO_804 (O_804,N_18702,N_15539);
xor UO_805 (O_805,N_15091,N_16892);
and UO_806 (O_806,N_17542,N_19231);
nand UO_807 (O_807,N_19184,N_15445);
xor UO_808 (O_808,N_16043,N_16668);
or UO_809 (O_809,N_19279,N_15305);
nand UO_810 (O_810,N_19312,N_16302);
nor UO_811 (O_811,N_19454,N_19615);
nand UO_812 (O_812,N_19130,N_15770);
or UO_813 (O_813,N_18615,N_16793);
and UO_814 (O_814,N_19975,N_17121);
nor UO_815 (O_815,N_15231,N_16669);
xor UO_816 (O_816,N_19719,N_17860);
or UO_817 (O_817,N_16572,N_15627);
and UO_818 (O_818,N_17113,N_18598);
nor UO_819 (O_819,N_19293,N_18382);
xnor UO_820 (O_820,N_18625,N_17297);
nand UO_821 (O_821,N_17750,N_15046);
and UO_822 (O_822,N_16614,N_15524);
and UO_823 (O_823,N_18437,N_16483);
or UO_824 (O_824,N_19129,N_18654);
or UO_825 (O_825,N_18127,N_16432);
nand UO_826 (O_826,N_16904,N_18797);
nor UO_827 (O_827,N_19961,N_19827);
xnor UO_828 (O_828,N_17077,N_19393);
nand UO_829 (O_829,N_15342,N_18709);
nand UO_830 (O_830,N_19244,N_16557);
and UO_831 (O_831,N_19792,N_19338);
or UO_832 (O_832,N_18032,N_19316);
xor UO_833 (O_833,N_17623,N_16498);
or UO_834 (O_834,N_19382,N_19902);
nor UO_835 (O_835,N_17232,N_16114);
nand UO_836 (O_836,N_17998,N_15107);
and UO_837 (O_837,N_16881,N_16202);
xor UO_838 (O_838,N_18920,N_17500);
xnor UO_839 (O_839,N_16592,N_17727);
xor UO_840 (O_840,N_19152,N_18858);
or UO_841 (O_841,N_15855,N_16349);
nand UO_842 (O_842,N_15755,N_15053);
nor UO_843 (O_843,N_18294,N_17026);
nand UO_844 (O_844,N_19807,N_18517);
xnor UO_845 (O_845,N_19065,N_15841);
or UO_846 (O_846,N_19121,N_17448);
nor UO_847 (O_847,N_16406,N_16584);
and UO_848 (O_848,N_17105,N_17901);
and UO_849 (O_849,N_15099,N_16083);
nor UO_850 (O_850,N_18980,N_18751);
nand UO_851 (O_851,N_18154,N_15896);
xor UO_852 (O_852,N_17370,N_19743);
and UO_853 (O_853,N_15034,N_18843);
and UO_854 (O_854,N_15814,N_15598);
and UO_855 (O_855,N_15196,N_15128);
or UO_856 (O_856,N_15614,N_19070);
nor UO_857 (O_857,N_19923,N_17677);
and UO_858 (O_858,N_18680,N_19260);
xor UO_859 (O_859,N_16839,N_15477);
xor UO_860 (O_860,N_18798,N_18534);
xor UO_861 (O_861,N_16509,N_17261);
xor UO_862 (O_862,N_17071,N_15594);
nor UO_863 (O_863,N_15070,N_19375);
nand UO_864 (O_864,N_19373,N_15167);
xor UO_865 (O_865,N_17101,N_15179);
or UO_866 (O_866,N_19344,N_18522);
and UO_867 (O_867,N_15491,N_15561);
xnor UO_868 (O_868,N_16587,N_16896);
nor UO_869 (O_869,N_16947,N_16968);
xor UO_870 (O_870,N_15674,N_16961);
nand UO_871 (O_871,N_16946,N_19290);
xor UO_872 (O_872,N_15406,N_16333);
nor UO_873 (O_873,N_18609,N_15323);
nor UO_874 (O_874,N_18093,N_15464);
nand UO_875 (O_875,N_17395,N_16988);
nor UO_876 (O_876,N_18363,N_17330);
and UO_877 (O_877,N_19791,N_19829);
nand UO_878 (O_878,N_19095,N_17011);
and UO_879 (O_879,N_16973,N_17656);
and UO_880 (O_880,N_16508,N_17737);
nand UO_881 (O_881,N_19416,N_17343);
or UO_882 (O_882,N_18830,N_17541);
or UO_883 (O_883,N_19466,N_18962);
nor UO_884 (O_884,N_19544,N_19226);
nor UO_885 (O_885,N_15708,N_18794);
nand UO_886 (O_886,N_15988,N_16201);
xnor UO_887 (O_887,N_15475,N_19083);
nand UO_888 (O_888,N_15736,N_17535);
nand UO_889 (O_889,N_17049,N_15281);
nor UO_890 (O_890,N_15276,N_16034);
nand UO_891 (O_891,N_18678,N_18141);
xor UO_892 (O_892,N_17183,N_17501);
nand UO_893 (O_893,N_16780,N_15870);
nor UO_894 (O_894,N_19157,N_16594);
xnor UO_895 (O_895,N_16328,N_19880);
and UO_896 (O_896,N_16936,N_15335);
xnor UO_897 (O_897,N_16801,N_16253);
nand UO_898 (O_898,N_18039,N_16764);
or UO_899 (O_899,N_17752,N_15527);
nor UO_900 (O_900,N_16922,N_15018);
and UO_901 (O_901,N_15493,N_16659);
xor UO_902 (O_902,N_16756,N_16234);
nor UO_903 (O_903,N_16672,N_18208);
nor UO_904 (O_904,N_18545,N_16284);
xnor UO_905 (O_905,N_17647,N_19712);
and UO_906 (O_906,N_16758,N_16611);
nand UO_907 (O_907,N_17663,N_15069);
and UO_908 (O_908,N_17734,N_18988);
and UO_909 (O_909,N_17908,N_16293);
and UO_910 (O_910,N_15169,N_19357);
nor UO_911 (O_911,N_19297,N_18847);
nand UO_912 (O_912,N_19607,N_19705);
nor UO_913 (O_913,N_15631,N_18010);
xnor UO_914 (O_914,N_15775,N_18960);
and UO_915 (O_915,N_15283,N_16751);
and UO_916 (O_916,N_18423,N_16179);
and UO_917 (O_917,N_15636,N_18533);
nor UO_918 (O_918,N_17880,N_19543);
xnor UO_919 (O_919,N_16266,N_15992);
nor UO_920 (O_920,N_18077,N_15158);
and UO_921 (O_921,N_18318,N_19469);
xor UO_922 (O_922,N_17824,N_19850);
or UO_923 (O_923,N_18277,N_15471);
or UO_924 (O_924,N_15014,N_15517);
and UO_925 (O_925,N_15122,N_19541);
nand UO_926 (O_926,N_16272,N_15583);
xor UO_927 (O_927,N_15425,N_18190);
xnor UO_928 (O_928,N_15585,N_18210);
or UO_929 (O_929,N_19202,N_15774);
nand UO_930 (O_930,N_17721,N_19608);
xnor UO_931 (O_931,N_16790,N_17828);
nand UO_932 (O_932,N_19846,N_17872);
nand UO_933 (O_933,N_19433,N_16775);
xor UO_934 (O_934,N_16919,N_19761);
xnor UO_935 (O_935,N_15207,N_19573);
nand UO_936 (O_936,N_18354,N_16560);
and UO_937 (O_937,N_18506,N_19593);
nand UO_938 (O_938,N_17340,N_15498);
and UO_939 (O_939,N_17227,N_18105);
nor UO_940 (O_940,N_16914,N_15489);
or UO_941 (O_941,N_16479,N_19535);
and UO_942 (O_942,N_19872,N_17382);
and UO_943 (O_943,N_19664,N_15463);
xor UO_944 (O_944,N_17772,N_17711);
nor UO_945 (O_945,N_17948,N_16390);
xor UO_946 (O_946,N_19139,N_19032);
nand UO_947 (O_947,N_18540,N_16870);
nor UO_948 (O_948,N_17970,N_19217);
nor UO_949 (O_949,N_17947,N_17103);
and UO_950 (O_950,N_17745,N_19740);
nor UO_951 (O_951,N_16236,N_19909);
xor UO_952 (O_952,N_19612,N_18645);
or UO_953 (O_953,N_16727,N_15726);
nand UO_954 (O_954,N_18705,N_17950);
or UO_955 (O_955,N_18547,N_17225);
nor UO_956 (O_956,N_16216,N_15468);
nand UO_957 (O_957,N_19163,N_19966);
xor UO_958 (O_958,N_18582,N_17076);
xor UO_959 (O_959,N_15738,N_17669);
and UO_960 (O_960,N_19181,N_19303);
and UO_961 (O_961,N_17248,N_15579);
nand UO_962 (O_962,N_15852,N_19528);
nor UO_963 (O_963,N_18358,N_17314);
nor UO_964 (O_964,N_15356,N_15634);
nor UO_965 (O_965,N_15237,N_16139);
xnor UO_966 (O_966,N_19765,N_15876);
or UO_967 (O_967,N_15613,N_15209);
xnor UO_968 (O_968,N_15548,N_19890);
nand UO_969 (O_969,N_17632,N_19845);
xnor UO_970 (O_970,N_16232,N_19061);
nand UO_971 (O_971,N_18739,N_15590);
xor UO_972 (O_972,N_15671,N_19549);
and UO_973 (O_973,N_18052,N_16393);
or UO_974 (O_974,N_18725,N_19762);
nand UO_975 (O_975,N_15824,N_17637);
nand UO_976 (O_976,N_19747,N_19955);
and UO_977 (O_977,N_17786,N_18332);
nor UO_978 (O_978,N_15721,N_18163);
nor UO_979 (O_979,N_19572,N_17853);
xnor UO_980 (O_980,N_15080,N_16753);
nand UO_981 (O_981,N_15624,N_18882);
xnor UO_982 (O_982,N_18050,N_18964);
or UO_983 (O_983,N_18014,N_15448);
xor UO_984 (O_984,N_16425,N_17132);
or UO_985 (O_985,N_18670,N_15520);
or UO_986 (O_986,N_16290,N_15991);
or UO_987 (O_987,N_16813,N_16917);
nand UO_988 (O_988,N_16007,N_18630);
and UO_989 (O_989,N_19863,N_15905);
nor UO_990 (O_990,N_19349,N_15998);
nand UO_991 (O_991,N_19113,N_18424);
or UO_992 (O_992,N_19328,N_18969);
xor UO_993 (O_993,N_16589,N_16000);
and UO_994 (O_994,N_18375,N_18450);
and UO_995 (O_995,N_17384,N_17461);
xor UO_996 (O_996,N_16597,N_16399);
xnor UO_997 (O_997,N_18472,N_18513);
and UO_998 (O_998,N_18419,N_15089);
xor UO_999 (O_999,N_18950,N_19320);
or UO_1000 (O_1000,N_16860,N_16426);
nand UO_1001 (O_1001,N_16830,N_18155);
and UO_1002 (O_1002,N_16834,N_15414);
xor UO_1003 (O_1003,N_19686,N_16182);
xor UO_1004 (O_1004,N_15143,N_16803);
and UO_1005 (O_1005,N_15939,N_18114);
or UO_1006 (O_1006,N_17344,N_18011);
xor UO_1007 (O_1007,N_15482,N_18777);
and UO_1008 (O_1008,N_18917,N_19158);
nor UO_1009 (O_1009,N_19232,N_15055);
and UO_1010 (O_1010,N_19949,N_15581);
and UO_1011 (O_1011,N_17349,N_18930);
nor UO_1012 (O_1012,N_18410,N_18306);
and UO_1013 (O_1013,N_17381,N_16056);
and UO_1014 (O_1014,N_17223,N_17989);
and UO_1015 (O_1015,N_19336,N_18990);
or UO_1016 (O_1016,N_18662,N_18180);
and UO_1017 (O_1017,N_15252,N_19259);
and UO_1018 (O_1018,N_16348,N_15150);
nand UO_1019 (O_1019,N_15325,N_16313);
nand UO_1020 (O_1020,N_16605,N_15102);
nand UO_1021 (O_1021,N_16409,N_15470);
nor UO_1022 (O_1022,N_17457,N_18465);
and UO_1023 (O_1023,N_19206,N_19894);
nand UO_1024 (O_1024,N_16174,N_15981);
xor UO_1025 (O_1025,N_16879,N_16228);
xor UO_1026 (O_1026,N_16222,N_15591);
xnor UO_1027 (O_1027,N_17226,N_16488);
nor UO_1028 (O_1028,N_16543,N_16356);
nor UO_1029 (O_1029,N_19697,N_18688);
and UO_1030 (O_1030,N_16271,N_17058);
and UO_1031 (O_1031,N_19402,N_16503);
xor UO_1032 (O_1032,N_19471,N_16658);
or UO_1033 (O_1033,N_19892,N_15433);
xnor UO_1034 (O_1034,N_17775,N_16020);
nand UO_1035 (O_1035,N_17014,N_15078);
nor UO_1036 (O_1036,N_18649,N_15519);
nor UO_1037 (O_1037,N_15156,N_17267);
nor UO_1038 (O_1038,N_15168,N_17117);
xnor UO_1039 (O_1039,N_16452,N_15229);
nand UO_1040 (O_1040,N_19049,N_18242);
and UO_1041 (O_1041,N_17654,N_16583);
xnor UO_1042 (O_1042,N_15555,N_18311);
or UO_1043 (O_1043,N_15236,N_17886);
nor UO_1044 (O_1044,N_15329,N_15390);
xor UO_1045 (O_1045,N_15742,N_17466);
nor UO_1046 (O_1046,N_15479,N_19138);
and UO_1047 (O_1047,N_18096,N_18000);
or UO_1048 (O_1048,N_16623,N_17450);
nand UO_1049 (O_1049,N_19150,N_15601);
xor UO_1050 (O_1050,N_17488,N_18925);
and UO_1051 (O_1051,N_15866,N_15880);
xor UO_1052 (O_1052,N_16700,N_19614);
nand UO_1053 (O_1053,N_18362,N_17976);
or UO_1054 (O_1054,N_18507,N_15444);
nor UO_1055 (O_1055,N_18284,N_19748);
or UO_1056 (O_1056,N_19701,N_18133);
and UO_1057 (O_1057,N_17847,N_19005);
xnor UO_1058 (O_1058,N_19822,N_19929);
xor UO_1059 (O_1059,N_19502,N_18408);
nor UO_1060 (O_1060,N_15637,N_16207);
xnor UO_1061 (O_1061,N_19207,N_19302);
nor UO_1062 (O_1062,N_18291,N_18302);
nand UO_1063 (O_1063,N_15077,N_19795);
nand UO_1064 (O_1064,N_16646,N_15419);
nand UO_1065 (O_1065,N_17510,N_17763);
and UO_1066 (O_1066,N_15759,N_18906);
nor UO_1067 (O_1067,N_15881,N_16256);
xor UO_1068 (O_1068,N_17498,N_17433);
xnor UO_1069 (O_1069,N_16847,N_18549);
xor UO_1070 (O_1070,N_18309,N_19453);
and UO_1071 (O_1071,N_15370,N_17741);
or UO_1072 (O_1072,N_18585,N_16492);
or UO_1073 (O_1073,N_15871,N_19209);
nor UO_1074 (O_1074,N_15542,N_16633);
nor UO_1075 (O_1075,N_15819,N_19492);
nand UO_1076 (O_1076,N_16603,N_18085);
xor UO_1077 (O_1077,N_15451,N_19988);
nand UO_1078 (O_1078,N_17797,N_15182);
and UO_1079 (O_1079,N_15353,N_15452);
or UO_1080 (O_1080,N_19034,N_18862);
nand UO_1081 (O_1081,N_17164,N_15768);
xnor UO_1082 (O_1082,N_19505,N_16921);
or UO_1083 (O_1083,N_15037,N_16436);
xor UO_1084 (O_1084,N_19621,N_18653);
or UO_1085 (O_1085,N_15084,N_15973);
xnor UO_1086 (O_1086,N_19048,N_18918);
nor UO_1087 (O_1087,N_18453,N_19201);
nand UO_1088 (O_1088,N_15668,N_18167);
nand UO_1089 (O_1089,N_16317,N_19948);
or UO_1090 (O_1090,N_16023,N_18477);
nand UO_1091 (O_1091,N_16855,N_17923);
and UO_1092 (O_1092,N_17126,N_19383);
nor UO_1093 (O_1093,N_17547,N_17980);
nand UO_1094 (O_1094,N_16143,N_18198);
xnor UO_1095 (O_1095,N_18479,N_19893);
xor UO_1096 (O_1096,N_18162,N_18861);
xnor UO_1097 (O_1097,N_15563,N_16146);
nand UO_1098 (O_1098,N_19436,N_17645);
nor UO_1099 (O_1099,N_16048,N_16277);
and UO_1100 (O_1100,N_15690,N_18560);
xnor UO_1101 (O_1101,N_18787,N_17746);
nor UO_1102 (O_1102,N_19465,N_18772);
nand UO_1103 (O_1103,N_16883,N_18024);
nor UO_1104 (O_1104,N_16598,N_16631);
nand UO_1105 (O_1105,N_15667,N_16463);
or UO_1106 (O_1106,N_17086,N_19831);
nor UO_1107 (O_1107,N_18812,N_18824);
xor UO_1108 (O_1108,N_17325,N_19749);
nor UO_1109 (O_1109,N_19233,N_19084);
xnor UO_1110 (O_1110,N_15183,N_16838);
nor UO_1111 (O_1111,N_15974,N_17486);
nor UO_1112 (O_1112,N_17821,N_16794);
nand UO_1113 (O_1113,N_16131,N_15632);
nor UO_1114 (O_1114,N_18983,N_18002);
nand UO_1115 (O_1115,N_17881,N_19932);
or UO_1116 (O_1116,N_16829,N_16325);
nand UO_1117 (O_1117,N_16677,N_16036);
or UO_1118 (O_1118,N_15743,N_15017);
nand UO_1119 (O_1119,N_17707,N_19325);
nand UO_1120 (O_1120,N_18381,N_19945);
nor UO_1121 (O_1121,N_15154,N_17037);
and UO_1122 (O_1122,N_17258,N_17303);
nor UO_1123 (O_1123,N_17211,N_18360);
nand UO_1124 (O_1124,N_15515,N_19509);
nand UO_1125 (O_1125,N_18215,N_16215);
or UO_1126 (O_1126,N_16342,N_15427);
or UO_1127 (O_1127,N_17822,N_19801);
or UO_1128 (O_1128,N_15560,N_18744);
nor UO_1129 (O_1129,N_15707,N_15541);
nand UO_1130 (O_1130,N_15567,N_16826);
nand UO_1131 (O_1131,N_15199,N_16809);
nor UO_1132 (O_1132,N_17666,N_16501);
xor UO_1133 (O_1133,N_18632,N_15002);
and UO_1134 (O_1134,N_17359,N_15205);
or UO_1135 (O_1135,N_17360,N_17548);
nor UO_1136 (O_1136,N_17570,N_18758);
or UO_1137 (O_1137,N_17658,N_19114);
xnor UO_1138 (O_1138,N_17725,N_18345);
nor UO_1139 (O_1139,N_18737,N_18552);
nand UO_1140 (O_1140,N_18855,N_15417);
or UO_1141 (O_1141,N_16270,N_15983);
nor UO_1142 (O_1142,N_18958,N_16496);
nor UO_1143 (O_1143,N_17405,N_16774);
xnor UO_1144 (O_1144,N_16440,N_18699);
or UO_1145 (O_1145,N_19703,N_15165);
and UO_1146 (O_1146,N_17338,N_17865);
and UO_1147 (O_1147,N_16943,N_18218);
nor UO_1148 (O_1148,N_19261,N_17852);
or UO_1149 (O_1149,N_17525,N_19307);
nor UO_1150 (O_1150,N_18884,N_15339);
nor UO_1151 (O_1151,N_17933,N_16730);
nor UO_1152 (O_1152,N_16104,N_18780);
and UO_1153 (O_1153,N_19778,N_15027);
nand UO_1154 (O_1154,N_19334,N_19364);
nor UO_1155 (O_1155,N_19603,N_16552);
or UO_1156 (O_1156,N_18188,N_17459);
and UO_1157 (O_1157,N_17116,N_17172);
or UO_1158 (O_1158,N_18836,N_18264);
nand UO_1159 (O_1159,N_17141,N_17412);
or UO_1160 (O_1160,N_19560,N_19311);
xor UO_1161 (O_1161,N_18658,N_15103);
nand UO_1162 (O_1162,N_17604,N_15431);
xor UO_1163 (O_1163,N_17699,N_15731);
nor UO_1164 (O_1164,N_19913,N_17608);
nor UO_1165 (O_1165,N_18495,N_18359);
and UO_1166 (O_1166,N_17504,N_16541);
or UO_1167 (O_1167,N_17877,N_16147);
nand UO_1168 (O_1168,N_15617,N_15009);
nor UO_1169 (O_1169,N_19933,N_18687);
nand UO_1170 (O_1170,N_16637,N_16856);
nand UO_1171 (O_1171,N_18765,N_17205);
nor UO_1172 (O_1172,N_16084,N_15801);
xor UO_1173 (O_1173,N_16949,N_18579);
and UO_1174 (O_1174,N_17455,N_15054);
and UO_1175 (O_1175,N_17562,N_18225);
xnor UO_1176 (O_1176,N_17252,N_15476);
nor UO_1177 (O_1177,N_15639,N_15337);
nand UO_1178 (O_1178,N_17911,N_17035);
nor UO_1179 (O_1179,N_19636,N_18279);
xor UO_1180 (O_1180,N_19927,N_19797);
and UO_1181 (O_1181,N_19039,N_18216);
xnor UO_1182 (O_1182,N_19881,N_18939);
nand UO_1183 (O_1183,N_15132,N_19766);
or UO_1184 (O_1184,N_18400,N_17512);
and UO_1185 (O_1185,N_19663,N_16863);
or UO_1186 (O_1186,N_18500,N_19346);
xor UO_1187 (O_1187,N_15823,N_18546);
and UO_1188 (O_1188,N_16169,N_17144);
nor UO_1189 (O_1189,N_15589,N_17897);
nor UO_1190 (O_1190,N_19128,N_15809);
xnor UO_1191 (O_1191,N_16959,N_19851);
xnor UO_1192 (O_1192,N_17476,N_15095);
or UO_1193 (O_1193,N_16088,N_16175);
and UO_1194 (O_1194,N_18987,N_15380);
and UO_1195 (O_1195,N_16705,N_15288);
nand UO_1196 (O_1196,N_15502,N_19109);
nand UO_1197 (O_1197,N_19006,N_18961);
nand UO_1198 (O_1198,N_19737,N_19524);
nor UO_1199 (O_1199,N_18727,N_17157);
or UO_1200 (O_1200,N_18738,N_15457);
nand UO_1201 (O_1201,N_15267,N_16227);
xor UO_1202 (O_1202,N_15206,N_18110);
or UO_1203 (O_1203,N_19815,N_19639);
xor UO_1204 (O_1204,N_19626,N_19370);
nor UO_1205 (O_1205,N_18704,N_18827);
nor UO_1206 (O_1206,N_19286,N_15623);
xor UO_1207 (O_1207,N_15928,N_15028);
xor UO_1208 (O_1208,N_17366,N_18721);
and UO_1209 (O_1209,N_19627,N_19101);
nand UO_1210 (O_1210,N_17365,N_18017);
and UO_1211 (O_1211,N_19814,N_18045);
or UO_1212 (O_1212,N_15269,N_15782);
nor UO_1213 (O_1213,N_16442,N_18568);
or UO_1214 (O_1214,N_17792,N_17129);
and UO_1215 (O_1215,N_17981,N_16989);
and UO_1216 (O_1216,N_15246,N_18327);
nor UO_1217 (O_1217,N_17095,N_15320);
and UO_1218 (O_1218,N_15754,N_19584);
nand UO_1219 (O_1219,N_18171,N_19180);
and UO_1220 (O_1220,N_16868,N_19921);
or UO_1221 (O_1221,N_17618,N_16080);
nor UO_1222 (O_1222,N_15075,N_16815);
nand UO_1223 (O_1223,N_18636,N_16206);
and UO_1224 (O_1224,N_17316,N_19732);
xnor UO_1225 (O_1225,N_19027,N_15024);
or UO_1226 (O_1226,N_18185,N_16076);
or UO_1227 (O_1227,N_18931,N_18514);
nand UO_1228 (O_1228,N_19448,N_16511);
nor UO_1229 (O_1229,N_17464,N_18569);
xor UO_1230 (O_1230,N_16945,N_18676);
nand UO_1231 (O_1231,N_18607,N_19640);
or UO_1232 (O_1232,N_18624,N_18539);
or UO_1233 (O_1233,N_18489,N_15728);
or UO_1234 (O_1234,N_17791,N_15593);
xor UO_1235 (O_1235,N_16733,N_16335);
xnor UO_1236 (O_1236,N_19272,N_15399);
or UO_1237 (O_1237,N_18908,N_19973);
or UO_1238 (O_1238,N_16345,N_18429);
nand UO_1239 (O_1239,N_15659,N_15604);
xor UO_1240 (O_1240,N_18061,N_18016);
nand UO_1241 (O_1241,N_15716,N_19854);
nor UO_1242 (O_1242,N_17867,N_15180);
or UO_1243 (O_1243,N_18432,N_18250);
and UO_1244 (O_1244,N_19915,N_18951);
or UO_1245 (O_1245,N_18092,N_15582);
xnor UO_1246 (O_1246,N_17633,N_19106);
nand UO_1247 (O_1247,N_18456,N_19722);
xnor UO_1248 (O_1248,N_16570,N_19437);
xor UO_1249 (O_1249,N_15646,N_18063);
nor UO_1250 (O_1250,N_17044,N_16453);
or UO_1251 (O_1251,N_19193,N_15830);
and UO_1252 (O_1252,N_17507,N_19043);
nand UO_1253 (O_1253,N_16515,N_15277);
nor UO_1254 (O_1254,N_16151,N_17875);
xnor UO_1255 (O_1255,N_16622,N_19353);
nand UO_1256 (O_1256,N_18055,N_19836);
nor UO_1257 (O_1257,N_18244,N_18563);
nor UO_1258 (O_1258,N_19819,N_15840);
or UO_1259 (O_1259,N_15450,N_18722);
or UO_1260 (O_1260,N_16299,N_19029);
and UO_1261 (O_1261,N_17426,N_15874);
nor UO_1262 (O_1262,N_18257,N_16510);
nor UO_1263 (O_1263,N_15971,N_16021);
nor UO_1264 (O_1264,N_17145,N_17566);
and UO_1265 (O_1265,N_15480,N_17761);
xor UO_1266 (O_1266,N_16723,N_15447);
and UO_1267 (O_1267,N_18018,N_19745);
and UO_1268 (O_1268,N_15836,N_15923);
nor UO_1269 (O_1269,N_19162,N_16739);
and UO_1270 (O_1270,N_19990,N_16233);
nand UO_1271 (O_1271,N_19310,N_17490);
nand UO_1272 (O_1272,N_19753,N_19658);
nand UO_1273 (O_1273,N_16337,N_19266);
and UO_1274 (O_1274,N_15995,N_16639);
or UO_1275 (O_1275,N_17057,N_18700);
xor UO_1276 (O_1276,N_19728,N_15739);
or UO_1277 (O_1277,N_17776,N_17094);
or UO_1278 (O_1278,N_17479,N_15332);
nor UO_1279 (O_1279,N_16231,N_16185);
or UO_1280 (O_1280,N_17928,N_17973);
and UO_1281 (O_1281,N_15678,N_19940);
and UO_1282 (O_1282,N_15114,N_19003);
nand UO_1283 (O_1283,N_16297,N_19687);
nand UO_1284 (O_1284,N_18131,N_19442);
and UO_1285 (O_1285,N_18746,N_16199);
and UO_1286 (O_1286,N_16858,N_15577);
nor UO_1287 (O_1287,N_16473,N_16565);
and UO_1288 (O_1288,N_18668,N_19361);
nor UO_1289 (O_1289,N_15313,N_17055);
or UO_1290 (O_1290,N_19016,N_16599);
and UO_1291 (O_1291,N_16443,N_15235);
or UO_1292 (O_1292,N_16708,N_15007);
or UO_1293 (O_1293,N_17373,N_17758);
and UO_1294 (O_1294,N_18926,N_19969);
or UO_1295 (O_1295,N_17703,N_15174);
or UO_1296 (O_1296,N_17481,N_15592);
nor UO_1297 (O_1297,N_15255,N_18895);
nand UO_1298 (O_1298,N_18519,N_17323);
nand UO_1299 (O_1299,N_17528,N_15105);
nand UO_1300 (O_1300,N_16003,N_18415);
or UO_1301 (O_1301,N_17447,N_16951);
or UO_1302 (O_1302,N_17944,N_18669);
and UO_1303 (O_1303,N_18246,N_18864);
or UO_1304 (O_1304,N_16689,N_17100);
or UO_1305 (O_1305,N_15779,N_16156);
xor UO_1306 (O_1306,N_19562,N_15061);
and UO_1307 (O_1307,N_16983,N_17091);
nand UO_1308 (O_1308,N_18191,N_18068);
and UO_1309 (O_1309,N_18335,N_18778);
xor UO_1310 (O_1310,N_16491,N_18165);
or UO_1311 (O_1311,N_17807,N_15750);
and UO_1312 (O_1312,N_16817,N_18605);
nand UO_1313 (O_1313,N_16528,N_17904);
xor UO_1314 (O_1314,N_18719,N_16853);
nand UO_1315 (O_1315,N_18071,N_16183);
or UO_1316 (O_1316,N_16872,N_18828);
nor UO_1317 (O_1317,N_15748,N_15499);
nor UO_1318 (O_1318,N_16517,N_16602);
nand UO_1319 (O_1319,N_16549,N_18305);
xor UO_1320 (O_1320,N_16279,N_15386);
and UO_1321 (O_1321,N_17945,N_16991);
and UO_1322 (O_1322,N_15241,N_18809);
or UO_1323 (O_1323,N_19799,N_18852);
or UO_1324 (O_1324,N_15740,N_15571);
xnor UO_1325 (O_1325,N_16307,N_17719);
xor UO_1326 (O_1326,N_16068,N_15794);
and UO_1327 (O_1327,N_16025,N_19110);
xnor UO_1328 (O_1328,N_15556,N_19425);
nand UO_1329 (O_1329,N_16682,N_16091);
and UO_1330 (O_1330,N_19362,N_18151);
nor UO_1331 (O_1331,N_16451,N_19980);
and UO_1332 (O_1332,N_19684,N_18175);
xor UO_1333 (O_1333,N_19729,N_18435);
xnor UO_1334 (O_1334,N_16726,N_16519);
nand UO_1335 (O_1335,N_19715,N_18020);
nor UO_1336 (O_1336,N_19995,N_17787);
and UO_1337 (O_1337,N_15647,N_16367);
nand UO_1338 (O_1338,N_15818,N_19159);
nand UO_1339 (O_1339,N_18732,N_19280);
and UO_1340 (O_1340,N_17031,N_15799);
nor UO_1341 (O_1341,N_19657,N_16229);
nand UO_1342 (O_1342,N_19622,N_15820);
nor UO_1343 (O_1343,N_17723,N_19726);
and UO_1344 (O_1344,N_17681,N_19585);
xnor UO_1345 (O_1345,N_19178,N_18119);
and UO_1346 (O_1346,N_19936,N_17919);
nand UO_1347 (O_1347,N_15978,N_18095);
or UO_1348 (O_1348,N_16851,N_17827);
xnor UO_1349 (O_1349,N_15272,N_19784);
nand UO_1350 (O_1350,N_16777,N_15397);
and UO_1351 (O_1351,N_17846,N_18252);
or UO_1352 (O_1352,N_19452,N_16346);
or UO_1353 (O_1353,N_16166,N_18583);
nand UO_1354 (O_1354,N_18057,N_15426);
xnor UO_1355 (O_1355,N_19154,N_19494);
nand UO_1356 (O_1356,N_16280,N_19495);
and UO_1357 (O_1357,N_18430,N_17657);
or UO_1358 (O_1358,N_19389,N_18112);
nand UO_1359 (O_1359,N_18526,N_15945);
or UO_1360 (O_1360,N_16818,N_18278);
and UO_1361 (O_1361,N_17109,N_19675);
nand UO_1362 (O_1362,N_19885,N_16164);
or UO_1363 (O_1363,N_18745,N_15603);
and UO_1364 (O_1364,N_19853,N_16136);
xnor UO_1365 (O_1365,N_17870,N_18361);
nor UO_1366 (O_1366,N_18388,N_18285);
and UO_1367 (O_1367,N_15652,N_18044);
xnor UO_1368 (O_1368,N_15893,N_19323);
nand UO_1369 (O_1369,N_18066,N_18234);
or UO_1370 (O_1370,N_16294,N_19472);
and UO_1371 (O_1371,N_19671,N_16703);
xor UO_1372 (O_1372,N_19708,N_18083);
nand UO_1373 (O_1373,N_18879,N_18281);
nor UO_1374 (O_1374,N_16548,N_19886);
or UO_1375 (O_1375,N_17063,N_17364);
nand UO_1376 (O_1376,N_19176,N_16619);
or UO_1377 (O_1377,N_15975,N_15643);
nor UO_1378 (O_1378,N_15878,N_15977);
nand UO_1379 (O_1379,N_16380,N_16357);
xor UO_1380 (O_1380,N_17783,N_16165);
nor UO_1381 (O_1381,N_17371,N_16741);
nor UO_1382 (O_1382,N_17648,N_17659);
or UO_1383 (O_1383,N_18570,N_19276);
xnor UO_1384 (O_1384,N_16529,N_17683);
and UO_1385 (O_1385,N_18174,N_16447);
nor UO_1386 (O_1386,N_15403,N_17046);
or UO_1387 (O_1387,N_17760,N_18788);
xnor UO_1388 (O_1388,N_18621,N_17435);
or UO_1389 (O_1389,N_15172,N_18697);
or UO_1390 (O_1390,N_19835,N_15648);
and UO_1391 (O_1391,N_18089,N_19077);
nand UO_1392 (O_1392,N_18074,N_18548);
nand UO_1393 (O_1393,N_17219,N_17644);
and UO_1394 (O_1394,N_15789,N_16445);
nor UO_1395 (O_1395,N_16467,N_15268);
and UO_1396 (O_1396,N_15472,N_18994);
nor UO_1397 (O_1397,N_19910,N_15553);
and UO_1398 (O_1398,N_15687,N_17573);
or UO_1399 (O_1399,N_15620,N_17762);
or UO_1400 (O_1400,N_15986,N_16050);
and UO_1401 (O_1401,N_16814,N_16109);
nor UO_1402 (O_1402,N_17417,N_19660);
xnor UO_1403 (O_1403,N_19212,N_18850);
nor UO_1404 (O_1404,N_17237,N_18265);
and UO_1405 (O_1405,N_18325,N_17269);
nor UO_1406 (O_1406,N_18130,N_19263);
or UO_1407 (O_1407,N_17194,N_15215);
nand UO_1408 (O_1408,N_18613,N_17423);
nor UO_1409 (O_1409,N_15270,N_17108);
nand UO_1410 (O_1410,N_19857,N_15221);
xnor UO_1411 (O_1411,N_15308,N_17887);
xnor UO_1412 (O_1412,N_19960,N_18028);
and UO_1413 (O_1413,N_15724,N_18554);
nor UO_1414 (O_1414,N_18385,N_17967);
or UO_1415 (O_1415,N_17446,N_16250);
or UO_1416 (O_1416,N_15757,N_16181);
or UO_1417 (O_1417,N_18713,N_15412);
and UO_1418 (O_1418,N_15837,N_17087);
and UO_1419 (O_1419,N_17590,N_16049);
nor UO_1420 (O_1420,N_15352,N_17240);
or UO_1421 (O_1421,N_19305,N_18004);
nand UO_1422 (O_1422,N_18301,N_16567);
nand UO_1423 (O_1423,N_15997,N_16374);
and UO_1424 (O_1424,N_18647,N_16251);
nand UO_1425 (O_1425,N_19390,N_17819);
or UO_1426 (O_1426,N_19074,N_18340);
and UO_1427 (O_1427,N_18946,N_17442);
and UO_1428 (O_1428,N_15512,N_16985);
xor UO_1429 (O_1429,N_19558,N_17820);
and UO_1430 (O_1430,N_16663,N_19444);
xnor UO_1431 (O_1431,N_18976,N_17487);
and UO_1432 (O_1432,N_17151,N_15217);
nor UO_1433 (O_1433,N_16286,N_17168);
and UO_1434 (O_1434,N_16681,N_18091);
nand UO_1435 (O_1435,N_15164,N_17122);
nand UO_1436 (O_1436,N_19713,N_19707);
or UO_1437 (O_1437,N_19610,N_19752);
nor UO_1438 (O_1438,N_18528,N_18874);
xor UO_1439 (O_1439,N_15056,N_15140);
xnor UO_1440 (O_1440,N_17032,N_15081);
and UO_1441 (O_1441,N_15733,N_16836);
or UO_1442 (O_1442,N_15171,N_18937);
nand UO_1443 (O_1443,N_17052,N_16009);
nor UO_1444 (O_1444,N_15212,N_19050);
nand UO_1445 (O_1445,N_19211,N_16287);
or UO_1446 (O_1446,N_15416,N_15612);
and UO_1447 (O_1447,N_19224,N_15901);
nand UO_1448 (O_1448,N_15429,N_18104);
nor UO_1449 (O_1449,N_19288,N_18589);
nor UO_1450 (O_1450,N_15347,N_19776);
xor UO_1451 (O_1451,N_18557,N_18860);
xor UO_1452 (O_1452,N_15894,N_17759);
or UO_1453 (O_1453,N_15996,N_18577);
and UO_1454 (O_1454,N_15137,N_18815);
nor UO_1455 (O_1455,N_15796,N_19840);
or UO_1456 (O_1456,N_17672,N_15919);
nor UO_1457 (O_1457,N_16397,N_19592);
nand UO_1458 (O_1458,N_16265,N_19556);
or UO_1459 (O_1459,N_16075,N_16965);
and UO_1460 (O_1460,N_19257,N_15946);
or UO_1461 (O_1461,N_15800,N_18455);
nor UO_1462 (O_1462,N_17273,N_17453);
or UO_1463 (O_1463,N_17784,N_19283);
or UO_1464 (O_1464,N_17934,N_16784);
and UO_1465 (O_1465,N_15848,N_17634);
nor UO_1466 (O_1466,N_17859,N_15496);
xnor UO_1467 (O_1467,N_19643,N_19462);
xor UO_1468 (O_1468,N_15683,N_19142);
and UO_1469 (O_1469,N_15500,N_19539);
or UO_1470 (O_1470,N_16470,N_19059);
nand UO_1471 (O_1471,N_17996,N_15661);
nand UO_1472 (O_1472,N_15341,N_18086);
or UO_1473 (O_1473,N_19837,N_15899);
xor UO_1474 (O_1474,N_17613,N_19324);
and UO_1475 (O_1475,N_17213,N_19952);
and UO_1476 (O_1476,N_15948,N_17009);
nor UO_1477 (O_1477,N_18610,N_15552);
nand UO_1478 (O_1478,N_17309,N_16832);
or UO_1479 (O_1479,N_17697,N_17438);
xnor UO_1480 (O_1480,N_15638,N_18681);
nand UO_1481 (O_1481,N_15322,N_18551);
nand UO_1482 (O_1482,N_16670,N_15259);
nand UO_1483 (O_1483,N_18675,N_18356);
nand UO_1484 (O_1484,N_15665,N_17722);
nand UO_1485 (O_1485,N_18849,N_19754);
and UO_1486 (O_1486,N_18352,N_16208);
nor UO_1487 (O_1487,N_18527,N_16433);
and UO_1488 (O_1488,N_19458,N_17241);
and UO_1489 (O_1489,N_19542,N_16477);
xnor UO_1490 (O_1490,N_18573,N_15503);
and UO_1491 (O_1491,N_16095,N_16320);
xor UO_1492 (O_1492,N_17575,N_15467);
or UO_1493 (O_1493,N_19522,N_19694);
nor UO_1494 (O_1494,N_16173,N_16059);
nand UO_1495 (O_1495,N_16420,N_17885);
xor UO_1496 (O_1496,N_18351,N_15835);
or UO_1497 (O_1497,N_19939,N_17445);
nand UO_1498 (O_1498,N_16435,N_19734);
nor UO_1499 (O_1499,N_18715,N_19699);
or UO_1500 (O_1500,N_18261,N_16089);
nor UO_1501 (O_1501,N_18530,N_17197);
or UO_1502 (O_1502,N_16754,N_18397);
or UO_1503 (O_1503,N_18232,N_16057);
or UO_1504 (O_1504,N_17704,N_17220);
or UO_1505 (O_1505,N_17061,N_17767);
nand UO_1506 (O_1506,N_15357,N_18789);
and UO_1507 (O_1507,N_17257,N_16062);
xor UO_1508 (O_1508,N_18897,N_18475);
or UO_1509 (O_1509,N_16535,N_18844);
or UO_1510 (O_1510,N_15495,N_16124);
and UO_1511 (O_1511,N_19733,N_17532);
nor UO_1512 (O_1512,N_18505,N_16046);
nor UO_1513 (O_1513,N_16107,N_18978);
and UO_1514 (O_1514,N_17114,N_16353);
nand UO_1515 (O_1515,N_15405,N_19906);
or UO_1516 (O_1516,N_15437,N_17798);
nor UO_1517 (O_1517,N_15574,N_19935);
or UO_1518 (O_1518,N_19887,N_17766);
nor UO_1519 (O_1519,N_19637,N_15159);
or UO_1520 (O_1520,N_19062,N_16113);
nand UO_1521 (O_1521,N_16071,N_16369);
and UO_1522 (O_1522,N_19993,N_18001);
or UO_1523 (O_1523,N_19218,N_19587);
or UO_1524 (O_1524,N_16874,N_17831);
or UO_1525 (O_1525,N_16993,N_15815);
nor UO_1526 (O_1526,N_15684,N_16717);
and UO_1527 (O_1527,N_19379,N_19816);
or UO_1528 (O_1528,N_17869,N_15376);
nor UO_1529 (O_1529,N_17986,N_15596);
nor UO_1530 (O_1530,N_19696,N_19804);
and UO_1531 (O_1531,N_17339,N_17208);
nor UO_1532 (O_1532,N_19264,N_17298);
or UO_1533 (O_1533,N_18942,N_19552);
and UO_1534 (O_1534,N_15963,N_16422);
and UO_1535 (O_1535,N_17354,N_17616);
nor UO_1536 (O_1536,N_15501,N_16039);
xnor UO_1537 (O_1537,N_18030,N_15669);
xor UO_1538 (O_1538,N_17209,N_15243);
nand UO_1539 (O_1539,N_17367,N_19104);
or UO_1540 (O_1540,N_19790,N_15569);
nor UO_1541 (O_1541,N_17042,N_17533);
nor UO_1542 (O_1542,N_16913,N_19931);
xnor UO_1543 (O_1543,N_19038,N_18690);
xnor UO_1544 (O_1544,N_15149,N_15635);
and UO_1545 (O_1545,N_18434,N_17250);
xnor UO_1546 (O_1546,N_19717,N_19239);
and UO_1547 (O_1547,N_19073,N_15202);
or UO_1548 (O_1548,N_16984,N_15798);
and UO_1549 (O_1549,N_19096,N_19229);
xnor UO_1550 (O_1550,N_16016,N_19818);
nor UO_1551 (O_1551,N_19908,N_17743);
xnor UO_1552 (O_1552,N_16632,N_18922);
nor UO_1553 (O_1553,N_16366,N_15810);
or UO_1554 (O_1554,N_18757,N_15769);
and UO_1555 (O_1555,N_16408,N_19230);
nand UO_1556 (O_1556,N_17586,N_17977);
nand UO_1557 (O_1557,N_17664,N_16635);
nor UO_1558 (O_1558,N_15629,N_18866);
nand UO_1559 (O_1559,N_15979,N_18896);
nor UO_1560 (O_1560,N_19371,N_18241);
nand UO_1561 (O_1561,N_15857,N_16108);
and UO_1562 (O_1562,N_18590,N_17801);
xnor UO_1563 (O_1563,N_18040,N_18679);
or UO_1564 (O_1564,N_19911,N_15924);
nor UO_1565 (O_1565,N_16937,N_15872);
or UO_1566 (O_1566,N_15278,N_15004);
or UO_1567 (O_1567,N_17018,N_18134);
or UO_1568 (O_1568,N_15381,N_16563);
or UO_1569 (O_1569,N_19185,N_19978);
nor UO_1570 (O_1570,N_15248,N_19559);
or UO_1571 (O_1571,N_18288,N_15008);
nand UO_1572 (O_1572,N_15575,N_18298);
nand UO_1573 (O_1573,N_15696,N_15440);
nand UO_1574 (O_1574,N_16464,N_16953);
nand UO_1575 (O_1575,N_17834,N_16258);
and UO_1576 (O_1576,N_16055,N_18462);
nand UO_1577 (O_1577,N_15558,N_15127);
nand UO_1578 (O_1578,N_19015,N_17428);
xor UO_1579 (O_1579,N_16634,N_19493);
and UO_1580 (O_1580,N_15792,N_17617);
xor UO_1581 (O_1581,N_19313,N_19962);
xnor UO_1582 (O_1582,N_15521,N_18510);
nor UO_1583 (O_1583,N_16375,N_18837);
nand UO_1584 (O_1584,N_16540,N_18321);
nor UO_1585 (O_1585,N_15929,N_18145);
nand UO_1586 (O_1586,N_19868,N_15826);
and UO_1587 (O_1587,N_17010,N_16779);
and UO_1588 (O_1588,N_15767,N_19485);
nor UO_1589 (O_1589,N_17913,N_15642);
nor UO_1590 (O_1590,N_15967,N_15285);
or UO_1591 (O_1591,N_15066,N_17650);
nor UO_1592 (O_1592,N_16763,N_19235);
or UO_1593 (O_1593,N_18779,N_19506);
xnor UO_1594 (O_1594,N_18164,N_19826);
nand UO_1595 (O_1595,N_16970,N_18829);
or UO_1596 (O_1596,N_17306,N_16295);
nor UO_1597 (O_1597,N_18243,N_17917);
nand UO_1598 (O_1598,N_18531,N_16476);
or UO_1599 (O_1599,N_19964,N_18859);
nand UO_1600 (O_1600,N_18013,N_18023);
nand UO_1601 (O_1601,N_17099,N_19475);
nand UO_1602 (O_1602,N_16239,N_15065);
and UO_1603 (O_1603,N_15294,N_18233);
or UO_1604 (O_1604,N_16264,N_18115);
nand UO_1605 (O_1605,N_15890,N_18608);
xor UO_1606 (O_1606,N_19574,N_17667);
nor UO_1607 (O_1607,N_17685,N_16805);
nand UO_1608 (O_1608,N_16273,N_19794);
or UO_1609 (O_1609,N_17983,N_16962);
nor UO_1610 (O_1610,N_18894,N_19376);
xnor UO_1611 (O_1611,N_16792,N_15219);
or UO_1612 (O_1612,N_15562,N_15984);
nor UO_1613 (O_1613,N_17131,N_19459);
nor UO_1614 (O_1614,N_15486,N_15564);
or UO_1615 (O_1615,N_19268,N_15507);
and UO_1616 (O_1616,N_17710,N_19198);
nand UO_1617 (O_1617,N_18807,N_17795);
nand UO_1618 (O_1618,N_19957,N_17202);
and UO_1619 (O_1619,N_17134,N_19463);
xnor UO_1620 (O_1620,N_17378,N_16687);
nor UO_1621 (O_1621,N_19319,N_17075);
and UO_1622 (O_1622,N_19982,N_16030);
and UO_1623 (O_1623,N_16267,N_17287);
xor UO_1624 (O_1624,N_18696,N_19987);
nor UO_1625 (O_1625,N_18186,N_19407);
or UO_1626 (O_1626,N_19760,N_17735);
xor UO_1627 (O_1627,N_18876,N_16938);
or UO_1628 (O_1628,N_16861,N_15976);
nor UO_1629 (O_1629,N_16954,N_16322);
or UO_1630 (O_1630,N_16383,N_16680);
nand UO_1631 (O_1631,N_16666,N_15811);
nand UO_1632 (O_1632,N_15383,N_18695);
and UO_1633 (O_1633,N_19600,N_17551);
and UO_1634 (O_1634,N_19258,N_19631);
or UO_1635 (O_1635,N_18661,N_17192);
xnor UO_1636 (O_1636,N_16224,N_15694);
nand UO_1637 (O_1637,N_19331,N_16499);
xor UO_1638 (O_1638,N_18957,N_16261);
xnor UO_1639 (O_1639,N_15134,N_16986);
nand UO_1640 (O_1640,N_15864,N_16462);
xor UO_1641 (O_1641,N_18328,N_19786);
nand UO_1642 (O_1642,N_19332,N_16158);
nand UO_1643 (O_1643,N_15019,N_15295);
or UO_1644 (O_1644,N_19435,N_18888);
and UO_1645 (O_1645,N_17436,N_16331);
and UO_1646 (O_1646,N_18307,N_19650);
xor UO_1647 (O_1647,N_17652,N_16291);
xnor UO_1648 (O_1648,N_16033,N_18529);
nand UO_1649 (O_1649,N_17352,N_18207);
or UO_1650 (O_1650,N_15898,N_17691);
nand UO_1651 (O_1651,N_16246,N_16539);
nor UO_1652 (O_1652,N_18945,N_16760);
and UO_1653 (O_1653,N_15947,N_16417);
nor UO_1654 (O_1654,N_19689,N_16578);
xnor UO_1655 (O_1655,N_15304,N_19068);
nor UO_1656 (O_1656,N_15413,N_15943);
xor UO_1657 (O_1657,N_15658,N_15969);
xor UO_1658 (O_1658,N_19812,N_19291);
xnor UO_1659 (O_1659,N_15224,N_16198);
nand UO_1660 (O_1660,N_19691,N_17495);
or UO_1661 (O_1661,N_19731,N_18790);
or UO_1662 (O_1662,N_17556,N_17830);
or UO_1663 (O_1663,N_15485,N_18588);
or UO_1664 (O_1664,N_16423,N_18667);
nor UO_1665 (O_1665,N_17876,N_17764);
and UO_1666 (O_1666,N_17660,N_19525);
or UO_1667 (O_1667,N_17062,N_15328);
xor UO_1668 (O_1668,N_17754,N_17096);
nand UO_1669 (O_1669,N_19195,N_19339);
xnor UO_1670 (O_1670,N_17408,N_19397);
xor UO_1671 (O_1671,N_19971,N_19479);
xnor UO_1672 (O_1672,N_15239,N_16038);
and UO_1673 (O_1673,N_17612,N_18544);
nor UO_1674 (O_1674,N_16209,N_15922);
xnor UO_1675 (O_1675,N_18179,N_18364);
nand UO_1676 (O_1676,N_17499,N_19309);
nand UO_1677 (O_1677,N_17537,N_15968);
or UO_1678 (O_1678,N_17385,N_16073);
xnor UO_1679 (O_1679,N_19820,N_17315);
xnor UO_1680 (O_1680,N_15958,N_15402);
and UO_1681 (O_1681,N_18932,N_17511);
xnor UO_1682 (O_1682,N_16816,N_19582);
and UO_1683 (O_1683,N_15373,N_19270);
and UO_1684 (O_1684,N_16469,N_19787);
or UO_1685 (O_1685,N_19221,N_17160);
or UO_1686 (O_1686,N_18981,N_15155);
nand UO_1687 (O_1687,N_17655,N_16742);
or UO_1688 (O_1688,N_16843,N_15584);
xor UO_1689 (O_1689,N_16897,N_15194);
nor UO_1690 (O_1690,N_19924,N_19031);
xor UO_1691 (O_1691,N_19174,N_18447);
xnor UO_1692 (O_1692,N_16456,N_17592);
or UO_1693 (O_1693,N_16886,N_19183);
xor UO_1694 (O_1694,N_17778,N_19624);
xor UO_1695 (O_1695,N_16630,N_18124);
or UO_1696 (O_1696,N_18486,N_17369);
nor UO_1697 (O_1697,N_18716,N_16283);
and UO_1698 (O_1698,N_17376,N_17794);
nand UO_1699 (O_1699,N_18685,N_16933);
and UO_1700 (O_1700,N_15015,N_18532);
or UO_1701 (O_1701,N_15942,N_16618);
xor UO_1702 (O_1702,N_15238,N_18775);
nand UO_1703 (O_1703,N_19922,N_19418);
xnor UO_1704 (O_1704,N_16192,N_19087);
or UO_1705 (O_1705,N_19409,N_16781);
xnor UO_1706 (O_1706,N_16707,N_15640);
nand UO_1707 (O_1707,N_19849,N_16791);
xor UO_1708 (O_1708,N_18635,N_18481);
and UO_1709 (O_1709,N_15825,N_17070);
nor UO_1710 (O_1710,N_19879,N_18223);
xor UO_1711 (O_1711,N_16194,N_15211);
xnor UO_1712 (O_1712,N_19605,N_15725);
xor UO_1713 (O_1713,N_17965,N_17610);
nor UO_1714 (O_1714,N_18973,N_17627);
nand UO_1715 (O_1715,N_17628,N_15365);
xor UO_1716 (O_1716,N_18136,N_18955);
or UO_1717 (O_1717,N_16765,N_17918);
and UO_1718 (O_1718,N_16186,N_17574);
xnor UO_1719 (O_1719,N_17207,N_16398);
nor UO_1720 (O_1720,N_18072,N_18806);
xnor UO_1721 (O_1721,N_16262,N_19300);
nor UO_1722 (O_1722,N_17584,N_17804);
xor UO_1723 (O_1723,N_19199,N_15186);
and UO_1724 (O_1724,N_15955,N_16292);
nand UO_1725 (O_1725,N_17024,N_17638);
xor UO_1726 (O_1726,N_18899,N_17670);
xnor UO_1727 (O_1727,N_17215,N_16728);
and UO_1728 (O_1728,N_15326,N_17388);
and UO_1729 (O_1729,N_17093,N_17079);
and UO_1730 (O_1730,N_16650,N_16604);
or UO_1731 (O_1731,N_18042,N_15096);
nor UO_1732 (O_1732,N_17004,N_15732);
and UO_1733 (O_1733,N_17529,N_17788);
and UO_1734 (O_1734,N_15068,N_15868);
nand UO_1735 (O_1735,N_19363,N_19351);
and UO_1736 (O_1736,N_19255,N_17770);
or UO_1737 (O_1737,N_15324,N_19970);
xor UO_1738 (O_1738,N_15954,N_15385);
nor UO_1739 (O_1739,N_19738,N_19182);
or UO_1740 (O_1740,N_19372,N_16906);
nor UO_1741 (O_1741,N_17348,N_19688);
nand UO_1742 (O_1742,N_18293,N_18538);
nor UO_1743 (O_1743,N_18442,N_16651);
and UO_1744 (O_1744,N_16750,N_15401);
nand UO_1745 (O_1745,N_16384,N_17133);
and UO_1746 (O_1746,N_15952,N_15481);
nand UO_1747 (O_1747,N_17571,N_17694);
nor UO_1748 (O_1748,N_15907,N_16558);
xnor UO_1749 (O_1749,N_17631,N_19078);
nor UO_1750 (O_1750,N_18648,N_19811);
or UO_1751 (O_1751,N_17708,N_16720);
nor UO_1752 (O_1752,N_17726,N_16862);
xnor UO_1753 (O_1753,N_17149,N_15572);
or UO_1754 (O_1754,N_19000,N_19523);
or UO_1755 (O_1755,N_16189,N_19813);
xor UO_1756 (O_1756,N_19125,N_17199);
xnor UO_1757 (O_1757,N_19632,N_17054);
and UO_1758 (O_1758,N_19055,N_17731);
and UO_1759 (O_1759,N_19214,N_15273);
nor UO_1760 (O_1760,N_16301,N_19366);
xnor UO_1761 (O_1761,N_15985,N_19388);
xnor UO_1762 (O_1762,N_16340,N_19149);
nor UO_1763 (O_1763,N_19107,N_15616);
nor UO_1764 (O_1764,N_16371,N_16170);
and UO_1765 (O_1765,N_17098,N_17311);
or UO_1766 (O_1766,N_18691,N_15441);
or UO_1767 (O_1767,N_19695,N_19869);
and UO_1768 (O_1768,N_18126,N_17434);
or UO_1769 (O_1769,N_15067,N_17432);
and UO_1770 (O_1770,N_17687,N_16444);
nand UO_1771 (O_1771,N_15200,N_15438);
nor UO_1772 (O_1772,N_19531,N_18781);
nand UO_1773 (O_1773,N_17696,N_18350);
or UO_1774 (O_1774,N_18142,N_19026);
xnor UO_1775 (O_1775,N_17148,N_15816);
xnor UO_1776 (O_1776,N_17173,N_17294);
or UO_1777 (O_1777,N_18712,N_19861);
nand UO_1778 (O_1778,N_16226,N_16918);
nor UO_1779 (O_1779,N_18393,N_19155);
or UO_1780 (O_1780,N_17271,N_17903);
or UO_1781 (O_1781,N_18267,N_18553);
xnor UO_1782 (O_1782,N_18181,N_17469);
xnor UO_1783 (O_1783,N_16848,N_15987);
nor UO_1784 (O_1784,N_17410,N_19781);
nand UO_1785 (O_1785,N_18986,N_19275);
and UO_1786 (O_1786,N_17050,N_15052);
nand UO_1787 (O_1787,N_18012,N_15112);
or UO_1788 (O_1788,N_19172,N_18566);
nor UO_1789 (O_1789,N_15747,N_16952);
nand UO_1790 (O_1790,N_18616,N_16260);
and UO_1791 (O_1791,N_16015,N_18297);
or UO_1792 (O_1792,N_16051,N_16828);
nor UO_1793 (O_1793,N_19611,N_17621);
xnor UO_1794 (O_1794,N_18556,N_19758);
xor UO_1795 (O_1795,N_15458,N_17526);
nand UO_1796 (O_1796,N_18440,N_16240);
nor UO_1797 (O_1797,N_15530,N_19596);
xor UO_1798 (O_1798,N_18217,N_18256);
nand UO_1799 (O_1799,N_17489,N_15737);
xor UO_1800 (O_1800,N_15850,N_18484);
and UO_1801 (O_1801,N_17363,N_19066);
and UO_1802 (O_1802,N_15847,N_18521);
nand UO_1803 (O_1803,N_17599,N_19215);
xnor UO_1804 (O_1804,N_15735,N_19858);
or UO_1805 (O_1805,N_16376,N_18792);
xnor UO_1806 (O_1806,N_17429,N_19666);
nand UO_1807 (O_1807,N_15362,N_16827);
and UO_1808 (O_1808,N_18502,N_15041);
nand UO_1809 (O_1809,N_16172,N_18380);
and UO_1810 (O_1810,N_18341,N_19618);
xor UO_1811 (O_1811,N_17473,N_19374);
and UO_1812 (O_1812,N_17268,N_15511);
xnor UO_1813 (O_1813,N_16459,N_16487);
and UO_1814 (O_1814,N_19839,N_17962);
and UO_1815 (O_1815,N_16203,N_18594);
xor UO_1816 (O_1816,N_15916,N_19783);
xor UO_1817 (O_1817,N_17039,N_16054);
xnor UO_1818 (O_1818,N_15537,N_16795);
nand UO_1819 (O_1819,N_18856,N_16686);
and UO_1820 (O_1820,N_17676,N_17260);
or UO_1821 (O_1821,N_15702,N_16556);
or UO_1822 (O_1822,N_17286,N_15586);
nand UO_1823 (O_1823,N_16282,N_17393);
or UO_1824 (O_1824,N_18037,N_18541);
xor UO_1825 (O_1825,N_18599,N_17045);
and UO_1826 (O_1826,N_18572,N_17296);
and UO_1827 (O_1827,N_18392,N_17539);
xnor UO_1828 (O_1828,N_18161,N_16372);
or UO_1829 (O_1829,N_19998,N_16329);
xnor UO_1830 (O_1830,N_15266,N_19426);
or UO_1831 (O_1831,N_15071,N_15161);
nor UO_1832 (O_1832,N_16053,N_17679);
nand UO_1833 (O_1833,N_19315,N_16534);
nand UO_1834 (O_1834,N_15926,N_15010);
xor UO_1835 (O_1835,N_17012,N_15394);
or UO_1836 (O_1836,N_15606,N_15087);
or UO_1837 (O_1837,N_16505,N_19501);
and UO_1838 (O_1838,N_16799,N_17053);
xor UO_1839 (O_1839,N_16225,N_15846);
or UO_1840 (O_1840,N_17020,N_17629);
xnor UO_1841 (O_1841,N_17700,N_18927);
nor UO_1842 (O_1842,N_15263,N_19548);
nand UO_1843 (O_1843,N_19213,N_16506);
xnor UO_1844 (O_1844,N_18485,N_18079);
nand UO_1845 (O_1845,N_15776,N_18915);
or UO_1846 (O_1846,N_18022,N_16077);
xnor UO_1847 (O_1847,N_17646,N_15655);
nand UO_1848 (O_1848,N_16601,N_15117);
xnor UO_1849 (O_1849,N_17083,N_16600);
or UO_1850 (O_1850,N_19386,N_16311);
xnor UO_1851 (O_1851,N_18575,N_18172);
nand UO_1852 (O_1852,N_16212,N_16221);
and UO_1853 (O_1853,N_17245,N_17818);
nand UO_1854 (O_1854,N_15072,N_18593);
or UO_1855 (O_1855,N_19647,N_19974);
xnor UO_1856 (O_1856,N_18122,N_18120);
xor UO_1857 (O_1857,N_15003,N_19404);
or UO_1858 (O_1858,N_19986,N_17848);
or UO_1859 (O_1859,N_19333,N_15697);
nor UO_1860 (O_1860,N_16719,N_18840);
nand UO_1861 (O_1861,N_16500,N_19504);
nand UO_1862 (O_1862,N_19165,N_19284);
or UO_1863 (O_1863,N_15265,N_19991);
nor UO_1864 (O_1864,N_16338,N_19877);
and UO_1865 (O_1865,N_18169,N_19981);
nor UO_1866 (O_1866,N_18303,N_18317);
xnor UO_1867 (O_1867,N_17995,N_16466);
xnor UO_1868 (O_1868,N_15292,N_19097);
nor UO_1869 (O_1869,N_15626,N_18399);
nor UO_1870 (O_1870,N_19866,N_17021);
nor UO_1871 (O_1871,N_15966,N_18027);
nor UO_1872 (O_1872,N_16244,N_17753);
nand UO_1873 (O_1873,N_15817,N_15681);
nand UO_1874 (O_1874,N_19714,N_18749);
or UO_1875 (O_1875,N_19141,N_18997);
nor UO_1876 (O_1876,N_18839,N_19497);
nand UO_1877 (O_1877,N_16512,N_15630);
or UO_1878 (O_1878,N_19604,N_18763);
nand UO_1879 (O_1879,N_17921,N_16358);
or UO_1880 (O_1880,N_19100,N_17958);
nand UO_1881 (O_1881,N_19271,N_18211);
xnor UO_1882 (O_1882,N_15940,N_16568);
nand UO_1883 (O_1883,N_18907,N_17868);
or UO_1884 (O_1884,N_19555,N_16495);
nand UO_1885 (O_1885,N_18405,N_17301);
nor UO_1886 (O_1886,N_19400,N_15125);
nor UO_1887 (O_1887,N_17115,N_16571);
xor UO_1888 (O_1888,N_19422,N_17389);
and UO_1889 (O_1889,N_19512,N_19838);
or UO_1890 (O_1890,N_17295,N_15459);
xnor UO_1891 (O_1891,N_15279,N_19979);
xor UO_1892 (O_1892,N_16310,N_16330);
or UO_1893 (O_1893,N_16490,N_17729);
and UO_1894 (O_1894,N_15059,N_16732);
xor UO_1895 (O_1895,N_15889,N_19219);
or UO_1896 (O_1896,N_15264,N_17684);
xnor UO_1897 (O_1897,N_19716,N_19950);
and UO_1898 (O_1898,N_18674,N_18420);
nand UO_1899 (O_1899,N_15722,N_16351);
nand UO_1900 (O_1900,N_15844,N_17089);
nand UO_1901 (O_1901,N_17961,N_19403);
nor UO_1902 (O_1902,N_15856,N_18454);
and UO_1903 (O_1903,N_19337,N_15785);
xnor UO_1904 (O_1904,N_17188,N_15262);
xnor UO_1905 (O_1905,N_19763,N_15355);
nand UO_1906 (O_1906,N_18240,N_16060);
nand UO_1907 (O_1907,N_18773,N_15783);
nand UO_1908 (O_1908,N_17398,N_17284);
xnor UO_1909 (O_1909,N_15745,N_16135);
or UO_1910 (O_1910,N_16058,N_17582);
xnor UO_1911 (O_1911,N_17307,N_19777);
or UO_1912 (O_1912,N_17238,N_15628);
nand UO_1913 (O_1913,N_18374,N_18871);
or UO_1914 (O_1914,N_19105,N_16699);
nand UO_1915 (O_1915,N_17546,N_16696);
nand UO_1916 (O_1916,N_19796,N_15430);
nor UO_1917 (O_1917,N_16935,N_16928);
xnor UO_1918 (O_1918,N_17368,N_16901);
nand UO_1919 (O_1919,N_17403,N_19878);
and UO_1920 (O_1920,N_19296,N_15903);
nand UO_1921 (O_1921,N_18723,N_16701);
xor UO_1922 (O_1922,N_18718,N_18290);
or UO_1923 (O_1923,N_16220,N_16323);
nor UO_1924 (O_1924,N_17124,N_17835);
nor UO_1925 (O_1925,N_18646,N_19756);
and UO_1926 (O_1926,N_17332,N_15289);
nor UO_1927 (O_1927,N_18832,N_16882);
or UO_1928 (O_1928,N_15291,N_15260);
and UO_1929 (O_1929,N_17185,N_16654);
or UO_1930 (O_1930,N_17231,N_17243);
nand UO_1931 (O_1931,N_17107,N_19467);
or UO_1932 (O_1932,N_19116,N_17686);
xnor UO_1933 (O_1933,N_18426,N_15887);
or UO_1934 (O_1934,N_16671,N_17357);
nand UO_1935 (O_1935,N_18271,N_19601);
and UO_1936 (O_1936,N_18238,N_15185);
nand UO_1937 (O_1937,N_15957,N_16079);
xor UO_1938 (O_1938,N_18928,N_16418);
nand UO_1939 (O_1939,N_15549,N_19841);
nor UO_1940 (O_1940,N_18428,N_19730);
nand UO_1941 (O_1941,N_18421,N_16613);
xnor UO_1942 (O_1942,N_17462,N_18324);
nand UO_1943 (O_1943,N_19330,N_15372);
nor UO_1944 (O_1944,N_16343,N_18755);
and UO_1945 (O_1945,N_17255,N_17614);
nand UO_1946 (O_1946,N_15531,N_17397);
xor UO_1947 (O_1947,N_16716,N_16608);
nand UO_1948 (O_1948,N_19251,N_15605);
and UO_1949 (O_1949,N_17756,N_19412);
xnor UO_1950 (O_1950,N_17275,N_18717);
or UO_1951 (O_1951,N_15318,N_18338);
or UO_1952 (O_1952,N_17957,N_15098);
or UO_1953 (O_1953,N_16678,N_18892);
and UO_1954 (O_1954,N_17553,N_16546);
or UO_1955 (O_1955,N_19683,N_19586);
xnor UO_1956 (O_1956,N_18262,N_19685);
nand UO_1957 (O_1957,N_17482,N_16895);
nand UO_1958 (O_1958,N_18867,N_17987);
and UO_1959 (O_1959,N_16352,N_15097);
nor UO_1960 (O_1960,N_17415,N_17290);
and UO_1961 (O_1961,N_16341,N_18108);
or UO_1962 (O_1962,N_17597,N_18845);
or UO_1963 (O_1963,N_15330,N_17755);
nand UO_1964 (O_1964,N_18038,N_17347);
and UO_1965 (O_1965,N_16405,N_18121);
nor UO_1966 (O_1966,N_19450,N_19192);
nor UO_1967 (O_1967,N_15423,N_17137);
xor UO_1968 (O_1968,N_17942,N_16237);
or UO_1969 (O_1969,N_18348,N_15723);
xnor UO_1970 (O_1970,N_15317,N_16807);
nand UO_1971 (O_1971,N_16197,N_17793);
nor UO_1972 (O_1972,N_17118,N_16555);
or UO_1973 (O_1973,N_18900,N_17278);
xor UO_1974 (O_1974,N_17843,N_19746);
nor UO_1975 (O_1975,N_18496,N_17002);
xor UO_1976 (O_1976,N_17825,N_17990);
nand UO_1977 (O_1977,N_17939,N_15022);
xnor UO_1978 (O_1978,N_16070,N_15006);
xor UO_1979 (O_1979,N_16783,N_16833);
nor UO_1980 (O_1980,N_18910,N_16766);
or UO_1981 (O_1981,N_19958,N_16087);
nand UO_1982 (O_1982,N_16643,N_17175);
and UO_1983 (O_1983,N_19245,N_19281);
nor UO_1984 (O_1984,N_18236,N_17805);
and UO_1985 (O_1985,N_15424,N_17866);
xnor UO_1986 (O_1986,N_17001,N_16454);
or UO_1987 (O_1987,N_15453,N_17890);
nor UO_1988 (O_1988,N_15251,N_19238);
and UO_1989 (O_1989,N_19642,N_16638);
or UO_1990 (O_1990,N_16482,N_16722);
or UO_1991 (O_1991,N_16026,N_16526);
or UO_1992 (O_1992,N_18304,N_18222);
or UO_1993 (O_1993,N_18999,N_15677);
xnor UO_1994 (O_1994,N_19033,N_18343);
xor UO_1995 (O_1995,N_15895,N_17203);
and UO_1996 (O_1996,N_17276,N_17738);
or UO_1997 (O_1997,N_18873,N_18793);
or UO_1998 (O_1998,N_16504,N_16823);
nand UO_1999 (O_1999,N_19623,N_19487);
and UO_2000 (O_2000,N_17605,N_17059);
and UO_2001 (O_2001,N_19830,N_15029);
and UO_2002 (O_2002,N_15210,N_15366);
nor UO_2003 (O_2003,N_17718,N_16610);
and UO_2004 (O_2004,N_19380,N_19498);
or UO_2005 (O_2005,N_16072,N_15378);
nand UO_2006 (O_2006,N_19299,N_18893);
and UO_2007 (O_2007,N_17333,N_16411);
and UO_2008 (O_2008,N_16214,N_17842);
nor UO_2009 (O_2009,N_19956,N_17451);
and UO_2010 (O_2010,N_18657,N_18140);
or UO_2011 (O_2011,N_17609,N_17549);
and UO_2012 (O_2012,N_19490,N_17879);
or UO_2013 (O_2013,N_19588,N_16524);
xor UO_2014 (O_2014,N_16269,N_18220);
and UO_2015 (O_2015,N_17471,N_17266);
nor UO_2016 (O_2016,N_15528,N_17607);
xnor UO_2017 (O_2017,N_18846,N_18273);
xnor UO_2018 (O_2018,N_16485,N_19037);
nor UO_2019 (O_2019,N_19602,N_18159);
and UO_2020 (O_2020,N_18953,N_19907);
nand UO_2021 (O_2021,N_18369,N_18137);
and UO_2022 (O_2022,N_17502,N_16002);
nand UO_2023 (O_2023,N_16573,N_19123);
xnor UO_2024 (O_2024,N_15704,N_18659);
and UO_2025 (O_2025,N_16607,N_18735);
and UO_2026 (O_2026,N_17748,N_16905);
xnor UO_2027 (O_2027,N_17964,N_18558);
xor UO_2028 (O_2028,N_18084,N_16412);
xor UO_2029 (O_2029,N_17195,N_17739);
nor UO_2030 (O_2030,N_18673,N_17678);
nor UO_2031 (O_2031,N_18967,N_16743);
nand UO_2032 (O_2032,N_18923,N_16093);
nand UO_2033 (O_2033,N_15051,N_15141);
xnor UO_2034 (O_2034,N_16441,N_18748);
nand UO_2035 (O_2035,N_19044,N_18431);
nand UO_2036 (O_2036,N_17736,N_18665);
nor UO_2037 (O_2037,N_16626,N_17688);
and UO_2038 (O_2038,N_19222,N_15909);
nand UO_2039 (O_2039,N_15301,N_16757);
and UO_2040 (O_2040,N_17895,N_16513);
nand UO_2041 (O_2041,N_16259,N_18212);
and UO_2042 (O_2042,N_19035,N_15396);
nand UO_2043 (O_2043,N_19515,N_17265);
or UO_2044 (O_2044,N_16334,N_17724);
nor UO_2045 (O_2045,N_19870,N_16106);
or UO_2046 (O_2046,N_18869,N_19102);
nor UO_2047 (O_2047,N_18029,N_15761);
xnor UO_2048 (O_2048,N_17769,N_17212);
and UO_2049 (O_2049,N_19020,N_19401);
and UO_2050 (O_2050,N_15832,N_18082);
and UO_2051 (O_2051,N_16596,N_17234);
or UO_2052 (O_2052,N_16200,N_17949);
and UO_2053 (O_2053,N_15543,N_18387);
nor UO_2054 (O_2054,N_16747,N_18173);
xor UO_2055 (O_2055,N_19432,N_18443);
and UO_2056 (O_2056,N_17019,N_19018);
and UO_2057 (O_2057,N_18989,N_16955);
xnor UO_2058 (O_2058,N_19052,N_16969);
and UO_2059 (O_2059,N_19428,N_15040);
nand UO_2060 (O_2060,N_16875,N_16871);
nand UO_2061 (O_2061,N_18366,N_15363);
nand UO_2062 (O_2062,N_19012,N_17712);
or UO_2063 (O_2063,N_16789,N_19577);
and UO_2064 (O_2064,N_16465,N_18197);
and UO_2065 (O_2065,N_15302,N_18103);
nand UO_2066 (O_2066,N_16018,N_15160);
nor UO_2067 (O_2067,N_17938,N_19359);
or UO_2068 (O_2068,N_18493,N_15961);
nand UO_2069 (O_2069,N_17027,N_15118);
xor UO_2070 (O_2070,N_18603,N_19208);
nor UO_2071 (O_2071,N_15250,N_15764);
and UO_2072 (O_2072,N_18342,N_18898);
and UO_2073 (O_2073,N_19394,N_19147);
nand UO_2074 (O_2074,N_15703,N_18076);
nor UO_2075 (O_2075,N_17839,N_16305);
xor UO_2076 (O_2076,N_16714,N_17591);
nor UO_2077 (O_2077,N_18818,N_19706);
xnor UO_2078 (O_2078,N_19317,N_16006);
nor UO_2079 (O_2079,N_19530,N_18650);
nand UO_2080 (O_2080,N_17331,N_18640);
xnor UO_2081 (O_2081,N_19847,N_18365);
or UO_2082 (O_2082,N_18943,N_16923);
and UO_2083 (O_2083,N_15597,N_18878);
nand UO_2084 (O_2084,N_18300,N_19599);
nand UO_2085 (O_2085,N_16074,N_16457);
nor UO_2086 (O_2086,N_15578,N_17374);
and UO_2087 (O_2087,N_19546,N_16647);
nand UO_2088 (O_2088,N_15933,N_18184);
xnor UO_2089 (O_2089,N_15282,N_18734);
nand UO_2090 (O_2090,N_15193,N_15734);
nor UO_2091 (O_2091,N_19488,N_16776);
and UO_2092 (O_2092,N_18501,N_19508);
nand UO_2093 (O_2093,N_16191,N_18312);
nand UO_2094 (O_2094,N_18511,N_17682);
and UO_2095 (O_2095,N_15109,N_19387);
nor UO_2096 (O_2096,N_17228,N_17882);
and UO_2097 (O_2097,N_15338,N_17065);
or UO_2098 (O_2098,N_19625,N_18933);
nand UO_2099 (O_2099,N_19896,N_16484);
nand UO_2100 (O_2100,N_18965,N_18487);
nand UO_2101 (O_2101,N_15568,N_18384);
nand UO_2102 (O_2102,N_17443,N_18139);
or UO_2103 (O_2103,N_18296,N_19367);
nor UO_2104 (O_2104,N_19301,N_15361);
xor UO_2105 (O_2105,N_19692,N_15936);
and UO_2106 (O_2106,N_19117,N_18877);
or UO_2107 (O_2107,N_18168,N_18231);
xor UO_2108 (O_2108,N_17891,N_15650);
xnor UO_2109 (O_2109,N_17150,N_18054);
and UO_2110 (O_2110,N_17396,N_19491);
xor UO_2111 (O_2111,N_17817,N_15536);
and UO_2112 (O_2112,N_16999,N_18708);
nor UO_2113 (O_2113,N_17060,N_17138);
or UO_2114 (O_2114,N_16520,N_16497);
xor UO_2115 (O_2115,N_16434,N_17439);
xnor UO_2116 (O_2116,N_16648,N_18833);
or UO_2117 (O_2117,N_18726,N_19112);
or UO_2118 (O_2118,N_17387,N_15526);
xor UO_2119 (O_2119,N_15970,N_17680);
nor UO_2120 (O_2120,N_18620,N_19427);
xnor UO_2121 (O_2121,N_18398,N_16840);
and UO_2122 (O_2122,N_19996,N_18870);
nor UO_2123 (O_2123,N_19591,N_18634);
xnor UO_2124 (O_2124,N_19237,N_19925);
and UO_2125 (O_2125,N_19984,N_17630);
and UO_2126 (O_2126,N_17329,N_16013);
nand UO_2127 (O_2127,N_15364,N_18047);
xnor UO_2128 (O_2128,N_18459,N_17579);
and UO_2129 (O_2129,N_17809,N_15865);
nor UO_2130 (O_2130,N_19127,N_19616);
and UO_2131 (O_2131,N_19916,N_18612);
or UO_2132 (O_2132,N_15532,N_15410);
or UO_2133 (O_2133,N_19075,N_17906);
and UO_2134 (O_2134,N_17992,N_15662);
or UO_2135 (O_2135,N_16514,N_18642);
and UO_2136 (O_2136,N_17567,N_16825);
xnor UO_2137 (O_2137,N_18741,N_15348);
nand UO_2138 (O_2138,N_17930,N_17483);
and UO_2139 (O_2139,N_19486,N_15327);
or UO_2140 (O_2140,N_17785,N_15031);
xnor UO_2141 (O_2141,N_18150,N_19132);
xnor UO_2142 (O_2142,N_17530,N_16275);
and UO_2143 (O_2143,N_17170,N_16624);
nand UO_2144 (O_2144,N_15701,N_15711);
nand UO_2145 (O_2145,N_18026,N_18199);
xor UO_2146 (O_2146,N_15092,N_18633);
nor UO_2147 (O_2147,N_17178,N_19919);
nor UO_2148 (O_2148,N_19449,N_18153);
nor UO_2149 (O_2149,N_16019,N_18853);
or UO_2150 (O_2150,N_19164,N_19767);
or UO_2151 (O_2151,N_19205,N_17097);
nand UO_2152 (O_2152,N_15062,N_18982);
nor UO_2153 (O_2153,N_18390,N_18464);
and UO_2154 (O_2154,N_18916,N_17120);
nand UO_2155 (O_2155,N_18905,N_17936);
nor UO_2156 (O_2156,N_19041,N_15715);
and UO_2157 (O_2157,N_17304,N_18090);
nor UO_2158 (O_2158,N_15990,N_19292);
xnor UO_2159 (O_2159,N_18996,N_15455);
nor UO_2160 (O_2160,N_15786,N_19951);
and UO_2161 (O_2161,N_17221,N_15309);
nand UO_2162 (O_2162,N_16138,N_18148);
nand UO_2163 (O_2163,N_19568,N_17905);
nor UO_2164 (O_2164,N_19424,N_16925);
and UO_2165 (O_2165,N_18146,N_19824);
nor UO_2166 (O_2166,N_19825,N_18441);
or UO_2167 (O_2167,N_17177,N_16365);
xnor UO_2168 (O_2168,N_19720,N_16035);
and UO_2169 (O_2169,N_17668,N_18604);
or UO_2170 (O_2170,N_16575,N_19965);
nand UO_2171 (O_2171,N_16249,N_17952);
and UO_2172 (O_2172,N_16005,N_17673);
or UO_2173 (O_2173,N_16187,N_15375);
or UO_2174 (O_2174,N_17503,N_16694);
nand UO_2175 (O_2175,N_15388,N_15609);
and UO_2176 (O_2176,N_17979,N_15862);
nor UO_2177 (O_2177,N_18449,N_17968);
nor UO_2178 (O_2178,N_18107,N_16115);
and UO_2179 (O_2179,N_16939,N_19278);
and UO_2180 (O_2180,N_19977,N_18671);
nor UO_2181 (O_2181,N_18736,N_17598);
nand UO_2182 (O_2182,N_19322,N_17143);
nor UO_2183 (O_2183,N_16532,N_18201);
xnor UO_2184 (O_2184,N_17334,N_15001);
or UO_2185 (O_2185,N_19474,N_18189);
nand UO_2186 (O_2186,N_17902,N_16152);
nand UO_2187 (O_2187,N_19250,N_18515);
nor UO_2188 (O_2188,N_18622,N_15082);
and UO_2189 (O_2189,N_18731,N_18597);
and UO_2190 (O_2190,N_16866,N_18835);
nor UO_2191 (O_2191,N_17162,N_15060);
nand UO_2192 (O_2192,N_19447,N_15513);
nor UO_2193 (O_2193,N_16238,N_17444);
and UO_2194 (O_2194,N_18936,N_17068);
and UO_2195 (O_2195,N_17966,N_17305);
and UO_2196 (O_2196,N_17034,N_19304);
nand UO_2197 (O_2197,N_18249,N_19507);
or UO_2198 (O_2198,N_17492,N_17603);
nand UO_2199 (O_2199,N_19768,N_16403);
nor UO_2200 (O_2200,N_19669,N_16092);
and UO_2201 (O_2201,N_17006,N_18660);
xor UO_2202 (O_2202,N_18689,N_19976);
xnor UO_2203 (O_2203,N_16061,N_16154);
and UO_2204 (O_2204,N_17308,N_15675);
and UO_2205 (O_2205,N_17106,N_16767);
or UO_2206 (O_2206,N_19571,N_17572);
nor UO_2207 (O_2207,N_16787,N_17342);
nand UO_2208 (O_2208,N_16067,N_18006);
or UO_2209 (O_2209,N_17602,N_19800);
nor UO_2210 (O_2210,N_18394,N_17600);
xor UO_2211 (O_2211,N_15570,N_19254);
xnor UO_2212 (O_2212,N_15360,N_16296);
nand UO_2213 (O_2213,N_16692,N_19285);
and UO_2214 (O_2214,N_16362,N_16439);
nor UO_2215 (O_2215,N_19252,N_18911);
or UO_2216 (O_2216,N_18729,N_18993);
nand UO_2217 (O_2217,N_16298,N_15484);
and UO_2218 (O_2218,N_17441,N_18848);
xnor UO_2219 (O_2219,N_16037,N_18113);
nor UO_2220 (O_2220,N_16377,N_15162);
xor UO_2221 (O_2221,N_16217,N_15287);
xnor UO_2222 (O_2222,N_15139,N_18008);
xnor UO_2223 (O_2223,N_19860,N_18854);
nor UO_2224 (O_2224,N_17456,N_16471);
xor UO_2225 (O_2225,N_16319,N_16849);
and UO_2226 (O_2226,N_16438,N_17910);
nor UO_2227 (O_2227,N_17206,N_18263);
nand UO_2228 (O_2228,N_16942,N_15247);
xnor UO_2229 (O_2229,N_18287,N_18628);
nor UO_2230 (O_2230,N_17051,N_19277);
nand UO_2231 (O_2231,N_18299,N_17593);
or UO_2232 (O_2232,N_16123,N_19759);
and UO_2233 (O_2233,N_18760,N_15135);
nor UO_2234 (O_2234,N_18337,N_17595);
nand UO_2235 (O_2235,N_19661,N_19520);
nor UO_2236 (O_2236,N_16588,N_17587);
nand UO_2237 (O_2237,N_15679,N_17915);
nor UO_2238 (O_2238,N_16161,N_19145);
xnor UO_2239 (O_2239,N_17747,N_18823);
nor UO_2240 (O_2240,N_17000,N_18033);
or UO_2241 (O_2241,N_19354,N_17709);
or UO_2242 (O_2242,N_18182,N_16580);
nand UO_2243 (O_2243,N_19135,N_15191);
nor UO_2244 (O_2244,N_16063,N_19985);
xnor UO_2245 (O_2245,N_19067,N_17015);
or UO_2246 (O_2246,N_19938,N_16674);
or UO_2247 (O_2247,N_16893,N_17299);
or UO_2248 (O_2248,N_16128,N_15368);
xnor UO_2249 (O_2249,N_16693,N_17926);
and UO_2250 (O_2250,N_17732,N_19318);
xor UO_2251 (O_2251,N_16415,N_15950);
nor UO_2252 (O_2252,N_15803,N_16773);
and UO_2253 (O_2253,N_16612,N_16748);
and UO_2254 (O_2254,N_16315,N_16523);
nand UO_2255 (O_2255,N_19414,N_16288);
and UO_2256 (O_2256,N_18005,N_15941);
nand UO_2257 (O_2257,N_16582,N_15435);
or UO_2258 (O_2258,N_18330,N_17201);
xor UO_2259 (O_2259,N_15462,N_18480);
nor UO_2260 (O_2260,N_16027,N_16964);
nor UO_2261 (O_2261,N_15398,N_18156);
and UO_2262 (O_2262,N_19136,N_17757);
and UO_2263 (O_2263,N_16382,N_17564);
nand UO_2264 (O_2264,N_18542,N_19423);
xnor UO_2265 (O_2265,N_17943,N_15853);
xor UO_2266 (O_2266,N_17893,N_17372);
nand UO_2267 (O_2267,N_19098,N_19551);
and UO_2268 (O_2268,N_15699,N_15845);
or UO_2269 (O_2269,N_17653,N_16569);
nand UO_2270 (O_2270,N_19007,N_15312);
and UO_2271 (O_2271,N_15170,N_15917);
nor UO_2272 (O_2272,N_18938,N_15203);
nor UO_2273 (O_2273,N_19076,N_19828);
xor UO_2274 (O_2274,N_16982,N_18336);
nand UO_2275 (O_2275,N_16844,N_17837);
nand UO_2276 (O_2276,N_18227,N_18468);
or UO_2277 (O_2277,N_15510,N_15083);
or UO_2278 (O_2278,N_17534,N_17844);
and UO_2279 (O_2279,N_19072,N_15672);
or UO_2280 (O_2280,N_19086,N_19744);
nor UO_2281 (O_2281,N_19306,N_16911);
and UO_2282 (O_2282,N_15843,N_18147);
and UO_2283 (O_2283,N_15516,N_19091);
nor UO_2284 (O_2284,N_15807,N_16355);
or UO_2285 (O_2285,N_19079,N_19249);
or UO_2286 (O_2286,N_18498,N_16566);
nand UO_2287 (O_2287,N_18386,N_18275);
nor UO_2288 (O_2288,N_19204,N_16544);
nor UO_2289 (O_2289,N_17362,N_16160);
nor UO_2290 (O_2290,N_16586,N_15086);
xor UO_2291 (O_2291,N_15932,N_18567);
xor UO_2292 (O_2292,N_15371,N_18875);
and UO_2293 (O_2293,N_15925,N_19798);
or UO_2294 (O_2294,N_15093,N_17147);
xnor UO_2295 (O_2295,N_15315,N_16931);
and UO_2296 (O_2296,N_16029,N_16724);
and UO_2297 (O_2297,N_18703,N_19793);
or UO_2298 (O_2298,N_17300,N_18518);
or UO_2299 (O_2299,N_15130,N_16407);
or UO_2300 (O_2300,N_19169,N_18224);
nand UO_2301 (O_2301,N_16649,N_17740);
xor UO_2302 (O_2302,N_17611,N_15115);
nand UO_2303 (O_2303,N_18333,N_17156);
and UO_2304 (O_2304,N_16894,N_15622);
and UO_2305 (O_2305,N_19460,N_18952);
nand UO_2306 (O_2306,N_18509,N_17345);
or UO_2307 (O_2307,N_15254,N_16976);
nor UO_2308 (O_2308,N_18488,N_17335);
or UO_2309 (O_2309,N_16455,N_15494);
and UO_2310 (O_2310,N_17963,N_19678);
or UO_2311 (O_2311,N_19177,N_18041);
nand UO_2312 (O_2312,N_18776,N_17523);
xor UO_2313 (O_2313,N_18694,N_18389);
or UO_2314 (O_2314,N_15790,N_18260);
and UO_2315 (O_2315,N_15705,N_17182);
or UO_2316 (O_2316,N_16429,N_18058);
or UO_2317 (O_2317,N_19649,N_18707);
or UO_2318 (O_2318,N_17013,N_19681);
nand UO_2319 (O_2319,N_15351,N_16178);
xnor UO_2320 (O_2320,N_18280,N_15912);
nor UO_2321 (O_2321,N_16481,N_19821);
nand UO_2322 (O_2322,N_19679,N_19852);
xor UO_2323 (O_2323,N_18206,N_18523);
or UO_2324 (O_2324,N_18872,N_19808);
nor UO_2325 (O_2325,N_16736,N_16920);
or UO_2326 (O_2326,N_16852,N_19377);
xor UO_2327 (O_2327,N_19646,N_16709);
xor UO_2328 (O_2328,N_19789,N_19329);
nand UO_2329 (O_2329,N_19369,N_17802);
nand UO_2330 (O_2330,N_15944,N_16394);
xnor UO_2331 (O_2331,N_17715,N_16389);
nor UO_2332 (O_2332,N_15714,N_15111);
nand UO_2333 (O_2333,N_15188,N_16017);
nand UO_2334 (O_2334,N_16675,N_15076);
xor UO_2335 (O_2335,N_16975,N_15822);
and UO_2336 (O_2336,N_17321,N_17350);
nand UO_2337 (O_2337,N_17544,N_16137);
and UO_2338 (O_2338,N_15377,N_15712);
xor UO_2339 (O_2339,N_17920,N_15693);
nand UO_2340 (O_2340,N_15333,N_16045);
nand UO_2341 (O_2341,N_18947,N_18595);
xnor UO_2342 (O_2342,N_17216,N_15208);
nor UO_2343 (O_2343,N_15189,N_19672);
and UO_2344 (O_2344,N_17873,N_16142);
xor UO_2345 (O_2345,N_17999,N_17452);
xnor UO_2346 (O_2346,N_17814,N_18368);
nor UO_2347 (O_2347,N_16318,N_16078);
xor UO_2348 (O_2348,N_16144,N_17038);
nor UO_2349 (O_2349,N_15126,N_15225);
or UO_2350 (O_2350,N_16118,N_16621);
and UO_2351 (O_2351,N_16416,N_16903);
and UO_2352 (O_2352,N_15340,N_15296);
and UO_2353 (O_2353,N_18752,N_16044);
and UO_2354 (O_2354,N_18492,N_15891);
nand UO_2355 (O_2355,N_15346,N_18353);
and UO_2356 (O_2356,N_19589,N_17884);
nor UO_2357 (O_2357,N_18985,N_16252);
nand UO_2358 (O_2358,N_19704,N_19764);
or UO_2359 (O_2359,N_15244,N_18651);
and UO_2360 (O_2360,N_19124,N_17375);
nand UO_2361 (O_2361,N_17313,N_16008);
nor UO_2362 (O_2362,N_19200,N_16545);
or UO_2363 (O_2363,N_17390,N_18383);
or UO_2364 (O_2364,N_18470,N_19668);
xnor UO_2365 (O_2365,N_16527,N_19151);
or UO_2366 (O_2366,N_16098,N_15727);
nand UO_2367 (O_2367,N_19347,N_15691);
nor UO_2368 (O_2368,N_17198,N_17806);
nor UO_2369 (O_2369,N_16219,N_15314);
and UO_2370 (O_2370,N_19553,N_16878);
or UO_2371 (O_2371,N_19576,N_18482);
nand UO_2372 (O_2372,N_16321,N_18193);
nand UO_2373 (O_2373,N_19321,N_18334);
xor UO_2374 (O_2374,N_19855,N_16564);
or UO_2375 (O_2375,N_15709,N_19802);
or UO_2376 (O_2376,N_17180,N_16022);
nor UO_2377 (O_2377,N_15710,N_15044);
xnor UO_2378 (O_2378,N_16966,N_17912);
and UO_2379 (O_2379,N_19203,N_17472);
nor UO_2380 (O_2380,N_17861,N_18935);
or UO_2381 (O_2381,N_19175,N_15960);
or UO_2382 (O_2382,N_15245,N_19477);
nor UO_2383 (O_2383,N_18750,N_16660);
nand UO_2384 (O_2384,N_15849,N_15039);
and UO_2385 (O_2385,N_16802,N_16122);
nand UO_2386 (O_2386,N_15116,N_19521);
and UO_2387 (O_2387,N_17236,N_19274);
and UO_2388 (O_2388,N_15514,N_15509);
xor UO_2389 (O_2389,N_17857,N_17016);
nor UO_2390 (O_2390,N_19051,N_15649);
or UO_2391 (O_2391,N_15518,N_16040);
nand UO_2392 (O_2392,N_17380,N_16176);
or UO_2393 (O_2393,N_15124,N_18373);
xor UO_2394 (O_2394,N_15012,N_15119);
nand UO_2395 (O_2395,N_16664,N_17855);
xnor UO_2396 (O_2396,N_18851,N_18838);
and UO_2397 (O_2397,N_16428,N_19122);
and UO_2398 (O_2398,N_18129,N_19564);
nor UO_2399 (O_2399,N_15765,N_16972);
nand UO_2400 (O_2400,N_15888,N_16230);
or UO_2401 (O_2401,N_15369,N_18720);
xnor UO_2402 (O_2402,N_19352,N_17279);
nor UO_2403 (O_2403,N_18782,N_19482);
or UO_2404 (O_2404,N_19817,N_18816);
xnor UO_2405 (O_2405,N_18913,N_16012);
and UO_2406 (O_2406,N_18834,N_19578);
xor UO_2407 (O_2407,N_16616,N_18395);
nor UO_2408 (O_2408,N_18292,N_17136);
or UO_2409 (O_2409,N_15873,N_16241);
or UO_2410 (O_2410,N_15980,N_18059);
nor UO_2411 (O_2411,N_15956,N_19580);
or UO_2412 (O_2412,N_17789,N_17336);
nor UO_2413 (O_2413,N_19635,N_15763);
xor UO_2414 (O_2414,N_17900,N_15177);
and UO_2415 (O_2415,N_19081,N_17589);
and UO_2416 (O_2416,N_19954,N_19723);
and UO_2417 (O_2417,N_19241,N_18804);
nor UO_2418 (O_2418,N_19619,N_17519);
xor UO_2419 (O_2419,N_15190,N_18412);
nor UO_2420 (O_2420,N_15359,N_15930);
or UO_2421 (O_2421,N_17849,N_15787);
and UO_2422 (O_2422,N_15566,N_18666);
nor UO_2423 (O_2423,N_15343,N_15187);
and UO_2424 (O_2424,N_19399,N_19030);
and UO_2425 (O_2425,N_18433,N_18929);
nand UO_2426 (O_2426,N_19013,N_17552);
or UO_2427 (O_2427,N_16676,N_17554);
xor UO_2428 (O_2428,N_19429,N_18209);
or UO_2429 (O_2429,N_15290,N_15038);
xor UO_2430 (O_2430,N_19992,N_16927);
and UO_2431 (O_2431,N_16245,N_15540);
and UO_2432 (O_2432,N_16644,N_17563);
nand UO_2433 (O_2433,N_17320,N_16691);
and UO_2434 (O_2434,N_16554,N_19634);
nor UO_2435 (O_2435,N_15644,N_15148);
or UO_2436 (O_2436,N_16401,N_19160);
nor UO_2437 (O_2437,N_18149,N_19413);
xnor UO_2438 (O_2438,N_15213,N_19028);
nand UO_2439 (O_2439,N_19609,N_17971);
xnor UO_2440 (O_2440,N_17864,N_19566);
nand UO_2441 (O_2441,N_15682,N_16864);
or UO_2442 (O_2442,N_15409,N_16360);
or UO_2443 (O_2443,N_16581,N_18422);
or UO_2444 (O_2444,N_16450,N_17924);
or UO_2445 (O_2445,N_19298,N_19108);
or UO_2446 (O_2446,N_16458,N_16684);
or UO_2447 (O_2447,N_17803,N_18954);
xor UO_2448 (O_2448,N_17341,N_18714);
nand UO_2449 (O_2449,N_18771,N_18106);
nand UO_2450 (O_2450,N_17522,N_17082);
and UO_2451 (O_2451,N_15771,N_15802);
or UO_2452 (O_2452,N_18099,N_19934);
and UO_2453 (O_2453,N_18995,N_16711);
nor UO_2454 (O_2454,N_18458,N_15214);
nor UO_2455 (O_2455,N_19597,N_17242);
xor UO_2456 (O_2456,N_15927,N_17956);
nor UO_2457 (O_2457,N_17577,N_17351);
or UO_2458 (O_2458,N_19959,N_15791);
and UO_2459 (O_2459,N_17960,N_17856);
xor UO_2460 (O_2460,N_15043,N_17674);
or UO_2461 (O_2461,N_16916,N_16502);
nor UO_2462 (O_2462,N_17927,N_19994);
xnor UO_2463 (O_2463,N_16257,N_18768);
and UO_2464 (O_2464,N_18272,N_16963);
or UO_2465 (O_2465,N_16121,N_16308);
nand UO_2466 (O_2466,N_17317,N_16052);
and UO_2467 (O_2467,N_16507,N_16576);
nor UO_2468 (O_2468,N_18799,N_15358);
nor UO_2469 (O_2469,N_15222,N_16171);
and UO_2470 (O_2470,N_16771,N_16967);
or UO_2471 (O_2471,N_15813,N_19503);
nand UO_2472 (O_2472,N_16065,N_17531);
nor UO_2473 (O_2473,N_17073,N_17695);
xnor UO_2474 (O_2474,N_15885,N_17277);
or UO_2475 (O_2475,N_18049,N_16706);
xor UO_2476 (O_2476,N_16368,N_16960);
nor UO_2477 (O_2477,N_17833,N_16001);
xor UO_2478 (O_2478,N_16326,N_19667);
nand UO_2479 (O_2479,N_17291,N_17675);
xnor UO_2480 (O_2480,N_19071,N_19513);
or UO_2481 (O_2481,N_18601,N_19972);
nor UO_2482 (O_2482,N_17871,N_16752);
and UO_2483 (O_2483,N_17033,N_17560);
and UO_2484 (O_2484,N_17513,N_17496);
nor UO_2485 (O_2485,N_19021,N_19234);
or UO_2486 (O_2486,N_16031,N_18051);
or UO_2487 (O_2487,N_19532,N_16735);
or UO_2488 (O_2488,N_16887,N_19194);
nand UO_2489 (O_2489,N_19411,N_17744);
and UO_2490 (O_2490,N_17765,N_17988);
nand UO_2491 (O_2491,N_16082,N_18283);
nor UO_2492 (O_2492,N_16822,N_16655);
nand UO_2493 (O_2493,N_16615,N_18320);
nor UO_2494 (O_2494,N_19289,N_16086);
and UO_2495 (O_2495,N_15460,N_15133);
nand UO_2496 (O_2496,N_18402,N_16276);
nor UO_2497 (O_2497,N_15379,N_16309);
nor UO_2498 (O_2498,N_19210,N_15033);
nor UO_2499 (O_2499,N_16120,N_17565);
endmodule