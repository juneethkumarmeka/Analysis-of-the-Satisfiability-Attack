module basic_1500_15000_2000_10_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1339,In_63);
or U1 (N_1,In_187,In_224);
and U2 (N_2,In_1095,In_1157);
nand U3 (N_3,In_1014,In_194);
and U4 (N_4,In_1202,In_1269);
nor U5 (N_5,In_11,In_381);
nand U6 (N_6,In_825,In_1230);
or U7 (N_7,In_1008,In_765);
nand U8 (N_8,In_749,In_1305);
nor U9 (N_9,In_198,In_872);
nand U10 (N_10,In_1400,In_873);
nand U11 (N_11,In_239,In_984);
and U12 (N_12,In_4,In_1160);
nor U13 (N_13,In_318,In_550);
or U14 (N_14,In_479,In_946);
or U15 (N_15,In_1030,In_513);
and U16 (N_16,In_1348,In_635);
xor U17 (N_17,In_589,In_793);
or U18 (N_18,In_1231,In_1439);
nor U19 (N_19,In_499,In_469);
and U20 (N_20,In_1488,In_837);
and U21 (N_21,In_836,In_485);
nor U22 (N_22,In_493,In_387);
nand U23 (N_23,In_1407,In_990);
and U24 (N_24,In_29,In_1153);
nor U25 (N_25,In_445,In_710);
and U26 (N_26,In_476,In_920);
and U27 (N_27,In_1066,In_129);
nor U28 (N_28,In_788,In_721);
or U29 (N_29,In_1350,In_293);
nand U30 (N_30,In_933,In_1347);
nor U31 (N_31,In_1022,In_1);
nor U32 (N_32,In_160,In_794);
and U33 (N_33,In_256,In_929);
or U34 (N_34,In_13,In_746);
or U35 (N_35,In_264,In_983);
nor U36 (N_36,In_148,In_1482);
nor U37 (N_37,In_1408,In_636);
nand U38 (N_38,In_1227,In_491);
nor U39 (N_39,In_927,In_1221);
or U40 (N_40,In_847,In_146);
nand U41 (N_41,In_972,In_1459);
nand U42 (N_42,In_1322,In_511);
nand U43 (N_43,In_848,In_1416);
and U44 (N_44,In_1360,In_1499);
xnor U45 (N_45,In_1300,In_1009);
and U46 (N_46,In_377,In_1164);
and U47 (N_47,In_599,In_1148);
nor U48 (N_48,In_422,In_1229);
nor U49 (N_49,In_608,In_383);
and U50 (N_50,In_580,In_1070);
nor U51 (N_51,In_1471,In_219);
and U52 (N_52,In_945,In_1484);
and U53 (N_53,In_596,In_1122);
or U54 (N_54,In_628,In_309);
or U55 (N_55,In_542,In_565);
nand U56 (N_56,In_1051,In_1479);
nand U57 (N_57,In_1314,In_885);
and U58 (N_58,In_986,In_1295);
nor U59 (N_59,In_881,In_1494);
nor U60 (N_60,In_680,In_228);
nand U61 (N_61,In_522,In_151);
and U62 (N_62,In_405,In_649);
nor U63 (N_63,In_335,In_312);
or U64 (N_64,In_442,In_418);
and U65 (N_65,In_529,In_296);
and U66 (N_66,In_127,In_388);
nor U67 (N_67,In_800,In_435);
nand U68 (N_68,In_1282,In_1460);
nor U69 (N_69,In_1205,In_252);
nand U70 (N_70,In_1475,In_530);
nor U71 (N_71,In_532,In_475);
or U72 (N_72,In_423,In_366);
nand U73 (N_73,In_1316,In_327);
or U74 (N_74,In_997,In_1379);
xor U75 (N_75,In_1011,In_38);
or U76 (N_76,In_582,In_704);
nor U77 (N_77,In_560,In_1065);
xor U78 (N_78,In_334,In_55);
nor U79 (N_79,In_1150,In_541);
and U80 (N_80,In_1412,In_851);
nand U81 (N_81,In_254,In_1485);
and U82 (N_82,In_618,In_1369);
xnor U83 (N_83,In_1058,In_1478);
xnor U84 (N_84,In_735,In_954);
and U85 (N_85,In_1137,In_46);
nand U86 (N_86,In_1224,In_1077);
nor U87 (N_87,In_1085,In_152);
nand U88 (N_88,In_761,In_222);
nor U89 (N_89,In_128,In_22);
or U90 (N_90,In_263,In_1220);
nor U91 (N_91,In_1055,In_557);
xnor U92 (N_92,In_226,In_1012);
nor U93 (N_93,In_44,In_340);
nor U94 (N_94,In_901,In_826);
xor U95 (N_95,In_632,In_39);
nand U96 (N_96,In_780,In_451);
or U97 (N_97,In_890,In_189);
or U98 (N_98,In_783,In_938);
nand U99 (N_99,In_785,In_1223);
or U100 (N_100,In_1114,In_463);
nor U101 (N_101,In_401,In_1127);
nand U102 (N_102,In_584,In_120);
nand U103 (N_103,In_614,In_1287);
nor U104 (N_104,In_1024,In_47);
and U105 (N_105,In_1108,In_278);
nand U106 (N_106,In_303,In_80);
or U107 (N_107,In_270,In_611);
nand U108 (N_108,In_424,In_521);
nand U109 (N_109,In_601,In_1299);
and U110 (N_110,In_115,In_645);
and U111 (N_111,In_15,In_403);
or U112 (N_112,In_292,In_17);
nor U113 (N_113,In_1234,In_1358);
and U114 (N_114,In_571,In_70);
or U115 (N_115,In_354,In_573);
nor U116 (N_116,In_79,In_980);
nor U117 (N_117,In_86,In_755);
xor U118 (N_118,In_266,In_50);
or U119 (N_119,In_1423,In_164);
and U120 (N_120,In_496,In_594);
nand U121 (N_121,In_1431,In_1464);
and U122 (N_122,In_416,In_685);
and U123 (N_123,In_767,In_536);
nor U124 (N_124,In_974,In_360);
and U125 (N_125,In_1345,In_779);
nor U126 (N_126,In_1191,In_1063);
nor U127 (N_127,In_883,In_1173);
nor U128 (N_128,In_199,In_1332);
xor U129 (N_129,In_1483,In_1477);
or U130 (N_130,In_953,In_1125);
nand U131 (N_131,In_1487,In_668);
nand U132 (N_132,In_502,In_1243);
and U133 (N_133,In_300,In_1395);
nand U134 (N_134,In_1436,In_40);
or U135 (N_135,In_99,In_1178);
nor U136 (N_136,In_770,In_915);
xnor U137 (N_137,In_458,In_588);
or U138 (N_138,In_653,In_776);
and U139 (N_139,In_478,In_695);
nand U140 (N_140,In_899,In_287);
nor U141 (N_141,In_1073,In_210);
and U142 (N_142,In_42,In_877);
or U143 (N_143,In_1255,In_930);
xnor U144 (N_144,In_505,In_169);
nand U145 (N_145,In_1158,In_654);
and U146 (N_146,In_142,In_1414);
and U147 (N_147,In_1000,In_162);
or U148 (N_148,In_639,In_936);
nand U149 (N_149,In_864,In_1213);
nor U150 (N_150,In_1007,In_871);
nand U151 (N_151,In_205,In_677);
and U152 (N_152,In_248,In_208);
xnor U153 (N_153,In_659,In_1264);
and U154 (N_154,In_790,In_740);
or U155 (N_155,In_891,In_490);
nor U156 (N_156,In_437,In_359);
or U157 (N_157,In_1249,In_1207);
xor U158 (N_158,In_1432,In_839);
nor U159 (N_159,In_1111,In_1179);
or U160 (N_160,In_170,In_261);
nor U161 (N_161,In_1028,In_339);
or U162 (N_162,In_69,In_832);
nand U163 (N_163,In_430,In_981);
xor U164 (N_164,In_525,In_323);
nand U165 (N_165,In_213,In_1336);
nor U166 (N_166,In_688,In_736);
or U167 (N_167,In_904,In_1401);
or U168 (N_168,In_682,In_906);
and U169 (N_169,In_774,In_561);
and U170 (N_170,In_308,In_365);
nor U171 (N_171,In_868,In_1309);
nor U172 (N_172,In_1270,In_657);
and U173 (N_173,In_66,In_144);
and U174 (N_174,In_979,In_968);
nor U175 (N_175,In_1088,In_414);
nand U176 (N_176,In_1391,In_138);
or U177 (N_177,In_344,In_1129);
xor U178 (N_178,In_835,In_617);
or U179 (N_179,In_1184,In_1418);
nor U180 (N_180,In_674,In_861);
nand U181 (N_181,In_235,In_1294);
nand U182 (N_182,In_577,In_275);
nor U183 (N_183,In_1161,In_919);
or U184 (N_184,In_1372,In_268);
and U185 (N_185,In_1411,In_718);
nand U186 (N_186,In_712,In_1089);
and U187 (N_187,In_1349,In_955);
nor U188 (N_188,In_28,In_1242);
and U189 (N_189,In_364,In_1200);
xnor U190 (N_190,In_516,In_111);
nor U191 (N_191,In_326,In_14);
and U192 (N_192,In_1092,In_831);
nor U193 (N_193,In_691,In_526);
nand U194 (N_194,In_158,In_1476);
nand U195 (N_195,In_285,In_876);
xor U196 (N_196,In_562,In_552);
and U197 (N_197,In_139,In_1467);
and U198 (N_198,In_886,In_465);
and U199 (N_199,In_1225,In_937);
or U200 (N_200,In_1198,In_816);
and U201 (N_201,In_174,In_1363);
nor U202 (N_202,In_612,In_259);
nand U203 (N_203,In_1327,In_247);
nor U204 (N_204,In_1399,In_1465);
nor U205 (N_205,In_301,In_1235);
or U206 (N_206,In_1116,In_1183);
nor U207 (N_207,In_1132,In_775);
nor U208 (N_208,In_1035,In_528);
or U209 (N_209,In_1434,In_333);
nand U210 (N_210,In_587,In_400);
and U211 (N_211,In_362,In_484);
xor U212 (N_212,In_1123,In_313);
or U213 (N_213,In_1274,In_398);
xor U214 (N_214,In_1244,In_568);
nor U215 (N_215,In_41,In_21);
or U216 (N_216,In_1452,In_527);
xnor U217 (N_217,In_282,In_315);
or U218 (N_218,In_1013,In_1171);
and U219 (N_219,In_1373,In_1212);
nor U220 (N_220,In_507,In_45);
nor U221 (N_221,In_1119,In_1291);
or U222 (N_222,In_329,In_842);
xor U223 (N_223,In_1480,In_1142);
nand U224 (N_224,In_1446,In_503);
and U225 (N_225,In_1260,In_820);
or U226 (N_226,In_1091,In_1107);
nand U227 (N_227,In_778,In_638);
or U228 (N_228,In_923,In_616);
or U229 (N_229,In_743,In_808);
xnor U230 (N_230,In_67,In_1146);
or U231 (N_231,In_314,In_1417);
nand U232 (N_232,In_1343,In_209);
and U233 (N_233,In_633,In_595);
nand U234 (N_234,In_730,In_299);
or U235 (N_235,In_947,In_1147);
nand U236 (N_236,In_1440,In_1068);
nor U237 (N_237,In_384,In_578);
or U238 (N_238,In_1302,In_1115);
or U239 (N_239,In_1128,In_766);
nand U240 (N_240,In_626,In_420);
nor U241 (N_241,In_1381,In_108);
and U242 (N_242,In_351,In_593);
or U243 (N_243,In_944,In_902);
or U244 (N_244,In_630,In_773);
nor U245 (N_245,In_840,In_862);
and U246 (N_246,In_1096,In_1105);
nand U247 (N_247,In_348,In_466);
and U248 (N_248,In_1017,In_1004);
nand U249 (N_249,In_1313,In_581);
nor U250 (N_250,In_870,In_1236);
and U251 (N_251,In_548,In_952);
or U252 (N_252,In_1043,In_243);
and U253 (N_253,In_1232,In_62);
or U254 (N_254,In_1080,In_821);
xor U255 (N_255,In_6,In_830);
nor U256 (N_256,In_702,In_474);
or U257 (N_257,In_1172,In_179);
and U258 (N_258,In_846,In_670);
nor U259 (N_259,In_1099,In_1187);
nor U260 (N_260,In_1023,In_716);
and U261 (N_261,In_10,In_230);
and U262 (N_262,In_723,In_998);
nand U263 (N_263,In_903,In_1090);
and U264 (N_264,In_242,In_843);
nand U265 (N_265,In_1034,In_814);
nor U266 (N_266,In_345,In_544);
xnor U267 (N_267,In_1152,In_738);
and U268 (N_268,In_921,In_892);
xnor U269 (N_269,In_698,In_439);
nand U270 (N_270,In_1273,In_1312);
nand U271 (N_271,In_24,In_739);
nand U272 (N_272,In_368,In_23);
and U273 (N_273,In_176,In_1254);
or U274 (N_274,In_487,In_1199);
nand U275 (N_275,In_1126,In_1308);
nand U276 (N_276,In_196,In_33);
xnor U277 (N_277,In_336,In_163);
xnor U278 (N_278,In_1366,In_1292);
xor U279 (N_279,In_492,In_211);
and U280 (N_280,In_520,In_687);
and U281 (N_281,In_1344,In_855);
nor U282 (N_282,In_676,In_349);
or U283 (N_283,In_385,In_71);
and U284 (N_284,In_147,In_255);
nand U285 (N_285,In_762,In_1424);
nor U286 (N_286,In_456,In_1020);
nand U287 (N_287,In_184,In_605);
nor U288 (N_288,In_1040,In_1177);
or U289 (N_289,In_1176,In_271);
nor U290 (N_290,In_415,In_926);
nor U291 (N_291,In_647,In_1419);
nand U292 (N_292,In_1293,In_324);
and U293 (N_293,In_1303,In_887);
nand U294 (N_294,In_1056,In_438);
nand U295 (N_295,In_201,In_1331);
nand U296 (N_296,In_689,In_1057);
nor U297 (N_297,In_1272,In_760);
or U298 (N_298,In_566,In_707);
and U299 (N_299,In_711,In_1250);
nor U300 (N_300,In_1259,In_473);
nor U301 (N_301,In_995,In_481);
xnor U302 (N_302,In_1044,In_1193);
or U303 (N_303,In_273,In_1289);
or U304 (N_304,In_1319,In_965);
or U305 (N_305,In_534,In_796);
nand U306 (N_306,In_104,In_1237);
nor U307 (N_307,In_898,In_1496);
xnor U308 (N_308,In_43,In_1329);
nand U309 (N_309,In_123,In_655);
and U310 (N_310,In_833,In_823);
and U311 (N_311,In_662,In_1325);
or U312 (N_312,In_191,In_515);
or U313 (N_313,In_613,In_1490);
xnor U314 (N_314,In_1239,In_480);
nor U315 (N_315,In_854,In_126);
and U316 (N_316,In_1081,In_631);
or U317 (N_317,In_155,In_924);
and U318 (N_318,In_725,In_494);
and U319 (N_319,In_1385,In_1397);
xor U320 (N_320,In_913,In_203);
or U321 (N_321,In_894,In_1267);
nand U322 (N_322,In_1386,In_245);
nor U323 (N_323,In_787,In_686);
or U324 (N_324,In_461,In_810);
and U325 (N_325,In_234,In_48);
xor U326 (N_326,In_889,In_1268);
nand U327 (N_327,In_1357,In_1498);
nor U328 (N_328,In_1222,In_856);
or U329 (N_329,In_701,In_171);
nand U330 (N_330,In_1141,In_132);
and U331 (N_331,In_575,In_512);
or U332 (N_332,In_1365,In_1247);
and U333 (N_333,In_283,In_696);
and U334 (N_334,In_124,In_260);
nand U335 (N_335,In_1405,In_975);
nor U336 (N_336,In_102,In_1032);
nor U337 (N_337,In_1435,In_753);
nand U338 (N_338,In_1083,In_748);
nor U339 (N_339,In_1075,In_341);
nor U340 (N_340,In_1362,In_1135);
nand U341 (N_341,In_134,In_1371);
nor U342 (N_342,In_1437,In_533);
or U343 (N_343,In_238,In_625);
nand U344 (N_344,In_579,In_1493);
xor U345 (N_345,In_64,In_900);
and U346 (N_346,In_713,In_897);
or U347 (N_347,In_81,In_448);
and U348 (N_348,In_1280,In_824);
and U349 (N_349,In_1087,In_849);
nor U350 (N_350,In_715,In_1252);
and U351 (N_351,In_1136,In_1233);
nand U352 (N_352,In_462,In_1185);
nand U353 (N_353,In_295,In_841);
or U354 (N_354,In_150,In_1109);
nand U355 (N_355,In_1406,In_971);
and U356 (N_356,In_1265,In_1455);
or U357 (N_357,In_1206,In_1155);
and U358 (N_358,In_1311,In_782);
nand U359 (N_359,In_1276,In_133);
nor U360 (N_360,In_629,In_1402);
nand U361 (N_361,In_253,In_747);
nor U362 (N_362,In_1466,In_699);
nor U363 (N_363,In_1163,In_346);
nor U364 (N_364,In_720,In_942);
xor U365 (N_365,In_467,In_1338);
and U366 (N_366,In_413,In_429);
xnor U367 (N_367,In_281,In_225);
or U368 (N_368,In_697,In_118);
and U369 (N_369,In_985,In_621);
or U370 (N_370,In_1415,In_1156);
nor U371 (N_371,In_646,In_183);
and U372 (N_372,In_1328,In_912);
or U373 (N_373,In_386,In_272);
nand U374 (N_374,In_306,In_220);
or U375 (N_375,In_1442,In_370);
or U376 (N_376,In_1278,In_845);
and U377 (N_377,In_352,In_172);
or U378 (N_378,In_570,In_1100);
nor U379 (N_379,In_828,In_1469);
xnor U380 (N_380,In_978,In_969);
nor U381 (N_381,In_610,In_190);
nand U382 (N_382,In_1474,In_402);
nand U383 (N_383,In_1124,In_440);
nand U384 (N_384,In_408,In_1315);
nor U385 (N_385,In_1180,In_412);
nand U386 (N_386,In_1215,In_175);
and U387 (N_387,In_989,In_1421);
xor U388 (N_388,In_1489,In_962);
or U389 (N_389,In_551,In_1006);
or U390 (N_390,In_771,In_26);
or U391 (N_391,In_258,In_893);
or U392 (N_392,In_262,In_918);
or U393 (N_393,In_731,In_1266);
and U394 (N_394,In_811,In_1053);
nor U395 (N_395,In_666,In_165);
or U396 (N_396,In_813,In_1323);
xnor U397 (N_397,In_1097,In_369);
nor U398 (N_398,In_1016,In_1304);
or U399 (N_399,In_409,In_895);
xnor U400 (N_400,In_431,In_103);
or U401 (N_401,In_879,In_182);
and U402 (N_402,In_331,In_1041);
nor U403 (N_403,In_396,In_524);
nand U404 (N_404,In_49,In_432);
nand U405 (N_405,In_569,In_733);
nor U406 (N_406,In_1262,In_931);
and U407 (N_407,In_939,In_1226);
and U408 (N_408,In_591,In_585);
nand U409 (N_409,In_83,In_768);
or U410 (N_410,In_1082,In_193);
and U411 (N_411,In_497,In_991);
and U412 (N_412,In_156,In_453);
nand U413 (N_413,In_2,In_1048);
nor U414 (N_414,In_1258,In_727);
nand U415 (N_415,In_9,In_539);
and U416 (N_416,In_135,In_1015);
nor U417 (N_417,In_1413,In_609);
or U418 (N_418,In_1340,In_1102);
or U419 (N_419,In_880,In_1382);
nand U420 (N_420,In_865,In_1420);
nor U421 (N_421,In_316,In_1067);
nand U422 (N_422,In_664,In_56);
nor U423 (N_423,In_1166,In_819);
nor U424 (N_424,In_1429,In_592);
and U425 (N_425,In_1042,In_789);
or U426 (N_426,In_1447,In_241);
nand U427 (N_427,In_192,In_495);
nor U428 (N_428,In_648,In_844);
and U429 (N_429,In_708,In_322);
nand U430 (N_430,In_1398,In_31);
and U431 (N_431,In_1072,In_700);
nand U432 (N_432,In_276,In_119);
or U433 (N_433,In_1283,In_397);
nor U434 (N_434,In_237,In_358);
xor U435 (N_435,In_393,In_231);
nor U436 (N_436,In_84,In_1342);
xnor U437 (N_437,In_286,In_973);
or U438 (N_438,In_694,In_1364);
xor U439 (N_439,In_1021,In_131);
nor U440 (N_440,In_1454,In_643);
and U441 (N_441,In_443,In_317);
xor U442 (N_442,In_874,In_204);
nor U443 (N_443,In_54,In_1121);
and U444 (N_444,In_122,In_935);
or U445 (N_445,In_297,In_330);
nor U446 (N_446,In_1039,In_197);
nand U447 (N_447,In_1195,In_1174);
or U448 (N_448,In_215,In_858);
nand U449 (N_449,In_95,In_1359);
and U450 (N_450,In_818,In_624);
or U451 (N_451,In_321,In_1346);
nand U452 (N_452,In_141,In_1390);
xor U453 (N_453,In_987,In_1403);
nor U454 (N_454,In_112,In_1106);
or U455 (N_455,In_149,In_752);
nand U456 (N_456,In_357,In_284);
and U457 (N_457,In_1219,In_1367);
xnor U458 (N_458,In_1457,In_380);
nor U459 (N_459,In_428,In_310);
or U460 (N_460,In_168,In_1433);
nor U461 (N_461,In_1410,In_53);
and U462 (N_462,In_60,In_482);
and U463 (N_463,In_1201,In_294);
or U464 (N_464,In_620,In_722);
or U465 (N_465,In_291,In_449);
and U466 (N_466,In_1443,In_185);
or U467 (N_467,In_1361,In_1441);
nor U468 (N_468,In_1049,In_555);
nor U469 (N_469,In_289,In_371);
nor U470 (N_470,In_769,In_470);
or U471 (N_471,In_20,In_556);
or U472 (N_472,In_1154,In_140);
xnor U473 (N_473,In_1481,In_89);
xor U474 (N_474,In_732,In_1209);
xnor U475 (N_475,In_367,In_1353);
and U476 (N_476,In_1059,In_173);
nand U477 (N_477,In_399,In_269);
nand U478 (N_478,In_1182,In_1246);
or U479 (N_479,In_110,In_957);
xor U480 (N_480,In_543,In_615);
xor U481 (N_481,In_1029,In_1079);
and U482 (N_482,In_642,In_1117);
or U483 (N_483,In_1165,In_1240);
nor U484 (N_484,In_756,In_510);
or U485 (N_485,In_154,In_922);
nand U486 (N_486,In_602,In_1425);
nand U487 (N_487,In_867,In_1120);
nor U488 (N_488,In_390,In_454);
nand U489 (N_489,In_501,In_663);
or U490 (N_490,In_724,In_650);
and U491 (N_491,In_791,In_1389);
and U492 (N_492,In_1326,In_389);
or U493 (N_493,In_1378,In_457);
xnor U494 (N_494,In_717,In_640);
xor U495 (N_495,In_737,In_180);
nor U496 (N_496,In_65,In_1131);
nor U497 (N_497,In_658,In_1286);
nand U498 (N_498,In_709,In_1101);
and U499 (N_499,In_434,In_279);
nand U500 (N_500,In_153,In_540);
nor U501 (N_501,In_1409,In_909);
nand U502 (N_502,In_1170,In_407);
and U503 (N_503,In_1110,In_590);
or U504 (N_504,In_107,In_1281);
and U505 (N_505,In_667,In_372);
nand U506 (N_506,In_178,In_27);
and U507 (N_507,In_742,In_1027);
nand U508 (N_508,In_671,In_1470);
xor U509 (N_509,In_1256,In_159);
or U510 (N_510,In_355,In_1388);
nor U511 (N_511,In_436,In_483);
nor U512 (N_512,In_1317,In_274);
nor U513 (N_513,In_547,In_1143);
nand U514 (N_514,In_233,In_212);
nor U515 (N_515,In_859,In_12);
and U516 (N_516,In_433,In_1306);
nor U517 (N_517,In_186,In_1098);
nor U518 (N_518,In_934,In_116);
nand U519 (N_519,In_1375,In_290);
xnor U520 (N_520,In_227,In_719);
nand U521 (N_521,In_1194,In_419);
and U522 (N_522,In_459,In_328);
or U523 (N_523,In_1061,In_757);
or U524 (N_524,In_57,In_714);
or U525 (N_525,In_574,In_1054);
and U526 (N_526,In_940,In_106);
xnor U527 (N_527,In_93,In_1140);
nor U528 (N_528,In_745,In_232);
and U529 (N_529,In_932,In_1162);
and U530 (N_530,In_5,In_679);
xor U531 (N_531,In_280,In_206);
and U532 (N_532,In_896,In_32);
and U533 (N_533,In_797,In_754);
nor U534 (N_534,In_1341,In_363);
nor U535 (N_535,In_812,In_161);
xor U536 (N_536,In_97,In_18);
xor U537 (N_537,In_337,In_1451);
or U538 (N_538,In_195,In_598);
or U539 (N_539,In_250,In_523);
xnor U540 (N_540,In_1139,In_302);
xnor U541 (N_541,In_1279,In_1472);
nor U542 (N_542,In_907,In_257);
or U543 (N_543,In_37,In_244);
or U544 (N_544,In_1393,In_1210);
or U545 (N_545,In_1321,In_804);
or U546 (N_546,In_1253,In_802);
or U547 (N_547,In_741,In_690);
or U548 (N_548,In_1052,In_838);
xor U549 (N_549,In_1078,In_411);
nand U550 (N_550,In_267,In_1495);
nand U551 (N_551,In_852,In_125);
nor U552 (N_552,In_229,In_798);
nand U553 (N_553,In_1394,In_450);
nand U554 (N_554,In_759,In_683);
nor U555 (N_555,In_1103,In_1396);
nor U556 (N_556,In_607,In_817);
xnor U557 (N_557,In_693,In_1036);
nand U558 (N_558,In_744,In_559);
or U559 (N_559,In_1251,In_207);
and U560 (N_560,In_805,In_661);
or U561 (N_561,In_1175,In_519);
nor U562 (N_562,In_1005,In_1071);
or U563 (N_563,In_882,In_982);
and U564 (N_564,In_1430,In_1086);
and U565 (N_565,In_959,In_1190);
nor U566 (N_566,In_1189,In_1428);
nand U567 (N_567,In_16,In_1370);
or U568 (N_568,In_1228,In_1438);
or U569 (N_569,In_325,In_1324);
and U570 (N_570,In_1074,In_703);
or U571 (N_571,In_1218,In_311);
nor U572 (N_572,In_113,In_1355);
or U573 (N_573,In_684,In_251);
nand U574 (N_574,In_298,In_910);
nand U575 (N_575,In_1037,In_1019);
and U576 (N_576,In_35,In_406);
xor U577 (N_577,In_999,In_1130);
and U578 (N_578,In_656,In_100);
nor U579 (N_579,In_603,In_277);
and U580 (N_580,In_1351,In_1426);
nand U581 (N_581,In_600,In_382);
nor U582 (N_582,In_137,In_509);
nand U583 (N_583,In_1296,In_446);
or U584 (N_584,In_681,In_583);
nor U585 (N_585,In_249,In_988);
or U586 (N_586,In_1307,In_217);
nor U587 (N_587,In_884,In_378);
and U588 (N_588,In_1197,In_98);
xor U589 (N_589,In_72,In_374);
or U590 (N_590,In_1463,In_606);
or U591 (N_591,In_1167,In_531);
or U592 (N_592,In_1003,In_117);
nor U593 (N_593,In_517,In_1168);
or U594 (N_594,In_426,In_644);
nor U595 (N_595,In_3,In_1045);
or U596 (N_596,In_52,In_1214);
nand U597 (N_597,In_1380,In_1138);
or U598 (N_598,In_1263,In_1196);
nor U599 (N_599,In_976,In_1076);
and U600 (N_600,In_1384,In_1444);
nand U601 (N_601,In_1377,In_563);
and U602 (N_602,In_489,In_82);
nor U603 (N_603,In_966,In_375);
nor U604 (N_604,In_669,In_361);
nor U605 (N_605,In_221,In_356);
nor U606 (N_606,In_417,In_994);
or U607 (N_607,In_1335,In_1376);
and U608 (N_608,In_223,In_74);
nand U609 (N_609,In_202,In_964);
nand U610 (N_610,In_1151,In_34);
nand U611 (N_611,In_786,In_51);
nor U612 (N_612,In_729,In_427);
or U613 (N_613,In_834,In_806);
or U614 (N_614,In_705,In_958);
and U615 (N_615,In_1320,In_96);
nand U616 (N_616,In_19,In_307);
or U617 (N_617,In_1113,In_567);
and U618 (N_618,In_950,In_216);
xnor U619 (N_619,In_506,In_728);
nand U620 (N_620,In_908,In_1144);
nor U621 (N_621,In_1468,In_1337);
nand U622 (N_622,In_447,In_444);
nand U623 (N_623,In_827,In_1461);
nand U624 (N_624,In_807,In_518);
and U625 (N_625,In_218,In_1216);
nand U626 (N_626,In_1277,In_136);
and U627 (N_627,In_853,In_1288);
and U628 (N_628,In_338,In_869);
and U629 (N_629,In_92,In_1062);
nor U630 (N_630,In_343,In_1404);
or U631 (N_631,In_948,In_949);
nor U632 (N_632,In_77,In_863);
nand U633 (N_633,In_85,In_181);
or U634 (N_634,In_1064,In_675);
xnor U635 (N_635,In_1318,In_1010);
nand U636 (N_636,In_545,In_78);
nand U637 (N_637,In_7,In_1001);
or U638 (N_638,In_395,In_992);
nor U639 (N_639,In_1450,In_917);
or U640 (N_640,In_1297,In_777);
nand U641 (N_641,In_58,In_627);
nor U642 (N_642,In_815,In_36);
or U643 (N_643,In_332,In_916);
nand U644 (N_644,In_857,In_455);
nand U645 (N_645,In_236,In_860);
and U646 (N_646,In_319,In_1333);
nand U647 (N_647,In_993,In_101);
xnor U648 (N_648,In_764,In_1050);
nor U649 (N_649,In_672,In_1112);
xor U650 (N_650,In_379,In_392);
nand U651 (N_651,In_905,In_750);
nand U652 (N_652,In_734,In_866);
and U653 (N_653,In_941,In_960);
nor U654 (N_654,In_925,In_1383);
or U655 (N_655,In_809,In_59);
or U656 (N_656,In_265,In_1257);
nor U657 (N_657,In_1310,In_665);
and U658 (N_658,In_1133,In_1169);
and U659 (N_659,In_87,In_1186);
xnor U660 (N_660,In_758,In_441);
nor U661 (N_661,In_1334,In_394);
nor U662 (N_662,In_1134,In_1002);
nor U663 (N_663,In_996,In_500);
or U664 (N_664,In_145,In_486);
nand U665 (N_665,In_1453,In_1449);
nand U666 (N_666,In_1060,In_875);
or U667 (N_667,In_1188,In_1271);
nand U668 (N_668,In_1301,In_342);
nor U669 (N_669,In_1285,In_634);
nor U670 (N_670,In_967,In_1217);
nor U671 (N_671,In_726,In_498);
nor U672 (N_672,In_751,In_1181);
or U673 (N_673,In_803,In_1392);
xor U674 (N_674,In_1069,In_706);
and U675 (N_675,In_88,In_850);
and U676 (N_676,In_410,In_1486);
nor U677 (N_677,In_660,In_353);
xnor U678 (N_678,In_1033,In_1458);
nor U679 (N_679,In_576,In_1118);
nand U680 (N_680,In_376,In_977);
or U681 (N_681,In_1462,In_1145);
and U682 (N_682,In_214,In_1492);
and U683 (N_683,In_1374,In_373);
or U684 (N_684,In_792,In_477);
xor U685 (N_685,In_240,In_468);
nand U686 (N_686,In_1047,In_535);
and U687 (N_687,In_564,In_504);
xor U688 (N_688,In_1208,In_546);
xnor U689 (N_689,In_537,In_956);
nand U690 (N_690,In_304,In_829);
and U691 (N_691,In_801,In_1448);
or U692 (N_692,In_1497,In_1211);
nor U693 (N_693,In_1284,In_549);
xor U694 (N_694,In_90,In_200);
and U695 (N_695,In_763,In_784);
xor U696 (N_696,In_350,In_1352);
nor U697 (N_697,In_772,In_951);
and U698 (N_698,In_623,In_73);
and U699 (N_699,In_347,In_1368);
and U700 (N_700,In_464,In_0);
xnor U701 (N_701,In_1261,In_673);
xor U702 (N_702,In_911,In_586);
nand U703 (N_703,In_1046,In_452);
and U704 (N_704,In_1275,In_597);
and U705 (N_705,In_1025,In_114);
or U706 (N_706,In_914,In_320);
nand U707 (N_707,In_1238,In_305);
and U708 (N_708,In_75,In_288);
nor U709 (N_709,In_1422,In_94);
and U710 (N_710,In_822,In_651);
or U711 (N_711,In_472,In_943);
or U712 (N_712,In_637,In_25);
nand U713 (N_713,In_130,In_1248);
nand U714 (N_714,In_1038,In_692);
nor U715 (N_715,In_1084,In_1354);
nor U716 (N_716,In_514,In_167);
nor U717 (N_717,In_554,In_404);
and U718 (N_718,In_68,In_795);
and U719 (N_719,In_1094,In_471);
or U720 (N_720,In_1491,In_8);
nand U721 (N_721,In_888,In_1290);
nor U722 (N_722,In_1204,In_619);
nor U723 (N_723,In_1018,In_91);
nor U724 (N_724,In_1241,In_553);
and U725 (N_725,In_538,In_970);
nand U726 (N_726,In_781,In_1456);
and U727 (N_727,In_558,In_1192);
or U728 (N_728,In_604,In_961);
or U729 (N_729,In_188,In_1104);
xor U730 (N_730,In_799,In_1356);
and U731 (N_731,In_641,In_1159);
and U732 (N_732,In_157,In_1298);
and U733 (N_733,In_963,In_1203);
xor U734 (N_734,In_61,In_30);
and U735 (N_735,In_105,In_76);
or U736 (N_736,In_1427,In_391);
nand U737 (N_737,In_678,In_1473);
nor U738 (N_738,In_488,In_1093);
nor U739 (N_739,In_622,In_1026);
xor U740 (N_740,In_1031,In_109);
and U741 (N_741,In_572,In_425);
nand U742 (N_742,In_421,In_121);
and U743 (N_743,In_1245,In_1330);
or U744 (N_744,In_246,In_652);
and U745 (N_745,In_878,In_928);
or U746 (N_746,In_177,In_166);
or U747 (N_747,In_1445,In_508);
or U748 (N_748,In_460,In_1149);
or U749 (N_749,In_1387,In_143);
nor U750 (N_750,In_827,In_1111);
nand U751 (N_751,In_770,In_65);
nand U752 (N_752,In_176,In_429);
and U753 (N_753,In_1478,In_1451);
nand U754 (N_754,In_62,In_690);
nand U755 (N_755,In_395,In_973);
nor U756 (N_756,In_294,In_616);
xor U757 (N_757,In_975,In_1370);
nand U758 (N_758,In_1332,In_137);
and U759 (N_759,In_507,In_1224);
and U760 (N_760,In_999,In_79);
and U761 (N_761,In_1341,In_459);
nor U762 (N_762,In_1036,In_1420);
and U763 (N_763,In_1438,In_1050);
and U764 (N_764,In_1121,In_679);
nor U765 (N_765,In_1175,In_911);
nor U766 (N_766,In_904,In_41);
and U767 (N_767,In_1408,In_1467);
nand U768 (N_768,In_23,In_329);
xnor U769 (N_769,In_66,In_39);
or U770 (N_770,In_322,In_729);
and U771 (N_771,In_1155,In_984);
nand U772 (N_772,In_1055,In_373);
and U773 (N_773,In_742,In_1417);
or U774 (N_774,In_56,In_418);
and U775 (N_775,In_239,In_323);
or U776 (N_776,In_1225,In_672);
nor U777 (N_777,In_106,In_239);
and U778 (N_778,In_646,In_75);
nand U779 (N_779,In_479,In_632);
and U780 (N_780,In_990,In_763);
nor U781 (N_781,In_93,In_188);
or U782 (N_782,In_238,In_1313);
or U783 (N_783,In_673,In_655);
nor U784 (N_784,In_741,In_122);
nor U785 (N_785,In_400,In_1052);
or U786 (N_786,In_1441,In_341);
xor U787 (N_787,In_520,In_877);
and U788 (N_788,In_258,In_1326);
xnor U789 (N_789,In_222,In_553);
or U790 (N_790,In_1065,In_1120);
or U791 (N_791,In_704,In_710);
nor U792 (N_792,In_1016,In_449);
or U793 (N_793,In_499,In_1383);
or U794 (N_794,In_853,In_601);
and U795 (N_795,In_1470,In_165);
nand U796 (N_796,In_27,In_331);
nand U797 (N_797,In_487,In_1209);
nand U798 (N_798,In_441,In_1169);
or U799 (N_799,In_746,In_1484);
and U800 (N_800,In_213,In_438);
or U801 (N_801,In_13,In_624);
and U802 (N_802,In_1148,In_454);
and U803 (N_803,In_232,In_1344);
nor U804 (N_804,In_604,In_784);
and U805 (N_805,In_107,In_220);
nor U806 (N_806,In_962,In_790);
nand U807 (N_807,In_119,In_193);
or U808 (N_808,In_1289,In_1300);
nor U809 (N_809,In_1331,In_1386);
nor U810 (N_810,In_1482,In_0);
nor U811 (N_811,In_476,In_908);
or U812 (N_812,In_126,In_943);
and U813 (N_813,In_1098,In_1070);
or U814 (N_814,In_701,In_439);
nand U815 (N_815,In_1284,In_65);
and U816 (N_816,In_1095,In_1337);
or U817 (N_817,In_196,In_179);
or U818 (N_818,In_877,In_182);
and U819 (N_819,In_10,In_1162);
nand U820 (N_820,In_57,In_366);
nor U821 (N_821,In_1119,In_1315);
or U822 (N_822,In_1012,In_612);
or U823 (N_823,In_787,In_1128);
or U824 (N_824,In_1069,In_299);
and U825 (N_825,In_1145,In_380);
nor U826 (N_826,In_1230,In_247);
or U827 (N_827,In_655,In_766);
or U828 (N_828,In_1484,In_233);
nor U829 (N_829,In_296,In_350);
nand U830 (N_830,In_514,In_648);
nor U831 (N_831,In_947,In_379);
nand U832 (N_832,In_671,In_413);
and U833 (N_833,In_1036,In_487);
or U834 (N_834,In_398,In_1493);
xnor U835 (N_835,In_958,In_794);
nand U836 (N_836,In_236,In_302);
nand U837 (N_837,In_473,In_657);
or U838 (N_838,In_132,In_411);
and U839 (N_839,In_405,In_139);
and U840 (N_840,In_1476,In_287);
nor U841 (N_841,In_573,In_1250);
nor U842 (N_842,In_1258,In_1207);
and U843 (N_843,In_625,In_241);
nor U844 (N_844,In_1176,In_255);
and U845 (N_845,In_1462,In_1125);
or U846 (N_846,In_1271,In_1405);
nand U847 (N_847,In_306,In_1385);
nand U848 (N_848,In_391,In_860);
or U849 (N_849,In_1376,In_966);
and U850 (N_850,In_51,In_472);
nor U851 (N_851,In_1249,In_1433);
nand U852 (N_852,In_810,In_239);
and U853 (N_853,In_182,In_1302);
or U854 (N_854,In_1472,In_1003);
nor U855 (N_855,In_688,In_209);
or U856 (N_856,In_257,In_700);
or U857 (N_857,In_84,In_1472);
and U858 (N_858,In_882,In_746);
and U859 (N_859,In_1074,In_1498);
and U860 (N_860,In_686,In_1454);
and U861 (N_861,In_1445,In_651);
nand U862 (N_862,In_43,In_955);
nand U863 (N_863,In_917,In_516);
or U864 (N_864,In_345,In_1281);
nor U865 (N_865,In_392,In_1300);
or U866 (N_866,In_844,In_254);
or U867 (N_867,In_952,In_595);
nor U868 (N_868,In_1266,In_1022);
nand U869 (N_869,In_35,In_941);
or U870 (N_870,In_572,In_164);
and U871 (N_871,In_456,In_751);
nor U872 (N_872,In_963,In_613);
nand U873 (N_873,In_1106,In_425);
or U874 (N_874,In_409,In_781);
or U875 (N_875,In_291,In_936);
nor U876 (N_876,In_899,In_371);
nor U877 (N_877,In_1001,In_382);
or U878 (N_878,In_312,In_155);
or U879 (N_879,In_199,In_937);
or U880 (N_880,In_1439,In_1035);
nand U881 (N_881,In_474,In_359);
and U882 (N_882,In_307,In_255);
nand U883 (N_883,In_346,In_695);
nor U884 (N_884,In_595,In_750);
nor U885 (N_885,In_1057,In_1499);
nor U886 (N_886,In_343,In_49);
or U887 (N_887,In_1199,In_381);
nor U888 (N_888,In_1217,In_897);
nor U889 (N_889,In_284,In_821);
nand U890 (N_890,In_600,In_1275);
nand U891 (N_891,In_1472,In_314);
nor U892 (N_892,In_1133,In_787);
nor U893 (N_893,In_347,In_501);
nor U894 (N_894,In_1346,In_235);
xnor U895 (N_895,In_1395,In_284);
nand U896 (N_896,In_130,In_500);
xor U897 (N_897,In_569,In_611);
or U898 (N_898,In_1199,In_426);
nand U899 (N_899,In_204,In_567);
nor U900 (N_900,In_396,In_241);
nor U901 (N_901,In_1070,In_253);
xnor U902 (N_902,In_1015,In_303);
or U903 (N_903,In_1362,In_163);
and U904 (N_904,In_698,In_839);
and U905 (N_905,In_760,In_167);
and U906 (N_906,In_1308,In_752);
or U907 (N_907,In_38,In_649);
or U908 (N_908,In_1198,In_1034);
nor U909 (N_909,In_13,In_916);
and U910 (N_910,In_799,In_92);
and U911 (N_911,In_1457,In_882);
nor U912 (N_912,In_892,In_312);
nor U913 (N_913,In_316,In_564);
or U914 (N_914,In_73,In_807);
nand U915 (N_915,In_1014,In_463);
and U916 (N_916,In_853,In_945);
and U917 (N_917,In_372,In_774);
or U918 (N_918,In_1280,In_1374);
xor U919 (N_919,In_516,In_133);
or U920 (N_920,In_913,In_1058);
nand U921 (N_921,In_638,In_1332);
and U922 (N_922,In_82,In_519);
nand U923 (N_923,In_91,In_1491);
nand U924 (N_924,In_350,In_69);
or U925 (N_925,In_1455,In_83);
nand U926 (N_926,In_93,In_801);
nand U927 (N_927,In_214,In_971);
or U928 (N_928,In_923,In_929);
or U929 (N_929,In_803,In_922);
nor U930 (N_930,In_1216,In_938);
nand U931 (N_931,In_991,In_92);
or U932 (N_932,In_1231,In_1208);
nand U933 (N_933,In_805,In_849);
xnor U934 (N_934,In_1061,In_1282);
nand U935 (N_935,In_233,In_758);
or U936 (N_936,In_573,In_71);
or U937 (N_937,In_1281,In_380);
xor U938 (N_938,In_348,In_148);
nor U939 (N_939,In_1446,In_619);
or U940 (N_940,In_184,In_1183);
nor U941 (N_941,In_1414,In_648);
and U942 (N_942,In_1402,In_376);
or U943 (N_943,In_350,In_1134);
nor U944 (N_944,In_188,In_408);
or U945 (N_945,In_495,In_114);
nor U946 (N_946,In_1060,In_81);
nand U947 (N_947,In_1093,In_1182);
nor U948 (N_948,In_727,In_1312);
nand U949 (N_949,In_501,In_165);
nor U950 (N_950,In_441,In_202);
or U951 (N_951,In_516,In_1283);
or U952 (N_952,In_92,In_150);
or U953 (N_953,In_468,In_137);
nand U954 (N_954,In_550,In_236);
and U955 (N_955,In_383,In_94);
nor U956 (N_956,In_912,In_11);
and U957 (N_957,In_1019,In_1401);
nand U958 (N_958,In_12,In_1418);
nor U959 (N_959,In_590,In_1264);
nand U960 (N_960,In_837,In_199);
nor U961 (N_961,In_287,In_901);
and U962 (N_962,In_786,In_1085);
or U963 (N_963,In_1366,In_1043);
or U964 (N_964,In_661,In_1316);
xor U965 (N_965,In_1433,In_1169);
nand U966 (N_966,In_454,In_319);
nor U967 (N_967,In_1454,In_1414);
nand U968 (N_968,In_1250,In_1466);
or U969 (N_969,In_869,In_169);
nand U970 (N_970,In_595,In_829);
nor U971 (N_971,In_633,In_471);
and U972 (N_972,In_581,In_471);
and U973 (N_973,In_35,In_619);
nor U974 (N_974,In_503,In_1489);
nor U975 (N_975,In_1231,In_23);
and U976 (N_976,In_614,In_410);
nand U977 (N_977,In_589,In_691);
or U978 (N_978,In_1393,In_104);
xor U979 (N_979,In_1227,In_691);
or U980 (N_980,In_73,In_727);
nor U981 (N_981,In_163,In_1467);
and U982 (N_982,In_688,In_35);
or U983 (N_983,In_1465,In_617);
and U984 (N_984,In_656,In_1407);
or U985 (N_985,In_295,In_247);
xnor U986 (N_986,In_1352,In_861);
and U987 (N_987,In_1302,In_1215);
nor U988 (N_988,In_363,In_485);
nand U989 (N_989,In_410,In_345);
and U990 (N_990,In_700,In_784);
or U991 (N_991,In_1230,In_1345);
or U992 (N_992,In_70,In_534);
nand U993 (N_993,In_765,In_1223);
nor U994 (N_994,In_773,In_816);
or U995 (N_995,In_909,In_1043);
xnor U996 (N_996,In_233,In_289);
and U997 (N_997,In_1421,In_1229);
nor U998 (N_998,In_1102,In_795);
or U999 (N_999,In_38,In_448);
nor U1000 (N_1000,In_88,In_1358);
nand U1001 (N_1001,In_892,In_918);
nor U1002 (N_1002,In_803,In_35);
nand U1003 (N_1003,In_1113,In_727);
and U1004 (N_1004,In_297,In_419);
nor U1005 (N_1005,In_1055,In_247);
nor U1006 (N_1006,In_53,In_1408);
and U1007 (N_1007,In_477,In_590);
nor U1008 (N_1008,In_458,In_70);
and U1009 (N_1009,In_1250,In_110);
nand U1010 (N_1010,In_683,In_463);
xnor U1011 (N_1011,In_1448,In_923);
nor U1012 (N_1012,In_97,In_343);
nand U1013 (N_1013,In_70,In_1276);
and U1014 (N_1014,In_688,In_1112);
nor U1015 (N_1015,In_302,In_1248);
nand U1016 (N_1016,In_31,In_839);
nand U1017 (N_1017,In_1051,In_1251);
and U1018 (N_1018,In_831,In_827);
and U1019 (N_1019,In_488,In_306);
and U1020 (N_1020,In_1451,In_1177);
nand U1021 (N_1021,In_1425,In_875);
nor U1022 (N_1022,In_256,In_881);
nand U1023 (N_1023,In_183,In_1226);
nand U1024 (N_1024,In_251,In_90);
nor U1025 (N_1025,In_435,In_1231);
xnor U1026 (N_1026,In_751,In_1054);
or U1027 (N_1027,In_1171,In_259);
and U1028 (N_1028,In_715,In_758);
or U1029 (N_1029,In_1398,In_997);
or U1030 (N_1030,In_741,In_1013);
nand U1031 (N_1031,In_509,In_1409);
or U1032 (N_1032,In_1390,In_673);
xnor U1033 (N_1033,In_789,In_1339);
and U1034 (N_1034,In_312,In_1395);
nor U1035 (N_1035,In_266,In_329);
or U1036 (N_1036,In_1331,In_220);
and U1037 (N_1037,In_1259,In_1038);
and U1038 (N_1038,In_503,In_888);
and U1039 (N_1039,In_198,In_143);
xnor U1040 (N_1040,In_1482,In_1233);
nor U1041 (N_1041,In_1224,In_444);
and U1042 (N_1042,In_1350,In_442);
and U1043 (N_1043,In_1265,In_1403);
and U1044 (N_1044,In_1249,In_1160);
nand U1045 (N_1045,In_1430,In_1101);
nor U1046 (N_1046,In_145,In_548);
or U1047 (N_1047,In_1058,In_1263);
or U1048 (N_1048,In_955,In_74);
or U1049 (N_1049,In_40,In_1231);
or U1050 (N_1050,In_454,In_233);
and U1051 (N_1051,In_1335,In_806);
nand U1052 (N_1052,In_126,In_329);
or U1053 (N_1053,In_1283,In_722);
and U1054 (N_1054,In_1163,In_245);
or U1055 (N_1055,In_101,In_1283);
nor U1056 (N_1056,In_592,In_632);
and U1057 (N_1057,In_470,In_1169);
or U1058 (N_1058,In_923,In_477);
and U1059 (N_1059,In_1460,In_615);
and U1060 (N_1060,In_1170,In_49);
nand U1061 (N_1061,In_467,In_719);
or U1062 (N_1062,In_433,In_387);
or U1063 (N_1063,In_483,In_186);
and U1064 (N_1064,In_280,In_385);
nand U1065 (N_1065,In_1024,In_1376);
nor U1066 (N_1066,In_1142,In_1408);
xor U1067 (N_1067,In_76,In_266);
nor U1068 (N_1068,In_570,In_648);
nand U1069 (N_1069,In_1444,In_1026);
or U1070 (N_1070,In_149,In_920);
xor U1071 (N_1071,In_927,In_271);
nand U1072 (N_1072,In_382,In_266);
xor U1073 (N_1073,In_133,In_756);
or U1074 (N_1074,In_1043,In_1137);
and U1075 (N_1075,In_1317,In_437);
nand U1076 (N_1076,In_1125,In_1020);
or U1077 (N_1077,In_600,In_838);
nand U1078 (N_1078,In_1326,In_952);
and U1079 (N_1079,In_394,In_317);
xnor U1080 (N_1080,In_993,In_371);
and U1081 (N_1081,In_1266,In_697);
nand U1082 (N_1082,In_488,In_58);
nor U1083 (N_1083,In_1371,In_989);
xor U1084 (N_1084,In_1192,In_642);
or U1085 (N_1085,In_1420,In_859);
or U1086 (N_1086,In_780,In_131);
nor U1087 (N_1087,In_1473,In_1452);
or U1088 (N_1088,In_974,In_294);
or U1089 (N_1089,In_1106,In_706);
and U1090 (N_1090,In_869,In_254);
or U1091 (N_1091,In_706,In_355);
nand U1092 (N_1092,In_758,In_351);
and U1093 (N_1093,In_1244,In_1356);
xor U1094 (N_1094,In_36,In_1190);
and U1095 (N_1095,In_1389,In_1195);
nand U1096 (N_1096,In_457,In_1205);
nor U1097 (N_1097,In_302,In_241);
and U1098 (N_1098,In_1428,In_764);
nand U1099 (N_1099,In_362,In_118);
xnor U1100 (N_1100,In_571,In_956);
and U1101 (N_1101,In_903,In_1497);
or U1102 (N_1102,In_268,In_1138);
nor U1103 (N_1103,In_537,In_268);
nor U1104 (N_1104,In_164,In_1333);
and U1105 (N_1105,In_704,In_718);
nand U1106 (N_1106,In_681,In_1256);
nor U1107 (N_1107,In_772,In_1093);
and U1108 (N_1108,In_1391,In_369);
nand U1109 (N_1109,In_356,In_1470);
nor U1110 (N_1110,In_1167,In_950);
nor U1111 (N_1111,In_779,In_1025);
or U1112 (N_1112,In_41,In_228);
or U1113 (N_1113,In_959,In_724);
nand U1114 (N_1114,In_1446,In_206);
nand U1115 (N_1115,In_1372,In_782);
nor U1116 (N_1116,In_306,In_1210);
and U1117 (N_1117,In_1170,In_34);
and U1118 (N_1118,In_1014,In_1442);
or U1119 (N_1119,In_1047,In_1209);
xnor U1120 (N_1120,In_1230,In_384);
and U1121 (N_1121,In_1172,In_1144);
and U1122 (N_1122,In_933,In_1464);
nor U1123 (N_1123,In_460,In_1462);
xor U1124 (N_1124,In_1170,In_196);
nand U1125 (N_1125,In_407,In_892);
and U1126 (N_1126,In_126,In_10);
or U1127 (N_1127,In_1200,In_187);
nor U1128 (N_1128,In_684,In_374);
and U1129 (N_1129,In_350,In_534);
and U1130 (N_1130,In_825,In_364);
nor U1131 (N_1131,In_1487,In_907);
xnor U1132 (N_1132,In_748,In_1490);
nor U1133 (N_1133,In_830,In_1003);
or U1134 (N_1134,In_717,In_204);
and U1135 (N_1135,In_1441,In_1144);
and U1136 (N_1136,In_59,In_953);
nand U1137 (N_1137,In_466,In_1392);
xnor U1138 (N_1138,In_418,In_549);
nor U1139 (N_1139,In_444,In_1089);
nor U1140 (N_1140,In_465,In_910);
and U1141 (N_1141,In_1451,In_437);
and U1142 (N_1142,In_1405,In_605);
or U1143 (N_1143,In_435,In_948);
and U1144 (N_1144,In_932,In_712);
nand U1145 (N_1145,In_1475,In_71);
nor U1146 (N_1146,In_1016,In_42);
nor U1147 (N_1147,In_186,In_91);
nand U1148 (N_1148,In_559,In_675);
or U1149 (N_1149,In_1402,In_178);
nor U1150 (N_1150,In_824,In_1047);
nand U1151 (N_1151,In_1392,In_130);
xnor U1152 (N_1152,In_1384,In_888);
nor U1153 (N_1153,In_522,In_723);
nand U1154 (N_1154,In_860,In_909);
or U1155 (N_1155,In_857,In_170);
nand U1156 (N_1156,In_1033,In_484);
or U1157 (N_1157,In_1295,In_1456);
nor U1158 (N_1158,In_1051,In_816);
or U1159 (N_1159,In_290,In_633);
and U1160 (N_1160,In_1464,In_680);
nor U1161 (N_1161,In_176,In_63);
or U1162 (N_1162,In_1057,In_1316);
nor U1163 (N_1163,In_1320,In_25);
nor U1164 (N_1164,In_1182,In_1388);
nor U1165 (N_1165,In_931,In_1112);
or U1166 (N_1166,In_396,In_229);
nor U1167 (N_1167,In_1106,In_1031);
nor U1168 (N_1168,In_796,In_79);
nand U1169 (N_1169,In_1202,In_881);
nor U1170 (N_1170,In_82,In_1217);
or U1171 (N_1171,In_683,In_1218);
nand U1172 (N_1172,In_172,In_349);
and U1173 (N_1173,In_92,In_15);
nand U1174 (N_1174,In_729,In_174);
nand U1175 (N_1175,In_690,In_1296);
and U1176 (N_1176,In_748,In_75);
nand U1177 (N_1177,In_558,In_420);
nor U1178 (N_1178,In_885,In_247);
nor U1179 (N_1179,In_1096,In_678);
nor U1180 (N_1180,In_937,In_271);
nor U1181 (N_1181,In_620,In_20);
or U1182 (N_1182,In_191,In_967);
and U1183 (N_1183,In_1327,In_1236);
xnor U1184 (N_1184,In_1105,In_632);
xnor U1185 (N_1185,In_360,In_1084);
nor U1186 (N_1186,In_1329,In_1274);
or U1187 (N_1187,In_626,In_1459);
or U1188 (N_1188,In_107,In_1117);
xnor U1189 (N_1189,In_789,In_459);
xor U1190 (N_1190,In_549,In_1255);
or U1191 (N_1191,In_773,In_605);
or U1192 (N_1192,In_413,In_1463);
nor U1193 (N_1193,In_357,In_366);
and U1194 (N_1194,In_937,In_488);
or U1195 (N_1195,In_86,In_99);
nand U1196 (N_1196,In_965,In_1165);
or U1197 (N_1197,In_682,In_689);
xnor U1198 (N_1198,In_1108,In_914);
nor U1199 (N_1199,In_130,In_1237);
nand U1200 (N_1200,In_246,In_920);
xnor U1201 (N_1201,In_1088,In_108);
nand U1202 (N_1202,In_1045,In_25);
nor U1203 (N_1203,In_478,In_410);
nor U1204 (N_1204,In_575,In_528);
xnor U1205 (N_1205,In_1240,In_160);
and U1206 (N_1206,In_1008,In_1239);
nor U1207 (N_1207,In_1093,In_1313);
or U1208 (N_1208,In_392,In_728);
nor U1209 (N_1209,In_401,In_120);
nand U1210 (N_1210,In_304,In_411);
and U1211 (N_1211,In_960,In_1362);
and U1212 (N_1212,In_1395,In_165);
nand U1213 (N_1213,In_716,In_783);
or U1214 (N_1214,In_379,In_204);
nor U1215 (N_1215,In_46,In_653);
nor U1216 (N_1216,In_328,In_90);
nor U1217 (N_1217,In_111,In_1075);
nor U1218 (N_1218,In_317,In_395);
nand U1219 (N_1219,In_1300,In_1138);
nor U1220 (N_1220,In_1093,In_687);
or U1221 (N_1221,In_1306,In_118);
nor U1222 (N_1222,In_737,In_19);
nand U1223 (N_1223,In_1286,In_19);
and U1224 (N_1224,In_290,In_1311);
nand U1225 (N_1225,In_297,In_268);
nand U1226 (N_1226,In_237,In_174);
nor U1227 (N_1227,In_69,In_1309);
nor U1228 (N_1228,In_229,In_414);
and U1229 (N_1229,In_255,In_498);
or U1230 (N_1230,In_1311,In_11);
nand U1231 (N_1231,In_112,In_1318);
nor U1232 (N_1232,In_1136,In_1246);
and U1233 (N_1233,In_1409,In_167);
and U1234 (N_1234,In_783,In_869);
or U1235 (N_1235,In_724,In_353);
or U1236 (N_1236,In_56,In_120);
or U1237 (N_1237,In_1187,In_1207);
nand U1238 (N_1238,In_828,In_142);
nand U1239 (N_1239,In_835,In_1323);
xnor U1240 (N_1240,In_816,In_197);
nor U1241 (N_1241,In_280,In_501);
xor U1242 (N_1242,In_672,In_1444);
or U1243 (N_1243,In_508,In_1058);
or U1244 (N_1244,In_49,In_229);
nand U1245 (N_1245,In_495,In_1306);
or U1246 (N_1246,In_230,In_1470);
and U1247 (N_1247,In_944,In_449);
xnor U1248 (N_1248,In_432,In_1481);
nand U1249 (N_1249,In_1048,In_640);
nor U1250 (N_1250,In_590,In_514);
nor U1251 (N_1251,In_339,In_830);
and U1252 (N_1252,In_288,In_1242);
and U1253 (N_1253,In_1438,In_1324);
xor U1254 (N_1254,In_1064,In_425);
or U1255 (N_1255,In_991,In_1338);
nor U1256 (N_1256,In_1401,In_273);
and U1257 (N_1257,In_282,In_373);
or U1258 (N_1258,In_169,In_724);
xnor U1259 (N_1259,In_5,In_828);
and U1260 (N_1260,In_325,In_924);
nand U1261 (N_1261,In_1073,In_1346);
and U1262 (N_1262,In_619,In_465);
or U1263 (N_1263,In_1459,In_672);
and U1264 (N_1264,In_547,In_1223);
and U1265 (N_1265,In_1184,In_31);
or U1266 (N_1266,In_389,In_1397);
or U1267 (N_1267,In_408,In_724);
nor U1268 (N_1268,In_239,In_71);
and U1269 (N_1269,In_1497,In_1062);
or U1270 (N_1270,In_271,In_1432);
and U1271 (N_1271,In_1187,In_241);
nor U1272 (N_1272,In_481,In_1179);
or U1273 (N_1273,In_1484,In_1098);
xnor U1274 (N_1274,In_845,In_1251);
or U1275 (N_1275,In_480,In_149);
or U1276 (N_1276,In_81,In_910);
nand U1277 (N_1277,In_1191,In_57);
or U1278 (N_1278,In_628,In_356);
nor U1279 (N_1279,In_1239,In_801);
nand U1280 (N_1280,In_1023,In_967);
and U1281 (N_1281,In_173,In_1206);
nor U1282 (N_1282,In_208,In_1211);
nand U1283 (N_1283,In_724,In_683);
and U1284 (N_1284,In_292,In_72);
xnor U1285 (N_1285,In_1121,In_1455);
or U1286 (N_1286,In_969,In_1067);
nand U1287 (N_1287,In_487,In_1443);
nor U1288 (N_1288,In_258,In_176);
nor U1289 (N_1289,In_1093,In_862);
nand U1290 (N_1290,In_243,In_445);
and U1291 (N_1291,In_1063,In_551);
nor U1292 (N_1292,In_298,In_846);
and U1293 (N_1293,In_569,In_1434);
or U1294 (N_1294,In_1247,In_1272);
or U1295 (N_1295,In_76,In_150);
nor U1296 (N_1296,In_8,In_1191);
nor U1297 (N_1297,In_780,In_1391);
or U1298 (N_1298,In_477,In_969);
nand U1299 (N_1299,In_106,In_832);
and U1300 (N_1300,In_1403,In_400);
xor U1301 (N_1301,In_280,In_213);
and U1302 (N_1302,In_775,In_562);
nor U1303 (N_1303,In_221,In_1068);
nand U1304 (N_1304,In_882,In_1114);
nor U1305 (N_1305,In_1272,In_1016);
nor U1306 (N_1306,In_1454,In_757);
or U1307 (N_1307,In_834,In_1135);
nand U1308 (N_1308,In_727,In_688);
nand U1309 (N_1309,In_941,In_1361);
nor U1310 (N_1310,In_1064,In_405);
nor U1311 (N_1311,In_231,In_1299);
or U1312 (N_1312,In_1019,In_773);
nor U1313 (N_1313,In_1030,In_544);
or U1314 (N_1314,In_1396,In_406);
or U1315 (N_1315,In_1018,In_435);
nor U1316 (N_1316,In_257,In_101);
and U1317 (N_1317,In_198,In_477);
nand U1318 (N_1318,In_436,In_1400);
nor U1319 (N_1319,In_1498,In_83);
and U1320 (N_1320,In_701,In_955);
nand U1321 (N_1321,In_1389,In_84);
or U1322 (N_1322,In_802,In_658);
or U1323 (N_1323,In_1413,In_1255);
nor U1324 (N_1324,In_1031,In_110);
or U1325 (N_1325,In_201,In_257);
nand U1326 (N_1326,In_30,In_1142);
and U1327 (N_1327,In_1353,In_417);
nand U1328 (N_1328,In_1030,In_918);
and U1329 (N_1329,In_752,In_843);
nor U1330 (N_1330,In_1436,In_278);
xor U1331 (N_1331,In_1115,In_1470);
nor U1332 (N_1332,In_1391,In_1182);
nor U1333 (N_1333,In_890,In_1332);
and U1334 (N_1334,In_1104,In_300);
or U1335 (N_1335,In_1249,In_872);
and U1336 (N_1336,In_1276,In_1141);
nor U1337 (N_1337,In_1256,In_1249);
nor U1338 (N_1338,In_1163,In_1135);
and U1339 (N_1339,In_838,In_350);
or U1340 (N_1340,In_191,In_38);
nand U1341 (N_1341,In_588,In_726);
or U1342 (N_1342,In_403,In_540);
or U1343 (N_1343,In_571,In_175);
nor U1344 (N_1344,In_1035,In_249);
and U1345 (N_1345,In_918,In_318);
or U1346 (N_1346,In_222,In_448);
or U1347 (N_1347,In_1412,In_745);
nand U1348 (N_1348,In_465,In_326);
nand U1349 (N_1349,In_204,In_413);
xnor U1350 (N_1350,In_551,In_73);
nor U1351 (N_1351,In_329,In_362);
nand U1352 (N_1352,In_803,In_1381);
nor U1353 (N_1353,In_574,In_111);
nand U1354 (N_1354,In_211,In_490);
nand U1355 (N_1355,In_1314,In_1464);
or U1356 (N_1356,In_96,In_1425);
xnor U1357 (N_1357,In_562,In_1359);
xnor U1358 (N_1358,In_658,In_261);
or U1359 (N_1359,In_622,In_1366);
nor U1360 (N_1360,In_1084,In_707);
nand U1361 (N_1361,In_644,In_1478);
nor U1362 (N_1362,In_360,In_41);
or U1363 (N_1363,In_1166,In_509);
and U1364 (N_1364,In_717,In_837);
nor U1365 (N_1365,In_324,In_378);
nor U1366 (N_1366,In_1353,In_1464);
or U1367 (N_1367,In_23,In_340);
nand U1368 (N_1368,In_899,In_844);
nand U1369 (N_1369,In_913,In_231);
nor U1370 (N_1370,In_288,In_950);
nor U1371 (N_1371,In_93,In_608);
nand U1372 (N_1372,In_63,In_445);
nand U1373 (N_1373,In_1464,In_879);
or U1374 (N_1374,In_633,In_36);
or U1375 (N_1375,In_513,In_1475);
or U1376 (N_1376,In_678,In_1212);
or U1377 (N_1377,In_1329,In_806);
nand U1378 (N_1378,In_1281,In_434);
nand U1379 (N_1379,In_1177,In_393);
or U1380 (N_1380,In_1335,In_629);
or U1381 (N_1381,In_1209,In_869);
and U1382 (N_1382,In_740,In_96);
nor U1383 (N_1383,In_231,In_752);
nand U1384 (N_1384,In_347,In_244);
and U1385 (N_1385,In_620,In_567);
nand U1386 (N_1386,In_147,In_238);
and U1387 (N_1387,In_297,In_593);
nor U1388 (N_1388,In_597,In_1379);
nand U1389 (N_1389,In_1109,In_236);
or U1390 (N_1390,In_1420,In_1366);
nor U1391 (N_1391,In_1081,In_58);
nand U1392 (N_1392,In_183,In_267);
nor U1393 (N_1393,In_945,In_1058);
nand U1394 (N_1394,In_377,In_666);
nor U1395 (N_1395,In_1076,In_600);
nand U1396 (N_1396,In_85,In_268);
nand U1397 (N_1397,In_1273,In_737);
nor U1398 (N_1398,In_538,In_384);
nand U1399 (N_1399,In_597,In_420);
and U1400 (N_1400,In_137,In_1097);
and U1401 (N_1401,In_438,In_277);
and U1402 (N_1402,In_231,In_349);
or U1403 (N_1403,In_1445,In_1124);
or U1404 (N_1404,In_54,In_472);
and U1405 (N_1405,In_1263,In_1233);
nand U1406 (N_1406,In_1398,In_1149);
nor U1407 (N_1407,In_1109,In_800);
and U1408 (N_1408,In_1206,In_1006);
nor U1409 (N_1409,In_287,In_655);
xnor U1410 (N_1410,In_1118,In_1021);
and U1411 (N_1411,In_1405,In_375);
nor U1412 (N_1412,In_364,In_1428);
and U1413 (N_1413,In_330,In_248);
or U1414 (N_1414,In_500,In_1038);
xnor U1415 (N_1415,In_264,In_1250);
or U1416 (N_1416,In_275,In_523);
nor U1417 (N_1417,In_510,In_892);
nor U1418 (N_1418,In_181,In_973);
nor U1419 (N_1419,In_879,In_609);
nor U1420 (N_1420,In_1150,In_1231);
nor U1421 (N_1421,In_1359,In_719);
nand U1422 (N_1422,In_797,In_300);
or U1423 (N_1423,In_918,In_1158);
or U1424 (N_1424,In_402,In_308);
or U1425 (N_1425,In_669,In_806);
or U1426 (N_1426,In_1125,In_158);
and U1427 (N_1427,In_357,In_394);
or U1428 (N_1428,In_569,In_1018);
or U1429 (N_1429,In_162,In_806);
nand U1430 (N_1430,In_739,In_1472);
xnor U1431 (N_1431,In_200,In_392);
xor U1432 (N_1432,In_809,In_1171);
or U1433 (N_1433,In_920,In_1448);
or U1434 (N_1434,In_829,In_816);
xor U1435 (N_1435,In_386,In_1052);
nor U1436 (N_1436,In_352,In_989);
and U1437 (N_1437,In_608,In_316);
or U1438 (N_1438,In_953,In_307);
nor U1439 (N_1439,In_989,In_884);
nor U1440 (N_1440,In_276,In_1446);
xnor U1441 (N_1441,In_335,In_650);
and U1442 (N_1442,In_656,In_173);
or U1443 (N_1443,In_404,In_463);
xnor U1444 (N_1444,In_911,In_149);
or U1445 (N_1445,In_801,In_647);
and U1446 (N_1446,In_46,In_61);
and U1447 (N_1447,In_1036,In_1320);
xor U1448 (N_1448,In_241,In_919);
nand U1449 (N_1449,In_831,In_158);
or U1450 (N_1450,In_1110,In_832);
nand U1451 (N_1451,In_463,In_105);
nor U1452 (N_1452,In_837,In_1352);
nor U1453 (N_1453,In_944,In_453);
nand U1454 (N_1454,In_74,In_283);
or U1455 (N_1455,In_1342,In_795);
nor U1456 (N_1456,In_642,In_1059);
and U1457 (N_1457,In_1155,In_955);
xnor U1458 (N_1458,In_822,In_1474);
nand U1459 (N_1459,In_534,In_571);
or U1460 (N_1460,In_686,In_645);
xnor U1461 (N_1461,In_1163,In_1194);
nor U1462 (N_1462,In_1449,In_1408);
xnor U1463 (N_1463,In_1484,In_1287);
nand U1464 (N_1464,In_1314,In_771);
and U1465 (N_1465,In_305,In_1368);
nor U1466 (N_1466,In_289,In_701);
nor U1467 (N_1467,In_991,In_1335);
nor U1468 (N_1468,In_1485,In_886);
or U1469 (N_1469,In_1076,In_1010);
nand U1470 (N_1470,In_1140,In_1190);
nor U1471 (N_1471,In_1308,In_396);
xnor U1472 (N_1472,In_137,In_217);
nor U1473 (N_1473,In_249,In_758);
nand U1474 (N_1474,In_1258,In_923);
nor U1475 (N_1475,In_1093,In_698);
and U1476 (N_1476,In_459,In_651);
nand U1477 (N_1477,In_704,In_382);
or U1478 (N_1478,In_960,In_1256);
nand U1479 (N_1479,In_1448,In_376);
nor U1480 (N_1480,In_139,In_384);
or U1481 (N_1481,In_809,In_749);
and U1482 (N_1482,In_1397,In_922);
or U1483 (N_1483,In_631,In_1395);
or U1484 (N_1484,In_3,In_1223);
or U1485 (N_1485,In_1480,In_490);
or U1486 (N_1486,In_863,In_1084);
or U1487 (N_1487,In_1381,In_1128);
or U1488 (N_1488,In_657,In_784);
and U1489 (N_1489,In_535,In_492);
or U1490 (N_1490,In_112,In_1242);
or U1491 (N_1491,In_741,In_472);
nand U1492 (N_1492,In_8,In_887);
nand U1493 (N_1493,In_1095,In_244);
and U1494 (N_1494,In_886,In_1132);
nand U1495 (N_1495,In_1367,In_199);
xor U1496 (N_1496,In_1308,In_1095);
and U1497 (N_1497,In_852,In_1145);
xnor U1498 (N_1498,In_62,In_626);
nor U1499 (N_1499,In_899,In_1386);
or U1500 (N_1500,N_923,N_223);
nand U1501 (N_1501,N_1302,N_1121);
nand U1502 (N_1502,N_236,N_1448);
nor U1503 (N_1503,N_621,N_186);
nand U1504 (N_1504,N_619,N_1422);
nor U1505 (N_1505,N_1069,N_1096);
nor U1506 (N_1506,N_44,N_22);
and U1507 (N_1507,N_154,N_951);
or U1508 (N_1508,N_1040,N_1081);
or U1509 (N_1509,N_1166,N_513);
nor U1510 (N_1510,N_294,N_1375);
or U1511 (N_1511,N_1046,N_651);
and U1512 (N_1512,N_784,N_815);
and U1513 (N_1513,N_773,N_208);
nand U1514 (N_1514,N_311,N_293);
nand U1515 (N_1515,N_939,N_347);
nor U1516 (N_1516,N_893,N_1215);
or U1517 (N_1517,N_1473,N_234);
or U1518 (N_1518,N_827,N_216);
or U1519 (N_1519,N_752,N_662);
nand U1520 (N_1520,N_864,N_1167);
or U1521 (N_1521,N_47,N_252);
or U1522 (N_1522,N_366,N_681);
nor U1523 (N_1523,N_887,N_181);
nand U1524 (N_1524,N_788,N_1230);
and U1525 (N_1525,N_429,N_30);
or U1526 (N_1526,N_356,N_20);
and U1527 (N_1527,N_903,N_944);
nand U1528 (N_1528,N_885,N_1218);
nor U1529 (N_1529,N_1184,N_221);
nand U1530 (N_1530,N_1074,N_1236);
or U1531 (N_1531,N_574,N_861);
or U1532 (N_1532,N_1350,N_835);
or U1533 (N_1533,N_1283,N_858);
nor U1534 (N_1534,N_37,N_174);
nand U1535 (N_1535,N_1421,N_488);
nor U1536 (N_1536,N_1367,N_1151);
and U1537 (N_1537,N_904,N_1177);
xor U1538 (N_1538,N_1106,N_510);
nor U1539 (N_1539,N_1005,N_557);
nor U1540 (N_1540,N_355,N_516);
nand U1541 (N_1541,N_563,N_1010);
and U1542 (N_1542,N_1150,N_29);
nand U1543 (N_1543,N_363,N_1254);
nor U1544 (N_1544,N_799,N_1045);
or U1545 (N_1545,N_1039,N_1414);
xnor U1546 (N_1546,N_1057,N_793);
and U1547 (N_1547,N_258,N_484);
or U1548 (N_1548,N_1424,N_1380);
nand U1549 (N_1549,N_260,N_834);
or U1550 (N_1550,N_928,N_1337);
nor U1551 (N_1551,N_988,N_1193);
or U1552 (N_1552,N_105,N_712);
or U1553 (N_1553,N_612,N_1373);
xnor U1554 (N_1554,N_532,N_714);
nor U1555 (N_1555,N_359,N_1468);
and U1556 (N_1556,N_1044,N_756);
nand U1557 (N_1557,N_897,N_239);
nor U1558 (N_1558,N_1396,N_1155);
nand U1559 (N_1559,N_685,N_1338);
nand U1560 (N_1560,N_1162,N_1029);
nand U1561 (N_1561,N_1488,N_556);
or U1562 (N_1562,N_1273,N_1312);
or U1563 (N_1563,N_704,N_880);
nor U1564 (N_1564,N_1111,N_760);
or U1565 (N_1565,N_933,N_1371);
nand U1566 (N_1566,N_503,N_671);
and U1567 (N_1567,N_411,N_164);
or U1568 (N_1568,N_200,N_110);
nand U1569 (N_1569,N_640,N_241);
or U1570 (N_1570,N_423,N_1159);
and U1571 (N_1571,N_505,N_1058);
nor U1572 (N_1572,N_1209,N_1353);
nand U1573 (N_1573,N_322,N_1191);
nand U1574 (N_1574,N_298,N_713);
nor U1575 (N_1575,N_531,N_1282);
nor U1576 (N_1576,N_1387,N_2);
and U1577 (N_1577,N_1087,N_768);
nand U1578 (N_1578,N_907,N_843);
xor U1579 (N_1579,N_661,N_916);
or U1580 (N_1580,N_1319,N_68);
and U1581 (N_1581,N_462,N_909);
nor U1582 (N_1582,N_1153,N_971);
xnor U1583 (N_1583,N_314,N_419);
or U1584 (N_1584,N_300,N_1298);
nand U1585 (N_1585,N_1031,N_1059);
or U1586 (N_1586,N_1052,N_1126);
nor U1587 (N_1587,N_286,N_1496);
and U1588 (N_1588,N_1118,N_1103);
xnor U1589 (N_1589,N_213,N_740);
and U1590 (N_1590,N_833,N_1133);
nor U1591 (N_1591,N_1013,N_986);
nor U1592 (N_1592,N_689,N_1024);
nor U1593 (N_1593,N_635,N_36);
xor U1594 (N_1594,N_228,N_570);
or U1595 (N_1595,N_587,N_425);
and U1596 (N_1596,N_1214,N_395);
and U1597 (N_1597,N_70,N_401);
nand U1598 (N_1598,N_472,N_708);
nor U1599 (N_1599,N_614,N_1169);
or U1600 (N_1600,N_962,N_109);
and U1601 (N_1601,N_977,N_999);
nand U1602 (N_1602,N_1378,N_1480);
nand U1603 (N_1603,N_95,N_480);
or U1604 (N_1604,N_1123,N_232);
and U1605 (N_1605,N_1347,N_1038);
or U1606 (N_1606,N_1016,N_1385);
or U1607 (N_1607,N_968,N_950);
or U1608 (N_1608,N_953,N_348);
or U1609 (N_1609,N_894,N_1438);
and U1610 (N_1610,N_371,N_309);
and U1611 (N_1611,N_987,N_895);
nand U1612 (N_1612,N_508,N_633);
nor U1613 (N_1613,N_1134,N_1394);
xnor U1614 (N_1614,N_757,N_1355);
and U1615 (N_1615,N_1291,N_952);
and U1616 (N_1616,N_1474,N_892);
xor U1617 (N_1617,N_1293,N_645);
or U1618 (N_1618,N_1322,N_1237);
nor U1619 (N_1619,N_278,N_440);
and U1620 (N_1620,N_726,N_1275);
and U1621 (N_1621,N_137,N_1444);
nor U1622 (N_1622,N_749,N_433);
nand U1623 (N_1623,N_1303,N_1374);
and U1624 (N_1624,N_447,N_468);
nor U1625 (N_1625,N_1416,N_461);
nand U1626 (N_1626,N_1075,N_1120);
and U1627 (N_1627,N_1182,N_1221);
or U1628 (N_1628,N_736,N_634);
or U1629 (N_1629,N_1,N_402);
nor U1630 (N_1630,N_945,N_924);
or U1631 (N_1631,N_1195,N_703);
xor U1632 (N_1632,N_869,N_99);
nor U1633 (N_1633,N_1160,N_828);
nor U1634 (N_1634,N_1464,N_600);
or U1635 (N_1635,N_343,N_394);
xnor U1636 (N_1636,N_1112,N_504);
and U1637 (N_1637,N_1135,N_731);
nand U1638 (N_1638,N_568,N_1241);
or U1639 (N_1639,N_195,N_459);
or U1640 (N_1640,N_1170,N_849);
xnor U1641 (N_1641,N_1430,N_1128);
xor U1642 (N_1642,N_1261,N_418);
and U1643 (N_1643,N_997,N_791);
nor U1644 (N_1644,N_1203,N_1376);
nor U1645 (N_1645,N_872,N_350);
nand U1646 (N_1646,N_98,N_1392);
nand U1647 (N_1647,N_145,N_360);
nor U1648 (N_1648,N_1107,N_9);
and U1649 (N_1649,N_812,N_1406);
nand U1650 (N_1650,N_1099,N_352);
and U1651 (N_1651,N_1475,N_1346);
nor U1652 (N_1652,N_1239,N_474);
or U1653 (N_1653,N_400,N_61);
or U1654 (N_1654,N_535,N_1379);
nor U1655 (N_1655,N_1307,N_1117);
xor U1656 (N_1656,N_743,N_437);
nand U1657 (N_1657,N_850,N_390);
nor U1658 (N_1658,N_375,N_1130);
and U1659 (N_1659,N_798,N_284);
nand U1660 (N_1660,N_163,N_1043);
and U1661 (N_1661,N_744,N_617);
and U1662 (N_1662,N_450,N_102);
nand U1663 (N_1663,N_644,N_540);
nand U1664 (N_1664,N_1328,N_1268);
and U1665 (N_1665,N_478,N_18);
or U1666 (N_1666,N_72,N_1274);
nor U1667 (N_1667,N_122,N_1369);
nand U1668 (N_1668,N_1224,N_1455);
and U1669 (N_1669,N_1090,N_1255);
nand U1670 (N_1670,N_615,N_76);
nand U1671 (N_1671,N_193,N_285);
nor U1672 (N_1672,N_603,N_762);
or U1673 (N_1673,N_1484,N_1101);
nor U1674 (N_1674,N_959,N_1073);
and U1675 (N_1675,N_1469,N_638);
or U1676 (N_1676,N_316,N_441);
nor U1677 (N_1677,N_697,N_595);
nor U1678 (N_1678,N_995,N_591);
nor U1679 (N_1679,N_514,N_722);
or U1680 (N_1680,N_1427,N_3);
nor U1681 (N_1681,N_1290,N_248);
nor U1682 (N_1682,N_1051,N_807);
xor U1683 (N_1683,N_367,N_761);
xor U1684 (N_1684,N_976,N_1356);
nand U1685 (N_1685,N_203,N_659);
nor U1686 (N_1686,N_583,N_982);
xnor U1687 (N_1687,N_702,N_271);
or U1688 (N_1688,N_111,N_874);
or U1689 (N_1689,N_463,N_1233);
and U1690 (N_1690,N_1381,N_1127);
nand U1691 (N_1691,N_868,N_106);
nand U1692 (N_1692,N_179,N_1026);
and U1693 (N_1693,N_1390,N_1110);
nor U1694 (N_1694,N_158,N_627);
or U1695 (N_1695,N_281,N_144);
nand U1696 (N_1696,N_911,N_139);
or U1697 (N_1697,N_149,N_270);
nand U1698 (N_1698,N_104,N_1078);
nor U1699 (N_1699,N_739,N_1194);
nand U1700 (N_1700,N_431,N_166);
xor U1701 (N_1701,N_1272,N_732);
and U1702 (N_1702,N_225,N_1345);
and U1703 (N_1703,N_1143,N_51);
or U1704 (N_1704,N_707,N_862);
nor U1705 (N_1705,N_1049,N_1401);
or U1706 (N_1706,N_1494,N_209);
nor U1707 (N_1707,N_940,N_1316);
nand U1708 (N_1708,N_1163,N_918);
and U1709 (N_1709,N_1242,N_597);
nor U1710 (N_1710,N_94,N_994);
nand U1711 (N_1711,N_27,N_175);
nand U1712 (N_1712,N_912,N_1451);
nor U1713 (N_1713,N_191,N_667);
nand U1714 (N_1714,N_866,N_368);
nand U1715 (N_1715,N_1186,N_1459);
and U1716 (N_1716,N_335,N_444);
nand U1717 (N_1717,N_771,N_253);
and U1718 (N_1718,N_683,N_491);
and U1719 (N_1719,N_1084,N_86);
and U1720 (N_1720,N_721,N_1048);
and U1721 (N_1721,N_879,N_21);
or U1722 (N_1722,N_160,N_465);
nand U1723 (N_1723,N_124,N_738);
or U1724 (N_1724,N_454,N_929);
or U1725 (N_1725,N_416,N_1280);
nand U1726 (N_1726,N_1364,N_292);
or U1727 (N_1727,N_1413,N_753);
or U1728 (N_1728,N_782,N_1253);
nand U1729 (N_1729,N_679,N_1433);
nand U1730 (N_1730,N_471,N_1093);
or U1731 (N_1731,N_1020,N_63);
and U1732 (N_1732,N_1113,N_1011);
xnor U1733 (N_1733,N_764,N_825);
nor U1734 (N_1734,N_631,N_1348);
and U1735 (N_1735,N_1157,N_351);
and U1736 (N_1736,N_1384,N_935);
and U1737 (N_1737,N_943,N_1300);
and U1738 (N_1738,N_1012,N_930);
xor U1739 (N_1739,N_15,N_746);
nor U1740 (N_1740,N_674,N_985);
nand U1741 (N_1741,N_0,N_318);
nand U1742 (N_1742,N_1228,N_565);
or U1743 (N_1743,N_846,N_12);
nor U1744 (N_1744,N_646,N_1165);
nor U1745 (N_1745,N_1262,N_654);
nand U1746 (N_1746,N_1440,N_536);
or U1747 (N_1747,N_1426,N_1419);
nand U1748 (N_1748,N_259,N_448);
or U1749 (N_1749,N_677,N_134);
xnor U1750 (N_1750,N_837,N_628);
nor U1751 (N_1751,N_1004,N_1311);
nor U1752 (N_1752,N_177,N_1340);
or U1753 (N_1753,N_544,N_388);
and U1754 (N_1754,N_657,N_665);
xor U1755 (N_1755,N_446,N_1267);
or U1756 (N_1756,N_436,N_291);
and U1757 (N_1757,N_150,N_792);
or U1758 (N_1758,N_1377,N_715);
and U1759 (N_1759,N_129,N_676);
and U1760 (N_1760,N_1471,N_219);
xnor U1761 (N_1761,N_204,N_428);
nand U1762 (N_1762,N_80,N_1343);
or U1763 (N_1763,N_17,N_374);
and U1764 (N_1764,N_496,N_687);
nand U1765 (N_1765,N_955,N_641);
and U1766 (N_1766,N_967,N_970);
nand U1767 (N_1767,N_1017,N_485);
xor U1768 (N_1768,N_716,N_533);
or U1769 (N_1769,N_908,N_865);
nor U1770 (N_1770,N_1320,N_307);
and U1771 (N_1771,N_24,N_282);
and U1772 (N_1772,N_1189,N_362);
and U1773 (N_1773,N_1225,N_40);
and U1774 (N_1774,N_821,N_332);
xnor U1775 (N_1775,N_421,N_691);
nor U1776 (N_1776,N_148,N_915);
or U1777 (N_1777,N_1206,N_289);
nor U1778 (N_1778,N_336,N_1144);
nor U1779 (N_1779,N_519,N_117);
nor U1780 (N_1780,N_571,N_1349);
or U1781 (N_1781,N_706,N_888);
nand U1782 (N_1782,N_1313,N_1139);
nor U1783 (N_1783,N_1244,N_647);
nand U1784 (N_1784,N_590,N_247);
or U1785 (N_1785,N_1014,N_413);
or U1786 (N_1786,N_408,N_460);
nor U1787 (N_1787,N_1372,N_1063);
nor U1788 (N_1788,N_701,N_430);
or U1789 (N_1789,N_919,N_594);
nand U1790 (N_1790,N_178,N_656);
xor U1791 (N_1791,N_1247,N_1131);
nor U1792 (N_1792,N_1257,N_73);
nand U1793 (N_1793,N_1327,N_487);
nor U1794 (N_1794,N_1173,N_32);
nor U1795 (N_1795,N_304,N_1216);
or U1796 (N_1796,N_1076,N_189);
nor U1797 (N_1797,N_1080,N_1007);
or U1798 (N_1798,N_1138,N_1095);
and U1799 (N_1799,N_121,N_1407);
nor U1800 (N_1800,N_517,N_153);
or U1801 (N_1801,N_720,N_1124);
nand U1802 (N_1802,N_1083,N_475);
or U1803 (N_1803,N_69,N_1466);
or U1804 (N_1804,N_1066,N_141);
and U1805 (N_1805,N_1408,N_758);
xnor U1806 (N_1806,N_1476,N_884);
nand U1807 (N_1807,N_42,N_183);
nand U1808 (N_1808,N_306,N_1399);
nor U1809 (N_1809,N_1329,N_1070);
nor U1810 (N_1810,N_123,N_507);
nand U1811 (N_1811,N_1270,N_326);
nor U1812 (N_1812,N_1425,N_339);
xor U1813 (N_1813,N_582,N_48);
nand U1814 (N_1814,N_1217,N_992);
and U1815 (N_1815,N_1091,N_1418);
and U1816 (N_1816,N_576,N_1437);
or U1817 (N_1817,N_422,N_1411);
nand U1818 (N_1818,N_599,N_287);
and U1819 (N_1819,N_1212,N_966);
or U1820 (N_1820,N_1287,N_692);
nand U1821 (N_1821,N_205,N_206);
xor U1822 (N_1822,N_337,N_776);
nand U1823 (N_1823,N_58,N_1019);
and U1824 (N_1824,N_56,N_1008);
or U1825 (N_1825,N_1188,N_804);
and U1826 (N_1826,N_10,N_1116);
and U1827 (N_1827,N_592,N_948);
nand U1828 (N_1828,N_1149,N_787);
nand U1829 (N_1829,N_639,N_853);
and U1830 (N_1830,N_1202,N_381);
or U1831 (N_1831,N_564,N_1449);
or U1832 (N_1832,N_878,N_1092);
nand U1833 (N_1833,N_13,N_1285);
nand U1834 (N_1834,N_949,N_957);
nor U1835 (N_1835,N_303,N_1428);
nor U1836 (N_1836,N_1393,N_663);
nor U1837 (N_1837,N_584,N_373);
nor U1838 (N_1838,N_1432,N_876);
or U1839 (N_1839,N_889,N_192);
or U1840 (N_1840,N_115,N_1317);
nor U1841 (N_1841,N_295,N_705);
and U1842 (N_1842,N_280,N_700);
nor U1843 (N_1843,N_742,N_328);
nor U1844 (N_1844,N_152,N_477);
nand U1845 (N_1845,N_710,N_856);
or U1846 (N_1846,N_389,N_509);
and U1847 (N_1847,N_473,N_6);
nand U1848 (N_1848,N_937,N_1132);
nand U1849 (N_1849,N_101,N_755);
nor U1850 (N_1850,N_523,N_699);
or U1851 (N_1851,N_308,N_1243);
or U1852 (N_1852,N_978,N_1382);
and U1853 (N_1853,N_218,N_142);
or U1854 (N_1854,N_1315,N_66);
nand U1855 (N_1855,N_763,N_156);
or U1856 (N_1856,N_396,N_860);
or U1857 (N_1857,N_873,N_824);
and U1858 (N_1858,N_1219,N_1006);
xor U1859 (N_1859,N_397,N_961);
xor U1860 (N_1860,N_172,N_385);
nor U1861 (N_1861,N_1079,N_745);
or U1862 (N_1862,N_1276,N_201);
or U1863 (N_1863,N_759,N_1478);
xnor U1864 (N_1864,N_890,N_62);
nand U1865 (N_1865,N_1023,N_197);
or U1866 (N_1866,N_1498,N_386);
nor U1867 (N_1867,N_341,N_1154);
and U1868 (N_1868,N_1325,N_35);
or U1869 (N_1869,N_524,N_684);
nor U1870 (N_1870,N_1213,N_1234);
or U1871 (N_1871,N_1050,N_1199);
and U1872 (N_1872,N_242,N_266);
nor U1873 (N_1873,N_1077,N_767);
or U1874 (N_1874,N_273,N_159);
and U1875 (N_1875,N_991,N_558);
or U1876 (N_1876,N_1002,N_1477);
nor U1877 (N_1877,N_354,N_1062);
and U1878 (N_1878,N_1022,N_1196);
and U1879 (N_1879,N_613,N_136);
nand U1880 (N_1880,N_493,N_596);
or U1881 (N_1881,N_1339,N_1391);
xor U1882 (N_1882,N_237,N_83);
nand U1883 (N_1883,N_1171,N_457);
and U1884 (N_1884,N_727,N_648);
or U1885 (N_1885,N_199,N_182);
or U1886 (N_1886,N_1210,N_905);
and U1887 (N_1887,N_254,N_901);
nor U1888 (N_1888,N_276,N_777);
nand U1889 (N_1889,N_1483,N_1447);
and U1890 (N_1890,N_979,N_211);
and U1891 (N_1891,N_1457,N_364);
xor U1892 (N_1892,N_79,N_766);
and U1893 (N_1893,N_800,N_891);
nor U1894 (N_1894,N_451,N_649);
or U1895 (N_1895,N_1493,N_1067);
and U1896 (N_1896,N_906,N_358);
nand U1897 (N_1897,N_1208,N_652);
nand U1898 (N_1898,N_403,N_551);
nor U1899 (N_1899,N_1492,N_658);
nor U1900 (N_1900,N_1088,N_795);
nand U1901 (N_1901,N_1129,N_476);
or U1902 (N_1902,N_1140,N_820);
nand U1903 (N_1903,N_1487,N_226);
xor U1904 (N_1904,N_67,N_954);
nor U1905 (N_1905,N_511,N_165);
nor U1906 (N_1906,N_779,N_575);
nand U1907 (N_1907,N_747,N_775);
and U1908 (N_1908,N_1174,N_1305);
or U1909 (N_1909,N_859,N_1299);
and U1910 (N_1910,N_902,N_816);
nand U1911 (N_1911,N_481,N_187);
xnor U1912 (N_1912,N_855,N_1489);
or U1913 (N_1913,N_1495,N_857);
and U1914 (N_1914,N_817,N_1003);
nand U1915 (N_1915,N_434,N_1156);
and U1916 (N_1916,N_97,N_313);
and U1917 (N_1917,N_1042,N_606);
or U1918 (N_1918,N_604,N_624);
and U1919 (N_1919,N_301,N_369);
nand U1920 (N_1920,N_718,N_1297);
or U1921 (N_1921,N_409,N_882);
nand U1922 (N_1922,N_1248,N_1161);
and U1923 (N_1923,N_632,N_113);
nor U1924 (N_1924,N_668,N_729);
or U1925 (N_1925,N_642,N_1086);
nand U1926 (N_1926,N_1398,N_126);
and U1927 (N_1927,N_1145,N_161);
and U1928 (N_1928,N_1168,N_499);
or U1929 (N_1929,N_1324,N_1064);
and U1930 (N_1930,N_1175,N_806);
nand U1931 (N_1931,N_841,N_1061);
or U1932 (N_1932,N_494,N_666);
and U1933 (N_1933,N_1470,N_1400);
or U1934 (N_1934,N_334,N_378);
xor U1935 (N_1935,N_31,N_464);
or U1936 (N_1936,N_1352,N_682);
and U1937 (N_1937,N_1001,N_370);
and U1938 (N_1938,N_1366,N_1310);
nor U1939 (N_1939,N_1085,N_439);
and U1940 (N_1940,N_1289,N_57);
nor U1941 (N_1941,N_1402,N_1190);
and U1942 (N_1942,N_789,N_1370);
xor U1943 (N_1943,N_498,N_809);
or U1944 (N_1944,N_60,N_424);
or U1945 (N_1945,N_1486,N_1205);
nand U1946 (N_1946,N_393,N_989);
nor U1947 (N_1947,N_610,N_321);
or U1948 (N_1948,N_342,N_735);
or U1949 (N_1949,N_8,N_100);
nand U1950 (N_1950,N_327,N_405);
nor U1951 (N_1951,N_1114,N_1499);
or U1952 (N_1952,N_169,N_412);
and U1953 (N_1953,N_840,N_251);
nor U1954 (N_1954,N_826,N_696);
or U1955 (N_1955,N_1431,N_215);
or U1956 (N_1956,N_1223,N_217);
nand U1957 (N_1957,N_936,N_340);
nor U1958 (N_1958,N_1397,N_754);
nor U1959 (N_1959,N_1410,N_618);
xnor U1960 (N_1960,N_1238,N_780);
and U1961 (N_1961,N_210,N_808);
nor U1962 (N_1962,N_543,N_1357);
nand U1963 (N_1963,N_709,N_751);
nand U1964 (N_1964,N_176,N_297);
and U1965 (N_1965,N_1259,N_686);
nand U1966 (N_1966,N_1220,N_1054);
or U1967 (N_1967,N_1441,N_87);
nor U1968 (N_1968,N_1028,N_1265);
and U1969 (N_1969,N_728,N_25);
nand U1970 (N_1970,N_814,N_1009);
nor U1971 (N_1971,N_1141,N_1197);
nor U1972 (N_1972,N_49,N_1122);
nor U1973 (N_1973,N_90,N_778);
and U1974 (N_1974,N_1335,N_427);
nand U1975 (N_1975,N_693,N_711);
xnor U1976 (N_1976,N_1445,N_625);
or U1977 (N_1977,N_1232,N_863);
and U1978 (N_1978,N_553,N_781);
nand U1979 (N_1979,N_1472,N_458);
and U1980 (N_1980,N_1341,N_675);
nand U1981 (N_1981,N_445,N_609);
and U1982 (N_1982,N_14,N_973);
nand U1983 (N_1983,N_325,N_1462);
xor U1984 (N_1984,N_53,N_1211);
nor U1985 (N_1985,N_1035,N_1331);
nor U1986 (N_1986,N_796,N_65);
xor U1987 (N_1987,N_1423,N_264);
nor U1988 (N_1988,N_1231,N_1458);
xnor U1989 (N_1989,N_1249,N_695);
and U1990 (N_1990,N_19,N_1294);
nand U1991 (N_1991,N_93,N_4);
xor U1992 (N_1992,N_1227,N_803);
or U1993 (N_1993,N_34,N_832);
and U1994 (N_1994,N_794,N_250);
nor U1995 (N_1995,N_222,N_956);
nand U1996 (N_1996,N_772,N_1108);
or U1997 (N_1997,N_622,N_1089);
or U1998 (N_1998,N_229,N_1342);
or U1999 (N_1999,N_567,N_518);
and U2000 (N_2000,N_1229,N_492);
and U2001 (N_2001,N_542,N_224);
nand U2002 (N_2002,N_82,N_1446);
and U2003 (N_2003,N_733,N_190);
xor U2004 (N_2004,N_143,N_1201);
and U2005 (N_2005,N_1187,N_1460);
and U2006 (N_2006,N_630,N_1260);
or U2007 (N_2007,N_184,N_108);
and U2008 (N_2008,N_453,N_257);
and U2009 (N_2009,N_1235,N_830);
and U2010 (N_2010,N_566,N_1256);
or U2011 (N_2011,N_1146,N_233);
and U2012 (N_2012,N_678,N_456);
or U2013 (N_2013,N_406,N_520);
nor U2014 (N_2014,N_1176,N_921);
nand U2015 (N_2015,N_883,N_398);
xor U2016 (N_2016,N_530,N_1333);
nor U2017 (N_2017,N_415,N_650);
xor U2018 (N_2018,N_914,N_960);
or U2019 (N_2019,N_410,N_1252);
xor U2020 (N_2020,N_797,N_585);
nor U2021 (N_2021,N_925,N_848);
nor U2022 (N_2022,N_1060,N_214);
nand U2023 (N_2023,N_1389,N_1318);
nand U2024 (N_2024,N_1222,N_317);
or U2025 (N_2025,N_330,N_133);
nand U2026 (N_2026,N_896,N_391);
xor U2027 (N_2027,N_277,N_120);
nor U2028 (N_2028,N_1358,N_1296);
nand U2029 (N_2029,N_435,N_361);
nand U2030 (N_2030,N_1395,N_502);
or U2031 (N_2031,N_196,N_265);
and U2032 (N_2032,N_1497,N_938);
or U2033 (N_2033,N_1180,N_33);
nor U2034 (N_2034,N_579,N_188);
nand U2035 (N_2035,N_107,N_512);
and U2036 (N_2036,N_212,N_443);
nand U2037 (N_2037,N_1158,N_338);
or U2038 (N_2038,N_984,N_823);
or U2039 (N_2039,N_268,N_765);
or U2040 (N_2040,N_1036,N_96);
and U2041 (N_2041,N_399,N_877);
nand U2042 (N_2042,N_1125,N_92);
nand U2043 (N_2043,N_1015,N_1207);
nor U2044 (N_2044,N_1344,N_934);
or U2045 (N_2045,N_324,N_231);
xor U2046 (N_2046,N_495,N_947);
or U2047 (N_2047,N_1362,N_500);
nor U2048 (N_2048,N_140,N_1456);
nor U2049 (N_2049,N_578,N_900);
nand U2050 (N_2050,N_1368,N_1304);
or U2051 (N_2051,N_546,N_554);
nor U2052 (N_2052,N_331,N_220);
nand U2053 (N_2053,N_1250,N_1271);
or U2054 (N_2054,N_5,N_312);
and U2055 (N_2055,N_917,N_547);
nor U2056 (N_2056,N_741,N_1109);
and U2057 (N_2057,N_1442,N_238);
or U2058 (N_2058,N_1306,N_1295);
or U2059 (N_2059,N_1485,N_515);
or U2060 (N_2060,N_1403,N_1415);
nand U2061 (N_2061,N_941,N_555);
and U2062 (N_2062,N_147,N_333);
and U2063 (N_2063,N_71,N_1490);
nand U2064 (N_2064,N_842,N_611);
nand U2065 (N_2065,N_1025,N_151);
xor U2066 (N_2066,N_41,N_1292);
or U2067 (N_2067,N_886,N_414);
nand U2068 (N_2068,N_871,N_572);
and U2069 (N_2069,N_64,N_269);
nor U2070 (N_2070,N_698,N_963);
nand U2071 (N_2071,N_819,N_466);
nor U2072 (N_2072,N_1030,N_1412);
or U2073 (N_2073,N_975,N_1192);
nor U2074 (N_2074,N_246,N_50);
and U2075 (N_2075,N_673,N_240);
and U2076 (N_2076,N_931,N_1068);
nand U2077 (N_2077,N_1251,N_75);
or U2078 (N_2078,N_1047,N_527);
nand U2079 (N_2079,N_724,N_1266);
and U2080 (N_2080,N_854,N_1033);
nor U2081 (N_2081,N_302,N_379);
and U2082 (N_2082,N_168,N_867);
or U2083 (N_2083,N_1027,N_1263);
nor U2084 (N_2084,N_561,N_586);
nand U2085 (N_2085,N_1467,N_1147);
xnor U2086 (N_2086,N_1308,N_1281);
and U2087 (N_2087,N_84,N_1443);
or U2088 (N_2088,N_349,N_1481);
or U2089 (N_2089,N_1336,N_483);
nor U2090 (N_2090,N_932,N_1098);
and U2091 (N_2091,N_1269,N_1258);
nand U2092 (N_2092,N_942,N_881);
or U2093 (N_2093,N_655,N_998);
or U2094 (N_2094,N_521,N_1104);
nor U2095 (N_2095,N_1326,N_382);
or U2096 (N_2096,N_103,N_89);
or U2097 (N_2097,N_690,N_972);
or U2098 (N_2098,N_55,N_227);
and U2099 (N_2099,N_275,N_417);
or U2100 (N_2100,N_245,N_602);
and U2101 (N_2101,N_620,N_323);
or U2102 (N_2102,N_501,N_244);
nor U2103 (N_2103,N_114,N_1491);
xor U2104 (N_2104,N_847,N_1181);
xnor U2105 (N_2105,N_875,N_545);
nor U2106 (N_2106,N_1071,N_1082);
and U2107 (N_2107,N_958,N_643);
and U2108 (N_2108,N_243,N_1204);
and U2109 (N_2109,N_927,N_497);
xnor U2110 (N_2110,N_7,N_489);
or U2111 (N_2111,N_1360,N_734);
xnor U2112 (N_2112,N_790,N_922);
nand U2113 (N_2113,N_490,N_783);
xnor U2114 (N_2114,N_608,N_125);
nor U2115 (N_2115,N_822,N_946);
and U2116 (N_2116,N_346,N_580);
or U2117 (N_2117,N_1332,N_1434);
nand U2118 (N_2118,N_964,N_1100);
xor U2119 (N_2119,N_77,N_1200);
nand U2120 (N_2120,N_1359,N_1179);
or U2121 (N_2121,N_249,N_1277);
or U2122 (N_2122,N_506,N_1321);
or U2123 (N_2123,N_965,N_980);
nand U2124 (N_2124,N_290,N_601);
nand U2125 (N_2125,N_1334,N_353);
nand U2126 (N_2126,N_59,N_329);
nor U2127 (N_2127,N_538,N_470);
and U2128 (N_2128,N_455,N_1436);
nand U2129 (N_2129,N_1439,N_670);
or U2130 (N_2130,N_852,N_1450);
nor U2131 (N_2131,N_380,N_319);
and U2132 (N_2132,N_629,N_1032);
and U2133 (N_2133,N_810,N_845);
and U2134 (N_2134,N_719,N_1279);
nand U2135 (N_2135,N_279,N_1018);
nand U2136 (N_2136,N_1136,N_235);
or U2137 (N_2137,N_526,N_46);
or U2138 (N_2138,N_1240,N_750);
and U2139 (N_2139,N_831,N_263);
nor U2140 (N_2140,N_785,N_157);
nand U2141 (N_2141,N_1094,N_1288);
nand U2142 (N_2142,N_479,N_320);
or U2143 (N_2143,N_315,N_774);
nor U2144 (N_2144,N_1330,N_119);
nand U2145 (N_2145,N_256,N_387);
and U2146 (N_2146,N_541,N_28);
xor U2147 (N_2147,N_267,N_283);
nand U2148 (N_2148,N_534,N_376);
or U2149 (N_2149,N_1482,N_1429);
and U2150 (N_2150,N_1178,N_1365);
nand U2151 (N_2151,N_469,N_805);
nor U2152 (N_2152,N_1137,N_198);
or U2153 (N_2153,N_420,N_230);
and U2154 (N_2154,N_426,N_1361);
nor U2155 (N_2155,N_131,N_528);
or U2156 (N_2156,N_272,N_786);
or U2157 (N_2157,N_1278,N_844);
and U2158 (N_2158,N_1034,N_274);
nand U2159 (N_2159,N_569,N_717);
or U2160 (N_2160,N_1383,N_1454);
and U2161 (N_2161,N_372,N_636);
and U2162 (N_2162,N_345,N_288);
and U2163 (N_2163,N_138,N_1323);
nand U2164 (N_2164,N_725,N_1102);
nor U2165 (N_2165,N_1000,N_1301);
nor U2166 (N_2166,N_467,N_870);
or U2167 (N_2167,N_432,N_1115);
and U2168 (N_2168,N_43,N_112);
or U2169 (N_2169,N_926,N_377);
nor U2170 (N_2170,N_920,N_680);
and U2171 (N_2171,N_913,N_616);
nor U2172 (N_2172,N_559,N_588);
nor U2173 (N_2173,N_653,N_85);
nand U2174 (N_2174,N_1053,N_128);
nand U2175 (N_2175,N_74,N_537);
and U2176 (N_2176,N_132,N_623);
and U2177 (N_2177,N_851,N_1097);
nor U2178 (N_2178,N_1479,N_1072);
nor U2179 (N_2179,N_748,N_983);
and U2180 (N_2180,N_1152,N_1065);
or U2181 (N_2181,N_769,N_801);
nor U2182 (N_2182,N_660,N_438);
and U2183 (N_2183,N_261,N_118);
nor U2184 (N_2184,N_770,N_1465);
nor U2185 (N_2185,N_1309,N_836);
nand U2186 (N_2186,N_482,N_813);
nand U2187 (N_2187,N_1056,N_1264);
xor U2188 (N_2188,N_88,N_996);
and U2189 (N_2189,N_26,N_1148);
nand U2190 (N_2190,N_255,N_170);
and U2191 (N_2191,N_1286,N_1185);
nor U2192 (N_2192,N_78,N_552);
or U2193 (N_2193,N_1404,N_1246);
or U2194 (N_2194,N_1172,N_990);
or U2195 (N_2195,N_299,N_1055);
or U2196 (N_2196,N_664,N_548);
or U2197 (N_2197,N_1463,N_1351);
and U2198 (N_2198,N_310,N_818);
and U2199 (N_2199,N_146,N_296);
and U2200 (N_2200,N_173,N_607);
nor U2201 (N_2201,N_11,N_560);
and U2202 (N_2202,N_357,N_802);
and U2203 (N_2203,N_1417,N_974);
and U2204 (N_2204,N_1388,N_344);
or U2205 (N_2205,N_442,N_162);
and U2206 (N_2206,N_525,N_1041);
xnor U2207 (N_2207,N_898,N_839);
nor U2208 (N_2208,N_39,N_1435);
nor U2209 (N_2209,N_185,N_672);
and U2210 (N_2210,N_23,N_993);
nor U2211 (N_2211,N_737,N_1198);
nor U2212 (N_2212,N_598,N_1245);
or U2213 (N_2213,N_838,N_593);
xor U2214 (N_2214,N_1105,N_38);
nand U2215 (N_2215,N_116,N_392);
or U2216 (N_2216,N_365,N_981);
or U2217 (N_2217,N_1142,N_383);
and U2218 (N_2218,N_171,N_52);
nor U2219 (N_2219,N_130,N_969);
or U2220 (N_2220,N_910,N_577);
or U2221 (N_2221,N_1386,N_1021);
nor U2222 (N_2222,N_1314,N_1452);
nor U2223 (N_2223,N_1183,N_1405);
xnor U2224 (N_2224,N_127,N_581);
and U2225 (N_2225,N_262,N_194);
nand U2226 (N_2226,N_1409,N_550);
nor U2227 (N_2227,N_135,N_305);
nor U2228 (N_2228,N_549,N_730);
nand U2229 (N_2229,N_669,N_539);
or U2230 (N_2230,N_407,N_180);
xnor U2231 (N_2231,N_1037,N_522);
nand U2232 (N_2232,N_1453,N_449);
and U2233 (N_2233,N_829,N_1354);
nor U2234 (N_2234,N_202,N_404);
xnor U2235 (N_2235,N_562,N_1119);
nor U2236 (N_2236,N_1461,N_452);
nor U2237 (N_2237,N_54,N_637);
nand U2238 (N_2238,N_899,N_573);
or U2239 (N_2239,N_91,N_1420);
nor U2240 (N_2240,N_626,N_1164);
and U2241 (N_2241,N_1363,N_1226);
and U2242 (N_2242,N_589,N_688);
nor U2243 (N_2243,N_207,N_155);
nor U2244 (N_2244,N_723,N_694);
and U2245 (N_2245,N_486,N_45);
or U2246 (N_2246,N_167,N_529);
or U2247 (N_2247,N_81,N_384);
nand U2248 (N_2248,N_811,N_1284);
nor U2249 (N_2249,N_605,N_16);
or U2250 (N_2250,N_1267,N_1054);
nor U2251 (N_2251,N_377,N_109);
nand U2252 (N_2252,N_32,N_772);
nand U2253 (N_2253,N_810,N_1379);
nor U2254 (N_2254,N_598,N_1031);
and U2255 (N_2255,N_1101,N_708);
or U2256 (N_2256,N_1037,N_1498);
and U2257 (N_2257,N_1465,N_1218);
and U2258 (N_2258,N_757,N_1483);
and U2259 (N_2259,N_646,N_208);
nand U2260 (N_2260,N_840,N_1085);
xnor U2261 (N_2261,N_1067,N_310);
nor U2262 (N_2262,N_539,N_1338);
nand U2263 (N_2263,N_951,N_1054);
nor U2264 (N_2264,N_697,N_1096);
xnor U2265 (N_2265,N_627,N_602);
or U2266 (N_2266,N_712,N_39);
or U2267 (N_2267,N_1238,N_1279);
nor U2268 (N_2268,N_532,N_323);
and U2269 (N_2269,N_1326,N_1223);
or U2270 (N_2270,N_1211,N_1174);
or U2271 (N_2271,N_360,N_699);
and U2272 (N_2272,N_715,N_291);
and U2273 (N_2273,N_534,N_784);
or U2274 (N_2274,N_125,N_138);
or U2275 (N_2275,N_482,N_1360);
or U2276 (N_2276,N_955,N_33);
or U2277 (N_2277,N_538,N_252);
and U2278 (N_2278,N_1085,N_772);
and U2279 (N_2279,N_91,N_199);
or U2280 (N_2280,N_1065,N_683);
or U2281 (N_2281,N_381,N_26);
nand U2282 (N_2282,N_1006,N_300);
nor U2283 (N_2283,N_363,N_475);
nand U2284 (N_2284,N_784,N_686);
xnor U2285 (N_2285,N_244,N_705);
nand U2286 (N_2286,N_182,N_488);
nand U2287 (N_2287,N_1423,N_734);
xnor U2288 (N_2288,N_1069,N_580);
nand U2289 (N_2289,N_1408,N_448);
nor U2290 (N_2290,N_899,N_985);
or U2291 (N_2291,N_741,N_920);
nand U2292 (N_2292,N_495,N_159);
xor U2293 (N_2293,N_731,N_358);
or U2294 (N_2294,N_619,N_620);
nand U2295 (N_2295,N_1001,N_318);
xor U2296 (N_2296,N_393,N_957);
and U2297 (N_2297,N_410,N_1464);
or U2298 (N_2298,N_1206,N_1062);
nor U2299 (N_2299,N_987,N_1370);
nand U2300 (N_2300,N_900,N_1294);
nor U2301 (N_2301,N_1342,N_1080);
nand U2302 (N_2302,N_1146,N_393);
or U2303 (N_2303,N_1022,N_285);
and U2304 (N_2304,N_661,N_645);
nand U2305 (N_2305,N_466,N_113);
and U2306 (N_2306,N_614,N_502);
xnor U2307 (N_2307,N_870,N_1210);
nand U2308 (N_2308,N_1350,N_983);
nand U2309 (N_2309,N_543,N_551);
or U2310 (N_2310,N_701,N_354);
nor U2311 (N_2311,N_70,N_894);
nand U2312 (N_2312,N_601,N_1422);
and U2313 (N_2313,N_54,N_1000);
xnor U2314 (N_2314,N_1240,N_123);
nand U2315 (N_2315,N_1158,N_466);
and U2316 (N_2316,N_1393,N_762);
nor U2317 (N_2317,N_542,N_125);
nor U2318 (N_2318,N_651,N_142);
or U2319 (N_2319,N_1089,N_1026);
nand U2320 (N_2320,N_24,N_423);
nand U2321 (N_2321,N_886,N_665);
nor U2322 (N_2322,N_198,N_1143);
nor U2323 (N_2323,N_236,N_206);
and U2324 (N_2324,N_1472,N_784);
or U2325 (N_2325,N_387,N_779);
or U2326 (N_2326,N_43,N_660);
and U2327 (N_2327,N_111,N_361);
xor U2328 (N_2328,N_1434,N_1253);
and U2329 (N_2329,N_395,N_110);
nor U2330 (N_2330,N_170,N_3);
or U2331 (N_2331,N_61,N_482);
nor U2332 (N_2332,N_974,N_1164);
or U2333 (N_2333,N_1369,N_329);
nand U2334 (N_2334,N_392,N_1477);
and U2335 (N_2335,N_889,N_105);
nor U2336 (N_2336,N_730,N_95);
nand U2337 (N_2337,N_810,N_194);
nor U2338 (N_2338,N_823,N_150);
nand U2339 (N_2339,N_6,N_450);
nor U2340 (N_2340,N_307,N_755);
and U2341 (N_2341,N_389,N_1022);
or U2342 (N_2342,N_267,N_1425);
and U2343 (N_2343,N_892,N_493);
or U2344 (N_2344,N_464,N_261);
nor U2345 (N_2345,N_18,N_374);
or U2346 (N_2346,N_556,N_570);
nand U2347 (N_2347,N_1142,N_503);
or U2348 (N_2348,N_395,N_956);
or U2349 (N_2349,N_537,N_82);
nand U2350 (N_2350,N_260,N_860);
xor U2351 (N_2351,N_1128,N_1066);
nor U2352 (N_2352,N_1084,N_442);
and U2353 (N_2353,N_312,N_163);
nand U2354 (N_2354,N_93,N_1341);
nor U2355 (N_2355,N_358,N_977);
or U2356 (N_2356,N_501,N_612);
nand U2357 (N_2357,N_778,N_335);
nand U2358 (N_2358,N_832,N_114);
nor U2359 (N_2359,N_13,N_1311);
or U2360 (N_2360,N_35,N_970);
or U2361 (N_2361,N_212,N_1144);
or U2362 (N_2362,N_1283,N_392);
or U2363 (N_2363,N_157,N_557);
nand U2364 (N_2364,N_115,N_17);
nor U2365 (N_2365,N_1444,N_1093);
or U2366 (N_2366,N_74,N_1290);
nor U2367 (N_2367,N_1113,N_851);
xor U2368 (N_2368,N_1299,N_350);
or U2369 (N_2369,N_390,N_1434);
and U2370 (N_2370,N_649,N_1057);
and U2371 (N_2371,N_1419,N_1177);
nor U2372 (N_2372,N_578,N_227);
or U2373 (N_2373,N_738,N_1106);
and U2374 (N_2374,N_964,N_1020);
xor U2375 (N_2375,N_232,N_1012);
xor U2376 (N_2376,N_1345,N_1);
and U2377 (N_2377,N_33,N_624);
and U2378 (N_2378,N_1289,N_1365);
and U2379 (N_2379,N_739,N_364);
nor U2380 (N_2380,N_194,N_1335);
nor U2381 (N_2381,N_532,N_1428);
nor U2382 (N_2382,N_342,N_1158);
or U2383 (N_2383,N_1380,N_912);
or U2384 (N_2384,N_972,N_794);
or U2385 (N_2385,N_1241,N_588);
or U2386 (N_2386,N_1245,N_1459);
nor U2387 (N_2387,N_1077,N_509);
and U2388 (N_2388,N_1141,N_329);
xor U2389 (N_2389,N_928,N_1095);
and U2390 (N_2390,N_537,N_1216);
xnor U2391 (N_2391,N_1035,N_567);
nand U2392 (N_2392,N_1246,N_1149);
nand U2393 (N_2393,N_332,N_642);
or U2394 (N_2394,N_211,N_131);
or U2395 (N_2395,N_1201,N_400);
nand U2396 (N_2396,N_180,N_486);
nor U2397 (N_2397,N_1402,N_115);
nand U2398 (N_2398,N_423,N_455);
and U2399 (N_2399,N_459,N_608);
or U2400 (N_2400,N_385,N_779);
nor U2401 (N_2401,N_1070,N_1325);
xnor U2402 (N_2402,N_19,N_767);
and U2403 (N_2403,N_1384,N_611);
nand U2404 (N_2404,N_109,N_1321);
nor U2405 (N_2405,N_680,N_187);
and U2406 (N_2406,N_970,N_329);
xor U2407 (N_2407,N_1440,N_780);
nand U2408 (N_2408,N_579,N_518);
nand U2409 (N_2409,N_114,N_1068);
nor U2410 (N_2410,N_922,N_608);
or U2411 (N_2411,N_1271,N_878);
xor U2412 (N_2412,N_337,N_585);
and U2413 (N_2413,N_498,N_106);
or U2414 (N_2414,N_312,N_1358);
nor U2415 (N_2415,N_444,N_486);
or U2416 (N_2416,N_1131,N_527);
nand U2417 (N_2417,N_213,N_1103);
or U2418 (N_2418,N_762,N_738);
xor U2419 (N_2419,N_1262,N_1486);
or U2420 (N_2420,N_318,N_805);
or U2421 (N_2421,N_999,N_1446);
nor U2422 (N_2422,N_423,N_364);
and U2423 (N_2423,N_515,N_933);
and U2424 (N_2424,N_5,N_1181);
nor U2425 (N_2425,N_142,N_205);
and U2426 (N_2426,N_966,N_604);
nor U2427 (N_2427,N_487,N_927);
nand U2428 (N_2428,N_557,N_1471);
nor U2429 (N_2429,N_1154,N_965);
nor U2430 (N_2430,N_101,N_636);
and U2431 (N_2431,N_139,N_1201);
or U2432 (N_2432,N_1426,N_752);
nand U2433 (N_2433,N_608,N_212);
nand U2434 (N_2434,N_1060,N_991);
and U2435 (N_2435,N_774,N_199);
or U2436 (N_2436,N_190,N_221);
nand U2437 (N_2437,N_273,N_1348);
nor U2438 (N_2438,N_510,N_1298);
nand U2439 (N_2439,N_1309,N_583);
and U2440 (N_2440,N_875,N_784);
xor U2441 (N_2441,N_857,N_396);
nand U2442 (N_2442,N_910,N_1366);
and U2443 (N_2443,N_56,N_1200);
and U2444 (N_2444,N_1152,N_104);
and U2445 (N_2445,N_1175,N_778);
and U2446 (N_2446,N_365,N_620);
nor U2447 (N_2447,N_669,N_750);
or U2448 (N_2448,N_766,N_35);
xnor U2449 (N_2449,N_566,N_339);
nor U2450 (N_2450,N_901,N_1447);
or U2451 (N_2451,N_664,N_764);
or U2452 (N_2452,N_512,N_326);
nor U2453 (N_2453,N_253,N_1404);
nand U2454 (N_2454,N_441,N_519);
xnor U2455 (N_2455,N_742,N_17);
or U2456 (N_2456,N_878,N_503);
or U2457 (N_2457,N_518,N_123);
and U2458 (N_2458,N_1466,N_272);
nor U2459 (N_2459,N_875,N_1144);
nor U2460 (N_2460,N_332,N_1194);
nand U2461 (N_2461,N_959,N_657);
and U2462 (N_2462,N_75,N_783);
nand U2463 (N_2463,N_374,N_496);
nor U2464 (N_2464,N_976,N_426);
nor U2465 (N_2465,N_1214,N_166);
nor U2466 (N_2466,N_758,N_1072);
nand U2467 (N_2467,N_1373,N_792);
nor U2468 (N_2468,N_1114,N_1360);
or U2469 (N_2469,N_1430,N_1192);
nand U2470 (N_2470,N_1109,N_922);
and U2471 (N_2471,N_61,N_777);
or U2472 (N_2472,N_394,N_487);
or U2473 (N_2473,N_1235,N_1060);
xnor U2474 (N_2474,N_587,N_864);
nor U2475 (N_2475,N_887,N_976);
and U2476 (N_2476,N_661,N_316);
or U2477 (N_2477,N_1187,N_1420);
nand U2478 (N_2478,N_837,N_1413);
or U2479 (N_2479,N_1022,N_1278);
nor U2480 (N_2480,N_1428,N_1373);
or U2481 (N_2481,N_124,N_642);
or U2482 (N_2482,N_282,N_514);
and U2483 (N_2483,N_1454,N_1217);
or U2484 (N_2484,N_123,N_470);
xor U2485 (N_2485,N_938,N_891);
nor U2486 (N_2486,N_241,N_306);
or U2487 (N_2487,N_631,N_415);
nor U2488 (N_2488,N_502,N_1038);
xnor U2489 (N_2489,N_1269,N_889);
or U2490 (N_2490,N_1045,N_350);
and U2491 (N_2491,N_1303,N_972);
nor U2492 (N_2492,N_362,N_1434);
nor U2493 (N_2493,N_265,N_697);
nand U2494 (N_2494,N_580,N_731);
nor U2495 (N_2495,N_747,N_358);
nand U2496 (N_2496,N_1212,N_861);
or U2497 (N_2497,N_663,N_1236);
xnor U2498 (N_2498,N_267,N_393);
xnor U2499 (N_2499,N_1041,N_9);
or U2500 (N_2500,N_882,N_512);
nor U2501 (N_2501,N_655,N_1372);
xnor U2502 (N_2502,N_1184,N_263);
nand U2503 (N_2503,N_937,N_866);
nand U2504 (N_2504,N_101,N_336);
xnor U2505 (N_2505,N_452,N_426);
and U2506 (N_2506,N_1452,N_592);
xnor U2507 (N_2507,N_145,N_759);
or U2508 (N_2508,N_108,N_334);
or U2509 (N_2509,N_946,N_1200);
and U2510 (N_2510,N_103,N_1309);
or U2511 (N_2511,N_931,N_1055);
nor U2512 (N_2512,N_926,N_98);
xor U2513 (N_2513,N_996,N_310);
and U2514 (N_2514,N_339,N_404);
nand U2515 (N_2515,N_11,N_942);
and U2516 (N_2516,N_577,N_211);
or U2517 (N_2517,N_1240,N_1472);
or U2518 (N_2518,N_613,N_470);
and U2519 (N_2519,N_592,N_189);
and U2520 (N_2520,N_965,N_924);
nor U2521 (N_2521,N_1478,N_1342);
and U2522 (N_2522,N_579,N_465);
nand U2523 (N_2523,N_416,N_396);
or U2524 (N_2524,N_13,N_267);
and U2525 (N_2525,N_451,N_975);
or U2526 (N_2526,N_859,N_1042);
nor U2527 (N_2527,N_954,N_688);
and U2528 (N_2528,N_331,N_469);
or U2529 (N_2529,N_19,N_1157);
or U2530 (N_2530,N_754,N_1477);
nand U2531 (N_2531,N_118,N_567);
nand U2532 (N_2532,N_377,N_895);
or U2533 (N_2533,N_306,N_922);
xor U2534 (N_2534,N_1453,N_117);
xor U2535 (N_2535,N_1399,N_482);
nand U2536 (N_2536,N_46,N_946);
nand U2537 (N_2537,N_1050,N_1022);
and U2538 (N_2538,N_1292,N_1478);
nand U2539 (N_2539,N_625,N_254);
nor U2540 (N_2540,N_1026,N_1468);
or U2541 (N_2541,N_1034,N_633);
nor U2542 (N_2542,N_977,N_654);
and U2543 (N_2543,N_495,N_1091);
or U2544 (N_2544,N_477,N_94);
or U2545 (N_2545,N_421,N_835);
nor U2546 (N_2546,N_865,N_1229);
nor U2547 (N_2547,N_1142,N_778);
nor U2548 (N_2548,N_1166,N_1167);
nand U2549 (N_2549,N_1424,N_1389);
or U2550 (N_2550,N_1332,N_153);
or U2551 (N_2551,N_540,N_1337);
or U2552 (N_2552,N_989,N_620);
or U2553 (N_2553,N_245,N_772);
and U2554 (N_2554,N_51,N_1451);
nor U2555 (N_2555,N_379,N_1347);
or U2556 (N_2556,N_730,N_875);
or U2557 (N_2557,N_943,N_85);
or U2558 (N_2558,N_1254,N_477);
or U2559 (N_2559,N_1443,N_500);
and U2560 (N_2560,N_819,N_903);
or U2561 (N_2561,N_920,N_671);
or U2562 (N_2562,N_818,N_507);
or U2563 (N_2563,N_57,N_1433);
or U2564 (N_2564,N_636,N_792);
xor U2565 (N_2565,N_814,N_560);
or U2566 (N_2566,N_366,N_182);
or U2567 (N_2567,N_1351,N_411);
nand U2568 (N_2568,N_664,N_796);
or U2569 (N_2569,N_1491,N_976);
xnor U2570 (N_2570,N_1219,N_430);
or U2571 (N_2571,N_325,N_1479);
xnor U2572 (N_2572,N_1463,N_129);
and U2573 (N_2573,N_869,N_140);
nand U2574 (N_2574,N_889,N_731);
nor U2575 (N_2575,N_1113,N_45);
nand U2576 (N_2576,N_114,N_1073);
and U2577 (N_2577,N_1065,N_1153);
and U2578 (N_2578,N_1472,N_1467);
nor U2579 (N_2579,N_673,N_1080);
and U2580 (N_2580,N_328,N_488);
nand U2581 (N_2581,N_1221,N_476);
and U2582 (N_2582,N_861,N_783);
nor U2583 (N_2583,N_1222,N_16);
nor U2584 (N_2584,N_243,N_1486);
nand U2585 (N_2585,N_899,N_857);
or U2586 (N_2586,N_20,N_54);
or U2587 (N_2587,N_254,N_59);
or U2588 (N_2588,N_882,N_1437);
or U2589 (N_2589,N_390,N_894);
or U2590 (N_2590,N_458,N_1363);
and U2591 (N_2591,N_307,N_655);
nand U2592 (N_2592,N_826,N_1285);
nor U2593 (N_2593,N_909,N_1474);
or U2594 (N_2594,N_977,N_647);
nand U2595 (N_2595,N_1241,N_725);
or U2596 (N_2596,N_880,N_940);
xor U2597 (N_2597,N_785,N_1451);
xor U2598 (N_2598,N_1418,N_1);
or U2599 (N_2599,N_1237,N_823);
and U2600 (N_2600,N_210,N_413);
xor U2601 (N_2601,N_934,N_1323);
and U2602 (N_2602,N_1432,N_508);
or U2603 (N_2603,N_865,N_1036);
nand U2604 (N_2604,N_192,N_249);
nand U2605 (N_2605,N_1170,N_113);
xnor U2606 (N_2606,N_736,N_527);
or U2607 (N_2607,N_503,N_475);
nor U2608 (N_2608,N_1325,N_955);
nor U2609 (N_2609,N_712,N_154);
nand U2610 (N_2610,N_5,N_504);
and U2611 (N_2611,N_546,N_742);
nand U2612 (N_2612,N_623,N_521);
nor U2613 (N_2613,N_174,N_934);
nand U2614 (N_2614,N_469,N_40);
or U2615 (N_2615,N_263,N_462);
and U2616 (N_2616,N_926,N_998);
nand U2617 (N_2617,N_1337,N_820);
nand U2618 (N_2618,N_1126,N_343);
nor U2619 (N_2619,N_1382,N_820);
or U2620 (N_2620,N_346,N_1057);
nor U2621 (N_2621,N_655,N_119);
nand U2622 (N_2622,N_958,N_1082);
nor U2623 (N_2623,N_650,N_144);
nor U2624 (N_2624,N_296,N_556);
nor U2625 (N_2625,N_1491,N_708);
nand U2626 (N_2626,N_771,N_1326);
or U2627 (N_2627,N_170,N_497);
nand U2628 (N_2628,N_746,N_258);
xnor U2629 (N_2629,N_681,N_1412);
nand U2630 (N_2630,N_636,N_1057);
and U2631 (N_2631,N_1045,N_955);
nor U2632 (N_2632,N_1466,N_884);
nand U2633 (N_2633,N_70,N_554);
nand U2634 (N_2634,N_489,N_852);
nor U2635 (N_2635,N_697,N_56);
and U2636 (N_2636,N_1128,N_565);
nand U2637 (N_2637,N_224,N_1322);
and U2638 (N_2638,N_1029,N_818);
or U2639 (N_2639,N_1339,N_1028);
or U2640 (N_2640,N_1434,N_1100);
nor U2641 (N_2641,N_1455,N_1452);
or U2642 (N_2642,N_1344,N_549);
or U2643 (N_2643,N_569,N_847);
nor U2644 (N_2644,N_1045,N_877);
or U2645 (N_2645,N_1061,N_1376);
and U2646 (N_2646,N_1235,N_673);
nand U2647 (N_2647,N_155,N_759);
xor U2648 (N_2648,N_622,N_1358);
nand U2649 (N_2649,N_1135,N_5);
or U2650 (N_2650,N_1255,N_484);
nor U2651 (N_2651,N_1462,N_1370);
nand U2652 (N_2652,N_1298,N_770);
and U2653 (N_2653,N_1376,N_807);
nand U2654 (N_2654,N_1043,N_262);
and U2655 (N_2655,N_1000,N_129);
or U2656 (N_2656,N_770,N_518);
xnor U2657 (N_2657,N_1246,N_1451);
or U2658 (N_2658,N_1471,N_955);
nor U2659 (N_2659,N_185,N_291);
and U2660 (N_2660,N_465,N_120);
nand U2661 (N_2661,N_1161,N_98);
and U2662 (N_2662,N_507,N_977);
xor U2663 (N_2663,N_849,N_1235);
nor U2664 (N_2664,N_264,N_191);
nand U2665 (N_2665,N_1138,N_632);
xor U2666 (N_2666,N_970,N_1457);
and U2667 (N_2667,N_583,N_644);
or U2668 (N_2668,N_723,N_688);
nand U2669 (N_2669,N_738,N_580);
and U2670 (N_2670,N_900,N_726);
and U2671 (N_2671,N_1080,N_871);
or U2672 (N_2672,N_748,N_76);
and U2673 (N_2673,N_73,N_908);
nand U2674 (N_2674,N_975,N_596);
and U2675 (N_2675,N_612,N_1401);
nor U2676 (N_2676,N_217,N_1454);
nand U2677 (N_2677,N_834,N_637);
or U2678 (N_2678,N_963,N_414);
nand U2679 (N_2679,N_628,N_172);
nor U2680 (N_2680,N_779,N_907);
nor U2681 (N_2681,N_714,N_564);
nand U2682 (N_2682,N_1168,N_885);
nand U2683 (N_2683,N_501,N_416);
xnor U2684 (N_2684,N_570,N_428);
and U2685 (N_2685,N_81,N_329);
nor U2686 (N_2686,N_1337,N_732);
nor U2687 (N_2687,N_243,N_1345);
and U2688 (N_2688,N_315,N_303);
and U2689 (N_2689,N_452,N_1466);
or U2690 (N_2690,N_1290,N_755);
and U2691 (N_2691,N_69,N_678);
and U2692 (N_2692,N_1101,N_787);
nand U2693 (N_2693,N_16,N_1495);
and U2694 (N_2694,N_1388,N_1453);
and U2695 (N_2695,N_973,N_1091);
xnor U2696 (N_2696,N_676,N_715);
nand U2697 (N_2697,N_811,N_754);
and U2698 (N_2698,N_2,N_880);
xor U2699 (N_2699,N_1357,N_622);
nor U2700 (N_2700,N_1385,N_148);
and U2701 (N_2701,N_635,N_1484);
and U2702 (N_2702,N_145,N_1210);
nand U2703 (N_2703,N_281,N_1161);
nand U2704 (N_2704,N_1182,N_389);
and U2705 (N_2705,N_629,N_818);
and U2706 (N_2706,N_390,N_1152);
or U2707 (N_2707,N_1331,N_364);
nand U2708 (N_2708,N_68,N_843);
or U2709 (N_2709,N_1448,N_323);
nor U2710 (N_2710,N_563,N_989);
nand U2711 (N_2711,N_1388,N_701);
xor U2712 (N_2712,N_1006,N_496);
or U2713 (N_2713,N_87,N_1284);
and U2714 (N_2714,N_719,N_180);
xnor U2715 (N_2715,N_395,N_251);
and U2716 (N_2716,N_287,N_973);
and U2717 (N_2717,N_676,N_76);
and U2718 (N_2718,N_1253,N_442);
or U2719 (N_2719,N_1318,N_761);
or U2720 (N_2720,N_216,N_876);
or U2721 (N_2721,N_1087,N_616);
and U2722 (N_2722,N_239,N_797);
nand U2723 (N_2723,N_1249,N_596);
nand U2724 (N_2724,N_1417,N_667);
and U2725 (N_2725,N_1061,N_1423);
and U2726 (N_2726,N_1278,N_537);
or U2727 (N_2727,N_202,N_634);
nand U2728 (N_2728,N_938,N_211);
or U2729 (N_2729,N_1462,N_114);
nand U2730 (N_2730,N_465,N_1341);
nor U2731 (N_2731,N_423,N_249);
xnor U2732 (N_2732,N_95,N_409);
nor U2733 (N_2733,N_101,N_397);
nand U2734 (N_2734,N_1154,N_1315);
nand U2735 (N_2735,N_74,N_566);
nand U2736 (N_2736,N_1260,N_1126);
and U2737 (N_2737,N_1003,N_640);
nor U2738 (N_2738,N_61,N_1162);
or U2739 (N_2739,N_1304,N_237);
and U2740 (N_2740,N_49,N_1151);
and U2741 (N_2741,N_770,N_459);
or U2742 (N_2742,N_1398,N_1203);
nor U2743 (N_2743,N_745,N_970);
nand U2744 (N_2744,N_352,N_1383);
nand U2745 (N_2745,N_266,N_166);
or U2746 (N_2746,N_322,N_1433);
nor U2747 (N_2747,N_989,N_631);
nand U2748 (N_2748,N_912,N_465);
and U2749 (N_2749,N_885,N_104);
xnor U2750 (N_2750,N_369,N_193);
and U2751 (N_2751,N_271,N_728);
or U2752 (N_2752,N_1432,N_772);
or U2753 (N_2753,N_1348,N_949);
and U2754 (N_2754,N_450,N_56);
nor U2755 (N_2755,N_1166,N_694);
or U2756 (N_2756,N_1294,N_1201);
nand U2757 (N_2757,N_944,N_58);
and U2758 (N_2758,N_1455,N_526);
nor U2759 (N_2759,N_147,N_512);
or U2760 (N_2760,N_926,N_1064);
nor U2761 (N_2761,N_28,N_1103);
and U2762 (N_2762,N_122,N_63);
or U2763 (N_2763,N_253,N_400);
or U2764 (N_2764,N_1152,N_623);
nand U2765 (N_2765,N_46,N_171);
nor U2766 (N_2766,N_86,N_111);
nand U2767 (N_2767,N_1152,N_571);
nor U2768 (N_2768,N_554,N_1166);
or U2769 (N_2769,N_1489,N_34);
and U2770 (N_2770,N_481,N_659);
nor U2771 (N_2771,N_602,N_905);
nand U2772 (N_2772,N_1,N_1332);
nor U2773 (N_2773,N_629,N_834);
nand U2774 (N_2774,N_420,N_561);
nand U2775 (N_2775,N_1219,N_1118);
or U2776 (N_2776,N_785,N_1134);
xnor U2777 (N_2777,N_382,N_44);
and U2778 (N_2778,N_435,N_58);
nor U2779 (N_2779,N_110,N_287);
nor U2780 (N_2780,N_368,N_97);
nor U2781 (N_2781,N_883,N_764);
nor U2782 (N_2782,N_481,N_496);
and U2783 (N_2783,N_635,N_289);
nand U2784 (N_2784,N_127,N_1063);
nor U2785 (N_2785,N_1481,N_742);
nand U2786 (N_2786,N_46,N_136);
nor U2787 (N_2787,N_698,N_1387);
xnor U2788 (N_2788,N_1139,N_183);
or U2789 (N_2789,N_775,N_1232);
nor U2790 (N_2790,N_651,N_475);
or U2791 (N_2791,N_1296,N_825);
or U2792 (N_2792,N_279,N_692);
nand U2793 (N_2793,N_110,N_1369);
nand U2794 (N_2794,N_1015,N_1387);
xnor U2795 (N_2795,N_852,N_238);
and U2796 (N_2796,N_944,N_124);
and U2797 (N_2797,N_313,N_470);
and U2798 (N_2798,N_363,N_1161);
nand U2799 (N_2799,N_1377,N_42);
or U2800 (N_2800,N_9,N_1474);
or U2801 (N_2801,N_1299,N_361);
nand U2802 (N_2802,N_857,N_1421);
nor U2803 (N_2803,N_42,N_280);
or U2804 (N_2804,N_777,N_578);
nand U2805 (N_2805,N_457,N_1261);
nor U2806 (N_2806,N_1131,N_586);
nand U2807 (N_2807,N_89,N_1073);
and U2808 (N_2808,N_1110,N_1067);
or U2809 (N_2809,N_847,N_846);
or U2810 (N_2810,N_801,N_1205);
and U2811 (N_2811,N_1100,N_966);
and U2812 (N_2812,N_1326,N_1488);
or U2813 (N_2813,N_1415,N_369);
nor U2814 (N_2814,N_817,N_1246);
and U2815 (N_2815,N_1163,N_491);
xnor U2816 (N_2816,N_575,N_774);
and U2817 (N_2817,N_818,N_524);
xor U2818 (N_2818,N_857,N_327);
nand U2819 (N_2819,N_312,N_760);
nand U2820 (N_2820,N_303,N_495);
and U2821 (N_2821,N_1358,N_765);
and U2822 (N_2822,N_1193,N_686);
and U2823 (N_2823,N_800,N_899);
and U2824 (N_2824,N_632,N_942);
and U2825 (N_2825,N_7,N_247);
and U2826 (N_2826,N_141,N_604);
nand U2827 (N_2827,N_76,N_486);
xnor U2828 (N_2828,N_797,N_275);
or U2829 (N_2829,N_385,N_923);
or U2830 (N_2830,N_668,N_111);
nand U2831 (N_2831,N_1399,N_1236);
and U2832 (N_2832,N_604,N_1311);
nand U2833 (N_2833,N_311,N_1449);
or U2834 (N_2834,N_857,N_1021);
nor U2835 (N_2835,N_257,N_970);
nor U2836 (N_2836,N_1043,N_74);
and U2837 (N_2837,N_823,N_304);
and U2838 (N_2838,N_477,N_844);
nor U2839 (N_2839,N_546,N_91);
nand U2840 (N_2840,N_4,N_600);
xor U2841 (N_2841,N_1291,N_1184);
or U2842 (N_2842,N_1111,N_457);
or U2843 (N_2843,N_462,N_248);
and U2844 (N_2844,N_1195,N_1472);
nor U2845 (N_2845,N_1467,N_425);
nor U2846 (N_2846,N_21,N_623);
or U2847 (N_2847,N_642,N_743);
nor U2848 (N_2848,N_409,N_146);
nand U2849 (N_2849,N_681,N_885);
and U2850 (N_2850,N_1101,N_1375);
nand U2851 (N_2851,N_621,N_289);
nor U2852 (N_2852,N_535,N_151);
nand U2853 (N_2853,N_553,N_1056);
nor U2854 (N_2854,N_85,N_288);
or U2855 (N_2855,N_83,N_944);
xnor U2856 (N_2856,N_670,N_794);
or U2857 (N_2857,N_1209,N_1333);
or U2858 (N_2858,N_899,N_301);
and U2859 (N_2859,N_355,N_1053);
and U2860 (N_2860,N_1327,N_226);
xor U2861 (N_2861,N_768,N_1481);
nor U2862 (N_2862,N_673,N_417);
nand U2863 (N_2863,N_884,N_1372);
nand U2864 (N_2864,N_1160,N_38);
and U2865 (N_2865,N_743,N_1308);
nor U2866 (N_2866,N_1112,N_1101);
or U2867 (N_2867,N_964,N_572);
or U2868 (N_2868,N_1299,N_334);
and U2869 (N_2869,N_331,N_283);
and U2870 (N_2870,N_1403,N_614);
nand U2871 (N_2871,N_402,N_1007);
nor U2872 (N_2872,N_309,N_1354);
nor U2873 (N_2873,N_692,N_300);
nor U2874 (N_2874,N_1408,N_1306);
nor U2875 (N_2875,N_1221,N_434);
nand U2876 (N_2876,N_1409,N_1440);
or U2877 (N_2877,N_791,N_311);
and U2878 (N_2878,N_588,N_613);
nand U2879 (N_2879,N_1391,N_939);
xor U2880 (N_2880,N_1068,N_1271);
and U2881 (N_2881,N_114,N_1373);
and U2882 (N_2882,N_175,N_908);
and U2883 (N_2883,N_65,N_427);
nand U2884 (N_2884,N_1471,N_571);
and U2885 (N_2885,N_1210,N_1419);
nor U2886 (N_2886,N_1070,N_725);
nand U2887 (N_2887,N_707,N_1421);
nor U2888 (N_2888,N_1422,N_919);
nand U2889 (N_2889,N_1157,N_317);
nand U2890 (N_2890,N_878,N_637);
nand U2891 (N_2891,N_682,N_24);
nor U2892 (N_2892,N_829,N_196);
nand U2893 (N_2893,N_1420,N_339);
nand U2894 (N_2894,N_309,N_708);
nand U2895 (N_2895,N_1339,N_111);
nor U2896 (N_2896,N_161,N_496);
nor U2897 (N_2897,N_563,N_983);
or U2898 (N_2898,N_1202,N_1125);
nor U2899 (N_2899,N_603,N_915);
nand U2900 (N_2900,N_296,N_54);
nand U2901 (N_2901,N_495,N_726);
or U2902 (N_2902,N_1239,N_544);
nor U2903 (N_2903,N_836,N_1145);
or U2904 (N_2904,N_114,N_213);
or U2905 (N_2905,N_1208,N_616);
nor U2906 (N_2906,N_685,N_656);
and U2907 (N_2907,N_25,N_1490);
nand U2908 (N_2908,N_141,N_981);
or U2909 (N_2909,N_107,N_248);
xor U2910 (N_2910,N_37,N_1073);
and U2911 (N_2911,N_899,N_226);
and U2912 (N_2912,N_279,N_231);
nor U2913 (N_2913,N_64,N_985);
nor U2914 (N_2914,N_1122,N_376);
or U2915 (N_2915,N_1158,N_394);
nor U2916 (N_2916,N_787,N_123);
and U2917 (N_2917,N_291,N_1263);
or U2918 (N_2918,N_1151,N_64);
and U2919 (N_2919,N_1300,N_1114);
or U2920 (N_2920,N_670,N_748);
or U2921 (N_2921,N_565,N_1050);
nor U2922 (N_2922,N_917,N_1350);
nand U2923 (N_2923,N_504,N_524);
or U2924 (N_2924,N_948,N_545);
or U2925 (N_2925,N_40,N_123);
nor U2926 (N_2926,N_45,N_483);
nor U2927 (N_2927,N_1225,N_1317);
and U2928 (N_2928,N_1361,N_532);
nand U2929 (N_2929,N_1248,N_1097);
nor U2930 (N_2930,N_409,N_1341);
xor U2931 (N_2931,N_916,N_541);
and U2932 (N_2932,N_1174,N_901);
and U2933 (N_2933,N_759,N_162);
nand U2934 (N_2934,N_1347,N_164);
nor U2935 (N_2935,N_671,N_1083);
and U2936 (N_2936,N_1240,N_239);
nand U2937 (N_2937,N_1104,N_1274);
and U2938 (N_2938,N_591,N_421);
nor U2939 (N_2939,N_43,N_354);
nand U2940 (N_2940,N_633,N_1137);
nor U2941 (N_2941,N_1033,N_868);
nand U2942 (N_2942,N_93,N_1366);
and U2943 (N_2943,N_418,N_138);
nor U2944 (N_2944,N_600,N_704);
xnor U2945 (N_2945,N_85,N_24);
and U2946 (N_2946,N_766,N_1235);
nor U2947 (N_2947,N_4,N_717);
or U2948 (N_2948,N_71,N_615);
nand U2949 (N_2949,N_750,N_336);
nor U2950 (N_2950,N_200,N_1155);
and U2951 (N_2951,N_1145,N_1461);
or U2952 (N_2952,N_782,N_1174);
and U2953 (N_2953,N_661,N_504);
or U2954 (N_2954,N_826,N_28);
and U2955 (N_2955,N_1389,N_1317);
and U2956 (N_2956,N_1163,N_1338);
nand U2957 (N_2957,N_852,N_81);
or U2958 (N_2958,N_1196,N_831);
nand U2959 (N_2959,N_513,N_1275);
nor U2960 (N_2960,N_592,N_734);
xnor U2961 (N_2961,N_1291,N_16);
and U2962 (N_2962,N_370,N_67);
xnor U2963 (N_2963,N_559,N_700);
nor U2964 (N_2964,N_190,N_777);
or U2965 (N_2965,N_1454,N_223);
and U2966 (N_2966,N_1189,N_1015);
and U2967 (N_2967,N_1128,N_145);
xor U2968 (N_2968,N_1107,N_1073);
and U2969 (N_2969,N_49,N_713);
nand U2970 (N_2970,N_1060,N_857);
xnor U2971 (N_2971,N_607,N_1090);
nand U2972 (N_2972,N_1104,N_826);
nor U2973 (N_2973,N_1269,N_276);
xnor U2974 (N_2974,N_166,N_65);
nor U2975 (N_2975,N_752,N_1153);
and U2976 (N_2976,N_1114,N_130);
nor U2977 (N_2977,N_944,N_1240);
xor U2978 (N_2978,N_668,N_1197);
and U2979 (N_2979,N_834,N_308);
nor U2980 (N_2980,N_761,N_883);
xor U2981 (N_2981,N_124,N_42);
nand U2982 (N_2982,N_1417,N_717);
nor U2983 (N_2983,N_919,N_209);
nor U2984 (N_2984,N_1456,N_1113);
nand U2985 (N_2985,N_1287,N_1129);
and U2986 (N_2986,N_1456,N_261);
xor U2987 (N_2987,N_1214,N_78);
nand U2988 (N_2988,N_886,N_1014);
and U2989 (N_2989,N_546,N_187);
and U2990 (N_2990,N_981,N_785);
nor U2991 (N_2991,N_1409,N_758);
and U2992 (N_2992,N_1105,N_475);
nor U2993 (N_2993,N_181,N_407);
and U2994 (N_2994,N_1195,N_402);
xnor U2995 (N_2995,N_618,N_1186);
nand U2996 (N_2996,N_1263,N_195);
nand U2997 (N_2997,N_996,N_197);
or U2998 (N_2998,N_1147,N_445);
nor U2999 (N_2999,N_615,N_1466);
nor U3000 (N_3000,N_2832,N_2968);
nor U3001 (N_3001,N_1659,N_2355);
and U3002 (N_3002,N_2530,N_1935);
nand U3003 (N_3003,N_1875,N_2063);
and U3004 (N_3004,N_1547,N_2563);
xnor U3005 (N_3005,N_2744,N_2792);
xnor U3006 (N_3006,N_1534,N_1780);
and U3007 (N_3007,N_1689,N_2922);
nor U3008 (N_3008,N_1690,N_2948);
nand U3009 (N_3009,N_1785,N_2532);
nor U3010 (N_3010,N_2011,N_2859);
and U3011 (N_3011,N_1632,N_1900);
and U3012 (N_3012,N_1673,N_1643);
nor U3013 (N_3013,N_2220,N_1624);
nand U3014 (N_3014,N_2136,N_2880);
and U3015 (N_3015,N_1837,N_1969);
nand U3016 (N_3016,N_2644,N_2902);
or U3017 (N_3017,N_1599,N_2677);
and U3018 (N_3018,N_2152,N_2358);
and U3019 (N_3019,N_2335,N_2754);
nor U3020 (N_3020,N_2997,N_1866);
nand U3021 (N_3021,N_1561,N_2021);
xnor U3022 (N_3022,N_2056,N_2099);
nor U3023 (N_3023,N_2651,N_2264);
nor U3024 (N_3024,N_2764,N_2741);
nand U3025 (N_3025,N_2830,N_2248);
or U3026 (N_3026,N_1579,N_2661);
nor U3027 (N_3027,N_2680,N_2747);
and U3028 (N_3028,N_2267,N_2628);
nand U3029 (N_3029,N_1538,N_1545);
nor U3030 (N_3030,N_2779,N_2894);
nand U3031 (N_3031,N_2102,N_2391);
or U3032 (N_3032,N_1899,N_2175);
and U3033 (N_3033,N_2447,N_2582);
xor U3034 (N_3034,N_1539,N_2460);
nor U3035 (N_3035,N_2124,N_2929);
nand U3036 (N_3036,N_2983,N_1505);
and U3037 (N_3037,N_1551,N_2345);
nand U3038 (N_3038,N_2446,N_2996);
xor U3039 (N_3039,N_2611,N_2521);
nand U3040 (N_3040,N_2626,N_2994);
or U3041 (N_3041,N_2957,N_2573);
nand U3042 (N_3042,N_2024,N_1711);
nand U3043 (N_3043,N_1628,N_2203);
nand U3044 (N_3044,N_1881,N_2614);
nand U3045 (N_3045,N_1509,N_2616);
nor U3046 (N_3046,N_1773,N_1824);
xor U3047 (N_3047,N_2462,N_2486);
nand U3048 (N_3048,N_1989,N_2960);
and U3049 (N_3049,N_2972,N_1640);
xor U3050 (N_3050,N_1993,N_2468);
nor U3051 (N_3051,N_2535,N_2854);
nand U3052 (N_3052,N_2751,N_2827);
or U3053 (N_3053,N_2978,N_2890);
and U3054 (N_3054,N_1915,N_2726);
nand U3055 (N_3055,N_2674,N_2520);
nor U3056 (N_3056,N_2459,N_1590);
and U3057 (N_3057,N_2867,N_2129);
and U3058 (N_3058,N_1734,N_1829);
nand U3059 (N_3059,N_2705,N_2756);
nand U3060 (N_3060,N_2128,N_2042);
and U3061 (N_3061,N_2720,N_2898);
nor U3062 (N_3062,N_2163,N_2612);
or U3063 (N_3063,N_2541,N_1654);
nand U3064 (N_3064,N_2966,N_2742);
nor U3065 (N_3065,N_2495,N_2185);
nor U3066 (N_3066,N_2760,N_2740);
nand U3067 (N_3067,N_1582,N_1563);
nor U3068 (N_3068,N_1980,N_1691);
nand U3069 (N_3069,N_2947,N_2246);
and U3070 (N_3070,N_1774,N_2667);
and U3071 (N_3071,N_1905,N_2334);
nand U3072 (N_3072,N_1975,N_2800);
and U3073 (N_3073,N_2875,N_2234);
or U3074 (N_3074,N_2378,N_2695);
and U3075 (N_3075,N_2684,N_2593);
xor U3076 (N_3076,N_2017,N_2080);
or U3077 (N_3077,N_2539,N_2901);
xor U3078 (N_3078,N_2002,N_2869);
nor U3079 (N_3079,N_2725,N_2911);
nor U3080 (N_3080,N_1944,N_2167);
and U3081 (N_3081,N_2383,N_2610);
nor U3082 (N_3082,N_2399,N_1849);
and U3083 (N_3083,N_1750,N_2314);
or U3084 (N_3084,N_2157,N_2476);
or U3085 (N_3085,N_2835,N_1612);
nand U3086 (N_3086,N_2665,N_2602);
nand U3087 (N_3087,N_2696,N_2503);
and U3088 (N_3088,N_2138,N_1834);
nand U3089 (N_3089,N_2678,N_2496);
nor U3090 (N_3090,N_1788,N_2207);
and U3091 (N_3091,N_1816,N_1540);
nor U3092 (N_3092,N_1621,N_1648);
and U3093 (N_3093,N_1857,N_1922);
and U3094 (N_3094,N_2150,N_2638);
nor U3095 (N_3095,N_2955,N_2753);
and U3096 (N_3096,N_1603,N_2022);
nor U3097 (N_3097,N_2219,N_2064);
or U3098 (N_3098,N_2950,N_2082);
and U3099 (N_3099,N_1636,N_2689);
nand U3100 (N_3100,N_1737,N_1615);
nand U3101 (N_3101,N_1808,N_2111);
nor U3102 (N_3102,N_2261,N_2072);
or U3103 (N_3103,N_2373,N_2896);
nand U3104 (N_3104,N_1946,N_2904);
xnor U3105 (N_3105,N_2653,N_2804);
nor U3106 (N_3106,N_2778,N_1833);
nor U3107 (N_3107,N_2328,N_1665);
and U3108 (N_3108,N_2492,N_2572);
nor U3109 (N_3109,N_2096,N_2538);
nand U3110 (N_3110,N_2595,N_2518);
xor U3111 (N_3111,N_2192,N_2784);
and U3112 (N_3112,N_1928,N_2599);
xnor U3113 (N_3113,N_2162,N_1790);
or U3114 (N_3114,N_2088,N_1646);
nor U3115 (N_3115,N_2473,N_2502);
nor U3116 (N_3116,N_2629,N_2666);
nor U3117 (N_3117,N_2151,N_2389);
and U3118 (N_3118,N_2853,N_1525);
xnor U3119 (N_3119,N_2078,N_1637);
xor U3120 (N_3120,N_1960,N_1838);
or U3121 (N_3121,N_2132,N_1544);
and U3122 (N_3122,N_2144,N_2316);
xor U3123 (N_3123,N_2304,N_1569);
nor U3124 (N_3124,N_1672,N_2380);
or U3125 (N_3125,N_2632,N_2103);
and U3126 (N_3126,N_2525,N_1543);
or U3127 (N_3127,N_2015,N_1508);
or U3128 (N_3128,N_1731,N_1642);
and U3129 (N_3129,N_2231,N_1766);
nor U3130 (N_3130,N_2286,N_2810);
nor U3131 (N_3131,N_2359,N_2750);
nand U3132 (N_3132,N_2336,N_2193);
nand U3133 (N_3133,N_2953,N_1608);
nand U3134 (N_3134,N_2449,N_2197);
nand U3135 (N_3135,N_2297,N_1645);
or U3136 (N_3136,N_2782,N_1797);
or U3137 (N_3137,N_2165,N_1822);
or U3138 (N_3138,N_1761,N_2196);
nor U3139 (N_3139,N_2243,N_2554);
nor U3140 (N_3140,N_2868,N_2937);
or U3141 (N_3141,N_2457,N_2637);
or U3142 (N_3142,N_1854,N_2509);
or U3143 (N_3143,N_2049,N_2499);
xnor U3144 (N_3144,N_2183,N_2608);
nand U3145 (N_3145,N_2475,N_1613);
nand U3146 (N_3146,N_2065,N_2850);
and U3147 (N_3147,N_1730,N_2491);
nand U3148 (N_3148,N_1681,N_2719);
and U3149 (N_3149,N_1572,N_1784);
nand U3150 (N_3150,N_1552,N_2642);
and U3151 (N_3151,N_2098,N_1864);
or U3152 (N_3152,N_1933,N_1943);
nand U3153 (N_3153,N_2101,N_2487);
nor U3154 (N_3154,N_2237,N_2069);
nor U3155 (N_3155,N_1717,N_2480);
nor U3156 (N_3156,N_2958,N_2250);
and U3157 (N_3157,N_2621,N_2673);
nor U3158 (N_3158,N_1546,N_2382);
nand U3159 (N_3159,N_2055,N_1977);
and U3160 (N_3160,N_1592,N_2117);
or U3161 (N_3161,N_1666,N_2092);
and U3162 (N_3162,N_1616,N_1846);
and U3163 (N_3163,N_1957,N_2836);
and U3164 (N_3164,N_2419,N_2450);
nand U3165 (N_3165,N_1853,N_2242);
and U3166 (N_3166,N_2766,N_1707);
or U3167 (N_3167,N_2870,N_2155);
and U3168 (N_3168,N_2565,N_2856);
xor U3169 (N_3169,N_1757,N_1815);
nor U3170 (N_3170,N_1671,N_2149);
nor U3171 (N_3171,N_2815,N_2706);
nor U3172 (N_3172,N_2845,N_1956);
nand U3173 (N_3173,N_2395,N_2893);
nor U3174 (N_3174,N_2083,N_2801);
nor U3175 (N_3175,N_2600,N_2494);
or U3176 (N_3176,N_2374,N_1502);
nor U3177 (N_3177,N_2089,N_2488);
nor U3178 (N_3178,N_2062,N_1716);
nor U3179 (N_3179,N_1722,N_2370);
or U3180 (N_3180,N_2321,N_1804);
and U3181 (N_3181,N_1715,N_2523);
nor U3182 (N_3182,N_2592,N_1823);
and U3183 (N_3183,N_2936,N_1680);
nand U3184 (N_3184,N_2570,N_2732);
and U3185 (N_3185,N_2174,N_2161);
xnor U3186 (N_3186,N_2915,N_1655);
nor U3187 (N_3187,N_1658,N_2033);
nand U3188 (N_3188,N_2551,N_2453);
nand U3189 (N_3189,N_1775,N_2189);
nor U3190 (N_3190,N_1990,N_2657);
nand U3191 (N_3191,N_2356,N_2390);
nor U3192 (N_3192,N_1811,N_1500);
or U3193 (N_3193,N_2445,N_1634);
and U3194 (N_3194,N_2851,N_2195);
nor U3195 (N_3195,N_2385,N_2240);
nor U3196 (N_3196,N_2202,N_1503);
nor U3197 (N_3197,N_1760,N_2553);
xnor U3198 (N_3198,N_2817,N_2353);
xor U3199 (N_3199,N_2709,N_2458);
or U3200 (N_3200,N_2077,N_2262);
or U3201 (N_3201,N_1988,N_2405);
nand U3202 (N_3202,N_2109,N_1562);
nand U3203 (N_3203,N_1950,N_2591);
or U3204 (N_3204,N_2692,N_2552);
and U3205 (N_3205,N_1511,N_2012);
xor U3206 (N_3206,N_1868,N_2364);
xnor U3207 (N_3207,N_1852,N_2333);
nor U3208 (N_3208,N_1515,N_2041);
nor U3209 (N_3209,N_1553,N_2107);
and U3210 (N_3210,N_1937,N_2464);
nor U3211 (N_3211,N_2376,N_1639);
or U3212 (N_3212,N_1945,N_2338);
nand U3213 (N_3213,N_1979,N_2433);
xor U3214 (N_3214,N_1843,N_2545);
or U3215 (N_3215,N_2799,N_2230);
or U3216 (N_3216,N_1991,N_1754);
nor U3217 (N_3217,N_2694,N_1926);
nand U3218 (N_3218,N_2342,N_1588);
nand U3219 (N_3219,N_2319,N_2886);
or U3220 (N_3220,N_2609,N_2131);
nor U3221 (N_3221,N_2797,N_1759);
nor U3222 (N_3222,N_2933,N_1949);
or U3223 (N_3223,N_1651,N_2580);
or U3224 (N_3224,N_1878,N_2635);
and U3225 (N_3225,N_1941,N_2897);
nand U3226 (N_3226,N_2420,N_2299);
xor U3227 (N_3227,N_1657,N_2474);
xnor U3228 (N_3228,N_2914,N_2825);
nand U3229 (N_3229,N_1530,N_1598);
nor U3230 (N_3230,N_1869,N_1894);
xor U3231 (N_3231,N_2222,N_1647);
nor U3232 (N_3232,N_2806,N_2302);
nor U3233 (N_3233,N_2723,N_2618);
nor U3234 (N_3234,N_2998,N_1653);
nor U3235 (N_3235,N_2829,N_1898);
nand U3236 (N_3236,N_1695,N_2871);
and U3237 (N_3237,N_2170,N_2498);
nor U3238 (N_3238,N_1524,N_2278);
nor U3239 (N_3239,N_2104,N_1789);
xor U3240 (N_3240,N_2985,N_2921);
nor U3241 (N_3241,N_1676,N_1510);
nor U3242 (N_3242,N_2884,N_2989);
or U3243 (N_3243,N_2030,N_2895);
nor U3244 (N_3244,N_1669,N_2605);
and U3245 (N_3245,N_2993,N_2862);
nand U3246 (N_3246,N_2187,N_2959);
nor U3247 (N_3247,N_1581,N_2841);
xnor U3248 (N_3248,N_2500,N_2350);
nor U3249 (N_3249,N_1858,N_2137);
or U3250 (N_3250,N_2479,N_1710);
xnor U3251 (N_3251,N_2965,N_2349);
nor U3252 (N_3252,N_2512,N_2838);
or U3253 (N_3253,N_2418,N_1606);
xnor U3254 (N_3254,N_2035,N_1519);
nor U3255 (N_3255,N_2351,N_2463);
nor U3256 (N_3256,N_2823,N_2014);
or U3257 (N_3257,N_2735,N_2718);
and U3258 (N_3258,N_2905,N_2354);
nand U3259 (N_3259,N_1549,N_2430);
xor U3260 (N_3260,N_2992,N_2566);
xor U3261 (N_3261,N_2690,N_2422);
and U3262 (N_3262,N_2038,N_1913);
nor U3263 (N_3263,N_2507,N_1924);
xor U3264 (N_3264,N_1693,N_2313);
or U3265 (N_3265,N_2180,N_1507);
nand U3266 (N_3266,N_2567,N_1968);
nor U3267 (N_3267,N_1587,N_2906);
nor U3268 (N_3268,N_1638,N_2141);
xnor U3269 (N_3269,N_2326,N_2006);
nand U3270 (N_3270,N_2415,N_2210);
or U3271 (N_3271,N_2171,N_2606);
nand U3272 (N_3272,N_1622,N_1840);
xnor U3273 (N_3273,N_2587,N_2847);
nand U3274 (N_3274,N_2544,N_1954);
nand U3275 (N_3275,N_2352,N_2279);
nand U3276 (N_3276,N_2483,N_2774);
or U3277 (N_3277,N_2848,N_2037);
nand U3278 (N_3278,N_2623,N_1712);
and U3279 (N_3279,N_1664,N_2622);
nand U3280 (N_3280,N_2182,N_1805);
nor U3281 (N_3281,N_1832,N_2659);
and U3282 (N_3282,N_2652,N_1863);
or U3283 (N_3283,N_1912,N_2821);
nand U3284 (N_3284,N_2110,N_1847);
nor U3285 (N_3285,N_1597,N_1802);
and U3286 (N_3286,N_2504,N_2036);
or U3287 (N_3287,N_2324,N_2467);
xor U3288 (N_3288,N_2477,N_1872);
nor U3289 (N_3289,N_2882,N_1542);
and U3290 (N_3290,N_2004,N_2687);
nor U3291 (N_3291,N_2057,N_1910);
nor U3292 (N_3292,N_1777,N_2771);
nand U3293 (N_3293,N_2394,N_2633);
nand U3294 (N_3294,N_1620,N_1981);
or U3295 (N_3295,N_2040,N_2236);
and U3296 (N_3296,N_1533,N_2400);
and U3297 (N_3297,N_2721,N_2999);
xor U3298 (N_3298,N_1541,N_2685);
nor U3299 (N_3299,N_2758,N_2414);
or U3300 (N_3300,N_1794,N_1874);
xnor U3301 (N_3301,N_1882,N_2942);
and U3302 (N_3302,N_2613,N_2100);
or U3303 (N_3303,N_1778,N_1674);
or U3304 (N_3304,N_2067,N_2927);
and U3305 (N_3305,N_2888,N_2232);
or U3306 (N_3306,N_2068,N_2013);
and U3307 (N_3307,N_2752,N_2925);
or U3308 (N_3308,N_1914,N_2146);
nand U3309 (N_3309,N_2786,N_1577);
xor U3310 (N_3310,N_2179,N_1629);
and U3311 (N_3311,N_1893,N_1678);
xnor U3312 (N_3312,N_1663,N_2497);
nand U3313 (N_3313,N_2408,N_2258);
nor U3314 (N_3314,N_2917,N_2931);
nand U3315 (N_3315,N_1535,N_2026);
or U3316 (N_3316,N_2926,N_2839);
or U3317 (N_3317,N_1818,N_1633);
nand U3318 (N_3318,N_2975,N_1504);
or U3319 (N_3319,N_2300,N_1756);
and U3320 (N_3320,N_2625,N_2048);
or U3321 (N_3321,N_2332,N_2700);
nand U3322 (N_3322,N_2974,N_1885);
nor U3323 (N_3323,N_2777,N_2537);
nor U3324 (N_3324,N_2003,N_2485);
or U3325 (N_3325,N_2007,N_2436);
nor U3326 (N_3326,N_1953,N_2676);
or U3327 (N_3327,N_1791,N_2987);
nor U3328 (N_3328,N_2118,N_1890);
nor U3329 (N_3329,N_2964,N_1527);
xnor U3330 (N_3330,N_1936,N_2416);
and U3331 (N_3331,N_2578,N_2791);
nand U3332 (N_3332,N_2670,N_1521);
nor U3333 (N_3333,N_2861,N_2995);
and U3334 (N_3334,N_1995,N_1531);
and U3335 (N_3335,N_2543,N_2619);
nor U3336 (N_3336,N_1744,N_2951);
or U3337 (N_3337,N_1770,N_1518);
or U3338 (N_3338,N_2401,N_1801);
or U3339 (N_3339,N_2780,N_1948);
nor U3340 (N_3340,N_2071,N_1512);
nor U3341 (N_3341,N_2424,N_1812);
nor U3342 (N_3342,N_1656,N_1548);
nor U3343 (N_3343,N_2233,N_1951);
nor U3344 (N_3344,N_2019,N_2688);
nor U3345 (N_3345,N_2820,N_2273);
xor U3346 (N_3346,N_1994,N_2548);
nand U3347 (N_3347,N_1558,N_1865);
or U3348 (N_3348,N_1699,N_1903);
or U3349 (N_3349,N_2770,N_2431);
nor U3350 (N_3350,N_1559,N_2181);
nor U3351 (N_3351,N_2051,N_2941);
nand U3352 (N_3352,N_2533,N_1571);
nand U3353 (N_3353,N_1880,N_2166);
or U3354 (N_3354,N_2075,N_1554);
and U3355 (N_3355,N_1595,N_2133);
xnor U3356 (N_3356,N_2112,N_1862);
nor U3357 (N_3357,N_1795,N_1850);
nor U3358 (N_3358,N_1618,N_2627);
or U3359 (N_3359,N_2158,N_2263);
or U3360 (N_3360,N_2768,N_2172);
or U3361 (N_3361,N_2793,N_1700);
xnor U3362 (N_3362,N_2361,N_1904);
xnor U3363 (N_3363,N_1746,N_1703);
or U3364 (N_3364,N_2887,N_2409);
nor U3365 (N_3365,N_1747,N_2268);
nand U3366 (N_3366,N_1641,N_2177);
nor U3367 (N_3367,N_2346,N_2298);
nand U3368 (N_3368,N_1568,N_1704);
or U3369 (N_3369,N_2643,N_1564);
nand U3370 (N_3370,N_2864,N_1723);
or U3371 (N_3371,N_2270,N_2675);
or U3372 (N_3372,N_1537,N_2191);
xnor U3373 (N_3373,N_2200,N_2034);
nor U3374 (N_3374,N_2369,N_1825);
nor U3375 (N_3375,N_2442,N_2879);
or U3376 (N_3376,N_2506,N_2227);
nand U3377 (N_3377,N_2224,N_2142);
xor U3378 (N_3378,N_2822,N_2682);
and U3379 (N_3379,N_2511,N_1826);
or U3380 (N_3380,N_1749,N_2287);
or U3381 (N_3381,N_2812,N_1842);
xor U3382 (N_3382,N_1844,N_1907);
nand U3383 (N_3383,N_2686,N_2074);
and U3384 (N_3384,N_2108,N_1961);
and U3385 (N_3385,N_1679,N_1803);
nand U3386 (N_3386,N_1614,N_2434);
or U3387 (N_3387,N_2814,N_2365);
xnor U3388 (N_3388,N_2586,N_2145);
and U3389 (N_3389,N_1719,N_1986);
xor U3390 (N_3390,N_1758,N_2818);
nand U3391 (N_3391,N_2954,N_1861);
and U3392 (N_3392,N_2315,N_2773);
nor U3393 (N_3393,N_1708,N_2226);
and U3394 (N_3394,N_2367,N_2106);
nor U3395 (N_3395,N_2844,N_2594);
and U3396 (N_3396,N_2765,N_2683);
nand U3397 (N_3397,N_2023,N_2148);
and U3398 (N_3398,N_1999,N_2935);
and U3399 (N_3399,N_2647,N_2976);
or U3400 (N_3400,N_1876,N_2546);
and U3401 (N_3401,N_2562,N_1983);
and U3402 (N_3402,N_2490,N_2788);
nand U3403 (N_3403,N_2199,N_2282);
or U3404 (N_3404,N_2245,N_1619);
nand U3405 (N_3405,N_1560,N_2481);
and U3406 (N_3406,N_2920,N_2849);
nand U3407 (N_3407,N_2748,N_2008);
xor U3408 (N_3408,N_2878,N_2428);
nor U3409 (N_3409,N_2484,N_2945);
nand U3410 (N_3410,N_2427,N_1817);
nor U3411 (N_3411,N_1532,N_2729);
xnor U3412 (N_3412,N_2501,N_2482);
or U3413 (N_3413,N_1567,N_2990);
and U3414 (N_3414,N_1520,N_2663);
and U3415 (N_3415,N_2009,N_2589);
nand U3416 (N_3416,N_1781,N_1660);
nand U3417 (N_3417,N_1729,N_2076);
or U3418 (N_3418,N_2962,N_2568);
nand U3419 (N_3419,N_2697,N_2411);
nor U3420 (N_3420,N_2872,N_2607);
or U3421 (N_3421,N_2769,N_2783);
xor U3422 (N_3422,N_2301,N_2113);
or U3423 (N_3423,N_2889,N_2842);
nand U3424 (N_3424,N_2930,N_1930);
nor U3425 (N_3425,N_1709,N_2432);
xor U3426 (N_3426,N_1902,N_2560);
or U3427 (N_3427,N_2824,N_2241);
or U3428 (N_3428,N_2981,N_1895);
xor U3429 (N_3429,N_2127,N_2259);
nor U3430 (N_3430,N_2636,N_1917);
nor U3431 (N_3431,N_2899,N_2362);
or U3432 (N_3432,N_1685,N_2239);
or U3433 (N_3433,N_2406,N_1809);
or U3434 (N_3434,N_2775,N_1600);
and U3435 (N_3435,N_1556,N_1783);
and U3436 (N_3436,N_2343,N_2603);
or U3437 (N_3437,N_2840,N_2249);
or U3438 (N_3438,N_2536,N_1997);
xnor U3439 (N_3439,N_1831,N_1786);
and U3440 (N_3440,N_1735,N_1896);
and U3441 (N_3441,N_2429,N_2455);
and U3442 (N_3442,N_2826,N_1740);
nand U3443 (N_3443,N_2846,N_2761);
nor U3444 (N_3444,N_1867,N_2357);
nand U3445 (N_3445,N_2216,N_1589);
and U3446 (N_3446,N_2253,N_2519);
nand U3447 (N_3447,N_2265,N_2341);
nor U3448 (N_3448,N_1574,N_1776);
nor U3449 (N_3449,N_2679,N_2646);
or U3450 (N_3450,N_2472,N_2918);
or U3451 (N_3451,N_1934,N_1884);
and U3452 (N_3452,N_2767,N_1819);
nand U3453 (N_3453,N_1630,N_1940);
nor U3454 (N_3454,N_2081,N_1771);
nor U3455 (N_3455,N_1738,N_1725);
xor U3456 (N_3456,N_2090,N_1984);
nand U3457 (N_3457,N_1836,N_2293);
and U3458 (N_3458,N_1557,N_1779);
or U3459 (N_3459,N_2423,N_2296);
nor U3460 (N_3460,N_2522,N_2816);
and U3461 (N_3461,N_2620,N_2097);
and U3462 (N_3462,N_2807,N_2542);
or U3463 (N_3463,N_2701,N_2513);
xnor U3464 (N_3464,N_2198,N_2215);
and U3465 (N_3465,N_2585,N_2303);
and U3466 (N_3466,N_1952,N_2309);
and U3467 (N_3467,N_2662,N_2787);
nor U3468 (N_3468,N_2808,N_2244);
xor U3469 (N_3469,N_2387,N_2514);
xnor U3470 (N_3470,N_1752,N_2439);
or U3471 (N_3471,N_1835,N_2274);
or U3472 (N_3472,N_2084,N_1967);
xnor U3473 (N_3473,N_2907,N_2714);
and U3474 (N_3474,N_2973,N_2208);
nand U3475 (N_3475,N_2311,N_2755);
nand U3476 (N_3476,N_2991,N_2698);
nor U3477 (N_3477,N_2883,N_2631);
nor U3478 (N_3478,N_2437,N_1701);
nor U3479 (N_3479,N_1586,N_2308);
or U3480 (N_3480,N_1570,N_2634);
nand U3481 (N_3481,N_1526,N_2704);
nand U3482 (N_3482,N_2272,N_1631);
and U3483 (N_3483,N_2122,N_2489);
and U3484 (N_3484,N_2223,N_1767);
nor U3485 (N_3485,N_2360,N_2288);
nor U3486 (N_3486,N_2079,N_1683);
nand U3487 (N_3487,N_1516,N_1684);
nor U3488 (N_3488,N_1787,N_1929);
and U3489 (N_3489,N_2256,N_2702);
or U3490 (N_3490,N_1886,N_2251);
and U3491 (N_3491,N_2443,N_1726);
and U3492 (N_3492,N_1923,N_2252);
nand U3493 (N_3493,N_1652,N_2178);
nand U3494 (N_3494,N_2798,N_2120);
and U3495 (N_3495,N_2440,N_1764);
or U3496 (N_3496,N_2596,N_2763);
and U3497 (N_3497,N_2577,N_1860);
nand U3498 (N_3498,N_2528,N_2323);
and U3499 (N_3499,N_2404,N_2255);
nand U3500 (N_3500,N_2329,N_2156);
nand U3501 (N_3501,N_1727,N_2703);
or U3502 (N_3502,N_1939,N_2873);
and U3503 (N_3503,N_1605,N_2348);
or U3504 (N_3504,N_1921,N_2205);
or U3505 (N_3505,N_1964,N_2866);
or U3506 (N_3506,N_2715,N_1743);
or U3507 (N_3507,N_2912,N_2949);
and U3508 (N_3508,N_2320,N_2837);
nand U3509 (N_3509,N_1649,N_1814);
and U3510 (N_3510,N_2734,N_2331);
nand U3511 (N_3511,N_2461,N_2159);
or U3512 (N_3512,N_2209,N_1827);
and U3513 (N_3513,N_2781,N_2052);
and U3514 (N_3514,N_1796,N_2843);
nor U3515 (N_3515,N_2691,N_2671);
nand U3516 (N_3516,N_1728,N_2368);
or U3517 (N_3517,N_1739,N_2441);
nor U3518 (N_3518,N_1611,N_2669);
nand U3519 (N_3519,N_2206,N_2087);
xor U3520 (N_3520,N_2561,N_2184);
xor U3521 (N_3521,N_2668,N_1959);
nand U3522 (N_3522,N_1536,N_2852);
or U3523 (N_3523,N_1602,N_2366);
xor U3524 (N_3524,N_1839,N_1974);
nand U3525 (N_3525,N_1845,N_1911);
nand U3526 (N_3526,N_2050,N_2834);
nor U3527 (N_3527,N_1798,N_1682);
nand U3528 (N_3528,N_2160,N_2564);
nor U3529 (N_3529,N_2271,N_2574);
and U3530 (N_3530,N_2053,N_1617);
or U3531 (N_3531,N_1765,N_2337);
nand U3532 (N_3532,N_2982,N_2307);
or U3533 (N_3533,N_2016,N_2276);
and U3534 (N_3534,N_2289,N_1987);
nor U3535 (N_3535,N_2010,N_1963);
nand U3536 (N_3536,N_2143,N_1751);
nand U3537 (N_3537,N_1670,N_2813);
nor U3538 (N_3538,N_2169,N_2970);
or U3539 (N_3539,N_2952,N_2295);
nor U3540 (N_3540,N_1585,N_2590);
or U3541 (N_3541,N_2325,N_1732);
xor U3542 (N_3542,N_1667,N_1573);
and U3543 (N_3543,N_2743,N_2785);
nor U3544 (N_3544,N_1978,N_2737);
and U3545 (N_3545,N_2280,N_2645);
nand U3546 (N_3546,N_1820,N_1856);
xnor U3547 (N_3547,N_2749,N_1593);
or U3548 (N_3548,N_2549,N_2534);
xor U3549 (N_3549,N_1870,N_1601);
xnor U3550 (N_3550,N_2527,N_2043);
and U3551 (N_3551,N_2738,N_2091);
or U3552 (N_3552,N_2713,N_2407);
xor U3553 (N_3553,N_2377,N_2386);
nand U3554 (N_3554,N_2794,N_2547);
nand U3555 (N_3555,N_2290,N_2550);
and U3556 (N_3556,N_2066,N_2860);
nor U3557 (N_3557,N_2858,N_2001);
nor U3558 (N_3558,N_1782,N_2005);
nor U3559 (N_3559,N_2517,N_2986);
nand U3560 (N_3560,N_1763,N_2292);
nor U3561 (N_3561,N_1768,N_1576);
or U3562 (N_3562,N_2044,N_2190);
or U3563 (N_3563,N_1938,N_2556);
nor U3564 (N_3564,N_2699,N_1821);
and U3565 (N_3565,N_2126,N_2803);
nor U3566 (N_3566,N_2865,N_1851);
nor U3567 (N_3567,N_1565,N_1799);
and U3568 (N_3568,N_2712,N_1748);
and U3569 (N_3569,N_1627,N_2515);
nand U3570 (N_3570,N_2371,N_1706);
and U3571 (N_3571,N_1566,N_2796);
or U3572 (N_3572,N_1800,N_2153);
and U3573 (N_3573,N_1887,N_1982);
nor U3574 (N_3574,N_1769,N_1909);
xnor U3575 (N_3575,N_2540,N_2649);
and U3576 (N_3576,N_2790,N_2617);
nor U3577 (N_3577,N_2655,N_1550);
nor U3578 (N_3578,N_2805,N_2397);
xnor U3579 (N_3579,N_2863,N_2967);
xnor U3580 (N_3580,N_2444,N_2641);
xnor U3581 (N_3581,N_2412,N_2648);
and U3582 (N_3582,N_2584,N_2508);
nand U3583 (N_3583,N_1908,N_1591);
or U3584 (N_3584,N_2093,N_2857);
or U3585 (N_3585,N_1692,N_2828);
nor U3586 (N_3586,N_2615,N_1916);
nand U3587 (N_3587,N_2294,N_1609);
nand U3588 (N_3588,N_2168,N_2588);
and U3589 (N_3589,N_1992,N_1879);
and U3590 (N_3590,N_2094,N_2254);
or U3591 (N_3591,N_2438,N_2940);
nand U3592 (N_3592,N_1897,N_2469);
and U3593 (N_3593,N_2330,N_2876);
nor U3594 (N_3594,N_2027,N_1931);
and U3595 (N_3595,N_2031,N_1555);
xnor U3596 (N_3596,N_2913,N_2123);
nor U3597 (N_3597,N_2392,N_1971);
nor U3598 (N_3598,N_1810,N_2891);
nor U3599 (N_3599,N_2347,N_2085);
nand U3600 (N_3600,N_1705,N_1918);
nor U3601 (N_3601,N_2597,N_2681);
nor U3602 (N_3602,N_2291,N_2213);
or U3603 (N_3603,N_2221,N_2322);
nand U3604 (N_3604,N_2581,N_1883);
or U3605 (N_3605,N_1919,N_2116);
nor U3606 (N_3606,N_1668,N_2928);
nand U3607 (N_3607,N_2448,N_1859);
nand U3608 (N_3608,N_1514,N_1635);
or U3609 (N_3609,N_2672,N_1976);
nor U3610 (N_3610,N_2710,N_1906);
nor U3611 (N_3611,N_2086,N_2025);
or U3612 (N_3612,N_2557,N_1947);
and U3613 (N_3613,N_1830,N_1714);
nor U3614 (N_3614,N_1650,N_1927);
or U3615 (N_3615,N_2154,N_2576);
and U3616 (N_3616,N_2526,N_2047);
nor U3617 (N_3617,N_2789,N_2885);
and U3618 (N_3618,N_2327,N_2961);
xnor U3619 (N_3619,N_2664,N_2963);
and U3620 (N_3620,N_1855,N_2257);
xor U3621 (N_3621,N_1688,N_2909);
and U3622 (N_3622,N_2121,N_1528);
nand U3623 (N_3623,N_1942,N_1755);
nand U3624 (N_3624,N_2795,N_2531);
xor U3625 (N_3625,N_2363,N_2266);
nand U3626 (N_3626,N_2139,N_2776);
nand U3627 (N_3627,N_2910,N_2946);
nand U3628 (N_3628,N_2939,N_1580);
nor U3629 (N_3629,N_2410,N_2114);
xnor U3630 (N_3630,N_1972,N_2658);
or U3631 (N_3631,N_1698,N_2140);
nand U3632 (N_3632,N_2529,N_2579);
nor U3633 (N_3633,N_2384,N_2656);
nand U3634 (N_3634,N_2654,N_2312);
nor U3635 (N_3635,N_1578,N_1575);
or U3636 (N_3636,N_2283,N_1607);
nor U3637 (N_3637,N_2717,N_1958);
and U3638 (N_3638,N_1807,N_2451);
nor U3639 (N_3639,N_2061,N_2235);
nor U3640 (N_3640,N_2173,N_2772);
nand U3641 (N_3641,N_2046,N_1529);
nand U3642 (N_3642,N_2381,N_1702);
nand U3643 (N_3643,N_2211,N_1662);
and U3644 (N_3644,N_2604,N_1848);
and U3645 (N_3645,N_2516,N_2029);
and U3646 (N_3646,N_2456,N_2650);
nand U3647 (N_3647,N_2711,N_2435);
nand U3648 (N_3648,N_2186,N_2938);
nor U3649 (N_3649,N_2934,N_1720);
nand U3650 (N_3650,N_2762,N_2733);
nor U3651 (N_3651,N_2317,N_2147);
nor U3652 (N_3652,N_1501,N_2730);
or U3653 (N_3653,N_2728,N_1873);
or U3654 (N_3654,N_2188,N_1686);
or U3655 (N_3655,N_2340,N_1522);
xor U3656 (N_3656,N_1762,N_2569);
xor U3657 (N_3657,N_2923,N_1891);
or U3658 (N_3658,N_1625,N_2130);
or U3659 (N_3659,N_2238,N_2707);
nand U3660 (N_3660,N_2969,N_1661);
nand U3661 (N_3661,N_1583,N_2214);
nand U3662 (N_3662,N_2212,N_1724);
and U3663 (N_3663,N_1584,N_2731);
nand U3664 (N_3664,N_2413,N_1925);
nor U3665 (N_3665,N_2465,N_1932);
nand U3666 (N_3666,N_1996,N_2454);
or U3667 (N_3667,N_2054,N_2125);
and U3668 (N_3668,N_2135,N_1753);
xor U3669 (N_3669,N_2217,N_1962);
nand U3670 (N_3670,N_2943,N_2831);
nand U3671 (N_3671,N_2285,N_2379);
xnor U3672 (N_3672,N_2372,N_2305);
nand U3673 (N_3673,N_1742,N_2559);
or U3674 (N_3674,N_2716,N_1506);
or U3675 (N_3675,N_2402,N_2903);
nand U3676 (N_3676,N_2470,N_2000);
nand U3677 (N_3677,N_2919,N_2524);
nand U3678 (N_3678,N_2575,N_1806);
and U3679 (N_3679,N_1718,N_1985);
nor U3680 (N_3680,N_1517,N_2493);
and U3681 (N_3681,N_2318,N_2045);
and U3682 (N_3682,N_2932,N_2059);
and U3683 (N_3683,N_2070,N_2693);
xnor U3684 (N_3684,N_2819,N_2275);
xnor U3685 (N_3685,N_1626,N_2624);
nand U3686 (N_3686,N_2944,N_2421);
nand U3687 (N_3687,N_1623,N_2058);
xor U3688 (N_3688,N_1687,N_2425);
nor U3689 (N_3689,N_2640,N_2281);
xor U3690 (N_3690,N_2979,N_2403);
nand U3691 (N_3691,N_2916,N_1694);
xor U3692 (N_3692,N_2727,N_1736);
xnor U3693 (N_3693,N_2977,N_2452);
nand U3694 (N_3694,N_2881,N_2375);
nor U3695 (N_3695,N_1889,N_2736);
and U3696 (N_3696,N_2510,N_2971);
nand U3697 (N_3697,N_2396,N_2176);
and U3698 (N_3698,N_2759,N_1973);
or U3699 (N_3699,N_2095,N_2228);
and U3700 (N_3700,N_1610,N_1675);
or U3701 (N_3701,N_2722,N_1644);
and U3702 (N_3702,N_2855,N_2583);
or U3703 (N_3703,N_2809,N_2339);
and U3704 (N_3704,N_1772,N_2204);
nand U3705 (N_3705,N_1888,N_2134);
and U3706 (N_3706,N_2892,N_1892);
or U3707 (N_3707,N_1792,N_2811);
nand U3708 (N_3708,N_2284,N_1955);
or U3709 (N_3709,N_2956,N_1965);
xnor U3710 (N_3710,N_2388,N_2988);
or U3711 (N_3711,N_2218,N_1877);
nor U3712 (N_3712,N_2225,N_1733);
nor U3713 (N_3713,N_2639,N_2060);
and U3714 (N_3714,N_1813,N_2471);
nand U3715 (N_3715,N_2194,N_1970);
xor U3716 (N_3716,N_2018,N_1696);
nor U3717 (N_3717,N_1596,N_2201);
nor U3718 (N_3718,N_2164,N_2708);
and U3719 (N_3719,N_1713,N_2032);
or U3720 (N_3720,N_2119,N_2398);
nand U3721 (N_3721,N_1677,N_2980);
nand U3722 (N_3722,N_2660,N_2020);
nand U3723 (N_3723,N_2306,N_2630);
nand U3724 (N_3724,N_2073,N_2555);
nand U3725 (N_3725,N_1828,N_1920);
or U3726 (N_3726,N_1998,N_1966);
or U3727 (N_3727,N_1604,N_2105);
or U3728 (N_3728,N_2571,N_2745);
nor U3729 (N_3729,N_2833,N_2877);
or U3730 (N_3730,N_1513,N_2984);
and U3731 (N_3731,N_1741,N_2802);
and U3732 (N_3732,N_2393,N_2277);
nor U3733 (N_3733,N_2039,N_2724);
and U3734 (N_3734,N_2310,N_1745);
or U3735 (N_3735,N_2260,N_2746);
nand U3736 (N_3736,N_1594,N_2115);
and U3737 (N_3737,N_2739,N_2757);
xnor U3738 (N_3738,N_2417,N_1793);
or U3739 (N_3739,N_1697,N_1871);
nand U3740 (N_3740,N_2229,N_2924);
and U3741 (N_3741,N_2505,N_2247);
nand U3742 (N_3742,N_2900,N_2598);
and U3743 (N_3743,N_1901,N_2028);
and U3744 (N_3744,N_2558,N_1721);
and U3745 (N_3745,N_1523,N_2269);
and U3746 (N_3746,N_2601,N_2466);
and U3747 (N_3747,N_1841,N_2426);
or U3748 (N_3748,N_2874,N_2478);
xnor U3749 (N_3749,N_2344,N_2908);
or U3750 (N_3750,N_2969,N_2626);
nor U3751 (N_3751,N_2459,N_1882);
nor U3752 (N_3752,N_2578,N_2922);
xor U3753 (N_3753,N_2486,N_2393);
and U3754 (N_3754,N_2405,N_2875);
nand U3755 (N_3755,N_2819,N_2347);
nor U3756 (N_3756,N_2456,N_2973);
and U3757 (N_3757,N_1716,N_2724);
and U3758 (N_3758,N_1564,N_2809);
nor U3759 (N_3759,N_2195,N_1557);
or U3760 (N_3760,N_1595,N_1895);
nor U3761 (N_3761,N_2736,N_2507);
nand U3762 (N_3762,N_1737,N_2428);
and U3763 (N_3763,N_2336,N_2837);
nor U3764 (N_3764,N_2884,N_2081);
nor U3765 (N_3765,N_2141,N_2147);
nor U3766 (N_3766,N_2420,N_1695);
and U3767 (N_3767,N_1823,N_1780);
and U3768 (N_3768,N_1870,N_2511);
nand U3769 (N_3769,N_2791,N_2716);
or U3770 (N_3770,N_2934,N_1673);
nor U3771 (N_3771,N_2858,N_2626);
xnor U3772 (N_3772,N_2776,N_1572);
xnor U3773 (N_3773,N_2395,N_2532);
or U3774 (N_3774,N_2117,N_2703);
or U3775 (N_3775,N_2817,N_2470);
nor U3776 (N_3776,N_2735,N_2218);
or U3777 (N_3777,N_1501,N_2824);
or U3778 (N_3778,N_2125,N_2222);
and U3779 (N_3779,N_1607,N_2510);
or U3780 (N_3780,N_1534,N_1524);
nand U3781 (N_3781,N_1658,N_2248);
nand U3782 (N_3782,N_2161,N_1777);
or U3783 (N_3783,N_2653,N_2550);
nor U3784 (N_3784,N_2091,N_2926);
nand U3785 (N_3785,N_2675,N_1732);
and U3786 (N_3786,N_2790,N_2758);
or U3787 (N_3787,N_1548,N_1872);
nand U3788 (N_3788,N_1768,N_2759);
nor U3789 (N_3789,N_2518,N_2571);
or U3790 (N_3790,N_1610,N_2094);
nand U3791 (N_3791,N_1949,N_1999);
nand U3792 (N_3792,N_2536,N_1923);
nor U3793 (N_3793,N_2727,N_2960);
and U3794 (N_3794,N_2735,N_1704);
and U3795 (N_3795,N_1788,N_2899);
and U3796 (N_3796,N_2837,N_1921);
nand U3797 (N_3797,N_2280,N_2643);
or U3798 (N_3798,N_1978,N_2192);
nor U3799 (N_3799,N_2066,N_2947);
nand U3800 (N_3800,N_1788,N_2372);
xnor U3801 (N_3801,N_1858,N_2720);
nor U3802 (N_3802,N_2564,N_2790);
or U3803 (N_3803,N_2988,N_2462);
or U3804 (N_3804,N_1601,N_1928);
nor U3805 (N_3805,N_2418,N_2956);
xor U3806 (N_3806,N_2227,N_1636);
and U3807 (N_3807,N_2513,N_2029);
nor U3808 (N_3808,N_2119,N_1974);
nand U3809 (N_3809,N_2981,N_2919);
nor U3810 (N_3810,N_2361,N_2941);
xor U3811 (N_3811,N_2941,N_1667);
nand U3812 (N_3812,N_1883,N_1704);
or U3813 (N_3813,N_2170,N_1834);
nand U3814 (N_3814,N_2953,N_1562);
and U3815 (N_3815,N_2452,N_2811);
or U3816 (N_3816,N_2635,N_2379);
nor U3817 (N_3817,N_1690,N_2622);
nor U3818 (N_3818,N_2567,N_2594);
or U3819 (N_3819,N_2468,N_2736);
nor U3820 (N_3820,N_2515,N_2889);
or U3821 (N_3821,N_2983,N_2602);
nor U3822 (N_3822,N_2149,N_2918);
nand U3823 (N_3823,N_1807,N_2890);
and U3824 (N_3824,N_2800,N_2117);
nor U3825 (N_3825,N_1666,N_2725);
and U3826 (N_3826,N_1596,N_2377);
nand U3827 (N_3827,N_2446,N_1870);
nand U3828 (N_3828,N_2124,N_2640);
or U3829 (N_3829,N_2203,N_2712);
xnor U3830 (N_3830,N_2322,N_2537);
or U3831 (N_3831,N_2091,N_2505);
xnor U3832 (N_3832,N_1851,N_2959);
and U3833 (N_3833,N_1949,N_1505);
nand U3834 (N_3834,N_1958,N_1698);
or U3835 (N_3835,N_2546,N_2633);
nor U3836 (N_3836,N_2812,N_2238);
and U3837 (N_3837,N_2055,N_1540);
nand U3838 (N_3838,N_2453,N_2838);
xnor U3839 (N_3839,N_2541,N_2846);
and U3840 (N_3840,N_2308,N_1975);
nand U3841 (N_3841,N_2473,N_2187);
nand U3842 (N_3842,N_2800,N_2861);
and U3843 (N_3843,N_2414,N_1618);
nand U3844 (N_3844,N_2723,N_2806);
nor U3845 (N_3845,N_1712,N_2518);
and U3846 (N_3846,N_2948,N_1662);
nor U3847 (N_3847,N_2730,N_2561);
nor U3848 (N_3848,N_1597,N_1576);
or U3849 (N_3849,N_2033,N_2464);
and U3850 (N_3850,N_2321,N_2387);
nor U3851 (N_3851,N_2979,N_1976);
xnor U3852 (N_3852,N_1758,N_1671);
or U3853 (N_3853,N_1623,N_1878);
or U3854 (N_3854,N_1716,N_1890);
or U3855 (N_3855,N_2623,N_2080);
nand U3856 (N_3856,N_2915,N_2498);
and U3857 (N_3857,N_1623,N_1816);
nor U3858 (N_3858,N_2951,N_1517);
or U3859 (N_3859,N_2592,N_2610);
nand U3860 (N_3860,N_1520,N_1564);
nand U3861 (N_3861,N_1616,N_1630);
and U3862 (N_3862,N_1553,N_2767);
or U3863 (N_3863,N_2490,N_2735);
nand U3864 (N_3864,N_2610,N_2478);
nor U3865 (N_3865,N_2607,N_2608);
or U3866 (N_3866,N_2281,N_2978);
and U3867 (N_3867,N_1516,N_2128);
nand U3868 (N_3868,N_1902,N_1615);
nor U3869 (N_3869,N_2308,N_1633);
or U3870 (N_3870,N_2878,N_2671);
or U3871 (N_3871,N_2558,N_1519);
nor U3872 (N_3872,N_2478,N_1521);
nand U3873 (N_3873,N_2121,N_2168);
or U3874 (N_3874,N_2837,N_1971);
nand U3875 (N_3875,N_2137,N_1565);
nand U3876 (N_3876,N_1942,N_2189);
nand U3877 (N_3877,N_1953,N_2090);
nand U3878 (N_3878,N_2377,N_1912);
or U3879 (N_3879,N_2971,N_1931);
nor U3880 (N_3880,N_2046,N_2978);
nor U3881 (N_3881,N_2695,N_2453);
nor U3882 (N_3882,N_2955,N_2121);
xnor U3883 (N_3883,N_2669,N_2378);
xnor U3884 (N_3884,N_1965,N_2609);
nand U3885 (N_3885,N_1700,N_2532);
and U3886 (N_3886,N_1853,N_2435);
nor U3887 (N_3887,N_2427,N_1786);
nor U3888 (N_3888,N_2213,N_2719);
or U3889 (N_3889,N_1643,N_2388);
nand U3890 (N_3890,N_1639,N_2950);
nand U3891 (N_3891,N_2120,N_1761);
or U3892 (N_3892,N_2789,N_2098);
and U3893 (N_3893,N_1835,N_2884);
or U3894 (N_3894,N_2986,N_2476);
or U3895 (N_3895,N_2207,N_1897);
xor U3896 (N_3896,N_2613,N_2938);
or U3897 (N_3897,N_2424,N_2865);
or U3898 (N_3898,N_2867,N_2433);
or U3899 (N_3899,N_1859,N_2681);
nand U3900 (N_3900,N_2547,N_2697);
nor U3901 (N_3901,N_2054,N_1662);
or U3902 (N_3902,N_2667,N_2644);
nand U3903 (N_3903,N_1863,N_1515);
and U3904 (N_3904,N_1702,N_1555);
xor U3905 (N_3905,N_2814,N_2279);
nor U3906 (N_3906,N_2981,N_2468);
nor U3907 (N_3907,N_2142,N_2679);
xor U3908 (N_3908,N_2522,N_1845);
nand U3909 (N_3909,N_1954,N_1984);
and U3910 (N_3910,N_2126,N_1671);
and U3911 (N_3911,N_1933,N_2909);
nand U3912 (N_3912,N_2758,N_2354);
or U3913 (N_3913,N_2121,N_2002);
and U3914 (N_3914,N_1712,N_2885);
nand U3915 (N_3915,N_2872,N_2681);
or U3916 (N_3916,N_2496,N_1857);
xnor U3917 (N_3917,N_2453,N_2421);
nor U3918 (N_3918,N_2115,N_2548);
and U3919 (N_3919,N_2687,N_1996);
nand U3920 (N_3920,N_2727,N_2858);
or U3921 (N_3921,N_1528,N_2163);
and U3922 (N_3922,N_2302,N_2574);
and U3923 (N_3923,N_1838,N_1630);
xor U3924 (N_3924,N_2282,N_1877);
nand U3925 (N_3925,N_2432,N_2852);
or U3926 (N_3926,N_2620,N_2212);
nor U3927 (N_3927,N_1977,N_2630);
nor U3928 (N_3928,N_2438,N_2373);
or U3929 (N_3929,N_1838,N_2635);
nand U3930 (N_3930,N_2901,N_2391);
and U3931 (N_3931,N_2812,N_1871);
and U3932 (N_3932,N_2813,N_1709);
and U3933 (N_3933,N_2490,N_2474);
nand U3934 (N_3934,N_2687,N_2786);
nor U3935 (N_3935,N_2224,N_2182);
nor U3936 (N_3936,N_2811,N_2429);
nor U3937 (N_3937,N_2167,N_2293);
nand U3938 (N_3938,N_2230,N_1604);
nand U3939 (N_3939,N_2443,N_2325);
nand U3940 (N_3940,N_1726,N_2771);
nor U3941 (N_3941,N_2043,N_2765);
and U3942 (N_3942,N_2361,N_2194);
or U3943 (N_3943,N_2530,N_2051);
nand U3944 (N_3944,N_2713,N_1832);
and U3945 (N_3945,N_2331,N_2472);
and U3946 (N_3946,N_2827,N_1776);
nand U3947 (N_3947,N_1704,N_1808);
nand U3948 (N_3948,N_2138,N_2560);
or U3949 (N_3949,N_1961,N_2354);
nand U3950 (N_3950,N_1632,N_1765);
nor U3951 (N_3951,N_2062,N_2171);
and U3952 (N_3952,N_2218,N_2043);
and U3953 (N_3953,N_2912,N_2782);
nor U3954 (N_3954,N_1607,N_2336);
nand U3955 (N_3955,N_2997,N_1898);
and U3956 (N_3956,N_1566,N_1840);
and U3957 (N_3957,N_1734,N_2860);
nor U3958 (N_3958,N_2452,N_2737);
or U3959 (N_3959,N_2594,N_1509);
xor U3960 (N_3960,N_1578,N_2315);
or U3961 (N_3961,N_1718,N_2542);
nor U3962 (N_3962,N_2594,N_1628);
nor U3963 (N_3963,N_1605,N_2421);
or U3964 (N_3964,N_1979,N_1807);
nor U3965 (N_3965,N_2793,N_2009);
or U3966 (N_3966,N_2203,N_2284);
nor U3967 (N_3967,N_2252,N_2891);
or U3968 (N_3968,N_1957,N_1564);
or U3969 (N_3969,N_1734,N_2917);
xor U3970 (N_3970,N_2059,N_2676);
or U3971 (N_3971,N_2866,N_2521);
nor U3972 (N_3972,N_1956,N_2852);
and U3973 (N_3973,N_2759,N_1567);
nor U3974 (N_3974,N_2768,N_2920);
nand U3975 (N_3975,N_2729,N_1714);
xnor U3976 (N_3976,N_1787,N_1713);
and U3977 (N_3977,N_1596,N_1848);
nand U3978 (N_3978,N_2660,N_2867);
and U3979 (N_3979,N_2745,N_2331);
xnor U3980 (N_3980,N_2097,N_2210);
or U3981 (N_3981,N_1742,N_1517);
or U3982 (N_3982,N_2970,N_1648);
nand U3983 (N_3983,N_2334,N_2205);
nor U3984 (N_3984,N_2236,N_1560);
or U3985 (N_3985,N_2127,N_1972);
and U3986 (N_3986,N_2715,N_2648);
xnor U3987 (N_3987,N_2389,N_2908);
nor U3988 (N_3988,N_1516,N_1674);
xor U3989 (N_3989,N_2657,N_1529);
or U3990 (N_3990,N_2698,N_1890);
nor U3991 (N_3991,N_2171,N_2722);
nor U3992 (N_3992,N_1948,N_1690);
and U3993 (N_3993,N_1693,N_2019);
or U3994 (N_3994,N_1841,N_2352);
nand U3995 (N_3995,N_2580,N_1993);
nand U3996 (N_3996,N_2074,N_2860);
or U3997 (N_3997,N_2388,N_2044);
nand U3998 (N_3998,N_2390,N_1967);
and U3999 (N_3999,N_2994,N_1635);
and U4000 (N_4000,N_2710,N_1811);
or U4001 (N_4001,N_2779,N_2799);
nand U4002 (N_4002,N_2962,N_2193);
nor U4003 (N_4003,N_2483,N_2312);
nand U4004 (N_4004,N_2570,N_2493);
or U4005 (N_4005,N_1536,N_2387);
nor U4006 (N_4006,N_2491,N_2741);
or U4007 (N_4007,N_1895,N_2295);
or U4008 (N_4008,N_2340,N_2309);
and U4009 (N_4009,N_1853,N_2551);
nor U4010 (N_4010,N_2613,N_2533);
or U4011 (N_4011,N_2010,N_2069);
nand U4012 (N_4012,N_2830,N_1849);
xor U4013 (N_4013,N_2022,N_2409);
nor U4014 (N_4014,N_2257,N_1541);
or U4015 (N_4015,N_1795,N_1743);
and U4016 (N_4016,N_2113,N_2870);
nand U4017 (N_4017,N_1502,N_1846);
or U4018 (N_4018,N_2781,N_2244);
nor U4019 (N_4019,N_1967,N_1833);
and U4020 (N_4020,N_2487,N_2843);
or U4021 (N_4021,N_2386,N_2743);
nor U4022 (N_4022,N_2852,N_2697);
or U4023 (N_4023,N_2002,N_2000);
nand U4024 (N_4024,N_2848,N_2858);
and U4025 (N_4025,N_1698,N_2034);
nand U4026 (N_4026,N_2542,N_2001);
and U4027 (N_4027,N_2303,N_2627);
or U4028 (N_4028,N_1593,N_2345);
nand U4029 (N_4029,N_1632,N_1815);
or U4030 (N_4030,N_1851,N_1691);
xnor U4031 (N_4031,N_2551,N_2082);
nor U4032 (N_4032,N_2401,N_1996);
nor U4033 (N_4033,N_2281,N_2547);
or U4034 (N_4034,N_2968,N_2747);
or U4035 (N_4035,N_1645,N_1576);
nand U4036 (N_4036,N_1674,N_2209);
or U4037 (N_4037,N_2188,N_2521);
nand U4038 (N_4038,N_2995,N_1955);
and U4039 (N_4039,N_1958,N_1942);
and U4040 (N_4040,N_1754,N_2412);
nand U4041 (N_4041,N_2370,N_2250);
or U4042 (N_4042,N_2812,N_1854);
nand U4043 (N_4043,N_2317,N_1503);
or U4044 (N_4044,N_1887,N_2737);
and U4045 (N_4045,N_1731,N_2104);
or U4046 (N_4046,N_2942,N_2915);
nor U4047 (N_4047,N_2633,N_2473);
or U4048 (N_4048,N_1707,N_2467);
xnor U4049 (N_4049,N_2975,N_1975);
nor U4050 (N_4050,N_2852,N_1519);
or U4051 (N_4051,N_2410,N_2881);
or U4052 (N_4052,N_2495,N_2991);
and U4053 (N_4053,N_1710,N_2439);
nor U4054 (N_4054,N_1598,N_2206);
nor U4055 (N_4055,N_2971,N_1723);
nand U4056 (N_4056,N_2639,N_2729);
and U4057 (N_4057,N_2524,N_1668);
and U4058 (N_4058,N_2711,N_2387);
and U4059 (N_4059,N_2771,N_1868);
xnor U4060 (N_4060,N_2608,N_1967);
or U4061 (N_4061,N_1690,N_1524);
or U4062 (N_4062,N_1701,N_1807);
or U4063 (N_4063,N_2637,N_1888);
nand U4064 (N_4064,N_2304,N_1865);
nand U4065 (N_4065,N_2438,N_1710);
and U4066 (N_4066,N_2374,N_1992);
nor U4067 (N_4067,N_2973,N_2833);
nor U4068 (N_4068,N_1698,N_2168);
and U4069 (N_4069,N_2678,N_2878);
or U4070 (N_4070,N_1628,N_1728);
and U4071 (N_4071,N_1694,N_2239);
nand U4072 (N_4072,N_2495,N_2138);
nand U4073 (N_4073,N_2866,N_2125);
xnor U4074 (N_4074,N_1531,N_2298);
and U4075 (N_4075,N_1868,N_2772);
or U4076 (N_4076,N_1982,N_2304);
nand U4077 (N_4077,N_2809,N_1773);
nor U4078 (N_4078,N_1992,N_2019);
nand U4079 (N_4079,N_2364,N_2411);
nor U4080 (N_4080,N_2671,N_2752);
and U4081 (N_4081,N_2171,N_2441);
and U4082 (N_4082,N_2968,N_1514);
nand U4083 (N_4083,N_1627,N_1802);
or U4084 (N_4084,N_1507,N_2608);
xor U4085 (N_4085,N_2281,N_2886);
nor U4086 (N_4086,N_1791,N_1542);
nor U4087 (N_4087,N_2195,N_2249);
and U4088 (N_4088,N_1884,N_1629);
xnor U4089 (N_4089,N_1641,N_1895);
nand U4090 (N_4090,N_1979,N_2832);
nor U4091 (N_4091,N_2634,N_2516);
and U4092 (N_4092,N_2151,N_2548);
xor U4093 (N_4093,N_1946,N_1581);
nand U4094 (N_4094,N_2254,N_2241);
nor U4095 (N_4095,N_2638,N_2678);
or U4096 (N_4096,N_1996,N_2818);
or U4097 (N_4097,N_2521,N_2034);
nor U4098 (N_4098,N_2326,N_2922);
nand U4099 (N_4099,N_2998,N_1766);
nand U4100 (N_4100,N_2031,N_2735);
nor U4101 (N_4101,N_2036,N_2055);
and U4102 (N_4102,N_1960,N_2804);
nor U4103 (N_4103,N_1779,N_1899);
nor U4104 (N_4104,N_1762,N_2285);
and U4105 (N_4105,N_2376,N_1614);
nand U4106 (N_4106,N_2287,N_1741);
and U4107 (N_4107,N_1590,N_2114);
or U4108 (N_4108,N_1684,N_2683);
xor U4109 (N_4109,N_2716,N_2429);
xnor U4110 (N_4110,N_1802,N_1861);
or U4111 (N_4111,N_2083,N_1537);
and U4112 (N_4112,N_1534,N_2610);
or U4113 (N_4113,N_1530,N_2458);
nand U4114 (N_4114,N_1690,N_2048);
or U4115 (N_4115,N_2746,N_2467);
nor U4116 (N_4116,N_1508,N_2039);
nand U4117 (N_4117,N_2831,N_2470);
nor U4118 (N_4118,N_2586,N_2743);
or U4119 (N_4119,N_2799,N_1598);
nor U4120 (N_4120,N_2413,N_2758);
nor U4121 (N_4121,N_1789,N_2100);
nor U4122 (N_4122,N_2534,N_2552);
nand U4123 (N_4123,N_1695,N_1654);
nor U4124 (N_4124,N_1716,N_1735);
nand U4125 (N_4125,N_2862,N_1744);
nor U4126 (N_4126,N_2993,N_2206);
or U4127 (N_4127,N_1742,N_1593);
nand U4128 (N_4128,N_2013,N_2553);
and U4129 (N_4129,N_2364,N_1907);
and U4130 (N_4130,N_2360,N_1793);
nand U4131 (N_4131,N_2957,N_2736);
and U4132 (N_4132,N_2860,N_2557);
or U4133 (N_4133,N_2868,N_1961);
nand U4134 (N_4134,N_1753,N_2656);
xor U4135 (N_4135,N_2750,N_2542);
nand U4136 (N_4136,N_2308,N_1507);
xor U4137 (N_4137,N_2049,N_2962);
nand U4138 (N_4138,N_1757,N_1758);
or U4139 (N_4139,N_2882,N_2838);
or U4140 (N_4140,N_1800,N_2693);
nand U4141 (N_4141,N_2361,N_2460);
nand U4142 (N_4142,N_1921,N_2088);
nor U4143 (N_4143,N_2014,N_2806);
nor U4144 (N_4144,N_2016,N_2216);
or U4145 (N_4145,N_1927,N_1987);
nor U4146 (N_4146,N_2677,N_2030);
or U4147 (N_4147,N_1703,N_1539);
nor U4148 (N_4148,N_1672,N_2789);
and U4149 (N_4149,N_2324,N_2794);
and U4150 (N_4150,N_2603,N_2294);
nand U4151 (N_4151,N_1516,N_2083);
or U4152 (N_4152,N_2434,N_2416);
and U4153 (N_4153,N_2006,N_2404);
xor U4154 (N_4154,N_1711,N_1709);
or U4155 (N_4155,N_2129,N_2063);
nand U4156 (N_4156,N_2714,N_2540);
or U4157 (N_4157,N_2544,N_1983);
xor U4158 (N_4158,N_2193,N_2517);
or U4159 (N_4159,N_2800,N_2218);
or U4160 (N_4160,N_2944,N_2036);
and U4161 (N_4161,N_2950,N_2500);
or U4162 (N_4162,N_2624,N_2246);
xnor U4163 (N_4163,N_1548,N_2321);
xor U4164 (N_4164,N_2553,N_2675);
nor U4165 (N_4165,N_2916,N_2285);
nand U4166 (N_4166,N_2032,N_2017);
or U4167 (N_4167,N_1803,N_2510);
nand U4168 (N_4168,N_2140,N_1985);
nor U4169 (N_4169,N_2480,N_2086);
nor U4170 (N_4170,N_2884,N_2816);
or U4171 (N_4171,N_1954,N_2911);
and U4172 (N_4172,N_1727,N_1775);
xnor U4173 (N_4173,N_1507,N_2711);
or U4174 (N_4174,N_2005,N_2315);
or U4175 (N_4175,N_2073,N_2708);
or U4176 (N_4176,N_1942,N_2845);
or U4177 (N_4177,N_2720,N_2044);
nand U4178 (N_4178,N_2325,N_1914);
nand U4179 (N_4179,N_2318,N_2479);
nand U4180 (N_4180,N_1799,N_2700);
xnor U4181 (N_4181,N_2611,N_2392);
or U4182 (N_4182,N_2080,N_2130);
nand U4183 (N_4183,N_2916,N_2137);
nor U4184 (N_4184,N_2838,N_2247);
nand U4185 (N_4185,N_1693,N_2427);
nand U4186 (N_4186,N_2613,N_2546);
and U4187 (N_4187,N_1853,N_2864);
or U4188 (N_4188,N_2155,N_2715);
nand U4189 (N_4189,N_2497,N_1702);
nand U4190 (N_4190,N_2478,N_2396);
or U4191 (N_4191,N_1969,N_1825);
nand U4192 (N_4192,N_2263,N_2644);
or U4193 (N_4193,N_1638,N_1888);
nor U4194 (N_4194,N_2514,N_2736);
nor U4195 (N_4195,N_1566,N_1859);
and U4196 (N_4196,N_1935,N_2205);
or U4197 (N_4197,N_2560,N_1582);
or U4198 (N_4198,N_1642,N_2980);
nand U4199 (N_4199,N_2190,N_1649);
nor U4200 (N_4200,N_2507,N_2328);
nor U4201 (N_4201,N_2592,N_2954);
nand U4202 (N_4202,N_1574,N_2633);
xor U4203 (N_4203,N_2494,N_1515);
or U4204 (N_4204,N_1812,N_2988);
and U4205 (N_4205,N_1984,N_2851);
nor U4206 (N_4206,N_1566,N_2433);
nor U4207 (N_4207,N_1755,N_2038);
xor U4208 (N_4208,N_1559,N_1992);
nand U4209 (N_4209,N_1821,N_2466);
and U4210 (N_4210,N_2186,N_2060);
nand U4211 (N_4211,N_1550,N_2967);
nor U4212 (N_4212,N_2465,N_1578);
xor U4213 (N_4213,N_2458,N_2465);
or U4214 (N_4214,N_1629,N_2911);
and U4215 (N_4215,N_2088,N_1739);
and U4216 (N_4216,N_2006,N_2078);
and U4217 (N_4217,N_2713,N_2898);
nor U4218 (N_4218,N_1878,N_2815);
or U4219 (N_4219,N_2349,N_2905);
nand U4220 (N_4220,N_1765,N_2703);
nand U4221 (N_4221,N_2017,N_2029);
xnor U4222 (N_4222,N_1539,N_2540);
nand U4223 (N_4223,N_1556,N_2190);
and U4224 (N_4224,N_2008,N_2381);
nand U4225 (N_4225,N_1578,N_1726);
or U4226 (N_4226,N_2243,N_2626);
nor U4227 (N_4227,N_2984,N_2415);
or U4228 (N_4228,N_2839,N_2514);
nand U4229 (N_4229,N_1518,N_2754);
nand U4230 (N_4230,N_2214,N_1518);
nor U4231 (N_4231,N_1648,N_2390);
or U4232 (N_4232,N_2417,N_1729);
and U4233 (N_4233,N_1538,N_2966);
xnor U4234 (N_4234,N_2138,N_2974);
nor U4235 (N_4235,N_2007,N_1502);
xor U4236 (N_4236,N_2798,N_2351);
or U4237 (N_4237,N_2866,N_1739);
or U4238 (N_4238,N_1577,N_2560);
or U4239 (N_4239,N_2560,N_2012);
nor U4240 (N_4240,N_1552,N_2291);
xnor U4241 (N_4241,N_2612,N_2776);
or U4242 (N_4242,N_1998,N_2419);
or U4243 (N_4243,N_2595,N_2794);
nor U4244 (N_4244,N_2372,N_1747);
nor U4245 (N_4245,N_2487,N_2472);
or U4246 (N_4246,N_1875,N_2125);
xor U4247 (N_4247,N_2337,N_1946);
nand U4248 (N_4248,N_2255,N_2592);
nand U4249 (N_4249,N_2525,N_1804);
nor U4250 (N_4250,N_2833,N_2862);
xnor U4251 (N_4251,N_2638,N_1737);
nor U4252 (N_4252,N_2103,N_1939);
nor U4253 (N_4253,N_1660,N_2148);
nor U4254 (N_4254,N_1542,N_2341);
nand U4255 (N_4255,N_1778,N_2220);
and U4256 (N_4256,N_1697,N_1723);
nand U4257 (N_4257,N_1672,N_1932);
nor U4258 (N_4258,N_2211,N_2592);
nand U4259 (N_4259,N_2340,N_1914);
or U4260 (N_4260,N_2934,N_2603);
nand U4261 (N_4261,N_2408,N_2087);
nand U4262 (N_4262,N_1578,N_2825);
xor U4263 (N_4263,N_2507,N_2546);
nor U4264 (N_4264,N_2235,N_2065);
nand U4265 (N_4265,N_2604,N_2739);
nand U4266 (N_4266,N_1882,N_1821);
or U4267 (N_4267,N_1932,N_1933);
xor U4268 (N_4268,N_2107,N_2407);
and U4269 (N_4269,N_2228,N_1786);
and U4270 (N_4270,N_2562,N_2398);
nor U4271 (N_4271,N_2684,N_2162);
or U4272 (N_4272,N_1785,N_1692);
xor U4273 (N_4273,N_2375,N_2035);
and U4274 (N_4274,N_2163,N_2425);
xor U4275 (N_4275,N_1809,N_2154);
or U4276 (N_4276,N_2710,N_2669);
xnor U4277 (N_4277,N_1671,N_2880);
and U4278 (N_4278,N_2977,N_2784);
or U4279 (N_4279,N_2727,N_2123);
nor U4280 (N_4280,N_2040,N_2248);
or U4281 (N_4281,N_1788,N_2292);
nand U4282 (N_4282,N_2650,N_2125);
or U4283 (N_4283,N_2672,N_2306);
xor U4284 (N_4284,N_2690,N_1789);
nand U4285 (N_4285,N_2859,N_2229);
and U4286 (N_4286,N_2646,N_2455);
nand U4287 (N_4287,N_2151,N_2675);
nor U4288 (N_4288,N_1920,N_2395);
xnor U4289 (N_4289,N_2393,N_1837);
nand U4290 (N_4290,N_1501,N_2998);
nor U4291 (N_4291,N_2242,N_1907);
and U4292 (N_4292,N_1816,N_1820);
nand U4293 (N_4293,N_1855,N_1998);
nand U4294 (N_4294,N_1937,N_1876);
nor U4295 (N_4295,N_2775,N_2432);
and U4296 (N_4296,N_1827,N_1602);
or U4297 (N_4297,N_1788,N_2492);
nor U4298 (N_4298,N_2532,N_2296);
nor U4299 (N_4299,N_2572,N_1740);
and U4300 (N_4300,N_2317,N_1621);
nor U4301 (N_4301,N_1699,N_2321);
and U4302 (N_4302,N_2803,N_2897);
nor U4303 (N_4303,N_2422,N_2118);
and U4304 (N_4304,N_2814,N_2444);
nand U4305 (N_4305,N_2016,N_1661);
nand U4306 (N_4306,N_1981,N_1896);
nand U4307 (N_4307,N_2141,N_2456);
and U4308 (N_4308,N_1686,N_2550);
or U4309 (N_4309,N_1733,N_1691);
nor U4310 (N_4310,N_2634,N_2211);
or U4311 (N_4311,N_1974,N_2736);
and U4312 (N_4312,N_2540,N_1778);
nor U4313 (N_4313,N_2418,N_2592);
nor U4314 (N_4314,N_2269,N_2946);
and U4315 (N_4315,N_2712,N_2266);
or U4316 (N_4316,N_2839,N_2545);
and U4317 (N_4317,N_1896,N_2340);
or U4318 (N_4318,N_1737,N_2561);
and U4319 (N_4319,N_2868,N_1671);
and U4320 (N_4320,N_2969,N_2827);
nor U4321 (N_4321,N_1982,N_2004);
or U4322 (N_4322,N_2785,N_2907);
xor U4323 (N_4323,N_2078,N_1574);
nor U4324 (N_4324,N_2131,N_2330);
nor U4325 (N_4325,N_2746,N_2663);
nand U4326 (N_4326,N_2825,N_2429);
nand U4327 (N_4327,N_2063,N_2387);
and U4328 (N_4328,N_2754,N_2685);
nand U4329 (N_4329,N_1840,N_2171);
nand U4330 (N_4330,N_2935,N_1695);
and U4331 (N_4331,N_1843,N_2974);
or U4332 (N_4332,N_2969,N_2105);
nor U4333 (N_4333,N_2456,N_2098);
xnor U4334 (N_4334,N_1712,N_2984);
or U4335 (N_4335,N_2651,N_2344);
nor U4336 (N_4336,N_2548,N_2701);
nor U4337 (N_4337,N_2709,N_2231);
or U4338 (N_4338,N_2554,N_2083);
nand U4339 (N_4339,N_1611,N_1963);
or U4340 (N_4340,N_1968,N_2064);
nand U4341 (N_4341,N_2057,N_2730);
and U4342 (N_4342,N_2724,N_2224);
and U4343 (N_4343,N_1841,N_2043);
and U4344 (N_4344,N_1694,N_2227);
and U4345 (N_4345,N_2047,N_2484);
nand U4346 (N_4346,N_2393,N_2597);
nand U4347 (N_4347,N_2287,N_2131);
or U4348 (N_4348,N_2278,N_2671);
and U4349 (N_4349,N_1763,N_2961);
xor U4350 (N_4350,N_2972,N_1821);
nor U4351 (N_4351,N_2721,N_2398);
xor U4352 (N_4352,N_2512,N_1993);
nor U4353 (N_4353,N_1542,N_2274);
or U4354 (N_4354,N_2537,N_2296);
nor U4355 (N_4355,N_2549,N_2407);
and U4356 (N_4356,N_1974,N_1859);
xor U4357 (N_4357,N_2283,N_2349);
or U4358 (N_4358,N_2106,N_2254);
nor U4359 (N_4359,N_2402,N_2848);
or U4360 (N_4360,N_2028,N_2177);
or U4361 (N_4361,N_2012,N_2147);
nand U4362 (N_4362,N_2975,N_2823);
nand U4363 (N_4363,N_1954,N_2191);
or U4364 (N_4364,N_2870,N_1996);
and U4365 (N_4365,N_2979,N_1602);
xor U4366 (N_4366,N_1763,N_2859);
nand U4367 (N_4367,N_1936,N_2360);
nand U4368 (N_4368,N_1709,N_2416);
nand U4369 (N_4369,N_1975,N_2394);
nand U4370 (N_4370,N_2427,N_1725);
and U4371 (N_4371,N_2414,N_2382);
or U4372 (N_4372,N_1790,N_2446);
nand U4373 (N_4373,N_2955,N_1689);
and U4374 (N_4374,N_2002,N_2041);
and U4375 (N_4375,N_1624,N_2766);
nand U4376 (N_4376,N_2253,N_2099);
and U4377 (N_4377,N_2085,N_2414);
nor U4378 (N_4378,N_1626,N_1526);
nand U4379 (N_4379,N_2492,N_1581);
or U4380 (N_4380,N_2548,N_2489);
and U4381 (N_4381,N_2477,N_2386);
nand U4382 (N_4382,N_2633,N_2889);
nor U4383 (N_4383,N_2119,N_2773);
and U4384 (N_4384,N_2735,N_2519);
nor U4385 (N_4385,N_2964,N_1755);
nor U4386 (N_4386,N_1907,N_2603);
nor U4387 (N_4387,N_1838,N_2041);
or U4388 (N_4388,N_2905,N_2856);
and U4389 (N_4389,N_2115,N_1743);
and U4390 (N_4390,N_2748,N_1681);
nor U4391 (N_4391,N_2388,N_1807);
and U4392 (N_4392,N_2640,N_2931);
and U4393 (N_4393,N_1870,N_2738);
xor U4394 (N_4394,N_2755,N_2725);
nand U4395 (N_4395,N_2587,N_1537);
or U4396 (N_4396,N_2747,N_2216);
or U4397 (N_4397,N_2641,N_2559);
nand U4398 (N_4398,N_1947,N_1529);
nor U4399 (N_4399,N_1943,N_2518);
and U4400 (N_4400,N_1754,N_2832);
nand U4401 (N_4401,N_2577,N_1917);
xor U4402 (N_4402,N_1661,N_2103);
nand U4403 (N_4403,N_2647,N_2956);
xor U4404 (N_4404,N_1632,N_2910);
nor U4405 (N_4405,N_2832,N_2145);
nor U4406 (N_4406,N_1947,N_1658);
nand U4407 (N_4407,N_2619,N_1859);
nor U4408 (N_4408,N_2222,N_1763);
or U4409 (N_4409,N_2875,N_2364);
nand U4410 (N_4410,N_1665,N_1817);
and U4411 (N_4411,N_2946,N_2849);
or U4412 (N_4412,N_2713,N_1703);
and U4413 (N_4413,N_2173,N_2862);
xor U4414 (N_4414,N_2555,N_1739);
nand U4415 (N_4415,N_2153,N_2236);
and U4416 (N_4416,N_2773,N_1508);
nor U4417 (N_4417,N_2884,N_2785);
nor U4418 (N_4418,N_2095,N_2992);
and U4419 (N_4419,N_1923,N_1736);
and U4420 (N_4420,N_1741,N_2739);
or U4421 (N_4421,N_2240,N_2410);
nor U4422 (N_4422,N_2914,N_1710);
xnor U4423 (N_4423,N_2314,N_2727);
nand U4424 (N_4424,N_2259,N_2950);
or U4425 (N_4425,N_1982,N_1737);
nand U4426 (N_4426,N_2978,N_2031);
xor U4427 (N_4427,N_1589,N_2082);
nor U4428 (N_4428,N_2986,N_1526);
or U4429 (N_4429,N_2212,N_2226);
and U4430 (N_4430,N_1599,N_1780);
and U4431 (N_4431,N_2929,N_2902);
nor U4432 (N_4432,N_2294,N_2472);
or U4433 (N_4433,N_1904,N_2693);
nor U4434 (N_4434,N_2420,N_2289);
or U4435 (N_4435,N_1677,N_2103);
nand U4436 (N_4436,N_1776,N_2928);
nor U4437 (N_4437,N_2764,N_2265);
or U4438 (N_4438,N_2058,N_1591);
nor U4439 (N_4439,N_1923,N_2641);
or U4440 (N_4440,N_1970,N_1944);
and U4441 (N_4441,N_1673,N_2370);
or U4442 (N_4442,N_1866,N_2221);
and U4443 (N_4443,N_1724,N_1877);
and U4444 (N_4444,N_2920,N_2254);
or U4445 (N_4445,N_2735,N_2607);
nor U4446 (N_4446,N_2277,N_2840);
nor U4447 (N_4447,N_2498,N_2443);
nand U4448 (N_4448,N_2424,N_2932);
nand U4449 (N_4449,N_1819,N_1540);
or U4450 (N_4450,N_1558,N_2045);
nand U4451 (N_4451,N_2094,N_1515);
nor U4452 (N_4452,N_1782,N_1923);
xnor U4453 (N_4453,N_1592,N_2164);
nor U4454 (N_4454,N_2941,N_1821);
nand U4455 (N_4455,N_2352,N_2552);
nand U4456 (N_4456,N_2810,N_1821);
nand U4457 (N_4457,N_2104,N_2272);
nand U4458 (N_4458,N_2937,N_2285);
nand U4459 (N_4459,N_2770,N_2010);
nand U4460 (N_4460,N_2220,N_2313);
nor U4461 (N_4461,N_2342,N_2659);
and U4462 (N_4462,N_1668,N_1958);
and U4463 (N_4463,N_1614,N_2119);
xnor U4464 (N_4464,N_2752,N_1873);
nor U4465 (N_4465,N_1761,N_2642);
or U4466 (N_4466,N_2853,N_2307);
nand U4467 (N_4467,N_1894,N_2284);
nor U4468 (N_4468,N_1632,N_2751);
and U4469 (N_4469,N_2281,N_2987);
nand U4470 (N_4470,N_1813,N_2338);
nor U4471 (N_4471,N_1913,N_2077);
nor U4472 (N_4472,N_2063,N_2266);
nor U4473 (N_4473,N_2676,N_2166);
nand U4474 (N_4474,N_1586,N_2537);
nor U4475 (N_4475,N_1863,N_2097);
nor U4476 (N_4476,N_2112,N_1903);
and U4477 (N_4477,N_1957,N_2319);
and U4478 (N_4478,N_2744,N_1712);
xnor U4479 (N_4479,N_2479,N_1626);
nand U4480 (N_4480,N_1787,N_2950);
and U4481 (N_4481,N_1507,N_1658);
nor U4482 (N_4482,N_2428,N_1791);
or U4483 (N_4483,N_1715,N_1815);
nand U4484 (N_4484,N_1544,N_1515);
or U4485 (N_4485,N_2493,N_1564);
or U4486 (N_4486,N_2158,N_1718);
and U4487 (N_4487,N_1919,N_2669);
nand U4488 (N_4488,N_2471,N_2808);
nand U4489 (N_4489,N_2674,N_1672);
or U4490 (N_4490,N_2658,N_1923);
nand U4491 (N_4491,N_2422,N_2897);
xnor U4492 (N_4492,N_2011,N_1953);
nand U4493 (N_4493,N_2951,N_2994);
and U4494 (N_4494,N_1988,N_2439);
and U4495 (N_4495,N_1579,N_1843);
and U4496 (N_4496,N_2834,N_1873);
and U4497 (N_4497,N_1722,N_2562);
xor U4498 (N_4498,N_2065,N_2138);
nand U4499 (N_4499,N_2801,N_2638);
nor U4500 (N_4500,N_3176,N_4015);
or U4501 (N_4501,N_3350,N_3718);
or U4502 (N_4502,N_3550,N_3390);
nor U4503 (N_4503,N_3192,N_3293);
or U4504 (N_4504,N_3609,N_3997);
nand U4505 (N_4505,N_3150,N_3715);
nand U4506 (N_4506,N_3043,N_3860);
nand U4507 (N_4507,N_3213,N_4049);
nand U4508 (N_4508,N_4076,N_4370);
and U4509 (N_4509,N_3976,N_3931);
and U4510 (N_4510,N_4089,N_3786);
nor U4511 (N_4511,N_4483,N_3728);
or U4512 (N_4512,N_3606,N_4428);
or U4513 (N_4513,N_3086,N_3926);
nor U4514 (N_4514,N_4338,N_4197);
or U4515 (N_4515,N_3536,N_3713);
nand U4516 (N_4516,N_4423,N_4010);
nand U4517 (N_4517,N_3085,N_3358);
or U4518 (N_4518,N_3189,N_3287);
and U4519 (N_4519,N_4401,N_4119);
xor U4520 (N_4520,N_3450,N_3357);
nor U4521 (N_4521,N_4218,N_3765);
and U4522 (N_4522,N_3615,N_3511);
nor U4523 (N_4523,N_3842,N_3826);
nor U4524 (N_4524,N_3468,N_4219);
or U4525 (N_4525,N_4053,N_4103);
and U4526 (N_4526,N_3971,N_4486);
or U4527 (N_4527,N_3201,N_3968);
nor U4528 (N_4528,N_4395,N_3092);
nor U4529 (N_4529,N_4029,N_4140);
nor U4530 (N_4530,N_3636,N_4208);
or U4531 (N_4531,N_3344,N_4324);
or U4532 (N_4532,N_3366,N_3809);
xor U4533 (N_4533,N_3608,N_3584);
nand U4534 (N_4534,N_4356,N_3900);
nor U4535 (N_4535,N_3214,N_3649);
or U4536 (N_4536,N_3046,N_3736);
nor U4537 (N_4537,N_3423,N_3061);
nand U4538 (N_4538,N_3072,N_3701);
or U4539 (N_4539,N_4038,N_3682);
nor U4540 (N_4540,N_4367,N_3578);
nor U4541 (N_4541,N_4259,N_3633);
nand U4542 (N_4542,N_3370,N_4052);
and U4543 (N_4543,N_3671,N_3603);
nor U4544 (N_4544,N_3879,N_3784);
or U4545 (N_4545,N_4333,N_4144);
nand U4546 (N_4546,N_3074,N_4037);
or U4547 (N_4547,N_3021,N_3805);
nand U4548 (N_4548,N_4301,N_3726);
and U4549 (N_4549,N_3032,N_3979);
nor U4550 (N_4550,N_4105,N_3022);
nor U4551 (N_4551,N_4067,N_3241);
or U4552 (N_4552,N_3017,N_3735);
and U4553 (N_4553,N_4439,N_3652);
or U4554 (N_4554,N_3434,N_4148);
nand U4555 (N_4555,N_3980,N_3400);
and U4556 (N_4556,N_3588,N_4080);
and U4557 (N_4557,N_3693,N_3523);
nor U4558 (N_4558,N_4388,N_3013);
nand U4559 (N_4559,N_3310,N_3121);
and U4560 (N_4560,N_4143,N_4255);
and U4561 (N_4561,N_3932,N_3525);
nand U4562 (N_4562,N_4109,N_4203);
xnor U4563 (N_4563,N_3341,N_3385);
nor U4564 (N_4564,N_3600,N_3903);
xor U4565 (N_4565,N_3650,N_3493);
and U4566 (N_4566,N_4350,N_3079);
nor U4567 (N_4567,N_3747,N_3259);
and U4568 (N_4568,N_4344,N_3955);
or U4569 (N_4569,N_3462,N_3300);
and U4570 (N_4570,N_3484,N_3863);
and U4571 (N_4571,N_3597,N_4481);
xor U4572 (N_4572,N_3379,N_3730);
and U4573 (N_4573,N_3539,N_3200);
nand U4574 (N_4574,N_3772,N_4434);
nand U4575 (N_4575,N_3054,N_3948);
and U4576 (N_4576,N_4376,N_3263);
nor U4577 (N_4577,N_4045,N_3995);
nor U4578 (N_4578,N_4251,N_3570);
and U4579 (N_4579,N_3288,N_3031);
nor U4580 (N_4580,N_3965,N_3224);
or U4581 (N_4581,N_4149,N_3655);
xnor U4582 (N_4582,N_3449,N_4393);
and U4583 (N_4583,N_4059,N_3299);
nor U4584 (N_4584,N_4195,N_3937);
and U4585 (N_4585,N_4378,N_3365);
nor U4586 (N_4586,N_4377,N_3210);
or U4587 (N_4587,N_4025,N_4297);
nor U4588 (N_4588,N_4436,N_3676);
and U4589 (N_4589,N_3376,N_3482);
and U4590 (N_4590,N_3729,N_4207);
and U4591 (N_4591,N_4491,N_3590);
or U4592 (N_4592,N_4249,N_3537);
nand U4593 (N_4593,N_3262,N_4005);
or U4594 (N_4594,N_3993,N_3977);
xor U4595 (N_4595,N_3549,N_3292);
nor U4596 (N_4596,N_4294,N_4346);
xnor U4597 (N_4597,N_3798,N_3432);
nor U4598 (N_4598,N_4232,N_3489);
nor U4599 (N_4599,N_3301,N_4335);
or U4600 (N_4600,N_3131,N_3561);
nor U4601 (N_4601,N_4159,N_4134);
and U4602 (N_4602,N_3169,N_3834);
nand U4603 (N_4603,N_3488,N_3473);
nand U4604 (N_4604,N_3795,N_4183);
nand U4605 (N_4605,N_3720,N_3741);
xor U4606 (N_4606,N_3198,N_4492);
xnor U4607 (N_4607,N_3972,N_3982);
nand U4608 (N_4608,N_3497,N_3235);
and U4609 (N_4609,N_3424,N_3229);
and U4610 (N_4610,N_4222,N_3501);
nand U4611 (N_4611,N_4457,N_3068);
nand U4612 (N_4612,N_3643,N_3986);
or U4613 (N_4613,N_3148,N_4090);
nor U4614 (N_4614,N_4055,N_3315);
or U4615 (N_4615,N_4343,N_4156);
and U4616 (N_4616,N_3311,N_3757);
or U4617 (N_4617,N_3388,N_3081);
and U4618 (N_4618,N_4086,N_3771);
nand U4619 (N_4619,N_3743,N_3058);
nand U4620 (N_4620,N_4136,N_3605);
or U4621 (N_4621,N_4215,N_3094);
nor U4622 (N_4622,N_4058,N_3167);
nor U4623 (N_4623,N_4050,N_3958);
nand U4624 (N_4624,N_3408,N_3171);
nand U4625 (N_4625,N_3125,N_4276);
nand U4626 (N_4626,N_3375,N_3815);
and U4627 (N_4627,N_3711,N_3732);
nand U4628 (N_4628,N_4360,N_3967);
nor U4629 (N_4629,N_4016,N_3279);
or U4630 (N_4630,N_3440,N_3604);
nor U4631 (N_4631,N_3969,N_4469);
nand U4632 (N_4632,N_4027,N_3250);
nand U4633 (N_4633,N_3897,N_3245);
nor U4634 (N_4634,N_3395,N_3999);
or U4635 (N_4635,N_4204,N_3923);
and U4636 (N_4636,N_4001,N_3869);
nor U4637 (N_4637,N_4456,N_3251);
and U4638 (N_4638,N_3779,N_3182);
xor U4639 (N_4639,N_3499,N_4072);
nor U4640 (N_4640,N_3875,N_4319);
or U4641 (N_4641,N_3822,N_3752);
nand U4642 (N_4642,N_3005,N_4274);
nand U4643 (N_4643,N_4328,N_3268);
or U4644 (N_4644,N_3446,N_4437);
or U4645 (N_4645,N_4235,N_4479);
nor U4646 (N_4646,N_3304,N_4092);
nor U4647 (N_4647,N_4230,N_4011);
or U4648 (N_4648,N_3707,N_3545);
and U4649 (N_4649,N_4310,N_3951);
nor U4650 (N_4650,N_4233,N_4252);
nand U4651 (N_4651,N_4246,N_3373);
xnor U4652 (N_4652,N_4336,N_3808);
xor U4653 (N_4653,N_3409,N_4403);
nand U4654 (N_4654,N_3099,N_3625);
nor U4655 (N_4655,N_4044,N_3952);
nor U4656 (N_4656,N_3254,N_3509);
and U4657 (N_4657,N_4443,N_3269);
nor U4658 (N_4658,N_3060,N_3233);
nor U4659 (N_4659,N_3194,N_3981);
xnor U4660 (N_4660,N_3885,N_4409);
nor U4661 (N_4661,N_3616,N_4490);
xnor U4662 (N_4662,N_4014,N_3048);
and U4663 (N_4663,N_4345,N_3964);
nor U4664 (N_4664,N_3249,N_4322);
nor U4665 (N_4665,N_3621,N_4305);
or U4666 (N_4666,N_3316,N_4163);
xnor U4667 (N_4667,N_3108,N_3890);
nor U4668 (N_4668,N_3016,N_3896);
nor U4669 (N_4669,N_3744,N_3832);
and U4670 (N_4670,N_3402,N_4146);
or U4671 (N_4671,N_3003,N_3789);
or U4672 (N_4672,N_4226,N_3295);
nand U4673 (N_4673,N_3338,N_3028);
nor U4674 (N_4674,N_3356,N_3168);
and U4675 (N_4675,N_4325,N_4300);
nand U4676 (N_4676,N_3800,N_4024);
or U4677 (N_4677,N_4426,N_4266);
and U4678 (N_4678,N_4341,N_4467);
nand U4679 (N_4679,N_4279,N_4416);
nand U4680 (N_4680,N_3510,N_3371);
nor U4681 (N_4681,N_4224,N_4242);
and U4682 (N_4682,N_3810,N_3697);
or U4683 (N_4683,N_3159,N_3565);
and U4684 (N_4684,N_3502,N_4497);
nor U4685 (N_4685,N_4002,N_3215);
nor U4686 (N_4686,N_3023,N_3666);
nand U4687 (N_4687,N_4361,N_4402);
and U4688 (N_4688,N_4422,N_4135);
and U4689 (N_4689,N_3612,N_3846);
and U4690 (N_4690,N_4308,N_4172);
xor U4691 (N_4691,N_3645,N_3983);
and U4692 (N_4692,N_3725,N_3817);
and U4693 (N_4693,N_4141,N_3394);
nand U4694 (N_4694,N_3107,N_3406);
nand U4695 (N_4695,N_3374,N_4243);
or U4696 (N_4696,N_3533,N_3833);
or U4697 (N_4697,N_3583,N_3345);
xnor U4698 (N_4698,N_3586,N_3466);
and U4699 (N_4699,N_3447,N_3769);
nor U4700 (N_4700,N_4462,N_3208);
or U4701 (N_4701,N_3332,N_3346);
nor U4702 (N_4702,N_3853,N_3975);
nor U4703 (N_4703,N_4220,N_4309);
and U4704 (N_4704,N_3524,N_3296);
nor U4705 (N_4705,N_4006,N_4284);
nand U4706 (N_4706,N_3962,N_3839);
nand U4707 (N_4707,N_4031,N_3640);
and U4708 (N_4708,N_4099,N_3688);
nand U4709 (N_4709,N_4406,N_4464);
nor U4710 (N_4710,N_3467,N_4093);
nand U4711 (N_4711,N_4091,N_3378);
and U4712 (N_4712,N_3631,N_4245);
nand U4713 (N_4713,N_4494,N_4033);
nand U4714 (N_4714,N_3333,N_3360);
and U4715 (N_4715,N_3258,N_3738);
or U4716 (N_4716,N_4124,N_3188);
nand U4717 (N_4717,N_3038,N_3690);
or U4718 (N_4718,N_4064,N_3252);
xnor U4719 (N_4719,N_3754,N_3567);
or U4720 (N_4720,N_3337,N_3443);
nor U4721 (N_4721,N_3270,N_4263);
nand U4722 (N_4722,N_3639,N_3909);
and U4723 (N_4723,N_4267,N_4234);
xor U4724 (N_4724,N_3289,N_3522);
nand U4725 (N_4725,N_3191,N_3414);
and U4726 (N_4726,N_3963,N_4487);
nor U4727 (N_4727,N_3889,N_3859);
and U4728 (N_4728,N_3246,N_3911);
and U4729 (N_4729,N_3824,N_4213);
nor U4730 (N_4730,N_3577,N_3929);
xnor U4731 (N_4731,N_3696,N_4285);
xnor U4732 (N_4732,N_3922,N_4188);
nand U4733 (N_4733,N_3542,N_3381);
and U4734 (N_4734,N_3437,N_4147);
xnor U4735 (N_4735,N_4270,N_4355);
or U4736 (N_4736,N_4066,N_3303);
nand U4737 (N_4737,N_3227,N_3905);
and U4738 (N_4738,N_4201,N_4168);
xor U4739 (N_4739,N_4244,N_3663);
and U4740 (N_4740,N_4400,N_4162);
or U4741 (N_4741,N_3284,N_4435);
nor U4742 (N_4742,N_3598,N_3156);
nor U4743 (N_4743,N_3740,N_3899);
nand U4744 (N_4744,N_3122,N_4290);
nand U4745 (N_4745,N_4191,N_3461);
and U4746 (N_4746,N_4100,N_3996);
and U4747 (N_4747,N_3844,N_3687);
nand U4748 (N_4748,N_4110,N_3543);
xnor U4749 (N_4749,N_4394,N_4190);
and U4750 (N_4750,N_3610,N_4181);
or U4751 (N_4751,N_3401,N_3307);
nor U4752 (N_4752,N_4392,N_3410);
or U4753 (N_4753,N_4003,N_4068);
nand U4754 (N_4754,N_4292,N_3788);
nor U4755 (N_4755,N_4206,N_4211);
and U4756 (N_4756,N_4425,N_4106);
or U4757 (N_4757,N_3681,N_4177);
or U4758 (N_4758,N_3018,N_3508);
and U4759 (N_4759,N_3430,N_3165);
and U4760 (N_4760,N_4169,N_3849);
or U4761 (N_4761,N_4164,N_3065);
or U4762 (N_4762,N_3796,N_3780);
or U4763 (N_4763,N_3143,N_4069);
nor U4764 (N_4764,N_4199,N_4421);
nand U4765 (N_4765,N_3298,N_3731);
or U4766 (N_4766,N_4414,N_3441);
or U4767 (N_4767,N_3277,N_3513);
and U4768 (N_4768,N_4381,N_3668);
or U4769 (N_4769,N_3185,N_4484);
nand U4770 (N_4770,N_4445,N_3248);
nor U4771 (N_4771,N_3193,N_4432);
nand U4772 (N_4772,N_3044,N_4042);
or U4773 (N_4773,N_4465,N_3564);
and U4774 (N_4774,N_3998,N_3405);
and U4775 (N_4775,N_3451,N_3893);
or U4776 (N_4776,N_3002,N_3827);
nor U4777 (N_4777,N_3175,N_4009);
xnor U4778 (N_4778,N_3566,N_3935);
nor U4779 (N_4779,N_3945,N_4209);
or U4780 (N_4780,N_3618,N_3212);
and U4781 (N_4781,N_3271,N_3053);
and U4782 (N_4782,N_4396,N_4241);
nor U4783 (N_4783,N_3211,N_3877);
and U4784 (N_4784,N_3925,N_4133);
nor U4785 (N_4785,N_3392,N_3367);
and U4786 (N_4786,N_3762,N_3538);
and U4787 (N_4787,N_3840,N_3276);
xor U4788 (N_4788,N_3010,N_3642);
nand U4789 (N_4789,N_4048,N_3514);
or U4790 (N_4790,N_3110,N_4200);
nand U4791 (N_4791,N_3033,N_3705);
or U4792 (N_4792,N_3572,N_3009);
nand U4793 (N_4793,N_3674,N_3455);
or U4794 (N_4794,N_4295,N_4289);
and U4795 (N_4795,N_3847,N_4374);
and U4796 (N_4796,N_3596,N_3576);
and U4797 (N_4797,N_3314,N_3129);
or U4798 (N_4798,N_3563,N_3097);
nand U4799 (N_4799,N_3217,N_3049);
and U4800 (N_4800,N_3628,N_4035);
nand U4801 (N_4801,N_3237,N_3095);
and U4802 (N_4802,N_4303,N_3286);
or U4803 (N_4803,N_3988,N_3943);
nor U4804 (N_4804,N_3419,N_3149);
and U4805 (N_4805,N_4461,N_4283);
or U4806 (N_4806,N_3954,N_4180);
and U4807 (N_4807,N_4253,N_3758);
nor U4808 (N_4808,N_3664,N_3120);
xnor U4809 (N_4809,N_3921,N_3727);
nand U4810 (N_4810,N_4485,N_3944);
nand U4811 (N_4811,N_3070,N_3222);
nor U4812 (N_4812,N_4030,N_3851);
or U4813 (N_4813,N_3126,N_3861);
xnor U4814 (N_4814,N_4454,N_3876);
nor U4815 (N_4815,N_3721,N_3843);
or U4816 (N_4816,N_4123,N_4313);
and U4817 (N_4817,N_3912,N_3359);
xnor U4818 (N_4818,N_3179,N_3920);
or U4819 (N_4819,N_4412,N_3580);
and U4820 (N_4820,N_3627,N_3490);
and U4821 (N_4821,N_3329,N_4250);
nand U4822 (N_4822,N_3763,N_4017);
nand U4823 (N_4823,N_3783,N_3858);
or U4824 (N_4824,N_3313,N_3936);
nor U4825 (N_4825,N_3012,N_3158);
and U4826 (N_4826,N_4137,N_3238);
or U4827 (N_4827,N_4228,N_3326);
and U4828 (N_4828,N_4473,N_3928);
xnor U4829 (N_4829,N_4413,N_3506);
or U4830 (N_4830,N_4311,N_3398);
nor U4831 (N_4831,N_3544,N_3101);
or U4832 (N_4832,N_3723,N_3892);
nor U4833 (N_4833,N_4386,N_3585);
nand U4834 (N_4834,N_4475,N_4020);
nor U4835 (N_4835,N_4185,N_4111);
or U4836 (N_4836,N_3066,N_3914);
and U4837 (N_4837,N_3090,N_4132);
xor U4838 (N_4838,N_3904,N_3865);
or U4839 (N_4839,N_4061,N_4306);
nor U4840 (N_4840,N_3464,N_4471);
or U4841 (N_4841,N_4216,N_3813);
nor U4842 (N_4842,N_4281,N_3742);
nand U4843 (N_4843,N_3775,N_3614);
nor U4844 (N_4844,N_4095,N_3647);
or U4845 (N_4845,N_3515,N_4021);
nand U4846 (N_4846,N_3884,N_3807);
nor U4847 (N_4847,N_3946,N_4463);
and U4848 (N_4848,N_3966,N_3794);
and U4849 (N_4849,N_3700,N_3327);
nand U4850 (N_4850,N_3051,N_3816);
and U4851 (N_4851,N_3679,N_4258);
nand U4852 (N_4852,N_3540,N_3716);
nand U4853 (N_4853,N_4107,N_3651);
or U4854 (N_4854,N_3646,N_4419);
xor U4855 (N_4855,N_4271,N_4451);
xnor U4856 (N_4856,N_3294,N_4450);
or U4857 (N_4857,N_3117,N_3624);
nor U4858 (N_4858,N_4417,N_3818);
nor U4859 (N_4859,N_3504,N_4430);
and U4860 (N_4860,N_3334,N_3868);
or U4861 (N_4861,N_3112,N_3138);
and U4862 (N_4862,N_3103,N_3848);
nand U4863 (N_4863,N_3137,N_4126);
or U4864 (N_4864,N_4117,N_3562);
or U4865 (N_4865,N_3582,N_3825);
or U4866 (N_4866,N_3302,N_3695);
nand U4867 (N_4867,N_4348,N_3280);
xnor U4868 (N_4868,N_4165,N_3617);
or U4869 (N_4869,N_4476,N_3427);
or U4870 (N_4870,N_4247,N_3069);
xnor U4871 (N_4871,N_3113,N_4314);
nand U4872 (N_4872,N_3234,N_3089);
nand U4873 (N_4873,N_3037,N_4125);
nand U4874 (N_4874,N_3426,N_4299);
xnor U4875 (N_4875,N_3672,N_3421);
nor U4876 (N_4876,N_4438,N_3555);
nand U4877 (N_4877,N_3760,N_3654);
nor U4878 (N_4878,N_3355,N_4366);
nand U4879 (N_4879,N_3384,N_4418);
nor U4880 (N_4880,N_4214,N_3556);
and U4881 (N_4881,N_4362,N_3759);
nor U4882 (N_4882,N_3014,N_4282);
nor U4883 (N_4883,N_3181,N_3199);
and U4884 (N_4884,N_3665,N_3559);
xor U4885 (N_4885,N_4223,N_3106);
nand U4886 (N_4886,N_3866,N_3613);
nor U4887 (N_4887,N_3494,N_3096);
or U4888 (N_4888,N_3218,N_4130);
and U4889 (N_4889,N_4411,N_3821);
or U4890 (N_4890,N_3080,N_3253);
nand U4891 (N_4891,N_3829,N_4187);
or U4892 (N_4892,N_4070,N_4329);
nor U4893 (N_4893,N_3147,N_3006);
and U4894 (N_4894,N_3749,N_4151);
nand U4895 (N_4895,N_4262,N_3008);
or U4896 (N_4896,N_3855,N_4018);
nand U4897 (N_4897,N_3476,N_4264);
nand U4898 (N_4898,N_3841,N_3084);
nand U4899 (N_4899,N_4154,N_3036);
and U4900 (N_4900,N_3990,N_3281);
nand U4901 (N_4901,N_3104,N_3052);
nor U4902 (N_4902,N_4028,N_3433);
nor U4903 (N_4903,N_4179,N_3452);
nand U4904 (N_4904,N_3236,N_4317);
or U4905 (N_4905,N_3871,N_3706);
and U4906 (N_4906,N_3264,N_4470);
nand U4907 (N_4907,N_3240,N_3267);
or U4908 (N_4908,N_4398,N_3418);
or U4909 (N_4909,N_4065,N_3256);
or U4910 (N_4910,N_3934,N_4122);
xnor U4911 (N_4911,N_3527,N_3644);
or U4912 (N_4912,N_3232,N_4036);
nand U4913 (N_4913,N_4007,N_4382);
and U4914 (N_4914,N_3734,N_4269);
or U4915 (N_4915,N_3802,N_3694);
nor U4916 (N_4916,N_3660,N_4458);
nor U4917 (N_4917,N_4293,N_3205);
nand U4918 (N_4918,N_3692,N_3656);
or U4919 (N_4919,N_4440,N_3261);
and U4920 (N_4920,N_3907,N_3026);
nor U4921 (N_4921,N_4210,N_3413);
and U4922 (N_4922,N_4442,N_3109);
xor U4923 (N_4923,N_3152,N_3611);
xor U4924 (N_4924,N_4073,N_3436);
nor U4925 (N_4925,N_3465,N_3431);
and U4926 (N_4926,N_3093,N_4145);
or U4927 (N_4927,N_4118,N_3776);
nand U4928 (N_4928,N_4040,N_4198);
and U4929 (N_4929,N_4189,N_4318);
nand U4930 (N_4930,N_3579,N_3919);
or U4931 (N_4931,N_3857,N_3130);
xnor U4932 (N_4932,N_3291,N_3278);
or U4933 (N_4933,N_3746,N_3891);
nand U4934 (N_4934,N_3630,N_3174);
nand U4935 (N_4935,N_3778,N_3994);
nor U4936 (N_4936,N_3056,N_3075);
nor U4937 (N_4937,N_4157,N_3220);
nor U4938 (N_4938,N_4408,N_3819);
or U4939 (N_4939,N_3231,N_3047);
nand U4940 (N_4940,N_4433,N_3751);
and U4941 (N_4941,N_3924,N_4171);
nor U4942 (N_4942,N_4205,N_4272);
nor U4943 (N_4943,N_3391,N_3675);
and U4944 (N_4944,N_4369,N_3098);
and U4945 (N_4945,N_4373,N_4477);
nor U4946 (N_4946,N_4217,N_3417);
and U4947 (N_4947,N_3685,N_3260);
nor U4948 (N_4948,N_3163,N_3034);
nor U4949 (N_4949,N_4129,N_4173);
nor U4950 (N_4950,N_3867,N_3351);
nor U4951 (N_4951,N_4323,N_4176);
or U4952 (N_4952,N_3386,N_3872);
nor U4953 (N_4953,N_3856,N_4221);
nor U4954 (N_4954,N_3407,N_3767);
nand U4955 (N_4955,N_4371,N_3535);
or U4956 (N_4956,N_4291,N_3161);
or U4957 (N_4957,N_3140,N_4212);
nor U4958 (N_4958,N_3349,N_4085);
nand U4959 (N_4959,N_3546,N_3242);
and U4960 (N_4960,N_3811,N_3145);
and U4961 (N_4961,N_3773,N_4460);
and U4962 (N_4962,N_3067,N_3471);
or U4963 (N_4963,N_3042,N_3330);
or U4964 (N_4964,N_4261,N_4420);
nand U4965 (N_4965,N_4225,N_3837);
xnor U4966 (N_4966,N_3393,N_3938);
or U4967 (N_4967,N_4287,N_3852);
and U4968 (N_4968,N_4448,N_3342);
nand U4969 (N_4969,N_4094,N_4256);
nand U4970 (N_4970,N_4365,N_3883);
or U4971 (N_4971,N_4041,N_3836);
nor U4972 (N_4972,N_3162,N_3714);
or U4973 (N_4973,N_3698,N_3463);
or U4974 (N_4974,N_4321,N_3335);
and U4975 (N_4975,N_4375,N_4431);
nor U4976 (N_4976,N_3274,N_3551);
nor U4977 (N_4977,N_3602,N_3530);
nor U4978 (N_4978,N_3753,N_4482);
nand U4979 (N_4979,N_4062,N_3364);
nor U4980 (N_4980,N_3331,N_3532);
and U4981 (N_4981,N_3166,N_3790);
and U4982 (N_4982,N_3321,N_4056);
nor U4983 (N_4983,N_3453,N_4280);
nand U4984 (N_4984,N_4184,N_3219);
or U4985 (N_4985,N_3071,N_3146);
and U4986 (N_4986,N_3623,N_3957);
nand U4987 (N_4987,N_4391,N_4158);
nand U4988 (N_4988,N_3265,N_3915);
xor U4989 (N_4989,N_3244,N_4452);
xor U4990 (N_4990,N_3136,N_3560);
or U4991 (N_4991,N_3448,N_4000);
nand U4992 (N_4992,N_4468,N_3702);
nor U4993 (N_4993,N_3412,N_3989);
and U4994 (N_4994,N_3474,N_3500);
and U4995 (N_4995,N_3638,N_4273);
nor U4996 (N_4996,N_3141,N_4131);
nor U4997 (N_4997,N_4196,N_3626);
or U4998 (N_4998,N_4127,N_3312);
xor U4999 (N_4999,N_3282,N_3491);
nor U5000 (N_5000,N_3803,N_3272);
or U5001 (N_5001,N_4496,N_4466);
nor U5002 (N_5002,N_3797,N_4240);
nand U5003 (N_5003,N_3480,N_3216);
nand U5004 (N_5004,N_3128,N_3571);
and U5005 (N_5005,N_3710,N_3083);
nor U5006 (N_5006,N_3257,N_4054);
nand U5007 (N_5007,N_3641,N_3403);
nand U5008 (N_5008,N_4012,N_3336);
nand U5009 (N_5009,N_4459,N_3823);
and U5010 (N_5010,N_4112,N_4342);
nand U5011 (N_5011,N_3428,N_3206);
nand U5012 (N_5012,N_4363,N_3686);
nor U5013 (N_5013,N_4139,N_4254);
nand U5014 (N_5014,N_3160,N_3173);
and U5015 (N_5015,N_3956,N_4453);
or U5016 (N_5016,N_3634,N_3678);
and U5017 (N_5017,N_3011,N_3362);
or U5018 (N_5018,N_3172,N_3661);
or U5019 (N_5019,N_3186,N_3558);
and U5020 (N_5020,N_4429,N_4104);
and U5021 (N_5021,N_4077,N_3170);
or U5022 (N_5022,N_3607,N_3416);
or U5023 (N_5023,N_3197,N_3133);
nand U5024 (N_5024,N_4032,N_4286);
xor U5025 (N_5025,N_3111,N_3323);
xnor U5026 (N_5026,N_3547,N_3063);
nor U5027 (N_5027,N_4115,N_3930);
nor U5028 (N_5028,N_3953,N_3970);
and U5029 (N_5029,N_4304,N_4167);
or U5030 (N_5030,N_4278,N_3704);
nor U5031 (N_5031,N_4083,N_3035);
nor U5032 (N_5032,N_4142,N_3458);
or U5033 (N_5033,N_3709,N_4316);
nand U5034 (N_5034,N_4379,N_3902);
and U5035 (N_5035,N_3040,N_3007);
or U5036 (N_5036,N_4298,N_3518);
nand U5037 (N_5037,N_4397,N_3781);
or U5038 (N_5038,N_3087,N_4170);
xor U5039 (N_5039,N_3230,N_4354);
or U5040 (N_5040,N_3838,N_3318);
and U5041 (N_5041,N_3961,N_4178);
nand U5042 (N_5042,N_4120,N_4495);
nand U5043 (N_5043,N_4113,N_3910);
or U5044 (N_5044,N_4034,N_3397);
and U5045 (N_5045,N_3139,N_3673);
or U5046 (N_5046,N_4236,N_3239);
nor U5047 (N_5047,N_4023,N_4096);
xnor U5048 (N_5048,N_3680,N_3528);
nand U5049 (N_5049,N_3503,N_3132);
xor U5050 (N_5050,N_3908,N_4257);
nor U5051 (N_5051,N_3155,N_3456);
xor U5052 (N_5052,N_4071,N_4330);
nor U5053 (N_5053,N_4192,N_3459);
nor U5054 (N_5054,N_4315,N_3862);
and U5055 (N_5055,N_4268,N_3939);
and U5056 (N_5056,N_3552,N_3203);
xnor U5057 (N_5057,N_3144,N_3348);
or U5058 (N_5058,N_3404,N_3498);
xor U5059 (N_5059,N_3870,N_3830);
or U5060 (N_5060,N_3756,N_4060);
nand U5061 (N_5061,N_3755,N_4153);
xor U5062 (N_5062,N_3435,N_3573);
and U5063 (N_5063,N_4022,N_4353);
or U5064 (N_5064,N_4277,N_3782);
or U5065 (N_5065,N_3768,N_3519);
and U5066 (N_5066,N_3873,N_3062);
nor U5067 (N_5067,N_4160,N_3479);
nor U5068 (N_5068,N_3933,N_3226);
and U5069 (N_5069,N_3512,N_4427);
and U5070 (N_5070,N_4116,N_3592);
or U5071 (N_5071,N_4493,N_3116);
xnor U5072 (N_5072,N_3309,N_3526);
or U5073 (N_5073,N_3761,N_3880);
nand U5074 (N_5074,N_4488,N_3273);
xor U5075 (N_5075,N_3180,N_4057);
nor U5076 (N_5076,N_3667,N_3082);
and U5077 (N_5077,N_4447,N_4446);
or U5078 (N_5078,N_3420,N_3669);
nand U5079 (N_5079,N_3801,N_3594);
and U5080 (N_5080,N_3442,N_3941);
xnor U5081 (N_5081,N_4352,N_4227);
or U5082 (N_5082,N_4357,N_4238);
nor U5083 (N_5083,N_4455,N_3835);
or U5084 (N_5084,N_4364,N_4296);
or U5085 (N_5085,N_4098,N_3712);
nor U5086 (N_5086,N_3454,N_3411);
nor U5087 (N_5087,N_3470,N_3699);
and U5088 (N_5088,N_3347,N_4334);
and U5089 (N_5089,N_3225,N_4087);
and U5090 (N_5090,N_3377,N_3888);
and U5091 (N_5091,N_3308,N_3799);
xnor U5092 (N_5092,N_3658,N_3100);
and U5093 (N_5093,N_3978,N_3534);
xor U5094 (N_5094,N_3025,N_3305);
nand U5095 (N_5095,N_3064,N_3045);
xor U5096 (N_5096,N_3619,N_3283);
and U5097 (N_5097,N_3019,N_4152);
nand U5098 (N_5098,N_4340,N_3599);
or U5099 (N_5099,N_3057,N_3196);
or U5100 (N_5100,N_4102,N_4351);
nand U5101 (N_5101,N_4019,N_3221);
xnor U5102 (N_5102,N_3387,N_4265);
or U5103 (N_5103,N_3195,N_4327);
nand U5104 (N_5104,N_3190,N_3505);
and U5105 (N_5105,N_4489,N_3372);
nand U5106 (N_5106,N_3881,N_3266);
nand U5107 (N_5107,N_4441,N_3724);
xor U5108 (N_5108,N_3950,N_3396);
and U5109 (N_5109,N_3659,N_4404);
nor U5110 (N_5110,N_3142,N_3322);
and U5111 (N_5111,N_3831,N_3864);
nand U5112 (N_5112,N_3820,N_4079);
nand U5113 (N_5113,N_4385,N_3785);
or U5114 (N_5114,N_4182,N_3992);
nor U5115 (N_5115,N_3845,N_3548);
nand U5116 (N_5116,N_4082,N_3854);
and U5117 (N_5117,N_4088,N_4202);
xor U5118 (N_5118,N_4288,N_3306);
xor U5119 (N_5119,N_4424,N_4444);
nor U5120 (N_5120,N_3806,N_3354);
xor U5121 (N_5121,N_3460,N_3317);
nand U5122 (N_5122,N_3439,N_4193);
nand U5123 (N_5123,N_3119,N_3425);
nor U5124 (N_5124,N_3557,N_3275);
nand U5125 (N_5125,N_4407,N_4499);
or U5126 (N_5126,N_4084,N_3737);
nand U5127 (N_5127,N_3593,N_3115);
nand U5128 (N_5128,N_3483,N_3153);
or U5129 (N_5129,N_4138,N_3529);
nand U5130 (N_5130,N_3733,N_3874);
or U5131 (N_5131,N_3828,N_3581);
or U5132 (N_5132,N_3328,N_4046);
nand U5133 (N_5133,N_3917,N_3444);
xor U5134 (N_5134,N_4174,N_3088);
or U5135 (N_5135,N_3648,N_3297);
xor U5136 (N_5136,N_3077,N_3792);
nand U5137 (N_5137,N_3475,N_3574);
or U5138 (N_5138,N_4332,N_3708);
xnor U5139 (N_5139,N_4175,N_3457);
nand U5140 (N_5140,N_3496,N_3587);
xnor U5141 (N_5141,N_3520,N_3554);
nor U5142 (N_5142,N_3091,N_3123);
and U5143 (N_5143,N_3793,N_3255);
or U5144 (N_5144,N_3207,N_4372);
or U5145 (N_5145,N_3927,N_3622);
nor U5146 (N_5146,N_3684,N_3114);
and U5147 (N_5147,N_4004,N_4161);
or U5148 (N_5148,N_4166,N_4326);
and U5149 (N_5149,N_3485,N_3882);
xor U5150 (N_5150,N_3154,N_3055);
nor U5151 (N_5151,N_4078,N_3399);
nand U5152 (N_5152,N_4383,N_3748);
and U5153 (N_5153,N_3368,N_3177);
nand U5154 (N_5154,N_3812,N_4410);
xor U5155 (N_5155,N_3601,N_3029);
and U5156 (N_5156,N_4349,N_3247);
or U5157 (N_5157,N_3670,N_4231);
and U5158 (N_5158,N_3531,N_4359);
or U5159 (N_5159,N_4337,N_3102);
or U5160 (N_5160,N_3486,N_4399);
and U5161 (N_5161,N_3164,N_3507);
and U5162 (N_5162,N_3020,N_4275);
nand U5163 (N_5163,N_3553,N_3974);
nor U5164 (N_5164,N_3947,N_3415);
and U5165 (N_5165,N_3913,N_3517);
nand U5166 (N_5166,N_3127,N_3050);
nor U5167 (N_5167,N_3662,N_4472);
or U5168 (N_5168,N_3134,N_3987);
nand U5169 (N_5169,N_3791,N_3887);
nand U5170 (N_5170,N_4498,N_4043);
and U5171 (N_5171,N_3777,N_3689);
nor U5172 (N_5172,N_3677,N_3595);
nand U5173 (N_5173,N_3487,N_3569);
or U5174 (N_5174,N_4347,N_4387);
nand U5175 (N_5175,N_3886,N_3438);
nor U5176 (N_5176,N_3481,N_3683);
nor U5177 (N_5177,N_4390,N_3942);
nor U5178 (N_5178,N_4229,N_3178);
nor U5179 (N_5179,N_4128,N_3906);
nand U5180 (N_5180,N_3209,N_3320);
xnor U5181 (N_5181,N_3575,N_3620);
nand U5182 (N_5182,N_3151,N_3750);
and U5183 (N_5183,N_4331,N_4474);
nor U5184 (N_5184,N_3445,N_3073);
nand U5185 (N_5185,N_3324,N_3657);
nor U5186 (N_5186,N_3898,N_3691);
nor U5187 (N_5187,N_4047,N_4380);
nor U5188 (N_5188,N_4101,N_4194);
nor U5189 (N_5189,N_3703,N_3878);
nor U5190 (N_5190,N_4074,N_3774);
nor U5191 (N_5191,N_4150,N_4081);
and U5192 (N_5192,N_3940,N_3541);
xnor U5193 (N_5193,N_4114,N_3653);
or U5194 (N_5194,N_3635,N_3243);
xor U5195 (N_5195,N_3389,N_4312);
and U5196 (N_5196,N_4039,N_4248);
nor U5197 (N_5197,N_3991,N_3984);
nor U5198 (N_5198,N_3039,N_3183);
nor U5199 (N_5199,N_3004,N_3429);
or U5200 (N_5200,N_4307,N_3422);
or U5201 (N_5201,N_3472,N_3591);
nand U5202 (N_5202,N_3719,N_3319);
or U5203 (N_5203,N_3361,N_3363);
and U5204 (N_5204,N_3202,N_3030);
and U5205 (N_5205,N_3959,N_3325);
or U5206 (N_5206,N_3015,N_4186);
nor U5207 (N_5207,N_4389,N_3353);
or U5208 (N_5208,N_4449,N_4026);
or U5209 (N_5209,N_3901,N_3918);
nand U5210 (N_5210,N_4302,N_3895);
nand U5211 (N_5211,N_3383,N_4051);
or U5212 (N_5212,N_3078,N_3027);
and U5213 (N_5213,N_3568,N_4237);
nand U5214 (N_5214,N_4155,N_4415);
nand U5215 (N_5215,N_3764,N_4013);
nor U5216 (N_5216,N_4097,N_4121);
nor U5217 (N_5217,N_3118,N_3973);
nand U5218 (N_5218,N_3382,N_3000);
or U5219 (N_5219,N_3041,N_3024);
or U5220 (N_5220,N_4405,N_4008);
or U5221 (N_5221,N_3340,N_3632);
and U5222 (N_5222,N_3492,N_3380);
or U5223 (N_5223,N_3369,N_3352);
nor U5224 (N_5224,N_4478,N_3478);
nand U5225 (N_5225,N_3477,N_3157);
nor U5226 (N_5226,N_3916,N_3469);
nor U5227 (N_5227,N_3285,N_3637);
or U5228 (N_5228,N_3204,N_3495);
or U5229 (N_5229,N_3516,N_3804);
nand U5230 (N_5230,N_4239,N_3589);
and U5231 (N_5231,N_4108,N_3184);
and U5232 (N_5232,N_3343,N_3629);
or U5233 (N_5233,N_3814,N_3745);
xnor U5234 (N_5234,N_4339,N_4075);
or U5235 (N_5235,N_3787,N_3001);
or U5236 (N_5236,N_3187,N_3722);
nand U5237 (N_5237,N_3770,N_3960);
and U5238 (N_5238,N_4358,N_3059);
nand U5239 (N_5239,N_4320,N_3228);
nand U5240 (N_5240,N_4368,N_3124);
and U5241 (N_5241,N_4063,N_3766);
or U5242 (N_5242,N_3850,N_3949);
nand U5243 (N_5243,N_3105,N_4260);
nor U5244 (N_5244,N_4480,N_3985);
nor U5245 (N_5245,N_3135,N_3521);
xnor U5246 (N_5246,N_3290,N_4384);
and U5247 (N_5247,N_3223,N_3339);
nand U5248 (N_5248,N_3717,N_3894);
nand U5249 (N_5249,N_3739,N_3076);
or U5250 (N_5250,N_3399,N_3400);
or U5251 (N_5251,N_4444,N_4335);
nand U5252 (N_5252,N_3297,N_3607);
nor U5253 (N_5253,N_4163,N_4147);
nand U5254 (N_5254,N_3906,N_3392);
or U5255 (N_5255,N_3010,N_3689);
nor U5256 (N_5256,N_3970,N_3377);
nand U5257 (N_5257,N_4277,N_3173);
nand U5258 (N_5258,N_3308,N_3598);
and U5259 (N_5259,N_3063,N_3621);
and U5260 (N_5260,N_4440,N_4277);
nor U5261 (N_5261,N_4311,N_3686);
nor U5262 (N_5262,N_3751,N_3226);
and U5263 (N_5263,N_4415,N_4177);
nor U5264 (N_5264,N_3221,N_3066);
or U5265 (N_5265,N_3774,N_3835);
and U5266 (N_5266,N_4277,N_3997);
or U5267 (N_5267,N_3423,N_4078);
or U5268 (N_5268,N_3455,N_4437);
and U5269 (N_5269,N_4458,N_3948);
and U5270 (N_5270,N_4277,N_4466);
or U5271 (N_5271,N_3197,N_3641);
xnor U5272 (N_5272,N_4396,N_4014);
nand U5273 (N_5273,N_3289,N_3319);
and U5274 (N_5274,N_3733,N_4440);
nor U5275 (N_5275,N_3540,N_3992);
or U5276 (N_5276,N_3028,N_3520);
nor U5277 (N_5277,N_3083,N_3317);
nor U5278 (N_5278,N_3410,N_3394);
and U5279 (N_5279,N_3431,N_3562);
nand U5280 (N_5280,N_3112,N_3562);
or U5281 (N_5281,N_3456,N_3855);
and U5282 (N_5282,N_4245,N_3892);
nor U5283 (N_5283,N_3356,N_3980);
nand U5284 (N_5284,N_4420,N_4287);
and U5285 (N_5285,N_3717,N_3789);
and U5286 (N_5286,N_3598,N_3442);
xnor U5287 (N_5287,N_3037,N_3434);
or U5288 (N_5288,N_3971,N_4106);
nand U5289 (N_5289,N_4239,N_3815);
nor U5290 (N_5290,N_4013,N_4051);
and U5291 (N_5291,N_3918,N_3762);
and U5292 (N_5292,N_3135,N_4273);
and U5293 (N_5293,N_3786,N_3880);
and U5294 (N_5294,N_4233,N_3180);
nand U5295 (N_5295,N_3532,N_3929);
and U5296 (N_5296,N_4148,N_3667);
and U5297 (N_5297,N_3166,N_3531);
nand U5298 (N_5298,N_3171,N_3927);
nand U5299 (N_5299,N_3455,N_3059);
nor U5300 (N_5300,N_3905,N_3330);
or U5301 (N_5301,N_3542,N_4114);
xor U5302 (N_5302,N_3790,N_3953);
nor U5303 (N_5303,N_4155,N_3545);
nand U5304 (N_5304,N_3969,N_4146);
nor U5305 (N_5305,N_4251,N_3469);
nand U5306 (N_5306,N_4383,N_3632);
nor U5307 (N_5307,N_3741,N_3240);
nor U5308 (N_5308,N_4338,N_3802);
or U5309 (N_5309,N_3789,N_3167);
or U5310 (N_5310,N_3302,N_4112);
and U5311 (N_5311,N_3294,N_3308);
and U5312 (N_5312,N_3851,N_4389);
or U5313 (N_5313,N_4224,N_4110);
and U5314 (N_5314,N_3345,N_4421);
xnor U5315 (N_5315,N_3329,N_4477);
and U5316 (N_5316,N_4353,N_4319);
nand U5317 (N_5317,N_4494,N_3385);
or U5318 (N_5318,N_3111,N_4380);
or U5319 (N_5319,N_4422,N_3535);
nor U5320 (N_5320,N_3360,N_4216);
nor U5321 (N_5321,N_3270,N_3573);
or U5322 (N_5322,N_3489,N_4484);
and U5323 (N_5323,N_3934,N_3917);
and U5324 (N_5324,N_3938,N_4046);
nor U5325 (N_5325,N_3699,N_3213);
or U5326 (N_5326,N_3006,N_3607);
nor U5327 (N_5327,N_3829,N_4071);
or U5328 (N_5328,N_3770,N_3512);
or U5329 (N_5329,N_3555,N_3905);
or U5330 (N_5330,N_3537,N_3950);
nor U5331 (N_5331,N_4460,N_3151);
xnor U5332 (N_5332,N_3004,N_3339);
or U5333 (N_5333,N_3939,N_4035);
or U5334 (N_5334,N_3102,N_3330);
and U5335 (N_5335,N_3358,N_3910);
nand U5336 (N_5336,N_3274,N_3618);
nor U5337 (N_5337,N_3732,N_3934);
nor U5338 (N_5338,N_3220,N_3319);
nand U5339 (N_5339,N_3359,N_4417);
or U5340 (N_5340,N_3280,N_3939);
nor U5341 (N_5341,N_3195,N_3105);
or U5342 (N_5342,N_3087,N_3937);
nor U5343 (N_5343,N_3797,N_3067);
or U5344 (N_5344,N_3516,N_4297);
or U5345 (N_5345,N_4244,N_3556);
nor U5346 (N_5346,N_3573,N_3394);
xnor U5347 (N_5347,N_3920,N_3711);
nor U5348 (N_5348,N_3137,N_3812);
nand U5349 (N_5349,N_3607,N_3983);
nor U5350 (N_5350,N_4477,N_4160);
and U5351 (N_5351,N_3278,N_3461);
or U5352 (N_5352,N_4478,N_3926);
nor U5353 (N_5353,N_3732,N_3350);
nand U5354 (N_5354,N_4345,N_4107);
or U5355 (N_5355,N_4254,N_3805);
nand U5356 (N_5356,N_4237,N_4478);
or U5357 (N_5357,N_3260,N_3266);
nand U5358 (N_5358,N_4149,N_4122);
nand U5359 (N_5359,N_4243,N_3013);
nand U5360 (N_5360,N_4048,N_3922);
or U5361 (N_5361,N_3726,N_4462);
nor U5362 (N_5362,N_3919,N_3058);
xnor U5363 (N_5363,N_3619,N_3229);
or U5364 (N_5364,N_3914,N_3002);
or U5365 (N_5365,N_4278,N_4448);
or U5366 (N_5366,N_3252,N_3367);
and U5367 (N_5367,N_4429,N_4318);
nand U5368 (N_5368,N_3635,N_3707);
and U5369 (N_5369,N_3416,N_4222);
and U5370 (N_5370,N_4260,N_3230);
or U5371 (N_5371,N_3147,N_4042);
or U5372 (N_5372,N_3181,N_3694);
nor U5373 (N_5373,N_3427,N_3951);
and U5374 (N_5374,N_3985,N_3253);
nand U5375 (N_5375,N_3991,N_4117);
nor U5376 (N_5376,N_3500,N_3948);
nand U5377 (N_5377,N_4452,N_3569);
or U5378 (N_5378,N_3609,N_4396);
and U5379 (N_5379,N_3575,N_4065);
xnor U5380 (N_5380,N_3095,N_3880);
and U5381 (N_5381,N_3180,N_3159);
nor U5382 (N_5382,N_3974,N_3478);
and U5383 (N_5383,N_4246,N_3079);
nor U5384 (N_5384,N_3793,N_3691);
and U5385 (N_5385,N_3091,N_4237);
or U5386 (N_5386,N_4155,N_3926);
or U5387 (N_5387,N_4135,N_3461);
or U5388 (N_5388,N_3016,N_4046);
nand U5389 (N_5389,N_3029,N_4121);
and U5390 (N_5390,N_4477,N_3998);
and U5391 (N_5391,N_3628,N_3263);
or U5392 (N_5392,N_3554,N_4260);
or U5393 (N_5393,N_4013,N_3362);
and U5394 (N_5394,N_4399,N_4075);
and U5395 (N_5395,N_3085,N_3156);
and U5396 (N_5396,N_3430,N_3639);
or U5397 (N_5397,N_3157,N_3774);
nor U5398 (N_5398,N_3451,N_4044);
or U5399 (N_5399,N_3770,N_4122);
nor U5400 (N_5400,N_3119,N_4351);
or U5401 (N_5401,N_4123,N_4278);
nor U5402 (N_5402,N_3109,N_4180);
and U5403 (N_5403,N_3620,N_3804);
nor U5404 (N_5404,N_3511,N_3469);
or U5405 (N_5405,N_4084,N_3439);
nor U5406 (N_5406,N_3986,N_3506);
nand U5407 (N_5407,N_4369,N_4370);
or U5408 (N_5408,N_3513,N_3858);
and U5409 (N_5409,N_4342,N_3137);
or U5410 (N_5410,N_4145,N_4493);
and U5411 (N_5411,N_4479,N_4393);
or U5412 (N_5412,N_4062,N_3062);
nand U5413 (N_5413,N_3401,N_3377);
and U5414 (N_5414,N_4304,N_4445);
xnor U5415 (N_5415,N_3967,N_3466);
or U5416 (N_5416,N_3485,N_3109);
nor U5417 (N_5417,N_3712,N_3038);
or U5418 (N_5418,N_3810,N_4071);
and U5419 (N_5419,N_3786,N_3471);
nor U5420 (N_5420,N_4182,N_4486);
nor U5421 (N_5421,N_4363,N_3175);
or U5422 (N_5422,N_3515,N_3017);
and U5423 (N_5423,N_3945,N_3272);
nand U5424 (N_5424,N_3726,N_3796);
or U5425 (N_5425,N_3372,N_4063);
and U5426 (N_5426,N_3118,N_4034);
nor U5427 (N_5427,N_3211,N_3579);
nor U5428 (N_5428,N_3689,N_4382);
nor U5429 (N_5429,N_3468,N_3648);
and U5430 (N_5430,N_3296,N_4280);
nor U5431 (N_5431,N_3010,N_4303);
or U5432 (N_5432,N_3205,N_4018);
and U5433 (N_5433,N_3465,N_3069);
nor U5434 (N_5434,N_3286,N_3238);
or U5435 (N_5435,N_3396,N_3295);
and U5436 (N_5436,N_3704,N_3169);
and U5437 (N_5437,N_3828,N_4298);
or U5438 (N_5438,N_3112,N_3120);
and U5439 (N_5439,N_4374,N_4486);
and U5440 (N_5440,N_3999,N_4384);
and U5441 (N_5441,N_3954,N_4219);
and U5442 (N_5442,N_4343,N_3401);
and U5443 (N_5443,N_3955,N_3420);
or U5444 (N_5444,N_3105,N_3352);
nor U5445 (N_5445,N_3951,N_3093);
nor U5446 (N_5446,N_3683,N_4323);
and U5447 (N_5447,N_4166,N_3117);
or U5448 (N_5448,N_3885,N_4018);
and U5449 (N_5449,N_4322,N_4171);
nor U5450 (N_5450,N_3314,N_3340);
xor U5451 (N_5451,N_3059,N_3767);
nand U5452 (N_5452,N_3364,N_3854);
nor U5453 (N_5453,N_4207,N_3353);
or U5454 (N_5454,N_3478,N_3588);
nor U5455 (N_5455,N_3716,N_3538);
or U5456 (N_5456,N_3329,N_3944);
or U5457 (N_5457,N_3798,N_3325);
nand U5458 (N_5458,N_3860,N_3174);
or U5459 (N_5459,N_4378,N_4441);
xnor U5460 (N_5460,N_3876,N_3503);
nand U5461 (N_5461,N_4479,N_4340);
xor U5462 (N_5462,N_3282,N_4407);
nand U5463 (N_5463,N_3249,N_4004);
or U5464 (N_5464,N_3747,N_3156);
nor U5465 (N_5465,N_3551,N_4472);
nor U5466 (N_5466,N_3329,N_3062);
or U5467 (N_5467,N_3758,N_3552);
xor U5468 (N_5468,N_3694,N_4278);
nor U5469 (N_5469,N_4448,N_3558);
and U5470 (N_5470,N_3815,N_4054);
nor U5471 (N_5471,N_4192,N_3816);
xnor U5472 (N_5472,N_3697,N_4077);
nor U5473 (N_5473,N_4365,N_4252);
and U5474 (N_5474,N_3947,N_4234);
nand U5475 (N_5475,N_3927,N_4328);
xnor U5476 (N_5476,N_3528,N_3905);
or U5477 (N_5477,N_3198,N_3788);
or U5478 (N_5478,N_3970,N_3666);
or U5479 (N_5479,N_3294,N_4383);
nand U5480 (N_5480,N_4331,N_4343);
nor U5481 (N_5481,N_3734,N_3743);
and U5482 (N_5482,N_3610,N_3341);
nor U5483 (N_5483,N_4154,N_4123);
and U5484 (N_5484,N_3442,N_3659);
nand U5485 (N_5485,N_3152,N_3001);
and U5486 (N_5486,N_3882,N_3602);
nand U5487 (N_5487,N_4420,N_4369);
xor U5488 (N_5488,N_3590,N_4170);
and U5489 (N_5489,N_4165,N_4392);
nor U5490 (N_5490,N_4406,N_4438);
nor U5491 (N_5491,N_3848,N_3376);
and U5492 (N_5492,N_3812,N_4460);
nor U5493 (N_5493,N_4287,N_4338);
and U5494 (N_5494,N_3448,N_3931);
nand U5495 (N_5495,N_3448,N_4270);
or U5496 (N_5496,N_3358,N_4052);
or U5497 (N_5497,N_3303,N_3188);
or U5498 (N_5498,N_3590,N_3397);
or U5499 (N_5499,N_3939,N_3473);
xnor U5500 (N_5500,N_4411,N_4322);
or U5501 (N_5501,N_4092,N_4043);
nor U5502 (N_5502,N_4437,N_3832);
or U5503 (N_5503,N_3305,N_3389);
nor U5504 (N_5504,N_3386,N_3043);
nor U5505 (N_5505,N_3877,N_3703);
and U5506 (N_5506,N_4111,N_3126);
and U5507 (N_5507,N_3329,N_4442);
or U5508 (N_5508,N_3089,N_3724);
and U5509 (N_5509,N_4011,N_4357);
and U5510 (N_5510,N_3132,N_3153);
nand U5511 (N_5511,N_4078,N_4189);
xor U5512 (N_5512,N_4108,N_4166);
nand U5513 (N_5513,N_3286,N_4060);
and U5514 (N_5514,N_3144,N_3435);
or U5515 (N_5515,N_3360,N_3532);
nand U5516 (N_5516,N_3352,N_4398);
or U5517 (N_5517,N_3981,N_3628);
nor U5518 (N_5518,N_4456,N_4298);
nor U5519 (N_5519,N_3827,N_3437);
and U5520 (N_5520,N_4355,N_3104);
nand U5521 (N_5521,N_3312,N_4133);
and U5522 (N_5522,N_3799,N_4235);
or U5523 (N_5523,N_3754,N_3187);
or U5524 (N_5524,N_3211,N_3530);
and U5525 (N_5525,N_3332,N_3408);
or U5526 (N_5526,N_3189,N_3844);
or U5527 (N_5527,N_4149,N_3006);
xnor U5528 (N_5528,N_3882,N_3717);
nand U5529 (N_5529,N_4368,N_3557);
and U5530 (N_5530,N_4431,N_3984);
and U5531 (N_5531,N_3136,N_3748);
and U5532 (N_5532,N_4308,N_3653);
nor U5533 (N_5533,N_3110,N_3738);
nand U5534 (N_5534,N_4316,N_3999);
or U5535 (N_5535,N_3333,N_3714);
xor U5536 (N_5536,N_3920,N_3753);
or U5537 (N_5537,N_4354,N_3977);
nor U5538 (N_5538,N_3918,N_3274);
and U5539 (N_5539,N_3895,N_3360);
nor U5540 (N_5540,N_4227,N_3372);
nor U5541 (N_5541,N_4212,N_3673);
or U5542 (N_5542,N_3328,N_3938);
xnor U5543 (N_5543,N_3118,N_4464);
nor U5544 (N_5544,N_3664,N_4431);
nand U5545 (N_5545,N_3203,N_3980);
or U5546 (N_5546,N_3532,N_4371);
nand U5547 (N_5547,N_4199,N_4418);
nand U5548 (N_5548,N_4399,N_3626);
and U5549 (N_5549,N_3559,N_3793);
or U5550 (N_5550,N_3636,N_4146);
nor U5551 (N_5551,N_4324,N_4235);
and U5552 (N_5552,N_3669,N_3150);
nor U5553 (N_5553,N_4375,N_3927);
nand U5554 (N_5554,N_3631,N_4246);
and U5555 (N_5555,N_3027,N_3363);
or U5556 (N_5556,N_3651,N_3975);
and U5557 (N_5557,N_3983,N_3179);
and U5558 (N_5558,N_3374,N_4418);
nor U5559 (N_5559,N_3623,N_3597);
nor U5560 (N_5560,N_3646,N_3635);
and U5561 (N_5561,N_3773,N_3385);
xnor U5562 (N_5562,N_3487,N_3874);
or U5563 (N_5563,N_3491,N_3152);
nor U5564 (N_5564,N_3913,N_4214);
nor U5565 (N_5565,N_4395,N_4225);
nor U5566 (N_5566,N_3493,N_3155);
and U5567 (N_5567,N_3914,N_4313);
nor U5568 (N_5568,N_4223,N_3887);
nand U5569 (N_5569,N_3852,N_4071);
nor U5570 (N_5570,N_3782,N_4483);
nor U5571 (N_5571,N_3993,N_3341);
xnor U5572 (N_5572,N_3993,N_3215);
or U5573 (N_5573,N_3695,N_4302);
and U5574 (N_5574,N_3227,N_3488);
and U5575 (N_5575,N_3970,N_3018);
nor U5576 (N_5576,N_4475,N_3795);
nand U5577 (N_5577,N_3218,N_4189);
nand U5578 (N_5578,N_4351,N_4173);
xor U5579 (N_5579,N_4101,N_3859);
nand U5580 (N_5580,N_4482,N_3741);
nor U5581 (N_5581,N_3576,N_3453);
nand U5582 (N_5582,N_3733,N_3862);
nor U5583 (N_5583,N_4441,N_4271);
nor U5584 (N_5584,N_3856,N_4201);
xor U5585 (N_5585,N_4131,N_3436);
nand U5586 (N_5586,N_4288,N_3227);
or U5587 (N_5587,N_3350,N_3081);
and U5588 (N_5588,N_4024,N_3406);
or U5589 (N_5589,N_3340,N_4218);
and U5590 (N_5590,N_3537,N_4487);
or U5591 (N_5591,N_4463,N_3713);
or U5592 (N_5592,N_3403,N_4300);
or U5593 (N_5593,N_3066,N_3184);
nor U5594 (N_5594,N_4172,N_3620);
nand U5595 (N_5595,N_4474,N_3323);
or U5596 (N_5596,N_3705,N_4081);
and U5597 (N_5597,N_3428,N_3989);
xnor U5598 (N_5598,N_3427,N_3351);
nor U5599 (N_5599,N_3962,N_3595);
nor U5600 (N_5600,N_3155,N_3637);
or U5601 (N_5601,N_3123,N_4161);
xor U5602 (N_5602,N_3774,N_3789);
or U5603 (N_5603,N_3011,N_3486);
and U5604 (N_5604,N_3180,N_3107);
or U5605 (N_5605,N_4180,N_4259);
nor U5606 (N_5606,N_3471,N_3707);
or U5607 (N_5607,N_3171,N_4109);
and U5608 (N_5608,N_3520,N_3038);
and U5609 (N_5609,N_3912,N_4335);
and U5610 (N_5610,N_3071,N_3712);
xnor U5611 (N_5611,N_3092,N_3208);
nor U5612 (N_5612,N_4316,N_3595);
xnor U5613 (N_5613,N_4477,N_4451);
nand U5614 (N_5614,N_3582,N_3652);
xor U5615 (N_5615,N_4008,N_4296);
nor U5616 (N_5616,N_3713,N_3179);
nor U5617 (N_5617,N_4061,N_3689);
and U5618 (N_5618,N_3939,N_4471);
nor U5619 (N_5619,N_3342,N_3315);
nor U5620 (N_5620,N_3871,N_4171);
nand U5621 (N_5621,N_3605,N_4267);
xor U5622 (N_5622,N_3167,N_3003);
nand U5623 (N_5623,N_3105,N_3007);
nor U5624 (N_5624,N_3043,N_3655);
xor U5625 (N_5625,N_3083,N_4412);
or U5626 (N_5626,N_4008,N_3634);
and U5627 (N_5627,N_3949,N_3463);
or U5628 (N_5628,N_4022,N_3824);
and U5629 (N_5629,N_3485,N_4316);
or U5630 (N_5630,N_3889,N_3045);
and U5631 (N_5631,N_3856,N_3099);
nand U5632 (N_5632,N_4459,N_3176);
nor U5633 (N_5633,N_4350,N_3650);
nor U5634 (N_5634,N_3385,N_4460);
and U5635 (N_5635,N_3279,N_3552);
xnor U5636 (N_5636,N_3249,N_4131);
nor U5637 (N_5637,N_3135,N_3490);
and U5638 (N_5638,N_3726,N_3042);
and U5639 (N_5639,N_3637,N_3921);
and U5640 (N_5640,N_3404,N_3640);
or U5641 (N_5641,N_3521,N_3098);
nand U5642 (N_5642,N_3295,N_4035);
or U5643 (N_5643,N_3227,N_3932);
or U5644 (N_5644,N_3094,N_3411);
nor U5645 (N_5645,N_3007,N_3051);
nand U5646 (N_5646,N_4197,N_4486);
nor U5647 (N_5647,N_4487,N_4319);
nor U5648 (N_5648,N_4462,N_3062);
and U5649 (N_5649,N_3367,N_3100);
and U5650 (N_5650,N_4213,N_3459);
and U5651 (N_5651,N_3602,N_3560);
xor U5652 (N_5652,N_4391,N_4455);
or U5653 (N_5653,N_3070,N_3531);
or U5654 (N_5654,N_4295,N_4046);
nor U5655 (N_5655,N_3229,N_4121);
xor U5656 (N_5656,N_4430,N_3899);
nand U5657 (N_5657,N_3279,N_4003);
or U5658 (N_5658,N_4070,N_4169);
nand U5659 (N_5659,N_3510,N_3866);
nand U5660 (N_5660,N_3072,N_3369);
nand U5661 (N_5661,N_3543,N_3798);
and U5662 (N_5662,N_3311,N_4076);
or U5663 (N_5663,N_4253,N_3094);
nor U5664 (N_5664,N_4093,N_3026);
nor U5665 (N_5665,N_3619,N_4438);
xnor U5666 (N_5666,N_3794,N_3011);
or U5667 (N_5667,N_4126,N_3649);
and U5668 (N_5668,N_3653,N_4066);
nand U5669 (N_5669,N_4499,N_4183);
nand U5670 (N_5670,N_3011,N_3968);
nand U5671 (N_5671,N_3169,N_3811);
and U5672 (N_5672,N_3487,N_4145);
nand U5673 (N_5673,N_3206,N_3495);
nand U5674 (N_5674,N_3024,N_3410);
or U5675 (N_5675,N_3008,N_4163);
nor U5676 (N_5676,N_3691,N_3157);
and U5677 (N_5677,N_3863,N_3651);
nor U5678 (N_5678,N_4085,N_3875);
or U5679 (N_5679,N_3474,N_3840);
nor U5680 (N_5680,N_3375,N_4445);
nor U5681 (N_5681,N_3295,N_3149);
and U5682 (N_5682,N_4278,N_3862);
or U5683 (N_5683,N_3831,N_4332);
or U5684 (N_5684,N_4362,N_3887);
nand U5685 (N_5685,N_3505,N_3716);
and U5686 (N_5686,N_3028,N_3595);
nand U5687 (N_5687,N_3114,N_3189);
and U5688 (N_5688,N_4183,N_4280);
xnor U5689 (N_5689,N_3790,N_4408);
nand U5690 (N_5690,N_4478,N_3580);
nor U5691 (N_5691,N_4328,N_3889);
nor U5692 (N_5692,N_4267,N_3697);
or U5693 (N_5693,N_3987,N_3789);
nand U5694 (N_5694,N_4190,N_4006);
nor U5695 (N_5695,N_4288,N_3617);
and U5696 (N_5696,N_3802,N_3925);
and U5697 (N_5697,N_3260,N_3588);
nor U5698 (N_5698,N_4432,N_4061);
xor U5699 (N_5699,N_3473,N_3726);
or U5700 (N_5700,N_3240,N_4122);
nand U5701 (N_5701,N_3596,N_3180);
and U5702 (N_5702,N_3678,N_3369);
and U5703 (N_5703,N_3871,N_3307);
nand U5704 (N_5704,N_3015,N_3299);
nand U5705 (N_5705,N_3516,N_3692);
or U5706 (N_5706,N_3638,N_3961);
nor U5707 (N_5707,N_3867,N_3531);
nor U5708 (N_5708,N_3789,N_4280);
nor U5709 (N_5709,N_3311,N_3777);
xnor U5710 (N_5710,N_4257,N_3347);
nand U5711 (N_5711,N_3738,N_3126);
nand U5712 (N_5712,N_4374,N_4315);
nand U5713 (N_5713,N_3639,N_4132);
nand U5714 (N_5714,N_3430,N_3195);
or U5715 (N_5715,N_3064,N_4241);
and U5716 (N_5716,N_3823,N_4305);
xor U5717 (N_5717,N_3861,N_3510);
nand U5718 (N_5718,N_4150,N_3322);
nand U5719 (N_5719,N_3781,N_3438);
or U5720 (N_5720,N_4327,N_3199);
nor U5721 (N_5721,N_3891,N_4066);
nand U5722 (N_5722,N_3108,N_4119);
or U5723 (N_5723,N_4470,N_3223);
xnor U5724 (N_5724,N_4484,N_4322);
nand U5725 (N_5725,N_4405,N_4152);
nor U5726 (N_5726,N_3897,N_4242);
and U5727 (N_5727,N_4028,N_3092);
or U5728 (N_5728,N_4391,N_4223);
and U5729 (N_5729,N_3208,N_3413);
xor U5730 (N_5730,N_3271,N_3753);
nand U5731 (N_5731,N_3327,N_4260);
nand U5732 (N_5732,N_3218,N_3143);
nand U5733 (N_5733,N_3700,N_4101);
xor U5734 (N_5734,N_4359,N_4258);
xor U5735 (N_5735,N_4288,N_4495);
and U5736 (N_5736,N_4472,N_3920);
or U5737 (N_5737,N_3226,N_3356);
nand U5738 (N_5738,N_3258,N_3139);
nor U5739 (N_5739,N_4473,N_3431);
xnor U5740 (N_5740,N_3171,N_3756);
nor U5741 (N_5741,N_4354,N_3596);
or U5742 (N_5742,N_3799,N_3507);
nor U5743 (N_5743,N_3442,N_3449);
nand U5744 (N_5744,N_3182,N_3103);
nor U5745 (N_5745,N_3576,N_3944);
nand U5746 (N_5746,N_3827,N_3139);
nand U5747 (N_5747,N_3031,N_3030);
nor U5748 (N_5748,N_3092,N_4150);
and U5749 (N_5749,N_4293,N_3130);
and U5750 (N_5750,N_4497,N_4451);
and U5751 (N_5751,N_3261,N_3316);
and U5752 (N_5752,N_4255,N_3903);
and U5753 (N_5753,N_4461,N_3353);
nor U5754 (N_5754,N_3970,N_3102);
and U5755 (N_5755,N_4013,N_3811);
nand U5756 (N_5756,N_3221,N_3644);
and U5757 (N_5757,N_3526,N_3655);
nand U5758 (N_5758,N_3476,N_3129);
or U5759 (N_5759,N_3726,N_3203);
or U5760 (N_5760,N_3358,N_3052);
nor U5761 (N_5761,N_4462,N_4329);
nand U5762 (N_5762,N_3917,N_3836);
nor U5763 (N_5763,N_3452,N_4198);
nor U5764 (N_5764,N_4033,N_4497);
or U5765 (N_5765,N_3903,N_3770);
and U5766 (N_5766,N_4154,N_3448);
nand U5767 (N_5767,N_4460,N_3669);
nand U5768 (N_5768,N_4077,N_4120);
nand U5769 (N_5769,N_3090,N_4348);
nor U5770 (N_5770,N_3328,N_3307);
and U5771 (N_5771,N_4302,N_4300);
nand U5772 (N_5772,N_4370,N_3697);
and U5773 (N_5773,N_3099,N_3287);
nor U5774 (N_5774,N_3055,N_3875);
or U5775 (N_5775,N_3976,N_4253);
nand U5776 (N_5776,N_3186,N_3755);
or U5777 (N_5777,N_3115,N_3783);
or U5778 (N_5778,N_3446,N_4026);
nor U5779 (N_5779,N_3005,N_3368);
or U5780 (N_5780,N_3075,N_3055);
or U5781 (N_5781,N_3985,N_4204);
or U5782 (N_5782,N_3508,N_3223);
or U5783 (N_5783,N_3271,N_3385);
or U5784 (N_5784,N_4471,N_4026);
xnor U5785 (N_5785,N_3603,N_4108);
and U5786 (N_5786,N_4454,N_4206);
nand U5787 (N_5787,N_3488,N_3532);
nor U5788 (N_5788,N_4487,N_3592);
nor U5789 (N_5789,N_4293,N_4035);
and U5790 (N_5790,N_4238,N_3610);
or U5791 (N_5791,N_3698,N_3986);
xor U5792 (N_5792,N_3859,N_3237);
nor U5793 (N_5793,N_3923,N_3672);
xnor U5794 (N_5794,N_4447,N_3453);
or U5795 (N_5795,N_3996,N_3864);
or U5796 (N_5796,N_3508,N_3997);
xnor U5797 (N_5797,N_3011,N_3316);
or U5798 (N_5798,N_4055,N_4376);
nor U5799 (N_5799,N_3684,N_3889);
nand U5800 (N_5800,N_4455,N_3248);
and U5801 (N_5801,N_4275,N_3910);
and U5802 (N_5802,N_3693,N_3921);
nor U5803 (N_5803,N_3517,N_4360);
or U5804 (N_5804,N_4324,N_3202);
and U5805 (N_5805,N_3466,N_3413);
or U5806 (N_5806,N_3487,N_3673);
and U5807 (N_5807,N_3809,N_4275);
nor U5808 (N_5808,N_3952,N_3074);
nor U5809 (N_5809,N_3224,N_3588);
nor U5810 (N_5810,N_4008,N_3718);
nor U5811 (N_5811,N_3551,N_3028);
nor U5812 (N_5812,N_3681,N_3061);
and U5813 (N_5813,N_4075,N_4346);
nand U5814 (N_5814,N_3201,N_3415);
xnor U5815 (N_5815,N_4468,N_3367);
nor U5816 (N_5816,N_3438,N_3140);
xor U5817 (N_5817,N_4136,N_3214);
and U5818 (N_5818,N_4156,N_4065);
and U5819 (N_5819,N_3918,N_3534);
nand U5820 (N_5820,N_3812,N_3481);
and U5821 (N_5821,N_3249,N_3092);
xnor U5822 (N_5822,N_3296,N_4498);
nand U5823 (N_5823,N_3766,N_4080);
nand U5824 (N_5824,N_3420,N_4341);
nand U5825 (N_5825,N_4040,N_3071);
and U5826 (N_5826,N_4317,N_3333);
or U5827 (N_5827,N_4446,N_3190);
nand U5828 (N_5828,N_3184,N_3140);
nor U5829 (N_5829,N_4228,N_4036);
and U5830 (N_5830,N_3148,N_3616);
nand U5831 (N_5831,N_4118,N_3393);
nor U5832 (N_5832,N_3547,N_3005);
and U5833 (N_5833,N_3777,N_4036);
nor U5834 (N_5834,N_4236,N_4274);
or U5835 (N_5835,N_4015,N_4296);
or U5836 (N_5836,N_4254,N_3060);
nor U5837 (N_5837,N_3290,N_3780);
and U5838 (N_5838,N_4328,N_3209);
or U5839 (N_5839,N_4428,N_3024);
and U5840 (N_5840,N_3880,N_4092);
nor U5841 (N_5841,N_3069,N_4254);
xor U5842 (N_5842,N_3179,N_3032);
nand U5843 (N_5843,N_4104,N_3931);
or U5844 (N_5844,N_3284,N_3400);
nor U5845 (N_5845,N_4240,N_3157);
nor U5846 (N_5846,N_4272,N_3518);
nor U5847 (N_5847,N_3871,N_3888);
xor U5848 (N_5848,N_4357,N_3574);
and U5849 (N_5849,N_3739,N_3008);
nor U5850 (N_5850,N_4097,N_3642);
and U5851 (N_5851,N_3547,N_3227);
and U5852 (N_5852,N_3397,N_3894);
or U5853 (N_5853,N_3097,N_3916);
xnor U5854 (N_5854,N_3111,N_3781);
and U5855 (N_5855,N_3006,N_4005);
nand U5856 (N_5856,N_4241,N_4080);
or U5857 (N_5857,N_4405,N_3744);
or U5858 (N_5858,N_3775,N_3611);
nand U5859 (N_5859,N_4273,N_3626);
and U5860 (N_5860,N_3983,N_4459);
nand U5861 (N_5861,N_3316,N_4084);
nand U5862 (N_5862,N_3412,N_4128);
and U5863 (N_5863,N_3269,N_3270);
nor U5864 (N_5864,N_3269,N_4342);
and U5865 (N_5865,N_3781,N_4405);
nor U5866 (N_5866,N_3010,N_4000);
nor U5867 (N_5867,N_3181,N_3758);
nor U5868 (N_5868,N_3627,N_3357);
xor U5869 (N_5869,N_3858,N_3673);
nor U5870 (N_5870,N_3699,N_3184);
or U5871 (N_5871,N_4100,N_3002);
or U5872 (N_5872,N_3289,N_3100);
and U5873 (N_5873,N_3909,N_3802);
or U5874 (N_5874,N_3286,N_3324);
nor U5875 (N_5875,N_4045,N_3633);
and U5876 (N_5876,N_4189,N_3178);
nor U5877 (N_5877,N_3014,N_3423);
nor U5878 (N_5878,N_4223,N_3607);
nand U5879 (N_5879,N_3180,N_4038);
nor U5880 (N_5880,N_3876,N_4083);
nand U5881 (N_5881,N_4376,N_4495);
or U5882 (N_5882,N_4466,N_3331);
or U5883 (N_5883,N_4458,N_3552);
xnor U5884 (N_5884,N_3106,N_3338);
nor U5885 (N_5885,N_3678,N_4366);
nor U5886 (N_5886,N_4440,N_4142);
and U5887 (N_5887,N_4469,N_3771);
nor U5888 (N_5888,N_3455,N_4041);
nor U5889 (N_5889,N_3631,N_3488);
xnor U5890 (N_5890,N_4206,N_4056);
xnor U5891 (N_5891,N_3511,N_3101);
nand U5892 (N_5892,N_4426,N_4004);
or U5893 (N_5893,N_4155,N_4058);
xnor U5894 (N_5894,N_3703,N_3412);
or U5895 (N_5895,N_4028,N_3059);
or U5896 (N_5896,N_3067,N_3900);
xor U5897 (N_5897,N_3238,N_3764);
and U5898 (N_5898,N_3641,N_4350);
or U5899 (N_5899,N_3500,N_3056);
and U5900 (N_5900,N_3220,N_4042);
or U5901 (N_5901,N_4228,N_4048);
or U5902 (N_5902,N_4477,N_3152);
nand U5903 (N_5903,N_3544,N_4442);
or U5904 (N_5904,N_3861,N_4254);
nand U5905 (N_5905,N_3311,N_3830);
and U5906 (N_5906,N_4497,N_3410);
nor U5907 (N_5907,N_3862,N_4095);
or U5908 (N_5908,N_3711,N_4316);
or U5909 (N_5909,N_3780,N_3800);
xor U5910 (N_5910,N_4398,N_4173);
nand U5911 (N_5911,N_4277,N_3737);
or U5912 (N_5912,N_3246,N_3593);
and U5913 (N_5913,N_4029,N_3985);
nand U5914 (N_5914,N_4269,N_3257);
or U5915 (N_5915,N_3316,N_3989);
nor U5916 (N_5916,N_4423,N_3505);
nand U5917 (N_5917,N_3308,N_3111);
nand U5918 (N_5918,N_3354,N_3704);
xnor U5919 (N_5919,N_3401,N_4055);
xor U5920 (N_5920,N_4388,N_3461);
and U5921 (N_5921,N_4105,N_3961);
nand U5922 (N_5922,N_3390,N_3144);
or U5923 (N_5923,N_4280,N_4437);
and U5924 (N_5924,N_4306,N_4496);
nor U5925 (N_5925,N_4215,N_4104);
and U5926 (N_5926,N_4042,N_4413);
nand U5927 (N_5927,N_3703,N_3804);
nor U5928 (N_5928,N_3679,N_3933);
nor U5929 (N_5929,N_3491,N_3448);
nor U5930 (N_5930,N_3389,N_3398);
or U5931 (N_5931,N_3976,N_3031);
and U5932 (N_5932,N_4432,N_3534);
or U5933 (N_5933,N_3837,N_4199);
and U5934 (N_5934,N_3826,N_4248);
and U5935 (N_5935,N_4381,N_3364);
nand U5936 (N_5936,N_3962,N_3665);
and U5937 (N_5937,N_3523,N_4252);
or U5938 (N_5938,N_4304,N_3662);
nand U5939 (N_5939,N_3060,N_3828);
and U5940 (N_5940,N_3379,N_3054);
nand U5941 (N_5941,N_4343,N_3220);
nand U5942 (N_5942,N_4295,N_4268);
or U5943 (N_5943,N_3401,N_3272);
xnor U5944 (N_5944,N_3633,N_3561);
or U5945 (N_5945,N_3219,N_4095);
and U5946 (N_5946,N_3357,N_3610);
and U5947 (N_5947,N_4148,N_4007);
nand U5948 (N_5948,N_3256,N_4090);
and U5949 (N_5949,N_3328,N_4000);
or U5950 (N_5950,N_4112,N_3436);
nor U5951 (N_5951,N_4179,N_4454);
or U5952 (N_5952,N_3307,N_3832);
nor U5953 (N_5953,N_3894,N_4342);
and U5954 (N_5954,N_4293,N_3828);
or U5955 (N_5955,N_4059,N_4091);
xor U5956 (N_5956,N_3669,N_4326);
nand U5957 (N_5957,N_3112,N_4280);
xnor U5958 (N_5958,N_4358,N_4258);
xor U5959 (N_5959,N_3881,N_3893);
nor U5960 (N_5960,N_3644,N_3388);
and U5961 (N_5961,N_4104,N_3508);
nand U5962 (N_5962,N_3440,N_4348);
nor U5963 (N_5963,N_4055,N_3816);
or U5964 (N_5964,N_4076,N_3772);
xnor U5965 (N_5965,N_3372,N_3053);
or U5966 (N_5966,N_3122,N_3424);
or U5967 (N_5967,N_4283,N_3840);
nand U5968 (N_5968,N_3522,N_4410);
nor U5969 (N_5969,N_3785,N_4037);
nor U5970 (N_5970,N_3925,N_4359);
or U5971 (N_5971,N_3460,N_3250);
nor U5972 (N_5972,N_3013,N_4115);
xor U5973 (N_5973,N_3519,N_4312);
nand U5974 (N_5974,N_3373,N_3976);
xor U5975 (N_5975,N_3865,N_3888);
xor U5976 (N_5976,N_3465,N_3244);
and U5977 (N_5977,N_3766,N_4451);
and U5978 (N_5978,N_3587,N_3775);
or U5979 (N_5979,N_3722,N_3851);
xnor U5980 (N_5980,N_3230,N_4155);
and U5981 (N_5981,N_4353,N_4232);
and U5982 (N_5982,N_3951,N_3480);
nand U5983 (N_5983,N_3923,N_4497);
or U5984 (N_5984,N_3989,N_3462);
or U5985 (N_5985,N_3740,N_3237);
nand U5986 (N_5986,N_4187,N_3703);
xor U5987 (N_5987,N_4294,N_3605);
and U5988 (N_5988,N_3682,N_3905);
and U5989 (N_5989,N_4000,N_3593);
nor U5990 (N_5990,N_4188,N_3847);
nor U5991 (N_5991,N_4480,N_4044);
nand U5992 (N_5992,N_4121,N_3672);
and U5993 (N_5993,N_3101,N_3879);
and U5994 (N_5994,N_4070,N_4067);
and U5995 (N_5995,N_4449,N_3156);
nand U5996 (N_5996,N_3023,N_4426);
nand U5997 (N_5997,N_3539,N_3691);
nand U5998 (N_5998,N_4057,N_4285);
xnor U5999 (N_5999,N_4044,N_4051);
or U6000 (N_6000,N_5271,N_5555);
xor U6001 (N_6001,N_5575,N_5835);
or U6002 (N_6002,N_4983,N_5206);
nand U6003 (N_6003,N_5549,N_4929);
and U6004 (N_6004,N_5726,N_5881);
or U6005 (N_6005,N_5043,N_5189);
nor U6006 (N_6006,N_5802,N_5940);
xnor U6007 (N_6007,N_5755,N_5606);
nor U6008 (N_6008,N_5197,N_5527);
nor U6009 (N_6009,N_5548,N_5706);
nor U6010 (N_6010,N_4877,N_5348);
and U6011 (N_6011,N_5041,N_5459);
or U6012 (N_6012,N_4910,N_5897);
and U6013 (N_6013,N_5398,N_5418);
xor U6014 (N_6014,N_5986,N_4536);
and U6015 (N_6015,N_5462,N_4559);
nand U6016 (N_6016,N_5784,N_5499);
nand U6017 (N_6017,N_5878,N_5998);
and U6018 (N_6018,N_4567,N_5336);
or U6019 (N_6019,N_4750,N_5050);
or U6020 (N_6020,N_5617,N_4915);
and U6021 (N_6021,N_4964,N_4534);
nand U6022 (N_6022,N_5656,N_4936);
nand U6023 (N_6023,N_4800,N_5852);
nand U6024 (N_6024,N_5437,N_5036);
or U6025 (N_6025,N_5038,N_5746);
nor U6026 (N_6026,N_5853,N_5566);
or U6027 (N_6027,N_5821,N_5521);
xnor U6028 (N_6028,N_5754,N_4587);
nor U6029 (N_6029,N_5449,N_5004);
nor U6030 (N_6030,N_4789,N_4869);
and U6031 (N_6031,N_5049,N_5352);
xor U6032 (N_6032,N_5309,N_5299);
or U6033 (N_6033,N_4514,N_4957);
nor U6034 (N_6034,N_4631,N_5236);
and U6035 (N_6035,N_4668,N_5910);
nand U6036 (N_6036,N_5035,N_5778);
or U6037 (N_6037,N_5861,N_4844);
and U6038 (N_6038,N_5423,N_4732);
nor U6039 (N_6039,N_5296,N_5481);
nand U6040 (N_6040,N_5615,N_5364);
nor U6041 (N_6041,N_4933,N_5490);
and U6042 (N_6042,N_4935,N_4865);
nor U6043 (N_6043,N_5612,N_4535);
nand U6044 (N_6044,N_5845,N_5228);
nand U6045 (N_6045,N_4526,N_5938);
nor U6046 (N_6046,N_4589,N_5900);
nor U6047 (N_6047,N_5609,N_5401);
or U6048 (N_6048,N_5948,N_5472);
nor U6049 (N_6049,N_5922,N_4878);
nor U6050 (N_6050,N_5077,N_5984);
nand U6051 (N_6051,N_5086,N_5993);
xnor U6052 (N_6052,N_5536,N_4576);
xor U6053 (N_6053,N_5582,N_4947);
and U6054 (N_6054,N_4902,N_5719);
nor U6055 (N_6055,N_4613,N_4709);
or U6056 (N_6056,N_5457,N_4760);
nor U6057 (N_6057,N_4773,N_4999);
nand U6058 (N_6058,N_5955,N_5093);
or U6059 (N_6059,N_4508,N_4585);
and U6060 (N_6060,N_4724,N_5742);
nor U6061 (N_6061,N_4956,N_4806);
or U6062 (N_6062,N_5202,N_4655);
nand U6063 (N_6063,N_5648,N_5087);
and U6064 (N_6064,N_4903,N_4620);
xnor U6065 (N_6065,N_5862,N_4510);
nand U6066 (N_6066,N_4867,N_4977);
or U6067 (N_6067,N_5048,N_5316);
nand U6068 (N_6068,N_4688,N_5338);
nor U6069 (N_6069,N_4890,N_5892);
or U6070 (N_6070,N_5935,N_5427);
nor U6071 (N_6071,N_5539,N_5693);
or U6072 (N_6072,N_5397,N_5244);
or U6073 (N_6073,N_5126,N_5903);
or U6074 (N_6074,N_5468,N_5221);
nor U6075 (N_6075,N_5239,N_5107);
or U6076 (N_6076,N_5252,N_5996);
nand U6077 (N_6077,N_5321,N_4808);
or U6078 (N_6078,N_4636,N_5332);
nor U6079 (N_6079,N_5240,N_4539);
and U6080 (N_6080,N_5194,N_5592);
nand U6081 (N_6081,N_5127,N_5392);
or U6082 (N_6082,N_4893,N_5629);
and U6083 (N_6083,N_4676,N_5760);
and U6084 (N_6084,N_5085,N_5602);
xnor U6085 (N_6085,N_5226,N_5762);
or U6086 (N_6086,N_4687,N_5285);
xnor U6087 (N_6087,N_5017,N_5353);
or U6088 (N_6088,N_4812,N_4594);
or U6089 (N_6089,N_5911,N_4777);
nand U6090 (N_6090,N_5010,N_5820);
nor U6091 (N_6091,N_5400,N_4522);
nand U6092 (N_6092,N_5979,N_4985);
nand U6093 (N_6093,N_4914,N_4794);
nor U6094 (N_6094,N_5789,N_5689);
or U6095 (N_6095,N_5956,N_4928);
and U6096 (N_6096,N_4811,N_4911);
and U6097 (N_6097,N_4930,N_5920);
and U6098 (N_6098,N_4775,N_5524);
nor U6099 (N_6099,N_5435,N_5088);
and U6100 (N_6100,N_5764,N_4931);
and U6101 (N_6101,N_4504,N_4669);
nand U6102 (N_6102,N_5070,N_4849);
or U6103 (N_6103,N_5937,N_5745);
and U6104 (N_6104,N_4634,N_5385);
and U6105 (N_6105,N_5003,N_4718);
and U6106 (N_6106,N_5395,N_4719);
nand U6107 (N_6107,N_4897,N_5894);
and U6108 (N_6108,N_5672,N_5219);
or U6109 (N_6109,N_5734,N_5058);
nor U6110 (N_6110,N_5696,N_5276);
nand U6111 (N_6111,N_5443,N_5618);
or U6112 (N_6112,N_5171,N_5924);
nor U6113 (N_6113,N_4916,N_5214);
nand U6114 (N_6114,N_5112,N_5224);
nand U6115 (N_6115,N_5512,N_5941);
nand U6116 (N_6116,N_5474,N_5812);
or U6117 (N_6117,N_5770,N_5039);
nor U6118 (N_6118,N_4828,N_5717);
nor U6119 (N_6119,N_5517,N_5664);
nor U6120 (N_6120,N_5703,N_5119);
nand U6121 (N_6121,N_4846,N_5500);
nand U6122 (N_6122,N_4638,N_4656);
or U6123 (N_6123,N_4778,N_5857);
and U6124 (N_6124,N_4689,N_5008);
nor U6125 (N_6125,N_5094,N_5558);
nand U6126 (N_6126,N_5439,N_5560);
nor U6127 (N_6127,N_5268,N_4934);
and U6128 (N_6128,N_5936,N_4619);
and U6129 (N_6129,N_4745,N_5367);
nor U6130 (N_6130,N_5836,N_5595);
nand U6131 (N_6131,N_4954,N_4521);
and U6132 (N_6132,N_5947,N_5181);
and U6133 (N_6133,N_5139,N_5415);
nor U6134 (N_6134,N_5626,N_4974);
xor U6135 (N_6135,N_5078,N_5972);
and U6136 (N_6136,N_4949,N_4894);
nand U6137 (N_6137,N_5889,N_5037);
xnor U6138 (N_6138,N_5767,N_4793);
and U6139 (N_6139,N_5799,N_5954);
or U6140 (N_6140,N_5263,N_4734);
nand U6141 (N_6141,N_4994,N_5649);
and U6142 (N_6142,N_5636,N_5893);
and U6143 (N_6143,N_5318,N_4829);
xnor U6144 (N_6144,N_5756,N_4838);
nand U6145 (N_6145,N_4986,N_4660);
nor U6146 (N_6146,N_5982,N_5045);
nor U6147 (N_6147,N_5934,N_5383);
or U6148 (N_6148,N_5773,N_4998);
nor U6149 (N_6149,N_4976,N_5442);
nor U6150 (N_6150,N_5682,N_5844);
nand U6151 (N_6151,N_5670,N_5559);
or U6152 (N_6152,N_4888,N_5735);
nand U6153 (N_6153,N_4663,N_5033);
and U6154 (N_6154,N_5780,N_5776);
and U6155 (N_6155,N_5229,N_5959);
and U6156 (N_6156,N_4607,N_5528);
nor U6157 (N_6157,N_5628,N_4713);
and U6158 (N_6158,N_4992,N_4770);
and U6159 (N_6159,N_5644,N_5065);
and U6160 (N_6160,N_5794,N_4917);
nand U6161 (N_6161,N_5104,N_4978);
nand U6162 (N_6162,N_4755,N_5025);
nor U6163 (N_6163,N_5200,N_5804);
and U6164 (N_6164,N_5064,N_5319);
nand U6165 (N_6165,N_5515,N_5402);
nor U6166 (N_6166,N_5391,N_4802);
xor U6167 (N_6167,N_5300,N_4747);
nand U6168 (N_6168,N_4905,N_5495);
or U6169 (N_6169,N_5619,N_5850);
nor U6170 (N_6170,N_5024,N_4795);
nor U6171 (N_6171,N_4749,N_5710);
nand U6172 (N_6172,N_4600,N_4881);
nor U6173 (N_6173,N_5198,N_5180);
or U6174 (N_6174,N_4898,N_5151);
nor U6175 (N_6175,N_4762,N_5311);
nand U6176 (N_6176,N_4809,N_5394);
and U6177 (N_6177,N_4791,N_4783);
and U6178 (N_6178,N_5054,N_4548);
nor U6179 (N_6179,N_4590,N_4624);
nor U6180 (N_6180,N_5218,N_5326);
nor U6181 (N_6181,N_5568,N_5456);
and U6182 (N_6182,N_5080,N_4782);
or U6183 (N_6183,N_5469,N_5262);
nand U6184 (N_6184,N_5019,N_5284);
xor U6185 (N_6185,N_4561,N_5409);
or U6186 (N_6186,N_4603,N_5665);
nand U6187 (N_6187,N_5368,N_5733);
and U6188 (N_6188,N_5494,N_4675);
and U6189 (N_6189,N_5953,N_4907);
nand U6190 (N_6190,N_5950,N_5795);
or U6191 (N_6191,N_5021,N_4835);
and U6192 (N_6192,N_5393,N_5883);
and U6193 (N_6193,N_5526,N_4546);
xnor U6194 (N_6194,N_5382,N_5987);
nor U6195 (N_6195,N_5115,N_4651);
and U6196 (N_6196,N_4637,N_5165);
nor U6197 (N_6197,N_5123,N_5491);
or U6198 (N_6198,N_5546,N_5057);
nor U6199 (N_6199,N_5818,N_5623);
nor U6200 (N_6200,N_5583,N_4908);
or U6201 (N_6201,N_5062,N_4784);
and U6202 (N_6202,N_4695,N_5563);
and U6203 (N_6203,N_5854,N_5106);
nor U6204 (N_6204,N_4579,N_5514);
or U6205 (N_6205,N_5729,N_4737);
nor U6206 (N_6206,N_5809,N_4609);
xnor U6207 (N_6207,N_5662,N_5258);
xor U6208 (N_6208,N_5012,N_4913);
nor U6209 (N_6209,N_4761,N_5334);
and U6210 (N_6210,N_5621,N_5846);
nand U6211 (N_6211,N_4971,N_5961);
nand U6212 (N_6212,N_5807,N_5369);
nor U6213 (N_6213,N_5339,N_4602);
and U6214 (N_6214,N_5371,N_5275);
and U6215 (N_6215,N_5637,N_5158);
xnor U6216 (N_6216,N_5376,N_5387);
and U6217 (N_6217,N_5440,N_4923);
and U6218 (N_6218,N_4601,N_5341);
nor U6219 (N_6219,N_5425,N_5305);
or U6220 (N_6220,N_5925,N_4950);
and U6221 (N_6221,N_5463,N_4593);
and U6222 (N_6222,N_4804,N_5731);
or U6223 (N_6223,N_5650,N_5335);
nor U6224 (N_6224,N_5831,N_4925);
or U6225 (N_6225,N_5390,N_4840);
nand U6226 (N_6226,N_4618,N_5128);
and U6227 (N_6227,N_5969,N_5859);
and U6228 (N_6228,N_5408,N_4738);
and U6229 (N_6229,N_5906,N_5660);
or U6230 (N_6230,N_5134,N_5686);
nand U6231 (N_6231,N_5028,N_5960);
nand U6232 (N_6232,N_4818,N_4845);
xor U6233 (N_6233,N_4513,N_5215);
xnor U6234 (N_6234,N_5446,N_5014);
and U6235 (N_6235,N_5205,N_5243);
xnor U6236 (N_6236,N_4815,N_5225);
nor U6237 (N_6237,N_5089,N_5797);
nor U6238 (N_6238,N_4884,N_5470);
and U6239 (N_6239,N_5248,N_5709);
or U6240 (N_6240,N_5360,N_4509);
and U6241 (N_6241,N_5242,N_5148);
or U6242 (N_6242,N_5504,N_4952);
nor U6243 (N_6243,N_4735,N_4507);
nand U6244 (N_6244,N_4757,N_5105);
nand U6245 (N_6245,N_5355,N_4906);
and U6246 (N_6246,N_5365,N_5673);
xor U6247 (N_6247,N_5531,N_4501);
and U6248 (N_6248,N_5381,N_4988);
and U6249 (N_6249,N_5000,N_5994);
or U6250 (N_6250,N_4683,N_4754);
and U6251 (N_6251,N_4856,N_5523);
and U6252 (N_6252,N_5677,N_5075);
or U6253 (N_6253,N_5034,N_4940);
nor U6254 (N_6254,N_5654,N_4944);
nand U6255 (N_6255,N_4855,N_4831);
nand U6256 (N_6256,N_5209,N_5805);
nor U6257 (N_6257,N_5161,N_4643);
nand U6258 (N_6258,N_4705,N_4573);
nor U6259 (N_6259,N_5542,N_4505);
nand U6260 (N_6260,N_5287,N_5980);
nand U6261 (N_6261,N_4690,N_5183);
and U6262 (N_6262,N_4604,N_5479);
or U6263 (N_6263,N_5758,N_5416);
or U6264 (N_6264,N_5052,N_4671);
or U6265 (N_6265,N_4662,N_5018);
or U6266 (N_6266,N_4725,N_5538);
xor U6267 (N_6267,N_5858,N_5641);
or U6268 (N_6268,N_5154,N_5145);
or U6269 (N_6269,N_4805,N_5477);
nand U6270 (N_6270,N_5149,N_4771);
and U6271 (N_6271,N_5988,N_4623);
nor U6272 (N_6272,N_4550,N_4642);
xnor U6273 (N_6273,N_5051,N_5480);
or U6274 (N_6274,N_5507,N_4541);
or U6275 (N_6275,N_5781,N_5405);
or U6276 (N_6276,N_5557,N_5482);
or U6277 (N_6277,N_5567,N_5066);
nor U6278 (N_6278,N_5044,N_4730);
and U6279 (N_6279,N_4969,N_5995);
nand U6280 (N_6280,N_5485,N_5337);
nand U6281 (N_6281,N_5902,N_4617);
nor U6282 (N_6282,N_4584,N_5722);
nor U6283 (N_6283,N_4799,N_5997);
xor U6284 (N_6284,N_5532,N_5247);
and U6285 (N_6285,N_5848,N_4598);
and U6286 (N_6286,N_5574,N_4571);
xnor U6287 (N_6287,N_5964,N_5289);
nor U6288 (N_6288,N_4707,N_5785);
and U6289 (N_6289,N_4736,N_4785);
nor U6290 (N_6290,N_5331,N_5674);
or U6291 (N_6291,N_5260,N_5905);
nand U6292 (N_6292,N_5740,N_4648);
nand U6293 (N_6293,N_5346,N_4659);
nor U6294 (N_6294,N_4583,N_5417);
and U6295 (N_6295,N_5868,N_5071);
nor U6296 (N_6296,N_5493,N_4901);
or U6297 (N_6297,N_4622,N_5297);
nand U6298 (N_6298,N_4728,N_4722);
and U6299 (N_6299,N_5201,N_4666);
or U6300 (N_6300,N_5274,N_4502);
xor U6301 (N_6301,N_4699,N_5830);
nor U6302 (N_6302,N_4834,N_4551);
nand U6303 (N_6303,N_4547,N_4922);
nor U6304 (N_6304,N_4863,N_4970);
or U6305 (N_6305,N_4765,N_5235);
nor U6306 (N_6306,N_5187,N_4615);
and U6307 (N_6307,N_5779,N_5904);
nand U6308 (N_6308,N_5506,N_4560);
xnor U6309 (N_6309,N_5102,N_4552);
nor U6310 (N_6310,N_4595,N_5915);
nand U6311 (N_6311,N_4825,N_4955);
nor U6312 (N_6312,N_5736,N_5492);
nand U6313 (N_6313,N_5359,N_4640);
and U6314 (N_6314,N_5109,N_4591);
nor U6315 (N_6315,N_4821,N_4766);
and U6316 (N_6316,N_5810,N_5720);
or U6317 (N_6317,N_4946,N_5073);
nor U6318 (N_6318,N_5537,N_4715);
or U6319 (N_6319,N_5222,N_4817);
or U6320 (N_6320,N_5097,N_5651);
and U6321 (N_6321,N_5645,N_4562);
nand U6322 (N_6322,N_5403,N_5627);
nand U6323 (N_6323,N_5203,N_5261);
nand U6324 (N_6324,N_5256,N_5687);
nor U6325 (N_6325,N_5324,N_5315);
nand U6326 (N_6326,N_5631,N_5032);
or U6327 (N_6327,N_5678,N_4532);
and U6328 (N_6328,N_5738,N_5138);
and U6329 (N_6329,N_5535,N_5730);
and U6330 (N_6330,N_5728,N_5529);
or U6331 (N_6331,N_5386,N_4810);
nand U6332 (N_6332,N_5130,N_5047);
nor U6333 (N_6333,N_5281,N_5308);
nor U6334 (N_6334,N_5697,N_5949);
nand U6335 (N_6335,N_4774,N_5101);
nand U6336 (N_6336,N_5223,N_4506);
nor U6337 (N_6337,N_5272,N_5843);
nand U6338 (N_6338,N_4610,N_4706);
nand U6339 (N_6339,N_5976,N_5020);
xor U6340 (N_6340,N_4684,N_5570);
or U6341 (N_6341,N_5023,N_5632);
nor U6342 (N_6342,N_5565,N_5658);
nand U6343 (N_6343,N_5759,N_5452);
and U6344 (N_6344,N_5136,N_4565);
nand U6345 (N_6345,N_5152,N_5354);
and U6346 (N_6346,N_4652,N_5188);
xor U6347 (N_6347,N_5639,N_4698);
and U6348 (N_6348,N_5162,N_5292);
nor U6349 (N_6349,N_5562,N_5550);
nor U6350 (N_6350,N_5552,N_5067);
or U6351 (N_6351,N_5839,N_5554);
nor U6352 (N_6352,N_5884,N_4945);
or U6353 (N_6353,N_4837,N_5486);
nand U6354 (N_6354,N_5384,N_4939);
and U6355 (N_6355,N_4592,N_5692);
nand U6356 (N_6356,N_5450,N_4580);
and U6357 (N_6357,N_5667,N_4667);
or U6358 (N_6358,N_5144,N_5520);
and U6359 (N_6359,N_5766,N_5815);
or U6360 (N_6360,N_5471,N_5834);
and U6361 (N_6361,N_5793,N_5840);
or U6362 (N_6362,N_5569,N_5159);
and U6363 (N_6363,N_5646,N_5833);
nand U6364 (N_6364,N_5137,N_5864);
nand U6365 (N_6365,N_5573,N_5399);
or U6366 (N_6366,N_5842,N_5847);
nor U6367 (N_6367,N_5788,N_4861);
nand U6368 (N_6368,N_5156,N_5304);
or U6369 (N_6369,N_5505,N_5330);
and U6370 (N_6370,N_5195,N_4596);
and U6371 (N_6371,N_5026,N_4870);
or U6372 (N_6372,N_5313,N_5543);
or U6373 (N_6373,N_5002,N_5921);
xnor U6374 (N_6374,N_5973,N_5798);
nand U6375 (N_6375,N_4720,N_5173);
and U6376 (N_6376,N_4941,N_4892);
nor U6377 (N_6377,N_4826,N_5120);
nor U6378 (N_6378,N_5027,N_5340);
nand U6379 (N_6379,N_5741,N_4544);
nor U6380 (N_6380,N_5931,N_4721);
nor U6381 (N_6381,N_5928,N_5791);
or U6382 (N_6382,N_5761,N_5060);
or U6383 (N_6383,N_5061,N_4768);
and U6384 (N_6384,N_5556,N_5663);
and U6385 (N_6385,N_4696,N_4927);
xnor U6386 (N_6386,N_5613,N_5129);
nand U6387 (N_6387,N_4899,N_5282);
or U6388 (N_6388,N_5962,N_5497);
nand U6389 (N_6389,N_5977,N_4554);
nand U6390 (N_6390,N_5370,N_4980);
or U6391 (N_6391,N_5875,N_5255);
and U6392 (N_6392,N_4932,N_5022);
and U6393 (N_6393,N_5428,N_5978);
and U6394 (N_6394,N_5429,N_5966);
or U6395 (N_6395,N_5561,N_5607);
nand U6396 (N_6396,N_5763,N_5460);
nand U6397 (N_6397,N_4540,N_4758);
or U6398 (N_6398,N_5625,N_5204);
and U6399 (N_6399,N_4597,N_5942);
or U6400 (N_6400,N_4860,N_4751);
xor U6401 (N_6401,N_4752,N_5388);
nand U6402 (N_6402,N_5808,N_4919);
nor U6403 (N_6403,N_5882,N_5769);
xor U6404 (N_6404,N_5679,N_4876);
nand U6405 (N_6405,N_4852,N_4864);
and U6406 (N_6406,N_5916,N_4926);
nor U6407 (N_6407,N_5691,N_4886);
nor U6408 (N_6408,N_5633,N_4674);
and U6409 (N_6409,N_5185,N_5431);
or U6410 (N_6410,N_5851,N_5074);
nor U6411 (N_6411,N_5212,N_4883);
or U6412 (N_6412,N_4871,N_5142);
or U6413 (N_6413,N_4649,N_5251);
or U6414 (N_6414,N_5898,N_5208);
nand U6415 (N_6415,N_4909,N_5207);
and U6416 (N_6416,N_5886,N_5965);
or U6417 (N_6417,N_5293,N_5099);
or U6418 (N_6418,N_4836,N_4827);
nor U6419 (N_6419,N_4527,N_5362);
nand U6420 (N_6420,N_5153,N_5917);
and U6421 (N_6421,N_4608,N_5877);
nor U6422 (N_6422,N_4972,N_4630);
nand U6423 (N_6423,N_4851,N_4518);
xor U6424 (N_6424,N_4632,N_5519);
or U6425 (N_6425,N_4606,N_5466);
xor U6426 (N_6426,N_4966,N_5266);
nor U6427 (N_6427,N_4543,N_5705);
or U6428 (N_6428,N_5675,N_5981);
xor U6429 (N_6429,N_5991,N_5895);
xor U6430 (N_6430,N_4556,N_5118);
and U6431 (N_6431,N_5192,N_5455);
xor U6432 (N_6432,N_4672,N_5193);
nor U6433 (N_6433,N_5343,N_5880);
nor U6434 (N_6434,N_4965,N_5042);
nand U6435 (N_6435,N_5683,N_5600);
or U6436 (N_6436,N_5611,N_4664);
and U6437 (N_6437,N_4570,N_5744);
and U6438 (N_6438,N_4680,N_5908);
nor U6439 (N_6439,N_5551,N_4553);
xnor U6440 (N_6440,N_5501,N_5737);
or U6441 (N_6441,N_5347,N_5301);
xor U6442 (N_6442,N_5856,N_4830);
nor U6443 (N_6443,N_4896,N_4989);
nor U6444 (N_6444,N_4797,N_5680);
or U6445 (N_6445,N_5992,N_5622);
nand U6446 (N_6446,N_5420,N_5259);
xor U6447 (N_6447,N_5098,N_4519);
nand U6448 (N_6448,N_5467,N_4767);
or U6449 (N_6449,N_4731,N_4517);
or U6450 (N_6450,N_4764,N_5787);
xor U6451 (N_6451,N_4753,N_4895);
and U6452 (N_6452,N_4963,N_5860);
or U6453 (N_6453,N_4853,N_5453);
nand U6454 (N_6454,N_5930,N_5841);
nand U6455 (N_6455,N_5001,N_5312);
or U6456 (N_6456,N_5015,N_5342);
or U6457 (N_6457,N_5872,N_4739);
nor U6458 (N_6458,N_5957,N_5454);
nand U6459 (N_6459,N_4924,N_5748);
and U6460 (N_6460,N_4990,N_5344);
nor U6461 (N_6461,N_5438,N_5092);
nand U6462 (N_6462,N_5747,N_5765);
nor U6463 (N_6463,N_4748,N_4918);
or U6464 (N_6464,N_5540,N_4833);
nand U6465 (N_6465,N_5863,N_5488);
nor U6466 (N_6466,N_4657,N_5356);
and U6467 (N_6467,N_4780,N_5306);
xor U6468 (N_6468,N_4900,N_4704);
xnor U6469 (N_6469,N_5451,N_5919);
nor U6470 (N_6470,N_5170,N_4530);
nor U6471 (N_6471,N_5135,N_5184);
nand U6472 (N_6472,N_4943,N_4612);
or U6473 (N_6473,N_4528,N_4962);
nor U6474 (N_6474,N_4621,N_5320);
and U6475 (N_6475,N_5707,N_4880);
nor U6476 (N_6476,N_5907,N_5484);
nor U6477 (N_6477,N_5116,N_5752);
or U6478 (N_6478,N_5874,N_5166);
nor U6479 (N_6479,N_5909,N_5676);
or U6480 (N_6480,N_4807,N_4968);
and U6481 (N_6481,N_5605,N_5952);
and U6482 (N_6482,N_4563,N_5213);
or U6483 (N_6483,N_4645,N_4733);
or U6484 (N_6484,N_4700,N_5597);
nand U6485 (N_6485,N_5110,N_5530);
nand U6486 (N_6486,N_5122,N_5246);
nand U6487 (N_6487,N_5076,N_4790);
or U6488 (N_6488,N_5286,N_5140);
nand U6489 (N_6489,N_5489,N_4813);
nand U6490 (N_6490,N_5661,N_5714);
and U6491 (N_6491,N_5314,N_4520);
nand U6492 (N_6492,N_5939,N_5768);
and U6493 (N_6493,N_5604,N_5870);
nor U6494 (N_6494,N_5361,N_5175);
nor U6495 (N_6495,N_4500,N_4549);
or U6496 (N_6496,N_5375,N_5329);
nand U6497 (N_6497,N_5124,N_5587);
nor U6498 (N_6498,N_5434,N_4575);
nor U6499 (N_6499,N_5544,N_5056);
and U6500 (N_6500,N_5350,N_5718);
and U6501 (N_6501,N_4996,N_5458);
and U6502 (N_6502,N_5389,N_5775);
nand U6503 (N_6503,N_5422,N_4686);
and U6504 (N_6504,N_5885,N_5141);
or U6505 (N_6505,N_5503,N_5147);
nor U6506 (N_6506,N_5414,N_5704);
nor U6507 (N_6507,N_4626,N_4889);
nand U6508 (N_6508,N_5576,N_5594);
nand U6509 (N_6509,N_5114,N_5708);
and U6510 (N_6510,N_5891,N_5216);
and U6511 (N_6511,N_5250,N_5826);
and U6512 (N_6512,N_5445,N_4564);
nor U6513 (N_6513,N_4647,N_5516);
nor U6514 (N_6514,N_5743,N_5081);
nand U6515 (N_6515,N_5578,N_5819);
nand U6516 (N_6516,N_5837,N_4788);
nand U6517 (N_6517,N_5943,N_5441);
xor U6518 (N_6518,N_4697,N_5100);
or U6519 (N_6519,N_4658,N_5534);
nor U6520 (N_6520,N_4824,N_5241);
and U6521 (N_6521,N_4742,N_5133);
nor U6522 (N_6522,N_4912,N_5178);
xor U6523 (N_6523,N_5063,N_4814);
or U6524 (N_6524,N_4982,N_4665);
nand U6525 (N_6525,N_4566,N_5774);
nor U6526 (N_6526,N_5095,N_4525);
and U6527 (N_6527,N_4858,N_5143);
xnor U6528 (N_6528,N_5473,N_5406);
and U6529 (N_6529,N_4820,N_5975);
or U6530 (N_6530,N_5912,N_4691);
and U6531 (N_6531,N_5866,N_5777);
or U6532 (N_6532,N_5896,N_4673);
nand U6533 (N_6533,N_5279,N_4717);
nand U6534 (N_6534,N_5411,N_5410);
nand U6535 (N_6535,N_4729,N_5155);
xor U6536 (N_6536,N_5476,N_4537);
xor U6537 (N_6537,N_4850,N_5307);
xnor U6538 (N_6538,N_5584,N_4979);
and U6539 (N_6539,N_4967,N_5509);
and U6540 (N_6540,N_5684,N_5933);
and U6541 (N_6541,N_4542,N_5822);
and U6542 (N_6542,N_5227,N_5377);
or U6543 (N_6543,N_4568,N_5553);
xnor U6544 (N_6544,N_5444,N_5513);
nor U6545 (N_6545,N_5111,N_5055);
nand U6546 (N_6546,N_5404,N_5525);
nor U6547 (N_6547,N_4531,N_5378);
nand U6548 (N_6548,N_4650,N_5508);
or U6549 (N_6549,N_4857,N_4938);
nand U6550 (N_6550,N_5190,N_5873);
nand U6551 (N_6551,N_5751,N_5652);
and U6552 (N_6552,N_5031,N_5083);
nand U6553 (N_6553,N_5254,N_5614);
or U6554 (N_6554,N_4555,N_4942);
and U6555 (N_6555,N_5832,N_4875);
and U6556 (N_6556,N_5069,N_5890);
xor U6557 (N_6557,N_4981,N_4512);
and U6558 (N_6558,N_4644,N_5169);
xnor U6559 (N_6559,N_4708,N_5725);
nand U6560 (N_6560,N_5541,N_5269);
and U6561 (N_6561,N_4639,N_5635);
or U6562 (N_6562,N_4787,N_5958);
and U6563 (N_6563,N_5721,N_5322);
xor U6564 (N_6564,N_4569,N_5599);
and U6565 (N_6565,N_5946,N_4616);
xor U6566 (N_6566,N_4792,N_5571);
nand U6567 (N_6567,N_4997,N_5412);
nand U6568 (N_6568,N_5783,N_5273);
and U6569 (N_6569,N_5298,N_4874);
nor U6570 (N_6570,N_5712,N_5951);
and U6571 (N_6571,N_4633,N_4693);
or U6572 (N_6572,N_5999,N_5217);
nor U6573 (N_6573,N_5125,N_4823);
nand U6574 (N_6574,N_5029,N_5379);
nand U6575 (N_6575,N_5270,N_5096);
xnor U6576 (N_6576,N_4756,N_5006);
nand U6577 (N_6577,N_4803,N_5817);
nor U6578 (N_6578,N_5245,N_5753);
or U6579 (N_6579,N_5572,N_5828);
nand U6580 (N_6580,N_5869,N_5825);
xor U6581 (N_6581,N_5968,N_5659);
or U6582 (N_6582,N_4953,N_5723);
nand U6583 (N_6583,N_5030,N_4727);
nor U6584 (N_6584,N_5210,N_5989);
or U6585 (N_6585,N_4887,N_5816);
or U6586 (N_6586,N_5580,N_4746);
or U6587 (N_6587,N_4991,N_5913);
nand U6588 (N_6588,N_4984,N_5046);
nand U6589 (N_6589,N_5823,N_4653);
or U6590 (N_6590,N_5630,N_5447);
and U6591 (N_6591,N_5586,N_5624);
or U6592 (N_6592,N_5727,N_4772);
and U6593 (N_6593,N_5640,N_5433);
or U6594 (N_6594,N_5160,N_5323);
and U6595 (N_6595,N_5829,N_5283);
nor U6596 (N_6596,N_5963,N_4581);
and U6597 (N_6597,N_5666,N_4816);
xor U6598 (N_6598,N_5699,N_5772);
or U6599 (N_6599,N_5108,N_5811);
and U6600 (N_6600,N_4533,N_5168);
nand U6601 (N_6601,N_4641,N_5803);
and U6602 (N_6602,N_4885,N_4681);
nand U6603 (N_6603,N_5887,N_5610);
and U6604 (N_6604,N_4958,N_5545);
nand U6605 (N_6605,N_5724,N_4635);
nor U6606 (N_6606,N_5518,N_5163);
and U6607 (N_6607,N_5131,N_5478);
xnor U6608 (N_6608,N_5653,N_4776);
and U6609 (N_6609,N_5317,N_5011);
and U6610 (N_6610,N_4685,N_5814);
xor U6611 (N_6611,N_4702,N_5264);
or U6612 (N_6612,N_5496,N_4801);
xnor U6613 (N_6613,N_4628,N_5291);
or U6614 (N_6614,N_5588,N_5970);
xnor U6615 (N_6615,N_5009,N_5237);
or U6616 (N_6616,N_5590,N_5234);
xor U6617 (N_6617,N_5487,N_5333);
and U6618 (N_6618,N_4714,N_5533);
or U6619 (N_6619,N_5374,N_5771);
or U6620 (N_6620,N_5090,N_5669);
or U6621 (N_6621,N_5351,N_4611);
and U6622 (N_6622,N_5827,N_5068);
and U6623 (N_6623,N_4832,N_4843);
nand U6624 (N_6624,N_5366,N_5603);
or U6625 (N_6625,N_5465,N_5564);
nor U6626 (N_6626,N_5310,N_5522);
and U6627 (N_6627,N_4798,N_5176);
xnor U6628 (N_6628,N_4646,N_4678);
or U6629 (N_6629,N_4605,N_5345);
nand U6630 (N_6630,N_5325,N_5694);
xnor U6631 (N_6631,N_4572,N_4574);
nor U6632 (N_6632,N_5464,N_5796);
nand U6633 (N_6633,N_4716,N_5876);
nor U6634 (N_6634,N_5899,N_5424);
or U6635 (N_6635,N_4586,N_5358);
or U6636 (N_6636,N_5690,N_5253);
nor U6637 (N_6637,N_5172,N_5983);
or U6638 (N_6638,N_4854,N_4959);
or U6639 (N_6639,N_4588,N_5357);
nand U6640 (N_6640,N_4859,N_4786);
and U6641 (N_6641,N_4866,N_5591);
nor U6642 (N_6642,N_5790,N_5929);
or U6643 (N_6643,N_4781,N_4670);
and U6644 (N_6644,N_5277,N_5871);
nor U6645 (N_6645,N_5581,N_4558);
nand U6646 (N_6646,N_4744,N_5713);
nor U6647 (N_6647,N_4712,N_5695);
and U6648 (N_6648,N_4503,N_5186);
and U6649 (N_6649,N_4993,N_5380);
nor U6650 (N_6650,N_4904,N_5121);
nand U6651 (N_6651,N_5824,N_4868);
nor U6652 (N_6652,N_5838,N_5328);
nand U6653 (N_6653,N_4987,N_4701);
and U6654 (N_6654,N_5249,N_5053);
nand U6655 (N_6655,N_5421,N_5257);
and U6656 (N_6656,N_4862,N_5593);
and U6657 (N_6657,N_5634,N_5585);
and U6658 (N_6658,N_5220,N_5547);
or U6659 (N_6659,N_5577,N_5865);
xor U6660 (N_6660,N_4677,N_5230);
nand U6661 (N_6661,N_5700,N_5373);
or U6662 (N_6662,N_5974,N_5007);
nand U6663 (N_6663,N_5985,N_5103);
and U6664 (N_6664,N_5914,N_5432);
and U6665 (N_6665,N_5177,N_4710);
xor U6666 (N_6666,N_5498,N_5786);
nor U6667 (N_6667,N_4726,N_5413);
xor U6668 (N_6668,N_5918,N_4577);
and U6669 (N_6669,N_4529,N_5647);
nand U6670 (N_6670,N_5589,N_5082);
or U6671 (N_6671,N_5598,N_4723);
or U6672 (N_6672,N_5502,N_4763);
nand U6673 (N_6673,N_5932,N_5132);
or U6674 (N_6674,N_5608,N_5196);
xnor U6675 (N_6675,N_5280,N_4692);
nor U6676 (N_6676,N_5146,N_5288);
xnor U6677 (N_6677,N_5849,N_5901);
nand U6678 (N_6678,N_4973,N_4545);
nand U6679 (N_6679,N_4842,N_5944);
nor U6680 (N_6680,N_5005,N_5396);
nand U6681 (N_6681,N_5150,N_5372);
or U6682 (N_6682,N_5601,N_5294);
and U6683 (N_6683,N_5167,N_5715);
nand U6684 (N_6684,N_4975,N_4682);
and U6685 (N_6685,N_5211,N_5182);
nor U6686 (N_6686,N_5302,N_4538);
nand U6687 (N_6687,N_5233,N_4796);
or U6688 (N_6688,N_4599,N_4995);
or U6689 (N_6689,N_4524,N_4847);
and U6690 (N_6690,N_5855,N_5800);
or U6691 (N_6691,N_5419,N_5349);
nor U6692 (N_6692,N_4951,N_5117);
nor U6693 (N_6693,N_4578,N_4625);
nand U6694 (N_6694,N_4873,N_5113);
and U6695 (N_6695,N_4848,N_5750);
nand U6696 (N_6696,N_5967,N_4627);
xnor U6697 (N_6697,N_5716,N_5671);
or U6698 (N_6698,N_5638,N_5174);
nand U6699 (N_6699,N_4679,N_5179);
xnor U6700 (N_6700,N_5867,N_5265);
and U6701 (N_6701,N_5681,N_5739);
nand U6702 (N_6702,N_4882,N_5363);
xnor U6703 (N_6703,N_5059,N_4937);
nand U6704 (N_6704,N_5685,N_5079);
or U6705 (N_6705,N_5668,N_5926);
nand U6706 (N_6706,N_5971,N_5511);
nor U6707 (N_6707,N_4511,N_5657);
nor U6708 (N_6708,N_5232,N_5579);
nor U6709 (N_6709,N_4961,N_4743);
nor U6710 (N_6710,N_4629,N_5698);
nor U6711 (N_6711,N_5278,N_4769);
xnor U6712 (N_6712,N_5701,N_5475);
or U6713 (N_6713,N_5461,N_4523);
xnor U6714 (N_6714,N_5732,N_4614);
or U6715 (N_6715,N_5711,N_5888);
and U6716 (N_6716,N_4741,N_5191);
nand U6717 (N_6717,N_5013,N_5290);
or U6718 (N_6718,N_5303,N_5616);
and U6719 (N_6719,N_5157,N_5231);
nor U6720 (N_6720,N_5945,N_5688);
nand U6721 (N_6721,N_4960,N_4921);
nor U6722 (N_6722,N_5510,N_4740);
nand U6723 (N_6723,N_4920,N_4879);
and U6724 (N_6724,N_5792,N_5927);
xnor U6725 (N_6725,N_5267,N_5879);
xor U6726 (N_6726,N_5407,N_5643);
and U6727 (N_6727,N_4654,N_5084);
and U6728 (N_6728,N_4661,N_5596);
or U6729 (N_6729,N_5923,N_5436);
nor U6730 (N_6730,N_5199,N_4515);
nand U6731 (N_6731,N_4557,N_4779);
and U6732 (N_6732,N_4822,N_5757);
xnor U6733 (N_6733,N_4759,N_5072);
nor U6734 (N_6734,N_4891,N_4872);
or U6735 (N_6735,N_4694,N_4841);
nand U6736 (N_6736,N_5164,N_4516);
or U6737 (N_6737,N_4819,N_4839);
and U6738 (N_6738,N_4948,N_5091);
xor U6739 (N_6739,N_5295,N_5430);
and U6740 (N_6740,N_5016,N_5806);
and U6741 (N_6741,N_5801,N_5327);
nand U6742 (N_6742,N_5426,N_5990);
and U6743 (N_6743,N_5655,N_4703);
xor U6744 (N_6744,N_5238,N_5702);
nand U6745 (N_6745,N_4711,N_5642);
and U6746 (N_6746,N_5813,N_5749);
and U6747 (N_6747,N_5040,N_4582);
or U6748 (N_6748,N_5483,N_5620);
or U6749 (N_6749,N_5782,N_5448);
nor U6750 (N_6750,N_4511,N_5524);
and U6751 (N_6751,N_5141,N_5380);
xor U6752 (N_6752,N_5441,N_5749);
xnor U6753 (N_6753,N_5188,N_5686);
and U6754 (N_6754,N_5233,N_5213);
and U6755 (N_6755,N_4987,N_5129);
nand U6756 (N_6756,N_5940,N_5869);
nor U6757 (N_6757,N_4953,N_5073);
nor U6758 (N_6758,N_4934,N_5652);
nor U6759 (N_6759,N_5973,N_5996);
nand U6760 (N_6760,N_4556,N_5650);
or U6761 (N_6761,N_5862,N_5179);
or U6762 (N_6762,N_4969,N_5075);
nor U6763 (N_6763,N_5128,N_5601);
nor U6764 (N_6764,N_4871,N_5411);
and U6765 (N_6765,N_4596,N_4940);
nand U6766 (N_6766,N_5956,N_5708);
nand U6767 (N_6767,N_5560,N_5570);
or U6768 (N_6768,N_5120,N_4953);
nor U6769 (N_6769,N_5722,N_5383);
nor U6770 (N_6770,N_4606,N_5954);
nand U6771 (N_6771,N_5464,N_5185);
nand U6772 (N_6772,N_5625,N_5858);
nand U6773 (N_6773,N_5733,N_4660);
and U6774 (N_6774,N_4690,N_5170);
nor U6775 (N_6775,N_4962,N_5020);
nor U6776 (N_6776,N_5828,N_5911);
nor U6777 (N_6777,N_4825,N_4981);
nor U6778 (N_6778,N_4591,N_4628);
nand U6779 (N_6779,N_5188,N_5285);
or U6780 (N_6780,N_5998,N_4925);
or U6781 (N_6781,N_5151,N_5383);
nand U6782 (N_6782,N_4556,N_4595);
nor U6783 (N_6783,N_4552,N_5281);
or U6784 (N_6784,N_5813,N_5600);
or U6785 (N_6785,N_4528,N_5067);
nor U6786 (N_6786,N_4632,N_4978);
nand U6787 (N_6787,N_4543,N_5223);
xnor U6788 (N_6788,N_5049,N_4848);
or U6789 (N_6789,N_4550,N_5462);
nor U6790 (N_6790,N_4971,N_4927);
nand U6791 (N_6791,N_5093,N_5934);
or U6792 (N_6792,N_5461,N_5583);
and U6793 (N_6793,N_5285,N_5903);
xnor U6794 (N_6794,N_4947,N_5967);
nand U6795 (N_6795,N_4857,N_5151);
nor U6796 (N_6796,N_5008,N_4704);
and U6797 (N_6797,N_5095,N_4922);
nor U6798 (N_6798,N_5370,N_5660);
nand U6799 (N_6799,N_4962,N_5840);
xnor U6800 (N_6800,N_5057,N_4865);
nand U6801 (N_6801,N_5608,N_5182);
and U6802 (N_6802,N_4603,N_4529);
nand U6803 (N_6803,N_5002,N_5845);
or U6804 (N_6804,N_5708,N_5719);
or U6805 (N_6805,N_5149,N_4834);
or U6806 (N_6806,N_5922,N_5771);
xor U6807 (N_6807,N_5193,N_5116);
nand U6808 (N_6808,N_5265,N_5525);
nand U6809 (N_6809,N_5279,N_5284);
xor U6810 (N_6810,N_4724,N_4564);
xor U6811 (N_6811,N_4711,N_5969);
and U6812 (N_6812,N_5101,N_4922);
and U6813 (N_6813,N_4987,N_5016);
xor U6814 (N_6814,N_5245,N_5365);
nand U6815 (N_6815,N_5542,N_4678);
or U6816 (N_6816,N_5004,N_4831);
nand U6817 (N_6817,N_5087,N_4947);
nand U6818 (N_6818,N_5633,N_5305);
nand U6819 (N_6819,N_4584,N_5477);
or U6820 (N_6820,N_5562,N_4964);
xor U6821 (N_6821,N_4937,N_5336);
xor U6822 (N_6822,N_5868,N_5999);
xnor U6823 (N_6823,N_5747,N_4913);
or U6824 (N_6824,N_4645,N_5863);
xnor U6825 (N_6825,N_5625,N_5127);
xor U6826 (N_6826,N_5136,N_5081);
and U6827 (N_6827,N_5976,N_5828);
or U6828 (N_6828,N_5798,N_5342);
xnor U6829 (N_6829,N_4829,N_4664);
nand U6830 (N_6830,N_4886,N_4799);
and U6831 (N_6831,N_4526,N_5643);
and U6832 (N_6832,N_4751,N_5555);
or U6833 (N_6833,N_5858,N_5395);
nand U6834 (N_6834,N_5410,N_4724);
and U6835 (N_6835,N_5043,N_4540);
nor U6836 (N_6836,N_5229,N_5843);
nand U6837 (N_6837,N_4645,N_4684);
or U6838 (N_6838,N_4652,N_5781);
xnor U6839 (N_6839,N_5717,N_5822);
nand U6840 (N_6840,N_4675,N_5011);
nand U6841 (N_6841,N_5029,N_4905);
nand U6842 (N_6842,N_4739,N_5210);
or U6843 (N_6843,N_5235,N_5091);
or U6844 (N_6844,N_5752,N_4990);
xor U6845 (N_6845,N_4741,N_4892);
nand U6846 (N_6846,N_5332,N_5717);
nand U6847 (N_6847,N_5735,N_5277);
nand U6848 (N_6848,N_5427,N_4554);
or U6849 (N_6849,N_4997,N_5329);
nand U6850 (N_6850,N_4975,N_5023);
or U6851 (N_6851,N_4535,N_5921);
nand U6852 (N_6852,N_4774,N_5668);
and U6853 (N_6853,N_4883,N_4501);
or U6854 (N_6854,N_5750,N_5662);
nor U6855 (N_6855,N_5355,N_4532);
and U6856 (N_6856,N_5336,N_4859);
nor U6857 (N_6857,N_5322,N_4551);
or U6858 (N_6858,N_4685,N_5079);
and U6859 (N_6859,N_4765,N_5864);
and U6860 (N_6860,N_4850,N_5150);
or U6861 (N_6861,N_5511,N_5537);
nand U6862 (N_6862,N_5523,N_5608);
and U6863 (N_6863,N_5714,N_4820);
and U6864 (N_6864,N_5766,N_5131);
nand U6865 (N_6865,N_4935,N_5408);
nand U6866 (N_6866,N_5388,N_5127);
and U6867 (N_6867,N_5025,N_5278);
xnor U6868 (N_6868,N_4565,N_5799);
nor U6869 (N_6869,N_4729,N_5399);
or U6870 (N_6870,N_5531,N_5503);
and U6871 (N_6871,N_5052,N_4570);
xor U6872 (N_6872,N_4869,N_4572);
nor U6873 (N_6873,N_5667,N_5613);
and U6874 (N_6874,N_4973,N_4816);
xnor U6875 (N_6875,N_5106,N_5323);
or U6876 (N_6876,N_5033,N_5924);
or U6877 (N_6877,N_5741,N_4559);
and U6878 (N_6878,N_5503,N_5839);
and U6879 (N_6879,N_4601,N_5867);
nor U6880 (N_6880,N_4658,N_5685);
nand U6881 (N_6881,N_4510,N_5400);
and U6882 (N_6882,N_5953,N_4670);
or U6883 (N_6883,N_4755,N_5841);
or U6884 (N_6884,N_4620,N_5411);
nor U6885 (N_6885,N_5214,N_4591);
nor U6886 (N_6886,N_5402,N_4889);
or U6887 (N_6887,N_5715,N_5233);
or U6888 (N_6888,N_5027,N_4742);
and U6889 (N_6889,N_5168,N_4699);
nand U6890 (N_6890,N_5707,N_5680);
nand U6891 (N_6891,N_5086,N_5262);
nor U6892 (N_6892,N_4867,N_5500);
nor U6893 (N_6893,N_5684,N_5611);
or U6894 (N_6894,N_5453,N_5379);
nor U6895 (N_6895,N_5215,N_5789);
or U6896 (N_6896,N_5697,N_5059);
and U6897 (N_6897,N_4577,N_5157);
nor U6898 (N_6898,N_5892,N_5368);
and U6899 (N_6899,N_5207,N_5349);
nand U6900 (N_6900,N_5353,N_5943);
nand U6901 (N_6901,N_4995,N_5001);
xor U6902 (N_6902,N_5420,N_5998);
or U6903 (N_6903,N_5280,N_5071);
nand U6904 (N_6904,N_5149,N_5028);
or U6905 (N_6905,N_5150,N_5505);
nand U6906 (N_6906,N_5802,N_4509);
xnor U6907 (N_6907,N_4527,N_4737);
or U6908 (N_6908,N_5240,N_5467);
or U6909 (N_6909,N_5528,N_5451);
nor U6910 (N_6910,N_5402,N_5188);
nor U6911 (N_6911,N_4594,N_5255);
or U6912 (N_6912,N_5612,N_4943);
and U6913 (N_6913,N_4664,N_5426);
and U6914 (N_6914,N_5630,N_4799);
nand U6915 (N_6915,N_4803,N_4811);
nand U6916 (N_6916,N_5958,N_4552);
nand U6917 (N_6917,N_5702,N_4864);
and U6918 (N_6918,N_5072,N_5834);
nor U6919 (N_6919,N_4774,N_5822);
nand U6920 (N_6920,N_4657,N_4546);
or U6921 (N_6921,N_5582,N_5003);
nor U6922 (N_6922,N_4715,N_5749);
nor U6923 (N_6923,N_4532,N_5476);
or U6924 (N_6924,N_4586,N_5832);
nor U6925 (N_6925,N_5157,N_5046);
or U6926 (N_6926,N_5198,N_5687);
nor U6927 (N_6927,N_4507,N_5992);
xor U6928 (N_6928,N_5469,N_5280);
and U6929 (N_6929,N_5783,N_4976);
nand U6930 (N_6930,N_5335,N_5670);
and U6931 (N_6931,N_5467,N_5156);
and U6932 (N_6932,N_4836,N_5029);
or U6933 (N_6933,N_4782,N_5222);
nand U6934 (N_6934,N_4701,N_5561);
nand U6935 (N_6935,N_5820,N_5206);
nand U6936 (N_6936,N_4631,N_5049);
nand U6937 (N_6937,N_5090,N_5461);
or U6938 (N_6938,N_4624,N_5503);
xnor U6939 (N_6939,N_5862,N_5913);
nor U6940 (N_6940,N_5701,N_5642);
nor U6941 (N_6941,N_5076,N_5558);
nor U6942 (N_6942,N_5202,N_5695);
or U6943 (N_6943,N_5083,N_5650);
and U6944 (N_6944,N_5644,N_5136);
nor U6945 (N_6945,N_5186,N_5791);
nor U6946 (N_6946,N_5123,N_5675);
and U6947 (N_6947,N_4989,N_5909);
and U6948 (N_6948,N_5030,N_4846);
nor U6949 (N_6949,N_5912,N_5925);
nand U6950 (N_6950,N_5343,N_4581);
or U6951 (N_6951,N_5100,N_5516);
xnor U6952 (N_6952,N_4955,N_5370);
nand U6953 (N_6953,N_5849,N_4530);
or U6954 (N_6954,N_5053,N_5515);
xor U6955 (N_6955,N_4973,N_5432);
and U6956 (N_6956,N_5727,N_4886);
nand U6957 (N_6957,N_5881,N_4742);
nor U6958 (N_6958,N_4595,N_4506);
and U6959 (N_6959,N_4790,N_5039);
or U6960 (N_6960,N_4934,N_5487);
xor U6961 (N_6961,N_4894,N_5672);
nor U6962 (N_6962,N_4737,N_5249);
or U6963 (N_6963,N_4607,N_5813);
and U6964 (N_6964,N_4827,N_5831);
or U6965 (N_6965,N_5715,N_4875);
nand U6966 (N_6966,N_4850,N_5821);
or U6967 (N_6967,N_5147,N_5184);
and U6968 (N_6968,N_4930,N_5642);
and U6969 (N_6969,N_4586,N_5908);
and U6970 (N_6970,N_4659,N_5325);
or U6971 (N_6971,N_5172,N_5616);
nand U6972 (N_6972,N_4913,N_5774);
or U6973 (N_6973,N_4737,N_5059);
and U6974 (N_6974,N_4853,N_5907);
or U6975 (N_6975,N_5892,N_5432);
xor U6976 (N_6976,N_5911,N_5688);
nand U6977 (N_6977,N_5132,N_5177);
nor U6978 (N_6978,N_5914,N_4763);
and U6979 (N_6979,N_4766,N_4986);
nor U6980 (N_6980,N_4793,N_5738);
and U6981 (N_6981,N_4803,N_5625);
nor U6982 (N_6982,N_5224,N_4887);
or U6983 (N_6983,N_5396,N_5940);
xnor U6984 (N_6984,N_5723,N_4755);
or U6985 (N_6985,N_5607,N_4684);
nand U6986 (N_6986,N_5293,N_4920);
xnor U6987 (N_6987,N_5357,N_5959);
and U6988 (N_6988,N_4895,N_5371);
and U6989 (N_6989,N_5618,N_5671);
nand U6990 (N_6990,N_5965,N_5953);
and U6991 (N_6991,N_5152,N_4670);
or U6992 (N_6992,N_5001,N_4949);
or U6993 (N_6993,N_5641,N_4961);
or U6994 (N_6994,N_4603,N_4637);
nor U6995 (N_6995,N_4587,N_5002);
nand U6996 (N_6996,N_5732,N_5718);
and U6997 (N_6997,N_4584,N_4893);
nand U6998 (N_6998,N_4702,N_5544);
nand U6999 (N_6999,N_5646,N_5130);
nand U7000 (N_7000,N_5819,N_4611);
nor U7001 (N_7001,N_4794,N_4887);
nand U7002 (N_7002,N_5763,N_4768);
nor U7003 (N_7003,N_5468,N_5569);
and U7004 (N_7004,N_4714,N_5171);
and U7005 (N_7005,N_5866,N_5895);
nor U7006 (N_7006,N_5342,N_5099);
xor U7007 (N_7007,N_5955,N_5683);
and U7008 (N_7008,N_4963,N_4896);
nor U7009 (N_7009,N_5609,N_4604);
nor U7010 (N_7010,N_5619,N_5043);
nor U7011 (N_7011,N_5782,N_4539);
nand U7012 (N_7012,N_4865,N_5455);
nor U7013 (N_7013,N_5395,N_5526);
nand U7014 (N_7014,N_5548,N_5396);
or U7015 (N_7015,N_4624,N_5360);
and U7016 (N_7016,N_4847,N_5531);
or U7017 (N_7017,N_4506,N_5836);
or U7018 (N_7018,N_4602,N_4654);
or U7019 (N_7019,N_5121,N_4987);
nand U7020 (N_7020,N_5835,N_5258);
and U7021 (N_7021,N_4785,N_5221);
or U7022 (N_7022,N_5673,N_5819);
and U7023 (N_7023,N_5577,N_5607);
nand U7024 (N_7024,N_5360,N_5359);
and U7025 (N_7025,N_5686,N_5358);
or U7026 (N_7026,N_4869,N_5374);
nor U7027 (N_7027,N_4802,N_4695);
and U7028 (N_7028,N_5051,N_5315);
nand U7029 (N_7029,N_5760,N_4912);
or U7030 (N_7030,N_5675,N_5967);
or U7031 (N_7031,N_4737,N_4717);
nand U7032 (N_7032,N_5912,N_5286);
nor U7033 (N_7033,N_5144,N_4709);
nor U7034 (N_7034,N_5711,N_5101);
nor U7035 (N_7035,N_4696,N_5228);
nand U7036 (N_7036,N_5059,N_5906);
nand U7037 (N_7037,N_5204,N_5801);
nor U7038 (N_7038,N_5462,N_4658);
nor U7039 (N_7039,N_5378,N_5524);
nand U7040 (N_7040,N_5842,N_4900);
and U7041 (N_7041,N_4855,N_4680);
nor U7042 (N_7042,N_5347,N_4507);
nor U7043 (N_7043,N_5806,N_5664);
and U7044 (N_7044,N_5620,N_5900);
nor U7045 (N_7045,N_4770,N_5572);
and U7046 (N_7046,N_5502,N_4807);
nor U7047 (N_7047,N_4616,N_4691);
nor U7048 (N_7048,N_5416,N_4869);
nand U7049 (N_7049,N_5896,N_4593);
and U7050 (N_7050,N_4533,N_4792);
or U7051 (N_7051,N_5864,N_5102);
nand U7052 (N_7052,N_5522,N_5797);
nand U7053 (N_7053,N_5053,N_4838);
and U7054 (N_7054,N_5396,N_5896);
or U7055 (N_7055,N_5622,N_5896);
xnor U7056 (N_7056,N_5654,N_5229);
or U7057 (N_7057,N_5454,N_4638);
nand U7058 (N_7058,N_5673,N_5063);
and U7059 (N_7059,N_5758,N_5158);
nand U7060 (N_7060,N_5271,N_5587);
or U7061 (N_7061,N_4881,N_5845);
or U7062 (N_7062,N_5184,N_5241);
xor U7063 (N_7063,N_5133,N_5963);
or U7064 (N_7064,N_4728,N_5146);
nand U7065 (N_7065,N_4798,N_4959);
nand U7066 (N_7066,N_4829,N_4967);
nor U7067 (N_7067,N_5482,N_5516);
nor U7068 (N_7068,N_5117,N_5539);
and U7069 (N_7069,N_5556,N_4692);
xor U7070 (N_7070,N_5754,N_5785);
nand U7071 (N_7071,N_5261,N_5959);
or U7072 (N_7072,N_4857,N_5180);
nand U7073 (N_7073,N_4529,N_4722);
nand U7074 (N_7074,N_5622,N_5724);
or U7075 (N_7075,N_5385,N_4676);
and U7076 (N_7076,N_5769,N_5735);
nor U7077 (N_7077,N_4563,N_5594);
nor U7078 (N_7078,N_5290,N_5475);
and U7079 (N_7079,N_4856,N_5352);
nor U7080 (N_7080,N_4799,N_4846);
and U7081 (N_7081,N_4638,N_4863);
nor U7082 (N_7082,N_5143,N_5223);
nand U7083 (N_7083,N_5343,N_5356);
nand U7084 (N_7084,N_4708,N_5230);
or U7085 (N_7085,N_5230,N_4648);
or U7086 (N_7086,N_5469,N_5391);
and U7087 (N_7087,N_5605,N_5342);
xnor U7088 (N_7088,N_5403,N_5379);
or U7089 (N_7089,N_5297,N_5266);
nand U7090 (N_7090,N_5423,N_5778);
and U7091 (N_7091,N_5015,N_5320);
nand U7092 (N_7092,N_5812,N_5938);
nand U7093 (N_7093,N_5634,N_5904);
or U7094 (N_7094,N_5591,N_4913);
and U7095 (N_7095,N_5001,N_5448);
and U7096 (N_7096,N_4529,N_4996);
nand U7097 (N_7097,N_5252,N_5755);
xor U7098 (N_7098,N_4545,N_4855);
or U7099 (N_7099,N_5923,N_5660);
or U7100 (N_7100,N_5979,N_5006);
and U7101 (N_7101,N_4930,N_5338);
nor U7102 (N_7102,N_4994,N_5389);
xor U7103 (N_7103,N_5281,N_5086);
nor U7104 (N_7104,N_4629,N_4835);
xor U7105 (N_7105,N_5518,N_5800);
or U7106 (N_7106,N_5892,N_5094);
nand U7107 (N_7107,N_4713,N_4574);
nand U7108 (N_7108,N_4642,N_5240);
nand U7109 (N_7109,N_5936,N_5037);
or U7110 (N_7110,N_4847,N_5608);
and U7111 (N_7111,N_5677,N_5564);
nor U7112 (N_7112,N_5154,N_4970);
nor U7113 (N_7113,N_4505,N_4694);
nor U7114 (N_7114,N_5090,N_4944);
or U7115 (N_7115,N_5084,N_5757);
nand U7116 (N_7116,N_5994,N_4842);
and U7117 (N_7117,N_4943,N_5699);
nor U7118 (N_7118,N_5882,N_5540);
or U7119 (N_7119,N_5348,N_4981);
nand U7120 (N_7120,N_4709,N_4525);
nand U7121 (N_7121,N_5543,N_5587);
and U7122 (N_7122,N_5401,N_5356);
nand U7123 (N_7123,N_4652,N_5811);
nor U7124 (N_7124,N_5036,N_4845);
or U7125 (N_7125,N_4889,N_5648);
nand U7126 (N_7126,N_5165,N_4762);
and U7127 (N_7127,N_5042,N_5801);
nor U7128 (N_7128,N_4742,N_5109);
and U7129 (N_7129,N_5544,N_4603);
or U7130 (N_7130,N_5199,N_5580);
nor U7131 (N_7131,N_5273,N_5078);
xor U7132 (N_7132,N_5917,N_5955);
and U7133 (N_7133,N_4702,N_4864);
nor U7134 (N_7134,N_5235,N_5198);
nand U7135 (N_7135,N_4633,N_5458);
or U7136 (N_7136,N_5580,N_5082);
or U7137 (N_7137,N_5288,N_5919);
nand U7138 (N_7138,N_5468,N_5220);
and U7139 (N_7139,N_5096,N_5475);
xnor U7140 (N_7140,N_5411,N_5613);
nor U7141 (N_7141,N_4714,N_5894);
nor U7142 (N_7142,N_4689,N_4982);
nand U7143 (N_7143,N_4984,N_5139);
and U7144 (N_7144,N_5076,N_5179);
nand U7145 (N_7145,N_5572,N_4667);
nand U7146 (N_7146,N_5645,N_4560);
or U7147 (N_7147,N_5075,N_4690);
or U7148 (N_7148,N_5914,N_4509);
and U7149 (N_7149,N_4970,N_5839);
xnor U7150 (N_7150,N_4691,N_4902);
and U7151 (N_7151,N_4673,N_5204);
nor U7152 (N_7152,N_5170,N_5758);
and U7153 (N_7153,N_4977,N_4759);
nor U7154 (N_7154,N_5379,N_5061);
and U7155 (N_7155,N_5779,N_4773);
nor U7156 (N_7156,N_4574,N_4657);
or U7157 (N_7157,N_4743,N_4664);
or U7158 (N_7158,N_5302,N_5441);
nand U7159 (N_7159,N_4969,N_5718);
xor U7160 (N_7160,N_5242,N_4843);
or U7161 (N_7161,N_5684,N_4602);
xor U7162 (N_7162,N_5496,N_5548);
nor U7163 (N_7163,N_5655,N_4873);
and U7164 (N_7164,N_4853,N_5832);
nand U7165 (N_7165,N_5659,N_4994);
or U7166 (N_7166,N_5298,N_4881);
and U7167 (N_7167,N_5603,N_4518);
nand U7168 (N_7168,N_4810,N_5725);
xnor U7169 (N_7169,N_5446,N_5339);
nand U7170 (N_7170,N_4728,N_4814);
and U7171 (N_7171,N_5556,N_5388);
nand U7172 (N_7172,N_5179,N_4954);
nand U7173 (N_7173,N_5579,N_4991);
nand U7174 (N_7174,N_4786,N_5409);
or U7175 (N_7175,N_4690,N_4906);
and U7176 (N_7176,N_5829,N_5519);
nand U7177 (N_7177,N_5799,N_5267);
nand U7178 (N_7178,N_5931,N_5435);
nand U7179 (N_7179,N_5197,N_5255);
nand U7180 (N_7180,N_4529,N_5906);
or U7181 (N_7181,N_5539,N_5731);
and U7182 (N_7182,N_4883,N_5227);
xor U7183 (N_7183,N_5473,N_4563);
nand U7184 (N_7184,N_5072,N_5299);
and U7185 (N_7185,N_4777,N_5178);
and U7186 (N_7186,N_5639,N_4699);
nand U7187 (N_7187,N_5184,N_4731);
nand U7188 (N_7188,N_5105,N_5283);
or U7189 (N_7189,N_4673,N_5604);
or U7190 (N_7190,N_5084,N_5469);
and U7191 (N_7191,N_5424,N_4548);
nand U7192 (N_7192,N_4941,N_5785);
and U7193 (N_7193,N_5214,N_5296);
xor U7194 (N_7194,N_4887,N_5858);
and U7195 (N_7195,N_4540,N_4732);
nand U7196 (N_7196,N_5409,N_5716);
xor U7197 (N_7197,N_5966,N_5882);
nor U7198 (N_7198,N_5374,N_4818);
xor U7199 (N_7199,N_5280,N_5276);
and U7200 (N_7200,N_5183,N_4873);
nor U7201 (N_7201,N_4688,N_4900);
nor U7202 (N_7202,N_5508,N_4542);
nor U7203 (N_7203,N_5253,N_5551);
nand U7204 (N_7204,N_5734,N_4547);
and U7205 (N_7205,N_5397,N_5085);
nand U7206 (N_7206,N_5898,N_5256);
nand U7207 (N_7207,N_5586,N_5718);
and U7208 (N_7208,N_5567,N_5338);
nor U7209 (N_7209,N_5478,N_5069);
nor U7210 (N_7210,N_4774,N_4904);
or U7211 (N_7211,N_5884,N_5588);
or U7212 (N_7212,N_5063,N_4516);
nor U7213 (N_7213,N_5523,N_4666);
and U7214 (N_7214,N_5211,N_5326);
nor U7215 (N_7215,N_5174,N_5365);
and U7216 (N_7216,N_4907,N_4839);
and U7217 (N_7217,N_5294,N_4795);
nor U7218 (N_7218,N_4747,N_5648);
or U7219 (N_7219,N_5641,N_4517);
nor U7220 (N_7220,N_5410,N_4764);
and U7221 (N_7221,N_4888,N_5479);
and U7222 (N_7222,N_5452,N_4997);
nor U7223 (N_7223,N_4664,N_5929);
and U7224 (N_7224,N_4721,N_4835);
and U7225 (N_7225,N_4594,N_5010);
and U7226 (N_7226,N_5364,N_5136);
or U7227 (N_7227,N_5408,N_4774);
nor U7228 (N_7228,N_5276,N_5311);
nand U7229 (N_7229,N_5279,N_4876);
and U7230 (N_7230,N_4593,N_5532);
nor U7231 (N_7231,N_5648,N_5017);
or U7232 (N_7232,N_4728,N_5478);
nand U7233 (N_7233,N_5980,N_5818);
nand U7234 (N_7234,N_4580,N_4739);
and U7235 (N_7235,N_4520,N_4708);
or U7236 (N_7236,N_5710,N_5399);
nor U7237 (N_7237,N_4876,N_5236);
or U7238 (N_7238,N_4525,N_5515);
nand U7239 (N_7239,N_5133,N_5651);
or U7240 (N_7240,N_5687,N_5854);
and U7241 (N_7241,N_4994,N_4704);
nor U7242 (N_7242,N_5069,N_5370);
or U7243 (N_7243,N_4805,N_5950);
or U7244 (N_7244,N_5649,N_5465);
and U7245 (N_7245,N_5087,N_5767);
nor U7246 (N_7246,N_4608,N_5477);
or U7247 (N_7247,N_5763,N_4854);
nand U7248 (N_7248,N_5712,N_4830);
and U7249 (N_7249,N_5431,N_5596);
nor U7250 (N_7250,N_4812,N_4842);
xor U7251 (N_7251,N_4694,N_5504);
or U7252 (N_7252,N_5822,N_5108);
nor U7253 (N_7253,N_4874,N_5364);
nand U7254 (N_7254,N_5952,N_5532);
or U7255 (N_7255,N_5997,N_5363);
nand U7256 (N_7256,N_4946,N_5453);
xor U7257 (N_7257,N_5432,N_4949);
nand U7258 (N_7258,N_5410,N_5154);
or U7259 (N_7259,N_5323,N_5637);
nor U7260 (N_7260,N_4692,N_4556);
nor U7261 (N_7261,N_4699,N_5992);
and U7262 (N_7262,N_4880,N_5376);
and U7263 (N_7263,N_5845,N_5244);
nor U7264 (N_7264,N_5903,N_5557);
nor U7265 (N_7265,N_5851,N_5154);
nor U7266 (N_7266,N_5493,N_5686);
nand U7267 (N_7267,N_4588,N_5111);
or U7268 (N_7268,N_5467,N_4977);
or U7269 (N_7269,N_5018,N_4910);
or U7270 (N_7270,N_4658,N_4947);
and U7271 (N_7271,N_5914,N_4507);
and U7272 (N_7272,N_5849,N_5075);
nand U7273 (N_7273,N_4907,N_4605);
and U7274 (N_7274,N_5042,N_5318);
nand U7275 (N_7275,N_4717,N_4881);
nand U7276 (N_7276,N_5549,N_5770);
or U7277 (N_7277,N_5000,N_5993);
nor U7278 (N_7278,N_5426,N_5980);
or U7279 (N_7279,N_5117,N_4833);
nor U7280 (N_7280,N_5269,N_4650);
and U7281 (N_7281,N_5745,N_5733);
and U7282 (N_7282,N_4536,N_5629);
nor U7283 (N_7283,N_5652,N_5094);
and U7284 (N_7284,N_5519,N_4705);
and U7285 (N_7285,N_4784,N_5575);
nor U7286 (N_7286,N_5472,N_5360);
nand U7287 (N_7287,N_4591,N_4981);
nor U7288 (N_7288,N_4595,N_5783);
nor U7289 (N_7289,N_5581,N_4520);
nor U7290 (N_7290,N_5991,N_5106);
xor U7291 (N_7291,N_4819,N_5694);
xor U7292 (N_7292,N_4504,N_5379);
and U7293 (N_7293,N_4806,N_4649);
or U7294 (N_7294,N_4593,N_5556);
nand U7295 (N_7295,N_5739,N_4683);
nor U7296 (N_7296,N_4896,N_5500);
nand U7297 (N_7297,N_4769,N_4764);
and U7298 (N_7298,N_5279,N_5086);
and U7299 (N_7299,N_5300,N_5243);
xor U7300 (N_7300,N_4568,N_4960);
or U7301 (N_7301,N_4673,N_5124);
xnor U7302 (N_7302,N_4638,N_5870);
or U7303 (N_7303,N_5375,N_5571);
and U7304 (N_7304,N_5487,N_5447);
or U7305 (N_7305,N_5377,N_4933);
nor U7306 (N_7306,N_4937,N_5125);
nand U7307 (N_7307,N_4662,N_4559);
or U7308 (N_7308,N_4918,N_4677);
and U7309 (N_7309,N_4623,N_5568);
nor U7310 (N_7310,N_4913,N_5336);
nor U7311 (N_7311,N_4903,N_4566);
nor U7312 (N_7312,N_5021,N_5166);
nor U7313 (N_7313,N_4809,N_4762);
xnor U7314 (N_7314,N_4736,N_5696);
or U7315 (N_7315,N_5963,N_5896);
or U7316 (N_7316,N_5048,N_4512);
nand U7317 (N_7317,N_5995,N_5900);
nor U7318 (N_7318,N_4611,N_4676);
or U7319 (N_7319,N_5228,N_5466);
nand U7320 (N_7320,N_5987,N_5081);
nor U7321 (N_7321,N_4869,N_5447);
xor U7322 (N_7322,N_5931,N_5411);
nor U7323 (N_7323,N_5226,N_4879);
nand U7324 (N_7324,N_5072,N_5747);
xnor U7325 (N_7325,N_5220,N_5229);
nand U7326 (N_7326,N_5429,N_5288);
nor U7327 (N_7327,N_4679,N_5699);
nor U7328 (N_7328,N_5865,N_5686);
and U7329 (N_7329,N_5111,N_5711);
nand U7330 (N_7330,N_4876,N_5772);
or U7331 (N_7331,N_5554,N_5399);
nor U7332 (N_7332,N_5085,N_5826);
nor U7333 (N_7333,N_5398,N_5739);
nor U7334 (N_7334,N_4558,N_4694);
nor U7335 (N_7335,N_5339,N_4846);
nor U7336 (N_7336,N_5957,N_5710);
or U7337 (N_7337,N_4756,N_4677);
and U7338 (N_7338,N_4765,N_4914);
nand U7339 (N_7339,N_5637,N_4711);
nor U7340 (N_7340,N_5138,N_5152);
nand U7341 (N_7341,N_5311,N_5934);
or U7342 (N_7342,N_5533,N_4711);
xnor U7343 (N_7343,N_4672,N_5577);
or U7344 (N_7344,N_5227,N_5560);
nor U7345 (N_7345,N_5931,N_5314);
and U7346 (N_7346,N_5590,N_5746);
nand U7347 (N_7347,N_4760,N_5982);
nand U7348 (N_7348,N_4733,N_5045);
and U7349 (N_7349,N_4678,N_4510);
and U7350 (N_7350,N_4610,N_5611);
and U7351 (N_7351,N_4969,N_5215);
and U7352 (N_7352,N_5315,N_5897);
and U7353 (N_7353,N_4822,N_4632);
nor U7354 (N_7354,N_4885,N_4964);
or U7355 (N_7355,N_5103,N_4837);
or U7356 (N_7356,N_5467,N_4554);
nor U7357 (N_7357,N_4993,N_5491);
and U7358 (N_7358,N_5946,N_5967);
nor U7359 (N_7359,N_4971,N_5542);
nor U7360 (N_7360,N_4829,N_5894);
xnor U7361 (N_7361,N_4990,N_5970);
or U7362 (N_7362,N_4524,N_4542);
nor U7363 (N_7363,N_5749,N_5903);
xor U7364 (N_7364,N_4511,N_5426);
and U7365 (N_7365,N_4607,N_5378);
or U7366 (N_7366,N_5229,N_4826);
or U7367 (N_7367,N_4627,N_4516);
or U7368 (N_7368,N_4804,N_4895);
nor U7369 (N_7369,N_4714,N_5603);
xnor U7370 (N_7370,N_4757,N_5353);
and U7371 (N_7371,N_5633,N_5556);
and U7372 (N_7372,N_5882,N_5803);
nor U7373 (N_7373,N_5040,N_5353);
or U7374 (N_7374,N_5558,N_4733);
xnor U7375 (N_7375,N_5855,N_5781);
nand U7376 (N_7376,N_5084,N_4847);
nand U7377 (N_7377,N_5031,N_5801);
nor U7378 (N_7378,N_4650,N_5373);
and U7379 (N_7379,N_4613,N_4886);
and U7380 (N_7380,N_5439,N_5295);
or U7381 (N_7381,N_4803,N_4576);
and U7382 (N_7382,N_5247,N_5599);
xnor U7383 (N_7383,N_5360,N_4962);
or U7384 (N_7384,N_5134,N_4789);
nor U7385 (N_7385,N_4917,N_5900);
and U7386 (N_7386,N_4552,N_5662);
nor U7387 (N_7387,N_4875,N_5376);
or U7388 (N_7388,N_5652,N_5571);
nand U7389 (N_7389,N_5194,N_5510);
or U7390 (N_7390,N_5881,N_5180);
and U7391 (N_7391,N_5310,N_4787);
nor U7392 (N_7392,N_5772,N_5648);
nor U7393 (N_7393,N_5603,N_5914);
nor U7394 (N_7394,N_4987,N_5539);
nand U7395 (N_7395,N_5954,N_4546);
or U7396 (N_7396,N_5745,N_5846);
and U7397 (N_7397,N_5965,N_4595);
or U7398 (N_7398,N_4783,N_5702);
or U7399 (N_7399,N_5373,N_5191);
and U7400 (N_7400,N_5212,N_5775);
and U7401 (N_7401,N_5896,N_5141);
xnor U7402 (N_7402,N_4767,N_5357);
and U7403 (N_7403,N_4511,N_4733);
and U7404 (N_7404,N_5451,N_5656);
nor U7405 (N_7405,N_5407,N_5141);
and U7406 (N_7406,N_5319,N_5479);
xor U7407 (N_7407,N_5421,N_5994);
nand U7408 (N_7408,N_4729,N_4684);
and U7409 (N_7409,N_4825,N_5350);
and U7410 (N_7410,N_4932,N_5742);
nand U7411 (N_7411,N_4503,N_4677);
and U7412 (N_7412,N_5322,N_5089);
or U7413 (N_7413,N_5119,N_5405);
xor U7414 (N_7414,N_5319,N_4591);
or U7415 (N_7415,N_4822,N_5018);
and U7416 (N_7416,N_5523,N_5929);
nor U7417 (N_7417,N_5935,N_5226);
and U7418 (N_7418,N_5749,N_5176);
and U7419 (N_7419,N_5954,N_5032);
nor U7420 (N_7420,N_4703,N_5001);
and U7421 (N_7421,N_4759,N_5518);
nand U7422 (N_7422,N_4739,N_5374);
and U7423 (N_7423,N_5733,N_5591);
nand U7424 (N_7424,N_4881,N_5209);
or U7425 (N_7425,N_4815,N_5296);
or U7426 (N_7426,N_4551,N_5409);
and U7427 (N_7427,N_5429,N_5427);
nor U7428 (N_7428,N_5918,N_5246);
nand U7429 (N_7429,N_5901,N_4780);
and U7430 (N_7430,N_5388,N_4870);
or U7431 (N_7431,N_4549,N_5719);
nand U7432 (N_7432,N_5437,N_5104);
or U7433 (N_7433,N_4504,N_5567);
and U7434 (N_7434,N_5524,N_5560);
nand U7435 (N_7435,N_5688,N_5017);
and U7436 (N_7436,N_4669,N_5649);
or U7437 (N_7437,N_4697,N_5629);
or U7438 (N_7438,N_5440,N_5475);
nor U7439 (N_7439,N_5631,N_5882);
nor U7440 (N_7440,N_5279,N_5940);
or U7441 (N_7441,N_5813,N_5474);
and U7442 (N_7442,N_5931,N_4657);
nand U7443 (N_7443,N_5235,N_4749);
and U7444 (N_7444,N_5131,N_5138);
nor U7445 (N_7445,N_5268,N_5829);
xnor U7446 (N_7446,N_5454,N_5159);
xnor U7447 (N_7447,N_5236,N_5654);
or U7448 (N_7448,N_5568,N_5324);
nand U7449 (N_7449,N_5820,N_5185);
xor U7450 (N_7450,N_5609,N_5513);
nand U7451 (N_7451,N_5078,N_4581);
nand U7452 (N_7452,N_5857,N_4802);
nand U7453 (N_7453,N_5612,N_5857);
and U7454 (N_7454,N_4510,N_5674);
or U7455 (N_7455,N_4573,N_5932);
and U7456 (N_7456,N_5859,N_4981);
or U7457 (N_7457,N_5699,N_4530);
nand U7458 (N_7458,N_5649,N_4791);
nand U7459 (N_7459,N_5757,N_5666);
or U7460 (N_7460,N_4551,N_4666);
xnor U7461 (N_7461,N_5862,N_4898);
and U7462 (N_7462,N_5725,N_5418);
nor U7463 (N_7463,N_5312,N_5686);
and U7464 (N_7464,N_4690,N_5913);
or U7465 (N_7465,N_4813,N_4811);
or U7466 (N_7466,N_4610,N_5925);
nand U7467 (N_7467,N_5101,N_4888);
nand U7468 (N_7468,N_4729,N_5814);
and U7469 (N_7469,N_4638,N_5575);
nand U7470 (N_7470,N_5055,N_4874);
and U7471 (N_7471,N_4679,N_5286);
and U7472 (N_7472,N_4978,N_5429);
or U7473 (N_7473,N_5799,N_5739);
nand U7474 (N_7474,N_5269,N_5368);
nor U7475 (N_7475,N_5966,N_5166);
nand U7476 (N_7476,N_5839,N_5101);
and U7477 (N_7477,N_4535,N_4898);
or U7478 (N_7478,N_4534,N_4740);
nor U7479 (N_7479,N_5001,N_5589);
nor U7480 (N_7480,N_5541,N_5984);
or U7481 (N_7481,N_4935,N_5556);
nor U7482 (N_7482,N_5983,N_5242);
nor U7483 (N_7483,N_5154,N_4554);
and U7484 (N_7484,N_5118,N_5113);
nor U7485 (N_7485,N_4803,N_5949);
or U7486 (N_7486,N_5976,N_5351);
nand U7487 (N_7487,N_5997,N_5309);
or U7488 (N_7488,N_5946,N_5153);
nor U7489 (N_7489,N_5726,N_4751);
xnor U7490 (N_7490,N_5567,N_4631);
nor U7491 (N_7491,N_5129,N_5705);
xnor U7492 (N_7492,N_4617,N_4569);
or U7493 (N_7493,N_5524,N_5362);
or U7494 (N_7494,N_5470,N_4693);
nand U7495 (N_7495,N_5484,N_4827);
xor U7496 (N_7496,N_5114,N_5220);
nand U7497 (N_7497,N_5426,N_5233);
nor U7498 (N_7498,N_4825,N_4993);
nor U7499 (N_7499,N_5651,N_4599);
or U7500 (N_7500,N_6329,N_6445);
nand U7501 (N_7501,N_6858,N_7438);
or U7502 (N_7502,N_7033,N_7404);
or U7503 (N_7503,N_6010,N_6394);
nor U7504 (N_7504,N_7274,N_6426);
and U7505 (N_7505,N_7419,N_6285);
nor U7506 (N_7506,N_7170,N_7396);
or U7507 (N_7507,N_7020,N_6692);
nor U7508 (N_7508,N_6875,N_7144);
nor U7509 (N_7509,N_6530,N_6458);
or U7510 (N_7510,N_7473,N_7221);
or U7511 (N_7511,N_7158,N_6415);
or U7512 (N_7512,N_6772,N_6263);
nand U7513 (N_7513,N_6702,N_7231);
and U7514 (N_7514,N_6178,N_6521);
xor U7515 (N_7515,N_6909,N_7393);
and U7516 (N_7516,N_7389,N_7101);
nor U7517 (N_7517,N_6659,N_7282);
nand U7518 (N_7518,N_6412,N_6274);
and U7519 (N_7519,N_6999,N_7115);
xnor U7520 (N_7520,N_6436,N_6947);
nand U7521 (N_7521,N_7229,N_7093);
nor U7522 (N_7522,N_6712,N_7041);
nand U7523 (N_7523,N_6163,N_6155);
nor U7524 (N_7524,N_7222,N_6189);
nor U7525 (N_7525,N_6810,N_6213);
nand U7526 (N_7526,N_7278,N_6481);
and U7527 (N_7527,N_6462,N_6707);
or U7528 (N_7528,N_6492,N_6850);
nand U7529 (N_7529,N_6349,N_6432);
or U7530 (N_7530,N_6759,N_6691);
nor U7531 (N_7531,N_7228,N_7431);
and U7532 (N_7532,N_6278,N_6228);
or U7533 (N_7533,N_7450,N_6761);
nand U7534 (N_7534,N_7487,N_7434);
nand U7535 (N_7535,N_6007,N_7053);
nor U7536 (N_7536,N_6685,N_7296);
and U7537 (N_7537,N_6244,N_6879);
or U7538 (N_7538,N_7232,N_7277);
or U7539 (N_7539,N_7412,N_6853);
nor U7540 (N_7540,N_6419,N_6201);
nand U7541 (N_7541,N_7360,N_7363);
or U7542 (N_7542,N_6636,N_6245);
nand U7543 (N_7543,N_7411,N_6605);
nand U7544 (N_7544,N_6096,N_6929);
nand U7545 (N_7545,N_6127,N_6825);
or U7546 (N_7546,N_6912,N_7392);
or U7547 (N_7547,N_7209,N_6491);
nand U7548 (N_7548,N_6723,N_7433);
xor U7549 (N_7549,N_6341,N_7082);
nor U7550 (N_7550,N_6113,N_6047);
nor U7551 (N_7551,N_6260,N_6430);
or U7552 (N_7552,N_6865,N_7356);
and U7553 (N_7553,N_6477,N_7202);
nand U7554 (N_7554,N_6955,N_7361);
and U7555 (N_7555,N_6240,N_6054);
or U7556 (N_7556,N_6264,N_6828);
nand U7557 (N_7557,N_6364,N_7444);
or U7558 (N_7558,N_6622,N_7315);
or U7559 (N_7559,N_6747,N_6442);
nor U7560 (N_7560,N_6627,N_7013);
nor U7561 (N_7561,N_6936,N_7416);
nor U7562 (N_7562,N_7448,N_6755);
and U7563 (N_7563,N_6934,N_7080);
and U7564 (N_7564,N_6181,N_6610);
nor U7565 (N_7565,N_6156,N_7178);
and U7566 (N_7566,N_6433,N_6558);
or U7567 (N_7567,N_7173,N_6637);
nand U7568 (N_7568,N_7475,N_6289);
nor U7569 (N_7569,N_7340,N_7186);
and U7570 (N_7570,N_7104,N_6124);
nor U7571 (N_7571,N_7148,N_7255);
and U7572 (N_7572,N_7204,N_6764);
and U7573 (N_7573,N_7388,N_6733);
and U7574 (N_7574,N_6215,N_6315);
or U7575 (N_7575,N_6719,N_6452);
nor U7576 (N_7576,N_6515,N_6149);
and U7577 (N_7577,N_7391,N_7370);
or U7578 (N_7578,N_6634,N_6486);
or U7579 (N_7579,N_6983,N_7409);
and U7580 (N_7580,N_6107,N_6261);
xnor U7581 (N_7581,N_7208,N_7156);
nand U7582 (N_7582,N_6055,N_6065);
nand U7583 (N_7583,N_7225,N_6669);
or U7584 (N_7584,N_6505,N_6922);
nor U7585 (N_7585,N_6941,N_6042);
nor U7586 (N_7586,N_7309,N_6701);
and U7587 (N_7587,N_6930,N_6147);
nor U7588 (N_7588,N_7179,N_6926);
nand U7589 (N_7589,N_7423,N_6802);
nor U7590 (N_7590,N_6880,N_6737);
and U7591 (N_7591,N_7332,N_6358);
and U7592 (N_7592,N_6200,N_7061);
nor U7593 (N_7593,N_6087,N_6104);
nor U7594 (N_7594,N_6205,N_7004);
or U7595 (N_7595,N_6496,N_6129);
nand U7596 (N_7596,N_6237,N_6175);
nor U7597 (N_7597,N_7137,N_6574);
and U7598 (N_7598,N_6561,N_6824);
or U7599 (N_7599,N_6427,N_6736);
xnor U7600 (N_7600,N_6949,N_6567);
nand U7601 (N_7601,N_6569,N_6478);
or U7602 (N_7602,N_7323,N_6413);
or U7603 (N_7603,N_7055,N_6956);
xor U7604 (N_7604,N_6467,N_6134);
xor U7605 (N_7605,N_6520,N_7031);
and U7606 (N_7606,N_7493,N_6804);
nand U7607 (N_7607,N_7210,N_6450);
xnor U7608 (N_7608,N_6706,N_6119);
or U7609 (N_7609,N_6892,N_7424);
xnor U7610 (N_7610,N_7163,N_6214);
and U7611 (N_7611,N_6722,N_7374);
nand U7612 (N_7612,N_6439,N_7140);
or U7613 (N_7613,N_6663,N_7422);
nand U7614 (N_7614,N_6958,N_7083);
nor U7615 (N_7615,N_6601,N_6696);
nor U7616 (N_7616,N_6385,N_6783);
nand U7617 (N_7617,N_7369,N_6826);
or U7618 (N_7618,N_6033,N_6500);
nand U7619 (N_7619,N_7014,N_6283);
nor U7620 (N_7620,N_6233,N_7086);
or U7621 (N_7621,N_6395,N_7220);
and U7622 (N_7622,N_7284,N_6079);
xnor U7623 (N_7623,N_6552,N_7472);
and U7624 (N_7624,N_6018,N_6418);
nor U7625 (N_7625,N_6877,N_7136);
or U7626 (N_7626,N_7261,N_7286);
nor U7627 (N_7627,N_7152,N_6356);
nand U7628 (N_7628,N_6580,N_6020);
nand U7629 (N_7629,N_6326,N_7149);
and U7630 (N_7630,N_6317,N_6230);
or U7631 (N_7631,N_6917,N_7212);
nand U7632 (N_7632,N_6840,N_7070);
or U7633 (N_7633,N_7197,N_6465);
nand U7634 (N_7634,N_6710,N_6307);
or U7635 (N_7635,N_6793,N_7474);
nor U7636 (N_7636,N_6689,N_6378);
and U7637 (N_7637,N_7485,N_6342);
nand U7638 (N_7638,N_6940,N_6298);
nor U7639 (N_7639,N_7265,N_6564);
nor U7640 (N_7640,N_6039,N_6453);
or U7641 (N_7641,N_6968,N_6391);
nor U7642 (N_7642,N_7239,N_6805);
or U7643 (N_7643,N_6670,N_7036);
or U7644 (N_7644,N_7470,N_6286);
nor U7645 (N_7645,N_6219,N_7216);
nand U7646 (N_7646,N_6197,N_7154);
and U7647 (N_7647,N_7445,N_6115);
nand U7648 (N_7648,N_6734,N_6075);
and U7649 (N_7649,N_6776,N_6015);
and U7650 (N_7650,N_7451,N_6125);
and U7651 (N_7651,N_6464,N_6526);
nand U7652 (N_7652,N_6550,N_6003);
and U7653 (N_7653,N_6517,N_7313);
xor U7654 (N_7654,N_7258,N_7453);
nand U7655 (N_7655,N_6847,N_6856);
and U7656 (N_7656,N_6456,N_7354);
nor U7657 (N_7657,N_7380,N_7100);
xnor U7658 (N_7658,N_7483,N_6203);
nor U7659 (N_7659,N_7147,N_6475);
and U7660 (N_7660,N_6488,N_6678);
nor U7661 (N_7661,N_6661,N_6998);
and U7662 (N_7662,N_6004,N_7234);
or U7663 (N_7663,N_7106,N_6231);
nand U7664 (N_7664,N_6906,N_7131);
and U7665 (N_7665,N_7290,N_7000);
or U7666 (N_7666,N_6294,N_6209);
or U7667 (N_7667,N_6221,N_7406);
or U7668 (N_7668,N_7492,N_7250);
and U7669 (N_7669,N_6619,N_6608);
xor U7670 (N_7670,N_7058,N_6292);
nand U7671 (N_7671,N_6861,N_7015);
nand U7672 (N_7672,N_7165,N_6752);
and U7673 (N_7673,N_7200,N_7477);
nor U7674 (N_7674,N_6891,N_6184);
or U7675 (N_7675,N_6153,N_7312);
nor U7676 (N_7676,N_6139,N_7267);
nor U7677 (N_7677,N_6207,N_7130);
and U7678 (N_7678,N_6196,N_6613);
or U7679 (N_7679,N_6083,N_6076);
nor U7680 (N_7680,N_6218,N_7349);
nand U7681 (N_7681,N_6206,N_7443);
and U7682 (N_7682,N_6437,N_7337);
nor U7683 (N_7683,N_6652,N_6551);
or U7684 (N_7684,N_6651,N_6604);
and U7685 (N_7685,N_6609,N_7213);
nand U7686 (N_7686,N_6069,N_7325);
or U7687 (N_7687,N_7283,N_6832);
and U7688 (N_7688,N_6674,N_7377);
nand U7689 (N_7689,N_6893,N_6760);
or U7690 (N_7690,N_7072,N_7375);
nand U7691 (N_7691,N_6607,N_7496);
nand U7692 (N_7692,N_6813,N_6643);
nor U7693 (N_7693,N_6672,N_7045);
or U7694 (N_7694,N_6962,N_6518);
and U7695 (N_7695,N_7460,N_7383);
and U7696 (N_7696,N_6165,N_6954);
xnor U7697 (N_7697,N_6910,N_6984);
xor U7698 (N_7698,N_6715,N_6351);
or U7699 (N_7699,N_6562,N_6186);
nor U7700 (N_7700,N_6781,N_6255);
nor U7701 (N_7701,N_7345,N_6754);
nor U7702 (N_7702,N_6835,N_7078);
and U7703 (N_7703,N_6368,N_6448);
nor U7704 (N_7704,N_7357,N_7010);
or U7705 (N_7705,N_6291,N_7067);
nor U7706 (N_7706,N_6660,N_7171);
nand U7707 (N_7707,N_7027,N_6673);
and U7708 (N_7708,N_6367,N_6318);
nand U7709 (N_7709,N_6690,N_6644);
or U7710 (N_7710,N_6822,N_6818);
and U7711 (N_7711,N_6282,N_7488);
and U7712 (N_7712,N_6797,N_7064);
and U7713 (N_7713,N_6100,N_6814);
nor U7714 (N_7714,N_6675,N_6820);
nor U7715 (N_7715,N_6277,N_6347);
xnor U7716 (N_7716,N_6308,N_6050);
and U7717 (N_7717,N_7056,N_6746);
or U7718 (N_7718,N_7246,N_6483);
nand U7719 (N_7719,N_6924,N_6421);
or U7720 (N_7720,N_7074,N_7235);
nor U7721 (N_7721,N_6350,N_7217);
and U7722 (N_7722,N_6111,N_6067);
nor U7723 (N_7723,N_7214,N_7047);
and U7724 (N_7724,N_6641,N_6498);
or U7725 (N_7725,N_6290,N_7457);
and U7726 (N_7726,N_6740,N_6322);
or U7727 (N_7727,N_6943,N_6928);
or U7728 (N_7728,N_7301,N_7128);
nand U7729 (N_7729,N_6687,N_7017);
nor U7730 (N_7730,N_6995,N_6226);
and U7731 (N_7731,N_6611,N_7317);
xnor U7732 (N_7732,N_7043,N_7242);
and U7733 (N_7733,N_6435,N_6332);
nor U7734 (N_7734,N_6679,N_6023);
nand U7735 (N_7735,N_7414,N_7376);
and U7736 (N_7736,N_6183,N_6868);
or U7737 (N_7737,N_6829,N_6117);
xor U7738 (N_7738,N_6172,N_6470);
or U7739 (N_7739,N_6757,N_6988);
nand U7740 (N_7740,N_6198,N_6946);
or U7741 (N_7741,N_6568,N_7300);
or U7742 (N_7742,N_6573,N_6137);
nand U7743 (N_7743,N_7440,N_6393);
nand U7744 (N_7744,N_7168,N_6036);
or U7745 (N_7745,N_7049,N_6204);
nand U7746 (N_7746,N_6589,N_7009);
nor U7747 (N_7747,N_6894,N_7192);
nor U7748 (N_7748,N_6586,N_7237);
or U7749 (N_7749,N_7191,N_6416);
nand U7750 (N_7750,N_7211,N_7099);
and U7751 (N_7751,N_6900,N_6774);
nand U7752 (N_7752,N_6817,N_6380);
nand U7753 (N_7753,N_6045,N_6299);
nor U7754 (N_7754,N_7341,N_6990);
and U7755 (N_7755,N_7159,N_6362);
nor U7756 (N_7756,N_6677,N_7395);
nand U7757 (N_7757,N_6638,N_7441);
xnor U7758 (N_7758,N_6720,N_7199);
nand U7759 (N_7759,N_7150,N_6250);
xnor U7760 (N_7760,N_6400,N_7001);
or U7761 (N_7761,N_6417,N_6058);
nand U7762 (N_7762,N_6281,N_6987);
and U7763 (N_7763,N_7166,N_6844);
xnor U7764 (N_7764,N_7198,N_6913);
nand U7765 (N_7765,N_7307,N_7127);
or U7766 (N_7766,N_6485,N_7111);
nor U7767 (N_7767,N_7418,N_6252);
nor U7768 (N_7768,N_6420,N_6506);
or U7769 (N_7769,N_6976,N_6503);
nand U7770 (N_7770,N_6837,N_7077);
nand U7771 (N_7771,N_7439,N_6208);
nand U7772 (N_7772,N_7091,N_6727);
nand U7773 (N_7773,N_6942,N_6938);
xnor U7774 (N_7774,N_6801,N_6376);
nand U7775 (N_7775,N_6251,N_6633);
nor U7776 (N_7776,N_7310,N_6616);
nand U7777 (N_7777,N_7461,N_6053);
nor U7778 (N_7778,N_6522,N_7069);
or U7779 (N_7779,N_6006,N_6310);
nand U7780 (N_7780,N_7291,N_7029);
and U7781 (N_7781,N_6105,N_7153);
nor U7782 (N_7782,N_6796,N_7138);
xor U7783 (N_7783,N_6901,N_6258);
nor U7784 (N_7784,N_6902,N_6484);
xor U7785 (N_7785,N_6262,N_6085);
nand U7786 (N_7786,N_7241,N_6920);
and U7787 (N_7787,N_7098,N_6787);
nor U7788 (N_7788,N_6533,N_7397);
and U7789 (N_7789,N_6345,N_6815);
nor U7790 (N_7790,N_7331,N_7121);
or U7791 (N_7791,N_7353,N_6867);
or U7792 (N_7792,N_7415,N_6549);
nor U7793 (N_7793,N_7366,N_6180);
nand U7794 (N_7794,N_7075,N_6753);
nor U7795 (N_7795,N_6973,N_7316);
nand U7796 (N_7796,N_6513,N_6431);
and U7797 (N_7797,N_6799,N_7203);
nor U7798 (N_7798,N_6883,N_6854);
nor U7799 (N_7799,N_6142,N_6528);
nand U7800 (N_7800,N_6676,N_6716);
or U7801 (N_7801,N_6092,N_6951);
nor U7802 (N_7802,N_7002,N_7481);
and U7803 (N_7803,N_6479,N_6583);
and U7804 (N_7804,N_7145,N_6664);
and U7805 (N_7805,N_6590,N_6306);
and U7806 (N_7806,N_7089,N_7103);
xnor U7807 (N_7807,N_6576,N_6164);
xnor U7808 (N_7808,N_7497,N_6236);
or U7809 (N_7809,N_6404,N_7062);
xor U7810 (N_7810,N_6771,N_6863);
nand U7811 (N_7811,N_6606,N_6831);
nand U7812 (N_7812,N_7046,N_7030);
nand U7813 (N_7813,N_7151,N_6642);
and U7814 (N_7814,N_6314,N_7458);
and U7815 (N_7815,N_7059,N_6238);
and U7816 (N_7816,N_6265,N_6494);
and U7817 (N_7817,N_6859,N_6786);
or U7818 (N_7818,N_7334,N_7037);
nor U7819 (N_7819,N_6031,N_6617);
or U7820 (N_7820,N_6195,N_7358);
or U7821 (N_7821,N_7355,N_6525);
or U7822 (N_7822,N_6584,N_7119);
or U7823 (N_7823,N_6749,N_6788);
xor U7824 (N_7824,N_7177,N_6108);
xor U7825 (N_7825,N_6037,N_6011);
or U7826 (N_7826,N_6009,N_6146);
or U7827 (N_7827,N_7328,N_6109);
or U7828 (N_7828,N_7379,N_6849);
xor U7829 (N_7829,N_7456,N_7215);
nor U7830 (N_7830,N_6560,N_6321);
or U7831 (N_7831,N_6680,N_6343);
nor U7832 (N_7832,N_6509,N_7096);
or U7833 (N_7833,N_6789,N_7126);
or U7834 (N_7834,N_6827,N_7245);
nand U7835 (N_7835,N_6013,N_7293);
and U7836 (N_7836,N_7436,N_7270);
and U7837 (N_7837,N_7134,N_7175);
xnor U7838 (N_7838,N_7048,N_7162);
nor U7839 (N_7839,N_7057,N_6460);
nor U7840 (N_7840,N_6846,N_6459);
xor U7841 (N_7841,N_6794,N_6425);
and U7842 (N_7842,N_7052,N_7187);
and U7843 (N_7843,N_6337,N_6192);
or U7844 (N_7844,N_7279,N_6199);
and U7845 (N_7845,N_6896,N_6571);
nor U7846 (N_7846,N_6592,N_6222);
and U7847 (N_7847,N_7188,N_6501);
xnor U7848 (N_7848,N_6565,N_6709);
nor U7849 (N_7849,N_7266,N_7303);
nand U7850 (N_7850,N_6945,N_6514);
nand U7851 (N_7851,N_7105,N_6148);
xor U7852 (N_7852,N_6235,N_6698);
nor U7853 (N_7853,N_7135,N_7275);
and U7854 (N_7854,N_7008,N_6961);
and U7855 (N_7855,N_6683,N_7367);
or U7856 (N_7856,N_6545,N_6708);
xnor U7857 (N_7857,N_6387,N_6792);
nand U7858 (N_7858,N_6296,N_7344);
or U7859 (N_7859,N_7176,N_6873);
and U7860 (N_7860,N_7318,N_7260);
xor U7861 (N_7861,N_6253,N_6171);
or U7862 (N_7862,N_6694,N_7011);
and U7863 (N_7863,N_6559,N_6414);
and U7864 (N_7864,N_7462,N_6741);
nor U7865 (N_7865,N_7452,N_7133);
or U7866 (N_7866,N_7343,N_6595);
nor U7867 (N_7867,N_6114,N_6798);
nand U7868 (N_7868,N_6102,N_6911);
nor U7869 (N_7869,N_6834,N_7063);
or U7870 (N_7870,N_6743,N_6331);
xnor U7871 (N_7871,N_6851,N_6327);
nor U7872 (N_7872,N_6950,N_7155);
nor U7873 (N_7873,N_6099,N_6081);
and U7874 (N_7874,N_6964,N_6038);
and U7875 (N_7875,N_6931,N_7003);
nor U7876 (N_7876,N_6908,N_6389);
nand U7877 (N_7877,N_6365,N_6889);
nand U7878 (N_7878,N_7464,N_6557);
nor U7879 (N_7879,N_7005,N_7182);
nor U7880 (N_7880,N_6572,N_6463);
nor U7881 (N_7881,N_6600,N_7193);
nand U7882 (N_7882,N_7259,N_7226);
xnor U7883 (N_7883,N_6110,N_6293);
or U7884 (N_7884,N_6493,N_6654);
or U7885 (N_7885,N_6088,N_7465);
nor U7886 (N_7886,N_7425,N_6202);
nor U7887 (N_7887,N_6048,N_6269);
nor U7888 (N_7888,N_6334,N_6193);
or U7889 (N_7889,N_7120,N_6980);
nor U7890 (N_7890,N_7421,N_6305);
and U7891 (N_7891,N_6800,N_7484);
nor U7892 (N_7892,N_7230,N_6136);
or U7893 (N_7893,N_6030,N_6126);
nor U7894 (N_7894,N_6027,N_6921);
or U7895 (N_7895,N_6591,N_7304);
and U7896 (N_7896,N_6937,N_6989);
nand U7897 (N_7897,N_6598,N_7160);
nand U7898 (N_7898,N_6457,N_6516);
xor U7899 (N_7899,N_6188,N_6537);
nand U7900 (N_7900,N_6275,N_6311);
or U7901 (N_7901,N_6991,N_6443);
xor U7902 (N_7902,N_7449,N_6071);
or U7903 (N_7903,N_7042,N_6735);
and U7904 (N_7904,N_6247,N_6978);
and U7905 (N_7905,N_6959,N_6535);
nor U7906 (N_7906,N_7482,N_7426);
nand U7907 (N_7907,N_6179,N_6090);
and U7908 (N_7908,N_6862,N_6823);
nor U7909 (N_7909,N_6790,N_6273);
or U7910 (N_7910,N_6451,N_6363);
nand U7911 (N_7911,N_6399,N_6684);
and U7912 (N_7912,N_6648,N_6532);
and U7913 (N_7913,N_7254,N_7066);
and U7914 (N_7914,N_7494,N_6848);
or U7915 (N_7915,N_7407,N_7342);
nand U7916 (N_7916,N_6512,N_7172);
nor U7917 (N_7917,N_6145,N_7142);
nand U7918 (N_7918,N_6700,N_6232);
nand U7919 (N_7919,N_6141,N_6768);
nor U7920 (N_7920,N_6975,N_6068);
nor U7921 (N_7921,N_6344,N_6070);
and U7922 (N_7922,N_6986,N_7026);
xor U7923 (N_7923,N_6403,N_7305);
and U7924 (N_7924,N_6507,N_6769);
or U7925 (N_7925,N_6182,N_6112);
xor U7926 (N_7926,N_6819,N_7139);
and U7927 (N_7927,N_6635,N_6878);
xor U7928 (N_7928,N_6185,N_6170);
nand U7929 (N_7929,N_7347,N_6061);
nor U7930 (N_7930,N_6581,N_6154);
or U7931 (N_7931,N_6072,N_6523);
xnor U7932 (N_7932,N_6836,N_7129);
and U7933 (N_7933,N_7073,N_6808);
nor U7934 (N_7934,N_6309,N_7194);
and U7935 (N_7935,N_6325,N_7382);
and U7936 (N_7936,N_6000,N_6080);
nand U7937 (N_7937,N_6150,N_6161);
and U7938 (N_7938,N_7195,N_6751);
nor U7939 (N_7939,N_6028,N_6135);
or U7940 (N_7940,N_6473,N_6021);
nand U7941 (N_7941,N_7403,N_6852);
and U7942 (N_7942,N_7264,N_7463);
nand U7943 (N_7943,N_6821,N_7044);
or U7944 (N_7944,N_7189,N_6718);
nand U7945 (N_7945,N_6194,N_6711);
or U7946 (N_7946,N_6773,N_6668);
nor U7947 (N_7947,N_7181,N_7320);
or U7948 (N_7948,N_6620,N_6035);
nor U7949 (N_7949,N_7206,N_7466);
or U7950 (N_7950,N_6686,N_6190);
nand U7951 (N_7951,N_6593,N_6907);
nor U7952 (N_7952,N_7132,N_7285);
or U7953 (N_7953,N_6739,N_6373);
nand U7954 (N_7954,N_7006,N_6248);
nor U7955 (N_7955,N_6952,N_6898);
or U7956 (N_7956,N_6122,N_6377);
nor U7957 (N_7957,N_6019,N_6131);
nor U7958 (N_7958,N_7102,N_7478);
and U7959 (N_7959,N_7196,N_6899);
and U7960 (N_7960,N_6704,N_6653);
nand U7961 (N_7961,N_6527,N_6697);
nand U7962 (N_7962,N_6548,N_6872);
nor U7963 (N_7963,N_7161,N_6953);
or U7964 (N_7964,N_6703,N_6220);
or U7965 (N_7965,N_7207,N_6257);
and U7966 (N_7966,N_7125,N_7427);
nand U7967 (N_7967,N_7372,N_6128);
nand U7968 (N_7968,N_6024,N_7302);
nor U7969 (N_7969,N_6531,N_7299);
xor U7970 (N_7970,N_6303,N_6052);
nor U7971 (N_7971,N_6402,N_7384);
or U7972 (N_7972,N_6650,N_7107);
and U7973 (N_7973,N_7034,N_6353);
nand U7974 (N_7974,N_6120,N_6504);
and U7975 (N_7975,N_6324,N_6313);
nand U7976 (N_7976,N_7257,N_7447);
and U7977 (N_7977,N_6992,N_7373);
nand U7978 (N_7978,N_6688,N_6816);
or U7979 (N_7979,N_6916,N_7420);
nand U7980 (N_7980,N_7248,N_7253);
or U7981 (N_7981,N_7114,N_6603);
nand U7982 (N_7982,N_6089,N_7365);
nand U7983 (N_7983,N_7294,N_6063);
and U7984 (N_7984,N_6588,N_6138);
nor U7985 (N_7985,N_6162,N_6328);
nor U7986 (N_7986,N_6046,N_7321);
nor U7987 (N_7987,N_6979,N_6434);
and U7988 (N_7988,N_6267,N_6428);
nand U7989 (N_7989,N_6152,N_7455);
or U7990 (N_7990,N_6167,N_6140);
or U7991 (N_7991,N_6887,N_7146);
nor U7992 (N_7992,N_6422,N_6682);
nand U7993 (N_7993,N_6499,N_7486);
and U7994 (N_7994,N_6410,N_7085);
xnor U7995 (N_7995,N_6996,N_7124);
xor U7996 (N_7996,N_6628,N_7019);
nand U7997 (N_7997,N_6730,N_6631);
nor U7998 (N_7998,N_7401,N_6423);
nand U7999 (N_7999,N_6782,N_6933);
xor U8000 (N_8000,N_6779,N_6316);
and U8001 (N_8001,N_7028,N_6246);
nor U8002 (N_8002,N_7256,N_6838);
nor U8003 (N_8003,N_6927,N_6217);
and U8004 (N_8004,N_6582,N_6330);
nand U8005 (N_8005,N_6312,N_6963);
xnor U8006 (N_8006,N_6374,N_6870);
nor U8007 (N_8007,N_7118,N_6919);
xnor U8008 (N_8008,N_7022,N_6855);
nand U8009 (N_8009,N_7288,N_7157);
or U8010 (N_8010,N_6173,N_6623);
and U8011 (N_8011,N_6519,N_7233);
nand U8012 (N_8012,N_6304,N_6082);
nor U8013 (N_8013,N_6807,N_7092);
nand U8014 (N_8014,N_7308,N_6508);
nand U8015 (N_8015,N_6287,N_6939);
nor U8016 (N_8016,N_6158,N_6438);
xnor U8017 (N_8017,N_6784,N_7292);
and U8018 (N_8018,N_6297,N_6091);
nor U8019 (N_8019,N_7035,N_7183);
nand U8020 (N_8020,N_6409,N_6918);
and U8021 (N_8021,N_6534,N_6666);
or U8022 (N_8022,N_6511,N_7263);
nand U8023 (N_8023,N_6812,N_6001);
or U8024 (N_8024,N_6064,N_6276);
and U8025 (N_8025,N_6721,N_6357);
nor U8026 (N_8026,N_7330,N_6594);
nand U8027 (N_8027,N_6765,N_7095);
or U8028 (N_8028,N_7499,N_6890);
and U8029 (N_8029,N_6775,N_6597);
or U8030 (N_8030,N_6002,N_6016);
nor U8031 (N_8031,N_6225,N_6914);
xor U8032 (N_8032,N_6270,N_7327);
and U8033 (N_8033,N_6383,N_6480);
or U8034 (N_8034,N_6602,N_7467);
nor U8035 (N_8035,N_7432,N_6541);
nand U8036 (N_8036,N_7410,N_6869);
nand U8037 (N_8037,N_6843,N_7262);
or U8038 (N_8038,N_7417,N_6407);
nor U8039 (N_8039,N_7480,N_7319);
or U8040 (N_8040,N_7268,N_7068);
nor U8041 (N_8041,N_6960,N_6970);
nand U8042 (N_8042,N_6585,N_6490);
xnor U8043 (N_8043,N_6043,N_7295);
or U8044 (N_8044,N_6626,N_6615);
nor U8045 (N_8045,N_7280,N_7251);
and U8046 (N_8046,N_7227,N_6806);
nand U8047 (N_8047,N_6731,N_7038);
nand U8048 (N_8048,N_6352,N_6717);
nor U8049 (N_8049,N_7180,N_6886);
nand U8050 (N_8050,N_6355,N_6529);
nand U8051 (N_8051,N_6791,N_6166);
and U8052 (N_8052,N_7169,N_7289);
nor U8053 (N_8053,N_6948,N_7476);
nor U8054 (N_8054,N_6044,N_6049);
or U8055 (N_8055,N_6742,N_6524);
nand U8056 (N_8056,N_7117,N_6424);
nor U8057 (N_8057,N_6130,N_6646);
and U8058 (N_8058,N_6234,N_6563);
nor U8059 (N_8059,N_6177,N_6441);
xor U8060 (N_8060,N_6728,N_6339);
or U8061 (N_8061,N_6360,N_6745);
nor U8062 (N_8062,N_6553,N_6369);
nor U8063 (N_8063,N_7339,N_6766);
nand U8064 (N_8064,N_6510,N_6780);
or U8065 (N_8065,N_6408,N_7348);
nor U8066 (N_8066,N_6216,N_6903);
or U8067 (N_8067,N_6026,N_7468);
nor U8068 (N_8068,N_6471,N_6864);
or U8069 (N_8069,N_6693,N_6833);
nor U8070 (N_8070,N_6025,N_6017);
or U8071 (N_8071,N_6372,N_6965);
and U8072 (N_8072,N_7371,N_6570);
nor U8073 (N_8073,N_7405,N_6132);
and U8074 (N_8074,N_6073,N_6060);
or U8075 (N_8075,N_6397,N_7032);
or U8076 (N_8076,N_7112,N_6323);
nand U8077 (N_8077,N_6884,N_6078);
and U8078 (N_8078,N_7122,N_7065);
nor U8079 (N_8079,N_7273,N_6981);
and U8080 (N_8080,N_6041,N_7495);
and U8081 (N_8081,N_6461,N_6012);
xnor U8082 (N_8082,N_6366,N_6106);
nor U8083 (N_8083,N_7324,N_7223);
or U8084 (N_8084,N_6778,N_6371);
or U8085 (N_8085,N_6904,N_6444);
nand U8086 (N_8086,N_6925,N_6699);
or U8087 (N_8087,N_6888,N_6575);
nor U8088 (N_8088,N_6333,N_6830);
xnor U8089 (N_8089,N_6390,N_6466);
and U8090 (N_8090,N_6982,N_7097);
nor U8091 (N_8091,N_7174,N_6577);
nor U8092 (N_8092,N_6762,N_6187);
and U8093 (N_8093,N_6587,N_6629);
or U8094 (N_8094,N_7333,N_7430);
xnor U8095 (N_8095,N_6487,N_7060);
nand U8096 (N_8096,N_6379,N_7113);
nor U8097 (N_8097,N_6502,N_6447);
xor U8098 (N_8098,N_7249,N_7071);
xor U8099 (N_8099,N_7094,N_7018);
and U8100 (N_8100,N_7116,N_7386);
nor U8101 (N_8101,N_6726,N_6476);
nand U8102 (N_8102,N_6118,N_6301);
or U8103 (N_8103,N_6384,N_7051);
nand U8104 (N_8104,N_6320,N_6094);
nor U8105 (N_8105,N_7269,N_7437);
and U8106 (N_8106,N_6489,N_7454);
or U8107 (N_8107,N_6667,N_7326);
nand U8108 (N_8108,N_6388,N_7336);
and U8109 (N_8109,N_6361,N_6280);
nor U8110 (N_8110,N_6845,N_7218);
or U8111 (N_8111,N_7398,N_6915);
and U8112 (N_8112,N_6621,N_6472);
or U8113 (N_8113,N_6544,N_6229);
or U8114 (N_8114,N_6546,N_6785);
nand U8115 (N_8115,N_7054,N_7385);
nand U8116 (N_8116,N_6168,N_6354);
nand U8117 (N_8117,N_7076,N_7399);
nand U8118 (N_8118,N_6985,N_7272);
nand U8119 (N_8119,N_7185,N_6335);
and U8120 (N_8120,N_6101,N_7297);
xor U8121 (N_8121,N_6429,N_6340);
or U8122 (N_8122,N_7446,N_6406);
nor U8123 (N_8123,N_7314,N_6116);
nand U8124 (N_8124,N_6121,N_7471);
nand U8125 (N_8125,N_6256,N_7362);
and U8126 (N_8126,N_6223,N_6066);
and U8127 (N_8127,N_6392,N_6866);
or U8128 (N_8128,N_6763,N_6935);
xnor U8129 (N_8129,N_7143,N_7024);
and U8130 (N_8130,N_7109,N_6243);
or U8131 (N_8131,N_7025,N_6645);
or U8132 (N_8132,N_6971,N_6239);
and U8133 (N_8133,N_6034,N_6614);
xor U8134 (N_8134,N_7252,N_7359);
and U8135 (N_8135,N_6098,N_7352);
xor U8136 (N_8136,N_7205,N_6649);
nor U8137 (N_8137,N_6860,N_6302);
nand U8138 (N_8138,N_6191,N_6640);
nand U8139 (N_8139,N_6446,N_7306);
nand U8140 (N_8140,N_6612,N_6336);
and U8141 (N_8141,N_6599,N_6618);
xor U8142 (N_8142,N_7039,N_7351);
and U8143 (N_8143,N_7408,N_7110);
or U8144 (N_8144,N_6750,N_6647);
nor U8145 (N_8145,N_6386,N_6536);
nor U8146 (N_8146,N_7081,N_7023);
nand U8147 (N_8147,N_6974,N_6625);
nor U8148 (N_8148,N_6871,N_6542);
and U8149 (N_8149,N_6074,N_6578);
or U8150 (N_8150,N_6174,N_6212);
and U8151 (N_8151,N_6022,N_6227);
nor U8152 (N_8152,N_6056,N_6295);
nand U8153 (N_8153,N_7123,N_6468);
xnor U8154 (N_8154,N_6695,N_6454);
nor U8155 (N_8155,N_7236,N_7364);
nand U8156 (N_8156,N_6540,N_6268);
nand U8157 (N_8157,N_6398,N_6469);
nor U8158 (N_8158,N_7442,N_6381);
and U8159 (N_8159,N_6271,N_6057);
nor U8160 (N_8160,N_6655,N_7090);
nor U8161 (N_8161,N_6639,N_7479);
xor U8162 (N_8162,N_6062,N_6396);
or U8163 (N_8163,N_6051,N_7243);
xnor U8164 (N_8164,N_6455,N_6596);
and U8165 (N_8165,N_7368,N_6905);
nand U8166 (N_8166,N_7381,N_6967);
or U8167 (N_8167,N_6732,N_6770);
and U8168 (N_8168,N_6997,N_6157);
nor U8169 (N_8169,N_6665,N_7276);
xor U8170 (N_8170,N_6969,N_6658);
nand U8171 (N_8171,N_6014,N_6482);
nand U8172 (N_8172,N_7298,N_7016);
and U8173 (N_8173,N_6839,N_7489);
nor U8174 (N_8174,N_6144,N_6210);
and U8175 (N_8175,N_7108,N_6169);
nor U8176 (N_8176,N_6032,N_7322);
xor U8177 (N_8177,N_6923,N_6103);
nand U8178 (N_8178,N_6440,N_6748);
nand U8179 (N_8179,N_7428,N_7164);
nor U8180 (N_8180,N_6547,N_7394);
xor U8181 (N_8181,N_7141,N_7167);
nor U8182 (N_8182,N_6972,N_6632);
xnor U8183 (N_8183,N_7190,N_6671);
nor U8184 (N_8184,N_6005,N_6795);
nor U8185 (N_8185,N_7184,N_7287);
or U8186 (N_8186,N_7079,N_6857);
or U8187 (N_8187,N_7335,N_6008);
or U8188 (N_8188,N_6249,N_6449);
and U8189 (N_8189,N_6405,N_6957);
xnor U8190 (N_8190,N_7238,N_6885);
or U8191 (N_8191,N_6259,N_6077);
nor U8192 (N_8192,N_7271,N_6411);
and U8193 (N_8193,N_6370,N_6348);
nand U8194 (N_8194,N_6375,N_6876);
and U8195 (N_8195,N_7490,N_6882);
or U8196 (N_8196,N_6543,N_7402);
nand U8197 (N_8197,N_6809,N_6359);
and U8198 (N_8198,N_6086,N_6159);
nor U8199 (N_8199,N_7201,N_7390);
nand U8200 (N_8200,N_7040,N_6133);
nand U8201 (N_8201,N_6284,N_6738);
nor U8202 (N_8202,N_6811,N_7469);
or U8203 (N_8203,N_6040,N_6059);
nand U8204 (N_8204,N_6497,N_7346);
or U8205 (N_8205,N_6176,N_6554);
or U8206 (N_8206,N_6993,N_7329);
nand U8207 (N_8207,N_6657,N_6725);
or U8208 (N_8208,N_6160,N_7387);
or U8209 (N_8209,N_6744,N_7413);
or U8210 (N_8210,N_7491,N_6241);
xnor U8211 (N_8211,N_6338,N_7219);
nand U8212 (N_8212,N_6994,N_6842);
or U8213 (N_8213,N_6279,N_6143);
or U8214 (N_8214,N_6495,N_6539);
or U8215 (N_8215,N_7311,N_6288);
and U8216 (N_8216,N_7459,N_7084);
and U8217 (N_8217,N_6756,N_6346);
and U8218 (N_8218,N_7050,N_6084);
nor U8219 (N_8219,N_6401,N_6724);
or U8220 (N_8220,N_6211,N_6254);
or U8221 (N_8221,N_6681,N_6729);
nand U8222 (N_8222,N_7435,N_7021);
nor U8223 (N_8223,N_6966,N_6758);
xor U8224 (N_8224,N_7007,N_6272);
nor U8225 (N_8225,N_6932,N_6777);
and U8226 (N_8226,N_6266,N_6895);
and U8227 (N_8227,N_7429,N_7378);
nand U8228 (N_8228,N_7350,N_6566);
or U8229 (N_8229,N_6097,N_6713);
or U8230 (N_8230,N_6897,N_7498);
or U8231 (N_8231,N_6319,N_6095);
and U8232 (N_8232,N_7224,N_7338);
nor U8233 (N_8233,N_6093,N_6714);
nand U8234 (N_8234,N_6123,N_7087);
nor U8235 (N_8235,N_7240,N_6662);
or U8236 (N_8236,N_7088,N_6944);
or U8237 (N_8237,N_6630,N_6300);
and U8238 (N_8238,N_6881,N_6841);
nor U8239 (N_8239,N_7012,N_6538);
and U8240 (N_8240,N_6803,N_6555);
and U8241 (N_8241,N_7400,N_6656);
nor U8242 (N_8242,N_6224,N_6382);
xnor U8243 (N_8243,N_6977,N_6874);
or U8244 (N_8244,N_6556,N_6151);
and U8245 (N_8245,N_7281,N_6767);
and U8246 (N_8246,N_6705,N_6474);
nor U8247 (N_8247,N_7244,N_7247);
xor U8248 (N_8248,N_6029,N_6579);
xnor U8249 (N_8249,N_6242,N_6624);
and U8250 (N_8250,N_6978,N_6202);
or U8251 (N_8251,N_6472,N_6352);
and U8252 (N_8252,N_6099,N_6527);
and U8253 (N_8253,N_6284,N_7338);
nor U8254 (N_8254,N_6842,N_7137);
or U8255 (N_8255,N_6257,N_6913);
or U8256 (N_8256,N_6973,N_6046);
or U8257 (N_8257,N_6057,N_6061);
nor U8258 (N_8258,N_7156,N_6548);
and U8259 (N_8259,N_6574,N_6304);
and U8260 (N_8260,N_6701,N_6395);
xnor U8261 (N_8261,N_7377,N_6893);
xnor U8262 (N_8262,N_6682,N_7397);
and U8263 (N_8263,N_6331,N_6259);
and U8264 (N_8264,N_6816,N_7008);
xnor U8265 (N_8265,N_6330,N_7413);
xor U8266 (N_8266,N_6745,N_6093);
and U8267 (N_8267,N_6087,N_6054);
or U8268 (N_8268,N_7469,N_6181);
nor U8269 (N_8269,N_6926,N_7061);
nor U8270 (N_8270,N_7135,N_6206);
and U8271 (N_8271,N_6411,N_7360);
nand U8272 (N_8272,N_6161,N_6090);
nor U8273 (N_8273,N_6677,N_6313);
nor U8274 (N_8274,N_6445,N_6142);
and U8275 (N_8275,N_6071,N_6559);
nand U8276 (N_8276,N_7467,N_7449);
nand U8277 (N_8277,N_6290,N_7372);
and U8278 (N_8278,N_6202,N_6613);
and U8279 (N_8279,N_6006,N_6422);
nand U8280 (N_8280,N_7463,N_7262);
nand U8281 (N_8281,N_6942,N_7261);
nand U8282 (N_8282,N_6359,N_6556);
and U8283 (N_8283,N_6139,N_6466);
or U8284 (N_8284,N_6675,N_6328);
or U8285 (N_8285,N_7195,N_7141);
and U8286 (N_8286,N_7130,N_7206);
and U8287 (N_8287,N_6092,N_6273);
and U8288 (N_8288,N_6781,N_6705);
nand U8289 (N_8289,N_7441,N_6136);
and U8290 (N_8290,N_6726,N_6284);
nor U8291 (N_8291,N_6950,N_7040);
and U8292 (N_8292,N_6647,N_6815);
or U8293 (N_8293,N_6989,N_7050);
nor U8294 (N_8294,N_7388,N_7101);
and U8295 (N_8295,N_6132,N_7368);
and U8296 (N_8296,N_6902,N_7066);
and U8297 (N_8297,N_6859,N_6874);
nor U8298 (N_8298,N_6359,N_7163);
nor U8299 (N_8299,N_6880,N_6936);
or U8300 (N_8300,N_7422,N_6795);
nand U8301 (N_8301,N_6457,N_6429);
nor U8302 (N_8302,N_7362,N_7218);
and U8303 (N_8303,N_6502,N_7086);
and U8304 (N_8304,N_6177,N_6603);
nand U8305 (N_8305,N_6495,N_6537);
nand U8306 (N_8306,N_7347,N_6119);
xnor U8307 (N_8307,N_7124,N_7015);
nor U8308 (N_8308,N_6560,N_7043);
and U8309 (N_8309,N_7172,N_6066);
and U8310 (N_8310,N_6673,N_6939);
nand U8311 (N_8311,N_6925,N_6092);
nor U8312 (N_8312,N_6786,N_6500);
nand U8313 (N_8313,N_6814,N_6498);
and U8314 (N_8314,N_6657,N_7059);
and U8315 (N_8315,N_6563,N_7261);
or U8316 (N_8316,N_6743,N_6181);
and U8317 (N_8317,N_6847,N_7362);
nor U8318 (N_8318,N_6953,N_6879);
or U8319 (N_8319,N_6070,N_7159);
and U8320 (N_8320,N_6055,N_6613);
or U8321 (N_8321,N_6792,N_7103);
or U8322 (N_8322,N_7156,N_6264);
or U8323 (N_8323,N_7404,N_6921);
or U8324 (N_8324,N_6719,N_7179);
or U8325 (N_8325,N_6623,N_6330);
or U8326 (N_8326,N_6223,N_7495);
and U8327 (N_8327,N_7043,N_7258);
nand U8328 (N_8328,N_6897,N_7311);
and U8329 (N_8329,N_6743,N_7069);
and U8330 (N_8330,N_6766,N_7320);
nand U8331 (N_8331,N_6356,N_7383);
nor U8332 (N_8332,N_7178,N_6900);
nand U8333 (N_8333,N_6312,N_6423);
xor U8334 (N_8334,N_6147,N_7485);
or U8335 (N_8335,N_6143,N_7165);
nand U8336 (N_8336,N_6617,N_6890);
nand U8337 (N_8337,N_6145,N_7454);
nor U8338 (N_8338,N_7440,N_6547);
and U8339 (N_8339,N_7241,N_6939);
and U8340 (N_8340,N_6079,N_6922);
or U8341 (N_8341,N_6292,N_7230);
xor U8342 (N_8342,N_6096,N_6392);
nor U8343 (N_8343,N_6991,N_6024);
xnor U8344 (N_8344,N_7288,N_6605);
nor U8345 (N_8345,N_6335,N_7142);
nor U8346 (N_8346,N_6570,N_7262);
or U8347 (N_8347,N_6875,N_7090);
or U8348 (N_8348,N_6985,N_6576);
nor U8349 (N_8349,N_6480,N_6715);
nor U8350 (N_8350,N_6036,N_7442);
nor U8351 (N_8351,N_7436,N_6023);
nand U8352 (N_8352,N_6608,N_6848);
nand U8353 (N_8353,N_6852,N_6220);
or U8354 (N_8354,N_6710,N_6464);
and U8355 (N_8355,N_6522,N_7281);
xor U8356 (N_8356,N_6755,N_6012);
and U8357 (N_8357,N_7302,N_6868);
or U8358 (N_8358,N_6738,N_7104);
or U8359 (N_8359,N_7283,N_7488);
and U8360 (N_8360,N_6135,N_6023);
nand U8361 (N_8361,N_6237,N_7101);
and U8362 (N_8362,N_6103,N_6937);
nor U8363 (N_8363,N_7329,N_7413);
and U8364 (N_8364,N_6909,N_7030);
nand U8365 (N_8365,N_7414,N_6639);
or U8366 (N_8366,N_6004,N_6171);
and U8367 (N_8367,N_6277,N_6454);
nand U8368 (N_8368,N_7038,N_6531);
nand U8369 (N_8369,N_6848,N_6471);
nand U8370 (N_8370,N_7494,N_7288);
nand U8371 (N_8371,N_6508,N_7289);
and U8372 (N_8372,N_7119,N_6460);
and U8373 (N_8373,N_6061,N_6785);
or U8374 (N_8374,N_6969,N_6608);
and U8375 (N_8375,N_6292,N_6368);
xor U8376 (N_8376,N_6094,N_6245);
or U8377 (N_8377,N_7224,N_6810);
or U8378 (N_8378,N_6092,N_7039);
nand U8379 (N_8379,N_6679,N_6986);
nor U8380 (N_8380,N_6404,N_6862);
and U8381 (N_8381,N_6640,N_6768);
nor U8382 (N_8382,N_6810,N_7021);
and U8383 (N_8383,N_6912,N_6784);
nand U8384 (N_8384,N_6550,N_6175);
or U8385 (N_8385,N_7474,N_7111);
nor U8386 (N_8386,N_6764,N_7403);
or U8387 (N_8387,N_6305,N_7342);
and U8388 (N_8388,N_7117,N_6999);
nor U8389 (N_8389,N_6832,N_6095);
nand U8390 (N_8390,N_7250,N_6875);
nand U8391 (N_8391,N_6880,N_7071);
or U8392 (N_8392,N_7397,N_6506);
or U8393 (N_8393,N_7182,N_7404);
and U8394 (N_8394,N_7149,N_6294);
nand U8395 (N_8395,N_6843,N_6703);
and U8396 (N_8396,N_6066,N_6807);
or U8397 (N_8397,N_6660,N_7473);
nor U8398 (N_8398,N_7179,N_6996);
nand U8399 (N_8399,N_7123,N_7441);
nor U8400 (N_8400,N_6001,N_6856);
nor U8401 (N_8401,N_6728,N_6421);
and U8402 (N_8402,N_6410,N_6778);
nand U8403 (N_8403,N_7070,N_6521);
nand U8404 (N_8404,N_7363,N_6651);
or U8405 (N_8405,N_6352,N_7282);
nand U8406 (N_8406,N_6083,N_7042);
nand U8407 (N_8407,N_7368,N_6323);
nor U8408 (N_8408,N_6312,N_7154);
xor U8409 (N_8409,N_6424,N_6749);
or U8410 (N_8410,N_6665,N_6759);
nor U8411 (N_8411,N_7179,N_6075);
and U8412 (N_8412,N_7348,N_6838);
nand U8413 (N_8413,N_6986,N_6291);
and U8414 (N_8414,N_6464,N_6599);
or U8415 (N_8415,N_6957,N_7052);
and U8416 (N_8416,N_6122,N_6908);
nor U8417 (N_8417,N_7010,N_7324);
nand U8418 (N_8418,N_6978,N_6075);
nand U8419 (N_8419,N_6636,N_7170);
nand U8420 (N_8420,N_7316,N_6842);
nor U8421 (N_8421,N_7203,N_7482);
or U8422 (N_8422,N_6384,N_6601);
nand U8423 (N_8423,N_6959,N_6616);
nand U8424 (N_8424,N_6684,N_6002);
nand U8425 (N_8425,N_6082,N_6245);
and U8426 (N_8426,N_7275,N_7084);
nor U8427 (N_8427,N_7477,N_6738);
nor U8428 (N_8428,N_6500,N_6049);
nand U8429 (N_8429,N_6318,N_6636);
and U8430 (N_8430,N_6665,N_6920);
or U8431 (N_8431,N_6555,N_6649);
or U8432 (N_8432,N_6104,N_6396);
and U8433 (N_8433,N_6167,N_6752);
nor U8434 (N_8434,N_7360,N_6479);
or U8435 (N_8435,N_6028,N_6677);
nand U8436 (N_8436,N_6438,N_6243);
nor U8437 (N_8437,N_6523,N_6334);
or U8438 (N_8438,N_7058,N_6223);
nand U8439 (N_8439,N_6643,N_7143);
or U8440 (N_8440,N_6973,N_7019);
nand U8441 (N_8441,N_7439,N_6872);
or U8442 (N_8442,N_7239,N_7447);
nand U8443 (N_8443,N_6557,N_6859);
or U8444 (N_8444,N_7319,N_7368);
nor U8445 (N_8445,N_6943,N_7443);
nand U8446 (N_8446,N_7264,N_6843);
and U8447 (N_8447,N_6698,N_6524);
xor U8448 (N_8448,N_6382,N_7022);
nand U8449 (N_8449,N_6234,N_6996);
or U8450 (N_8450,N_6549,N_6077);
xnor U8451 (N_8451,N_7218,N_6115);
and U8452 (N_8452,N_7390,N_6423);
nor U8453 (N_8453,N_7462,N_6119);
nand U8454 (N_8454,N_6770,N_7462);
nand U8455 (N_8455,N_7247,N_6183);
and U8456 (N_8456,N_6828,N_7223);
or U8457 (N_8457,N_7449,N_7333);
xor U8458 (N_8458,N_6722,N_7438);
nor U8459 (N_8459,N_7370,N_6936);
and U8460 (N_8460,N_6631,N_6689);
nand U8461 (N_8461,N_6430,N_6790);
nand U8462 (N_8462,N_7214,N_6765);
or U8463 (N_8463,N_6898,N_6975);
and U8464 (N_8464,N_6937,N_7046);
nand U8465 (N_8465,N_6499,N_6447);
or U8466 (N_8466,N_6269,N_6635);
nand U8467 (N_8467,N_6523,N_7175);
or U8468 (N_8468,N_7027,N_6469);
or U8469 (N_8469,N_6085,N_6176);
or U8470 (N_8470,N_6970,N_6397);
nor U8471 (N_8471,N_6249,N_6996);
and U8472 (N_8472,N_7188,N_6540);
nand U8473 (N_8473,N_7275,N_6447);
nand U8474 (N_8474,N_7373,N_6819);
and U8475 (N_8475,N_6614,N_6583);
nor U8476 (N_8476,N_6569,N_7100);
and U8477 (N_8477,N_6380,N_6778);
and U8478 (N_8478,N_6082,N_6767);
xor U8479 (N_8479,N_6091,N_7012);
xor U8480 (N_8480,N_7486,N_7117);
xnor U8481 (N_8481,N_7201,N_7081);
or U8482 (N_8482,N_6770,N_6027);
nor U8483 (N_8483,N_7388,N_6611);
nand U8484 (N_8484,N_6683,N_7152);
and U8485 (N_8485,N_6435,N_7388);
and U8486 (N_8486,N_6306,N_7049);
and U8487 (N_8487,N_6694,N_6663);
or U8488 (N_8488,N_6559,N_7465);
or U8489 (N_8489,N_6625,N_6806);
or U8490 (N_8490,N_7225,N_7238);
nor U8491 (N_8491,N_6238,N_6030);
nand U8492 (N_8492,N_7247,N_6842);
xnor U8493 (N_8493,N_6325,N_6927);
nor U8494 (N_8494,N_6858,N_6992);
nand U8495 (N_8495,N_6951,N_7013);
nor U8496 (N_8496,N_6224,N_6141);
or U8497 (N_8497,N_6107,N_6234);
xnor U8498 (N_8498,N_7311,N_6214);
or U8499 (N_8499,N_7015,N_6594);
nor U8500 (N_8500,N_7325,N_6042);
nor U8501 (N_8501,N_7037,N_6267);
nor U8502 (N_8502,N_6084,N_6844);
nor U8503 (N_8503,N_6643,N_6268);
and U8504 (N_8504,N_6753,N_6186);
nand U8505 (N_8505,N_6487,N_6630);
nor U8506 (N_8506,N_6544,N_6903);
xnor U8507 (N_8507,N_6122,N_7080);
or U8508 (N_8508,N_7380,N_6812);
nor U8509 (N_8509,N_6539,N_6905);
xnor U8510 (N_8510,N_6793,N_6687);
nor U8511 (N_8511,N_6604,N_6477);
or U8512 (N_8512,N_6486,N_6814);
nor U8513 (N_8513,N_6449,N_7473);
or U8514 (N_8514,N_7221,N_6859);
or U8515 (N_8515,N_6338,N_7252);
or U8516 (N_8516,N_6206,N_7141);
and U8517 (N_8517,N_6457,N_7376);
and U8518 (N_8518,N_7456,N_6206);
nand U8519 (N_8519,N_7087,N_6845);
xor U8520 (N_8520,N_6559,N_7071);
or U8521 (N_8521,N_7493,N_6901);
and U8522 (N_8522,N_7338,N_7171);
nand U8523 (N_8523,N_6837,N_6841);
or U8524 (N_8524,N_6255,N_6670);
and U8525 (N_8525,N_6986,N_7373);
nand U8526 (N_8526,N_6511,N_7013);
nor U8527 (N_8527,N_7183,N_6205);
or U8528 (N_8528,N_6477,N_6124);
nand U8529 (N_8529,N_7479,N_7130);
nand U8530 (N_8530,N_7239,N_7120);
nor U8531 (N_8531,N_7023,N_6201);
nand U8532 (N_8532,N_6075,N_7421);
xor U8533 (N_8533,N_6621,N_6720);
nand U8534 (N_8534,N_6412,N_6048);
nand U8535 (N_8535,N_7043,N_6335);
or U8536 (N_8536,N_6613,N_6836);
and U8537 (N_8537,N_6450,N_6770);
nor U8538 (N_8538,N_7317,N_6021);
nor U8539 (N_8539,N_7377,N_7104);
or U8540 (N_8540,N_6237,N_6797);
or U8541 (N_8541,N_6135,N_7226);
or U8542 (N_8542,N_7058,N_7113);
or U8543 (N_8543,N_6136,N_6245);
and U8544 (N_8544,N_6857,N_6746);
nor U8545 (N_8545,N_6644,N_6067);
or U8546 (N_8546,N_6180,N_7009);
nor U8547 (N_8547,N_6081,N_6323);
and U8548 (N_8548,N_6598,N_6868);
and U8549 (N_8549,N_7265,N_6110);
nor U8550 (N_8550,N_7467,N_6539);
nand U8551 (N_8551,N_6441,N_6506);
nor U8552 (N_8552,N_7366,N_6325);
nor U8553 (N_8553,N_6421,N_6829);
nor U8554 (N_8554,N_6684,N_6530);
nor U8555 (N_8555,N_7090,N_7025);
xnor U8556 (N_8556,N_6485,N_7119);
nor U8557 (N_8557,N_6994,N_7050);
and U8558 (N_8558,N_6070,N_7118);
nand U8559 (N_8559,N_6656,N_6669);
nor U8560 (N_8560,N_6521,N_6248);
or U8561 (N_8561,N_6640,N_6145);
xor U8562 (N_8562,N_6958,N_7256);
nand U8563 (N_8563,N_6944,N_6259);
or U8564 (N_8564,N_6863,N_6082);
xor U8565 (N_8565,N_6018,N_7243);
xor U8566 (N_8566,N_7333,N_7006);
or U8567 (N_8567,N_6891,N_6658);
and U8568 (N_8568,N_7229,N_6257);
nor U8569 (N_8569,N_6241,N_7356);
and U8570 (N_8570,N_6015,N_6584);
or U8571 (N_8571,N_6715,N_7159);
nand U8572 (N_8572,N_6528,N_7063);
nand U8573 (N_8573,N_6155,N_6987);
xor U8574 (N_8574,N_7169,N_6989);
nor U8575 (N_8575,N_6302,N_6300);
and U8576 (N_8576,N_6352,N_6277);
nand U8577 (N_8577,N_6911,N_6351);
or U8578 (N_8578,N_6447,N_6693);
or U8579 (N_8579,N_7115,N_7155);
nand U8580 (N_8580,N_7200,N_6321);
nor U8581 (N_8581,N_7313,N_7233);
xnor U8582 (N_8582,N_6658,N_6530);
and U8583 (N_8583,N_6475,N_6569);
or U8584 (N_8584,N_7485,N_7304);
xnor U8585 (N_8585,N_7022,N_6060);
xnor U8586 (N_8586,N_6224,N_7274);
or U8587 (N_8587,N_6470,N_6823);
or U8588 (N_8588,N_6504,N_7012);
nand U8589 (N_8589,N_6613,N_6770);
and U8590 (N_8590,N_7072,N_6240);
nand U8591 (N_8591,N_7040,N_6311);
nand U8592 (N_8592,N_6422,N_6705);
or U8593 (N_8593,N_6550,N_6553);
and U8594 (N_8594,N_7145,N_6565);
or U8595 (N_8595,N_6584,N_6031);
or U8596 (N_8596,N_6787,N_7392);
nand U8597 (N_8597,N_6627,N_6644);
xnor U8598 (N_8598,N_6372,N_6779);
or U8599 (N_8599,N_7222,N_6720);
nand U8600 (N_8600,N_6428,N_6233);
or U8601 (N_8601,N_7266,N_7255);
or U8602 (N_8602,N_7210,N_6223);
xor U8603 (N_8603,N_7250,N_6626);
xnor U8604 (N_8604,N_6758,N_6339);
nand U8605 (N_8605,N_6913,N_6804);
or U8606 (N_8606,N_6756,N_6250);
and U8607 (N_8607,N_6371,N_6515);
and U8608 (N_8608,N_6798,N_6655);
xnor U8609 (N_8609,N_6480,N_6868);
and U8610 (N_8610,N_6273,N_6047);
nand U8611 (N_8611,N_6594,N_6867);
and U8612 (N_8612,N_6088,N_7276);
nand U8613 (N_8613,N_6761,N_7056);
nor U8614 (N_8614,N_6600,N_6560);
or U8615 (N_8615,N_6908,N_6322);
nand U8616 (N_8616,N_6023,N_6645);
and U8617 (N_8617,N_7241,N_6411);
or U8618 (N_8618,N_6475,N_7376);
nand U8619 (N_8619,N_6744,N_6098);
or U8620 (N_8620,N_6498,N_6793);
or U8621 (N_8621,N_6137,N_6621);
or U8622 (N_8622,N_6936,N_7271);
nor U8623 (N_8623,N_6424,N_7192);
nor U8624 (N_8624,N_7253,N_6055);
nor U8625 (N_8625,N_7149,N_6205);
nand U8626 (N_8626,N_6130,N_7382);
and U8627 (N_8627,N_7036,N_7021);
nor U8628 (N_8628,N_7298,N_6771);
nor U8629 (N_8629,N_7068,N_6981);
nand U8630 (N_8630,N_6011,N_7210);
nor U8631 (N_8631,N_7196,N_6524);
nand U8632 (N_8632,N_6532,N_7152);
xnor U8633 (N_8633,N_7478,N_7452);
xnor U8634 (N_8634,N_6109,N_6589);
xnor U8635 (N_8635,N_7433,N_7254);
and U8636 (N_8636,N_6278,N_6989);
and U8637 (N_8637,N_6398,N_6273);
nor U8638 (N_8638,N_6162,N_6937);
nor U8639 (N_8639,N_7444,N_6920);
nand U8640 (N_8640,N_7439,N_6657);
nor U8641 (N_8641,N_6744,N_6596);
or U8642 (N_8642,N_7177,N_6713);
nor U8643 (N_8643,N_6874,N_6373);
and U8644 (N_8644,N_6264,N_6491);
nor U8645 (N_8645,N_7343,N_6729);
nor U8646 (N_8646,N_6570,N_6855);
nor U8647 (N_8647,N_6943,N_6865);
or U8648 (N_8648,N_6270,N_7364);
and U8649 (N_8649,N_6462,N_6890);
nor U8650 (N_8650,N_6769,N_7160);
or U8651 (N_8651,N_6750,N_6667);
nor U8652 (N_8652,N_6084,N_6314);
xnor U8653 (N_8653,N_7478,N_7134);
and U8654 (N_8654,N_7327,N_6955);
nand U8655 (N_8655,N_6063,N_6296);
nand U8656 (N_8656,N_6808,N_7250);
or U8657 (N_8657,N_6924,N_7197);
nor U8658 (N_8658,N_6447,N_6093);
or U8659 (N_8659,N_6292,N_6299);
or U8660 (N_8660,N_6633,N_6501);
nor U8661 (N_8661,N_6248,N_7403);
nor U8662 (N_8662,N_6070,N_6570);
nor U8663 (N_8663,N_7347,N_7455);
and U8664 (N_8664,N_6314,N_6320);
nor U8665 (N_8665,N_6689,N_6606);
nand U8666 (N_8666,N_7001,N_7140);
nand U8667 (N_8667,N_6505,N_6209);
nor U8668 (N_8668,N_7255,N_6213);
or U8669 (N_8669,N_6308,N_6452);
and U8670 (N_8670,N_6975,N_6992);
nand U8671 (N_8671,N_6213,N_7367);
or U8672 (N_8672,N_6147,N_6592);
nand U8673 (N_8673,N_6873,N_6287);
and U8674 (N_8674,N_6617,N_7312);
nand U8675 (N_8675,N_6203,N_6640);
nand U8676 (N_8676,N_6255,N_6268);
and U8677 (N_8677,N_7101,N_6218);
and U8678 (N_8678,N_6493,N_6807);
xor U8679 (N_8679,N_6971,N_6473);
xnor U8680 (N_8680,N_7155,N_6880);
nor U8681 (N_8681,N_6506,N_6315);
or U8682 (N_8682,N_7228,N_6628);
nand U8683 (N_8683,N_6571,N_6789);
and U8684 (N_8684,N_6025,N_7325);
nor U8685 (N_8685,N_7277,N_6673);
or U8686 (N_8686,N_6456,N_7124);
and U8687 (N_8687,N_6337,N_6559);
nand U8688 (N_8688,N_7484,N_7404);
and U8689 (N_8689,N_7219,N_6662);
and U8690 (N_8690,N_6741,N_6075);
nor U8691 (N_8691,N_6357,N_6162);
or U8692 (N_8692,N_7369,N_6801);
and U8693 (N_8693,N_6153,N_7175);
nand U8694 (N_8694,N_6657,N_6327);
nor U8695 (N_8695,N_6631,N_6903);
nor U8696 (N_8696,N_6324,N_6236);
nand U8697 (N_8697,N_6958,N_6454);
nor U8698 (N_8698,N_7093,N_7117);
nor U8699 (N_8699,N_7256,N_6027);
xor U8700 (N_8700,N_6647,N_6684);
nor U8701 (N_8701,N_7100,N_7388);
nor U8702 (N_8702,N_7313,N_6216);
and U8703 (N_8703,N_7348,N_6161);
nand U8704 (N_8704,N_6227,N_7114);
nand U8705 (N_8705,N_6092,N_6110);
or U8706 (N_8706,N_6677,N_7212);
and U8707 (N_8707,N_7210,N_7109);
nor U8708 (N_8708,N_6567,N_7132);
and U8709 (N_8709,N_6694,N_6786);
or U8710 (N_8710,N_7037,N_6213);
nand U8711 (N_8711,N_6107,N_6644);
and U8712 (N_8712,N_6524,N_6772);
nor U8713 (N_8713,N_7483,N_6439);
or U8714 (N_8714,N_7054,N_6069);
nand U8715 (N_8715,N_7379,N_7122);
or U8716 (N_8716,N_7489,N_6955);
nor U8717 (N_8717,N_6519,N_6207);
or U8718 (N_8718,N_6519,N_6040);
nand U8719 (N_8719,N_6996,N_6067);
nand U8720 (N_8720,N_6340,N_6560);
nor U8721 (N_8721,N_7258,N_6637);
and U8722 (N_8722,N_6390,N_6040);
or U8723 (N_8723,N_6786,N_6217);
nor U8724 (N_8724,N_7025,N_7437);
xnor U8725 (N_8725,N_6429,N_6718);
or U8726 (N_8726,N_6002,N_7327);
or U8727 (N_8727,N_6249,N_6533);
and U8728 (N_8728,N_7499,N_6986);
nand U8729 (N_8729,N_6404,N_6423);
and U8730 (N_8730,N_7401,N_6745);
xor U8731 (N_8731,N_6094,N_7329);
nor U8732 (N_8732,N_7420,N_6286);
or U8733 (N_8733,N_6469,N_6514);
or U8734 (N_8734,N_6174,N_7222);
and U8735 (N_8735,N_7421,N_6310);
nor U8736 (N_8736,N_7447,N_6863);
xnor U8737 (N_8737,N_6619,N_6302);
or U8738 (N_8738,N_7094,N_7076);
nor U8739 (N_8739,N_6441,N_6766);
or U8740 (N_8740,N_7402,N_7156);
and U8741 (N_8741,N_6733,N_6550);
nor U8742 (N_8742,N_6539,N_7379);
and U8743 (N_8743,N_6254,N_6577);
nor U8744 (N_8744,N_6108,N_6447);
nand U8745 (N_8745,N_6574,N_6393);
and U8746 (N_8746,N_7293,N_6531);
and U8747 (N_8747,N_6308,N_6087);
nor U8748 (N_8748,N_7030,N_7403);
nor U8749 (N_8749,N_6816,N_6975);
xnor U8750 (N_8750,N_7497,N_7415);
nor U8751 (N_8751,N_6388,N_6734);
nor U8752 (N_8752,N_7487,N_7058);
nand U8753 (N_8753,N_6088,N_6738);
xnor U8754 (N_8754,N_6973,N_6656);
or U8755 (N_8755,N_6688,N_6159);
nand U8756 (N_8756,N_7346,N_6193);
and U8757 (N_8757,N_6214,N_6479);
and U8758 (N_8758,N_6532,N_6261);
and U8759 (N_8759,N_7361,N_6561);
nor U8760 (N_8760,N_7369,N_6225);
or U8761 (N_8761,N_6959,N_7101);
xnor U8762 (N_8762,N_6045,N_6060);
nand U8763 (N_8763,N_6578,N_7305);
nand U8764 (N_8764,N_6913,N_6792);
nand U8765 (N_8765,N_7379,N_6971);
and U8766 (N_8766,N_6835,N_7371);
nand U8767 (N_8767,N_6661,N_6897);
nor U8768 (N_8768,N_6440,N_6195);
nor U8769 (N_8769,N_7448,N_7345);
nand U8770 (N_8770,N_7192,N_7476);
xnor U8771 (N_8771,N_7317,N_6397);
or U8772 (N_8772,N_6347,N_6718);
nor U8773 (N_8773,N_6536,N_7115);
nor U8774 (N_8774,N_6237,N_7084);
and U8775 (N_8775,N_6907,N_6808);
and U8776 (N_8776,N_6401,N_6384);
and U8777 (N_8777,N_6536,N_6519);
or U8778 (N_8778,N_6568,N_7309);
nand U8779 (N_8779,N_7333,N_6886);
nor U8780 (N_8780,N_6420,N_7387);
or U8781 (N_8781,N_6948,N_7130);
nor U8782 (N_8782,N_6810,N_7486);
nand U8783 (N_8783,N_6484,N_6945);
nor U8784 (N_8784,N_6204,N_7118);
or U8785 (N_8785,N_6572,N_6668);
and U8786 (N_8786,N_6853,N_6697);
or U8787 (N_8787,N_7136,N_6494);
nor U8788 (N_8788,N_6967,N_7034);
or U8789 (N_8789,N_6931,N_6308);
and U8790 (N_8790,N_6699,N_6775);
and U8791 (N_8791,N_6582,N_6807);
xnor U8792 (N_8792,N_6470,N_7493);
or U8793 (N_8793,N_6918,N_7424);
or U8794 (N_8794,N_6077,N_6137);
and U8795 (N_8795,N_7034,N_7100);
or U8796 (N_8796,N_7058,N_6462);
nand U8797 (N_8797,N_7496,N_7392);
nor U8798 (N_8798,N_7066,N_7334);
nand U8799 (N_8799,N_6176,N_6056);
xor U8800 (N_8800,N_7228,N_6795);
and U8801 (N_8801,N_6220,N_6873);
or U8802 (N_8802,N_6023,N_7074);
or U8803 (N_8803,N_6321,N_6329);
nor U8804 (N_8804,N_6876,N_7069);
xnor U8805 (N_8805,N_7455,N_6367);
and U8806 (N_8806,N_7170,N_6129);
or U8807 (N_8807,N_6185,N_7358);
or U8808 (N_8808,N_6936,N_6530);
or U8809 (N_8809,N_6535,N_6594);
and U8810 (N_8810,N_7070,N_7278);
xor U8811 (N_8811,N_6288,N_6739);
or U8812 (N_8812,N_6463,N_7078);
nor U8813 (N_8813,N_6175,N_6939);
nand U8814 (N_8814,N_6655,N_6170);
nor U8815 (N_8815,N_6491,N_6272);
xnor U8816 (N_8816,N_6560,N_6626);
or U8817 (N_8817,N_7228,N_7092);
and U8818 (N_8818,N_7138,N_6205);
nor U8819 (N_8819,N_7101,N_6870);
nand U8820 (N_8820,N_6661,N_6366);
nand U8821 (N_8821,N_6364,N_6021);
or U8822 (N_8822,N_6698,N_6718);
xor U8823 (N_8823,N_6059,N_7475);
nor U8824 (N_8824,N_6719,N_6690);
nor U8825 (N_8825,N_6827,N_7424);
and U8826 (N_8826,N_6343,N_6434);
xnor U8827 (N_8827,N_6431,N_7332);
and U8828 (N_8828,N_7118,N_7048);
or U8829 (N_8829,N_6635,N_7158);
nand U8830 (N_8830,N_6151,N_6978);
xnor U8831 (N_8831,N_6363,N_7256);
and U8832 (N_8832,N_6896,N_7163);
and U8833 (N_8833,N_6988,N_6687);
nor U8834 (N_8834,N_6453,N_6128);
or U8835 (N_8835,N_6860,N_6842);
nor U8836 (N_8836,N_6813,N_7101);
and U8837 (N_8837,N_7192,N_6668);
or U8838 (N_8838,N_7181,N_7156);
or U8839 (N_8839,N_6530,N_7022);
nor U8840 (N_8840,N_7255,N_6245);
and U8841 (N_8841,N_6424,N_6969);
and U8842 (N_8842,N_7399,N_7187);
and U8843 (N_8843,N_6925,N_7212);
nor U8844 (N_8844,N_6697,N_7264);
and U8845 (N_8845,N_7455,N_6959);
or U8846 (N_8846,N_7385,N_7275);
or U8847 (N_8847,N_6283,N_6648);
nor U8848 (N_8848,N_6591,N_6628);
nor U8849 (N_8849,N_6618,N_6117);
nor U8850 (N_8850,N_6855,N_6979);
and U8851 (N_8851,N_6781,N_6750);
nand U8852 (N_8852,N_6776,N_6823);
xnor U8853 (N_8853,N_6874,N_6764);
and U8854 (N_8854,N_7435,N_6124);
xnor U8855 (N_8855,N_7296,N_7076);
or U8856 (N_8856,N_6627,N_7097);
and U8857 (N_8857,N_6563,N_6762);
xnor U8858 (N_8858,N_7265,N_6466);
nand U8859 (N_8859,N_6855,N_6770);
and U8860 (N_8860,N_6412,N_6899);
nor U8861 (N_8861,N_7281,N_7291);
or U8862 (N_8862,N_6728,N_7328);
nor U8863 (N_8863,N_6399,N_6203);
nand U8864 (N_8864,N_7126,N_7452);
and U8865 (N_8865,N_7115,N_6561);
or U8866 (N_8866,N_6579,N_6409);
or U8867 (N_8867,N_7385,N_6509);
nand U8868 (N_8868,N_6398,N_6792);
or U8869 (N_8869,N_7130,N_7057);
xor U8870 (N_8870,N_6255,N_6485);
or U8871 (N_8871,N_7127,N_6485);
or U8872 (N_8872,N_6077,N_7043);
and U8873 (N_8873,N_7446,N_7257);
nand U8874 (N_8874,N_6302,N_6372);
nor U8875 (N_8875,N_6332,N_6396);
nand U8876 (N_8876,N_6515,N_7331);
or U8877 (N_8877,N_7146,N_7484);
nand U8878 (N_8878,N_6400,N_6565);
nand U8879 (N_8879,N_6786,N_6414);
and U8880 (N_8880,N_6792,N_6888);
or U8881 (N_8881,N_6340,N_7336);
and U8882 (N_8882,N_6836,N_6400);
xnor U8883 (N_8883,N_6794,N_6214);
or U8884 (N_8884,N_6086,N_6977);
nand U8885 (N_8885,N_7324,N_6339);
or U8886 (N_8886,N_7179,N_6088);
and U8887 (N_8887,N_6411,N_6868);
nor U8888 (N_8888,N_6462,N_6232);
and U8889 (N_8889,N_7148,N_7411);
nand U8890 (N_8890,N_6685,N_6955);
or U8891 (N_8891,N_6199,N_6798);
or U8892 (N_8892,N_6049,N_7047);
or U8893 (N_8893,N_6392,N_7299);
nor U8894 (N_8894,N_6480,N_7258);
nand U8895 (N_8895,N_6351,N_6129);
and U8896 (N_8896,N_6809,N_6076);
or U8897 (N_8897,N_7324,N_7253);
nand U8898 (N_8898,N_6603,N_7474);
and U8899 (N_8899,N_6278,N_6339);
nand U8900 (N_8900,N_7095,N_7254);
or U8901 (N_8901,N_6690,N_7225);
nor U8902 (N_8902,N_7313,N_6269);
nor U8903 (N_8903,N_7229,N_7015);
nand U8904 (N_8904,N_6149,N_6660);
nand U8905 (N_8905,N_7236,N_7355);
nor U8906 (N_8906,N_6881,N_6872);
nor U8907 (N_8907,N_6766,N_6018);
and U8908 (N_8908,N_6827,N_7172);
or U8909 (N_8909,N_6608,N_6684);
xor U8910 (N_8910,N_6101,N_7372);
nor U8911 (N_8911,N_6586,N_6132);
nand U8912 (N_8912,N_6647,N_7011);
and U8913 (N_8913,N_6868,N_6574);
xor U8914 (N_8914,N_6878,N_7381);
or U8915 (N_8915,N_6480,N_6767);
xnor U8916 (N_8916,N_6961,N_6757);
and U8917 (N_8917,N_6108,N_6432);
or U8918 (N_8918,N_6153,N_7432);
and U8919 (N_8919,N_6485,N_6288);
nand U8920 (N_8920,N_6645,N_7107);
or U8921 (N_8921,N_7201,N_6408);
or U8922 (N_8922,N_7013,N_6257);
and U8923 (N_8923,N_6494,N_7283);
and U8924 (N_8924,N_6754,N_6885);
or U8925 (N_8925,N_6144,N_6405);
nand U8926 (N_8926,N_6909,N_6140);
nor U8927 (N_8927,N_6590,N_7457);
nor U8928 (N_8928,N_6132,N_6133);
and U8929 (N_8929,N_6538,N_6864);
nor U8930 (N_8930,N_6018,N_6614);
nor U8931 (N_8931,N_6374,N_6051);
or U8932 (N_8932,N_7182,N_7469);
nand U8933 (N_8933,N_7012,N_6774);
xor U8934 (N_8934,N_7119,N_7313);
xnor U8935 (N_8935,N_6231,N_6298);
and U8936 (N_8936,N_7319,N_6879);
nand U8937 (N_8937,N_7334,N_6058);
and U8938 (N_8938,N_6402,N_6882);
and U8939 (N_8939,N_7133,N_7433);
or U8940 (N_8940,N_7197,N_7194);
xnor U8941 (N_8941,N_6727,N_6294);
nand U8942 (N_8942,N_6581,N_6819);
nand U8943 (N_8943,N_7247,N_7338);
or U8944 (N_8944,N_6442,N_7370);
or U8945 (N_8945,N_7443,N_6524);
xnor U8946 (N_8946,N_7008,N_6735);
and U8947 (N_8947,N_7402,N_6728);
or U8948 (N_8948,N_7391,N_6242);
and U8949 (N_8949,N_6989,N_6550);
nor U8950 (N_8950,N_6515,N_6129);
or U8951 (N_8951,N_7230,N_7266);
nor U8952 (N_8952,N_6942,N_7460);
nand U8953 (N_8953,N_6952,N_6441);
xnor U8954 (N_8954,N_7044,N_6615);
or U8955 (N_8955,N_6452,N_7491);
nor U8956 (N_8956,N_7166,N_6556);
nor U8957 (N_8957,N_7145,N_6409);
nand U8958 (N_8958,N_6101,N_6317);
nand U8959 (N_8959,N_7479,N_7052);
nand U8960 (N_8960,N_6298,N_7355);
and U8961 (N_8961,N_7138,N_6281);
xor U8962 (N_8962,N_6472,N_6716);
nand U8963 (N_8963,N_6154,N_6604);
and U8964 (N_8964,N_6244,N_6410);
nor U8965 (N_8965,N_7253,N_7105);
and U8966 (N_8966,N_6111,N_6010);
and U8967 (N_8967,N_6236,N_6150);
and U8968 (N_8968,N_7403,N_7101);
nor U8969 (N_8969,N_6625,N_6364);
xor U8970 (N_8970,N_7079,N_6429);
nand U8971 (N_8971,N_6416,N_7127);
nor U8972 (N_8972,N_6287,N_6177);
xor U8973 (N_8973,N_6364,N_6203);
nor U8974 (N_8974,N_6635,N_6937);
nor U8975 (N_8975,N_7039,N_7348);
and U8976 (N_8976,N_6548,N_6400);
xor U8977 (N_8977,N_7334,N_6149);
xnor U8978 (N_8978,N_6993,N_6238);
and U8979 (N_8979,N_7267,N_6238);
and U8980 (N_8980,N_6813,N_7061);
nor U8981 (N_8981,N_6338,N_7087);
or U8982 (N_8982,N_6446,N_7036);
nand U8983 (N_8983,N_6961,N_7283);
nor U8984 (N_8984,N_6693,N_7049);
nor U8985 (N_8985,N_6483,N_7444);
nor U8986 (N_8986,N_6257,N_6694);
nand U8987 (N_8987,N_6355,N_7235);
xnor U8988 (N_8988,N_6162,N_6016);
and U8989 (N_8989,N_6377,N_7452);
and U8990 (N_8990,N_6060,N_6406);
nand U8991 (N_8991,N_6571,N_7064);
and U8992 (N_8992,N_6556,N_7090);
and U8993 (N_8993,N_6261,N_7339);
xor U8994 (N_8994,N_6041,N_7327);
or U8995 (N_8995,N_7160,N_6949);
nor U8996 (N_8996,N_6602,N_6531);
and U8997 (N_8997,N_6384,N_7335);
xnor U8998 (N_8998,N_6980,N_6441);
xnor U8999 (N_8999,N_6492,N_6495);
and U9000 (N_9000,N_8192,N_7895);
nor U9001 (N_9001,N_8132,N_8812);
nor U9002 (N_9002,N_8633,N_7746);
or U9003 (N_9003,N_7534,N_7986);
nand U9004 (N_9004,N_8613,N_8223);
or U9005 (N_9005,N_7904,N_8968);
or U9006 (N_9006,N_8568,N_7772);
and U9007 (N_9007,N_7905,N_8660);
and U9008 (N_9008,N_7656,N_8564);
xor U9009 (N_9009,N_7714,N_7738);
xnor U9010 (N_9010,N_7813,N_8327);
and U9011 (N_9011,N_7950,N_8601);
xor U9012 (N_9012,N_8371,N_7901);
and U9013 (N_9013,N_8923,N_7575);
nor U9014 (N_9014,N_8958,N_7703);
nor U9015 (N_9015,N_8733,N_7624);
or U9016 (N_9016,N_7697,N_7885);
nor U9017 (N_9017,N_7934,N_7558);
nor U9018 (N_9018,N_8261,N_8838);
and U9019 (N_9019,N_8406,N_8070);
or U9020 (N_9020,N_7526,N_7594);
and U9021 (N_9021,N_8138,N_7958);
or U9022 (N_9022,N_8074,N_8494);
nor U9023 (N_9023,N_7936,N_7672);
xnor U9024 (N_9024,N_8403,N_8472);
nor U9025 (N_9025,N_7752,N_8875);
xnor U9026 (N_9026,N_8487,N_8753);
or U9027 (N_9027,N_7770,N_7541);
or U9028 (N_9028,N_8190,N_8298);
xor U9029 (N_9029,N_8974,N_8321);
nand U9030 (N_9030,N_7607,N_8609);
or U9031 (N_9031,N_7596,N_8685);
xor U9032 (N_9032,N_8067,N_7865);
nor U9033 (N_9033,N_7768,N_7787);
nor U9034 (N_9034,N_8393,N_8066);
or U9035 (N_9035,N_7573,N_7983);
xnor U9036 (N_9036,N_8616,N_8183);
or U9037 (N_9037,N_7852,N_8091);
and U9038 (N_9038,N_7891,N_7872);
or U9039 (N_9039,N_7828,N_8211);
nand U9040 (N_9040,N_8654,N_7667);
nor U9041 (N_9041,N_8804,N_8082);
xor U9042 (N_9042,N_7794,N_7991);
xor U9043 (N_9043,N_8763,N_7537);
nor U9044 (N_9044,N_8922,N_8554);
nand U9045 (N_9045,N_8398,N_8543);
nand U9046 (N_9046,N_8598,N_8892);
nor U9047 (N_9047,N_7643,N_7835);
and U9048 (N_9048,N_8129,N_7957);
and U9049 (N_9049,N_8786,N_8064);
nor U9050 (N_9050,N_8545,N_8574);
nor U9051 (N_9051,N_7825,N_8967);
nand U9052 (N_9052,N_8483,N_8374);
nand U9053 (N_9053,N_7932,N_8825);
nand U9054 (N_9054,N_8260,N_7941);
and U9055 (N_9055,N_8302,N_7887);
nor U9056 (N_9056,N_7733,N_8741);
nor U9057 (N_9057,N_8764,N_8796);
or U9058 (N_9058,N_8359,N_8397);
or U9059 (N_9059,N_7760,N_8936);
nand U9060 (N_9060,N_8788,N_7911);
or U9061 (N_9061,N_7559,N_8452);
and U9062 (N_9062,N_8384,N_7511);
nor U9063 (N_9063,N_8639,N_8336);
and U9064 (N_9064,N_7731,N_8760);
and U9065 (N_9065,N_8428,N_8048);
nand U9066 (N_9066,N_8343,N_8001);
nand U9067 (N_9067,N_8530,N_8439);
and U9068 (N_9068,N_7671,N_8556);
or U9069 (N_9069,N_7707,N_8592);
or U9070 (N_9070,N_7755,N_8931);
or U9071 (N_9071,N_8089,N_7786);
nand U9072 (N_9072,N_7871,N_8122);
and U9073 (N_9073,N_7664,N_8215);
nand U9074 (N_9074,N_8809,N_8293);
xnor U9075 (N_9075,N_8262,N_7778);
nor U9076 (N_9076,N_8068,N_8092);
and U9077 (N_9077,N_8345,N_8474);
and U9078 (N_9078,N_8444,N_8577);
xor U9079 (N_9079,N_8038,N_8532);
or U9080 (N_9080,N_8050,N_8843);
nand U9081 (N_9081,N_7970,N_7998);
and U9082 (N_9082,N_8940,N_8501);
and U9083 (N_9083,N_7613,N_8346);
and U9084 (N_9084,N_8728,N_8350);
xnor U9085 (N_9085,N_7536,N_8306);
or U9086 (N_9086,N_7879,N_8236);
and U9087 (N_9087,N_7914,N_8157);
nor U9088 (N_9088,N_8168,N_8593);
and U9089 (N_9089,N_8715,N_8954);
and U9090 (N_9090,N_8751,N_7732);
or U9091 (N_9091,N_7886,N_7681);
xnor U9092 (N_9092,N_8136,N_8959);
nand U9093 (N_9093,N_8789,N_8917);
nand U9094 (N_9094,N_7799,N_7706);
and U9095 (N_9095,N_7636,N_7845);
xnor U9096 (N_9096,N_7574,N_7780);
and U9097 (N_9097,N_8198,N_8857);
xnor U9098 (N_9098,N_8233,N_7759);
nand U9099 (N_9099,N_8182,N_8539);
nor U9100 (N_9100,N_8839,N_8106);
nand U9101 (N_9101,N_7723,N_8280);
nand U9102 (N_9102,N_8623,N_8755);
and U9103 (N_9103,N_8934,N_7682);
nor U9104 (N_9104,N_8188,N_7595);
or U9105 (N_9105,N_8228,N_8005);
or U9106 (N_9106,N_8746,N_8939);
nand U9107 (N_9107,N_8222,N_7603);
and U9108 (N_9108,N_8098,N_8322);
and U9109 (N_9109,N_8034,N_8110);
and U9110 (N_9110,N_8770,N_8376);
and U9111 (N_9111,N_8078,N_7884);
and U9112 (N_9112,N_7962,N_8480);
nor U9113 (N_9113,N_7629,N_7539);
or U9114 (N_9114,N_8982,N_7668);
nor U9115 (N_9115,N_8693,N_8818);
or U9116 (N_9116,N_8529,N_8295);
nor U9117 (N_9117,N_8705,N_7822);
and U9118 (N_9118,N_8666,N_8266);
and U9119 (N_9119,N_8737,N_8373);
and U9120 (N_9120,N_7517,N_8538);
or U9121 (N_9121,N_8077,N_7981);
nand U9122 (N_9122,N_8244,N_8862);
or U9123 (N_9123,N_7920,N_8535);
nor U9124 (N_9124,N_8853,N_8684);
nand U9125 (N_9125,N_8916,N_7652);
nand U9126 (N_9126,N_8665,N_8235);
nand U9127 (N_9127,N_8525,N_8097);
nand U9128 (N_9128,N_8015,N_8976);
nand U9129 (N_9129,N_8218,N_8184);
nor U9130 (N_9130,N_8987,N_8159);
nor U9131 (N_9131,N_8890,N_7561);
nor U9132 (N_9132,N_7639,N_8754);
and U9133 (N_9133,N_8863,N_8185);
nand U9134 (N_9134,N_7565,N_8929);
nand U9135 (N_9135,N_8012,N_8630);
and U9136 (N_9136,N_8626,N_8407);
or U9137 (N_9137,N_8200,N_8347);
nand U9138 (N_9138,N_7899,N_8986);
nand U9139 (N_9139,N_7586,N_8051);
or U9140 (N_9140,N_8793,N_8020);
nand U9141 (N_9141,N_7740,N_8411);
or U9142 (N_9142,N_7571,N_8820);
or U9143 (N_9143,N_8204,N_7698);
nand U9144 (N_9144,N_8632,N_7763);
or U9145 (N_9145,N_8864,N_7655);
nand U9146 (N_9146,N_7680,N_8169);
nor U9147 (N_9147,N_8978,N_8481);
xor U9148 (N_9148,N_8860,N_8251);
and U9149 (N_9149,N_8600,N_8305);
nand U9150 (N_9150,N_7519,N_8840);
and U9151 (N_9151,N_8166,N_7836);
or U9152 (N_9152,N_7612,N_8561);
nor U9153 (N_9153,N_8273,N_8769);
and U9154 (N_9154,N_7545,N_8844);
nor U9155 (N_9155,N_7720,N_8650);
nand U9156 (N_9156,N_8914,N_7583);
or U9157 (N_9157,N_8671,N_8477);
and U9158 (N_9158,N_8338,N_7789);
nand U9159 (N_9159,N_8714,N_8328);
nor U9160 (N_9160,N_8552,N_8674);
nor U9161 (N_9161,N_8387,N_8017);
nand U9162 (N_9162,N_8413,N_8022);
nor U9163 (N_9163,N_8207,N_7618);
or U9164 (N_9164,N_8563,N_8555);
nand U9165 (N_9165,N_8738,N_8856);
nor U9166 (N_9166,N_8093,N_8269);
nand U9167 (N_9167,N_8649,N_8283);
and U9168 (N_9168,N_8317,N_7555);
nand U9169 (N_9169,N_7873,N_8998);
nor U9170 (N_9170,N_8248,N_8203);
nand U9171 (N_9171,N_8622,N_8885);
nand U9172 (N_9172,N_8652,N_7843);
or U9173 (N_9173,N_8663,N_7966);
or U9174 (N_9174,N_8994,N_8794);
nand U9175 (N_9175,N_7553,N_7995);
nor U9176 (N_9176,N_8757,N_8697);
nand U9177 (N_9177,N_7666,N_8043);
nor U9178 (N_9178,N_7546,N_8526);
nor U9179 (N_9179,N_8915,N_8882);
or U9180 (N_9180,N_7951,N_8118);
nor U9181 (N_9181,N_7676,N_7600);
or U9182 (N_9182,N_8276,N_8055);
nand U9183 (N_9183,N_8320,N_7635);
nand U9184 (N_9184,N_8712,N_8806);
and U9185 (N_9185,N_7749,N_8523);
and U9186 (N_9186,N_8582,N_8502);
nand U9187 (N_9187,N_7501,N_8139);
or U9188 (N_9188,N_7520,N_7812);
xor U9189 (N_9189,N_8724,N_8807);
nor U9190 (N_9190,N_8509,N_8520);
and U9191 (N_9191,N_8521,N_8859);
nor U9192 (N_9192,N_8558,N_8517);
or U9193 (N_9193,N_7708,N_8165);
or U9194 (N_9194,N_8579,N_8114);
and U9195 (N_9195,N_7632,N_8516);
and U9196 (N_9196,N_8872,N_8960);
xnor U9197 (N_9197,N_7869,N_8816);
or U9198 (N_9198,N_7900,N_8268);
nand U9199 (N_9199,N_7971,N_8352);
or U9200 (N_9200,N_8656,N_7521);
or U9201 (N_9201,N_8101,N_8927);
and U9202 (N_9202,N_7599,N_7965);
or U9203 (N_9203,N_8057,N_8026);
and U9204 (N_9204,N_8636,N_8588);
nand U9205 (N_9205,N_8271,N_8478);
nand U9206 (N_9206,N_8498,N_8935);
nand U9207 (N_9207,N_8944,N_8108);
nor U9208 (N_9208,N_8435,N_8785);
and U9209 (N_9209,N_8158,N_7504);
or U9210 (N_9210,N_8175,N_8941);
and U9211 (N_9211,N_8572,N_7826);
nand U9212 (N_9212,N_8433,N_8044);
nor U9213 (N_9213,N_8833,N_8897);
or U9214 (N_9214,N_8979,N_7798);
or U9215 (N_9215,N_8379,N_7699);
or U9216 (N_9216,N_7592,N_7530);
and U9217 (N_9217,N_8135,N_8566);
nor U9218 (N_9218,N_8908,N_7633);
and U9219 (N_9219,N_8199,N_8596);
nand U9220 (N_9220,N_7771,N_7846);
nor U9221 (N_9221,N_7989,N_7975);
or U9222 (N_9222,N_8971,N_7518);
or U9223 (N_9223,N_8427,N_8725);
nand U9224 (N_9224,N_8606,N_7614);
nor U9225 (N_9225,N_8634,N_8454);
or U9226 (N_9226,N_7584,N_8670);
nor U9227 (N_9227,N_7711,N_8604);
nor U9228 (N_9228,N_7940,N_7510);
xnor U9229 (N_9229,N_7973,N_8515);
or U9230 (N_9230,N_7544,N_8750);
nand U9231 (N_9231,N_8469,N_7976);
nor U9232 (N_9232,N_8476,N_8581);
and U9233 (N_9233,N_7701,N_8446);
nand U9234 (N_9234,N_8732,N_7857);
xor U9235 (N_9235,N_7792,N_8086);
and U9236 (N_9236,N_8930,N_8599);
and U9237 (N_9237,N_8080,N_8434);
nand U9238 (N_9238,N_8676,N_8287);
and U9239 (N_9239,N_7999,N_7811);
and U9240 (N_9240,N_7921,N_7508);
nor U9241 (N_9241,N_7734,N_7619);
nor U9242 (N_9242,N_8368,N_7719);
and U9243 (N_9243,N_8042,N_7939);
nor U9244 (N_9244,N_8748,N_8881);
or U9245 (N_9245,N_8300,N_8871);
or U9246 (N_9246,N_7694,N_7834);
and U9247 (N_9247,N_7906,N_7659);
nor U9248 (N_9248,N_8422,N_8326);
nor U9249 (N_9249,N_8342,N_8528);
and U9250 (N_9250,N_8619,N_8717);
and U9251 (N_9251,N_8205,N_8194);
xor U9252 (N_9252,N_8401,N_7610);
nand U9253 (N_9253,N_8008,N_8292);
nand U9254 (N_9254,N_8332,N_7773);
or U9255 (N_9255,N_8255,N_7915);
nor U9256 (N_9256,N_8887,N_7809);
or U9257 (N_9257,N_8576,N_8800);
nor U9258 (N_9258,N_8551,N_7816);
or U9259 (N_9259,N_7867,N_7918);
or U9260 (N_9260,N_8756,N_8083);
and U9261 (N_9261,N_7882,N_8314);
xnor U9262 (N_9262,N_8220,N_7868);
nand U9263 (N_9263,N_7687,N_7754);
xnor U9264 (N_9264,N_7705,N_7827);
and U9265 (N_9265,N_7564,N_8503);
nor U9266 (N_9266,N_8865,N_8988);
nand U9267 (N_9267,N_8679,N_8729);
nor U9268 (N_9268,N_8720,N_8337);
nor U9269 (N_9269,N_7689,N_8781);
nor U9270 (N_9270,N_8821,N_7750);
nor U9271 (N_9271,N_7739,N_8285);
nand U9272 (N_9272,N_8615,N_8212);
and U9273 (N_9273,N_8040,N_8681);
nor U9274 (N_9274,N_8365,N_7551);
or U9275 (N_9275,N_8669,N_7590);
or U9276 (N_9276,N_7963,N_8814);
or U9277 (N_9277,N_7943,N_8824);
nand U9278 (N_9278,N_8873,N_7978);
nor U9279 (N_9279,N_7657,N_8226);
or U9280 (N_9280,N_8918,N_7888);
nand U9281 (N_9281,N_8363,N_8799);
nand U9282 (N_9282,N_8726,N_8851);
or U9283 (N_9283,N_8163,N_7937);
xor U9284 (N_9284,N_7729,N_8569);
nand U9285 (N_9285,N_7678,N_8229);
xnor U9286 (N_9286,N_8852,N_8969);
nor U9287 (N_9287,N_8698,N_8088);
nor U9288 (N_9288,N_8618,N_8062);
nand U9289 (N_9289,N_8178,N_8827);
nor U9290 (N_9290,N_8470,N_7540);
nand U9291 (N_9291,N_8497,N_8585);
nor U9292 (N_9292,N_8096,N_7529);
and U9293 (N_9293,N_8234,N_7806);
or U9294 (N_9294,N_8111,N_7945);
nand U9295 (N_9295,N_7721,N_8115);
nand U9296 (N_9296,N_8777,N_8531);
nor U9297 (N_9297,N_8339,N_8874);
and U9298 (N_9298,N_7860,N_8780);
nor U9299 (N_9299,N_8426,N_8399);
and U9300 (N_9300,N_7810,N_7982);
nand U9301 (N_9301,N_8404,N_8173);
and U9302 (N_9302,N_8016,N_8784);
or U9303 (N_9303,N_8107,N_8161);
and U9304 (N_9304,N_7985,N_8955);
and U9305 (N_9305,N_7647,N_8045);
nand U9306 (N_9306,N_8629,N_8683);
or U9307 (N_9307,N_8761,N_8471);
or U9308 (N_9308,N_8148,N_8488);
and U9309 (N_9309,N_8180,N_8113);
nand U9310 (N_9310,N_8191,N_8999);
or U9311 (N_9311,N_7912,N_7663);
and U9312 (N_9312,N_8032,N_8870);
nor U9313 (N_9313,N_8011,N_8625);
or U9314 (N_9314,N_8036,N_8484);
or U9315 (N_9315,N_8779,N_8217);
and U9316 (N_9316,N_7874,N_8239);
nor U9317 (N_9317,N_8252,N_8142);
nor U9318 (N_9318,N_8420,N_8993);
nand U9319 (N_9319,N_8854,N_7675);
or U9320 (N_9320,N_8430,N_8846);
xor U9321 (N_9321,N_7620,N_8962);
nor U9322 (N_9322,N_8928,N_7850);
and U9323 (N_9323,N_7777,N_8534);
or U9324 (N_9324,N_7820,N_8647);
nand U9325 (N_9325,N_8186,N_8297);
or U9326 (N_9326,N_8224,N_7690);
nor U9327 (N_9327,N_8721,N_8201);
or U9328 (N_9328,N_8391,N_8752);
and U9329 (N_9329,N_7829,N_7742);
nand U9330 (N_9330,N_8692,N_7863);
and U9331 (N_9331,N_8099,N_8637);
and U9332 (N_9332,N_7897,N_8948);
nor U9333 (N_9333,N_8541,N_8349);
or U9334 (N_9334,N_8522,N_7870);
nand U9335 (N_9335,N_7507,N_8855);
and U9336 (N_9336,N_8884,N_7830);
or U9337 (N_9337,N_7837,N_8004);
nand U9338 (N_9338,N_7696,N_8331);
nand U9339 (N_9339,N_8214,N_7929);
and U9340 (N_9340,N_8653,N_8858);
and U9341 (N_9341,N_7516,N_8586);
or U9342 (N_9342,N_8690,N_8208);
xnor U9343 (N_9343,N_7821,N_8803);
and U9344 (N_9344,N_8467,N_8571);
and U9345 (N_9345,N_8627,N_8731);
and U9346 (N_9346,N_7844,N_8776);
xnor U9347 (N_9347,N_8357,N_8258);
nand U9348 (N_9348,N_7737,N_7716);
nand U9349 (N_9349,N_7692,N_7758);
or U9350 (N_9350,N_8990,N_8787);
or U9351 (N_9351,N_8912,N_7992);
or U9352 (N_9352,N_8318,N_7726);
or U9353 (N_9353,N_7704,N_8952);
or U9354 (N_9354,N_8003,N_8354);
xor U9355 (N_9355,N_8805,N_8418);
nor U9356 (N_9356,N_8058,N_7700);
nand U9357 (N_9357,N_7621,N_8847);
xnor U9358 (N_9358,N_7557,N_8308);
or U9359 (N_9359,N_7500,N_8451);
xor U9360 (N_9360,N_8155,N_7823);
and U9361 (N_9361,N_8143,N_8028);
or U9362 (N_9362,N_7686,N_7762);
and U9363 (N_9363,N_8014,N_7515);
or U9364 (N_9364,N_8841,N_8176);
nand U9365 (N_9365,N_8270,N_8241);
and U9366 (N_9366,N_8826,N_7736);
nor U9367 (N_9367,N_7611,N_7572);
xnor U9368 (N_9368,N_8282,N_7630);
nor U9369 (N_9369,N_7741,N_8240);
nor U9370 (N_9370,N_7807,N_8395);
or U9371 (N_9371,N_8758,N_8723);
or U9372 (N_9372,N_8602,N_8673);
nor U9373 (N_9373,N_7935,N_7568);
or U9374 (N_9374,N_8675,N_7841);
nand U9375 (N_9375,N_8594,N_7925);
xnor U9376 (N_9376,N_8364,N_7566);
nor U9377 (N_9377,N_7684,N_8031);
nor U9378 (N_9378,N_7832,N_8035);
and U9379 (N_9379,N_8167,N_8333);
nand U9380 (N_9380,N_8655,N_7717);
or U9381 (N_9381,N_8866,N_8947);
nor U9382 (N_9382,N_7570,N_8059);
nor U9383 (N_9383,N_8878,N_7864);
xor U9384 (N_9384,N_8351,N_7604);
and U9385 (N_9385,N_8810,N_8313);
and U9386 (N_9386,N_8815,N_8583);
nor U9387 (N_9387,N_8834,N_8250);
nor U9388 (N_9388,N_8711,N_8025);
nand U9389 (N_9389,N_8938,N_8117);
nor U9390 (N_9390,N_8460,N_7964);
nand U9391 (N_9391,N_8791,N_8542);
nor U9392 (N_9392,N_8441,N_7756);
and U9393 (N_9393,N_7674,N_8053);
or U9394 (N_9394,N_7522,N_8464);
nand U9395 (N_9395,N_8975,N_7953);
and U9396 (N_9396,N_8970,N_8964);
and U9397 (N_9397,N_7783,N_8105);
nor U9398 (N_9398,N_8382,N_8390);
xor U9399 (N_9399,N_8850,N_8664);
nand U9400 (N_9400,N_8030,N_8849);
nand U9401 (N_9401,N_7990,N_8771);
and U9402 (N_9402,N_8249,N_8533);
nor U9403 (N_9403,N_7702,N_8473);
or U9404 (N_9404,N_8073,N_7679);
nand U9405 (N_9405,N_7875,N_8324);
nor U9406 (N_9406,N_8553,N_8450);
nand U9407 (N_9407,N_8801,N_8886);
or U9408 (N_9408,N_7877,N_8512);
nand U9409 (N_9409,N_7761,N_7858);
or U9410 (N_9410,N_8745,N_8272);
or U9411 (N_9411,N_8694,N_8876);
and U9412 (N_9412,N_8973,N_8047);
or U9413 (N_9413,N_8565,N_8486);
xnor U9414 (N_9414,N_7637,N_8701);
and U9415 (N_9415,N_8245,N_7903);
xor U9416 (N_9416,N_8680,N_7808);
nor U9417 (N_9417,N_7853,N_7889);
or U9418 (N_9418,N_7724,N_8150);
nand U9419 (N_9419,N_7550,N_8284);
or U9420 (N_9420,N_8505,N_8662);
xnor U9421 (N_9421,N_7993,N_8095);
nor U9422 (N_9422,N_8104,N_7974);
nand U9423 (N_9423,N_7556,N_8710);
nand U9424 (N_9424,N_8279,N_7948);
and U9425 (N_9425,N_7695,N_7790);
nand U9426 (N_9426,N_8511,N_7952);
nor U9427 (N_9427,N_8687,N_8274);
nor U9428 (N_9428,N_8485,N_8808);
nand U9429 (N_9429,N_8410,N_7803);
nand U9430 (N_9430,N_7959,N_8829);
nand U9431 (N_9431,N_7839,N_8232);
xnor U9432 (N_9432,N_7608,N_7597);
and U9433 (N_9433,N_8984,N_8490);
nor U9434 (N_9434,N_7523,N_8344);
and U9435 (N_9435,N_8628,N_7767);
nand U9436 (N_9436,N_8400,N_8310);
and U9437 (N_9437,N_8937,N_8432);
and U9438 (N_9438,N_8924,N_8951);
nand U9439 (N_9439,N_7956,N_7683);
and U9440 (N_9440,N_7650,N_8573);
nor U9441 (N_9441,N_8278,N_7693);
xor U9442 (N_9442,N_8767,N_8288);
and U9443 (N_9443,N_7972,N_7710);
or U9444 (N_9444,N_7745,N_8256);
and U9445 (N_9445,N_7961,N_8595);
or U9446 (N_9446,N_8703,N_7598);
nand U9447 (N_9447,N_8360,N_7791);
or U9448 (N_9448,N_7949,N_8304);
nor U9449 (N_9449,N_7649,N_7727);
nor U9450 (N_9450,N_8965,N_8037);
and U9451 (N_9451,N_7942,N_7751);
nand U9452 (N_9452,N_7960,N_8125);
and U9453 (N_9453,N_8883,N_7893);
and U9454 (N_9454,N_8880,N_8614);
nor U9455 (N_9455,N_7712,N_7585);
and U9456 (N_9456,N_7815,N_8549);
and U9457 (N_9457,N_7669,N_8216);
nor U9458 (N_9458,N_7634,N_8901);
nand U9459 (N_9459,N_8795,N_8635);
or U9460 (N_9460,N_8790,N_8286);
xor U9461 (N_9461,N_7641,N_8624);
nand U9462 (N_9462,N_8953,N_7902);
xor U9463 (N_9463,N_7856,N_8362);
and U9464 (N_9464,N_8130,N_8608);
and U9465 (N_9465,N_7642,N_8550);
and U9466 (N_9466,N_8029,N_7662);
nor U9467 (N_9467,N_8696,N_8296);
nand U9468 (N_9468,N_8380,N_8181);
nand U9469 (N_9469,N_8695,N_7548);
or U9470 (N_9470,N_7589,N_8879);
and U9471 (N_9471,N_8641,N_8455);
and U9472 (N_9472,N_8537,N_8638);
nand U9473 (N_9473,N_8926,N_8039);
or U9474 (N_9474,N_8195,N_7542);
nor U9475 (N_9475,N_8689,N_7769);
nand U9476 (N_9476,N_7797,N_8597);
nor U9477 (N_9477,N_8356,N_8742);
and U9478 (N_9478,N_7862,N_7543);
and U9479 (N_9479,N_8677,N_8506);
nor U9480 (N_9480,N_8891,N_8458);
nor U9481 (N_9481,N_8798,N_8991);
or U9482 (N_9482,N_8196,N_7503);
or U9483 (N_9483,N_7725,N_8997);
nor U9484 (N_9484,N_8699,N_8514);
nor U9485 (N_9485,N_8162,N_8479);
or U9486 (N_9486,N_8076,N_8792);
nand U9487 (N_9487,N_8831,N_7801);
or U9488 (N_9488,N_8465,N_7580);
nor U9489 (N_9489,N_7766,N_8154);
xor U9490 (N_9490,N_7660,N_8219);
and U9491 (N_9491,N_8303,N_7788);
and U9492 (N_9492,N_8686,N_7919);
xnor U9493 (N_9493,N_8981,N_7840);
nand U9494 (N_9494,N_7933,N_8449);
or U9495 (N_9495,N_8417,N_7824);
nand U9496 (N_9496,N_7718,N_7779);
nor U9497 (N_9497,N_8765,N_8943);
or U9498 (N_9498,N_8431,N_8348);
nor U9499 (N_9499,N_8837,N_8591);
xnor U9500 (N_9500,N_7554,N_8651);
nand U9501 (N_9501,N_7715,N_8645);
nor U9502 (N_9502,N_7563,N_8453);
nand U9503 (N_9503,N_8836,N_7833);
or U9504 (N_9504,N_8510,N_8559);
nand U9505 (N_9505,N_8567,N_8766);
nor U9506 (N_9506,N_7977,N_8193);
nand U9507 (N_9507,N_8797,N_7677);
nor U9508 (N_9508,N_8547,N_8919);
or U9509 (N_9509,N_7849,N_8768);
nor U9510 (N_9510,N_8963,N_8366);
and U9511 (N_9511,N_8519,N_8949);
or U9512 (N_9512,N_8445,N_7917);
and U9513 (N_9513,N_8457,N_8009);
nor U9514 (N_9514,N_8906,N_8440);
and U9515 (N_9515,N_7709,N_8772);
and U9516 (N_9516,N_8463,N_7562);
or U9517 (N_9517,N_7646,N_8749);
xor U9518 (N_9518,N_8312,N_8691);
or U9519 (N_9519,N_8492,N_8524);
or U9520 (N_9520,N_8740,N_8832);
and U9521 (N_9521,N_8416,N_7757);
nor U9522 (N_9522,N_8309,N_7800);
nor U9523 (N_9523,N_8747,N_8121);
nor U9524 (N_9524,N_7654,N_8461);
or U9525 (N_9525,N_7547,N_8315);
xnor U9526 (N_9526,N_8153,N_8835);
nor U9527 (N_9527,N_8299,N_7513);
nor U9528 (N_9528,N_8466,N_7617);
nand U9529 (N_9529,N_8081,N_8409);
or U9530 (N_9530,N_8277,N_8210);
and U9531 (N_9531,N_7688,N_7796);
nand U9532 (N_9532,N_8903,N_8065);
or U9533 (N_9533,N_8227,N_8396);
nand U9534 (N_9534,N_8145,N_8056);
nand U9535 (N_9535,N_7781,N_8961);
nor U9536 (N_9536,N_8713,N_8688);
xor U9537 (N_9537,N_8894,N_8358);
nand U9538 (N_9538,N_8932,N_8607);
nand U9539 (N_9539,N_8590,N_8709);
xor U9540 (N_9540,N_8383,N_8330);
xnor U9541 (N_9541,N_8972,N_8557);
nor U9542 (N_9542,N_8124,N_8657);
nor U9543 (N_9543,N_8072,N_7728);
and U9544 (N_9544,N_8718,N_8156);
or U9545 (N_9545,N_7691,N_7898);
or U9546 (N_9546,N_8319,N_8580);
nor U9547 (N_9547,N_8989,N_8775);
or U9548 (N_9548,N_7713,N_8773);
or U9549 (N_9549,N_8024,N_8508);
or U9550 (N_9550,N_7764,N_7665);
and U9551 (N_9551,N_8950,N_7593);
and U9552 (N_9552,N_7842,N_8075);
nand U9553 (N_9553,N_7626,N_8340);
and U9554 (N_9554,N_8079,N_8152);
xnor U9555 (N_9555,N_8722,N_8640);
nor U9556 (N_9556,N_7651,N_7549);
nor U9557 (N_9557,N_8019,N_8381);
nand U9558 (N_9558,N_8621,N_7954);
nand U9559 (N_9559,N_8744,N_7628);
and U9560 (N_9560,N_8378,N_8823);
xnor U9561 (N_9561,N_8783,N_7987);
nor U9562 (N_9562,N_7531,N_7776);
or U9563 (N_9563,N_8149,N_8540);
and U9564 (N_9564,N_7881,N_7930);
nor U9565 (N_9565,N_8617,N_8702);
nand U9566 (N_9566,N_8719,N_7640);
nor U9567 (N_9567,N_8289,N_8372);
and U9568 (N_9568,N_7994,N_8133);
nand U9569 (N_9569,N_8642,N_7876);
or U9570 (N_9570,N_7947,N_8489);
and U9571 (N_9571,N_8109,N_7980);
and U9572 (N_9572,N_7661,N_7908);
nor U9573 (N_9573,N_8762,N_8334);
nand U9574 (N_9574,N_7527,N_8341);
nor U9575 (N_9575,N_8736,N_8243);
nand U9576 (N_9576,N_8518,N_8237);
nand U9577 (N_9577,N_7880,N_7984);
nor U9578 (N_9578,N_8920,N_8323);
xor U9579 (N_9579,N_7805,N_8910);
nand U9580 (N_9580,N_8388,N_8739);
nor U9581 (N_9581,N_8027,N_8225);
nor U9582 (N_9582,N_8611,N_8238);
and U9583 (N_9583,N_7506,N_8706);
nand U9584 (N_9584,N_8405,N_8071);
and U9585 (N_9585,N_8727,N_7775);
nor U9586 (N_9586,N_8493,N_8570);
nand U9587 (N_9587,N_8377,N_8707);
or U9588 (N_9588,N_7627,N_7854);
nand U9589 (N_9589,N_8392,N_8589);
nor U9590 (N_9590,N_7817,N_7606);
xnor U9591 (N_9591,N_7533,N_7765);
or U9592 (N_9592,N_8221,N_8230);
and U9593 (N_9593,N_8909,N_7670);
or U9594 (N_9594,N_8819,N_8160);
or U9595 (N_9595,N_8033,N_7979);
nand U9596 (N_9596,N_8983,N_7855);
or U9597 (N_9597,N_8000,N_8902);
and U9598 (N_9598,N_8845,N_7535);
or U9599 (N_9599,N_8716,N_8456);
nor U9600 (N_9600,N_8049,N_8060);
nor U9601 (N_9601,N_7774,N_8367);
or U9602 (N_9602,N_7524,N_7512);
nand U9603 (N_9603,N_8209,N_8482);
and U9604 (N_9604,N_7944,N_8992);
nor U9605 (N_9605,N_8620,N_7744);
nor U9606 (N_9606,N_8151,N_8448);
or U9607 (N_9607,N_8868,N_7924);
and U9608 (N_9608,N_8010,N_7927);
and U9609 (N_9609,N_7502,N_8822);
or U9610 (N_9610,N_7928,N_8137);
xnor U9611 (N_9611,N_8782,N_7968);
or U9612 (N_9612,N_8375,N_8023);
and U9613 (N_9613,N_8259,N_8389);
nand U9614 (N_9614,N_8100,N_8197);
nor U9615 (N_9615,N_8896,N_8774);
and U9616 (N_9616,N_8500,N_8659);
or U9617 (N_9617,N_7883,N_8946);
and U9618 (N_9618,N_8462,N_7577);
nor U9619 (N_9619,N_8424,N_8667);
xnor U9620 (N_9620,N_7848,N_8899);
or U9621 (N_9621,N_8904,N_7722);
nor U9622 (N_9622,N_7505,N_7532);
xnor U9623 (N_9623,N_8021,N_8889);
or U9624 (N_9624,N_7988,N_7538);
and U9625 (N_9625,N_7591,N_7996);
nor U9626 (N_9626,N_8913,N_7653);
and U9627 (N_9627,N_8830,N_7748);
nand U9628 (N_9628,N_8144,N_8307);
and U9629 (N_9629,N_8504,N_8247);
nor U9630 (N_9630,N_8120,N_8877);
nand U9631 (N_9631,N_7969,N_7818);
xor U9632 (N_9632,N_8893,N_7638);
nand U9633 (N_9633,N_8842,N_8869);
or U9634 (N_9634,N_8447,N_7582);
nor U9635 (N_9635,N_8187,N_8301);
xnor U9636 (N_9636,N_8544,N_8644);
xnor U9637 (N_9637,N_8087,N_8985);
or U9638 (N_9638,N_7896,N_7605);
and U9639 (N_9639,N_7910,N_8164);
and U9640 (N_9640,N_8419,N_8848);
and U9641 (N_9641,N_8429,N_7525);
nor U9642 (N_9642,N_7907,N_8980);
nor U9643 (N_9643,N_8146,N_8646);
nand U9644 (N_9644,N_8933,N_8257);
and U9645 (N_9645,N_8172,N_8421);
nand U9646 (N_9646,N_8828,N_8921);
or U9647 (N_9647,N_7644,N_7866);
and U9648 (N_9648,N_8610,N_7847);
or U9649 (N_9649,N_8402,N_8562);
nand U9650 (N_9650,N_8996,N_8069);
nand U9651 (N_9651,N_7967,N_7923);
and U9652 (N_9652,N_7609,N_8605);
or U9653 (N_9653,N_7931,N_8054);
or U9654 (N_9654,N_7615,N_8900);
or U9655 (N_9655,N_8147,N_7631);
and U9656 (N_9656,N_8743,N_8475);
xor U9657 (N_9657,N_7785,N_7793);
xnor U9658 (N_9658,N_8294,N_8094);
xnor U9659 (N_9659,N_8905,N_8584);
nor U9660 (N_9660,N_8131,N_8867);
xor U9661 (N_9661,N_7997,N_8189);
xnor U9662 (N_9662,N_7509,N_7743);
nand U9663 (N_9663,N_8682,N_8548);
nor U9664 (N_9664,N_8394,N_8802);
nor U9665 (N_9665,N_8587,N_8370);
nor U9666 (N_9666,N_8438,N_8123);
xor U9667 (N_9667,N_8102,N_7890);
nor U9668 (N_9668,N_8275,N_8084);
xor U9669 (N_9669,N_7569,N_8700);
and U9670 (N_9670,N_8170,N_8246);
or U9671 (N_9671,N_8311,N_8668);
or U9672 (N_9672,N_8046,N_7601);
and U9673 (N_9673,N_7579,N_7955);
nor U9674 (N_9674,N_8513,N_8263);
and U9675 (N_9675,N_8202,N_7861);
and U9676 (N_9676,N_8578,N_7673);
or U9677 (N_9677,N_8658,N_8778);
or U9678 (N_9678,N_7814,N_7685);
nand U9679 (N_9679,N_7804,N_8385);
or U9680 (N_9680,N_8335,N_8052);
nand U9681 (N_9681,N_7913,N_8491);
or U9682 (N_9682,N_8995,N_8006);
and U9683 (N_9683,N_7588,N_8496);
or U9684 (N_9684,N_8386,N_8888);
nand U9685 (N_9685,N_8177,N_8468);
nand U9686 (N_9686,N_7560,N_8678);
nor U9687 (N_9687,N_8648,N_7892);
xor U9688 (N_9688,N_8231,N_8603);
nor U9689 (N_9689,N_8612,N_7795);
nand U9690 (N_9690,N_8291,N_7878);
nor U9691 (N_9691,N_7926,N_8325);
nor U9692 (N_9692,N_8361,N_7514);
or U9693 (N_9693,N_8907,N_7784);
and U9694 (N_9694,N_7602,N_8013);
or U9695 (N_9695,N_7578,N_8414);
or U9696 (N_9696,N_8128,N_8817);
and U9697 (N_9697,N_7747,N_8957);
nor U9698 (N_9698,N_8408,N_8316);
nor U9699 (N_9699,N_8442,N_8116);
and U9700 (N_9700,N_8412,N_7859);
or U9701 (N_9701,N_7567,N_8041);
or U9702 (N_9702,N_8174,N_8127);
and U9703 (N_9703,N_8119,N_8103);
or U9704 (N_9704,N_8134,N_8734);
nand U9705 (N_9705,N_7576,N_8672);
or U9706 (N_9706,N_8329,N_8536);
nor U9707 (N_9707,N_8423,N_7622);
nand U9708 (N_9708,N_7802,N_8643);
and U9709 (N_9709,N_8415,N_8735);
nor U9710 (N_9710,N_8575,N_7851);
nor U9711 (N_9711,N_8436,N_7946);
nand U9712 (N_9712,N_8499,N_8898);
or U9713 (N_9713,N_7658,N_8977);
nand U9714 (N_9714,N_8112,N_8281);
and U9715 (N_9715,N_7587,N_8560);
xor U9716 (N_9716,N_7528,N_8527);
nand U9717 (N_9717,N_8206,N_8459);
xor U9718 (N_9718,N_7625,N_8355);
nor U9719 (N_9719,N_7730,N_8495);
and U9720 (N_9720,N_7782,N_8425);
nor U9721 (N_9721,N_8126,N_8267);
xor U9722 (N_9722,N_7909,N_8861);
or U9723 (N_9723,N_8661,N_8171);
xnor U9724 (N_9724,N_7938,N_8002);
nor U9725 (N_9725,N_8140,N_8759);
or U9726 (N_9726,N_8730,N_8813);
nand U9727 (N_9727,N_8213,N_8141);
or U9728 (N_9728,N_8956,N_8443);
and U9729 (N_9729,N_8018,N_7916);
nand U9730 (N_9730,N_8085,N_8063);
nor U9731 (N_9731,N_8942,N_8007);
nand U9732 (N_9732,N_7581,N_7735);
or U9733 (N_9733,N_7894,N_8090);
nor U9734 (N_9734,N_8546,N_8179);
and U9735 (N_9735,N_8911,N_8631);
or U9736 (N_9736,N_8242,N_8966);
or U9737 (N_9737,N_7831,N_8945);
nand U9738 (N_9738,N_8925,N_8061);
nand U9739 (N_9739,N_7922,N_7648);
nor U9740 (N_9740,N_8369,N_8507);
nor U9741 (N_9741,N_8437,N_8265);
or U9742 (N_9742,N_8708,N_8353);
and U9743 (N_9743,N_8290,N_8811);
xnor U9744 (N_9744,N_7819,N_7623);
nor U9745 (N_9745,N_7645,N_8264);
nor U9746 (N_9746,N_7753,N_7552);
nor U9747 (N_9747,N_8254,N_8253);
or U9748 (N_9748,N_7616,N_8895);
nand U9749 (N_9749,N_8704,N_7838);
and U9750 (N_9750,N_8367,N_7685);
xor U9751 (N_9751,N_8892,N_7670);
and U9752 (N_9752,N_7573,N_8632);
xnor U9753 (N_9753,N_8908,N_8567);
nor U9754 (N_9754,N_7655,N_8521);
and U9755 (N_9755,N_8014,N_8800);
and U9756 (N_9756,N_8288,N_8976);
or U9757 (N_9757,N_8437,N_8001);
and U9758 (N_9758,N_7703,N_8679);
nor U9759 (N_9759,N_7936,N_7555);
xnor U9760 (N_9760,N_8037,N_8407);
and U9761 (N_9761,N_7723,N_8587);
or U9762 (N_9762,N_8830,N_8639);
xor U9763 (N_9763,N_7932,N_8285);
nand U9764 (N_9764,N_8401,N_8105);
and U9765 (N_9765,N_8322,N_8527);
or U9766 (N_9766,N_7798,N_8974);
and U9767 (N_9767,N_8970,N_8681);
and U9768 (N_9768,N_8099,N_7936);
nand U9769 (N_9769,N_8318,N_7802);
or U9770 (N_9770,N_7574,N_7599);
nand U9771 (N_9771,N_8099,N_8344);
nor U9772 (N_9772,N_7674,N_8187);
and U9773 (N_9773,N_8999,N_8581);
nand U9774 (N_9774,N_8897,N_7559);
or U9775 (N_9775,N_7642,N_8252);
and U9776 (N_9776,N_8434,N_8794);
nand U9777 (N_9777,N_8826,N_8355);
or U9778 (N_9778,N_8222,N_8190);
nor U9779 (N_9779,N_8513,N_7618);
nand U9780 (N_9780,N_8240,N_8803);
or U9781 (N_9781,N_7554,N_8841);
and U9782 (N_9782,N_8412,N_8387);
and U9783 (N_9783,N_7501,N_8243);
nand U9784 (N_9784,N_8151,N_7633);
nor U9785 (N_9785,N_8505,N_8297);
or U9786 (N_9786,N_7844,N_7970);
or U9787 (N_9787,N_8433,N_8012);
and U9788 (N_9788,N_7868,N_8609);
nor U9789 (N_9789,N_8730,N_8758);
and U9790 (N_9790,N_7792,N_7513);
nor U9791 (N_9791,N_8818,N_8113);
nor U9792 (N_9792,N_7606,N_8854);
and U9793 (N_9793,N_7720,N_8422);
nand U9794 (N_9794,N_7576,N_8951);
xor U9795 (N_9795,N_7979,N_8187);
or U9796 (N_9796,N_7741,N_8129);
xnor U9797 (N_9797,N_7604,N_8513);
or U9798 (N_9798,N_8024,N_7858);
xnor U9799 (N_9799,N_8825,N_8040);
xnor U9800 (N_9800,N_8393,N_8464);
and U9801 (N_9801,N_7634,N_8089);
nor U9802 (N_9802,N_8782,N_7840);
nor U9803 (N_9803,N_7580,N_7729);
nor U9804 (N_9804,N_8340,N_8842);
or U9805 (N_9805,N_7569,N_7527);
and U9806 (N_9806,N_8858,N_7857);
nor U9807 (N_9807,N_7859,N_7651);
and U9808 (N_9808,N_7911,N_8679);
xor U9809 (N_9809,N_7530,N_7926);
and U9810 (N_9810,N_8808,N_8886);
nand U9811 (N_9811,N_8273,N_8967);
nor U9812 (N_9812,N_8971,N_7777);
or U9813 (N_9813,N_8247,N_8969);
and U9814 (N_9814,N_8186,N_8053);
nand U9815 (N_9815,N_8125,N_8725);
and U9816 (N_9816,N_7652,N_8002);
nor U9817 (N_9817,N_8960,N_8258);
nor U9818 (N_9818,N_8397,N_7954);
nor U9819 (N_9819,N_7615,N_8979);
xor U9820 (N_9820,N_7888,N_8791);
nand U9821 (N_9821,N_8225,N_8471);
and U9822 (N_9822,N_8585,N_7967);
or U9823 (N_9823,N_7957,N_8852);
or U9824 (N_9824,N_8915,N_8007);
nand U9825 (N_9825,N_8212,N_8258);
nor U9826 (N_9826,N_8464,N_7752);
nand U9827 (N_9827,N_8448,N_7862);
and U9828 (N_9828,N_8817,N_8265);
xnor U9829 (N_9829,N_8898,N_8491);
nand U9830 (N_9830,N_7544,N_7531);
and U9831 (N_9831,N_7898,N_7513);
nand U9832 (N_9832,N_8227,N_8623);
or U9833 (N_9833,N_8014,N_7536);
nor U9834 (N_9834,N_7553,N_7979);
nand U9835 (N_9835,N_8364,N_8037);
nand U9836 (N_9836,N_8127,N_7837);
nor U9837 (N_9837,N_8672,N_7837);
and U9838 (N_9838,N_7830,N_8090);
nand U9839 (N_9839,N_8895,N_7958);
nor U9840 (N_9840,N_8456,N_8793);
nor U9841 (N_9841,N_7932,N_8925);
and U9842 (N_9842,N_7739,N_7576);
nor U9843 (N_9843,N_7576,N_8171);
or U9844 (N_9844,N_7861,N_8868);
nor U9845 (N_9845,N_8320,N_8283);
and U9846 (N_9846,N_7542,N_7522);
nand U9847 (N_9847,N_7759,N_8288);
nand U9848 (N_9848,N_8928,N_8938);
nand U9849 (N_9849,N_8035,N_8383);
xor U9850 (N_9850,N_8836,N_7619);
and U9851 (N_9851,N_8401,N_8893);
xor U9852 (N_9852,N_8067,N_8549);
nor U9853 (N_9853,N_8695,N_7747);
xor U9854 (N_9854,N_8680,N_8668);
or U9855 (N_9855,N_7639,N_8510);
nor U9856 (N_9856,N_8378,N_8006);
or U9857 (N_9857,N_8031,N_7896);
nand U9858 (N_9858,N_8690,N_8618);
or U9859 (N_9859,N_8587,N_8524);
nand U9860 (N_9860,N_8935,N_8567);
xnor U9861 (N_9861,N_8980,N_7903);
nand U9862 (N_9862,N_7612,N_8354);
or U9863 (N_9863,N_7996,N_7891);
nor U9864 (N_9864,N_7711,N_8311);
or U9865 (N_9865,N_7691,N_8549);
nand U9866 (N_9866,N_8012,N_7659);
nand U9867 (N_9867,N_8477,N_7879);
and U9868 (N_9868,N_8871,N_8616);
or U9869 (N_9869,N_7654,N_8702);
and U9870 (N_9870,N_8972,N_8699);
nand U9871 (N_9871,N_7717,N_8296);
and U9872 (N_9872,N_7905,N_7829);
and U9873 (N_9873,N_7611,N_8024);
nor U9874 (N_9874,N_7589,N_8397);
nor U9875 (N_9875,N_7942,N_7702);
or U9876 (N_9876,N_8215,N_8382);
and U9877 (N_9877,N_8196,N_7692);
nand U9878 (N_9878,N_7709,N_7831);
nand U9879 (N_9879,N_7581,N_7757);
or U9880 (N_9880,N_7903,N_7852);
and U9881 (N_9881,N_7911,N_8905);
or U9882 (N_9882,N_7623,N_7548);
nor U9883 (N_9883,N_8825,N_7744);
nor U9884 (N_9884,N_7689,N_8701);
nor U9885 (N_9885,N_7819,N_8565);
and U9886 (N_9886,N_7501,N_8928);
nor U9887 (N_9887,N_8454,N_7607);
nand U9888 (N_9888,N_7833,N_7932);
or U9889 (N_9889,N_8906,N_8403);
nor U9890 (N_9890,N_8436,N_8840);
or U9891 (N_9891,N_8983,N_7827);
nor U9892 (N_9892,N_8711,N_8745);
nor U9893 (N_9893,N_8573,N_8650);
nand U9894 (N_9894,N_8886,N_8859);
nand U9895 (N_9895,N_8893,N_8667);
and U9896 (N_9896,N_8604,N_8509);
nand U9897 (N_9897,N_8858,N_8681);
or U9898 (N_9898,N_7677,N_7546);
or U9899 (N_9899,N_8035,N_8227);
nand U9900 (N_9900,N_8791,N_7771);
nor U9901 (N_9901,N_8057,N_8937);
nand U9902 (N_9902,N_7990,N_8502);
or U9903 (N_9903,N_7950,N_8525);
nand U9904 (N_9904,N_7633,N_8631);
nor U9905 (N_9905,N_8244,N_8512);
nand U9906 (N_9906,N_8786,N_7518);
and U9907 (N_9907,N_8411,N_8414);
nand U9908 (N_9908,N_8882,N_8432);
nor U9909 (N_9909,N_8535,N_8243);
or U9910 (N_9910,N_8495,N_8574);
nand U9911 (N_9911,N_8293,N_8306);
nand U9912 (N_9912,N_7628,N_8067);
xor U9913 (N_9913,N_7548,N_7775);
nand U9914 (N_9914,N_7737,N_8355);
nand U9915 (N_9915,N_8687,N_8111);
nand U9916 (N_9916,N_7565,N_8967);
and U9917 (N_9917,N_8426,N_7728);
and U9918 (N_9918,N_7676,N_8304);
nand U9919 (N_9919,N_7919,N_8027);
nand U9920 (N_9920,N_7913,N_7938);
or U9921 (N_9921,N_7603,N_8540);
and U9922 (N_9922,N_8479,N_8427);
nor U9923 (N_9923,N_7891,N_8558);
nor U9924 (N_9924,N_8987,N_8587);
nor U9925 (N_9925,N_8423,N_8412);
xnor U9926 (N_9926,N_8901,N_8002);
and U9927 (N_9927,N_7668,N_8363);
nand U9928 (N_9928,N_8042,N_7750);
and U9929 (N_9929,N_8893,N_7995);
and U9930 (N_9930,N_8391,N_8314);
nor U9931 (N_9931,N_8490,N_8959);
nor U9932 (N_9932,N_7771,N_8228);
or U9933 (N_9933,N_8715,N_7968);
or U9934 (N_9934,N_7726,N_7698);
nor U9935 (N_9935,N_7594,N_8241);
and U9936 (N_9936,N_8439,N_8310);
nand U9937 (N_9937,N_7835,N_8887);
or U9938 (N_9938,N_8788,N_8261);
nand U9939 (N_9939,N_8151,N_8278);
or U9940 (N_9940,N_8124,N_8776);
or U9941 (N_9941,N_8066,N_8108);
and U9942 (N_9942,N_8090,N_7806);
and U9943 (N_9943,N_8724,N_8587);
nor U9944 (N_9944,N_8940,N_7589);
nand U9945 (N_9945,N_7559,N_7573);
and U9946 (N_9946,N_8283,N_8809);
and U9947 (N_9947,N_8131,N_8304);
nor U9948 (N_9948,N_8679,N_8523);
or U9949 (N_9949,N_8934,N_8878);
and U9950 (N_9950,N_8759,N_7676);
nand U9951 (N_9951,N_8116,N_7841);
or U9952 (N_9952,N_7985,N_8419);
nor U9953 (N_9953,N_8383,N_8515);
and U9954 (N_9954,N_8071,N_8047);
nand U9955 (N_9955,N_7800,N_8277);
or U9956 (N_9956,N_8696,N_7738);
nand U9957 (N_9957,N_8103,N_8022);
and U9958 (N_9958,N_8177,N_7818);
or U9959 (N_9959,N_8190,N_8270);
and U9960 (N_9960,N_8582,N_8583);
xnor U9961 (N_9961,N_8645,N_7668);
or U9962 (N_9962,N_8746,N_7992);
nand U9963 (N_9963,N_8296,N_7690);
nand U9964 (N_9964,N_8076,N_7637);
nor U9965 (N_9965,N_7723,N_8448);
nand U9966 (N_9966,N_7533,N_8277);
or U9967 (N_9967,N_7992,N_8905);
or U9968 (N_9968,N_8392,N_8823);
and U9969 (N_9969,N_8937,N_8804);
and U9970 (N_9970,N_7834,N_8682);
nand U9971 (N_9971,N_7776,N_7663);
nand U9972 (N_9972,N_8510,N_8785);
and U9973 (N_9973,N_8784,N_7937);
nand U9974 (N_9974,N_7942,N_7743);
or U9975 (N_9975,N_8689,N_7732);
and U9976 (N_9976,N_7603,N_8429);
nor U9977 (N_9977,N_8304,N_7748);
xor U9978 (N_9978,N_8803,N_8572);
nor U9979 (N_9979,N_8428,N_8252);
and U9980 (N_9980,N_7789,N_8947);
nor U9981 (N_9981,N_8100,N_7707);
nor U9982 (N_9982,N_7771,N_8294);
and U9983 (N_9983,N_7764,N_8638);
or U9984 (N_9984,N_8643,N_8642);
nor U9985 (N_9985,N_8920,N_7874);
nand U9986 (N_9986,N_8256,N_7839);
nand U9987 (N_9987,N_8729,N_8986);
nor U9988 (N_9988,N_7732,N_8861);
nand U9989 (N_9989,N_7628,N_7511);
or U9990 (N_9990,N_8137,N_7823);
xnor U9991 (N_9991,N_7933,N_8741);
nand U9992 (N_9992,N_7603,N_8436);
xor U9993 (N_9993,N_7672,N_8407);
xnor U9994 (N_9994,N_7835,N_8249);
and U9995 (N_9995,N_7938,N_8681);
or U9996 (N_9996,N_8253,N_8490);
and U9997 (N_9997,N_8739,N_8620);
nor U9998 (N_9998,N_8328,N_8476);
nor U9999 (N_9999,N_7637,N_8298);
nand U10000 (N_10000,N_7545,N_7805);
nand U10001 (N_10001,N_8125,N_7773);
and U10002 (N_10002,N_8515,N_8394);
or U10003 (N_10003,N_8218,N_8664);
nor U10004 (N_10004,N_8226,N_7705);
nor U10005 (N_10005,N_8532,N_8477);
and U10006 (N_10006,N_7780,N_8392);
and U10007 (N_10007,N_8597,N_8523);
nor U10008 (N_10008,N_8470,N_8635);
nand U10009 (N_10009,N_8033,N_8857);
and U10010 (N_10010,N_8090,N_7754);
nor U10011 (N_10011,N_7869,N_8627);
nand U10012 (N_10012,N_8076,N_8896);
nor U10013 (N_10013,N_8970,N_7817);
nand U10014 (N_10014,N_8322,N_7845);
xnor U10015 (N_10015,N_8114,N_8000);
and U10016 (N_10016,N_8244,N_8069);
xnor U10017 (N_10017,N_8346,N_8296);
and U10018 (N_10018,N_8466,N_8294);
nand U10019 (N_10019,N_8475,N_7886);
or U10020 (N_10020,N_7788,N_7787);
or U10021 (N_10021,N_8021,N_8309);
or U10022 (N_10022,N_7814,N_8048);
xor U10023 (N_10023,N_7603,N_8732);
and U10024 (N_10024,N_7791,N_8483);
nor U10025 (N_10025,N_8622,N_7908);
xor U10026 (N_10026,N_8522,N_7704);
or U10027 (N_10027,N_7791,N_7644);
nor U10028 (N_10028,N_8717,N_8888);
nor U10029 (N_10029,N_8958,N_8383);
or U10030 (N_10030,N_8419,N_7846);
nor U10031 (N_10031,N_8303,N_8697);
nor U10032 (N_10032,N_7831,N_7840);
nor U10033 (N_10033,N_7933,N_8376);
nand U10034 (N_10034,N_8174,N_8918);
xor U10035 (N_10035,N_8211,N_8578);
nor U10036 (N_10036,N_8876,N_8925);
or U10037 (N_10037,N_7561,N_7855);
and U10038 (N_10038,N_7700,N_8402);
nor U10039 (N_10039,N_7751,N_8202);
xnor U10040 (N_10040,N_8690,N_8172);
nand U10041 (N_10041,N_8571,N_7652);
nor U10042 (N_10042,N_8787,N_7827);
xnor U10043 (N_10043,N_8415,N_8712);
nor U10044 (N_10044,N_8162,N_8547);
nand U10045 (N_10045,N_7858,N_7895);
and U10046 (N_10046,N_8173,N_8092);
nor U10047 (N_10047,N_8754,N_8504);
nor U10048 (N_10048,N_8730,N_8694);
or U10049 (N_10049,N_7911,N_7936);
nand U10050 (N_10050,N_7733,N_7584);
and U10051 (N_10051,N_8070,N_8600);
and U10052 (N_10052,N_8661,N_8342);
and U10053 (N_10053,N_8585,N_8360);
and U10054 (N_10054,N_8313,N_7677);
nand U10055 (N_10055,N_8237,N_8661);
and U10056 (N_10056,N_8893,N_8654);
nor U10057 (N_10057,N_7553,N_8233);
nor U10058 (N_10058,N_7570,N_8157);
xnor U10059 (N_10059,N_8995,N_8707);
nor U10060 (N_10060,N_7507,N_7985);
nand U10061 (N_10061,N_8581,N_7787);
or U10062 (N_10062,N_7823,N_7689);
nor U10063 (N_10063,N_7850,N_7806);
or U10064 (N_10064,N_7883,N_8274);
nand U10065 (N_10065,N_8360,N_8920);
or U10066 (N_10066,N_7969,N_8630);
nor U10067 (N_10067,N_8737,N_8164);
nand U10068 (N_10068,N_7639,N_7673);
nor U10069 (N_10069,N_8527,N_7991);
nand U10070 (N_10070,N_8207,N_8335);
and U10071 (N_10071,N_8898,N_8433);
nor U10072 (N_10072,N_8487,N_8167);
or U10073 (N_10073,N_8778,N_7906);
nand U10074 (N_10074,N_8858,N_8943);
nand U10075 (N_10075,N_7718,N_8462);
and U10076 (N_10076,N_7721,N_8319);
and U10077 (N_10077,N_7553,N_8263);
and U10078 (N_10078,N_7681,N_8180);
nor U10079 (N_10079,N_8725,N_7716);
and U10080 (N_10080,N_8930,N_8013);
nor U10081 (N_10081,N_8359,N_8962);
xnor U10082 (N_10082,N_8084,N_8828);
nor U10083 (N_10083,N_8709,N_7907);
nor U10084 (N_10084,N_7974,N_8394);
or U10085 (N_10085,N_8159,N_7974);
and U10086 (N_10086,N_8351,N_8117);
and U10087 (N_10087,N_8948,N_8789);
and U10088 (N_10088,N_8265,N_8615);
nor U10089 (N_10089,N_8452,N_8749);
nand U10090 (N_10090,N_7930,N_8267);
or U10091 (N_10091,N_7976,N_7987);
and U10092 (N_10092,N_8475,N_8218);
or U10093 (N_10093,N_8058,N_8002);
nor U10094 (N_10094,N_8777,N_7663);
and U10095 (N_10095,N_7780,N_8923);
nor U10096 (N_10096,N_7605,N_7936);
or U10097 (N_10097,N_8841,N_8308);
and U10098 (N_10098,N_7795,N_8541);
and U10099 (N_10099,N_8772,N_8506);
or U10100 (N_10100,N_8567,N_7615);
nand U10101 (N_10101,N_8079,N_8289);
and U10102 (N_10102,N_7679,N_8388);
and U10103 (N_10103,N_8964,N_8734);
nand U10104 (N_10104,N_7547,N_8595);
and U10105 (N_10105,N_8081,N_8344);
nor U10106 (N_10106,N_7557,N_8004);
and U10107 (N_10107,N_8501,N_8410);
nand U10108 (N_10108,N_7819,N_7880);
nor U10109 (N_10109,N_7895,N_8754);
and U10110 (N_10110,N_7574,N_8764);
nor U10111 (N_10111,N_7565,N_8748);
xnor U10112 (N_10112,N_8853,N_8062);
or U10113 (N_10113,N_8551,N_7855);
nand U10114 (N_10114,N_8250,N_8882);
and U10115 (N_10115,N_8115,N_8271);
or U10116 (N_10116,N_8091,N_8461);
and U10117 (N_10117,N_7717,N_8793);
nor U10118 (N_10118,N_8320,N_7794);
and U10119 (N_10119,N_7898,N_8917);
and U10120 (N_10120,N_8966,N_8128);
nand U10121 (N_10121,N_8032,N_8165);
nand U10122 (N_10122,N_8224,N_7727);
nor U10123 (N_10123,N_8729,N_8894);
and U10124 (N_10124,N_8137,N_7710);
or U10125 (N_10125,N_8148,N_7658);
nand U10126 (N_10126,N_8446,N_8251);
and U10127 (N_10127,N_7680,N_8529);
nand U10128 (N_10128,N_7732,N_8362);
and U10129 (N_10129,N_7773,N_7588);
nand U10130 (N_10130,N_7755,N_8542);
and U10131 (N_10131,N_8546,N_8568);
or U10132 (N_10132,N_7511,N_8888);
and U10133 (N_10133,N_7698,N_7683);
and U10134 (N_10134,N_7873,N_8311);
and U10135 (N_10135,N_7634,N_8991);
nor U10136 (N_10136,N_7745,N_7591);
or U10137 (N_10137,N_8477,N_8909);
xor U10138 (N_10138,N_7673,N_8255);
nand U10139 (N_10139,N_8443,N_7542);
or U10140 (N_10140,N_8925,N_8479);
or U10141 (N_10141,N_8879,N_7654);
and U10142 (N_10142,N_7672,N_8476);
nor U10143 (N_10143,N_8453,N_8356);
nand U10144 (N_10144,N_7613,N_8834);
nand U10145 (N_10145,N_8334,N_8258);
or U10146 (N_10146,N_8173,N_8819);
xnor U10147 (N_10147,N_7553,N_8626);
nor U10148 (N_10148,N_8985,N_7937);
or U10149 (N_10149,N_8566,N_8564);
nor U10150 (N_10150,N_7609,N_8312);
nand U10151 (N_10151,N_8330,N_8069);
or U10152 (N_10152,N_7845,N_8042);
nor U10153 (N_10153,N_7883,N_7554);
nor U10154 (N_10154,N_8829,N_7948);
and U10155 (N_10155,N_8322,N_8272);
nor U10156 (N_10156,N_8715,N_7727);
and U10157 (N_10157,N_7696,N_8679);
and U10158 (N_10158,N_8999,N_8517);
nand U10159 (N_10159,N_8757,N_8563);
nor U10160 (N_10160,N_8905,N_8093);
or U10161 (N_10161,N_8357,N_8927);
or U10162 (N_10162,N_8380,N_8167);
and U10163 (N_10163,N_7676,N_8043);
nor U10164 (N_10164,N_8792,N_8233);
nand U10165 (N_10165,N_7965,N_8625);
and U10166 (N_10166,N_8908,N_8291);
nor U10167 (N_10167,N_8703,N_7533);
nand U10168 (N_10168,N_7525,N_8705);
xnor U10169 (N_10169,N_8805,N_8699);
nor U10170 (N_10170,N_8250,N_8361);
and U10171 (N_10171,N_8563,N_8264);
or U10172 (N_10172,N_8308,N_8290);
and U10173 (N_10173,N_7645,N_8645);
and U10174 (N_10174,N_7774,N_8131);
or U10175 (N_10175,N_7505,N_8347);
nor U10176 (N_10176,N_8192,N_8759);
or U10177 (N_10177,N_7727,N_8484);
nand U10178 (N_10178,N_8689,N_8421);
nand U10179 (N_10179,N_7768,N_8778);
or U10180 (N_10180,N_8768,N_8706);
nor U10181 (N_10181,N_8497,N_7933);
nor U10182 (N_10182,N_7951,N_8764);
xnor U10183 (N_10183,N_7983,N_8275);
and U10184 (N_10184,N_8607,N_7871);
nor U10185 (N_10185,N_7728,N_8107);
nor U10186 (N_10186,N_8827,N_8632);
and U10187 (N_10187,N_7619,N_7924);
or U10188 (N_10188,N_7593,N_7833);
nor U10189 (N_10189,N_8216,N_7546);
xnor U10190 (N_10190,N_8988,N_7515);
and U10191 (N_10191,N_8697,N_8606);
nand U10192 (N_10192,N_7929,N_8042);
and U10193 (N_10193,N_7977,N_8732);
nor U10194 (N_10194,N_8599,N_8479);
nor U10195 (N_10195,N_8228,N_8996);
and U10196 (N_10196,N_7522,N_8826);
nor U10197 (N_10197,N_7752,N_8056);
nand U10198 (N_10198,N_8198,N_8967);
and U10199 (N_10199,N_8234,N_7882);
or U10200 (N_10200,N_8643,N_8723);
nand U10201 (N_10201,N_7749,N_8464);
nor U10202 (N_10202,N_8112,N_8419);
xor U10203 (N_10203,N_8839,N_8760);
xnor U10204 (N_10204,N_7954,N_8936);
xnor U10205 (N_10205,N_8376,N_8941);
xor U10206 (N_10206,N_8376,N_8886);
nand U10207 (N_10207,N_7960,N_7824);
and U10208 (N_10208,N_7781,N_7663);
and U10209 (N_10209,N_7800,N_8606);
nand U10210 (N_10210,N_8693,N_7515);
nor U10211 (N_10211,N_7578,N_8939);
and U10212 (N_10212,N_7883,N_7614);
xnor U10213 (N_10213,N_7836,N_8795);
nand U10214 (N_10214,N_8240,N_8205);
xnor U10215 (N_10215,N_7705,N_8461);
or U10216 (N_10216,N_8819,N_8028);
and U10217 (N_10217,N_8189,N_7991);
or U10218 (N_10218,N_7887,N_8562);
and U10219 (N_10219,N_8346,N_7668);
and U10220 (N_10220,N_8917,N_8923);
nor U10221 (N_10221,N_7545,N_8362);
nand U10222 (N_10222,N_7509,N_7674);
nor U10223 (N_10223,N_7975,N_8357);
nor U10224 (N_10224,N_8306,N_8850);
and U10225 (N_10225,N_7822,N_8973);
and U10226 (N_10226,N_8946,N_8410);
or U10227 (N_10227,N_8821,N_7518);
or U10228 (N_10228,N_8153,N_7976);
and U10229 (N_10229,N_7557,N_7783);
nand U10230 (N_10230,N_8932,N_7970);
nand U10231 (N_10231,N_7844,N_7950);
and U10232 (N_10232,N_8306,N_8852);
nor U10233 (N_10233,N_8400,N_8235);
or U10234 (N_10234,N_8807,N_7593);
nor U10235 (N_10235,N_7782,N_8389);
nor U10236 (N_10236,N_7823,N_8954);
nand U10237 (N_10237,N_7527,N_8837);
nand U10238 (N_10238,N_7784,N_8477);
nand U10239 (N_10239,N_8285,N_8342);
nand U10240 (N_10240,N_8930,N_7533);
or U10241 (N_10241,N_8959,N_7942);
and U10242 (N_10242,N_8829,N_7966);
nand U10243 (N_10243,N_8286,N_8653);
or U10244 (N_10244,N_7614,N_8743);
and U10245 (N_10245,N_8554,N_7940);
and U10246 (N_10246,N_7846,N_8590);
or U10247 (N_10247,N_8891,N_8451);
and U10248 (N_10248,N_7934,N_7557);
or U10249 (N_10249,N_7948,N_7711);
nand U10250 (N_10250,N_7699,N_8175);
or U10251 (N_10251,N_8856,N_8731);
and U10252 (N_10252,N_7730,N_8683);
nand U10253 (N_10253,N_7554,N_7932);
nor U10254 (N_10254,N_7875,N_7596);
nand U10255 (N_10255,N_7795,N_8110);
nand U10256 (N_10256,N_8095,N_8107);
nor U10257 (N_10257,N_7788,N_8058);
nor U10258 (N_10258,N_7899,N_8479);
nand U10259 (N_10259,N_7900,N_8702);
and U10260 (N_10260,N_8119,N_8534);
xor U10261 (N_10261,N_8423,N_8251);
nor U10262 (N_10262,N_7903,N_8516);
or U10263 (N_10263,N_8303,N_8465);
or U10264 (N_10264,N_7933,N_8243);
or U10265 (N_10265,N_8715,N_8106);
nand U10266 (N_10266,N_7659,N_8046);
or U10267 (N_10267,N_8495,N_8909);
nand U10268 (N_10268,N_8138,N_8555);
or U10269 (N_10269,N_7945,N_8990);
and U10270 (N_10270,N_8635,N_7758);
xor U10271 (N_10271,N_7708,N_7845);
or U10272 (N_10272,N_7973,N_7641);
or U10273 (N_10273,N_8647,N_8535);
xnor U10274 (N_10274,N_8096,N_8619);
nand U10275 (N_10275,N_7884,N_8017);
nor U10276 (N_10276,N_8363,N_7782);
and U10277 (N_10277,N_8361,N_8385);
nand U10278 (N_10278,N_7646,N_8597);
or U10279 (N_10279,N_8734,N_8864);
or U10280 (N_10280,N_7571,N_7917);
xor U10281 (N_10281,N_8151,N_8550);
and U10282 (N_10282,N_7895,N_8099);
and U10283 (N_10283,N_7543,N_8140);
and U10284 (N_10284,N_7795,N_8608);
nand U10285 (N_10285,N_8139,N_8852);
nand U10286 (N_10286,N_7801,N_7881);
nand U10287 (N_10287,N_7766,N_8030);
or U10288 (N_10288,N_8211,N_7865);
and U10289 (N_10289,N_7914,N_8391);
nor U10290 (N_10290,N_8876,N_8797);
or U10291 (N_10291,N_8528,N_7957);
or U10292 (N_10292,N_8597,N_8577);
nor U10293 (N_10293,N_8739,N_8812);
nor U10294 (N_10294,N_7705,N_7782);
or U10295 (N_10295,N_8101,N_8234);
and U10296 (N_10296,N_8330,N_8842);
xor U10297 (N_10297,N_8509,N_8558);
nand U10298 (N_10298,N_7950,N_8555);
or U10299 (N_10299,N_8739,N_8881);
nand U10300 (N_10300,N_7855,N_8339);
and U10301 (N_10301,N_7920,N_7615);
nand U10302 (N_10302,N_8738,N_8750);
or U10303 (N_10303,N_8886,N_8489);
and U10304 (N_10304,N_8380,N_8140);
nor U10305 (N_10305,N_7668,N_8129);
and U10306 (N_10306,N_8657,N_8946);
or U10307 (N_10307,N_8796,N_8482);
nand U10308 (N_10308,N_8330,N_7777);
nor U10309 (N_10309,N_7951,N_8184);
nor U10310 (N_10310,N_7630,N_8662);
and U10311 (N_10311,N_8265,N_8587);
and U10312 (N_10312,N_7767,N_7818);
and U10313 (N_10313,N_8948,N_7919);
nand U10314 (N_10314,N_8406,N_7928);
or U10315 (N_10315,N_8809,N_8030);
or U10316 (N_10316,N_8671,N_8943);
and U10317 (N_10317,N_7588,N_7889);
nor U10318 (N_10318,N_8033,N_7822);
nor U10319 (N_10319,N_7741,N_8653);
nand U10320 (N_10320,N_8629,N_8959);
and U10321 (N_10321,N_8982,N_8543);
nor U10322 (N_10322,N_8761,N_8422);
or U10323 (N_10323,N_8584,N_8117);
and U10324 (N_10324,N_8737,N_7840);
nand U10325 (N_10325,N_8233,N_8348);
or U10326 (N_10326,N_8118,N_7851);
nand U10327 (N_10327,N_8456,N_8167);
and U10328 (N_10328,N_8956,N_7702);
or U10329 (N_10329,N_7822,N_8551);
and U10330 (N_10330,N_7535,N_8692);
xnor U10331 (N_10331,N_7972,N_7822);
or U10332 (N_10332,N_8000,N_8579);
xor U10333 (N_10333,N_8606,N_8155);
xnor U10334 (N_10334,N_8844,N_8079);
or U10335 (N_10335,N_7943,N_8917);
nor U10336 (N_10336,N_7861,N_7788);
nor U10337 (N_10337,N_7817,N_8489);
or U10338 (N_10338,N_8411,N_8236);
or U10339 (N_10339,N_8621,N_7604);
or U10340 (N_10340,N_7935,N_7872);
nand U10341 (N_10341,N_8440,N_8234);
xor U10342 (N_10342,N_8677,N_8478);
or U10343 (N_10343,N_8550,N_8682);
nor U10344 (N_10344,N_8322,N_7561);
and U10345 (N_10345,N_7777,N_7976);
and U10346 (N_10346,N_8510,N_8143);
and U10347 (N_10347,N_8063,N_8581);
and U10348 (N_10348,N_7588,N_8414);
nor U10349 (N_10349,N_8174,N_8092);
and U10350 (N_10350,N_8939,N_8294);
or U10351 (N_10351,N_7539,N_8217);
xor U10352 (N_10352,N_7634,N_8452);
nor U10353 (N_10353,N_8938,N_7993);
xor U10354 (N_10354,N_8898,N_7645);
nand U10355 (N_10355,N_7996,N_7875);
nor U10356 (N_10356,N_8914,N_7516);
nand U10357 (N_10357,N_8278,N_8722);
nand U10358 (N_10358,N_8927,N_8421);
nor U10359 (N_10359,N_8328,N_8300);
and U10360 (N_10360,N_7822,N_8304);
nand U10361 (N_10361,N_7779,N_8323);
nand U10362 (N_10362,N_8368,N_7758);
or U10363 (N_10363,N_7592,N_8819);
or U10364 (N_10364,N_7852,N_7632);
nor U10365 (N_10365,N_8186,N_7509);
nand U10366 (N_10366,N_7559,N_7560);
nand U10367 (N_10367,N_7850,N_8886);
and U10368 (N_10368,N_8064,N_7963);
nand U10369 (N_10369,N_7609,N_8564);
nor U10370 (N_10370,N_7932,N_8921);
xnor U10371 (N_10371,N_8203,N_8954);
or U10372 (N_10372,N_8360,N_7942);
xnor U10373 (N_10373,N_8045,N_8398);
or U10374 (N_10374,N_7919,N_7960);
nand U10375 (N_10375,N_7550,N_8183);
or U10376 (N_10376,N_7665,N_7993);
xor U10377 (N_10377,N_8343,N_8100);
nor U10378 (N_10378,N_7998,N_8454);
nand U10379 (N_10379,N_8859,N_8906);
or U10380 (N_10380,N_8935,N_7865);
and U10381 (N_10381,N_7707,N_8212);
and U10382 (N_10382,N_8432,N_8263);
and U10383 (N_10383,N_7928,N_8571);
nand U10384 (N_10384,N_8863,N_8259);
nor U10385 (N_10385,N_8219,N_8923);
and U10386 (N_10386,N_7890,N_7657);
nand U10387 (N_10387,N_7828,N_7820);
and U10388 (N_10388,N_8695,N_8875);
and U10389 (N_10389,N_8981,N_8895);
or U10390 (N_10390,N_8006,N_8385);
and U10391 (N_10391,N_7809,N_8409);
nor U10392 (N_10392,N_7757,N_8567);
xnor U10393 (N_10393,N_7604,N_8054);
and U10394 (N_10394,N_7783,N_7678);
and U10395 (N_10395,N_8212,N_7606);
or U10396 (N_10396,N_8771,N_7906);
nand U10397 (N_10397,N_8905,N_8263);
nand U10398 (N_10398,N_8713,N_7600);
xnor U10399 (N_10399,N_8706,N_8736);
nor U10400 (N_10400,N_8492,N_7917);
xnor U10401 (N_10401,N_8612,N_8026);
and U10402 (N_10402,N_8732,N_7841);
xnor U10403 (N_10403,N_8320,N_7501);
nand U10404 (N_10404,N_7866,N_8287);
xor U10405 (N_10405,N_7983,N_7594);
nor U10406 (N_10406,N_7518,N_8910);
or U10407 (N_10407,N_7890,N_8737);
nand U10408 (N_10408,N_7645,N_8234);
nand U10409 (N_10409,N_7927,N_8178);
or U10410 (N_10410,N_8110,N_8948);
and U10411 (N_10411,N_8597,N_8413);
nor U10412 (N_10412,N_8869,N_8934);
nand U10413 (N_10413,N_8478,N_8382);
nand U10414 (N_10414,N_8240,N_7706);
xor U10415 (N_10415,N_8995,N_8146);
xnor U10416 (N_10416,N_8812,N_7556);
nor U10417 (N_10417,N_7900,N_8561);
nor U10418 (N_10418,N_7960,N_8001);
and U10419 (N_10419,N_8356,N_8674);
or U10420 (N_10420,N_7901,N_8374);
nor U10421 (N_10421,N_8420,N_7897);
and U10422 (N_10422,N_8619,N_8012);
nor U10423 (N_10423,N_7613,N_8727);
nand U10424 (N_10424,N_8757,N_7660);
or U10425 (N_10425,N_7945,N_8432);
nand U10426 (N_10426,N_7616,N_8517);
nand U10427 (N_10427,N_8962,N_8546);
and U10428 (N_10428,N_8921,N_8097);
xnor U10429 (N_10429,N_8513,N_7593);
and U10430 (N_10430,N_7733,N_7667);
and U10431 (N_10431,N_8320,N_8326);
nor U10432 (N_10432,N_8045,N_8882);
or U10433 (N_10433,N_8438,N_8607);
nand U10434 (N_10434,N_8483,N_8141);
or U10435 (N_10435,N_8181,N_8407);
nand U10436 (N_10436,N_8338,N_7714);
or U10437 (N_10437,N_8450,N_7712);
xnor U10438 (N_10438,N_7613,N_7625);
and U10439 (N_10439,N_8518,N_8564);
and U10440 (N_10440,N_8426,N_8999);
and U10441 (N_10441,N_8776,N_8259);
or U10442 (N_10442,N_8754,N_8835);
nand U10443 (N_10443,N_8149,N_8924);
and U10444 (N_10444,N_8028,N_7805);
nand U10445 (N_10445,N_8595,N_8358);
nand U10446 (N_10446,N_7607,N_7520);
and U10447 (N_10447,N_8762,N_7641);
and U10448 (N_10448,N_8774,N_7516);
and U10449 (N_10449,N_7617,N_8725);
or U10450 (N_10450,N_7866,N_7923);
and U10451 (N_10451,N_8482,N_8004);
or U10452 (N_10452,N_8665,N_8351);
or U10453 (N_10453,N_8127,N_8574);
and U10454 (N_10454,N_8292,N_8813);
xnor U10455 (N_10455,N_8933,N_7834);
or U10456 (N_10456,N_8504,N_8679);
and U10457 (N_10457,N_7703,N_7537);
and U10458 (N_10458,N_8221,N_7994);
nand U10459 (N_10459,N_7743,N_8233);
xnor U10460 (N_10460,N_7769,N_7670);
nand U10461 (N_10461,N_8298,N_7855);
nor U10462 (N_10462,N_7943,N_7546);
nand U10463 (N_10463,N_8658,N_8895);
or U10464 (N_10464,N_8803,N_8396);
nand U10465 (N_10465,N_8210,N_7594);
nor U10466 (N_10466,N_8650,N_8964);
nor U10467 (N_10467,N_8907,N_8905);
or U10468 (N_10468,N_8273,N_8251);
nand U10469 (N_10469,N_8027,N_8955);
xnor U10470 (N_10470,N_8822,N_8424);
nor U10471 (N_10471,N_8709,N_7745);
nand U10472 (N_10472,N_8572,N_7942);
nor U10473 (N_10473,N_8096,N_7981);
nor U10474 (N_10474,N_8023,N_8458);
nor U10475 (N_10475,N_8200,N_8749);
nor U10476 (N_10476,N_8149,N_8601);
nand U10477 (N_10477,N_8270,N_8094);
nand U10478 (N_10478,N_8821,N_8974);
and U10479 (N_10479,N_7668,N_7725);
nand U10480 (N_10480,N_8737,N_8113);
nand U10481 (N_10481,N_8997,N_8270);
or U10482 (N_10482,N_8319,N_7928);
nand U10483 (N_10483,N_7652,N_8708);
nor U10484 (N_10484,N_7684,N_8925);
and U10485 (N_10485,N_7645,N_7755);
and U10486 (N_10486,N_8334,N_8255);
xor U10487 (N_10487,N_8195,N_7715);
nand U10488 (N_10488,N_8388,N_8843);
or U10489 (N_10489,N_8936,N_7857);
or U10490 (N_10490,N_8962,N_8506);
or U10491 (N_10491,N_8733,N_8480);
nand U10492 (N_10492,N_8822,N_7664);
nor U10493 (N_10493,N_7553,N_8569);
nor U10494 (N_10494,N_8040,N_7653);
nand U10495 (N_10495,N_8841,N_8074);
xnor U10496 (N_10496,N_8415,N_8982);
or U10497 (N_10497,N_7739,N_8506);
nor U10498 (N_10498,N_8273,N_8423);
xor U10499 (N_10499,N_8248,N_8825);
and U10500 (N_10500,N_9336,N_10471);
or U10501 (N_10501,N_9866,N_9019);
nand U10502 (N_10502,N_9579,N_9879);
xnor U10503 (N_10503,N_9631,N_10214);
and U10504 (N_10504,N_9832,N_10274);
or U10505 (N_10505,N_9556,N_9968);
nor U10506 (N_10506,N_9238,N_9734);
nand U10507 (N_10507,N_9739,N_9725);
nor U10508 (N_10508,N_9784,N_9664);
nor U10509 (N_10509,N_10244,N_9954);
nor U10510 (N_10510,N_9256,N_9440);
nand U10511 (N_10511,N_10251,N_9768);
and U10512 (N_10512,N_9048,N_9073);
nand U10513 (N_10513,N_10459,N_9609);
nand U10514 (N_10514,N_9641,N_9358);
or U10515 (N_10515,N_9466,N_9471);
or U10516 (N_10516,N_9240,N_10106);
xnor U10517 (N_10517,N_9665,N_9117);
nand U10518 (N_10518,N_9920,N_10256);
or U10519 (N_10519,N_9895,N_9494);
or U10520 (N_10520,N_9771,N_9708);
nor U10521 (N_10521,N_9165,N_10301);
nand U10522 (N_10522,N_9961,N_9473);
or U10523 (N_10523,N_9476,N_10325);
and U10524 (N_10524,N_9865,N_9569);
xnor U10525 (N_10525,N_9421,N_9963);
or U10526 (N_10526,N_10454,N_9026);
nor U10527 (N_10527,N_10169,N_9166);
nand U10528 (N_10528,N_10289,N_9416);
xnor U10529 (N_10529,N_9228,N_9255);
nand U10530 (N_10530,N_10223,N_9382);
xnor U10531 (N_10531,N_10424,N_9842);
or U10532 (N_10532,N_10047,N_9905);
nand U10533 (N_10533,N_9332,N_9044);
nand U10534 (N_10534,N_9038,N_9550);
nand U10535 (N_10535,N_9847,N_9236);
nor U10536 (N_10536,N_10347,N_9386);
nor U10537 (N_10537,N_9521,N_9083);
and U10538 (N_10538,N_9069,N_10282);
and U10539 (N_10539,N_9567,N_9837);
nand U10540 (N_10540,N_9425,N_9225);
nand U10541 (N_10541,N_10233,N_10364);
or U10542 (N_10542,N_9356,N_10401);
and U10543 (N_10543,N_9046,N_9405);
nor U10544 (N_10544,N_9605,N_9681);
xor U10545 (N_10545,N_10015,N_9156);
nand U10546 (N_10546,N_10435,N_9642);
nor U10547 (N_10547,N_9796,N_10438);
xnor U10548 (N_10548,N_9029,N_9031);
nor U10549 (N_10549,N_9063,N_9179);
and U10550 (N_10550,N_10068,N_9115);
nand U10551 (N_10551,N_10010,N_10283);
nand U10552 (N_10552,N_9946,N_9705);
nor U10553 (N_10553,N_9505,N_9517);
and U10554 (N_10554,N_9318,N_9120);
and U10555 (N_10555,N_9619,N_9223);
or U10556 (N_10556,N_9608,N_9465);
or U10557 (N_10557,N_9911,N_10292);
nand U10558 (N_10558,N_10490,N_9673);
or U10559 (N_10559,N_9390,N_9180);
or U10560 (N_10560,N_10241,N_9452);
or U10561 (N_10561,N_10120,N_10036);
nand U10562 (N_10562,N_9343,N_9350);
nand U10563 (N_10563,N_10048,N_9001);
nor U10564 (N_10564,N_9052,N_9259);
and U10565 (N_10565,N_9366,N_9597);
xnor U10566 (N_10566,N_9246,N_9233);
nor U10567 (N_10567,N_9629,N_9980);
or U10568 (N_10568,N_9338,N_9906);
and U10569 (N_10569,N_9330,N_10387);
or U10570 (N_10570,N_9649,N_10207);
nand U10571 (N_10571,N_9838,N_10163);
nand U10572 (N_10572,N_9174,N_9772);
xor U10573 (N_10573,N_10226,N_9541);
xnor U10574 (N_10574,N_9245,N_9017);
or U10575 (N_10575,N_10349,N_9387);
nor U10576 (N_10576,N_9827,N_10136);
nand U10577 (N_10577,N_10412,N_9442);
or U10578 (N_10578,N_9388,N_9977);
or U10579 (N_10579,N_9348,N_10185);
and U10580 (N_10580,N_9765,N_10477);
nor U10581 (N_10581,N_9430,N_10208);
nor U10582 (N_10582,N_10137,N_9474);
nand U10583 (N_10583,N_9939,N_10383);
or U10584 (N_10584,N_9114,N_9930);
xnor U10585 (N_10585,N_10355,N_9721);
and U10586 (N_10586,N_9902,N_9798);
nand U10587 (N_10587,N_9116,N_9611);
or U10588 (N_10588,N_10452,N_10055);
or U10589 (N_10589,N_9532,N_9242);
and U10590 (N_10590,N_9874,N_10118);
or U10591 (N_10591,N_9652,N_10427);
or U10592 (N_10592,N_10162,N_9620);
nand U10593 (N_10593,N_9250,N_10171);
nor U10594 (N_10594,N_9834,N_9081);
and U10595 (N_10595,N_10252,N_9618);
or U10596 (N_10596,N_9817,N_9821);
nand U10597 (N_10597,N_10455,N_9668);
or U10598 (N_10598,N_9857,N_9551);
nand U10599 (N_10599,N_9660,N_10192);
and U10600 (N_10600,N_10377,N_9185);
nand U10601 (N_10601,N_10307,N_9365);
or U10602 (N_10602,N_9970,N_9995);
nor U10603 (N_10603,N_10385,N_10341);
nor U10604 (N_10604,N_9441,N_10371);
and U10605 (N_10605,N_9379,N_10458);
or U10606 (N_10606,N_9923,N_9011);
nand U10607 (N_10607,N_10020,N_9399);
or U10608 (N_10608,N_9422,N_9484);
or U10609 (N_10609,N_9058,N_9858);
or U10610 (N_10610,N_9751,N_9310);
nor U10611 (N_10611,N_9791,N_10187);
or U10612 (N_10612,N_9439,N_10317);
or U10613 (N_10613,N_9105,N_10013);
or U10614 (N_10614,N_9919,N_10413);
and U10615 (N_10615,N_10161,N_9713);
and U10616 (N_10616,N_9186,N_9720);
and U10617 (N_10617,N_9872,N_9519);
or U10618 (N_10618,N_9061,N_9621);
and U10619 (N_10619,N_9414,N_9363);
xnor U10620 (N_10620,N_10021,N_9984);
nand U10621 (N_10621,N_10416,N_10132);
nor U10622 (N_10622,N_10334,N_9459);
nand U10623 (N_10623,N_10038,N_9071);
xor U10624 (N_10624,N_9764,N_10276);
or U10625 (N_10625,N_9632,N_9131);
or U10626 (N_10626,N_10428,N_10291);
nand U10627 (N_10627,N_10141,N_9563);
and U10628 (N_10628,N_9126,N_10303);
or U10629 (N_10629,N_10176,N_9106);
and U10630 (N_10630,N_10417,N_9633);
and U10631 (N_10631,N_10462,N_10243);
xnor U10632 (N_10632,N_9757,N_9364);
nand U10633 (N_10633,N_10389,N_10017);
and U10634 (N_10634,N_10343,N_9202);
nor U10635 (N_10635,N_9010,N_9997);
and U10636 (N_10636,N_9333,N_10384);
xor U10637 (N_10637,N_9254,N_9819);
nand U10638 (N_10638,N_9941,N_9004);
nand U10639 (N_10639,N_9142,N_10296);
nand U10640 (N_10640,N_10114,N_10356);
and U10641 (N_10641,N_10150,N_9362);
nor U10642 (N_10642,N_9731,N_9136);
nor U10643 (N_10643,N_9592,N_9373);
nand U10644 (N_10644,N_9215,N_10368);
or U10645 (N_10645,N_10367,N_10103);
nor U10646 (N_10646,N_9952,N_10066);
nor U10647 (N_10647,N_10202,N_10085);
nor U10648 (N_10648,N_10255,N_10016);
nor U10649 (N_10649,N_9098,N_9357);
xor U10650 (N_10650,N_9220,N_9654);
or U10651 (N_10651,N_9801,N_9383);
nor U10652 (N_10652,N_10219,N_10441);
and U10653 (N_10653,N_9637,N_9320);
nor U10654 (N_10654,N_9525,N_10266);
nor U10655 (N_10655,N_9898,N_9848);
or U10656 (N_10656,N_10045,N_9773);
xnor U10657 (N_10657,N_10101,N_10331);
nand U10658 (N_10658,N_10306,N_9229);
or U10659 (N_10659,N_9193,N_9710);
nand U10660 (N_10660,N_10362,N_10026);
nor U10661 (N_10661,N_10059,N_10105);
or U10662 (N_10662,N_10180,N_9475);
nor U10663 (N_10663,N_9574,N_9989);
nand U10664 (N_10664,N_9758,N_9403);
nor U10665 (N_10665,N_9045,N_9682);
nand U10666 (N_10666,N_9119,N_9750);
nor U10667 (N_10667,N_9639,N_10311);
or U10668 (N_10668,N_10472,N_9538);
nand U10669 (N_10669,N_10145,N_10217);
or U10670 (N_10670,N_10193,N_9766);
or U10671 (N_10671,N_9511,N_9337);
and U10672 (N_10672,N_9210,N_10314);
nor U10673 (N_10673,N_9718,N_10351);
nor U10674 (N_10674,N_9717,N_10337);
and U10675 (N_10675,N_9743,N_9354);
or U10676 (N_10676,N_9341,N_9149);
nand U10677 (N_10677,N_10155,N_9786);
nor U10678 (N_10678,N_10468,N_10429);
nand U10679 (N_10679,N_9581,N_9938);
or U10680 (N_10680,N_10405,N_10353);
nor U10681 (N_10681,N_9445,N_10330);
or U10682 (N_10682,N_9566,N_9686);
nand U10683 (N_10683,N_9868,N_9839);
nand U10684 (N_10684,N_9962,N_9985);
nor U10685 (N_10685,N_10445,N_9864);
nand U10686 (N_10686,N_10422,N_10482);
nor U10687 (N_10687,N_9092,N_9630);
or U10688 (N_10688,N_9303,N_9510);
and U10689 (N_10689,N_9378,N_9959);
nand U10690 (N_10690,N_9804,N_9208);
or U10691 (N_10691,N_9127,N_9507);
xor U10692 (N_10692,N_9779,N_10135);
nand U10693 (N_10693,N_10300,N_9072);
or U10694 (N_10694,N_9600,N_9109);
nand U10695 (N_10695,N_9774,N_10222);
or U10696 (N_10696,N_9204,N_9575);
and U10697 (N_10697,N_9509,N_9040);
nand U10698 (N_10698,N_10061,N_9643);
nand U10699 (N_10699,N_9716,N_9807);
or U10700 (N_10700,N_9896,N_9122);
and U10701 (N_10701,N_9340,N_9368);
nand U10702 (N_10702,N_9535,N_9274);
xnor U10703 (N_10703,N_10234,N_9140);
nor U10704 (N_10704,N_10495,N_9129);
nor U10705 (N_10705,N_9392,N_9900);
nor U10706 (N_10706,N_10130,N_10324);
xor U10707 (N_10707,N_9955,N_10464);
xor U10708 (N_10708,N_9612,N_10277);
or U10709 (N_10709,N_9104,N_9576);
and U10710 (N_10710,N_10081,N_9822);
nand U10711 (N_10711,N_9329,N_10379);
and U10712 (N_10712,N_9737,N_10295);
and U10713 (N_10713,N_9559,N_9171);
or U10714 (N_10714,N_9391,N_10370);
nand U10715 (N_10715,N_10211,N_9467);
or U10716 (N_10716,N_10000,N_9647);
nor U10717 (N_10717,N_9323,N_10394);
and U10718 (N_10718,N_10275,N_9067);
nor U10719 (N_10719,N_9049,N_9273);
xnor U10720 (N_10720,N_9570,N_9776);
nor U10721 (N_10721,N_9863,N_9258);
nand U10722 (N_10722,N_9079,N_9697);
and U10723 (N_10723,N_9317,N_9606);
or U10724 (N_10724,N_9160,N_9381);
nand U10725 (N_10725,N_9482,N_9146);
and U10726 (N_10726,N_9487,N_9132);
and U10727 (N_10727,N_9518,N_9824);
or U10728 (N_10728,N_9981,N_10284);
nand U10729 (N_10729,N_10125,N_9782);
and U10730 (N_10730,N_10160,N_10272);
and U10731 (N_10731,N_9881,N_9549);
and U10732 (N_10732,N_10231,N_9263);
xnor U10733 (N_10733,N_9808,N_9196);
nand U10734 (N_10734,N_9753,N_9723);
xor U10735 (N_10735,N_9489,N_9546);
nand U10736 (N_10736,N_9221,N_10200);
and U10737 (N_10737,N_9603,N_9172);
and U10738 (N_10738,N_9557,N_10086);
nand U10739 (N_10739,N_10260,N_9829);
nand U10740 (N_10740,N_10318,N_9170);
and U10741 (N_10741,N_10299,N_9385);
nand U10742 (N_10742,N_9501,N_9396);
and U10743 (N_10743,N_9926,N_9055);
and U10744 (N_10744,N_10236,N_9527);
nor U10745 (N_10745,N_9463,N_9704);
nand U10746 (N_10746,N_9491,N_9875);
nor U10747 (N_10747,N_9552,N_9400);
nor U10748 (N_10748,N_9740,N_9640);
and U10749 (N_10749,N_10258,N_10022);
and U10750 (N_10750,N_10040,N_9924);
and U10751 (N_10751,N_9878,N_10465);
nor U10752 (N_10752,N_9135,N_9094);
or U10753 (N_10753,N_9712,N_9588);
or U10754 (N_10754,N_9144,N_9907);
nor U10755 (N_10755,N_9932,N_9187);
or U10756 (N_10756,N_9614,N_10392);
xnor U10757 (N_10757,N_9714,N_10213);
nand U10758 (N_10758,N_9699,N_10328);
nand U10759 (N_10759,N_9111,N_9625);
or U10760 (N_10760,N_10184,N_9410);
or U10761 (N_10761,N_9455,N_9871);
or U10762 (N_10762,N_9976,N_9407);
nand U10763 (N_10763,N_9014,N_10238);
or U10764 (N_10764,N_9253,N_10131);
xor U10765 (N_10765,N_10375,N_9080);
xnor U10766 (N_10766,N_10407,N_10082);
nor U10767 (N_10767,N_9286,N_9082);
nor U10768 (N_10768,N_9792,N_9531);
or U10769 (N_10769,N_10496,N_10257);
nand U10770 (N_10770,N_9948,N_9277);
or U10771 (N_10771,N_9437,N_10411);
nand U10772 (N_10772,N_9522,N_9503);
xor U10773 (N_10773,N_9449,N_10304);
and U10774 (N_10774,N_9292,N_9683);
nand U10775 (N_10775,N_9086,N_9219);
nand U10776 (N_10776,N_9456,N_10391);
and U10777 (N_10777,N_9530,N_10425);
nor U10778 (N_10778,N_9065,N_10321);
and U10779 (N_10779,N_10240,N_9293);
and U10780 (N_10780,N_10206,N_9168);
nand U10781 (N_10781,N_9411,N_9921);
nand U10782 (N_10782,N_9666,N_9586);
and U10783 (N_10783,N_10003,N_10312);
and U10784 (N_10784,N_9852,N_10332);
nand U10785 (N_10785,N_10209,N_10363);
or U10786 (N_10786,N_9443,N_9481);
nand U10787 (N_10787,N_9423,N_10409);
nand U10788 (N_10788,N_9290,N_10002);
or U10789 (N_10789,N_9232,N_10067);
or U10790 (N_10790,N_10271,N_9755);
or U10791 (N_10791,N_9823,N_9599);
and U10792 (N_10792,N_10149,N_10358);
and U10793 (N_10793,N_9638,N_10108);
or U10794 (N_10794,N_9418,N_9982);
nand U10795 (N_10795,N_9913,N_9922);
and U10796 (N_10796,N_9369,N_9927);
nand U10797 (N_10797,N_9978,N_9595);
and U10798 (N_10798,N_9056,N_9690);
and U10799 (N_10799,N_9735,N_9685);
nor U10800 (N_10800,N_10220,N_10083);
nor U10801 (N_10801,N_10298,N_9536);
and U10802 (N_10802,N_10181,N_9584);
and U10803 (N_10803,N_9309,N_9175);
or U10804 (N_10804,N_9677,N_9585);
nand U10805 (N_10805,N_9793,N_9873);
xnor U10806 (N_10806,N_9280,N_9041);
and U10807 (N_10807,N_9653,N_10381);
or U10808 (N_10808,N_10457,N_10032);
nand U10809 (N_10809,N_9190,N_9085);
nand U10810 (N_10810,N_9862,N_10227);
nand U10811 (N_10811,N_9767,N_9667);
nand U10812 (N_10812,N_9313,N_9733);
and U10813 (N_10813,N_9153,N_9361);
nor U10814 (N_10814,N_9207,N_10119);
xor U10815 (N_10815,N_10323,N_9444);
or U10816 (N_10816,N_10097,N_9300);
and U10817 (N_10817,N_9248,N_10092);
and U10818 (N_10818,N_9433,N_9025);
nand U10819 (N_10819,N_9987,N_9562);
and U10820 (N_10820,N_9068,N_10342);
and U10821 (N_10821,N_9555,N_9892);
nor U10822 (N_10822,N_9213,N_9715);
nor U10823 (N_10823,N_9745,N_9870);
or U10824 (N_10824,N_9324,N_9591);
or U10825 (N_10825,N_9478,N_9684);
or U10826 (N_10826,N_9448,N_10474);
nor U10827 (N_10827,N_9741,N_9658);
or U10828 (N_10828,N_9006,N_9284);
nand U10829 (N_10829,N_9830,N_9943);
or U10830 (N_10830,N_9806,N_10210);
nor U10831 (N_10831,N_9209,N_9891);
and U10832 (N_10832,N_9030,N_10170);
and U10833 (N_10833,N_9543,N_9167);
and U10834 (N_10834,N_9601,N_10153);
nand U10835 (N_10835,N_9623,N_10124);
nand U10836 (N_10836,N_9093,N_9121);
nand U10837 (N_10837,N_9890,N_9626);
xor U10838 (N_10838,N_10398,N_9674);
nor U10839 (N_10839,N_9008,N_10448);
and U10840 (N_10840,N_9402,N_9222);
or U10841 (N_10841,N_9226,N_10144);
xnor U10842 (N_10842,N_9428,N_10094);
or U10843 (N_10843,N_9424,N_9724);
nor U10844 (N_10844,N_10397,N_9893);
or U10845 (N_10845,N_9972,N_9656);
nand U10846 (N_10846,N_9526,N_9617);
nand U10847 (N_10847,N_9059,N_9815);
or U10848 (N_10848,N_9088,N_9042);
or U10849 (N_10849,N_9188,N_10333);
nor U10850 (N_10850,N_9321,N_9427);
nand U10851 (N_10851,N_10478,N_9374);
and U10852 (N_10852,N_9298,N_9719);
nor U10853 (N_10853,N_9027,N_9636);
nor U10854 (N_10854,N_10463,N_9777);
nor U10855 (N_10855,N_9760,N_9053);
or U10856 (N_10856,N_9925,N_10313);
or U10857 (N_10857,N_10178,N_9787);
and U10858 (N_10858,N_9624,N_9050);
or U10859 (N_10859,N_9028,N_9021);
nor U10860 (N_10860,N_9498,N_9251);
xnor U10861 (N_10861,N_10286,N_10224);
and U10862 (N_10862,N_9602,N_10065);
or U10863 (N_10863,N_10268,N_9889);
or U10864 (N_10864,N_9752,N_9964);
or U10865 (N_10865,N_9814,N_9936);
or U10866 (N_10866,N_9593,N_10420);
and U10867 (N_10867,N_9988,N_9464);
nand U10868 (N_10868,N_10366,N_9840);
and U10869 (N_10869,N_9780,N_9375);
or U10870 (N_10870,N_10172,N_9537);
nor U10871 (N_10871,N_10027,N_10034);
nor U10872 (N_10872,N_9901,N_9012);
xor U10873 (N_10873,N_10221,N_9888);
and U10874 (N_10874,N_10175,N_10262);
and U10875 (N_10875,N_10091,N_9692);
nand U10876 (N_10876,N_9490,N_10476);
nor U10877 (N_10877,N_9853,N_9813);
or U10878 (N_10878,N_10090,N_9899);
and U10879 (N_10879,N_10338,N_10290);
nand U10880 (N_10880,N_9678,N_9472);
nand U10881 (N_10881,N_9876,N_9231);
or U10882 (N_10882,N_10044,N_9732);
nor U10883 (N_10883,N_9243,N_9470);
and U10884 (N_10884,N_10430,N_9176);
and U10885 (N_10885,N_9097,N_10031);
nor U10886 (N_10886,N_10089,N_9095);
nand U10887 (N_10887,N_9897,N_9159);
and U10888 (N_10888,N_10479,N_9534);
nand U10889 (N_10889,N_10339,N_10382);
or U10890 (N_10890,N_10467,N_10451);
nand U10891 (N_10891,N_9975,N_10431);
and U10892 (N_10892,N_9260,N_9070);
or U10893 (N_10893,N_9036,N_9763);
nand U10894 (N_10894,N_9074,N_9661);
or U10895 (N_10895,N_9296,N_9800);
or U10896 (N_10896,N_9130,N_9706);
xor U10897 (N_10897,N_10228,N_10029);
nor U10898 (N_10898,N_10461,N_10485);
and U10899 (N_10899,N_9492,N_10310);
nand U10900 (N_10900,N_10168,N_9308);
nand U10901 (N_10901,N_9194,N_9545);
nand U10902 (N_10902,N_10156,N_9687);
nor U10903 (N_10903,N_9211,N_9060);
and U10904 (N_10904,N_10245,N_9009);
or U10905 (N_10905,N_9299,N_9420);
and U10906 (N_10906,N_9331,N_9426);
or U10907 (N_10907,N_9802,N_9759);
and U10908 (N_10908,N_10100,N_9841);
nand U10909 (N_10909,N_9138,N_10203);
and U10910 (N_10910,N_9247,N_10437);
xnor U10911 (N_10911,N_10009,N_9504);
nand U10912 (N_10912,N_9991,N_9971);
and U10913 (N_10913,N_9903,N_10361);
nand U10914 (N_10914,N_9974,N_10080);
nor U10915 (N_10915,N_9650,N_10280);
nor U10916 (N_10916,N_9669,N_10189);
nor U10917 (N_10917,N_9276,N_10129);
or U10918 (N_10918,N_10302,N_10399);
nor U10919 (N_10919,N_10287,N_9191);
or U10920 (N_10920,N_9833,N_9347);
nand U10921 (N_10921,N_9880,N_10134);
xor U10922 (N_10922,N_9904,N_9281);
and U10923 (N_10923,N_9578,N_9744);
or U10924 (N_10924,N_10042,N_9147);
nor U10925 (N_10925,N_9198,N_9377);
and U10926 (N_10926,N_9957,N_9604);
and U10927 (N_10927,N_10166,N_9533);
nor U10928 (N_10928,N_9003,N_9596);
and U10929 (N_10929,N_10253,N_9528);
nand U10930 (N_10930,N_9000,N_10195);
or U10931 (N_10931,N_10374,N_9139);
and U10932 (N_10932,N_9370,N_9189);
and U10933 (N_10933,N_9200,N_9529);
xnor U10934 (N_10934,N_9432,N_10205);
nor U10935 (N_10935,N_9295,N_9613);
nor U10936 (N_10936,N_9412,N_9703);
xnor U10937 (N_10937,N_9785,N_9257);
or U10938 (N_10938,N_9769,N_10488);
nand U10939 (N_10939,N_10473,N_9458);
nor U10940 (N_10940,N_9124,N_9675);
and U10941 (N_10941,N_9707,N_9994);
xnor U10942 (N_10942,N_9990,N_9287);
nand U10943 (N_10943,N_10104,N_9746);
nor U10944 (N_10944,N_9212,N_9747);
and U10945 (N_10945,N_10225,N_9788);
nor U10946 (N_10946,N_9319,N_9886);
and U10947 (N_10947,N_10186,N_9195);
nor U10948 (N_10948,N_9197,N_10327);
or U10949 (N_10949,N_9949,N_9810);
or U10950 (N_10950,N_9325,N_9616);
nand U10951 (N_10951,N_10265,N_9169);
nor U10952 (N_10952,N_9181,N_9761);
or U10953 (N_10953,N_10201,N_9944);
and U10954 (N_10954,N_10491,N_9485);
or U10955 (N_10955,N_9016,N_10078);
nor U10956 (N_10956,N_9583,N_9966);
xnor U10957 (N_10957,N_9662,N_9770);
nor U10958 (N_10958,N_9457,N_9628);
and U10959 (N_10959,N_9043,N_10439);
nor U10960 (N_10960,N_9701,N_10426);
and U10961 (N_10961,N_9942,N_10400);
and U10962 (N_10962,N_9622,N_9327);
nand U10963 (N_10963,N_9516,N_10063);
nand U10964 (N_10964,N_9408,N_10133);
nor U10965 (N_10965,N_9726,N_9429);
or U10966 (N_10966,N_10076,N_10340);
and U10967 (N_10967,N_9883,N_10449);
nand U10968 (N_10968,N_10098,N_9154);
nor U10969 (N_10969,N_10115,N_10345);
nor U10970 (N_10970,N_9799,N_9587);
or U10971 (N_10971,N_10230,N_9230);
and U10972 (N_10972,N_9344,N_9345);
nand U10973 (N_10973,N_10126,N_9265);
nor U10974 (N_10974,N_9607,N_10281);
nand U10975 (N_10975,N_9334,N_10267);
and U10976 (N_10976,N_9571,N_10322);
nor U10977 (N_10977,N_9199,N_9217);
nor U10978 (N_10978,N_10365,N_9289);
nand U10979 (N_10979,N_10254,N_10147);
or U10980 (N_10980,N_9778,N_9355);
xnor U10981 (N_10981,N_10064,N_9502);
or U10982 (N_10982,N_10242,N_9267);
nor U10983 (N_10983,N_9520,N_9845);
nor U10984 (N_10984,N_9406,N_9173);
or U10985 (N_10985,N_9076,N_9148);
nand U10986 (N_10986,N_9998,N_9486);
and U10987 (N_10987,N_9203,N_9590);
nor U10988 (N_10988,N_9844,N_10259);
or U10989 (N_10989,N_10309,N_9118);
or U10990 (N_10990,N_9335,N_9655);
and U10991 (N_10991,N_9831,N_10099);
and U10992 (N_10992,N_9328,N_9326);
nor U10993 (N_10993,N_9695,N_9515);
and U10994 (N_10994,N_9820,N_9568);
and U10995 (N_10995,N_9161,N_10191);
and U10996 (N_10996,N_10456,N_10418);
or U10997 (N_10997,N_9496,N_9351);
nor U10998 (N_10998,N_9722,N_10025);
and U10999 (N_10999,N_10121,N_9615);
nand U11000 (N_11000,N_9024,N_9162);
and U11001 (N_11001,N_9506,N_9469);
nor U11002 (N_11002,N_9291,N_9380);
nand U11003 (N_11003,N_9956,N_9206);
xor U11004 (N_11004,N_9371,N_10188);
and U11005 (N_11005,N_9884,N_9311);
nor U11006 (N_11006,N_9635,N_10335);
and U11007 (N_11007,N_9315,N_10084);
xnor U11008 (N_11008,N_10110,N_10390);
or U11009 (N_11009,N_9032,N_9431);
xor U11010 (N_11010,N_9953,N_9680);
or U11011 (N_11011,N_10194,N_10232);
or U11012 (N_11012,N_9483,N_9133);
nand U11013 (N_11013,N_9384,N_9034);
xor U11014 (N_11014,N_10146,N_9102);
or U11015 (N_11015,N_10264,N_10037);
and U11016 (N_11016,N_10497,N_10079);
or U11017 (N_11017,N_9736,N_10249);
or U11018 (N_11018,N_9397,N_10483);
nand U11019 (N_11019,N_9730,N_9918);
nand U11020 (N_11020,N_10071,N_9855);
and U11021 (N_11021,N_9269,N_9882);
nand U11022 (N_11022,N_9275,N_10173);
or U11023 (N_11023,N_10329,N_9158);
or U11024 (N_11024,N_9645,N_10350);
nor U11025 (N_11025,N_9749,N_9762);
and U11026 (N_11026,N_10250,N_9182);
nor U11027 (N_11027,N_10419,N_10436);
and U11028 (N_11028,N_9013,N_9304);
xor U11029 (N_11029,N_10006,N_10096);
nor U11030 (N_11030,N_9672,N_9514);
and U11031 (N_11031,N_9224,N_10165);
and U11032 (N_11032,N_9007,N_9435);
and U11033 (N_11033,N_9100,N_9150);
and U11034 (N_11034,N_9698,N_9693);
nor U11035 (N_11035,N_9261,N_10159);
xnor U11036 (N_11036,N_9134,N_9945);
nor U11037 (N_11037,N_10247,N_9264);
or U11038 (N_11038,N_9054,N_10294);
nor U11039 (N_11039,N_9342,N_10442);
and U11040 (N_11040,N_9151,N_9500);
or U11041 (N_11041,N_9237,N_9818);
xor U11042 (N_11042,N_10285,N_9268);
and U11043 (N_11043,N_10023,N_10487);
xor U11044 (N_11044,N_9096,N_9419);
or U11045 (N_11045,N_10344,N_10388);
and U11046 (N_11046,N_10278,N_10434);
nand U11047 (N_11047,N_9434,N_9940);
xor U11048 (N_11048,N_9278,N_9497);
nor U11049 (N_11049,N_9748,N_9931);
or U11050 (N_11050,N_9960,N_9689);
xor U11051 (N_11051,N_10446,N_9033);
and U11052 (N_11052,N_9262,N_9288);
or U11053 (N_11053,N_9178,N_10348);
or U11054 (N_11054,N_9659,N_9524);
nor U11055 (N_11055,N_9346,N_9914);
nor U11056 (N_11056,N_10308,N_10288);
and U11057 (N_11057,N_9849,N_10140);
nor U11058 (N_11058,N_9312,N_10024);
xnor U11059 (N_11059,N_9861,N_10041);
and U11060 (N_11060,N_9241,N_9090);
xnor U11061 (N_11061,N_9670,N_9087);
nand U11062 (N_11062,N_9910,N_9123);
xnor U11063 (N_11063,N_10113,N_9022);
nand U11064 (N_11064,N_9580,N_10433);
or U11065 (N_11065,N_9558,N_10376);
nand U11066 (N_11066,N_9294,N_10018);
nor U11067 (N_11067,N_9803,N_9020);
and U11068 (N_11068,N_9547,N_10052);
xnor U11069 (N_11069,N_10215,N_10167);
or U11070 (N_11070,N_10111,N_10154);
xor U11071 (N_11071,N_10123,N_10152);
or U11072 (N_11072,N_9227,N_9163);
or U11073 (N_11073,N_10014,N_9937);
xnor U11074 (N_11074,N_10028,N_9417);
or U11075 (N_11075,N_10373,N_9999);
nand U11076 (N_11076,N_10177,N_9316);
nor U11077 (N_11077,N_9539,N_10480);
or U11078 (N_11078,N_9393,N_9376);
xor U11079 (N_11079,N_9646,N_10139);
and U11080 (N_11080,N_10062,N_9468);
xnor U11081 (N_11081,N_9152,N_9091);
nand U11082 (N_11082,N_9908,N_9573);
or U11083 (N_11083,N_9214,N_10432);
or U11084 (N_11084,N_10046,N_9239);
or U11085 (N_11085,N_9057,N_10073);
or U11086 (N_11086,N_10212,N_9836);
xnor U11087 (N_11087,N_9969,N_9950);
nor U11088 (N_11088,N_10011,N_9843);
or U11089 (N_11089,N_10492,N_9285);
or U11090 (N_11090,N_9002,N_10261);
nor U11091 (N_11091,N_10183,N_10049);
and U11092 (N_11092,N_9454,N_10246);
and U11093 (N_11093,N_9544,N_9349);
nor U11094 (N_11094,N_10057,N_10360);
nor U11095 (N_11095,N_9727,N_10199);
nand U11096 (N_11096,N_9729,N_9915);
nand U11097 (N_11097,N_10414,N_9409);
nand U11098 (N_11098,N_9851,N_9283);
xnor U11099 (N_11099,N_9967,N_9051);
xor U11100 (N_11100,N_9353,N_9679);
nand U11101 (N_11101,N_10386,N_10450);
and U11102 (N_11102,N_9446,N_9916);
nand U11103 (N_11103,N_9201,N_10198);
nand U11104 (N_11104,N_9453,N_9113);
and U11105 (N_11105,N_9917,N_9110);
or U11106 (N_11106,N_9477,N_9064);
nand U11107 (N_11107,N_9828,N_9781);
or U11108 (N_11108,N_10410,N_9572);
xor U11109 (N_11109,N_9018,N_9648);
or U11110 (N_11110,N_9244,N_9279);
and U11111 (N_11111,N_9634,N_9877);
xor U11112 (N_11112,N_10174,N_9935);
and U11113 (N_11113,N_10043,N_10102);
nor U11114 (N_11114,N_10007,N_10143);
nand U11115 (N_11115,N_10315,N_9023);
nor U11116 (N_11116,N_10336,N_9565);
or U11117 (N_11117,N_10088,N_10484);
nor U11118 (N_11118,N_10460,N_9598);
nand U11119 (N_11119,N_10164,N_10093);
or U11120 (N_11120,N_9495,N_10008);
nand U11121 (N_11121,N_9084,N_10402);
nand U11122 (N_11122,N_9218,N_9754);
or U11123 (N_11123,N_9307,N_10359);
and U11124 (N_11124,N_9493,N_10218);
nor U11125 (N_11125,N_10494,N_9794);
xor U11126 (N_11126,N_10486,N_9266);
and U11127 (N_11127,N_10444,N_9789);
nand U11128 (N_11128,N_9314,N_10369);
nor U11129 (N_11129,N_10326,N_10316);
and U11130 (N_11130,N_9322,N_9297);
or U11131 (N_11131,N_9461,N_9447);
nand U11132 (N_11132,N_9101,N_9594);
nand U11133 (N_11133,N_9005,N_9252);
and U11134 (N_11134,N_10109,N_10127);
and U11135 (N_11135,N_9436,N_10263);
nor U11136 (N_11136,N_9811,N_9996);
or U11137 (N_11137,N_9986,N_9846);
nand U11138 (N_11138,N_9928,N_9137);
and U11139 (N_11139,N_9554,N_10447);
and U11140 (N_11140,N_10269,N_9205);
and U11141 (N_11141,N_9479,N_9973);
nand U11142 (N_11142,N_10229,N_10122);
or U11143 (N_11143,N_9577,N_9644);
or U11144 (N_11144,N_9951,N_10406);
or U11145 (N_11145,N_10403,N_10196);
nor U11146 (N_11146,N_10116,N_9790);
nand U11147 (N_11147,N_10305,N_9037);
nand U11148 (N_11148,N_10142,N_10443);
nand U11149 (N_11149,N_9775,N_10475);
and U11150 (N_11150,N_9145,N_9125);
and U11151 (N_11151,N_9825,N_9460);
or U11152 (N_11152,N_9663,N_10466);
nand U11153 (N_11153,N_9965,N_10499);
or U11154 (N_11154,N_9271,N_9854);
and U11155 (N_11155,N_9306,N_9184);
or U11156 (N_11156,N_9850,N_9711);
nand U11157 (N_11157,N_10060,N_10204);
and U11158 (N_11158,N_9488,N_10050);
nor U11159 (N_11159,N_9983,N_9270);
and U11160 (N_11160,N_9499,N_9107);
nor U11161 (N_11161,N_10279,N_9415);
or U11162 (N_11162,N_10498,N_9869);
xnor U11163 (N_11163,N_9582,N_9993);
nand U11164 (N_11164,N_10158,N_9691);
or U11165 (N_11165,N_10197,N_9835);
and U11166 (N_11166,N_10070,N_9216);
or U11167 (N_11167,N_9360,N_9610);
nand U11168 (N_11168,N_9812,N_9235);
and U11169 (N_11169,N_9894,N_10056);
nand U11170 (N_11170,N_10005,N_10128);
nor U11171 (N_11171,N_9561,N_10319);
and U11172 (N_11172,N_9688,N_9395);
xor U11173 (N_11173,N_10393,N_9450);
and U11174 (N_11174,N_9164,N_9359);
xnor U11175 (N_11175,N_9401,N_9947);
and U11176 (N_11176,N_10004,N_10035);
and U11177 (N_11177,N_9112,N_10053);
and U11178 (N_11178,N_10138,N_9272);
and U11179 (N_11179,N_10012,N_9809);
nor U11180 (N_11180,N_9887,N_10239);
or U11181 (N_11181,N_9438,N_9738);
nor U11182 (N_11182,N_9480,N_9078);
and U11183 (N_11183,N_9508,N_10077);
nand U11184 (N_11184,N_9671,N_9035);
or U11185 (N_11185,N_9909,N_9540);
nor U11186 (N_11186,N_10297,N_10493);
nand U11187 (N_11187,N_9155,N_10001);
or U11188 (N_11188,N_10095,N_9389);
nor U11189 (N_11189,N_9856,N_9783);
or U11190 (N_11190,N_9451,N_9352);
nor U11191 (N_11191,N_9305,N_9192);
nor U11192 (N_11192,N_9958,N_9805);
nor U11193 (N_11193,N_10248,N_9795);
or U11194 (N_11194,N_10380,N_9301);
nor U11195 (N_11195,N_10489,N_9523);
nor U11196 (N_11196,N_9702,N_9934);
xor U11197 (N_11197,N_10117,N_9816);
nor U11198 (N_11198,N_9709,N_9249);
nor U11199 (N_11199,N_9553,N_9867);
nand U11200 (N_11200,N_10469,N_9077);
or U11201 (N_11201,N_9859,N_10157);
nor U11202 (N_11202,N_9885,N_9589);
nand U11203 (N_11203,N_9657,N_9128);
xor U11204 (N_11204,N_9099,N_10030);
and U11205 (N_11205,N_10182,N_9912);
xnor U11206 (N_11206,N_9282,N_10320);
xor U11207 (N_11207,N_10354,N_9742);
and U11208 (N_11208,N_10357,N_9183);
nor U11209 (N_11209,N_10352,N_10074);
nor U11210 (N_11210,N_10372,N_9075);
nand U11211 (N_11211,N_9929,N_9066);
or U11212 (N_11212,N_9992,N_9367);
nor U11213 (N_11213,N_10415,N_10470);
and U11214 (N_11214,N_9177,N_10148);
and U11215 (N_11215,N_10346,N_9548);
nand U11216 (N_11216,N_9141,N_9560);
nor U11217 (N_11217,N_9394,N_10378);
nor U11218 (N_11218,N_9651,N_9756);
nor U11219 (N_11219,N_10421,N_9302);
xor U11220 (N_11220,N_10395,N_10270);
xnor U11221 (N_11221,N_9339,N_9157);
or U11222 (N_11222,N_10190,N_9108);
nor U11223 (N_11223,N_10075,N_10453);
xnor U11224 (N_11224,N_10051,N_9513);
nor U11225 (N_11225,N_10151,N_9694);
xnor U11226 (N_11226,N_10293,N_9089);
nand U11227 (N_11227,N_9564,N_9728);
or U11228 (N_11228,N_9933,N_10404);
nor U11229 (N_11229,N_10058,N_9860);
nand U11230 (N_11230,N_10019,N_10235);
nand U11231 (N_11231,N_9413,N_10273);
nor U11232 (N_11232,N_9234,N_10408);
or U11233 (N_11233,N_9103,N_10039);
or U11234 (N_11234,N_10069,N_9143);
nor U11235 (N_11235,N_9700,N_10087);
nor U11236 (N_11236,N_10179,N_9372);
or U11237 (N_11237,N_10440,N_9062);
nand U11238 (N_11238,N_10072,N_10107);
and U11239 (N_11239,N_9015,N_10423);
and U11240 (N_11240,N_10112,N_9979);
nor U11241 (N_11241,N_10237,N_9462);
or U11242 (N_11242,N_9676,N_9627);
nor U11243 (N_11243,N_9039,N_9542);
and U11244 (N_11244,N_10396,N_10216);
nand U11245 (N_11245,N_9826,N_9404);
or U11246 (N_11246,N_10033,N_9398);
nor U11247 (N_11247,N_9047,N_10054);
and U11248 (N_11248,N_9797,N_9512);
nand U11249 (N_11249,N_9696,N_10481);
and U11250 (N_11250,N_10125,N_9462);
nand U11251 (N_11251,N_9168,N_9073);
or U11252 (N_11252,N_9717,N_9817);
or U11253 (N_11253,N_9408,N_10418);
or U11254 (N_11254,N_9390,N_10214);
nor U11255 (N_11255,N_9557,N_10033);
nor U11256 (N_11256,N_9068,N_9673);
nor U11257 (N_11257,N_10278,N_9351);
nor U11258 (N_11258,N_9380,N_9458);
nand U11259 (N_11259,N_10003,N_10110);
nor U11260 (N_11260,N_9876,N_10270);
or U11261 (N_11261,N_10044,N_9050);
or U11262 (N_11262,N_10069,N_10256);
or U11263 (N_11263,N_9335,N_9074);
or U11264 (N_11264,N_9953,N_9908);
nand U11265 (N_11265,N_9742,N_9967);
nor U11266 (N_11266,N_10496,N_9069);
or U11267 (N_11267,N_9663,N_10484);
and U11268 (N_11268,N_9583,N_9925);
or U11269 (N_11269,N_9854,N_9694);
xor U11270 (N_11270,N_10081,N_9966);
nor U11271 (N_11271,N_9907,N_9451);
nor U11272 (N_11272,N_9244,N_9007);
xnor U11273 (N_11273,N_9984,N_9757);
nor U11274 (N_11274,N_10482,N_10123);
nand U11275 (N_11275,N_10334,N_9397);
and U11276 (N_11276,N_9558,N_10481);
nor U11277 (N_11277,N_9015,N_9685);
nor U11278 (N_11278,N_9994,N_9810);
nor U11279 (N_11279,N_9564,N_10303);
nor U11280 (N_11280,N_10270,N_10190);
or U11281 (N_11281,N_10340,N_9154);
nand U11282 (N_11282,N_9230,N_9063);
or U11283 (N_11283,N_9310,N_9849);
xnor U11284 (N_11284,N_9278,N_9020);
and U11285 (N_11285,N_9591,N_9492);
nor U11286 (N_11286,N_9127,N_9383);
nor U11287 (N_11287,N_9722,N_9822);
nand U11288 (N_11288,N_9660,N_9183);
nor U11289 (N_11289,N_10007,N_10484);
or U11290 (N_11290,N_10470,N_9496);
nand U11291 (N_11291,N_9949,N_10397);
nor U11292 (N_11292,N_9329,N_10452);
nand U11293 (N_11293,N_9656,N_9819);
or U11294 (N_11294,N_9322,N_9354);
nor U11295 (N_11295,N_9754,N_10469);
nand U11296 (N_11296,N_10281,N_9227);
nand U11297 (N_11297,N_10458,N_9293);
xor U11298 (N_11298,N_9104,N_9019);
nand U11299 (N_11299,N_10005,N_10415);
and U11300 (N_11300,N_9600,N_10490);
nor U11301 (N_11301,N_10389,N_10076);
nand U11302 (N_11302,N_9822,N_9385);
nor U11303 (N_11303,N_9192,N_10321);
and U11304 (N_11304,N_9352,N_9474);
and U11305 (N_11305,N_9028,N_9869);
nand U11306 (N_11306,N_10195,N_10410);
and U11307 (N_11307,N_10471,N_10257);
nor U11308 (N_11308,N_10245,N_9318);
nor U11309 (N_11309,N_10056,N_9496);
or U11310 (N_11310,N_9494,N_9839);
and U11311 (N_11311,N_10101,N_10042);
nand U11312 (N_11312,N_10085,N_9134);
or U11313 (N_11313,N_9723,N_9708);
nor U11314 (N_11314,N_9501,N_9573);
nand U11315 (N_11315,N_9467,N_9022);
nand U11316 (N_11316,N_9143,N_9707);
nand U11317 (N_11317,N_9441,N_10434);
nor U11318 (N_11318,N_10145,N_9308);
or U11319 (N_11319,N_10086,N_9771);
and U11320 (N_11320,N_9726,N_9349);
nand U11321 (N_11321,N_9400,N_9723);
nor U11322 (N_11322,N_9831,N_9696);
nand U11323 (N_11323,N_10332,N_9414);
xnor U11324 (N_11324,N_9703,N_9928);
nand U11325 (N_11325,N_10117,N_10014);
and U11326 (N_11326,N_10259,N_10187);
xor U11327 (N_11327,N_9338,N_9516);
nor U11328 (N_11328,N_9274,N_9047);
xnor U11329 (N_11329,N_9313,N_9146);
nor U11330 (N_11330,N_10256,N_9061);
or U11331 (N_11331,N_9971,N_9810);
or U11332 (N_11332,N_10248,N_9312);
and U11333 (N_11333,N_10379,N_9860);
nand U11334 (N_11334,N_9594,N_10233);
nor U11335 (N_11335,N_9836,N_9622);
nand U11336 (N_11336,N_9148,N_9020);
and U11337 (N_11337,N_9537,N_9885);
nand U11338 (N_11338,N_10077,N_9910);
nor U11339 (N_11339,N_9241,N_10106);
nand U11340 (N_11340,N_9267,N_10446);
and U11341 (N_11341,N_10067,N_9546);
nand U11342 (N_11342,N_9257,N_9887);
nand U11343 (N_11343,N_10405,N_9555);
nand U11344 (N_11344,N_10370,N_10322);
or U11345 (N_11345,N_9647,N_9174);
nor U11346 (N_11346,N_10332,N_9174);
nor U11347 (N_11347,N_9543,N_10281);
and U11348 (N_11348,N_9076,N_9995);
nor U11349 (N_11349,N_10421,N_9461);
and U11350 (N_11350,N_10453,N_9748);
xnor U11351 (N_11351,N_9199,N_9680);
xor U11352 (N_11352,N_9812,N_10221);
nand U11353 (N_11353,N_10157,N_10096);
nand U11354 (N_11354,N_9086,N_10305);
and U11355 (N_11355,N_9143,N_10368);
xor U11356 (N_11356,N_9717,N_9362);
or U11357 (N_11357,N_10344,N_9185);
or U11358 (N_11358,N_9601,N_9639);
nand U11359 (N_11359,N_9822,N_9017);
or U11360 (N_11360,N_9114,N_10135);
and U11361 (N_11361,N_9280,N_10087);
nand U11362 (N_11362,N_9319,N_9604);
nand U11363 (N_11363,N_10261,N_9122);
and U11364 (N_11364,N_9272,N_9138);
nor U11365 (N_11365,N_9532,N_10332);
or U11366 (N_11366,N_10129,N_9716);
nor U11367 (N_11367,N_9595,N_9693);
or U11368 (N_11368,N_9359,N_10485);
nand U11369 (N_11369,N_9092,N_10183);
and U11370 (N_11370,N_9317,N_9415);
and U11371 (N_11371,N_9407,N_10466);
xor U11372 (N_11372,N_10048,N_9461);
nor U11373 (N_11373,N_9050,N_9977);
nor U11374 (N_11374,N_10059,N_9948);
nor U11375 (N_11375,N_9322,N_10027);
and U11376 (N_11376,N_9804,N_9227);
or U11377 (N_11377,N_9041,N_10402);
and U11378 (N_11378,N_9952,N_10269);
and U11379 (N_11379,N_9388,N_10422);
or U11380 (N_11380,N_9960,N_10096);
nand U11381 (N_11381,N_9018,N_10246);
xor U11382 (N_11382,N_9945,N_10445);
xnor U11383 (N_11383,N_10311,N_9199);
nor U11384 (N_11384,N_9319,N_9746);
or U11385 (N_11385,N_9342,N_10102);
and U11386 (N_11386,N_9288,N_10121);
or U11387 (N_11387,N_10485,N_9660);
or U11388 (N_11388,N_10407,N_10461);
and U11389 (N_11389,N_9188,N_9988);
or U11390 (N_11390,N_9351,N_10044);
or U11391 (N_11391,N_9272,N_9453);
nand U11392 (N_11392,N_10008,N_9343);
or U11393 (N_11393,N_9270,N_9718);
nor U11394 (N_11394,N_9268,N_9563);
nor U11395 (N_11395,N_9604,N_9306);
and U11396 (N_11396,N_10326,N_10012);
nand U11397 (N_11397,N_9657,N_10353);
and U11398 (N_11398,N_9017,N_9067);
nand U11399 (N_11399,N_9883,N_10206);
nor U11400 (N_11400,N_10484,N_10218);
nor U11401 (N_11401,N_9702,N_10281);
or U11402 (N_11402,N_10065,N_10034);
or U11403 (N_11403,N_9537,N_9848);
and U11404 (N_11404,N_10103,N_9452);
nor U11405 (N_11405,N_9424,N_9879);
nand U11406 (N_11406,N_9050,N_10455);
nor U11407 (N_11407,N_9126,N_9130);
nand U11408 (N_11408,N_9159,N_10384);
or U11409 (N_11409,N_10273,N_9390);
nand U11410 (N_11410,N_10323,N_9277);
and U11411 (N_11411,N_10480,N_9637);
nand U11412 (N_11412,N_9799,N_10328);
or U11413 (N_11413,N_9178,N_9878);
nand U11414 (N_11414,N_10075,N_9015);
xnor U11415 (N_11415,N_9923,N_9962);
nor U11416 (N_11416,N_9476,N_10377);
and U11417 (N_11417,N_10279,N_10444);
and U11418 (N_11418,N_10494,N_9342);
or U11419 (N_11419,N_9445,N_9457);
nor U11420 (N_11420,N_9927,N_9994);
or U11421 (N_11421,N_9815,N_9697);
nand U11422 (N_11422,N_9040,N_9279);
or U11423 (N_11423,N_9342,N_9696);
xnor U11424 (N_11424,N_9910,N_10066);
nand U11425 (N_11425,N_9848,N_10128);
nor U11426 (N_11426,N_9976,N_10006);
and U11427 (N_11427,N_9778,N_9133);
or U11428 (N_11428,N_10295,N_9899);
nand U11429 (N_11429,N_9574,N_10292);
or U11430 (N_11430,N_10213,N_9782);
and U11431 (N_11431,N_10122,N_9000);
xor U11432 (N_11432,N_9875,N_9975);
nor U11433 (N_11433,N_9752,N_10038);
or U11434 (N_11434,N_9524,N_9676);
nor U11435 (N_11435,N_9820,N_9458);
or U11436 (N_11436,N_10228,N_10105);
nor U11437 (N_11437,N_9880,N_9988);
and U11438 (N_11438,N_9397,N_9041);
and U11439 (N_11439,N_10178,N_10048);
or U11440 (N_11440,N_9527,N_9749);
nor U11441 (N_11441,N_9154,N_9621);
and U11442 (N_11442,N_9232,N_9599);
nand U11443 (N_11443,N_10306,N_9846);
or U11444 (N_11444,N_10436,N_9357);
or U11445 (N_11445,N_9814,N_9884);
nor U11446 (N_11446,N_9858,N_9946);
nand U11447 (N_11447,N_9016,N_10136);
nor U11448 (N_11448,N_10040,N_9368);
and U11449 (N_11449,N_10320,N_9235);
nand U11450 (N_11450,N_10084,N_9774);
nor U11451 (N_11451,N_9977,N_9613);
and U11452 (N_11452,N_9462,N_10491);
nand U11453 (N_11453,N_9188,N_9069);
nand U11454 (N_11454,N_10193,N_9868);
or U11455 (N_11455,N_10034,N_10476);
or U11456 (N_11456,N_9430,N_9864);
nor U11457 (N_11457,N_9571,N_9166);
nand U11458 (N_11458,N_9093,N_9593);
and U11459 (N_11459,N_10133,N_9498);
nor U11460 (N_11460,N_9108,N_9593);
or U11461 (N_11461,N_9080,N_9505);
nor U11462 (N_11462,N_10292,N_10408);
or U11463 (N_11463,N_9541,N_9074);
nor U11464 (N_11464,N_9474,N_9107);
nand U11465 (N_11465,N_10134,N_9718);
xor U11466 (N_11466,N_9772,N_10430);
and U11467 (N_11467,N_9863,N_9023);
or U11468 (N_11468,N_9483,N_10389);
and U11469 (N_11469,N_9541,N_9166);
or U11470 (N_11470,N_9578,N_10496);
or U11471 (N_11471,N_9106,N_10100);
xnor U11472 (N_11472,N_9879,N_9324);
or U11473 (N_11473,N_9072,N_9625);
nand U11474 (N_11474,N_10120,N_9981);
or U11475 (N_11475,N_9369,N_10423);
nor U11476 (N_11476,N_9566,N_9156);
xor U11477 (N_11477,N_9641,N_9436);
or U11478 (N_11478,N_10479,N_10463);
or U11479 (N_11479,N_9642,N_10079);
or U11480 (N_11480,N_9370,N_9294);
nor U11481 (N_11481,N_10032,N_9529);
nand U11482 (N_11482,N_9858,N_10431);
and U11483 (N_11483,N_9169,N_9651);
and U11484 (N_11484,N_9393,N_10285);
xor U11485 (N_11485,N_9818,N_9527);
or U11486 (N_11486,N_9495,N_9274);
or U11487 (N_11487,N_9351,N_9168);
nor U11488 (N_11488,N_9521,N_10468);
or U11489 (N_11489,N_9499,N_9899);
nand U11490 (N_11490,N_9834,N_9723);
and U11491 (N_11491,N_10073,N_9126);
or U11492 (N_11492,N_10300,N_9858);
nand U11493 (N_11493,N_10192,N_10376);
or U11494 (N_11494,N_10334,N_9043);
or U11495 (N_11495,N_10465,N_9471);
or U11496 (N_11496,N_10462,N_10361);
and U11497 (N_11497,N_9997,N_10185);
xor U11498 (N_11498,N_10061,N_9698);
nand U11499 (N_11499,N_9158,N_9667);
nand U11500 (N_11500,N_10447,N_9795);
xor U11501 (N_11501,N_9910,N_9327);
or U11502 (N_11502,N_9507,N_10258);
nor U11503 (N_11503,N_10197,N_9540);
xnor U11504 (N_11504,N_10489,N_9079);
xnor U11505 (N_11505,N_10142,N_9295);
or U11506 (N_11506,N_9247,N_9853);
or U11507 (N_11507,N_10263,N_9229);
nor U11508 (N_11508,N_9926,N_10082);
and U11509 (N_11509,N_10478,N_9591);
and U11510 (N_11510,N_9497,N_9200);
and U11511 (N_11511,N_9386,N_9766);
nor U11512 (N_11512,N_9903,N_10138);
or U11513 (N_11513,N_9211,N_9978);
and U11514 (N_11514,N_10476,N_9409);
nand U11515 (N_11515,N_10445,N_10436);
and U11516 (N_11516,N_9743,N_9017);
nand U11517 (N_11517,N_9008,N_9525);
and U11518 (N_11518,N_9430,N_9725);
nor U11519 (N_11519,N_10348,N_9512);
xor U11520 (N_11520,N_9783,N_9640);
nor U11521 (N_11521,N_9517,N_9084);
nand U11522 (N_11522,N_10363,N_10094);
nand U11523 (N_11523,N_10139,N_9270);
nor U11524 (N_11524,N_9828,N_10215);
and U11525 (N_11525,N_10396,N_10199);
or U11526 (N_11526,N_10286,N_9926);
and U11527 (N_11527,N_10211,N_9562);
or U11528 (N_11528,N_10350,N_9943);
or U11529 (N_11529,N_9886,N_10064);
or U11530 (N_11530,N_9097,N_9066);
or U11531 (N_11531,N_10495,N_10111);
and U11532 (N_11532,N_9475,N_9182);
or U11533 (N_11533,N_9166,N_9122);
xnor U11534 (N_11534,N_9851,N_9651);
nor U11535 (N_11535,N_9720,N_9581);
nor U11536 (N_11536,N_9213,N_9013);
nand U11537 (N_11537,N_10019,N_10151);
and U11538 (N_11538,N_9090,N_9716);
xnor U11539 (N_11539,N_9737,N_9436);
xnor U11540 (N_11540,N_9818,N_9781);
nand U11541 (N_11541,N_9495,N_9246);
nand U11542 (N_11542,N_9991,N_9757);
nand U11543 (N_11543,N_9277,N_9413);
and U11544 (N_11544,N_10457,N_10404);
and U11545 (N_11545,N_9381,N_9806);
or U11546 (N_11546,N_9743,N_10111);
and U11547 (N_11547,N_9486,N_10325);
or U11548 (N_11548,N_10236,N_10135);
nand U11549 (N_11549,N_9646,N_10438);
nor U11550 (N_11550,N_9052,N_9927);
or U11551 (N_11551,N_9432,N_9493);
nor U11552 (N_11552,N_9068,N_9204);
or U11553 (N_11553,N_9232,N_9143);
or U11554 (N_11554,N_10191,N_9230);
nor U11555 (N_11555,N_10151,N_9576);
or U11556 (N_11556,N_9540,N_9823);
nand U11557 (N_11557,N_10215,N_9980);
and U11558 (N_11558,N_9406,N_9032);
nand U11559 (N_11559,N_9266,N_9250);
nor U11560 (N_11560,N_9064,N_10488);
nand U11561 (N_11561,N_9496,N_9246);
nand U11562 (N_11562,N_10277,N_9065);
nor U11563 (N_11563,N_10060,N_10129);
nor U11564 (N_11564,N_10343,N_9379);
xnor U11565 (N_11565,N_9528,N_9618);
nor U11566 (N_11566,N_10271,N_10484);
nor U11567 (N_11567,N_10336,N_9319);
nor U11568 (N_11568,N_9496,N_9613);
nand U11569 (N_11569,N_10187,N_10319);
and U11570 (N_11570,N_9041,N_9504);
xor U11571 (N_11571,N_9420,N_10169);
or U11572 (N_11572,N_9774,N_9458);
xnor U11573 (N_11573,N_9182,N_10245);
nor U11574 (N_11574,N_9521,N_9898);
nor U11575 (N_11575,N_9023,N_9974);
xnor U11576 (N_11576,N_9870,N_9731);
xor U11577 (N_11577,N_9717,N_9350);
and U11578 (N_11578,N_10222,N_9556);
or U11579 (N_11579,N_10456,N_9675);
and U11580 (N_11580,N_9217,N_9444);
or U11581 (N_11581,N_9401,N_9413);
or U11582 (N_11582,N_9149,N_10121);
nand U11583 (N_11583,N_9856,N_9135);
and U11584 (N_11584,N_9411,N_9058);
nand U11585 (N_11585,N_9657,N_9308);
and U11586 (N_11586,N_10112,N_9946);
and U11587 (N_11587,N_9801,N_9123);
or U11588 (N_11588,N_10271,N_10396);
nand U11589 (N_11589,N_9270,N_10086);
or U11590 (N_11590,N_10236,N_9422);
and U11591 (N_11591,N_10332,N_9262);
and U11592 (N_11592,N_9865,N_10240);
or U11593 (N_11593,N_10253,N_10035);
and U11594 (N_11594,N_9020,N_10285);
nand U11595 (N_11595,N_10444,N_9649);
nor U11596 (N_11596,N_10413,N_9034);
xor U11597 (N_11597,N_9408,N_9516);
xor U11598 (N_11598,N_10487,N_9720);
nor U11599 (N_11599,N_9532,N_9983);
or U11600 (N_11600,N_9477,N_9555);
nand U11601 (N_11601,N_9635,N_9620);
nand U11602 (N_11602,N_9644,N_9929);
xnor U11603 (N_11603,N_9571,N_10098);
nand U11604 (N_11604,N_9915,N_10395);
or U11605 (N_11605,N_10129,N_9306);
and U11606 (N_11606,N_10431,N_9905);
and U11607 (N_11607,N_10424,N_9870);
and U11608 (N_11608,N_9803,N_10023);
or U11609 (N_11609,N_10308,N_9280);
and U11610 (N_11610,N_9300,N_9266);
nand U11611 (N_11611,N_10377,N_10306);
or U11612 (N_11612,N_9986,N_9027);
and U11613 (N_11613,N_9059,N_10173);
nand U11614 (N_11614,N_10488,N_9953);
nor U11615 (N_11615,N_9474,N_10210);
nand U11616 (N_11616,N_10326,N_9991);
or U11617 (N_11617,N_10444,N_9555);
or U11618 (N_11618,N_9868,N_9598);
or U11619 (N_11619,N_10435,N_10371);
or U11620 (N_11620,N_9474,N_9615);
and U11621 (N_11621,N_10355,N_9495);
nor U11622 (N_11622,N_10288,N_10227);
nor U11623 (N_11623,N_9846,N_9122);
nor U11624 (N_11624,N_10428,N_10426);
or U11625 (N_11625,N_9953,N_10429);
nor U11626 (N_11626,N_9135,N_9353);
xor U11627 (N_11627,N_9018,N_9853);
nand U11628 (N_11628,N_9877,N_9646);
xnor U11629 (N_11629,N_9052,N_10087);
or U11630 (N_11630,N_9765,N_9905);
nand U11631 (N_11631,N_9486,N_9352);
nand U11632 (N_11632,N_9715,N_10220);
nand U11633 (N_11633,N_9066,N_10017);
xnor U11634 (N_11634,N_9767,N_9648);
xor U11635 (N_11635,N_10278,N_9685);
and U11636 (N_11636,N_9214,N_9018);
and U11637 (N_11637,N_9912,N_10393);
and U11638 (N_11638,N_9254,N_9151);
xnor U11639 (N_11639,N_9389,N_9136);
or U11640 (N_11640,N_9303,N_9912);
nand U11641 (N_11641,N_10105,N_9550);
xor U11642 (N_11642,N_9585,N_9168);
xor U11643 (N_11643,N_9467,N_9217);
nor U11644 (N_11644,N_9505,N_9215);
nor U11645 (N_11645,N_9970,N_9118);
nor U11646 (N_11646,N_9191,N_10145);
and U11647 (N_11647,N_10138,N_10382);
nor U11648 (N_11648,N_9193,N_9753);
and U11649 (N_11649,N_10149,N_10421);
or U11650 (N_11650,N_9989,N_9411);
and U11651 (N_11651,N_9664,N_10045);
or U11652 (N_11652,N_10231,N_9607);
and U11653 (N_11653,N_9494,N_9727);
and U11654 (N_11654,N_10253,N_9538);
and U11655 (N_11655,N_10326,N_10207);
nand U11656 (N_11656,N_10291,N_9030);
nand U11657 (N_11657,N_9824,N_9696);
or U11658 (N_11658,N_9803,N_10263);
nand U11659 (N_11659,N_10191,N_10209);
and U11660 (N_11660,N_9694,N_9816);
nand U11661 (N_11661,N_10093,N_9461);
nand U11662 (N_11662,N_9503,N_9725);
and U11663 (N_11663,N_9238,N_9522);
nand U11664 (N_11664,N_9217,N_10095);
or U11665 (N_11665,N_10298,N_9847);
and U11666 (N_11666,N_10408,N_10446);
nor U11667 (N_11667,N_10435,N_9628);
nor U11668 (N_11668,N_9476,N_9928);
and U11669 (N_11669,N_9392,N_9525);
nor U11670 (N_11670,N_10413,N_10263);
and U11671 (N_11671,N_9397,N_9999);
nand U11672 (N_11672,N_9865,N_9612);
nor U11673 (N_11673,N_10232,N_9504);
xnor U11674 (N_11674,N_9981,N_10349);
or U11675 (N_11675,N_9096,N_10185);
or U11676 (N_11676,N_9318,N_9398);
nor U11677 (N_11677,N_10172,N_9689);
nor U11678 (N_11678,N_10146,N_10169);
nor U11679 (N_11679,N_9959,N_9673);
or U11680 (N_11680,N_9713,N_9013);
and U11681 (N_11681,N_10449,N_9186);
and U11682 (N_11682,N_10045,N_9707);
nor U11683 (N_11683,N_9046,N_9604);
and U11684 (N_11684,N_10396,N_9880);
xor U11685 (N_11685,N_9002,N_9290);
and U11686 (N_11686,N_9352,N_9555);
nand U11687 (N_11687,N_9343,N_9060);
xor U11688 (N_11688,N_10417,N_9245);
xnor U11689 (N_11689,N_10046,N_10325);
nand U11690 (N_11690,N_9500,N_9282);
nor U11691 (N_11691,N_9405,N_9908);
nor U11692 (N_11692,N_10178,N_9472);
and U11693 (N_11693,N_9331,N_9251);
or U11694 (N_11694,N_10199,N_9077);
and U11695 (N_11695,N_9167,N_9282);
and U11696 (N_11696,N_9364,N_10256);
and U11697 (N_11697,N_10120,N_10209);
xnor U11698 (N_11698,N_9458,N_10045);
and U11699 (N_11699,N_10210,N_9673);
xnor U11700 (N_11700,N_9346,N_9569);
and U11701 (N_11701,N_10118,N_9061);
nand U11702 (N_11702,N_9382,N_9156);
and U11703 (N_11703,N_10434,N_10446);
and U11704 (N_11704,N_9741,N_10372);
nor U11705 (N_11705,N_9724,N_9434);
nand U11706 (N_11706,N_9690,N_9072);
or U11707 (N_11707,N_9151,N_9489);
xor U11708 (N_11708,N_9400,N_9430);
xnor U11709 (N_11709,N_10172,N_9917);
nor U11710 (N_11710,N_9485,N_9000);
or U11711 (N_11711,N_9252,N_9869);
nor U11712 (N_11712,N_9559,N_9563);
and U11713 (N_11713,N_9135,N_10418);
nand U11714 (N_11714,N_9430,N_9682);
xnor U11715 (N_11715,N_10479,N_9813);
and U11716 (N_11716,N_9091,N_9325);
xor U11717 (N_11717,N_10075,N_9483);
nor U11718 (N_11718,N_9737,N_9318);
nand U11719 (N_11719,N_9821,N_9195);
nor U11720 (N_11720,N_9298,N_9123);
nand U11721 (N_11721,N_9961,N_10435);
and U11722 (N_11722,N_9866,N_9393);
or U11723 (N_11723,N_10279,N_9589);
or U11724 (N_11724,N_10015,N_10397);
or U11725 (N_11725,N_9591,N_9336);
and U11726 (N_11726,N_9391,N_10037);
and U11727 (N_11727,N_10089,N_9527);
nor U11728 (N_11728,N_9920,N_10075);
xor U11729 (N_11729,N_10282,N_10137);
nand U11730 (N_11730,N_9504,N_9982);
or U11731 (N_11731,N_10001,N_9788);
nand U11732 (N_11732,N_9851,N_9568);
nand U11733 (N_11733,N_9185,N_9402);
nor U11734 (N_11734,N_9811,N_9583);
nor U11735 (N_11735,N_9545,N_9872);
nor U11736 (N_11736,N_9925,N_9494);
nor U11737 (N_11737,N_9755,N_10233);
nor U11738 (N_11738,N_9985,N_9429);
or U11739 (N_11739,N_9258,N_9480);
and U11740 (N_11740,N_9726,N_9619);
or U11741 (N_11741,N_9810,N_9276);
or U11742 (N_11742,N_9884,N_10033);
nor U11743 (N_11743,N_9012,N_10209);
and U11744 (N_11744,N_9457,N_10128);
and U11745 (N_11745,N_9475,N_9548);
nor U11746 (N_11746,N_9429,N_9357);
xor U11747 (N_11747,N_9273,N_9203);
nor U11748 (N_11748,N_9771,N_9027);
or U11749 (N_11749,N_10390,N_10329);
and U11750 (N_11750,N_10383,N_9392);
nor U11751 (N_11751,N_9597,N_9850);
nand U11752 (N_11752,N_9363,N_10276);
xor U11753 (N_11753,N_9408,N_9207);
or U11754 (N_11754,N_9890,N_9747);
nand U11755 (N_11755,N_9916,N_10267);
nor U11756 (N_11756,N_9952,N_10162);
and U11757 (N_11757,N_9699,N_9740);
or U11758 (N_11758,N_9007,N_10175);
nor U11759 (N_11759,N_9225,N_9369);
nor U11760 (N_11760,N_9301,N_9038);
nor U11761 (N_11761,N_9376,N_9005);
nor U11762 (N_11762,N_9806,N_9784);
nand U11763 (N_11763,N_9610,N_10396);
xnor U11764 (N_11764,N_10229,N_10062);
xnor U11765 (N_11765,N_9621,N_9919);
or U11766 (N_11766,N_10438,N_9814);
nand U11767 (N_11767,N_9133,N_9148);
nor U11768 (N_11768,N_9721,N_9304);
or U11769 (N_11769,N_9359,N_10421);
or U11770 (N_11770,N_9460,N_10187);
nor U11771 (N_11771,N_10208,N_9503);
xnor U11772 (N_11772,N_9138,N_9685);
and U11773 (N_11773,N_9659,N_10406);
and U11774 (N_11774,N_9036,N_9290);
xor U11775 (N_11775,N_9490,N_10442);
nor U11776 (N_11776,N_10323,N_9058);
and U11777 (N_11777,N_9761,N_10182);
or U11778 (N_11778,N_9006,N_9272);
nor U11779 (N_11779,N_9219,N_9856);
nand U11780 (N_11780,N_9702,N_10285);
nor U11781 (N_11781,N_9347,N_9234);
nor U11782 (N_11782,N_9699,N_10014);
or U11783 (N_11783,N_9213,N_9906);
and U11784 (N_11784,N_10292,N_9228);
or U11785 (N_11785,N_9053,N_9701);
nand U11786 (N_11786,N_10186,N_9179);
nand U11787 (N_11787,N_9688,N_9712);
or U11788 (N_11788,N_9086,N_9760);
nor U11789 (N_11789,N_9016,N_9328);
nand U11790 (N_11790,N_9618,N_10028);
and U11791 (N_11791,N_9674,N_10362);
and U11792 (N_11792,N_9716,N_9341);
or U11793 (N_11793,N_10496,N_9932);
nor U11794 (N_11794,N_9092,N_9880);
nand U11795 (N_11795,N_9365,N_10007);
and U11796 (N_11796,N_10073,N_9208);
or U11797 (N_11797,N_10185,N_10330);
nor U11798 (N_11798,N_10138,N_9166);
nor U11799 (N_11799,N_10106,N_9217);
nand U11800 (N_11800,N_9142,N_9110);
and U11801 (N_11801,N_9416,N_9299);
or U11802 (N_11802,N_9181,N_9546);
nor U11803 (N_11803,N_9312,N_9558);
or U11804 (N_11804,N_9100,N_10357);
and U11805 (N_11805,N_9813,N_10294);
and U11806 (N_11806,N_9585,N_9719);
and U11807 (N_11807,N_9501,N_9451);
or U11808 (N_11808,N_9159,N_9351);
nor U11809 (N_11809,N_9795,N_10094);
and U11810 (N_11810,N_10316,N_10353);
nor U11811 (N_11811,N_9886,N_9671);
nand U11812 (N_11812,N_9892,N_9896);
nor U11813 (N_11813,N_10403,N_9551);
nand U11814 (N_11814,N_9387,N_10378);
and U11815 (N_11815,N_10108,N_10268);
nor U11816 (N_11816,N_9517,N_10194);
nor U11817 (N_11817,N_9116,N_10411);
xor U11818 (N_11818,N_10193,N_9665);
nand U11819 (N_11819,N_10317,N_9865);
nor U11820 (N_11820,N_9017,N_10333);
or U11821 (N_11821,N_9364,N_9922);
nand U11822 (N_11822,N_9058,N_9192);
nand U11823 (N_11823,N_10118,N_9744);
nor U11824 (N_11824,N_9278,N_9511);
or U11825 (N_11825,N_9853,N_10192);
nand U11826 (N_11826,N_10441,N_9075);
nor U11827 (N_11827,N_9562,N_9718);
nor U11828 (N_11828,N_9360,N_9769);
nor U11829 (N_11829,N_10301,N_9072);
nand U11830 (N_11830,N_9336,N_9933);
nand U11831 (N_11831,N_9321,N_10239);
nand U11832 (N_11832,N_10495,N_9402);
nand U11833 (N_11833,N_9639,N_10278);
or U11834 (N_11834,N_9079,N_9083);
nor U11835 (N_11835,N_9592,N_9276);
or U11836 (N_11836,N_9255,N_9998);
nand U11837 (N_11837,N_9669,N_9746);
xor U11838 (N_11838,N_9500,N_10329);
or U11839 (N_11839,N_9946,N_10298);
or U11840 (N_11840,N_10119,N_10105);
xor U11841 (N_11841,N_9387,N_9600);
or U11842 (N_11842,N_9021,N_9749);
and U11843 (N_11843,N_9011,N_10042);
or U11844 (N_11844,N_9801,N_9235);
nand U11845 (N_11845,N_10415,N_10338);
and U11846 (N_11846,N_9678,N_10212);
xnor U11847 (N_11847,N_10194,N_10381);
or U11848 (N_11848,N_10411,N_9884);
or U11849 (N_11849,N_9430,N_9300);
nand U11850 (N_11850,N_10049,N_9836);
nor U11851 (N_11851,N_10484,N_9938);
and U11852 (N_11852,N_9773,N_9734);
nand U11853 (N_11853,N_10424,N_10118);
or U11854 (N_11854,N_9659,N_9319);
nand U11855 (N_11855,N_9553,N_10344);
nor U11856 (N_11856,N_9847,N_9304);
and U11857 (N_11857,N_9159,N_9445);
xor U11858 (N_11858,N_9616,N_10129);
xnor U11859 (N_11859,N_10083,N_9598);
xor U11860 (N_11860,N_9135,N_9843);
or U11861 (N_11861,N_9990,N_9486);
nand U11862 (N_11862,N_9478,N_9422);
nand U11863 (N_11863,N_10398,N_9758);
nand U11864 (N_11864,N_9109,N_9346);
or U11865 (N_11865,N_9392,N_9305);
and U11866 (N_11866,N_9654,N_9513);
nor U11867 (N_11867,N_10130,N_9797);
nand U11868 (N_11868,N_10299,N_9914);
or U11869 (N_11869,N_9865,N_9824);
or U11870 (N_11870,N_10163,N_10059);
and U11871 (N_11871,N_9553,N_9459);
or U11872 (N_11872,N_9191,N_9547);
nand U11873 (N_11873,N_10413,N_9767);
and U11874 (N_11874,N_9641,N_9422);
nor U11875 (N_11875,N_9791,N_10385);
and U11876 (N_11876,N_10440,N_10106);
nand U11877 (N_11877,N_10075,N_9508);
nor U11878 (N_11878,N_10303,N_9640);
nor U11879 (N_11879,N_9980,N_10137);
nor U11880 (N_11880,N_9705,N_9212);
or U11881 (N_11881,N_9591,N_9166);
nand U11882 (N_11882,N_10483,N_10404);
nor U11883 (N_11883,N_9952,N_9269);
and U11884 (N_11884,N_10118,N_10336);
or U11885 (N_11885,N_9876,N_9277);
nor U11886 (N_11886,N_9872,N_9725);
and U11887 (N_11887,N_9540,N_9824);
or U11888 (N_11888,N_9311,N_9856);
xnor U11889 (N_11889,N_9428,N_9121);
nor U11890 (N_11890,N_10454,N_9959);
or U11891 (N_11891,N_10442,N_10082);
xor U11892 (N_11892,N_10477,N_9442);
nor U11893 (N_11893,N_10159,N_9715);
or U11894 (N_11894,N_9521,N_9441);
nor U11895 (N_11895,N_10225,N_9411);
nor U11896 (N_11896,N_10325,N_9595);
and U11897 (N_11897,N_9336,N_10179);
nor U11898 (N_11898,N_10471,N_9858);
or U11899 (N_11899,N_9724,N_9357);
xor U11900 (N_11900,N_9657,N_9421);
nand U11901 (N_11901,N_9249,N_10075);
xnor U11902 (N_11902,N_9105,N_9444);
nor U11903 (N_11903,N_10060,N_9169);
and U11904 (N_11904,N_9077,N_10299);
or U11905 (N_11905,N_9453,N_9613);
nor U11906 (N_11906,N_9705,N_10456);
and U11907 (N_11907,N_9613,N_10327);
nor U11908 (N_11908,N_9974,N_10158);
xnor U11909 (N_11909,N_9514,N_10175);
or U11910 (N_11910,N_9600,N_9807);
and U11911 (N_11911,N_9998,N_10279);
nand U11912 (N_11912,N_10247,N_9471);
nor U11913 (N_11913,N_9635,N_9318);
nand U11914 (N_11914,N_9718,N_9330);
nand U11915 (N_11915,N_9231,N_10172);
or U11916 (N_11916,N_9649,N_9931);
nand U11917 (N_11917,N_9838,N_10131);
nor U11918 (N_11918,N_10260,N_9808);
nor U11919 (N_11919,N_9019,N_9531);
nand U11920 (N_11920,N_9511,N_10340);
nand U11921 (N_11921,N_9672,N_9690);
nor U11922 (N_11922,N_9290,N_9949);
or U11923 (N_11923,N_9247,N_9185);
or U11924 (N_11924,N_9084,N_9773);
nor U11925 (N_11925,N_9295,N_9101);
xor U11926 (N_11926,N_9572,N_9561);
nor U11927 (N_11927,N_10295,N_9419);
nor U11928 (N_11928,N_9268,N_10118);
nor U11929 (N_11929,N_10357,N_10446);
and U11930 (N_11930,N_10104,N_9377);
nand U11931 (N_11931,N_10305,N_9717);
nand U11932 (N_11932,N_10207,N_9733);
or U11933 (N_11933,N_10406,N_9154);
nor U11934 (N_11934,N_9932,N_9224);
nor U11935 (N_11935,N_9569,N_9484);
and U11936 (N_11936,N_9892,N_9100);
or U11937 (N_11937,N_9492,N_9626);
nand U11938 (N_11938,N_10063,N_9243);
xnor U11939 (N_11939,N_9642,N_9634);
nor U11940 (N_11940,N_10198,N_9272);
xor U11941 (N_11941,N_9277,N_10263);
and U11942 (N_11942,N_9737,N_9094);
and U11943 (N_11943,N_9454,N_10400);
xor U11944 (N_11944,N_9457,N_9132);
nand U11945 (N_11945,N_9744,N_9160);
nor U11946 (N_11946,N_10166,N_9419);
or U11947 (N_11947,N_10213,N_9051);
or U11948 (N_11948,N_9242,N_9786);
nand U11949 (N_11949,N_9039,N_9471);
nand U11950 (N_11950,N_9968,N_9681);
nand U11951 (N_11951,N_9041,N_9531);
and U11952 (N_11952,N_9696,N_9478);
nor U11953 (N_11953,N_9682,N_9867);
nand U11954 (N_11954,N_10375,N_9917);
xor U11955 (N_11955,N_9535,N_9086);
and U11956 (N_11956,N_9255,N_10157);
nand U11957 (N_11957,N_9696,N_9368);
and U11958 (N_11958,N_9573,N_10480);
xor U11959 (N_11959,N_10177,N_10001);
nand U11960 (N_11960,N_10049,N_10298);
nor U11961 (N_11961,N_9677,N_9133);
nor U11962 (N_11962,N_9824,N_9204);
or U11963 (N_11963,N_9156,N_10395);
or U11964 (N_11964,N_10401,N_9470);
nand U11965 (N_11965,N_10035,N_10455);
and U11966 (N_11966,N_10463,N_10197);
or U11967 (N_11967,N_9730,N_9133);
nand U11968 (N_11968,N_9917,N_9848);
and U11969 (N_11969,N_9244,N_9339);
nor U11970 (N_11970,N_10129,N_9361);
nor U11971 (N_11971,N_10299,N_9612);
nand U11972 (N_11972,N_10191,N_9620);
nor U11973 (N_11973,N_9390,N_9485);
nor U11974 (N_11974,N_10016,N_9808);
nor U11975 (N_11975,N_9417,N_10215);
nand U11976 (N_11976,N_9094,N_9444);
nor U11977 (N_11977,N_9417,N_9600);
or U11978 (N_11978,N_9760,N_10288);
and U11979 (N_11979,N_9021,N_9123);
nand U11980 (N_11980,N_10265,N_9552);
or U11981 (N_11981,N_10036,N_10396);
and U11982 (N_11982,N_9464,N_9026);
nand U11983 (N_11983,N_9540,N_10016);
and U11984 (N_11984,N_9413,N_9498);
or U11985 (N_11985,N_10290,N_9998);
or U11986 (N_11986,N_10384,N_10087);
nor U11987 (N_11987,N_10439,N_9347);
or U11988 (N_11988,N_10289,N_9118);
nand U11989 (N_11989,N_10099,N_10221);
nor U11990 (N_11990,N_10474,N_9354);
or U11991 (N_11991,N_9658,N_10394);
nand U11992 (N_11992,N_10022,N_10144);
nand U11993 (N_11993,N_10273,N_10201);
and U11994 (N_11994,N_9295,N_10424);
or U11995 (N_11995,N_9433,N_10478);
nand U11996 (N_11996,N_9066,N_9754);
xnor U11997 (N_11997,N_10444,N_9087);
and U11998 (N_11998,N_9326,N_9845);
nor U11999 (N_11999,N_9375,N_10286);
xor U12000 (N_12000,N_10785,N_10530);
nor U12001 (N_12001,N_10841,N_11765);
and U12002 (N_12002,N_11528,N_11881);
and U12003 (N_12003,N_11076,N_11092);
nand U12004 (N_12004,N_11542,N_11417);
or U12005 (N_12005,N_11415,N_11554);
nand U12006 (N_12006,N_11886,N_10673);
nor U12007 (N_12007,N_10784,N_11123);
nor U12008 (N_12008,N_11357,N_10995);
nand U12009 (N_12009,N_10691,N_11520);
nand U12010 (N_12010,N_11572,N_11160);
nand U12011 (N_12011,N_11151,N_10652);
nor U12012 (N_12012,N_11606,N_11477);
and U12013 (N_12013,N_10651,N_11490);
nor U12014 (N_12014,N_11804,N_10952);
nor U12015 (N_12015,N_11124,N_10970);
nor U12016 (N_12016,N_10735,N_10982);
nand U12017 (N_12017,N_11799,N_11147);
nand U12018 (N_12018,N_10722,N_11228);
and U12019 (N_12019,N_11567,N_11855);
xor U12020 (N_12020,N_11494,N_11755);
nor U12021 (N_12021,N_10867,N_10806);
nand U12022 (N_12022,N_11717,N_11693);
nor U12023 (N_12023,N_11183,N_11125);
xnor U12024 (N_12024,N_11075,N_10762);
nor U12025 (N_12025,N_11743,N_11121);
nand U12026 (N_12026,N_11928,N_10829);
nor U12027 (N_12027,N_11847,N_10577);
nand U12028 (N_12028,N_10976,N_11229);
nand U12029 (N_12029,N_11396,N_11754);
nor U12030 (N_12030,N_11346,N_11029);
and U12031 (N_12031,N_11421,N_11940);
nand U12032 (N_12032,N_11858,N_10950);
nand U12033 (N_12033,N_10587,N_11478);
nand U12034 (N_12034,N_10925,N_11563);
or U12035 (N_12035,N_11500,N_11390);
nand U12036 (N_12036,N_11854,N_11335);
and U12037 (N_12037,N_11305,N_10749);
nand U12038 (N_12038,N_11319,N_11053);
nand U12039 (N_12039,N_11734,N_10921);
xor U12040 (N_12040,N_10707,N_11094);
nand U12041 (N_12041,N_11808,N_11742);
or U12042 (N_12042,N_10657,N_10541);
or U12043 (N_12043,N_11920,N_10716);
or U12044 (N_12044,N_11677,N_11973);
and U12045 (N_12045,N_11043,N_11317);
nor U12046 (N_12046,N_10932,N_10622);
or U12047 (N_12047,N_11988,N_11455);
and U12048 (N_12048,N_11785,N_11066);
nand U12049 (N_12049,N_10824,N_11543);
or U12050 (N_12050,N_11974,N_11087);
xnor U12051 (N_12051,N_11320,N_11152);
nor U12052 (N_12052,N_11877,N_10771);
or U12053 (N_12053,N_10708,N_10682);
or U12054 (N_12054,N_11897,N_11284);
and U12055 (N_12055,N_11458,N_11360);
nor U12056 (N_12056,N_11022,N_11459);
nor U12057 (N_12057,N_11081,N_11953);
or U12058 (N_12058,N_10635,N_11907);
or U12059 (N_12059,N_11442,N_11522);
nor U12060 (N_12060,N_11583,N_11084);
or U12061 (N_12061,N_11883,N_11800);
and U12062 (N_12062,N_11351,N_10798);
and U12063 (N_12063,N_10944,N_10947);
nor U12064 (N_12064,N_11828,N_11960);
or U12065 (N_12065,N_11185,N_10757);
nor U12066 (N_12066,N_10849,N_11986);
xor U12067 (N_12067,N_11674,N_11110);
nor U12068 (N_12068,N_11817,N_11611);
nor U12069 (N_12069,N_10594,N_10988);
or U12070 (N_12070,N_11336,N_10540);
or U12071 (N_12071,N_11873,N_11661);
or U12072 (N_12072,N_11392,N_11069);
nand U12073 (N_12073,N_10552,N_11777);
xnor U12074 (N_12074,N_11130,N_11689);
or U12075 (N_12075,N_11891,N_10667);
and U12076 (N_12076,N_10690,N_11451);
or U12077 (N_12077,N_10868,N_11599);
nand U12078 (N_12078,N_11719,N_10669);
nor U12079 (N_12079,N_10737,N_11802);
or U12080 (N_12080,N_10767,N_11238);
or U12081 (N_12081,N_11007,N_10583);
nor U12082 (N_12082,N_11795,N_11767);
xnor U12083 (N_12083,N_11791,N_11862);
nand U12084 (N_12084,N_11419,N_11837);
and U12085 (N_12085,N_10949,N_11105);
and U12086 (N_12086,N_10763,N_10775);
or U12087 (N_12087,N_11622,N_10608);
nor U12088 (N_12088,N_10980,N_10727);
nand U12089 (N_12089,N_11435,N_11996);
and U12090 (N_12090,N_11325,N_11958);
and U12091 (N_12091,N_11057,N_11656);
and U12092 (N_12092,N_11327,N_10968);
or U12093 (N_12093,N_11710,N_11385);
or U12094 (N_12094,N_11021,N_11954);
nor U12095 (N_12095,N_10693,N_11205);
and U12096 (N_12096,N_10686,N_11998);
or U12097 (N_12097,N_11863,N_11261);
nor U12098 (N_12098,N_10597,N_11736);
nand U12099 (N_12099,N_11727,N_10927);
or U12100 (N_12100,N_11722,N_11384);
nand U12101 (N_12101,N_11363,N_11010);
and U12102 (N_12102,N_11990,N_11332);
nor U12103 (N_12103,N_11356,N_10565);
nor U12104 (N_12104,N_11640,N_11507);
or U12105 (N_12105,N_10698,N_11602);
nand U12106 (N_12106,N_11341,N_11989);
or U12107 (N_12107,N_11673,N_11801);
nand U12108 (N_12108,N_11070,N_11564);
or U12109 (N_12109,N_11823,N_11516);
and U12110 (N_12110,N_11005,N_11546);
or U12111 (N_12111,N_10629,N_11790);
or U12112 (N_12112,N_11118,N_11184);
nand U12113 (N_12113,N_11927,N_10514);
and U12114 (N_12114,N_10604,N_10502);
and U12115 (N_12115,N_11334,N_11464);
nand U12116 (N_12116,N_11272,N_10788);
nor U12117 (N_12117,N_10526,N_10522);
or U12118 (N_12118,N_11950,N_11245);
nand U12119 (N_12119,N_11432,N_11333);
nand U12120 (N_12120,N_11864,N_11122);
xnor U12121 (N_12121,N_10518,N_11844);
nor U12122 (N_12122,N_11687,N_10534);
or U12123 (N_12123,N_11354,N_11294);
and U12124 (N_12124,N_11058,N_11046);
xnor U12125 (N_12125,N_10973,N_11174);
nor U12126 (N_12126,N_10853,N_10625);
and U12127 (N_12127,N_11951,N_11193);
and U12128 (N_12128,N_10825,N_10769);
xnor U12129 (N_12129,N_11575,N_11299);
and U12130 (N_12130,N_11904,N_11237);
and U12131 (N_12131,N_11461,N_11982);
or U12132 (N_12132,N_11283,N_11915);
or U12133 (N_12133,N_11665,N_11642);
nor U12134 (N_12134,N_10515,N_11222);
nand U12135 (N_12135,N_11439,N_10633);
or U12136 (N_12136,N_11582,N_11629);
xor U12137 (N_12137,N_11170,N_10566);
or U12138 (N_12138,N_11874,N_11530);
nor U12139 (N_12139,N_10679,N_10712);
nor U12140 (N_12140,N_11475,N_11579);
nand U12141 (N_12141,N_11977,N_11639);
nand U12142 (N_12142,N_11497,N_11890);
nand U12143 (N_12143,N_11078,N_10855);
or U12144 (N_12144,N_11524,N_11420);
nand U12145 (N_12145,N_10713,N_11924);
nand U12146 (N_12146,N_11779,N_10505);
nor U12147 (N_12147,N_11748,N_10555);
nand U12148 (N_12148,N_10850,N_10525);
and U12149 (N_12149,N_10974,N_11410);
or U12150 (N_12150,N_11379,N_11145);
and U12151 (N_12151,N_10744,N_11882);
nor U12152 (N_12152,N_11889,N_11538);
and U12153 (N_12153,N_11816,N_10766);
xor U12154 (N_12154,N_11428,N_10684);
or U12155 (N_12155,N_11342,N_11708);
nor U12156 (N_12156,N_11098,N_10787);
or U12157 (N_12157,N_10781,N_11782);
or U12158 (N_12158,N_11964,N_11600);
and U12159 (N_12159,N_10697,N_11408);
or U12160 (N_12160,N_11578,N_11389);
nand U12161 (N_12161,N_10613,N_10985);
xnor U12162 (N_12162,N_11252,N_10987);
nor U12163 (N_12163,N_10848,N_10902);
or U12164 (N_12164,N_11655,N_11565);
nand U12165 (N_12165,N_10998,N_10883);
and U12166 (N_12166,N_10827,N_10546);
or U12167 (N_12167,N_11702,N_11745);
and U12168 (N_12168,N_10562,N_11949);
or U12169 (N_12169,N_11993,N_11362);
nor U12170 (N_12170,N_11095,N_10695);
or U12171 (N_12171,N_10983,N_11654);
xor U12172 (N_12172,N_11116,N_11628);
or U12173 (N_12173,N_11444,N_11574);
nand U12174 (N_12174,N_11613,N_11171);
nor U12175 (N_12175,N_11047,N_11876);
and U12176 (N_12176,N_11248,N_11089);
nand U12177 (N_12177,N_10903,N_11287);
xor U12178 (N_12178,N_11310,N_11880);
and U12179 (N_12179,N_11285,N_11201);
or U12180 (N_12180,N_10680,N_11433);
nor U12181 (N_12181,N_10752,N_10551);
nor U12182 (N_12182,N_11418,N_11209);
or U12183 (N_12183,N_10646,N_11086);
or U12184 (N_12184,N_10598,N_11311);
or U12185 (N_12185,N_10705,N_10601);
nor U12186 (N_12186,N_10978,N_11840);
xnor U12187 (N_12187,N_11634,N_10586);
nor U12188 (N_12188,N_11371,N_11809);
or U12189 (N_12189,N_11407,N_10751);
or U12190 (N_12190,N_11853,N_11207);
nand U12191 (N_12191,N_11117,N_11741);
and U12192 (N_12192,N_10638,N_11593);
and U12193 (N_12193,N_10828,N_10731);
or U12194 (N_12194,N_10840,N_10585);
xnor U12195 (N_12195,N_11612,N_11120);
and U12196 (N_12196,N_11830,N_10563);
or U12197 (N_12197,N_11035,N_11902);
nor U12198 (N_12198,N_11644,N_11353);
nand U12199 (N_12199,N_10928,N_11377);
or U12200 (N_12200,N_11413,N_11769);
nor U12201 (N_12201,N_10797,N_10761);
xor U12202 (N_12202,N_11916,N_11825);
and U12203 (N_12203,N_11839,N_11023);
and U12204 (N_12204,N_10871,N_11957);
or U12205 (N_12205,N_10734,N_11188);
nor U12206 (N_12206,N_11537,N_10953);
and U12207 (N_12207,N_10723,N_11345);
or U12208 (N_12208,N_10627,N_10882);
nand U12209 (N_12209,N_11621,N_11426);
or U12210 (N_12210,N_10508,N_11848);
nand U12211 (N_12211,N_10663,N_11079);
xnor U12212 (N_12212,N_11859,N_11934);
or U12213 (N_12213,N_11939,N_11082);
nand U12214 (N_12214,N_11756,N_10821);
nand U12215 (N_12215,N_11908,N_10813);
or U12216 (N_12216,N_11618,N_11162);
nand U12217 (N_12217,N_11893,N_11725);
nand U12218 (N_12218,N_11187,N_11259);
and U12219 (N_12219,N_10802,N_11555);
and U12220 (N_12220,N_11318,N_10880);
or U12221 (N_12221,N_11309,N_11609);
xnor U12222 (N_12222,N_11256,N_10990);
nor U12223 (N_12223,N_10791,N_11774);
nand U12224 (N_12224,N_11994,N_10611);
nand U12225 (N_12225,N_11645,N_11393);
nor U12226 (N_12226,N_11922,N_11836);
nand U12227 (N_12227,N_11300,N_11324);
nand U12228 (N_12228,N_11894,N_11165);
xnor U12229 (N_12229,N_11589,N_11937);
xnor U12230 (N_12230,N_11941,N_11984);
nand U12231 (N_12231,N_10852,N_11368);
nor U12232 (N_12232,N_10847,N_10694);
nor U12233 (N_12233,N_10543,N_10794);
xor U12234 (N_12234,N_11868,N_10639);
and U12235 (N_12235,N_10864,N_11008);
xnor U12236 (N_12236,N_10873,N_10936);
and U12237 (N_12237,N_11040,N_10975);
nand U12238 (N_12238,N_10571,N_11995);
nand U12239 (N_12239,N_11210,N_10759);
or U12240 (N_12240,N_10897,N_11987);
and U12241 (N_12241,N_10659,N_11849);
nor U12242 (N_12242,N_11380,N_11753);
nand U12243 (N_12243,N_11322,N_11314);
or U12244 (N_12244,N_10596,N_11244);
nor U12245 (N_12245,N_11664,N_11587);
nor U12246 (N_12246,N_11813,N_11036);
nand U12247 (N_12247,N_11113,N_11153);
xnor U12248 (N_12248,N_10938,N_11293);
nand U12249 (N_12249,N_11780,N_11400);
or U12250 (N_12250,N_11714,N_10913);
nand U12251 (N_12251,N_11747,N_10881);
nand U12252 (N_12252,N_11107,N_11604);
nor U12253 (N_12253,N_10580,N_10736);
nor U12254 (N_12254,N_10959,N_10812);
nand U12255 (N_12255,N_10768,N_11879);
and U12256 (N_12256,N_11000,N_11292);
nor U12257 (N_12257,N_10689,N_11423);
xnor U12258 (N_12258,N_11221,N_10786);
nand U12259 (N_12259,N_11718,N_10600);
nor U12260 (N_12260,N_11189,N_11387);
and U12261 (N_12261,N_11649,N_11484);
nor U12262 (N_12262,N_11919,N_10636);
or U12263 (N_12263,N_11243,N_10529);
or U12264 (N_12264,N_10746,N_11097);
nor U12265 (N_12265,N_10656,N_10739);
nand U12266 (N_12266,N_10887,N_10780);
or U12267 (N_12267,N_11457,N_11493);
nor U12268 (N_12268,N_10892,N_11947);
nand U12269 (N_12269,N_11071,N_11447);
nor U12270 (N_12270,N_11898,N_11758);
and U12271 (N_12271,N_11626,N_11297);
or U12272 (N_12272,N_11044,N_11704);
nor U12273 (N_12273,N_11992,N_11946);
or U12274 (N_12274,N_10832,N_10889);
or U12275 (N_12275,N_11014,N_10618);
nand U12276 (N_12276,N_10547,N_10807);
nand U12277 (N_12277,N_11394,N_10803);
xnor U12278 (N_12278,N_11106,N_10750);
and U12279 (N_12279,N_10859,N_11503);
and U12280 (N_12280,N_11614,N_11899);
or U12281 (N_12281,N_10935,N_10896);
nor U12282 (N_12282,N_10733,N_11405);
or U12283 (N_12283,N_10623,N_10692);
nand U12284 (N_12284,N_11676,N_11531);
nand U12285 (N_12285,N_10632,N_11506);
xor U12286 (N_12286,N_11104,N_11139);
nor U12287 (N_12287,N_11340,N_11246);
xor U12288 (N_12288,N_10919,N_11486);
or U12289 (N_12289,N_10711,N_11111);
nand U12290 (N_12290,N_11647,N_11910);
nor U12291 (N_12291,N_11026,N_11195);
and U12292 (N_12292,N_10658,N_11527);
and U12293 (N_12293,N_11746,N_11250);
nor U12294 (N_12294,N_10992,N_11397);
nand U12295 (N_12295,N_11027,N_11766);
nor U12296 (N_12296,N_10612,N_10776);
or U12297 (N_12297,N_11502,N_11063);
nand U12298 (N_12298,N_11961,N_11279);
and U12299 (N_12299,N_10877,N_10875);
nand U12300 (N_12300,N_10719,N_11818);
nor U12301 (N_12301,N_10643,N_10854);
xor U12302 (N_12302,N_10810,N_11424);
or U12303 (N_12303,N_11257,N_11471);
nand U12304 (N_12304,N_10701,N_10677);
nor U12305 (N_12305,N_10537,N_11896);
nand U12306 (N_12306,N_11739,N_11381);
nor U12307 (N_12307,N_11892,N_10842);
and U12308 (N_12308,N_11338,N_11018);
xnor U12309 (N_12309,N_11675,N_11968);
and U12310 (N_12310,N_11487,N_10792);
and U12311 (N_12311,N_11306,N_11806);
or U12312 (N_12312,N_11573,N_11692);
or U12313 (N_12313,N_10557,N_10961);
nand U12314 (N_12314,N_11616,N_11406);
and U12315 (N_12315,N_10650,N_10564);
nand U12316 (N_12316,N_10614,N_10574);
and U12317 (N_12317,N_10939,N_11751);
and U12318 (N_12318,N_11048,N_10872);
and U12319 (N_12319,N_11814,N_10524);
nor U12320 (N_12320,N_10645,N_11607);
and U12321 (N_12321,N_11700,N_11921);
and U12322 (N_12322,N_11352,N_11277);
nand U12323 (N_12323,N_10581,N_11526);
and U12324 (N_12324,N_10815,N_10715);
and U12325 (N_12325,N_11196,N_11498);
nand U12326 (N_12326,N_11672,N_11878);
and U12327 (N_12327,N_11265,N_11776);
or U12328 (N_12328,N_11615,N_10906);
nor U12329 (N_12329,N_10706,N_11308);
or U12330 (N_12330,N_10826,N_11803);
or U12331 (N_12331,N_11476,N_11952);
nor U12332 (N_12332,N_11559,N_11138);
nor U12333 (N_12333,N_10642,N_11343);
xnor U12334 (N_12334,N_10703,N_10820);
or U12335 (N_12335,N_11370,N_10770);
and U12336 (N_12336,N_11128,N_10894);
xnor U12337 (N_12337,N_10989,N_11784);
nand U12338 (N_12338,N_11833,N_11824);
or U12339 (N_12339,N_10945,N_11796);
and U12340 (N_12340,N_11001,N_11942);
nand U12341 (N_12341,N_10589,N_11401);
or U12342 (N_12342,N_10620,N_11669);
and U12343 (N_12343,N_10640,N_10728);
and U12344 (N_12344,N_11594,N_11212);
xnor U12345 (N_12345,N_10899,N_11298);
nand U12346 (N_12346,N_10511,N_11083);
nand U12347 (N_12347,N_10649,N_11798);
xor U12348 (N_12348,N_10915,N_11180);
and U12349 (N_12349,N_10575,N_11545);
or U12350 (N_12350,N_11678,N_10923);
and U12351 (N_12351,N_11786,N_11101);
nor U12352 (N_12352,N_10777,N_10765);
and U12353 (N_12353,N_11970,N_11247);
or U12354 (N_12354,N_11025,N_11466);
nand U12355 (N_12355,N_11013,N_11096);
or U12356 (N_12356,N_10665,N_10683);
nor U12357 (N_12357,N_10929,N_11499);
nor U12358 (N_12358,N_11670,N_11686);
or U12359 (N_12359,N_10616,N_11763);
or U12360 (N_12360,N_10960,N_11489);
and U12361 (N_12361,N_10630,N_11701);
or U12362 (N_12362,N_11275,N_10972);
nor U12363 (N_12363,N_10800,N_11374);
nor U12364 (N_12364,N_11625,N_10560);
or U12365 (N_12365,N_11440,N_10696);
nor U12366 (N_12366,N_10941,N_10648);
nand U12367 (N_12367,N_11793,N_11659);
nand U12368 (N_12368,N_11268,N_11633);
and U12369 (N_12369,N_11636,N_11015);
nor U12370 (N_12370,N_11909,N_10957);
nand U12371 (N_12371,N_10940,N_10607);
nor U12372 (N_12372,N_11359,N_10861);
and U12373 (N_12373,N_10545,N_11684);
and U12374 (N_12374,N_10532,N_11286);
nor U12375 (N_12375,N_11382,N_11752);
or U12376 (N_12376,N_10822,N_10789);
and U12377 (N_12377,N_11826,N_11276);
nand U12378 (N_12378,N_10535,N_11652);
or U12379 (N_12379,N_11794,N_10879);
nor U12380 (N_12380,N_10724,N_11031);
nor U12381 (N_12381,N_11177,N_11263);
xor U12382 (N_12382,N_11350,N_11975);
xor U12383 (N_12383,N_10504,N_11258);
or U12384 (N_12384,N_11789,N_10742);
or U12385 (N_12385,N_10914,N_11006);
and U12386 (N_12386,N_11827,N_11775);
nand U12387 (N_12387,N_11635,N_11991);
nand U12388 (N_12388,N_11773,N_11491);
nand U12389 (N_12389,N_11561,N_11867);
or U12390 (N_12390,N_10671,N_11199);
nand U12391 (N_12391,N_10745,N_11845);
nor U12392 (N_12392,N_11835,N_10506);
nand U12393 (N_12393,N_11509,N_11884);
nor U12394 (N_12394,N_11289,N_11980);
nor U12395 (N_12395,N_11721,N_11099);
or U12396 (N_12396,N_10740,N_11398);
nor U12397 (N_12397,N_10678,N_10895);
or U12398 (N_12398,N_11938,N_10704);
or U12399 (N_12399,N_10835,N_10907);
and U12400 (N_12400,N_10602,N_11744);
nor U12401 (N_12401,N_11969,N_11792);
nand U12402 (N_12402,N_10674,N_11032);
nor U12403 (N_12403,N_10778,N_10661);
nand U12404 (N_12404,N_10933,N_11157);
or U12405 (N_12405,N_11731,N_10956);
and U12406 (N_12406,N_11365,N_11706);
and U12407 (N_12407,N_11166,N_11651);
nor U12408 (N_12408,N_11781,N_11638);
nand U12409 (N_12409,N_10592,N_11643);
and U12410 (N_12410,N_10609,N_11936);
nor U12411 (N_12411,N_11641,N_11935);
nor U12412 (N_12412,N_11846,N_10573);
xnor U12413 (N_12413,N_10603,N_11366);
nand U12414 (N_12414,N_11402,N_11278);
xor U12415 (N_12415,N_11208,N_11525);
nor U12416 (N_12416,N_11586,N_11255);
nor U12417 (N_12417,N_10517,N_11231);
nor U12418 (N_12418,N_10539,N_10918);
xor U12419 (N_12419,N_11161,N_11077);
nand U12420 (N_12420,N_10688,N_11553);
nand U12421 (N_12421,N_11778,N_10743);
or U12422 (N_12422,N_11930,N_11198);
or U12423 (N_12423,N_11197,N_11011);
and U12424 (N_12424,N_11566,N_11601);
and U12425 (N_12425,N_11115,N_11730);
or U12426 (N_12426,N_11557,N_10624);
or U12427 (N_12427,N_10748,N_11720);
nor U12428 (N_12428,N_11663,N_11811);
nor U12429 (N_12429,N_10503,N_11028);
nor U12430 (N_12430,N_11711,N_10631);
nor U12431 (N_12431,N_11054,N_11312);
and U12432 (N_12432,N_11933,N_11430);
nand U12433 (N_12433,N_11585,N_10977);
nor U12434 (N_12434,N_11073,N_11158);
and U12435 (N_12435,N_11033,N_10533);
or U12436 (N_12436,N_11979,N_11852);
or U12437 (N_12437,N_11544,N_10931);
nand U12438 (N_12438,N_10668,N_11925);
and U12439 (N_12439,N_11416,N_11216);
nand U12440 (N_12440,N_11705,N_11367);
and U12441 (N_12441,N_11962,N_10513);
xnor U12442 (N_12442,N_11103,N_11482);
nand U12443 (N_12443,N_11729,N_11313);
xnor U12444 (N_12444,N_11735,N_10898);
and U12445 (N_12445,N_11631,N_10863);
nor U12446 (N_12446,N_11141,N_11945);
or U12447 (N_12447,N_11972,N_11349);
and U12448 (N_12448,N_10570,N_10790);
nand U12449 (N_12449,N_11218,N_11978);
nand U12450 (N_12450,N_10910,N_11241);
nand U12451 (N_12451,N_10804,N_10991);
or U12452 (N_12452,N_10610,N_11473);
or U12453 (N_12453,N_11182,N_10996);
and U12454 (N_12454,N_11965,N_11667);
nand U12455 (N_12455,N_10866,N_11843);
or U12456 (N_12456,N_10579,N_11049);
nand U12457 (N_12457,N_10922,N_11732);
nand U12458 (N_12458,N_11728,N_11723);
and U12459 (N_12459,N_11167,N_11142);
xnor U12460 (N_12460,N_11020,N_10655);
nor U12461 (N_12461,N_10979,N_11829);
and U12462 (N_12462,N_10754,N_11067);
or U12463 (N_12463,N_11963,N_11861);
xnor U12464 (N_12464,N_10818,N_11211);
or U12465 (N_12465,N_10865,N_11932);
or U12466 (N_12466,N_11348,N_11326);
nand U12467 (N_12467,N_10676,N_10599);
or U12468 (N_12468,N_11966,N_11347);
nor U12469 (N_12469,N_11173,N_11004);
nand U12470 (N_12470,N_11911,N_11917);
nand U12471 (N_12471,N_11155,N_11517);
or U12472 (N_12472,N_10836,N_11403);
nand U12473 (N_12473,N_10901,N_10860);
and U12474 (N_12474,N_10549,N_11648);
and U12475 (N_12475,N_10654,N_10521);
nand U12476 (N_12476,N_11623,N_11290);
and U12477 (N_12477,N_11434,N_10582);
and U12478 (N_12478,N_10559,N_10799);
xnor U12479 (N_12479,N_11483,N_11468);
nor U12480 (N_12480,N_10756,N_10550);
and U12481 (N_12481,N_11699,N_11501);
and U12482 (N_12482,N_10946,N_11671);
and U12483 (N_12483,N_10981,N_11851);
nor U12484 (N_12484,N_11203,N_11232);
xnor U12485 (N_12485,N_10523,N_11630);
nand U12486 (N_12486,N_10793,N_11361);
and U12487 (N_12487,N_10730,N_10764);
nand U12488 (N_12488,N_11787,N_10912);
or U12489 (N_12489,N_11658,N_11186);
nor U12490 (N_12490,N_11558,N_10954);
or U12491 (N_12491,N_11301,N_11569);
nor U12492 (N_12492,N_11088,N_11445);
nor U12493 (N_12493,N_11871,N_10984);
nor U12494 (N_12494,N_11280,N_10905);
nand U12495 (N_12495,N_11913,N_11163);
xor U12496 (N_12496,N_11900,N_11330);
or U12497 (N_12497,N_10885,N_11596);
nor U12498 (N_12498,N_10548,N_10997);
and U12499 (N_12499,N_10760,N_11632);
and U12500 (N_12500,N_11449,N_10725);
nand U12501 (N_12501,N_11515,N_11514);
nand U12502 (N_12502,N_11108,N_11591);
and U12503 (N_12503,N_11997,N_11831);
xor U12504 (N_12504,N_11291,N_10726);
or U12505 (N_12505,N_10536,N_10634);
or U12506 (N_12506,N_10773,N_11682);
or U12507 (N_12507,N_11137,N_11412);
nor U12508 (N_12508,N_11039,N_11529);
nand U12509 (N_12509,N_11749,N_10870);
xor U12510 (N_12510,N_10685,N_11556);
nand U12511 (N_12511,N_11761,N_11129);
nor U12512 (N_12512,N_11610,N_11093);
or U12513 (N_12513,N_11552,N_11427);
and U12514 (N_12514,N_11019,N_10908);
nor U12515 (N_12515,N_11885,N_10569);
or U12516 (N_12516,N_11136,N_11102);
nand U12517 (N_12517,N_10542,N_11038);
nor U12518 (N_12518,N_11668,N_11905);
or U12519 (N_12519,N_10510,N_11955);
nand U12520 (N_12520,N_11832,N_10702);
nand U12521 (N_12521,N_11737,N_11119);
or U12522 (N_12522,N_11926,N_10966);
nand U12523 (N_12523,N_10831,N_10805);
and U12524 (N_12524,N_10856,N_11548);
xor U12525 (N_12525,N_11901,N_10924);
nand U12526 (N_12526,N_11536,N_11738);
and U12527 (N_12527,N_11695,N_10869);
nand U12528 (N_12528,N_11856,N_11030);
and U12529 (N_12529,N_11154,N_11404);
or U12530 (N_12530,N_11650,N_11262);
nor U12531 (N_12531,N_10709,N_11764);
xor U12532 (N_12532,N_10590,N_11109);
and U12533 (N_12533,N_11592,N_11488);
or U12534 (N_12534,N_11712,N_10862);
nand U12535 (N_12535,N_10779,N_11757);
nand U12536 (N_12536,N_11707,N_11653);
nor U12537 (N_12537,N_11304,N_11269);
nand U12538 (N_12538,N_11090,N_10834);
and U12539 (N_12539,N_11146,N_10617);
nand U12540 (N_12540,N_11091,N_11462);
nand U12541 (N_12541,N_10556,N_10911);
nand U12542 (N_12542,N_11303,N_10930);
nand U12543 (N_12543,N_11441,N_11438);
and U12544 (N_12544,N_10738,N_10553);
or U12545 (N_12545,N_11156,N_11369);
or U12546 (N_12546,N_11590,N_11857);
or U12547 (N_12547,N_10886,N_10593);
or U12548 (N_12548,N_10558,N_11144);
nor U12549 (N_12549,N_10637,N_10544);
or U12550 (N_12550,N_11168,N_11452);
and U12551 (N_12551,N_10660,N_11666);
nand U12552 (N_12552,N_11697,N_11260);
nand U12553 (N_12553,N_11422,N_11074);
nand U12554 (N_12554,N_11581,N_11172);
nor U12555 (N_12555,N_11254,N_11194);
nand U12556 (N_12556,N_11505,N_10962);
and U12557 (N_12557,N_11976,N_11560);
and U12558 (N_12558,N_10884,N_11914);
or U12559 (N_12559,N_11282,N_11399);
nor U12560 (N_12560,N_10538,N_11617);
xor U12561 (N_12561,N_11223,N_10969);
nand U12562 (N_12562,N_10591,N_10846);
nor U12563 (N_12563,N_11535,N_10948);
nor U12564 (N_12564,N_10891,N_11133);
or U12565 (N_12565,N_11034,N_11227);
xor U12566 (N_12566,N_10500,N_10666);
nor U12567 (N_12567,N_10888,N_11495);
nand U12568 (N_12568,N_10999,N_11456);
and U12569 (N_12569,N_10527,N_11637);
nor U12570 (N_12570,N_11472,N_11562);
and U12571 (N_12571,N_11580,N_11740);
or U12572 (N_12572,N_11431,N_11364);
nand U12573 (N_12573,N_11295,N_11045);
or U12574 (N_12574,N_11923,N_11783);
or U12575 (N_12575,N_11355,N_11042);
or U12576 (N_12576,N_11050,N_10516);
nand U12577 (N_12577,N_10838,N_11713);
and U12578 (N_12578,N_10584,N_11344);
and U12579 (N_12579,N_11395,N_10965);
nor U12580 (N_12580,N_11576,N_11956);
nor U12581 (N_12581,N_11518,N_10830);
and U12582 (N_12582,N_10837,N_11331);
nand U12583 (N_12583,N_10675,N_11056);
or U12584 (N_12584,N_10942,N_10554);
and U12585 (N_12585,N_11903,N_10717);
nand U12586 (N_12586,N_11204,N_10782);
xor U12587 (N_12587,N_10851,N_10528);
nor U12588 (N_12588,N_11372,N_11485);
nand U12589 (N_12589,N_11540,N_11584);
or U12590 (N_12590,N_11999,N_10672);
nand U12591 (N_12591,N_10641,N_10809);
nand U12592 (N_12592,N_10900,N_11465);
and U12593 (N_12593,N_11131,N_11888);
and U12594 (N_12594,N_10520,N_10839);
nor U12595 (N_12595,N_11819,N_11062);
xor U12596 (N_12596,N_11126,N_11726);
nand U12597 (N_12597,N_10700,N_11577);
or U12598 (N_12598,N_11270,N_11061);
or U12599 (N_12599,N_11009,N_11264);
and U12600 (N_12600,N_10811,N_11383);
nor U12601 (N_12601,N_11912,N_11760);
and U12602 (N_12602,N_11437,N_10904);
and U12603 (N_12603,N_11681,N_11508);
and U12604 (N_12604,N_11213,N_10512);
xor U12605 (N_12605,N_10937,N_10519);
nor U12606 (N_12606,N_11603,N_10774);
or U12607 (N_12607,N_11024,N_10595);
nor U12608 (N_12608,N_10986,N_11971);
and U12609 (N_12609,N_11810,N_11688);
nand U12610 (N_12610,N_11453,N_11454);
nor U12611 (N_12611,N_10878,N_11179);
xnor U12612 (N_12612,N_10967,N_10844);
and U12613 (N_12613,N_10833,N_11967);
and U12614 (N_12614,N_11541,N_11175);
and U12615 (N_12615,N_11240,N_11328);
or U12616 (N_12616,N_11230,N_11226);
nor U12617 (N_12617,N_11178,N_11251);
or U12618 (N_12618,N_11085,N_11450);
xor U12619 (N_12619,N_11944,N_10567);
and U12620 (N_12620,N_11429,N_10994);
and U12621 (N_12621,N_11065,N_10653);
xor U12622 (N_12622,N_11872,N_11239);
and U12623 (N_12623,N_11164,N_11834);
nand U12624 (N_12624,N_10816,N_11519);
or U12625 (N_12625,N_10721,N_11691);
and U12626 (N_12626,N_10732,N_11055);
nand U12627 (N_12627,N_11150,N_11698);
nand U12628 (N_12628,N_11869,N_11134);
and U12629 (N_12629,N_10958,N_11807);
nor U12630 (N_12630,N_11135,N_11215);
and U12631 (N_12631,N_11064,N_10720);
nor U12632 (N_12632,N_11772,N_11598);
or U12633 (N_12633,N_10509,N_11820);
nand U12634 (N_12634,N_11660,N_11337);
nor U12635 (N_12635,N_11470,N_11192);
or U12636 (N_12636,N_11224,N_11549);
or U12637 (N_12637,N_10578,N_11225);
nand U12638 (N_12638,N_10963,N_11547);
and U12639 (N_12639,N_10619,N_10890);
and U12640 (N_12640,N_11895,N_11875);
nand U12641 (N_12641,N_11414,N_11512);
nand U12642 (N_12642,N_11267,N_11679);
nor U12643 (N_12643,N_11296,N_11588);
and U12644 (N_12644,N_10501,N_11838);
and U12645 (N_12645,N_10955,N_11657);
and U12646 (N_12646,N_10588,N_11985);
nor U12647 (N_12647,N_11202,N_10801);
nand U12648 (N_12648,N_11378,N_11842);
and U12649 (N_12649,N_11865,N_11504);
or U12650 (N_12650,N_11771,N_10741);
or U12651 (N_12651,N_11948,N_11812);
nor U12652 (N_12652,N_11929,N_11112);
nand U12653 (N_12653,N_11100,N_11041);
nor U12654 (N_12654,N_10909,N_10664);
or U12655 (N_12655,N_11143,N_11918);
and U12656 (N_12656,N_10917,N_11206);
nand U12657 (N_12657,N_11436,N_10758);
and U12658 (N_12658,N_11460,N_11510);
nor U12659 (N_12659,N_10572,N_11411);
or U12660 (N_12660,N_11140,N_11373);
or U12661 (N_12661,N_11608,N_11570);
and U12662 (N_12662,N_11219,N_11887);
nand U12663 (N_12663,N_10971,N_11242);
nor U12664 (N_12664,N_10576,N_11409);
or U12665 (N_12665,N_10615,N_11624);
nor U12666 (N_12666,N_11690,N_11822);
or U12667 (N_12667,N_10605,N_10943);
and U12668 (N_12668,N_10626,N_11376);
nand U12669 (N_12669,N_11051,N_11080);
or U12670 (N_12670,N_11709,N_11149);
xnor U12671 (N_12671,N_10710,N_11797);
and U12672 (N_12672,N_10561,N_11959);
nand U12673 (N_12673,N_10621,N_11513);
nor U12674 (N_12674,N_11323,N_11037);
and U12675 (N_12675,N_11266,N_11481);
or U12676 (N_12676,N_11002,N_11870);
nand U12677 (N_12677,N_11425,N_11492);
or U12678 (N_12678,N_11249,N_11467);
and U12679 (N_12679,N_10747,N_11068);
xnor U12680 (N_12680,N_11759,N_11605);
xor U12681 (N_12681,N_11943,N_11358);
and U12682 (N_12682,N_11480,N_11533);
nand U12683 (N_12683,N_10993,N_11683);
or U12684 (N_12684,N_11235,N_11860);
nand U12685 (N_12685,N_11288,N_11316);
xor U12686 (N_12686,N_10783,N_10876);
and U12687 (N_12687,N_10755,N_11217);
nand U12688 (N_12688,N_11696,N_10857);
xnor U12689 (N_12689,N_10916,N_10817);
and U12690 (N_12690,N_10951,N_11571);
xnor U12691 (N_12691,N_11768,N_10814);
or U12692 (N_12692,N_10845,N_10819);
nand U12693 (N_12693,N_10795,N_11595);
xor U12694 (N_12694,N_11733,N_11169);
or U12695 (N_12695,N_11568,N_11329);
nor U12696 (N_12696,N_10934,N_11532);
nor U12697 (N_12697,N_11200,N_10843);
and U12698 (N_12698,N_11302,N_11321);
or U12699 (N_12699,N_10568,N_11620);
nor U12700 (N_12700,N_11012,N_10699);
or U12701 (N_12701,N_10920,N_11072);
nand U12702 (N_12702,N_10628,N_11805);
or U12703 (N_12703,N_11551,N_10858);
or U12704 (N_12704,N_10823,N_10507);
nor U12705 (N_12705,N_11017,N_10729);
nand U12706 (N_12706,N_11176,N_10926);
or U12707 (N_12707,N_11234,N_11539);
nand U12708 (N_12708,N_11060,N_11339);
nor U12709 (N_12709,N_11474,N_11521);
and U12710 (N_12710,N_10964,N_11534);
and U12711 (N_12711,N_11236,N_10808);
or U12712 (N_12712,N_11315,N_11597);
nor U12713 (N_12713,N_11463,N_11479);
or U12714 (N_12714,N_10681,N_11443);
or U12715 (N_12715,N_10606,N_11788);
xor U12716 (N_12716,N_11715,N_11724);
and U12717 (N_12717,N_11114,N_11003);
nand U12718 (N_12718,N_10718,N_11448);
or U12719 (N_12719,N_11181,N_11906);
nand U12720 (N_12720,N_11821,N_11750);
or U12721 (N_12721,N_11190,N_11059);
nand U12722 (N_12722,N_11627,N_11127);
or U12723 (N_12723,N_11866,N_11496);
xor U12724 (N_12724,N_11931,N_10662);
nor U12725 (N_12725,N_11762,N_11981);
and U12726 (N_12726,N_10531,N_10753);
nand U12727 (N_12727,N_11694,N_11148);
nand U12728 (N_12728,N_10687,N_11815);
and U12729 (N_12729,N_11191,N_11703);
xnor U12730 (N_12730,N_11391,N_10772);
and U12731 (N_12731,N_11214,N_11446);
or U12732 (N_12732,N_10670,N_11386);
and U12733 (N_12733,N_11375,N_11716);
or U12734 (N_12734,N_11680,N_10647);
nand U12735 (N_12735,N_11511,N_11253);
nand U12736 (N_12736,N_11619,N_11523);
nor U12737 (N_12737,N_11685,N_11850);
xnor U12738 (N_12738,N_11983,N_10644);
nand U12739 (N_12739,N_10796,N_11016);
nor U12740 (N_12740,N_10893,N_10874);
nand U12741 (N_12741,N_11052,N_11841);
nor U12742 (N_12742,N_11274,N_11132);
nor U12743 (N_12743,N_11388,N_11662);
xnor U12744 (N_12744,N_11307,N_11233);
and U12745 (N_12745,N_11469,N_11646);
nand U12746 (N_12746,N_11220,N_10714);
and U12747 (N_12747,N_11271,N_11770);
and U12748 (N_12748,N_11281,N_11159);
nand U12749 (N_12749,N_11273,N_11550);
xnor U12750 (N_12750,N_11404,N_11012);
xnor U12751 (N_12751,N_11637,N_11608);
nand U12752 (N_12752,N_10510,N_10654);
or U12753 (N_12753,N_10583,N_11049);
nand U12754 (N_12754,N_11313,N_11235);
or U12755 (N_12755,N_10600,N_11494);
nor U12756 (N_12756,N_10911,N_11488);
and U12757 (N_12757,N_11323,N_10618);
nor U12758 (N_12758,N_11929,N_11011);
nand U12759 (N_12759,N_10663,N_11244);
or U12760 (N_12760,N_11376,N_10776);
or U12761 (N_12761,N_10518,N_10917);
or U12762 (N_12762,N_11182,N_11606);
nand U12763 (N_12763,N_11282,N_11459);
nand U12764 (N_12764,N_11256,N_10615);
nand U12765 (N_12765,N_10702,N_11894);
and U12766 (N_12766,N_11320,N_11780);
and U12767 (N_12767,N_11153,N_10512);
and U12768 (N_12768,N_10678,N_11539);
or U12769 (N_12769,N_11096,N_11130);
nand U12770 (N_12770,N_11884,N_10634);
xnor U12771 (N_12771,N_11077,N_11424);
nand U12772 (N_12772,N_10822,N_11290);
and U12773 (N_12773,N_10785,N_10504);
or U12774 (N_12774,N_11373,N_10770);
nand U12775 (N_12775,N_11544,N_11993);
nor U12776 (N_12776,N_11478,N_10562);
nand U12777 (N_12777,N_10939,N_11959);
xor U12778 (N_12778,N_11432,N_11554);
and U12779 (N_12779,N_11641,N_11484);
nand U12780 (N_12780,N_11856,N_11419);
or U12781 (N_12781,N_10663,N_11471);
nand U12782 (N_12782,N_11859,N_11664);
xor U12783 (N_12783,N_10630,N_11014);
and U12784 (N_12784,N_11833,N_11223);
and U12785 (N_12785,N_11550,N_11656);
and U12786 (N_12786,N_11426,N_11519);
and U12787 (N_12787,N_11932,N_10611);
nand U12788 (N_12788,N_10633,N_11180);
or U12789 (N_12789,N_10988,N_11577);
nand U12790 (N_12790,N_10832,N_11634);
or U12791 (N_12791,N_11902,N_11288);
xor U12792 (N_12792,N_11625,N_11298);
or U12793 (N_12793,N_11237,N_10622);
and U12794 (N_12794,N_11591,N_10924);
and U12795 (N_12795,N_11810,N_11133);
and U12796 (N_12796,N_10843,N_11482);
nand U12797 (N_12797,N_11374,N_11291);
nor U12798 (N_12798,N_10856,N_10724);
xnor U12799 (N_12799,N_11551,N_11017);
and U12800 (N_12800,N_11135,N_10974);
and U12801 (N_12801,N_11600,N_11980);
xnor U12802 (N_12802,N_10683,N_10705);
xor U12803 (N_12803,N_10509,N_11117);
nand U12804 (N_12804,N_11628,N_11177);
nand U12805 (N_12805,N_11889,N_10917);
or U12806 (N_12806,N_11251,N_10706);
and U12807 (N_12807,N_10659,N_10516);
and U12808 (N_12808,N_11068,N_11585);
nand U12809 (N_12809,N_11446,N_10703);
and U12810 (N_12810,N_11626,N_11325);
nor U12811 (N_12811,N_11356,N_11578);
nand U12812 (N_12812,N_11676,N_11988);
or U12813 (N_12813,N_11329,N_11721);
nand U12814 (N_12814,N_11815,N_11926);
and U12815 (N_12815,N_10621,N_10624);
nand U12816 (N_12816,N_10548,N_11706);
nand U12817 (N_12817,N_11432,N_11740);
and U12818 (N_12818,N_11415,N_10858);
and U12819 (N_12819,N_11026,N_11048);
nand U12820 (N_12820,N_11605,N_10527);
nand U12821 (N_12821,N_10617,N_10565);
and U12822 (N_12822,N_11619,N_10928);
and U12823 (N_12823,N_11719,N_11304);
nand U12824 (N_12824,N_11250,N_11490);
and U12825 (N_12825,N_11499,N_10907);
nand U12826 (N_12826,N_11155,N_11494);
nand U12827 (N_12827,N_11062,N_11138);
nor U12828 (N_12828,N_10934,N_11238);
nand U12829 (N_12829,N_11020,N_11684);
nand U12830 (N_12830,N_10901,N_10556);
and U12831 (N_12831,N_11602,N_10677);
xnor U12832 (N_12832,N_11409,N_11048);
nand U12833 (N_12833,N_11485,N_10901);
nand U12834 (N_12834,N_10610,N_10658);
nor U12835 (N_12835,N_11812,N_11406);
nor U12836 (N_12836,N_10571,N_10890);
xnor U12837 (N_12837,N_11918,N_11300);
nand U12838 (N_12838,N_11972,N_11561);
xnor U12839 (N_12839,N_10826,N_11644);
nand U12840 (N_12840,N_11442,N_10790);
or U12841 (N_12841,N_10871,N_11584);
nor U12842 (N_12842,N_11043,N_11397);
or U12843 (N_12843,N_11458,N_11744);
or U12844 (N_12844,N_11768,N_10551);
nand U12845 (N_12845,N_11113,N_10849);
nor U12846 (N_12846,N_10659,N_11500);
or U12847 (N_12847,N_10718,N_10808);
nor U12848 (N_12848,N_10983,N_11854);
and U12849 (N_12849,N_10538,N_10776);
nand U12850 (N_12850,N_11050,N_11421);
or U12851 (N_12851,N_10815,N_11991);
nand U12852 (N_12852,N_11269,N_10707);
xor U12853 (N_12853,N_10887,N_11808);
nor U12854 (N_12854,N_11059,N_10639);
nand U12855 (N_12855,N_11305,N_11291);
or U12856 (N_12856,N_11040,N_11383);
nor U12857 (N_12857,N_11802,N_11958);
and U12858 (N_12858,N_10728,N_11582);
nand U12859 (N_12859,N_10684,N_10677);
nand U12860 (N_12860,N_11328,N_10772);
xnor U12861 (N_12861,N_11340,N_11344);
nand U12862 (N_12862,N_11139,N_11968);
or U12863 (N_12863,N_11549,N_11215);
and U12864 (N_12864,N_11743,N_11658);
and U12865 (N_12865,N_11288,N_11141);
or U12866 (N_12866,N_10556,N_11319);
or U12867 (N_12867,N_10894,N_10741);
or U12868 (N_12868,N_10851,N_11997);
and U12869 (N_12869,N_11918,N_11468);
and U12870 (N_12870,N_10762,N_11619);
and U12871 (N_12871,N_11373,N_11993);
nor U12872 (N_12872,N_11194,N_11912);
or U12873 (N_12873,N_10511,N_10698);
nand U12874 (N_12874,N_10588,N_10822);
nor U12875 (N_12875,N_10823,N_11823);
xnor U12876 (N_12876,N_11781,N_10537);
nor U12877 (N_12877,N_10616,N_11114);
xnor U12878 (N_12878,N_11132,N_11005);
nor U12879 (N_12879,N_10539,N_11908);
nand U12880 (N_12880,N_10569,N_11152);
and U12881 (N_12881,N_11130,N_11184);
or U12882 (N_12882,N_11618,N_10987);
nand U12883 (N_12883,N_11761,N_11105);
or U12884 (N_12884,N_10540,N_11632);
nand U12885 (N_12885,N_10937,N_11210);
or U12886 (N_12886,N_11981,N_10507);
nand U12887 (N_12887,N_11538,N_11062);
or U12888 (N_12888,N_11754,N_11870);
nor U12889 (N_12889,N_11478,N_11452);
nand U12890 (N_12890,N_10681,N_11915);
nand U12891 (N_12891,N_10810,N_10679);
nand U12892 (N_12892,N_11542,N_11490);
nor U12893 (N_12893,N_11697,N_11497);
and U12894 (N_12894,N_11483,N_11042);
or U12895 (N_12895,N_11511,N_10783);
or U12896 (N_12896,N_11853,N_11713);
or U12897 (N_12897,N_11121,N_11994);
xnor U12898 (N_12898,N_11977,N_11226);
and U12899 (N_12899,N_11898,N_10642);
nand U12900 (N_12900,N_11121,N_11608);
nor U12901 (N_12901,N_10792,N_11593);
and U12902 (N_12902,N_10606,N_10744);
or U12903 (N_12903,N_10621,N_10623);
and U12904 (N_12904,N_11290,N_11242);
nor U12905 (N_12905,N_10729,N_10743);
or U12906 (N_12906,N_11418,N_10504);
or U12907 (N_12907,N_10565,N_11085);
nor U12908 (N_12908,N_10850,N_11442);
or U12909 (N_12909,N_11249,N_11567);
nand U12910 (N_12910,N_10622,N_11089);
nand U12911 (N_12911,N_11849,N_11645);
nor U12912 (N_12912,N_11148,N_11274);
nor U12913 (N_12913,N_10976,N_11851);
nor U12914 (N_12914,N_11544,N_10630);
and U12915 (N_12915,N_11932,N_11344);
or U12916 (N_12916,N_11432,N_11239);
nor U12917 (N_12917,N_11166,N_11407);
and U12918 (N_12918,N_10917,N_10845);
nor U12919 (N_12919,N_11888,N_10721);
nor U12920 (N_12920,N_11564,N_11107);
nand U12921 (N_12921,N_10644,N_10558);
nor U12922 (N_12922,N_11821,N_11826);
xnor U12923 (N_12923,N_10817,N_10999);
nand U12924 (N_12924,N_11223,N_10881);
nor U12925 (N_12925,N_10720,N_11807);
nand U12926 (N_12926,N_11617,N_11856);
nand U12927 (N_12927,N_11837,N_11317);
nor U12928 (N_12928,N_10779,N_10518);
and U12929 (N_12929,N_11736,N_11494);
nand U12930 (N_12930,N_11492,N_10664);
or U12931 (N_12931,N_11266,N_11653);
or U12932 (N_12932,N_11393,N_11360);
and U12933 (N_12933,N_10727,N_11104);
nand U12934 (N_12934,N_11523,N_11592);
and U12935 (N_12935,N_11955,N_11420);
and U12936 (N_12936,N_10930,N_11487);
or U12937 (N_12937,N_11683,N_11843);
nor U12938 (N_12938,N_10509,N_10979);
nand U12939 (N_12939,N_10653,N_10550);
nor U12940 (N_12940,N_10780,N_11634);
nand U12941 (N_12941,N_10706,N_10892);
or U12942 (N_12942,N_11692,N_11886);
or U12943 (N_12943,N_11754,N_11842);
nand U12944 (N_12944,N_11095,N_10898);
and U12945 (N_12945,N_10672,N_10799);
and U12946 (N_12946,N_11184,N_11110);
and U12947 (N_12947,N_10817,N_10806);
or U12948 (N_12948,N_10582,N_10852);
or U12949 (N_12949,N_11589,N_10695);
nand U12950 (N_12950,N_11990,N_11262);
or U12951 (N_12951,N_11623,N_10720);
and U12952 (N_12952,N_11726,N_11696);
or U12953 (N_12953,N_10795,N_11046);
or U12954 (N_12954,N_11316,N_11339);
nand U12955 (N_12955,N_10633,N_10668);
xor U12956 (N_12956,N_11054,N_11225);
xnor U12957 (N_12957,N_10864,N_11031);
nand U12958 (N_12958,N_11364,N_10683);
and U12959 (N_12959,N_10820,N_11796);
nand U12960 (N_12960,N_10985,N_10971);
and U12961 (N_12961,N_11784,N_11278);
nor U12962 (N_12962,N_11462,N_11771);
nand U12963 (N_12963,N_11592,N_10564);
nand U12964 (N_12964,N_11589,N_10820);
nor U12965 (N_12965,N_10863,N_10821);
nor U12966 (N_12966,N_11089,N_11037);
nor U12967 (N_12967,N_11934,N_10840);
nand U12968 (N_12968,N_11389,N_11911);
nand U12969 (N_12969,N_11867,N_11625);
nand U12970 (N_12970,N_10694,N_10713);
or U12971 (N_12971,N_10691,N_11695);
nand U12972 (N_12972,N_10593,N_10660);
and U12973 (N_12973,N_11049,N_11238);
nor U12974 (N_12974,N_10708,N_11913);
nor U12975 (N_12975,N_11547,N_11806);
or U12976 (N_12976,N_10651,N_11329);
nor U12977 (N_12977,N_11165,N_10625);
or U12978 (N_12978,N_11013,N_11192);
nand U12979 (N_12979,N_11967,N_11852);
nand U12980 (N_12980,N_11465,N_10752);
and U12981 (N_12981,N_11036,N_11918);
nand U12982 (N_12982,N_10847,N_11201);
or U12983 (N_12983,N_10723,N_10710);
or U12984 (N_12984,N_11070,N_11237);
xor U12985 (N_12985,N_10843,N_10746);
and U12986 (N_12986,N_11351,N_11478);
and U12987 (N_12987,N_11804,N_10791);
nand U12988 (N_12988,N_10581,N_11087);
or U12989 (N_12989,N_11239,N_11167);
nor U12990 (N_12990,N_11331,N_11205);
nor U12991 (N_12991,N_10708,N_11537);
and U12992 (N_12992,N_11113,N_10698);
nor U12993 (N_12993,N_10607,N_11862);
nor U12994 (N_12994,N_10887,N_11829);
nand U12995 (N_12995,N_11867,N_11914);
nand U12996 (N_12996,N_10523,N_11044);
or U12997 (N_12997,N_10852,N_11835);
and U12998 (N_12998,N_10572,N_10845);
xnor U12999 (N_12999,N_10730,N_11305);
nor U13000 (N_13000,N_11876,N_11917);
or U13001 (N_13001,N_10977,N_11321);
nor U13002 (N_13002,N_11924,N_11875);
xnor U13003 (N_13003,N_11269,N_11915);
nand U13004 (N_13004,N_10772,N_10817);
nand U13005 (N_13005,N_11400,N_10780);
nor U13006 (N_13006,N_11139,N_10642);
or U13007 (N_13007,N_10912,N_11487);
nand U13008 (N_13008,N_10870,N_10911);
and U13009 (N_13009,N_11239,N_10574);
nand U13010 (N_13010,N_11547,N_11762);
and U13011 (N_13011,N_11299,N_11007);
nor U13012 (N_13012,N_10668,N_10877);
xnor U13013 (N_13013,N_10615,N_11216);
nand U13014 (N_13014,N_11708,N_10984);
nand U13015 (N_13015,N_11312,N_11251);
or U13016 (N_13016,N_11574,N_11163);
nand U13017 (N_13017,N_11933,N_11894);
and U13018 (N_13018,N_10715,N_11519);
nor U13019 (N_13019,N_11503,N_10781);
nor U13020 (N_13020,N_10689,N_11055);
or U13021 (N_13021,N_11668,N_11530);
or U13022 (N_13022,N_10650,N_11539);
and U13023 (N_13023,N_11310,N_11862);
or U13024 (N_13024,N_11442,N_11674);
and U13025 (N_13025,N_10879,N_11556);
nor U13026 (N_13026,N_11243,N_11310);
and U13027 (N_13027,N_11156,N_10671);
and U13028 (N_13028,N_10516,N_11936);
or U13029 (N_13029,N_11684,N_10524);
and U13030 (N_13030,N_10658,N_11251);
nor U13031 (N_13031,N_11392,N_11015);
nor U13032 (N_13032,N_11073,N_11794);
or U13033 (N_13033,N_11018,N_10663);
and U13034 (N_13034,N_10624,N_10844);
or U13035 (N_13035,N_11694,N_11884);
nor U13036 (N_13036,N_11970,N_11272);
nor U13037 (N_13037,N_11358,N_10923);
or U13038 (N_13038,N_11310,N_11104);
nor U13039 (N_13039,N_11437,N_10745);
nor U13040 (N_13040,N_11293,N_11334);
and U13041 (N_13041,N_10886,N_10800);
nor U13042 (N_13042,N_10986,N_10798);
nand U13043 (N_13043,N_10816,N_10835);
nor U13044 (N_13044,N_11118,N_10872);
nand U13045 (N_13045,N_11957,N_10658);
or U13046 (N_13046,N_11832,N_11746);
or U13047 (N_13047,N_11488,N_11299);
and U13048 (N_13048,N_11879,N_11981);
and U13049 (N_13049,N_10752,N_10859);
and U13050 (N_13050,N_10632,N_11351);
nand U13051 (N_13051,N_11508,N_11808);
and U13052 (N_13052,N_10601,N_11222);
and U13053 (N_13053,N_11648,N_11070);
nor U13054 (N_13054,N_10898,N_11066);
nand U13055 (N_13055,N_11379,N_11794);
nor U13056 (N_13056,N_11250,N_11115);
and U13057 (N_13057,N_11211,N_10866);
or U13058 (N_13058,N_10719,N_11984);
and U13059 (N_13059,N_11320,N_11071);
nor U13060 (N_13060,N_11031,N_11585);
and U13061 (N_13061,N_11088,N_10727);
and U13062 (N_13062,N_11493,N_10612);
or U13063 (N_13063,N_10714,N_10545);
nand U13064 (N_13064,N_11529,N_10813);
and U13065 (N_13065,N_11468,N_11462);
nor U13066 (N_13066,N_10665,N_11706);
nor U13067 (N_13067,N_11323,N_10735);
nor U13068 (N_13068,N_11394,N_11982);
nor U13069 (N_13069,N_11198,N_11598);
or U13070 (N_13070,N_11304,N_11137);
or U13071 (N_13071,N_10745,N_11653);
nor U13072 (N_13072,N_11334,N_11717);
or U13073 (N_13073,N_11624,N_11341);
nand U13074 (N_13074,N_11946,N_11181);
or U13075 (N_13075,N_10667,N_11258);
nand U13076 (N_13076,N_11143,N_11028);
nand U13077 (N_13077,N_11569,N_11144);
nand U13078 (N_13078,N_11978,N_11432);
nand U13079 (N_13079,N_10992,N_11078);
or U13080 (N_13080,N_10625,N_11484);
nor U13081 (N_13081,N_11137,N_11481);
xnor U13082 (N_13082,N_11803,N_10550);
and U13083 (N_13083,N_10990,N_10768);
nor U13084 (N_13084,N_10882,N_11346);
and U13085 (N_13085,N_10615,N_11541);
or U13086 (N_13086,N_11831,N_11970);
nand U13087 (N_13087,N_11021,N_10672);
and U13088 (N_13088,N_11587,N_10817);
and U13089 (N_13089,N_11073,N_11765);
nor U13090 (N_13090,N_11786,N_11273);
nor U13091 (N_13091,N_10883,N_11194);
nor U13092 (N_13092,N_10595,N_11903);
nor U13093 (N_13093,N_10806,N_11636);
xnor U13094 (N_13094,N_11683,N_11108);
nand U13095 (N_13095,N_11774,N_10838);
nor U13096 (N_13096,N_11606,N_11173);
and U13097 (N_13097,N_10695,N_11158);
and U13098 (N_13098,N_11234,N_11137);
or U13099 (N_13099,N_10847,N_11147);
xor U13100 (N_13100,N_11951,N_10849);
or U13101 (N_13101,N_10825,N_11008);
nor U13102 (N_13102,N_11599,N_11712);
xor U13103 (N_13103,N_11675,N_10724);
xnor U13104 (N_13104,N_10864,N_11167);
or U13105 (N_13105,N_10657,N_10870);
xor U13106 (N_13106,N_11795,N_10893);
and U13107 (N_13107,N_11717,N_11259);
or U13108 (N_13108,N_11104,N_10756);
and U13109 (N_13109,N_11294,N_10969);
and U13110 (N_13110,N_11801,N_10575);
nor U13111 (N_13111,N_11538,N_10844);
nor U13112 (N_13112,N_11349,N_11060);
or U13113 (N_13113,N_11121,N_10637);
or U13114 (N_13114,N_11985,N_11057);
nand U13115 (N_13115,N_10955,N_11997);
and U13116 (N_13116,N_11291,N_10870);
nand U13117 (N_13117,N_11498,N_11110);
xor U13118 (N_13118,N_11026,N_11128);
and U13119 (N_13119,N_10710,N_11025);
and U13120 (N_13120,N_10589,N_11353);
nand U13121 (N_13121,N_11788,N_11663);
or U13122 (N_13122,N_11451,N_11250);
and U13123 (N_13123,N_10839,N_11290);
and U13124 (N_13124,N_10868,N_11192);
and U13125 (N_13125,N_10502,N_10991);
nor U13126 (N_13126,N_11349,N_10954);
and U13127 (N_13127,N_11795,N_11983);
nor U13128 (N_13128,N_11326,N_10594);
and U13129 (N_13129,N_11707,N_11807);
nor U13130 (N_13130,N_11131,N_11597);
nand U13131 (N_13131,N_11343,N_11266);
or U13132 (N_13132,N_11355,N_11056);
nor U13133 (N_13133,N_11060,N_11473);
xor U13134 (N_13134,N_11994,N_11553);
or U13135 (N_13135,N_11948,N_11449);
xor U13136 (N_13136,N_10847,N_11386);
nand U13137 (N_13137,N_10848,N_10792);
and U13138 (N_13138,N_10539,N_10503);
nand U13139 (N_13139,N_11051,N_11257);
or U13140 (N_13140,N_11546,N_10582);
nor U13141 (N_13141,N_10704,N_10818);
nor U13142 (N_13142,N_11033,N_10571);
xnor U13143 (N_13143,N_11608,N_11382);
and U13144 (N_13144,N_11620,N_10500);
nor U13145 (N_13145,N_11742,N_11038);
or U13146 (N_13146,N_11189,N_11476);
or U13147 (N_13147,N_11157,N_10701);
or U13148 (N_13148,N_11702,N_10929);
nor U13149 (N_13149,N_11515,N_11389);
nor U13150 (N_13150,N_10700,N_11736);
or U13151 (N_13151,N_11115,N_11818);
or U13152 (N_13152,N_11891,N_11963);
and U13153 (N_13153,N_11413,N_11846);
or U13154 (N_13154,N_10705,N_11500);
or U13155 (N_13155,N_11148,N_11920);
nand U13156 (N_13156,N_11132,N_10873);
nand U13157 (N_13157,N_11571,N_11155);
or U13158 (N_13158,N_11146,N_10874);
or U13159 (N_13159,N_11323,N_11047);
or U13160 (N_13160,N_11786,N_10560);
and U13161 (N_13161,N_11990,N_10512);
nand U13162 (N_13162,N_11274,N_10840);
or U13163 (N_13163,N_10554,N_11652);
nand U13164 (N_13164,N_10873,N_11818);
or U13165 (N_13165,N_10851,N_10906);
nand U13166 (N_13166,N_11765,N_10842);
nand U13167 (N_13167,N_10866,N_11145);
nor U13168 (N_13168,N_10638,N_11023);
nor U13169 (N_13169,N_10568,N_10896);
or U13170 (N_13170,N_11873,N_11354);
nand U13171 (N_13171,N_11668,N_11794);
and U13172 (N_13172,N_11307,N_11923);
and U13173 (N_13173,N_11731,N_11944);
nand U13174 (N_13174,N_11752,N_11456);
nor U13175 (N_13175,N_11582,N_11005);
nor U13176 (N_13176,N_11239,N_11864);
nand U13177 (N_13177,N_10807,N_11722);
or U13178 (N_13178,N_11491,N_11787);
and U13179 (N_13179,N_11785,N_11853);
or U13180 (N_13180,N_11554,N_10961);
or U13181 (N_13181,N_10792,N_11988);
nand U13182 (N_13182,N_11637,N_10745);
nand U13183 (N_13183,N_11051,N_11021);
and U13184 (N_13184,N_11167,N_11193);
nor U13185 (N_13185,N_11066,N_11253);
nor U13186 (N_13186,N_10667,N_11182);
and U13187 (N_13187,N_11631,N_10674);
nor U13188 (N_13188,N_10647,N_10638);
nor U13189 (N_13189,N_10641,N_11206);
nor U13190 (N_13190,N_11411,N_11070);
nand U13191 (N_13191,N_10588,N_11223);
xor U13192 (N_13192,N_10538,N_11257);
and U13193 (N_13193,N_10704,N_11509);
and U13194 (N_13194,N_10731,N_11986);
nand U13195 (N_13195,N_11073,N_11543);
xor U13196 (N_13196,N_11857,N_10773);
nand U13197 (N_13197,N_11340,N_10963);
or U13198 (N_13198,N_11100,N_11366);
nor U13199 (N_13199,N_11992,N_11748);
or U13200 (N_13200,N_11340,N_10900);
nand U13201 (N_13201,N_11934,N_11686);
and U13202 (N_13202,N_11194,N_10877);
nor U13203 (N_13203,N_11769,N_11946);
or U13204 (N_13204,N_10854,N_11213);
or U13205 (N_13205,N_11495,N_11271);
nand U13206 (N_13206,N_11296,N_11510);
or U13207 (N_13207,N_10842,N_11726);
or U13208 (N_13208,N_11064,N_10539);
or U13209 (N_13209,N_11125,N_11157);
nor U13210 (N_13210,N_11071,N_10677);
and U13211 (N_13211,N_11917,N_10615);
or U13212 (N_13212,N_10936,N_11422);
or U13213 (N_13213,N_11200,N_11193);
or U13214 (N_13214,N_11291,N_10678);
nor U13215 (N_13215,N_11019,N_10637);
nor U13216 (N_13216,N_11812,N_11063);
nor U13217 (N_13217,N_10877,N_11783);
xnor U13218 (N_13218,N_11202,N_11399);
nand U13219 (N_13219,N_10984,N_11508);
nor U13220 (N_13220,N_11718,N_10688);
xnor U13221 (N_13221,N_11979,N_11936);
or U13222 (N_13222,N_10644,N_10526);
nand U13223 (N_13223,N_11190,N_10875);
xnor U13224 (N_13224,N_10549,N_10992);
nand U13225 (N_13225,N_10965,N_11951);
and U13226 (N_13226,N_11622,N_11364);
nand U13227 (N_13227,N_11971,N_10831);
or U13228 (N_13228,N_11757,N_10526);
nand U13229 (N_13229,N_11854,N_11151);
nor U13230 (N_13230,N_11395,N_11908);
and U13231 (N_13231,N_11913,N_11305);
nor U13232 (N_13232,N_11427,N_11892);
or U13233 (N_13233,N_10753,N_11559);
and U13234 (N_13234,N_11806,N_10645);
nand U13235 (N_13235,N_10679,N_11779);
xnor U13236 (N_13236,N_10917,N_10881);
and U13237 (N_13237,N_11220,N_10781);
and U13238 (N_13238,N_11834,N_11166);
and U13239 (N_13239,N_11839,N_10609);
or U13240 (N_13240,N_10903,N_10626);
and U13241 (N_13241,N_10658,N_10742);
nor U13242 (N_13242,N_10780,N_11981);
or U13243 (N_13243,N_11178,N_11431);
and U13244 (N_13244,N_10915,N_11997);
xor U13245 (N_13245,N_11372,N_11076);
nand U13246 (N_13246,N_11219,N_11313);
and U13247 (N_13247,N_10690,N_11658);
and U13248 (N_13248,N_11061,N_10652);
nand U13249 (N_13249,N_11288,N_11137);
nor U13250 (N_13250,N_11410,N_10671);
nand U13251 (N_13251,N_11061,N_10562);
nand U13252 (N_13252,N_11623,N_11054);
or U13253 (N_13253,N_11781,N_11928);
or U13254 (N_13254,N_11435,N_11012);
and U13255 (N_13255,N_11757,N_11135);
nand U13256 (N_13256,N_11179,N_11272);
nor U13257 (N_13257,N_11491,N_11541);
nand U13258 (N_13258,N_11638,N_11567);
nand U13259 (N_13259,N_11834,N_11601);
nor U13260 (N_13260,N_11254,N_11550);
nor U13261 (N_13261,N_10629,N_10838);
nand U13262 (N_13262,N_11430,N_10753);
and U13263 (N_13263,N_11517,N_11762);
nand U13264 (N_13264,N_11877,N_11470);
nor U13265 (N_13265,N_11530,N_11198);
xnor U13266 (N_13266,N_11327,N_11976);
nor U13267 (N_13267,N_11651,N_11785);
and U13268 (N_13268,N_11178,N_11848);
nor U13269 (N_13269,N_11282,N_11642);
nand U13270 (N_13270,N_10742,N_11546);
or U13271 (N_13271,N_10953,N_10588);
and U13272 (N_13272,N_11171,N_11741);
nand U13273 (N_13273,N_11466,N_11595);
nor U13274 (N_13274,N_11696,N_11963);
nand U13275 (N_13275,N_11823,N_11934);
xnor U13276 (N_13276,N_10978,N_10874);
xor U13277 (N_13277,N_11085,N_10684);
nand U13278 (N_13278,N_11156,N_11091);
and U13279 (N_13279,N_10568,N_10745);
and U13280 (N_13280,N_10593,N_11620);
and U13281 (N_13281,N_11040,N_11618);
and U13282 (N_13282,N_11199,N_11648);
xor U13283 (N_13283,N_11499,N_10660);
nand U13284 (N_13284,N_11821,N_10776);
nand U13285 (N_13285,N_11613,N_10729);
nand U13286 (N_13286,N_11756,N_10712);
nor U13287 (N_13287,N_11565,N_11796);
nand U13288 (N_13288,N_11655,N_10587);
xor U13289 (N_13289,N_10618,N_11712);
or U13290 (N_13290,N_11883,N_10864);
and U13291 (N_13291,N_11679,N_10772);
xnor U13292 (N_13292,N_11626,N_11391);
nand U13293 (N_13293,N_11116,N_10892);
or U13294 (N_13294,N_11217,N_11126);
nor U13295 (N_13295,N_11542,N_10885);
nand U13296 (N_13296,N_11706,N_11258);
xnor U13297 (N_13297,N_10539,N_11162);
nor U13298 (N_13298,N_10861,N_11924);
and U13299 (N_13299,N_10699,N_11601);
and U13300 (N_13300,N_10776,N_11556);
and U13301 (N_13301,N_10799,N_11632);
or U13302 (N_13302,N_11349,N_10844);
nand U13303 (N_13303,N_10629,N_11668);
xnor U13304 (N_13304,N_11111,N_11030);
nor U13305 (N_13305,N_11934,N_11939);
nor U13306 (N_13306,N_11159,N_11112);
nand U13307 (N_13307,N_11934,N_10688);
and U13308 (N_13308,N_11049,N_10906);
nor U13309 (N_13309,N_10675,N_11090);
or U13310 (N_13310,N_11934,N_11917);
and U13311 (N_13311,N_10672,N_10926);
nor U13312 (N_13312,N_10571,N_11358);
nand U13313 (N_13313,N_11978,N_10552);
nand U13314 (N_13314,N_10734,N_11944);
or U13315 (N_13315,N_11699,N_11775);
or U13316 (N_13316,N_10989,N_10521);
and U13317 (N_13317,N_10617,N_11156);
and U13318 (N_13318,N_11183,N_10820);
and U13319 (N_13319,N_10779,N_10860);
nand U13320 (N_13320,N_11278,N_10644);
xor U13321 (N_13321,N_11630,N_10956);
nor U13322 (N_13322,N_11415,N_11895);
nand U13323 (N_13323,N_10796,N_10965);
nand U13324 (N_13324,N_11079,N_11678);
and U13325 (N_13325,N_11427,N_10978);
nor U13326 (N_13326,N_11056,N_11910);
xnor U13327 (N_13327,N_11676,N_10959);
xnor U13328 (N_13328,N_11330,N_11128);
or U13329 (N_13329,N_11884,N_10781);
or U13330 (N_13330,N_10733,N_11660);
nor U13331 (N_13331,N_11334,N_11979);
or U13332 (N_13332,N_10625,N_11395);
or U13333 (N_13333,N_11247,N_10561);
nand U13334 (N_13334,N_11300,N_10926);
nand U13335 (N_13335,N_10934,N_11213);
nor U13336 (N_13336,N_10896,N_11464);
nor U13337 (N_13337,N_11021,N_10665);
or U13338 (N_13338,N_10963,N_11607);
or U13339 (N_13339,N_10881,N_11646);
and U13340 (N_13340,N_11390,N_11290);
nand U13341 (N_13341,N_10939,N_11964);
nor U13342 (N_13342,N_10945,N_10965);
or U13343 (N_13343,N_11202,N_11660);
nand U13344 (N_13344,N_11371,N_11464);
and U13345 (N_13345,N_10534,N_11620);
or U13346 (N_13346,N_10593,N_11933);
and U13347 (N_13347,N_11034,N_11103);
and U13348 (N_13348,N_11857,N_10583);
nor U13349 (N_13349,N_10912,N_10993);
nor U13350 (N_13350,N_11735,N_11175);
or U13351 (N_13351,N_11295,N_11959);
or U13352 (N_13352,N_10923,N_11457);
nand U13353 (N_13353,N_11224,N_10524);
nor U13354 (N_13354,N_10636,N_10797);
nor U13355 (N_13355,N_10749,N_11478);
and U13356 (N_13356,N_11227,N_11823);
nor U13357 (N_13357,N_11937,N_11414);
nand U13358 (N_13358,N_11850,N_10587);
or U13359 (N_13359,N_11762,N_10997);
nor U13360 (N_13360,N_11908,N_11448);
nand U13361 (N_13361,N_11355,N_11969);
xor U13362 (N_13362,N_10762,N_10997);
and U13363 (N_13363,N_11529,N_10762);
and U13364 (N_13364,N_11109,N_10692);
and U13365 (N_13365,N_11356,N_10602);
nand U13366 (N_13366,N_11549,N_11164);
nor U13367 (N_13367,N_10732,N_11421);
xor U13368 (N_13368,N_11254,N_11211);
nor U13369 (N_13369,N_10763,N_11788);
nor U13370 (N_13370,N_10949,N_11167);
or U13371 (N_13371,N_11260,N_11349);
or U13372 (N_13372,N_11035,N_10964);
nand U13373 (N_13373,N_11781,N_10973);
and U13374 (N_13374,N_11082,N_11720);
nand U13375 (N_13375,N_10873,N_10918);
or U13376 (N_13376,N_11718,N_11246);
and U13377 (N_13377,N_11358,N_10865);
nand U13378 (N_13378,N_10724,N_11770);
or U13379 (N_13379,N_10656,N_11558);
or U13380 (N_13380,N_11897,N_11144);
nor U13381 (N_13381,N_11693,N_11483);
and U13382 (N_13382,N_11557,N_11304);
nand U13383 (N_13383,N_10662,N_10781);
nor U13384 (N_13384,N_11676,N_10516);
nand U13385 (N_13385,N_11253,N_11011);
or U13386 (N_13386,N_11913,N_11984);
nand U13387 (N_13387,N_10872,N_11164);
and U13388 (N_13388,N_10941,N_11657);
nor U13389 (N_13389,N_11293,N_10830);
xor U13390 (N_13390,N_10542,N_11588);
and U13391 (N_13391,N_10846,N_10602);
or U13392 (N_13392,N_11915,N_11486);
nand U13393 (N_13393,N_10678,N_11808);
nand U13394 (N_13394,N_11987,N_11197);
nand U13395 (N_13395,N_11549,N_10859);
nand U13396 (N_13396,N_10516,N_10872);
nand U13397 (N_13397,N_10923,N_10805);
nand U13398 (N_13398,N_11620,N_10848);
nor U13399 (N_13399,N_11186,N_11366);
nor U13400 (N_13400,N_10790,N_11995);
nand U13401 (N_13401,N_10787,N_11655);
or U13402 (N_13402,N_11578,N_11311);
or U13403 (N_13403,N_11118,N_11518);
nand U13404 (N_13404,N_11356,N_10507);
nor U13405 (N_13405,N_11127,N_11970);
nor U13406 (N_13406,N_11674,N_11252);
or U13407 (N_13407,N_10718,N_11270);
and U13408 (N_13408,N_11176,N_11516);
and U13409 (N_13409,N_11405,N_11610);
and U13410 (N_13410,N_10927,N_10518);
nor U13411 (N_13411,N_10865,N_10695);
nor U13412 (N_13412,N_11702,N_10884);
or U13413 (N_13413,N_11955,N_10734);
xnor U13414 (N_13414,N_10650,N_11513);
and U13415 (N_13415,N_10586,N_11730);
or U13416 (N_13416,N_11044,N_11317);
or U13417 (N_13417,N_11588,N_10508);
nor U13418 (N_13418,N_11500,N_11996);
nor U13419 (N_13419,N_11738,N_11394);
nor U13420 (N_13420,N_11122,N_11804);
nor U13421 (N_13421,N_10956,N_11212);
or U13422 (N_13422,N_11187,N_10941);
or U13423 (N_13423,N_10808,N_10646);
xor U13424 (N_13424,N_11310,N_10961);
nor U13425 (N_13425,N_10981,N_11134);
xnor U13426 (N_13426,N_11863,N_11764);
and U13427 (N_13427,N_10915,N_11690);
and U13428 (N_13428,N_10969,N_11048);
xnor U13429 (N_13429,N_10579,N_11410);
nand U13430 (N_13430,N_10862,N_11030);
or U13431 (N_13431,N_11282,N_11611);
or U13432 (N_13432,N_10772,N_11981);
nand U13433 (N_13433,N_10627,N_10885);
and U13434 (N_13434,N_11958,N_11287);
nor U13435 (N_13435,N_10801,N_11917);
xor U13436 (N_13436,N_10501,N_11272);
nor U13437 (N_13437,N_10742,N_11116);
and U13438 (N_13438,N_11507,N_11260);
nor U13439 (N_13439,N_11388,N_11340);
and U13440 (N_13440,N_10767,N_11117);
nand U13441 (N_13441,N_11861,N_10598);
or U13442 (N_13442,N_11478,N_10608);
or U13443 (N_13443,N_10985,N_11452);
nand U13444 (N_13444,N_11053,N_10648);
xnor U13445 (N_13445,N_10887,N_11122);
nor U13446 (N_13446,N_11030,N_10647);
or U13447 (N_13447,N_11206,N_11487);
and U13448 (N_13448,N_11479,N_11417);
and U13449 (N_13449,N_11858,N_10539);
xnor U13450 (N_13450,N_11335,N_10615);
or U13451 (N_13451,N_11387,N_11930);
or U13452 (N_13452,N_11045,N_11118);
nand U13453 (N_13453,N_10866,N_11283);
or U13454 (N_13454,N_11318,N_10643);
nor U13455 (N_13455,N_10622,N_11793);
and U13456 (N_13456,N_10891,N_10802);
nand U13457 (N_13457,N_11102,N_10501);
or U13458 (N_13458,N_11995,N_10506);
nand U13459 (N_13459,N_10920,N_10876);
xor U13460 (N_13460,N_11487,N_10696);
nor U13461 (N_13461,N_10703,N_10904);
nand U13462 (N_13462,N_11187,N_10572);
or U13463 (N_13463,N_10777,N_11908);
nand U13464 (N_13464,N_11591,N_11029);
or U13465 (N_13465,N_11661,N_10947);
or U13466 (N_13466,N_11249,N_11454);
xnor U13467 (N_13467,N_11563,N_11727);
nor U13468 (N_13468,N_11083,N_10541);
nand U13469 (N_13469,N_11290,N_11158);
or U13470 (N_13470,N_10581,N_11485);
nand U13471 (N_13471,N_11383,N_11348);
or U13472 (N_13472,N_10851,N_11197);
xnor U13473 (N_13473,N_10519,N_11012);
nor U13474 (N_13474,N_11016,N_11233);
nand U13475 (N_13475,N_11378,N_11937);
and U13476 (N_13476,N_11188,N_11984);
xnor U13477 (N_13477,N_11247,N_11632);
and U13478 (N_13478,N_11455,N_11078);
xor U13479 (N_13479,N_11791,N_11545);
or U13480 (N_13480,N_11110,N_11193);
and U13481 (N_13481,N_11509,N_11848);
xor U13482 (N_13482,N_11828,N_11380);
nor U13483 (N_13483,N_11591,N_11330);
nand U13484 (N_13484,N_11235,N_11166);
nand U13485 (N_13485,N_11030,N_11798);
nand U13486 (N_13486,N_11016,N_10783);
nand U13487 (N_13487,N_11510,N_11005);
nor U13488 (N_13488,N_10942,N_11925);
nand U13489 (N_13489,N_11682,N_10769);
xor U13490 (N_13490,N_10926,N_11385);
xor U13491 (N_13491,N_11394,N_11783);
nor U13492 (N_13492,N_11384,N_10695);
nand U13493 (N_13493,N_10892,N_11110);
nor U13494 (N_13494,N_11572,N_11999);
xor U13495 (N_13495,N_11286,N_10773);
nand U13496 (N_13496,N_11587,N_11184);
nor U13497 (N_13497,N_10984,N_10712);
nor U13498 (N_13498,N_10696,N_11612);
or U13499 (N_13499,N_11917,N_11347);
or U13500 (N_13500,N_12398,N_12446);
nor U13501 (N_13501,N_13434,N_13076);
nand U13502 (N_13502,N_12751,N_13131);
nand U13503 (N_13503,N_12329,N_12132);
nor U13504 (N_13504,N_12306,N_12339);
xnor U13505 (N_13505,N_12813,N_12419);
xor U13506 (N_13506,N_13466,N_12817);
or U13507 (N_13507,N_12886,N_13493);
nor U13508 (N_13508,N_13471,N_12209);
and U13509 (N_13509,N_12349,N_12006);
and U13510 (N_13510,N_12159,N_12040);
nand U13511 (N_13511,N_12050,N_12982);
or U13512 (N_13512,N_12195,N_12334);
or U13513 (N_13513,N_12758,N_13109);
nor U13514 (N_13514,N_12024,N_12205);
or U13515 (N_13515,N_13314,N_12400);
nor U13516 (N_13516,N_12241,N_12512);
or U13517 (N_13517,N_12760,N_13064);
xor U13518 (N_13518,N_13407,N_13244);
and U13519 (N_13519,N_12181,N_13368);
and U13520 (N_13520,N_12738,N_12971);
and U13521 (N_13521,N_12098,N_12722);
or U13522 (N_13522,N_13106,N_12719);
and U13523 (N_13523,N_12773,N_12675);
and U13524 (N_13524,N_12154,N_12327);
or U13525 (N_13525,N_12853,N_12338);
nor U13526 (N_13526,N_12402,N_12492);
nor U13527 (N_13527,N_12005,N_13336);
nand U13528 (N_13528,N_13092,N_13155);
nor U13529 (N_13529,N_12753,N_13499);
nor U13530 (N_13530,N_12156,N_12915);
and U13531 (N_13531,N_12654,N_12038);
or U13532 (N_13532,N_12126,N_13192);
and U13533 (N_13533,N_12717,N_12097);
nand U13534 (N_13534,N_12810,N_12534);
and U13535 (N_13535,N_12876,N_12567);
and U13536 (N_13536,N_12527,N_13234);
and U13537 (N_13537,N_13325,N_12657);
or U13538 (N_13538,N_13366,N_12806);
xnor U13539 (N_13539,N_12069,N_12684);
nand U13540 (N_13540,N_12546,N_13068);
nor U13541 (N_13541,N_12574,N_12163);
and U13542 (N_13542,N_12433,N_12291);
nor U13543 (N_13543,N_13157,N_12371);
nor U13544 (N_13544,N_12083,N_12037);
nor U13545 (N_13545,N_13341,N_12228);
or U13546 (N_13546,N_13150,N_12002);
or U13547 (N_13547,N_12749,N_12352);
or U13548 (N_13548,N_13171,N_13271);
nand U13549 (N_13549,N_12214,N_12447);
or U13550 (N_13550,N_13470,N_13290);
nand U13551 (N_13551,N_12885,N_12413);
or U13552 (N_13552,N_13289,N_12443);
and U13553 (N_13553,N_13405,N_12514);
nand U13554 (N_13554,N_12939,N_13468);
and U13555 (N_13555,N_12252,N_13227);
nand U13556 (N_13556,N_12138,N_13221);
nand U13557 (N_13557,N_12149,N_13229);
nor U13558 (N_13558,N_12115,N_12369);
and U13559 (N_13559,N_12171,N_12118);
nor U13560 (N_13560,N_13112,N_13382);
or U13561 (N_13561,N_12128,N_12392);
or U13562 (N_13562,N_12755,N_12548);
nand U13563 (N_13563,N_12878,N_12862);
or U13564 (N_13564,N_12586,N_12643);
nand U13565 (N_13565,N_12461,N_12950);
or U13566 (N_13566,N_12135,N_12121);
nor U13567 (N_13567,N_13156,N_12966);
nand U13568 (N_13568,N_12350,N_12899);
nand U13569 (N_13569,N_12998,N_13272);
and U13570 (N_13570,N_12144,N_12609);
nor U13571 (N_13571,N_12639,N_12331);
or U13572 (N_13572,N_12343,N_12091);
xor U13573 (N_13573,N_13057,N_12078);
nand U13574 (N_13574,N_12636,N_12829);
and U13575 (N_13575,N_13189,N_12445);
or U13576 (N_13576,N_12290,N_12234);
xnor U13577 (N_13577,N_12564,N_12616);
and U13578 (N_13578,N_13310,N_13484);
or U13579 (N_13579,N_12945,N_12785);
and U13580 (N_13580,N_13404,N_12438);
xor U13581 (N_13581,N_13100,N_12698);
nor U13582 (N_13582,N_12559,N_13352);
xor U13583 (N_13583,N_12152,N_12624);
and U13584 (N_13584,N_12737,N_12417);
or U13585 (N_13585,N_13082,N_13108);
nor U13586 (N_13586,N_13004,N_12669);
nor U13587 (N_13587,N_12423,N_12047);
nand U13588 (N_13588,N_12380,N_13160);
and U13589 (N_13589,N_12049,N_12203);
nor U13590 (N_13590,N_12463,N_12911);
nand U13591 (N_13591,N_12418,N_12670);
xor U13592 (N_13592,N_12487,N_12439);
nor U13593 (N_13593,N_12300,N_13135);
nor U13594 (N_13594,N_13001,N_12520);
nor U13595 (N_13595,N_12803,N_13482);
nor U13596 (N_13596,N_13232,N_13473);
and U13597 (N_13597,N_13374,N_13426);
and U13598 (N_13598,N_12092,N_12648);
nor U13599 (N_13599,N_12781,N_13396);
and U13600 (N_13600,N_13365,N_12298);
and U13601 (N_13601,N_12724,N_12431);
and U13602 (N_13602,N_12099,N_12772);
nor U13603 (N_13603,N_13213,N_13452);
and U13604 (N_13604,N_12765,N_12304);
or U13605 (N_13605,N_13093,N_12686);
nor U13606 (N_13606,N_12688,N_12907);
xor U13607 (N_13607,N_12364,N_13191);
nand U13608 (N_13608,N_12776,N_12133);
and U13609 (N_13609,N_13320,N_12299);
or U13610 (N_13610,N_12844,N_12778);
nand U13611 (N_13611,N_12951,N_12936);
or U13612 (N_13612,N_12057,N_12690);
nor U13613 (N_13613,N_13427,N_12732);
nand U13614 (N_13614,N_12042,N_13007);
nor U13615 (N_13615,N_12986,N_12385);
xor U13616 (N_13616,N_12134,N_12613);
and U13617 (N_13617,N_12708,N_12615);
xnor U13618 (N_13618,N_12764,N_12190);
and U13619 (N_13619,N_12028,N_12265);
and U13620 (N_13620,N_13309,N_12797);
and U13621 (N_13621,N_12821,N_13152);
nand U13622 (N_13622,N_13167,N_12762);
nor U13623 (N_13623,N_12476,N_12943);
or U13624 (N_13624,N_12058,N_12632);
nor U13625 (N_13625,N_13023,N_12411);
nand U13626 (N_13626,N_12425,N_13377);
nor U13627 (N_13627,N_12905,N_13246);
nand U13628 (N_13628,N_12630,N_12856);
nand U13629 (N_13629,N_12235,N_13299);
nor U13630 (N_13630,N_12137,N_13169);
nor U13631 (N_13631,N_13292,N_12116);
nand U13632 (N_13632,N_12009,N_12680);
or U13633 (N_13633,N_13260,N_12901);
or U13634 (N_13634,N_12931,N_12977);
or U13635 (N_13635,N_12569,N_12964);
nand U13636 (N_13636,N_12896,N_12969);
nand U13637 (N_13637,N_13173,N_13187);
xnor U13638 (N_13638,N_12441,N_12714);
nor U13639 (N_13639,N_12279,N_12695);
nor U13640 (N_13640,N_13347,N_12308);
or U13641 (N_13641,N_12902,N_12168);
nand U13642 (N_13642,N_12830,N_12017);
nor U13643 (N_13643,N_12712,N_12633);
and U13644 (N_13644,N_13081,N_12250);
and U13645 (N_13645,N_13371,N_12281);
nor U13646 (N_13646,N_13038,N_12489);
or U13647 (N_13647,N_12594,N_12314);
and U13648 (N_13648,N_13099,N_13370);
nand U13649 (N_13649,N_12259,N_12027);
and U13650 (N_13650,N_13275,N_12916);
or U13651 (N_13651,N_13383,N_12972);
or U13652 (N_13652,N_12059,N_12917);
or U13653 (N_13653,N_12555,N_13021);
nor U13654 (N_13654,N_12434,N_12479);
or U13655 (N_13655,N_12472,N_12549);
xnor U13656 (N_13656,N_12868,N_13075);
nand U13657 (N_13657,N_12909,N_12715);
nand U13658 (N_13658,N_13350,N_12179);
nand U13659 (N_13659,N_12847,N_13199);
nor U13660 (N_13660,N_12544,N_13040);
nand U13661 (N_13661,N_13206,N_12061);
and U13662 (N_13662,N_12394,N_13019);
nor U13663 (N_13663,N_13318,N_12748);
and U13664 (N_13664,N_12540,N_12136);
nor U13665 (N_13665,N_12401,N_13334);
nor U13666 (N_13666,N_12730,N_12227);
or U13667 (N_13667,N_12991,N_12946);
nor U13668 (N_13668,N_12296,N_12677);
and U13669 (N_13669,N_13186,N_12303);
nand U13670 (N_13670,N_12612,N_12273);
nand U13671 (N_13671,N_12344,N_12824);
nor U13672 (N_13672,N_13486,N_12914);
nand U13673 (N_13673,N_13414,N_12302);
nand U13674 (N_13674,N_12311,N_12442);
nor U13675 (N_13675,N_13089,N_12562);
nand U13676 (N_13676,N_12860,N_12882);
and U13677 (N_13677,N_13280,N_13175);
nor U13678 (N_13678,N_12767,N_12183);
or U13679 (N_13679,N_12893,N_13312);
nor U13680 (N_13680,N_12837,N_13451);
and U13681 (N_13681,N_12805,N_12543);
nor U13682 (N_13682,N_12890,N_13011);
nor U13683 (N_13683,N_12211,N_13284);
nor U13684 (N_13684,N_12981,N_12359);
nor U13685 (N_13685,N_12952,N_13137);
nand U13686 (N_13686,N_12427,N_12828);
nor U13687 (N_13687,N_12275,N_12033);
nor U13688 (N_13688,N_13480,N_13070);
xor U13689 (N_13689,N_12561,N_12967);
nand U13690 (N_13690,N_12108,N_12879);
nand U13691 (N_13691,N_12827,N_13225);
or U13692 (N_13692,N_13307,N_12404);
xor U13693 (N_13693,N_12668,N_12146);
nor U13694 (N_13694,N_12535,N_12023);
nand U13695 (N_13695,N_12464,N_12382);
or U13696 (N_13696,N_13119,N_12774);
nand U13697 (N_13697,N_12623,N_12627);
nor U13698 (N_13698,N_13145,N_12603);
nor U13699 (N_13699,N_13020,N_12840);
nor U13700 (N_13700,N_13197,N_12052);
nand U13701 (N_13701,N_12683,N_12576);
or U13702 (N_13702,N_13339,N_12855);
and U13703 (N_13703,N_12449,N_12277);
nor U13704 (N_13704,N_12956,N_13429);
or U13705 (N_13705,N_12904,N_12485);
nor U13706 (N_13706,N_12645,N_13185);
xor U13707 (N_13707,N_12598,N_12510);
nand U13708 (N_13708,N_13250,N_12538);
nand U13709 (N_13709,N_12375,N_13375);
nand U13710 (N_13710,N_12409,N_12237);
nand U13711 (N_13711,N_12036,N_12416);
and U13712 (N_13712,N_12619,N_12330);
or U13713 (N_13713,N_12784,N_12383);
nor U13714 (N_13714,N_12110,N_12187);
xnor U13715 (N_13715,N_13154,N_13008);
nand U13716 (N_13716,N_12516,N_13378);
xnor U13717 (N_13717,N_12366,N_12353);
xnor U13718 (N_13718,N_12429,N_12617);
and U13719 (N_13719,N_12949,N_13442);
nand U13720 (N_13720,N_12701,N_12872);
or U13721 (N_13721,N_13379,N_12611);
nand U13722 (N_13722,N_13143,N_12333);
or U13723 (N_13723,N_12457,N_12955);
and U13724 (N_13724,N_13133,N_12924);
nand U13725 (N_13725,N_12505,N_12247);
nand U13726 (N_13726,N_13445,N_12269);
nor U13727 (N_13727,N_12158,N_12161);
or U13728 (N_13728,N_13005,N_12039);
and U13729 (N_13729,N_12859,N_13031);
xor U13730 (N_13730,N_12864,N_12260);
nor U13731 (N_13731,N_12808,N_13287);
nor U13732 (N_13732,N_12226,N_12809);
and U13733 (N_13733,N_12105,N_12846);
or U13734 (N_13734,N_12599,N_12565);
and U13735 (N_13735,N_12518,N_13303);
or U13736 (N_13736,N_13243,N_13411);
or U13737 (N_13737,N_12189,N_12528);
and U13738 (N_13738,N_12990,N_12096);
or U13739 (N_13739,N_13002,N_12139);
or U13740 (N_13740,N_13104,N_13276);
nor U13741 (N_13741,N_13277,N_13316);
nor U13742 (N_13742,N_12318,N_12248);
nor U13743 (N_13743,N_12356,N_13358);
or U13744 (N_13744,N_12880,N_12881);
and U13745 (N_13745,N_13326,N_12367);
nand U13746 (N_13746,N_13389,N_12022);
or U13747 (N_13747,N_12948,N_12975);
nor U13748 (N_13748,N_12974,N_12388);
or U13749 (N_13749,N_13422,N_13181);
nor U13750 (N_13750,N_12581,N_13380);
nand U13751 (N_13751,N_13144,N_13097);
nor U13752 (N_13752,N_12210,N_13297);
and U13753 (N_13753,N_12324,N_12093);
nand U13754 (N_13754,N_12166,N_12725);
or U13755 (N_13755,N_13338,N_12693);
and U13756 (N_13756,N_12676,N_12869);
nand U13757 (N_13757,N_12086,N_13009);
or U13758 (N_13758,N_13444,N_13054);
nor U13759 (N_13759,N_12585,N_12664);
or U13760 (N_13760,N_12511,N_12095);
nor U13761 (N_13761,N_13322,N_12362);
nand U13762 (N_13762,N_12845,N_12276);
nand U13763 (N_13763,N_12957,N_12889);
or U13764 (N_13764,N_13488,N_13130);
and U13765 (N_13765,N_13490,N_12048);
xnor U13766 (N_13766,N_12777,N_13311);
nor U13767 (N_13767,N_12120,N_12665);
or U13768 (N_13768,N_13215,N_12592);
nand U13769 (N_13769,N_12779,N_12376);
nand U13770 (N_13770,N_12787,N_13291);
or U13771 (N_13771,N_12460,N_13198);
nor U13772 (N_13772,N_13025,N_12874);
and U13773 (N_13773,N_12642,N_12321);
and U13774 (N_13774,N_12628,N_12794);
nor U13775 (N_13775,N_12703,N_13072);
nor U13776 (N_13776,N_12264,N_12201);
and U13777 (N_13777,N_13432,N_12621);
nor U13778 (N_13778,N_13469,N_12666);
nor U13779 (N_13779,N_12386,N_13464);
or U13780 (N_13780,N_12697,N_13263);
xor U13781 (N_13781,N_12151,N_12992);
nor U13782 (N_13782,N_12673,N_13298);
nor U13783 (N_13783,N_13050,N_12075);
nand U13784 (N_13784,N_12918,N_13035);
nor U13785 (N_13785,N_12572,N_13285);
or U13786 (N_13786,N_12537,N_13059);
nor U13787 (N_13787,N_13373,N_12900);
or U13788 (N_13788,N_12947,N_12925);
nand U13789 (N_13789,N_13301,N_12733);
or U13790 (N_13790,N_12125,N_12531);
nor U13791 (N_13791,N_12430,N_13400);
and U13792 (N_13792,N_13385,N_12953);
and U13793 (N_13793,N_13107,N_12727);
and U13794 (N_13794,N_12456,N_13086);
nor U13795 (N_13795,N_12157,N_13308);
nor U13796 (N_13796,N_12906,N_13136);
nor U13797 (N_13797,N_12176,N_12710);
and U13798 (N_13798,N_13182,N_12743);
and U13799 (N_13799,N_12626,N_12173);
nand U13800 (N_13800,N_12452,N_13321);
xnor U13801 (N_13801,N_12458,N_12508);
and U13802 (N_13802,N_12802,N_13448);
and U13803 (N_13803,N_12354,N_12658);
and U13804 (N_13804,N_12851,N_12519);
and U13805 (N_13805,N_12188,N_12494);
or U13806 (N_13806,N_13302,N_12542);
or U13807 (N_13807,N_12620,N_12937);
and U13808 (N_13808,N_13264,N_12556);
and U13809 (N_13809,N_12003,N_12007);
or U13810 (N_13810,N_12858,N_12721);
and U13811 (N_13811,N_12647,N_12313);
nor U13812 (N_13812,N_13265,N_13034);
nor U13813 (N_13813,N_12614,N_12903);
nand U13814 (N_13814,N_13036,N_13248);
or U13815 (N_13815,N_12877,N_12987);
xor U13816 (N_13816,N_13024,N_13257);
or U13817 (N_13817,N_13300,N_12122);
and U13818 (N_13818,N_13037,N_12496);
nand U13819 (N_13819,N_12068,N_13395);
and U13820 (N_13820,N_12888,N_12601);
and U13821 (N_13821,N_12497,N_12606);
or U13822 (N_13822,N_13372,N_12517);
nand U13823 (N_13823,N_13105,N_12471);
or U13824 (N_13824,N_12795,N_12174);
nor U13825 (N_13825,N_12034,N_12836);
or U13826 (N_13826,N_12346,N_12021);
nand U13827 (N_13827,N_13356,N_13134);
xor U13828 (N_13828,N_12713,N_12412);
or U13829 (N_13829,N_13386,N_13039);
nor U13830 (N_13830,N_12001,N_12408);
nand U13831 (N_13831,N_12570,N_12268);
nand U13832 (N_13832,N_12213,N_13164);
or U13833 (N_13833,N_12825,N_13481);
or U13834 (N_13834,N_12477,N_12397);
and U13835 (N_13835,N_12414,N_12728);
nand U13836 (N_13836,N_12744,N_12578);
nand U13837 (N_13837,N_13278,N_12072);
or U13838 (N_13838,N_12745,N_12088);
nor U13839 (N_13839,N_12605,N_13345);
nand U13840 (N_13840,N_13273,N_12652);
xor U13841 (N_13841,N_12832,N_13124);
or U13842 (N_13842,N_13438,N_12278);
nor U13843 (N_13843,N_13195,N_13419);
nand U13844 (N_13844,N_12965,N_13362);
and U13845 (N_13845,N_13237,N_12500);
and U13846 (N_13846,N_12271,N_12124);
and U13847 (N_13847,N_13162,N_12563);
or U13848 (N_13848,N_12554,N_13492);
nor U13849 (N_13849,N_12687,N_12493);
nand U13850 (N_13850,N_12220,N_12410);
and U13851 (N_13851,N_13259,N_13161);
nor U13852 (N_13852,N_12667,N_13000);
or U13853 (N_13853,N_12790,N_12257);
and U13854 (N_13854,N_12453,N_12080);
and U13855 (N_13855,N_13165,N_13006);
and U13856 (N_13856,N_12373,N_12345);
or U13857 (N_13857,N_12251,N_12884);
or U13858 (N_13858,N_12897,N_13026);
and U13859 (N_13859,N_12579,N_12782);
nor U13860 (N_13860,N_13067,N_12481);
and U13861 (N_13861,N_12085,N_13330);
or U13862 (N_13862,N_13283,N_13251);
or U13863 (N_13863,N_13217,N_13125);
or U13864 (N_13864,N_12326,N_12358);
nand U13865 (N_13865,N_13017,N_13032);
or U13866 (N_13866,N_12557,N_13483);
nor U13867 (N_13867,N_12524,N_13418);
and U13868 (N_13868,N_12076,N_13016);
nand U13869 (N_13869,N_13381,N_13044);
or U13870 (N_13870,N_13194,N_12301);
and U13871 (N_13871,N_12348,N_12186);
nor U13872 (N_13872,N_12140,N_12622);
nor U13873 (N_13873,N_12656,N_12145);
and U13874 (N_13874,N_12478,N_12335);
nor U13875 (N_13875,N_12734,N_13354);
or U13876 (N_13876,N_13399,N_12959);
or U13877 (N_13877,N_12451,N_12062);
nor U13878 (N_13878,N_12067,N_12499);
nor U13879 (N_13879,N_12046,N_12768);
nor U13880 (N_13880,N_13090,N_13048);
xor U13881 (N_13881,N_12978,N_13474);
nand U13882 (N_13882,N_12854,N_13061);
nand U13883 (N_13883,N_13274,N_12484);
xnor U13884 (N_13884,N_13477,N_12102);
or U13885 (N_13885,N_13228,N_12106);
and U13886 (N_13886,N_12054,N_12420);
nand U13887 (N_13887,N_12740,N_13113);
and U13888 (N_13888,N_12769,N_12663);
and U13889 (N_13889,N_12930,N_12466);
nor U13890 (N_13890,N_13074,N_13266);
nand U13891 (N_13891,N_12629,N_12739);
nor U13892 (N_13892,N_12454,N_12292);
nand U13893 (N_13893,N_13176,N_12440);
xor U13894 (N_13894,N_12010,N_12267);
nand U13895 (N_13895,N_12162,N_12233);
and U13896 (N_13896,N_13436,N_12056);
nand U13897 (N_13897,N_12651,N_12736);
nand U13898 (N_13898,N_13317,N_12910);
and U13899 (N_13899,N_12705,N_12104);
and U13900 (N_13900,N_13077,N_12455);
or U13901 (N_13901,N_12217,N_12087);
or U13902 (N_13902,N_12533,N_13360);
nand U13903 (N_13903,N_13397,N_13027);
nor U13904 (N_13904,N_13126,N_13421);
or U13905 (N_13905,N_12539,N_12256);
xor U13906 (N_13906,N_12509,N_12243);
and U13907 (N_13907,N_12399,N_12871);
nor U13908 (N_13908,N_12170,N_12222);
or U13909 (N_13909,N_12525,N_12141);
nor U13910 (N_13910,N_12026,N_13073);
xor U13911 (N_13911,N_12839,N_12490);
xnor U13912 (N_13912,N_12403,N_12604);
and U13913 (N_13913,N_12444,N_12699);
or U13914 (N_13914,N_12225,N_12835);
or U13915 (N_13915,N_12655,N_12566);
or U13916 (N_13916,N_12602,N_13030);
and U13917 (N_13917,N_12506,N_13494);
and U13918 (N_13918,N_12595,N_13286);
nor U13919 (N_13919,N_13462,N_12053);
or U13920 (N_13920,N_13458,N_12702);
and U13921 (N_13921,N_13179,N_12031);
and U13922 (N_13922,N_12789,N_12898);
nor U13923 (N_13923,N_13028,N_13410);
xor U13924 (N_13924,N_12185,N_12320);
nor U13925 (N_13925,N_13241,N_12661);
nand U13926 (N_13926,N_13367,N_12094);
nand U13927 (N_13927,N_12130,N_12766);
nor U13928 (N_13928,N_12997,N_12070);
or U13929 (N_13929,N_13049,N_13329);
and U13930 (N_13930,N_12689,N_13069);
nand U13931 (N_13931,N_13249,N_12694);
nand U13932 (N_13932,N_12560,N_12283);
or U13933 (N_13933,N_12029,N_12771);
or U13934 (N_13934,N_12985,N_13342);
nand U13935 (N_13935,N_12200,N_13268);
and U13936 (N_13936,N_12522,N_13417);
and U13937 (N_13937,N_12498,N_13029);
nand U13938 (N_13938,N_12913,N_12221);
xnor U13939 (N_13939,N_12631,N_12448);
nand U13940 (N_13940,N_13485,N_12610);
or U13941 (N_13941,N_13128,N_12491);
nor U13942 (N_13942,N_13423,N_12600);
nor U13943 (N_13943,N_13224,N_13333);
or U13944 (N_13944,N_12618,N_12261);
and U13945 (N_13945,N_12012,N_12501);
or U13946 (N_13946,N_13063,N_13315);
nor U13947 (N_13947,N_13256,N_12363);
nand U13948 (N_13948,N_13351,N_12014);
and U13949 (N_13949,N_13364,N_13435);
or U13950 (N_13950,N_13079,N_12090);
nor U13951 (N_13951,N_13212,N_12393);
nand U13952 (N_13952,N_13201,N_13253);
xnor U13953 (N_13953,N_13491,N_12515);
nor U13954 (N_13954,N_12008,N_13340);
or U13955 (N_13955,N_12377,N_12912);
and U13956 (N_13956,N_12142,N_13214);
nor U13957 (N_13957,N_13071,N_12148);
or U13958 (N_13958,N_12337,N_13420);
or U13959 (N_13959,N_12079,N_13168);
nand U13960 (N_13960,N_12984,N_12081);
or U13961 (N_13961,N_13242,N_12826);
and U13962 (N_13962,N_13218,N_12816);
nand U13963 (N_13963,N_13196,N_12820);
xnor U13964 (N_13964,N_12553,N_12341);
or U13965 (N_13965,N_13455,N_12597);
nand U13966 (N_13966,N_13121,N_13042);
or U13967 (N_13967,N_12266,N_12309);
nor U13968 (N_13968,N_13363,N_12424);
nand U13969 (N_13969,N_12378,N_13337);
or U13970 (N_13970,N_13387,N_12584);
and U13971 (N_13971,N_12263,N_12800);
or U13972 (N_13972,N_12020,N_13190);
or U13973 (N_13973,N_12043,N_13202);
and U13974 (N_13974,N_13098,N_13088);
or U13975 (N_13975,N_12747,N_13022);
and U13976 (N_13976,N_13149,N_12297);
and U13977 (N_13977,N_12866,N_13409);
nand U13978 (N_13978,N_13127,N_12796);
and U13979 (N_13979,N_12641,N_12198);
or U13980 (N_13980,N_12970,N_12191);
or U13981 (N_13981,N_12812,N_12045);
nand U13982 (N_13982,N_13465,N_12999);
or U13983 (N_13983,N_12541,N_13430);
nor U13984 (N_13984,N_12892,N_12368);
and U13985 (N_13985,N_13454,N_13296);
nor U13986 (N_13986,N_12938,N_12993);
and U13987 (N_13987,N_12396,N_12123);
and U13988 (N_13988,N_12089,N_13166);
nand U13989 (N_13989,N_12224,N_12025);
nand U13990 (N_13990,N_13060,N_12819);
or U13991 (N_13991,N_13233,N_12696);
and U13992 (N_13992,N_12178,N_12004);
nor U13993 (N_13993,N_12254,N_12249);
nor U13994 (N_13994,N_12150,N_12390);
or U13995 (N_13995,N_12019,N_12934);
nor U13996 (N_13996,N_13343,N_12550);
nor U13997 (N_13997,N_13348,N_13123);
nor U13998 (N_13998,N_13269,N_12775);
xnor U13999 (N_13999,N_13231,N_12274);
or U14000 (N_14000,N_13406,N_12976);
nor U14001 (N_14001,N_12927,N_13174);
and U14002 (N_14002,N_12634,N_12317);
or U14003 (N_14003,N_13335,N_12996);
nand U14004 (N_14004,N_13055,N_13172);
or U14005 (N_14005,N_12763,N_12202);
nand U14006 (N_14006,N_13349,N_12968);
xnor U14007 (N_14007,N_12757,N_12580);
or U14008 (N_14008,N_12799,N_13437);
and U14009 (N_14009,N_12842,N_13180);
nand U14010 (N_14010,N_12588,N_12849);
nand U14011 (N_14011,N_12482,N_13209);
or U14012 (N_14012,N_12246,N_13208);
nor U14013 (N_14013,N_13267,N_13449);
nand U14014 (N_14014,N_13095,N_13101);
and U14015 (N_14015,N_12044,N_13046);
and U14016 (N_14016,N_12625,N_12172);
nand U14017 (N_14017,N_12823,N_12215);
nor U14018 (N_14018,N_12143,N_12218);
and U14019 (N_14019,N_12328,N_12340);
or U14020 (N_14020,N_12834,N_12182);
or U14021 (N_14021,N_13497,N_12644);
or U14022 (N_14022,N_13230,N_12838);
or U14023 (N_14023,N_12272,N_12223);
nor U14024 (N_14024,N_13140,N_12316);
nor U14025 (N_14025,N_12582,N_13496);
and U14026 (N_14026,N_13216,N_13255);
and U14027 (N_14027,N_12973,N_12325);
and U14028 (N_14028,N_12459,N_13110);
nor U14029 (N_14029,N_12865,N_12653);
nor U14030 (N_14030,N_12175,N_12294);
nand U14031 (N_14031,N_12681,N_13391);
or U14032 (N_14032,N_12707,N_13461);
or U14033 (N_14033,N_12770,N_12100);
nand U14034 (N_14034,N_12422,N_13401);
or U14035 (N_14035,N_12196,N_12155);
or U14036 (N_14036,N_13440,N_12608);
nor U14037 (N_14037,N_12635,N_13047);
or U14038 (N_14038,N_12288,N_12841);
nor U14039 (N_14039,N_13254,N_12861);
and U14040 (N_14040,N_12018,N_13319);
and U14041 (N_14041,N_12117,N_13412);
nand U14042 (N_14042,N_12843,N_12486);
nand U14043 (N_14043,N_12607,N_12521);
nor U14044 (N_14044,N_12691,N_12160);
or U14045 (N_14045,N_13361,N_12674);
or U14046 (N_14046,N_12646,N_13078);
nor U14047 (N_14047,N_12783,N_12750);
and U14048 (N_14048,N_12193,N_13327);
nor U14049 (N_14049,N_12426,N_13091);
nand U14050 (N_14050,N_13293,N_12536);
xnor U14051 (N_14051,N_12206,N_12746);
and U14052 (N_14052,N_12640,N_13239);
xor U14053 (N_14053,N_13495,N_12583);
or U14054 (N_14054,N_13084,N_12289);
or U14055 (N_14055,N_12127,N_12908);
and U14056 (N_14056,N_12245,N_12682);
and U14057 (N_14057,N_12462,N_12718);
nor U14058 (N_14058,N_13294,N_12262);
nand U14059 (N_14059,N_13012,N_12405);
or U14060 (N_14060,N_12811,N_13183);
or U14061 (N_14061,N_12231,N_12685);
or U14062 (N_14062,N_13117,N_13398);
or U14063 (N_14063,N_13238,N_13013);
or U14064 (N_14064,N_12015,N_12063);
xor U14065 (N_14065,N_13460,N_13433);
or U14066 (N_14066,N_12147,N_13355);
nor U14067 (N_14067,N_12756,N_12204);
nand U14068 (N_14068,N_12255,N_13394);
and U14069 (N_14069,N_13115,N_13376);
nand U14070 (N_14070,N_12387,N_12084);
and U14071 (N_14071,N_12207,N_12979);
xnor U14072 (N_14072,N_13258,N_12852);
nor U14073 (N_14073,N_13313,N_12285);
nand U14074 (N_14074,N_12468,N_13252);
and U14075 (N_14075,N_12786,N_12895);
nor U14076 (N_14076,N_12280,N_12286);
or U14077 (N_14077,N_13439,N_12435);
nor U14078 (N_14078,N_13132,N_13003);
or U14079 (N_14079,N_12103,N_12384);
nand U14080 (N_14080,N_13207,N_13261);
nor U14081 (N_14081,N_13058,N_12372);
and U14082 (N_14082,N_12818,N_13033);
or U14083 (N_14083,N_12637,N_12219);
and U14084 (N_14084,N_12270,N_12184);
nor U14085 (N_14085,N_12436,N_13148);
nor U14086 (N_14086,N_12729,N_12488);
nand U14087 (N_14087,N_13282,N_12229);
nor U14088 (N_14088,N_12551,N_12983);
and U14089 (N_14089,N_12980,N_12523);
xor U14090 (N_14090,N_12815,N_12391);
and U14091 (N_14091,N_13103,N_12863);
or U14092 (N_14092,N_12513,N_12545);
xnor U14093 (N_14093,N_12473,N_13118);
nand U14094 (N_14094,N_13384,N_13393);
and U14095 (N_14095,N_13014,N_13159);
or U14096 (N_14096,N_12962,N_13062);
and U14097 (N_14097,N_12558,N_12071);
or U14098 (N_14098,N_12593,N_13203);
or U14099 (N_14099,N_12920,N_13323);
nand U14100 (N_14100,N_12530,N_12470);
nand U14101 (N_14101,N_12679,N_12994);
and U14102 (N_14102,N_12735,N_13188);
nor U14103 (N_14103,N_12504,N_12469);
and U14104 (N_14104,N_13472,N_12942);
nor U14105 (N_14105,N_12989,N_12822);
nand U14106 (N_14106,N_12192,N_12180);
nand U14107 (N_14107,N_12671,N_12064);
nor U14108 (N_14108,N_13139,N_13487);
nand U14109 (N_14109,N_13369,N_12232);
xor U14110 (N_14110,N_12659,N_12253);
xnor U14111 (N_14111,N_12926,N_12590);
nand U14112 (N_14112,N_12319,N_12723);
and U14113 (N_14113,N_12164,N_13184);
nand U14114 (N_14114,N_12107,N_13447);
or U14115 (N_14115,N_13279,N_13147);
nand U14116 (N_14116,N_12672,N_12407);
and U14117 (N_14117,N_13177,N_13450);
and U14118 (N_14118,N_12041,N_12483);
nand U14119 (N_14119,N_13295,N_12575);
nor U14120 (N_14120,N_12432,N_13453);
xnor U14121 (N_14121,N_12857,N_12305);
nor U14122 (N_14122,N_12238,N_13328);
and U14123 (N_14123,N_13463,N_13270);
nor U14124 (N_14124,N_12921,N_12503);
xor U14125 (N_14125,N_12587,N_13220);
or U14126 (N_14126,N_12284,N_12379);
or U14127 (N_14127,N_12596,N_12894);
nand U14128 (N_14128,N_13102,N_13141);
xnor U14129 (N_14129,N_12741,N_13211);
nor U14130 (N_14130,N_13235,N_12944);
nor U14131 (N_14131,N_13151,N_13262);
nor U14132 (N_14132,N_13304,N_12197);
nand U14133 (N_14133,N_12165,N_13415);
nand U14134 (N_14134,N_13178,N_13153);
and U14135 (N_14135,N_12109,N_12131);
nor U14136 (N_14136,N_12011,N_12475);
nor U14137 (N_14137,N_13245,N_12804);
nand U14138 (N_14138,N_13353,N_12923);
and U14139 (N_14139,N_12315,N_13403);
and U14140 (N_14140,N_13456,N_12678);
or U14141 (N_14141,N_13114,N_12360);
and U14142 (N_14142,N_12940,N_12709);
or U14143 (N_14143,N_13122,N_12032);
or U14144 (N_14144,N_12055,N_12831);
nand U14145 (N_14145,N_12437,N_12467);
nand U14146 (N_14146,N_12589,N_12258);
nor U14147 (N_14147,N_12351,N_12502);
and U14148 (N_14148,N_12706,N_13476);
nand U14149 (N_14149,N_13305,N_12850);
and U14150 (N_14150,N_13425,N_13498);
or U14151 (N_14151,N_12212,N_13120);
and U14152 (N_14152,N_12060,N_12428);
nand U14153 (N_14153,N_12875,N_12711);
xor U14154 (N_14154,N_12111,N_12323);
xor U14155 (N_14155,N_12035,N_13163);
and U14156 (N_14156,N_13051,N_12073);
or U14157 (N_14157,N_12389,N_12230);
nor U14158 (N_14158,N_13288,N_12112);
nand U14159 (N_14159,N_12129,N_12244);
nor U14160 (N_14160,N_13478,N_12935);
and U14161 (N_14161,N_12919,N_12995);
or U14162 (N_14162,N_12077,N_12573);
nor U14163 (N_14163,N_12082,N_12169);
xnor U14164 (N_14164,N_13080,N_13094);
and U14165 (N_14165,N_13200,N_13129);
nand U14166 (N_14166,N_12650,N_12312);
nor U14167 (N_14167,N_12887,N_12941);
and U14168 (N_14168,N_12933,N_13489);
nand U14169 (N_14169,N_12421,N_12883);
or U14170 (N_14170,N_13443,N_12552);
nand U14171 (N_14171,N_13142,N_13015);
xor U14172 (N_14172,N_13459,N_12065);
nand U14173 (N_14173,N_12752,N_12293);
xor U14174 (N_14174,N_13158,N_13018);
xnor U14175 (N_14175,N_12336,N_12833);
and U14176 (N_14176,N_12792,N_12591);
nor U14177 (N_14177,N_13441,N_12415);
and U14178 (N_14178,N_12960,N_12495);
nand U14179 (N_14179,N_12307,N_12988);
nand U14180 (N_14180,N_12704,N_12236);
nor U14181 (N_14181,N_12731,N_12720);
nand U14182 (N_14182,N_12759,N_12074);
nand U14183 (N_14183,N_13053,N_12929);
xor U14184 (N_14184,N_13346,N_12807);
and U14185 (N_14185,N_13357,N_13413);
nand U14186 (N_14186,N_12242,N_13359);
nor U14187 (N_14187,N_12754,N_13045);
or U14188 (N_14188,N_12814,N_12638);
or U14189 (N_14189,N_12101,N_12532);
xnor U14190 (N_14190,N_12287,N_12780);
and U14191 (N_14191,N_12013,N_13116);
and U14192 (N_14192,N_12577,N_12692);
nand U14193 (N_14193,N_13056,N_12798);
xnor U14194 (N_14194,N_13331,N_13457);
nand U14195 (N_14195,N_12177,N_12954);
nor U14196 (N_14196,N_12051,N_12791);
nand U14197 (N_14197,N_13111,N_12568);
nor U14198 (N_14198,N_12357,N_13223);
nand U14199 (N_14199,N_13408,N_13010);
and U14200 (N_14200,N_12848,N_12801);
or U14201 (N_14201,N_12347,N_12365);
or U14202 (N_14202,N_13222,N_12322);
nor U14203 (N_14203,N_13210,N_12480);
nor U14204 (N_14204,N_13087,N_13204);
nor U14205 (N_14205,N_12406,N_13066);
nand U14206 (N_14206,N_12194,N_13332);
or U14207 (N_14207,N_13431,N_12000);
and U14208 (N_14208,N_13306,N_12199);
nor U14209 (N_14209,N_12239,N_12216);
and U14210 (N_14210,N_12571,N_12891);
and U14211 (N_14211,N_12870,N_12113);
nor U14212 (N_14212,N_13041,N_12761);
nor U14213 (N_14213,N_12649,N_13424);
nand U14214 (N_14214,N_12793,N_12788);
or U14215 (N_14215,N_13052,N_13043);
or U14216 (N_14216,N_13085,N_12873);
or U14217 (N_14217,N_12374,N_12465);
nor U14218 (N_14218,N_12716,N_12114);
or U14219 (N_14219,N_12332,N_12529);
or U14220 (N_14220,N_12361,N_13146);
or U14221 (N_14221,N_13083,N_12282);
and U14222 (N_14222,N_13392,N_12726);
and U14223 (N_14223,N_12958,N_13281);
nor U14224 (N_14224,N_12153,N_12961);
nand U14225 (N_14225,N_12016,N_13324);
or U14226 (N_14226,N_13236,N_12450);
and U14227 (N_14227,N_12928,N_12119);
nand U14228 (N_14228,N_13065,N_12355);
nand U14229 (N_14229,N_13388,N_13446);
nand U14230 (N_14230,N_12507,N_12922);
or U14231 (N_14231,N_12547,N_12370);
nand U14232 (N_14232,N_13390,N_12208);
and U14233 (N_14233,N_12381,N_13193);
nor U14234 (N_14234,N_12066,N_13344);
nand U14235 (N_14235,N_13219,N_12662);
and U14236 (N_14236,N_12395,N_12700);
xnor U14237 (N_14237,N_13467,N_12167);
nor U14238 (N_14238,N_12240,N_12526);
nand U14239 (N_14239,N_12932,N_13416);
nor U14240 (N_14240,N_12310,N_13170);
xor U14241 (N_14241,N_13205,N_12030);
or U14242 (N_14242,N_12474,N_13402);
nand U14243 (N_14243,N_13479,N_12867);
and U14244 (N_14244,N_12295,N_13138);
nand U14245 (N_14245,N_13240,N_12742);
and U14246 (N_14246,N_13475,N_13428);
nand U14247 (N_14247,N_13096,N_13226);
and U14248 (N_14248,N_12660,N_13247);
and U14249 (N_14249,N_12342,N_12963);
and U14250 (N_14250,N_12670,N_12222);
nor U14251 (N_14251,N_12496,N_12986);
nand U14252 (N_14252,N_12334,N_12509);
xnor U14253 (N_14253,N_12954,N_13371);
xnor U14254 (N_14254,N_12795,N_13080);
nor U14255 (N_14255,N_13012,N_12577);
nor U14256 (N_14256,N_12063,N_13158);
and U14257 (N_14257,N_12130,N_12606);
nor U14258 (N_14258,N_12860,N_13329);
nand U14259 (N_14259,N_12398,N_12299);
nand U14260 (N_14260,N_13292,N_12212);
xor U14261 (N_14261,N_12115,N_13289);
and U14262 (N_14262,N_13206,N_13145);
and U14263 (N_14263,N_12344,N_13130);
or U14264 (N_14264,N_13285,N_12650);
or U14265 (N_14265,N_13026,N_12363);
nand U14266 (N_14266,N_12290,N_12665);
or U14267 (N_14267,N_12607,N_12612);
and U14268 (N_14268,N_13397,N_12665);
or U14269 (N_14269,N_13450,N_12191);
xnor U14270 (N_14270,N_12422,N_12912);
xor U14271 (N_14271,N_12859,N_13188);
and U14272 (N_14272,N_12871,N_13119);
and U14273 (N_14273,N_13473,N_12526);
and U14274 (N_14274,N_12491,N_13298);
nand U14275 (N_14275,N_12280,N_13152);
nor U14276 (N_14276,N_13347,N_12969);
nand U14277 (N_14277,N_13053,N_12396);
xor U14278 (N_14278,N_12492,N_12861);
and U14279 (N_14279,N_13277,N_13373);
and U14280 (N_14280,N_12923,N_12763);
or U14281 (N_14281,N_12582,N_13140);
or U14282 (N_14282,N_12102,N_13496);
and U14283 (N_14283,N_12088,N_12336);
and U14284 (N_14284,N_12720,N_12443);
and U14285 (N_14285,N_12321,N_12422);
nand U14286 (N_14286,N_12409,N_12358);
nand U14287 (N_14287,N_12094,N_12867);
or U14288 (N_14288,N_12088,N_12565);
nor U14289 (N_14289,N_13123,N_12237);
nor U14290 (N_14290,N_12748,N_12566);
nand U14291 (N_14291,N_12562,N_13003);
or U14292 (N_14292,N_12872,N_12867);
and U14293 (N_14293,N_12538,N_12132);
or U14294 (N_14294,N_12835,N_12320);
and U14295 (N_14295,N_13401,N_12272);
nand U14296 (N_14296,N_13335,N_12075);
and U14297 (N_14297,N_13229,N_12542);
nand U14298 (N_14298,N_13042,N_12883);
nor U14299 (N_14299,N_12694,N_12972);
and U14300 (N_14300,N_12239,N_12287);
or U14301 (N_14301,N_12347,N_12970);
xnor U14302 (N_14302,N_12774,N_12024);
nand U14303 (N_14303,N_13274,N_12088);
nor U14304 (N_14304,N_12978,N_13417);
and U14305 (N_14305,N_12986,N_12864);
xor U14306 (N_14306,N_12142,N_12823);
nor U14307 (N_14307,N_12855,N_13332);
and U14308 (N_14308,N_12181,N_12191);
xnor U14309 (N_14309,N_12731,N_13025);
nor U14310 (N_14310,N_13244,N_12822);
and U14311 (N_14311,N_13464,N_12536);
nor U14312 (N_14312,N_12108,N_13399);
nand U14313 (N_14313,N_13020,N_13310);
and U14314 (N_14314,N_12917,N_13297);
or U14315 (N_14315,N_12685,N_12316);
or U14316 (N_14316,N_13314,N_12930);
and U14317 (N_14317,N_13305,N_12308);
nand U14318 (N_14318,N_12591,N_12498);
or U14319 (N_14319,N_12048,N_12907);
or U14320 (N_14320,N_12784,N_12520);
or U14321 (N_14321,N_12751,N_12073);
nand U14322 (N_14322,N_13280,N_12722);
or U14323 (N_14323,N_12456,N_12963);
or U14324 (N_14324,N_12012,N_13105);
and U14325 (N_14325,N_12922,N_12187);
and U14326 (N_14326,N_12444,N_12599);
nor U14327 (N_14327,N_12615,N_13383);
nand U14328 (N_14328,N_12430,N_12311);
nand U14329 (N_14329,N_12636,N_13487);
xnor U14330 (N_14330,N_12685,N_12830);
nand U14331 (N_14331,N_13132,N_12149);
xor U14332 (N_14332,N_12205,N_13469);
nand U14333 (N_14333,N_12650,N_12409);
nand U14334 (N_14334,N_12230,N_13039);
and U14335 (N_14335,N_12685,N_12920);
or U14336 (N_14336,N_12606,N_12857);
nor U14337 (N_14337,N_12674,N_13054);
nor U14338 (N_14338,N_12262,N_12529);
or U14339 (N_14339,N_12980,N_12443);
nor U14340 (N_14340,N_13071,N_13091);
or U14341 (N_14341,N_12318,N_12055);
nor U14342 (N_14342,N_13381,N_13371);
and U14343 (N_14343,N_12151,N_13283);
nand U14344 (N_14344,N_12102,N_12206);
and U14345 (N_14345,N_13439,N_13173);
nor U14346 (N_14346,N_12381,N_12450);
nand U14347 (N_14347,N_12007,N_12874);
nor U14348 (N_14348,N_13084,N_13112);
and U14349 (N_14349,N_12842,N_12763);
and U14350 (N_14350,N_12897,N_13461);
and U14351 (N_14351,N_13352,N_12107);
nor U14352 (N_14352,N_12742,N_12404);
nor U14353 (N_14353,N_13357,N_13345);
or U14354 (N_14354,N_12813,N_12215);
or U14355 (N_14355,N_12685,N_12803);
nor U14356 (N_14356,N_12188,N_12548);
or U14357 (N_14357,N_13328,N_13491);
or U14358 (N_14358,N_12111,N_12623);
or U14359 (N_14359,N_13300,N_12383);
or U14360 (N_14360,N_12076,N_12978);
and U14361 (N_14361,N_12849,N_12819);
or U14362 (N_14362,N_12161,N_13046);
and U14363 (N_14363,N_12640,N_12818);
and U14364 (N_14364,N_12978,N_12698);
and U14365 (N_14365,N_12594,N_13323);
nor U14366 (N_14366,N_12412,N_13313);
nor U14367 (N_14367,N_12677,N_12384);
or U14368 (N_14368,N_12893,N_12344);
nand U14369 (N_14369,N_12781,N_12212);
xor U14370 (N_14370,N_12510,N_12887);
and U14371 (N_14371,N_13236,N_12941);
or U14372 (N_14372,N_13085,N_12538);
or U14373 (N_14373,N_12646,N_12997);
and U14374 (N_14374,N_13069,N_12996);
nor U14375 (N_14375,N_12450,N_13137);
and U14376 (N_14376,N_12547,N_12890);
or U14377 (N_14377,N_12572,N_12782);
or U14378 (N_14378,N_12337,N_13266);
nand U14379 (N_14379,N_13126,N_12000);
nand U14380 (N_14380,N_13220,N_13014);
nor U14381 (N_14381,N_13364,N_12848);
xor U14382 (N_14382,N_13217,N_13246);
xnor U14383 (N_14383,N_12942,N_13228);
nand U14384 (N_14384,N_13445,N_13206);
nor U14385 (N_14385,N_12365,N_12263);
nand U14386 (N_14386,N_12451,N_13029);
and U14387 (N_14387,N_12543,N_12333);
and U14388 (N_14388,N_12508,N_12526);
nor U14389 (N_14389,N_12093,N_12385);
or U14390 (N_14390,N_12103,N_12440);
and U14391 (N_14391,N_12552,N_13462);
nor U14392 (N_14392,N_13312,N_12869);
nand U14393 (N_14393,N_12637,N_13012);
nor U14394 (N_14394,N_12873,N_12649);
or U14395 (N_14395,N_12413,N_12198);
xor U14396 (N_14396,N_12592,N_12321);
or U14397 (N_14397,N_12758,N_12582);
nor U14398 (N_14398,N_13415,N_12057);
and U14399 (N_14399,N_12604,N_13468);
xor U14400 (N_14400,N_12664,N_13308);
and U14401 (N_14401,N_13161,N_13397);
or U14402 (N_14402,N_12500,N_12160);
nand U14403 (N_14403,N_13067,N_12562);
or U14404 (N_14404,N_13467,N_12298);
nand U14405 (N_14405,N_13356,N_13087);
nand U14406 (N_14406,N_12834,N_13202);
and U14407 (N_14407,N_12315,N_12682);
or U14408 (N_14408,N_12147,N_13208);
nor U14409 (N_14409,N_13421,N_12941);
or U14410 (N_14410,N_13210,N_13266);
and U14411 (N_14411,N_13497,N_12401);
nand U14412 (N_14412,N_12013,N_13439);
or U14413 (N_14413,N_12583,N_13189);
and U14414 (N_14414,N_13273,N_13005);
and U14415 (N_14415,N_12986,N_12972);
nor U14416 (N_14416,N_13356,N_13290);
xnor U14417 (N_14417,N_12946,N_12172);
and U14418 (N_14418,N_13196,N_12150);
or U14419 (N_14419,N_12096,N_13308);
or U14420 (N_14420,N_13156,N_12640);
or U14421 (N_14421,N_12964,N_12700);
and U14422 (N_14422,N_12524,N_13102);
or U14423 (N_14423,N_12639,N_12578);
or U14424 (N_14424,N_13060,N_12435);
nor U14425 (N_14425,N_13011,N_12482);
or U14426 (N_14426,N_12346,N_12131);
or U14427 (N_14427,N_12709,N_12057);
nor U14428 (N_14428,N_12030,N_13222);
xnor U14429 (N_14429,N_13098,N_13480);
nand U14430 (N_14430,N_13452,N_12434);
xor U14431 (N_14431,N_12085,N_13038);
and U14432 (N_14432,N_13147,N_12159);
and U14433 (N_14433,N_12844,N_13484);
or U14434 (N_14434,N_12371,N_12997);
nor U14435 (N_14435,N_12535,N_12472);
nor U14436 (N_14436,N_12554,N_13118);
or U14437 (N_14437,N_13354,N_13070);
or U14438 (N_14438,N_13007,N_12839);
or U14439 (N_14439,N_12412,N_13097);
nor U14440 (N_14440,N_12169,N_12533);
and U14441 (N_14441,N_12708,N_12267);
or U14442 (N_14442,N_13235,N_12966);
nand U14443 (N_14443,N_12206,N_13031);
and U14444 (N_14444,N_13013,N_12500);
and U14445 (N_14445,N_12731,N_12037);
xnor U14446 (N_14446,N_12992,N_12507);
or U14447 (N_14447,N_12811,N_12936);
nand U14448 (N_14448,N_13457,N_12224);
nor U14449 (N_14449,N_13251,N_12573);
nor U14450 (N_14450,N_12528,N_12611);
and U14451 (N_14451,N_12986,N_12772);
xnor U14452 (N_14452,N_13103,N_13387);
nand U14453 (N_14453,N_12190,N_12670);
nor U14454 (N_14454,N_12077,N_12979);
nor U14455 (N_14455,N_12171,N_12036);
or U14456 (N_14456,N_12995,N_13055);
or U14457 (N_14457,N_13428,N_12499);
nor U14458 (N_14458,N_13384,N_13482);
and U14459 (N_14459,N_13016,N_12834);
and U14460 (N_14460,N_13093,N_12102);
or U14461 (N_14461,N_12646,N_12472);
nor U14462 (N_14462,N_12618,N_12994);
or U14463 (N_14463,N_12106,N_13129);
nor U14464 (N_14464,N_12448,N_12896);
or U14465 (N_14465,N_13445,N_13180);
xor U14466 (N_14466,N_12183,N_12096);
nor U14467 (N_14467,N_12963,N_13044);
or U14468 (N_14468,N_13047,N_12302);
xnor U14469 (N_14469,N_12002,N_12653);
and U14470 (N_14470,N_13477,N_13225);
nor U14471 (N_14471,N_12248,N_12884);
nand U14472 (N_14472,N_12708,N_12145);
nor U14473 (N_14473,N_12824,N_13213);
and U14474 (N_14474,N_12530,N_12709);
and U14475 (N_14475,N_12464,N_12532);
nor U14476 (N_14476,N_12563,N_12561);
nand U14477 (N_14477,N_13197,N_12925);
nand U14478 (N_14478,N_12186,N_13419);
or U14479 (N_14479,N_12303,N_13170);
and U14480 (N_14480,N_13492,N_13296);
or U14481 (N_14481,N_12495,N_13210);
nor U14482 (N_14482,N_12518,N_12178);
or U14483 (N_14483,N_13061,N_12400);
xnor U14484 (N_14484,N_12928,N_13233);
and U14485 (N_14485,N_12091,N_13079);
nand U14486 (N_14486,N_12538,N_13069);
nor U14487 (N_14487,N_13103,N_12495);
and U14488 (N_14488,N_13195,N_12627);
nor U14489 (N_14489,N_13041,N_12778);
nor U14490 (N_14490,N_12176,N_12702);
nor U14491 (N_14491,N_12806,N_12079);
nand U14492 (N_14492,N_12766,N_12883);
xnor U14493 (N_14493,N_12472,N_12194);
or U14494 (N_14494,N_12785,N_13222);
nand U14495 (N_14495,N_13066,N_13295);
nor U14496 (N_14496,N_13254,N_12697);
and U14497 (N_14497,N_13474,N_13202);
nand U14498 (N_14498,N_13003,N_12614);
and U14499 (N_14499,N_12802,N_12621);
or U14500 (N_14500,N_12644,N_12363);
and U14501 (N_14501,N_12680,N_12746);
or U14502 (N_14502,N_12090,N_12866);
nand U14503 (N_14503,N_12949,N_12361);
or U14504 (N_14504,N_13125,N_12618);
nand U14505 (N_14505,N_13293,N_12194);
nand U14506 (N_14506,N_13398,N_12327);
nor U14507 (N_14507,N_13375,N_12348);
and U14508 (N_14508,N_12394,N_13211);
or U14509 (N_14509,N_12433,N_12835);
nor U14510 (N_14510,N_13152,N_13218);
or U14511 (N_14511,N_13083,N_12246);
and U14512 (N_14512,N_12573,N_12116);
nand U14513 (N_14513,N_13278,N_13266);
or U14514 (N_14514,N_12875,N_13064);
nor U14515 (N_14515,N_12994,N_13197);
nor U14516 (N_14516,N_12757,N_12526);
and U14517 (N_14517,N_12399,N_12542);
or U14518 (N_14518,N_13401,N_12942);
nor U14519 (N_14519,N_12582,N_12513);
and U14520 (N_14520,N_12107,N_13110);
and U14521 (N_14521,N_12351,N_12222);
nand U14522 (N_14522,N_13420,N_13307);
nor U14523 (N_14523,N_13031,N_12830);
and U14524 (N_14524,N_13064,N_12492);
nor U14525 (N_14525,N_12800,N_13325);
nor U14526 (N_14526,N_12497,N_13264);
and U14527 (N_14527,N_12445,N_12586);
xor U14528 (N_14528,N_12187,N_12890);
and U14529 (N_14529,N_12882,N_13050);
nand U14530 (N_14530,N_12766,N_12931);
or U14531 (N_14531,N_13308,N_13278);
and U14532 (N_14532,N_13232,N_12887);
and U14533 (N_14533,N_13462,N_13206);
and U14534 (N_14534,N_13150,N_12585);
and U14535 (N_14535,N_12005,N_12872);
or U14536 (N_14536,N_12402,N_12228);
and U14537 (N_14537,N_12005,N_12785);
nand U14538 (N_14538,N_12242,N_13033);
and U14539 (N_14539,N_12194,N_13097);
or U14540 (N_14540,N_12375,N_12786);
nand U14541 (N_14541,N_12925,N_12518);
or U14542 (N_14542,N_12191,N_12615);
or U14543 (N_14543,N_12877,N_12703);
or U14544 (N_14544,N_12450,N_12236);
nand U14545 (N_14545,N_12522,N_12333);
and U14546 (N_14546,N_13427,N_12712);
and U14547 (N_14547,N_12123,N_12233);
or U14548 (N_14548,N_12291,N_12884);
xor U14549 (N_14549,N_12864,N_12537);
and U14550 (N_14550,N_12461,N_13235);
nor U14551 (N_14551,N_12377,N_12602);
nor U14552 (N_14552,N_12614,N_13055);
and U14553 (N_14553,N_12016,N_13460);
and U14554 (N_14554,N_12946,N_13324);
or U14555 (N_14555,N_12520,N_13214);
or U14556 (N_14556,N_12273,N_12589);
xor U14557 (N_14557,N_13249,N_12068);
nand U14558 (N_14558,N_12906,N_12470);
nor U14559 (N_14559,N_13154,N_12255);
nor U14560 (N_14560,N_13136,N_12464);
nand U14561 (N_14561,N_12153,N_13021);
xnor U14562 (N_14562,N_12666,N_12191);
and U14563 (N_14563,N_13166,N_12934);
nand U14564 (N_14564,N_13059,N_12546);
or U14565 (N_14565,N_13169,N_12052);
or U14566 (N_14566,N_13345,N_12344);
xor U14567 (N_14567,N_12161,N_13334);
and U14568 (N_14568,N_13445,N_12205);
nor U14569 (N_14569,N_12209,N_12104);
nor U14570 (N_14570,N_13067,N_12307);
or U14571 (N_14571,N_12502,N_12860);
nand U14572 (N_14572,N_12083,N_12628);
or U14573 (N_14573,N_13137,N_12300);
nor U14574 (N_14574,N_12183,N_12574);
or U14575 (N_14575,N_12831,N_12243);
xor U14576 (N_14576,N_13293,N_12138);
or U14577 (N_14577,N_12819,N_13402);
or U14578 (N_14578,N_13025,N_12721);
nand U14579 (N_14579,N_13254,N_12777);
and U14580 (N_14580,N_13281,N_12646);
nor U14581 (N_14581,N_13007,N_12857);
nor U14582 (N_14582,N_12676,N_12379);
nor U14583 (N_14583,N_12297,N_12007);
or U14584 (N_14584,N_12890,N_12072);
and U14585 (N_14585,N_12309,N_12760);
and U14586 (N_14586,N_12649,N_13133);
and U14587 (N_14587,N_12595,N_13389);
or U14588 (N_14588,N_13155,N_13128);
or U14589 (N_14589,N_13314,N_12589);
nor U14590 (N_14590,N_12639,N_13359);
nor U14591 (N_14591,N_13152,N_13275);
nand U14592 (N_14592,N_12819,N_13162);
nor U14593 (N_14593,N_12739,N_13352);
xor U14594 (N_14594,N_12219,N_12684);
nor U14595 (N_14595,N_12413,N_12129);
and U14596 (N_14596,N_13119,N_12345);
nand U14597 (N_14597,N_12574,N_12394);
and U14598 (N_14598,N_12616,N_12280);
or U14599 (N_14599,N_13473,N_12931);
or U14600 (N_14600,N_12818,N_13013);
nand U14601 (N_14601,N_12859,N_12813);
and U14602 (N_14602,N_12761,N_12742);
or U14603 (N_14603,N_12170,N_12135);
or U14604 (N_14604,N_12766,N_12493);
nand U14605 (N_14605,N_12387,N_13428);
or U14606 (N_14606,N_12588,N_12006);
or U14607 (N_14607,N_12422,N_12057);
xor U14608 (N_14608,N_13326,N_12174);
nand U14609 (N_14609,N_12381,N_13375);
nand U14610 (N_14610,N_12118,N_12412);
nor U14611 (N_14611,N_13373,N_12878);
nor U14612 (N_14612,N_12347,N_12946);
nor U14613 (N_14613,N_12461,N_12649);
and U14614 (N_14614,N_13142,N_12564);
nor U14615 (N_14615,N_13336,N_12341);
xnor U14616 (N_14616,N_13453,N_12832);
nor U14617 (N_14617,N_12171,N_12245);
nor U14618 (N_14618,N_12594,N_13120);
nand U14619 (N_14619,N_13426,N_12657);
xnor U14620 (N_14620,N_12359,N_12601);
and U14621 (N_14621,N_13161,N_12284);
or U14622 (N_14622,N_13031,N_12783);
nand U14623 (N_14623,N_12883,N_12898);
nand U14624 (N_14624,N_13062,N_13158);
or U14625 (N_14625,N_12298,N_12223);
or U14626 (N_14626,N_12771,N_12429);
nor U14627 (N_14627,N_12478,N_13061);
nand U14628 (N_14628,N_13421,N_12706);
nor U14629 (N_14629,N_12664,N_13458);
and U14630 (N_14630,N_12179,N_13102);
nand U14631 (N_14631,N_12139,N_12576);
nand U14632 (N_14632,N_12887,N_12365);
nand U14633 (N_14633,N_12539,N_12835);
xnor U14634 (N_14634,N_12901,N_12260);
xor U14635 (N_14635,N_12313,N_12131);
nor U14636 (N_14636,N_12767,N_12049);
nand U14637 (N_14637,N_12395,N_13415);
and U14638 (N_14638,N_12731,N_13203);
or U14639 (N_14639,N_12720,N_12724);
nor U14640 (N_14640,N_12224,N_12655);
nor U14641 (N_14641,N_12143,N_13097);
nand U14642 (N_14642,N_13022,N_12358);
or U14643 (N_14643,N_13386,N_12335);
or U14644 (N_14644,N_13306,N_12741);
nand U14645 (N_14645,N_12501,N_13271);
xnor U14646 (N_14646,N_13447,N_13356);
nor U14647 (N_14647,N_13208,N_12031);
nor U14648 (N_14648,N_13219,N_12575);
nor U14649 (N_14649,N_13184,N_13083);
or U14650 (N_14650,N_12564,N_12103);
nor U14651 (N_14651,N_12451,N_13142);
nor U14652 (N_14652,N_12797,N_13193);
or U14653 (N_14653,N_13440,N_13009);
xor U14654 (N_14654,N_12411,N_13438);
and U14655 (N_14655,N_12256,N_12427);
or U14656 (N_14656,N_13310,N_12922);
nand U14657 (N_14657,N_12362,N_12338);
and U14658 (N_14658,N_13079,N_12648);
and U14659 (N_14659,N_12189,N_12951);
nand U14660 (N_14660,N_13300,N_12522);
nand U14661 (N_14661,N_12768,N_12262);
nor U14662 (N_14662,N_12477,N_12025);
nand U14663 (N_14663,N_12483,N_13271);
and U14664 (N_14664,N_12248,N_12681);
nor U14665 (N_14665,N_13481,N_12017);
or U14666 (N_14666,N_12861,N_13073);
nor U14667 (N_14667,N_13442,N_12983);
nor U14668 (N_14668,N_12261,N_12164);
nor U14669 (N_14669,N_12080,N_12634);
or U14670 (N_14670,N_12438,N_12029);
nor U14671 (N_14671,N_13196,N_13374);
nor U14672 (N_14672,N_13175,N_13088);
nand U14673 (N_14673,N_13452,N_13401);
nor U14674 (N_14674,N_12275,N_13054);
and U14675 (N_14675,N_13295,N_13296);
nand U14676 (N_14676,N_12873,N_12536);
nand U14677 (N_14677,N_13287,N_13384);
or U14678 (N_14678,N_12351,N_12376);
or U14679 (N_14679,N_12106,N_12038);
and U14680 (N_14680,N_13294,N_12160);
and U14681 (N_14681,N_12232,N_12102);
nor U14682 (N_14682,N_13314,N_12903);
xnor U14683 (N_14683,N_12424,N_12569);
nor U14684 (N_14684,N_12157,N_13168);
and U14685 (N_14685,N_12861,N_12364);
and U14686 (N_14686,N_13430,N_12343);
nand U14687 (N_14687,N_12458,N_12262);
or U14688 (N_14688,N_13180,N_13133);
nand U14689 (N_14689,N_12256,N_12472);
nand U14690 (N_14690,N_13337,N_12934);
or U14691 (N_14691,N_12483,N_13240);
nor U14692 (N_14692,N_13044,N_12852);
nand U14693 (N_14693,N_13249,N_12327);
xnor U14694 (N_14694,N_12350,N_12499);
or U14695 (N_14695,N_12741,N_12398);
xor U14696 (N_14696,N_13068,N_12492);
and U14697 (N_14697,N_12084,N_13362);
nor U14698 (N_14698,N_12837,N_12783);
nand U14699 (N_14699,N_12642,N_12326);
nand U14700 (N_14700,N_12082,N_13459);
nor U14701 (N_14701,N_12204,N_13411);
nand U14702 (N_14702,N_12829,N_13243);
and U14703 (N_14703,N_12706,N_12127);
and U14704 (N_14704,N_12543,N_12540);
nor U14705 (N_14705,N_13485,N_12695);
nand U14706 (N_14706,N_12969,N_12183);
nand U14707 (N_14707,N_13491,N_13079);
nand U14708 (N_14708,N_13014,N_12422);
xor U14709 (N_14709,N_13013,N_12269);
and U14710 (N_14710,N_13339,N_13479);
nor U14711 (N_14711,N_12443,N_12665);
nand U14712 (N_14712,N_13321,N_13296);
and U14713 (N_14713,N_12070,N_12344);
and U14714 (N_14714,N_13310,N_12636);
nand U14715 (N_14715,N_13404,N_12136);
and U14716 (N_14716,N_12106,N_12240);
nor U14717 (N_14717,N_13450,N_12846);
xnor U14718 (N_14718,N_12871,N_13038);
nand U14719 (N_14719,N_12190,N_13186);
nand U14720 (N_14720,N_13334,N_12185);
nand U14721 (N_14721,N_13474,N_12061);
or U14722 (N_14722,N_12595,N_13477);
and U14723 (N_14723,N_12888,N_13378);
nand U14724 (N_14724,N_12095,N_13143);
xnor U14725 (N_14725,N_12014,N_13380);
nand U14726 (N_14726,N_12906,N_13434);
and U14727 (N_14727,N_12521,N_12009);
nand U14728 (N_14728,N_13282,N_12358);
and U14729 (N_14729,N_13173,N_12964);
nand U14730 (N_14730,N_12752,N_12983);
or U14731 (N_14731,N_13275,N_13144);
xnor U14732 (N_14732,N_12194,N_13484);
nand U14733 (N_14733,N_13417,N_12708);
xnor U14734 (N_14734,N_12749,N_13081);
nand U14735 (N_14735,N_13227,N_12369);
nand U14736 (N_14736,N_12386,N_13295);
nand U14737 (N_14737,N_12558,N_13397);
or U14738 (N_14738,N_12578,N_13126);
nand U14739 (N_14739,N_12872,N_13413);
nor U14740 (N_14740,N_13459,N_12190);
nand U14741 (N_14741,N_12584,N_12548);
xnor U14742 (N_14742,N_13065,N_13352);
or U14743 (N_14743,N_12602,N_13317);
nor U14744 (N_14744,N_12924,N_12529);
xnor U14745 (N_14745,N_13207,N_12306);
and U14746 (N_14746,N_12230,N_12912);
nand U14747 (N_14747,N_12311,N_13242);
nand U14748 (N_14748,N_12375,N_12626);
nor U14749 (N_14749,N_12900,N_12765);
nor U14750 (N_14750,N_12157,N_13181);
nor U14751 (N_14751,N_13331,N_13283);
and U14752 (N_14752,N_12567,N_12007);
nand U14753 (N_14753,N_12713,N_12715);
xnor U14754 (N_14754,N_12272,N_12799);
or U14755 (N_14755,N_12844,N_13225);
nor U14756 (N_14756,N_13310,N_12566);
nand U14757 (N_14757,N_12588,N_12834);
nor U14758 (N_14758,N_13314,N_12531);
or U14759 (N_14759,N_12041,N_12128);
and U14760 (N_14760,N_12414,N_12286);
or U14761 (N_14761,N_13222,N_13484);
nor U14762 (N_14762,N_13127,N_12842);
xnor U14763 (N_14763,N_13241,N_13012);
nor U14764 (N_14764,N_12308,N_12865);
or U14765 (N_14765,N_12403,N_12696);
or U14766 (N_14766,N_12824,N_12806);
nand U14767 (N_14767,N_12911,N_12964);
or U14768 (N_14768,N_12453,N_12035);
or U14769 (N_14769,N_12768,N_12481);
xor U14770 (N_14770,N_12633,N_12980);
or U14771 (N_14771,N_12025,N_12597);
nor U14772 (N_14772,N_13424,N_13272);
nand U14773 (N_14773,N_13244,N_12837);
nand U14774 (N_14774,N_12362,N_13307);
and U14775 (N_14775,N_13132,N_12807);
nor U14776 (N_14776,N_12014,N_12132);
nor U14777 (N_14777,N_13414,N_13338);
nand U14778 (N_14778,N_12769,N_13028);
nor U14779 (N_14779,N_12448,N_13259);
and U14780 (N_14780,N_12720,N_12103);
or U14781 (N_14781,N_12721,N_12410);
and U14782 (N_14782,N_13268,N_12888);
and U14783 (N_14783,N_12313,N_12309);
nand U14784 (N_14784,N_13439,N_12543);
xor U14785 (N_14785,N_13402,N_13284);
or U14786 (N_14786,N_12426,N_13163);
and U14787 (N_14787,N_12721,N_12649);
and U14788 (N_14788,N_12622,N_12825);
and U14789 (N_14789,N_12110,N_13097);
nand U14790 (N_14790,N_13162,N_13288);
nor U14791 (N_14791,N_12572,N_12526);
or U14792 (N_14792,N_12742,N_12960);
or U14793 (N_14793,N_12873,N_12730);
nand U14794 (N_14794,N_12458,N_12735);
nor U14795 (N_14795,N_13290,N_12937);
xor U14796 (N_14796,N_13484,N_12166);
and U14797 (N_14797,N_12985,N_12672);
or U14798 (N_14798,N_13387,N_13161);
or U14799 (N_14799,N_13499,N_12125);
nand U14800 (N_14800,N_12918,N_13405);
xor U14801 (N_14801,N_12212,N_13080);
or U14802 (N_14802,N_12207,N_13479);
nor U14803 (N_14803,N_12964,N_12805);
or U14804 (N_14804,N_13005,N_13177);
xnor U14805 (N_14805,N_13010,N_12621);
nand U14806 (N_14806,N_12361,N_13482);
and U14807 (N_14807,N_12684,N_12763);
and U14808 (N_14808,N_12216,N_13241);
nor U14809 (N_14809,N_12470,N_13375);
nand U14810 (N_14810,N_12805,N_13250);
or U14811 (N_14811,N_12311,N_13196);
nand U14812 (N_14812,N_13238,N_12442);
nor U14813 (N_14813,N_12839,N_12627);
xnor U14814 (N_14814,N_12503,N_13382);
nand U14815 (N_14815,N_12756,N_12758);
or U14816 (N_14816,N_13488,N_12914);
or U14817 (N_14817,N_13209,N_12653);
nor U14818 (N_14818,N_13478,N_13331);
xnor U14819 (N_14819,N_12488,N_12138);
nor U14820 (N_14820,N_12919,N_12927);
nor U14821 (N_14821,N_13153,N_12186);
and U14822 (N_14822,N_13182,N_12397);
and U14823 (N_14823,N_13294,N_13026);
or U14824 (N_14824,N_13372,N_12283);
nand U14825 (N_14825,N_12347,N_13155);
or U14826 (N_14826,N_13407,N_12466);
nand U14827 (N_14827,N_13316,N_12540);
nor U14828 (N_14828,N_12215,N_12198);
and U14829 (N_14829,N_13023,N_12008);
nor U14830 (N_14830,N_12598,N_13003);
nand U14831 (N_14831,N_12646,N_12016);
or U14832 (N_14832,N_12755,N_12430);
and U14833 (N_14833,N_12799,N_13151);
nand U14834 (N_14834,N_12852,N_12414);
xnor U14835 (N_14835,N_12856,N_12054);
nand U14836 (N_14836,N_12122,N_12526);
nor U14837 (N_14837,N_12271,N_12997);
nand U14838 (N_14838,N_13486,N_12591);
nor U14839 (N_14839,N_12574,N_12365);
nand U14840 (N_14840,N_12348,N_12547);
xnor U14841 (N_14841,N_12738,N_12670);
nor U14842 (N_14842,N_12469,N_12753);
and U14843 (N_14843,N_12510,N_13011);
or U14844 (N_14844,N_13214,N_12640);
and U14845 (N_14845,N_12028,N_12532);
and U14846 (N_14846,N_12254,N_13463);
and U14847 (N_14847,N_12440,N_12989);
nand U14848 (N_14848,N_13048,N_13056);
or U14849 (N_14849,N_13473,N_12134);
or U14850 (N_14850,N_12625,N_12592);
nor U14851 (N_14851,N_13377,N_12187);
and U14852 (N_14852,N_13364,N_12506);
nor U14853 (N_14853,N_13130,N_12490);
nor U14854 (N_14854,N_12295,N_12237);
or U14855 (N_14855,N_13279,N_12640);
or U14856 (N_14856,N_12577,N_12376);
and U14857 (N_14857,N_12793,N_12370);
nand U14858 (N_14858,N_12537,N_12278);
nand U14859 (N_14859,N_12634,N_13431);
or U14860 (N_14860,N_13062,N_12975);
or U14861 (N_14861,N_12749,N_12617);
nor U14862 (N_14862,N_12096,N_12215);
or U14863 (N_14863,N_13322,N_12406);
nor U14864 (N_14864,N_12783,N_12288);
and U14865 (N_14865,N_12930,N_12363);
nor U14866 (N_14866,N_13215,N_13192);
or U14867 (N_14867,N_12592,N_13355);
or U14868 (N_14868,N_13019,N_13058);
nand U14869 (N_14869,N_13074,N_12567);
nor U14870 (N_14870,N_13490,N_12288);
nor U14871 (N_14871,N_12220,N_12304);
and U14872 (N_14872,N_13466,N_13024);
nor U14873 (N_14873,N_12130,N_12137);
and U14874 (N_14874,N_13422,N_12098);
nand U14875 (N_14875,N_12052,N_12025);
nand U14876 (N_14876,N_12639,N_12674);
nand U14877 (N_14877,N_12252,N_12857);
and U14878 (N_14878,N_12994,N_12218);
and U14879 (N_14879,N_12821,N_12441);
nand U14880 (N_14880,N_12569,N_13395);
nor U14881 (N_14881,N_13069,N_13478);
nand U14882 (N_14882,N_12083,N_12744);
nand U14883 (N_14883,N_13213,N_12322);
nand U14884 (N_14884,N_12593,N_13185);
nor U14885 (N_14885,N_13300,N_13450);
or U14886 (N_14886,N_12699,N_12051);
or U14887 (N_14887,N_13216,N_12444);
nor U14888 (N_14888,N_12747,N_13068);
nand U14889 (N_14889,N_12502,N_12124);
nor U14890 (N_14890,N_12604,N_12691);
nand U14891 (N_14891,N_13185,N_12905);
or U14892 (N_14892,N_12103,N_12615);
nor U14893 (N_14893,N_12836,N_12708);
or U14894 (N_14894,N_12030,N_12326);
or U14895 (N_14895,N_13015,N_13392);
nand U14896 (N_14896,N_13423,N_12255);
and U14897 (N_14897,N_13252,N_12696);
nor U14898 (N_14898,N_12387,N_12214);
nor U14899 (N_14899,N_12017,N_12475);
nor U14900 (N_14900,N_13278,N_12161);
and U14901 (N_14901,N_12501,N_12018);
and U14902 (N_14902,N_12980,N_13034);
nand U14903 (N_14903,N_12410,N_12070);
or U14904 (N_14904,N_12177,N_12665);
and U14905 (N_14905,N_12502,N_12437);
nor U14906 (N_14906,N_13491,N_12804);
nor U14907 (N_14907,N_12547,N_13264);
xnor U14908 (N_14908,N_12713,N_12522);
nor U14909 (N_14909,N_13102,N_12688);
or U14910 (N_14910,N_12934,N_13324);
xnor U14911 (N_14911,N_13335,N_12264);
nor U14912 (N_14912,N_13458,N_13142);
nand U14913 (N_14913,N_12452,N_13201);
nor U14914 (N_14914,N_13493,N_12167);
and U14915 (N_14915,N_13317,N_13369);
or U14916 (N_14916,N_12063,N_12830);
and U14917 (N_14917,N_12261,N_12673);
xnor U14918 (N_14918,N_12116,N_12845);
nor U14919 (N_14919,N_12684,N_12328);
or U14920 (N_14920,N_12340,N_12748);
or U14921 (N_14921,N_13404,N_12446);
nand U14922 (N_14922,N_12132,N_12152);
and U14923 (N_14923,N_12656,N_12341);
nor U14924 (N_14924,N_12718,N_12278);
nand U14925 (N_14925,N_13135,N_13065);
nor U14926 (N_14926,N_12003,N_12321);
or U14927 (N_14927,N_13352,N_13248);
or U14928 (N_14928,N_12083,N_12016);
or U14929 (N_14929,N_12463,N_12309);
or U14930 (N_14930,N_12166,N_13255);
or U14931 (N_14931,N_12111,N_12322);
nand U14932 (N_14932,N_12503,N_12507);
nand U14933 (N_14933,N_12209,N_13424);
and U14934 (N_14934,N_12092,N_13033);
or U14935 (N_14935,N_12474,N_13301);
or U14936 (N_14936,N_13213,N_12074);
nor U14937 (N_14937,N_12127,N_12914);
nand U14938 (N_14938,N_12532,N_12193);
nand U14939 (N_14939,N_12569,N_12699);
xnor U14940 (N_14940,N_12884,N_12797);
nand U14941 (N_14941,N_12984,N_12994);
nand U14942 (N_14942,N_13295,N_12915);
or U14943 (N_14943,N_12542,N_12506);
nor U14944 (N_14944,N_13209,N_13337);
or U14945 (N_14945,N_12387,N_13298);
or U14946 (N_14946,N_13453,N_13043);
nor U14947 (N_14947,N_12936,N_12529);
nor U14948 (N_14948,N_12393,N_12263);
and U14949 (N_14949,N_13015,N_12623);
and U14950 (N_14950,N_12226,N_12980);
and U14951 (N_14951,N_13099,N_12865);
nand U14952 (N_14952,N_13068,N_13282);
or U14953 (N_14953,N_12847,N_13217);
xnor U14954 (N_14954,N_12709,N_12722);
xor U14955 (N_14955,N_12435,N_12737);
nand U14956 (N_14956,N_12801,N_12387);
and U14957 (N_14957,N_12212,N_13032);
and U14958 (N_14958,N_13131,N_12778);
nor U14959 (N_14959,N_12973,N_12876);
nor U14960 (N_14960,N_12521,N_13112);
nand U14961 (N_14961,N_13260,N_12099);
nor U14962 (N_14962,N_12363,N_12166);
nor U14963 (N_14963,N_12725,N_12317);
or U14964 (N_14964,N_12437,N_12141);
and U14965 (N_14965,N_13341,N_12346);
nand U14966 (N_14966,N_12310,N_12785);
and U14967 (N_14967,N_12426,N_12668);
or U14968 (N_14968,N_12362,N_12156);
xnor U14969 (N_14969,N_12090,N_12790);
nand U14970 (N_14970,N_12530,N_12681);
or U14971 (N_14971,N_12412,N_13393);
and U14972 (N_14972,N_12644,N_13328);
and U14973 (N_14973,N_13128,N_12271);
nand U14974 (N_14974,N_13072,N_12430);
and U14975 (N_14975,N_13491,N_13166);
xnor U14976 (N_14976,N_12641,N_13473);
nor U14977 (N_14977,N_12783,N_12984);
or U14978 (N_14978,N_13124,N_12539);
and U14979 (N_14979,N_12818,N_12855);
and U14980 (N_14980,N_13389,N_13187);
and U14981 (N_14981,N_12676,N_12190);
nand U14982 (N_14982,N_12311,N_13246);
nor U14983 (N_14983,N_12618,N_13223);
nor U14984 (N_14984,N_12115,N_12282);
nand U14985 (N_14985,N_13490,N_13476);
nand U14986 (N_14986,N_12415,N_13452);
or U14987 (N_14987,N_12853,N_12850);
xor U14988 (N_14988,N_12995,N_12070);
or U14989 (N_14989,N_12945,N_12891);
xnor U14990 (N_14990,N_12657,N_12236);
nand U14991 (N_14991,N_12302,N_12548);
nor U14992 (N_14992,N_12107,N_12457);
and U14993 (N_14993,N_13403,N_13385);
or U14994 (N_14994,N_13287,N_13169);
nand U14995 (N_14995,N_12338,N_12778);
and U14996 (N_14996,N_12625,N_12639);
or U14997 (N_14997,N_13306,N_12069);
or U14998 (N_14998,N_12186,N_13397);
and U14999 (N_14999,N_12688,N_12220);
nand UO_0 (O_0,N_14885,N_13897);
xnor UO_1 (O_1,N_14379,N_14735);
nand UO_2 (O_2,N_13591,N_13501);
or UO_3 (O_3,N_14254,N_14375);
nand UO_4 (O_4,N_13988,N_13791);
nand UO_5 (O_5,N_14488,N_14427);
or UO_6 (O_6,N_14041,N_13911);
and UO_7 (O_7,N_14639,N_14596);
or UO_8 (O_8,N_13899,N_13901);
nor UO_9 (O_9,N_14408,N_13996);
nand UO_10 (O_10,N_14872,N_14274);
or UO_11 (O_11,N_13903,N_14657);
nand UO_12 (O_12,N_14925,N_13752);
and UO_13 (O_13,N_14163,N_13835);
or UO_14 (O_14,N_14996,N_14446);
xor UO_15 (O_15,N_14865,N_13548);
or UO_16 (O_16,N_14185,N_14043);
nor UO_17 (O_17,N_14524,N_13614);
or UO_18 (O_18,N_14636,N_14541);
nor UO_19 (O_19,N_14417,N_14745);
nand UO_20 (O_20,N_13886,N_14780);
or UO_21 (O_21,N_14281,N_14299);
nand UO_22 (O_22,N_13627,N_13601);
or UO_23 (O_23,N_13561,N_14268);
or UO_24 (O_24,N_14118,N_14309);
nor UO_25 (O_25,N_13979,N_13722);
and UO_26 (O_26,N_14455,N_14114);
nor UO_27 (O_27,N_14181,N_14791);
or UO_28 (O_28,N_14108,N_13829);
or UO_29 (O_29,N_14470,N_14969);
nor UO_30 (O_30,N_14562,N_13740);
xnor UO_31 (O_31,N_14617,N_14345);
nand UO_32 (O_32,N_14081,N_13851);
nor UO_33 (O_33,N_14390,N_14095);
nand UO_34 (O_34,N_14728,N_14710);
and UO_35 (O_35,N_14014,N_14863);
nor UO_36 (O_36,N_14204,N_13794);
xnor UO_37 (O_37,N_13852,N_14898);
nand UO_38 (O_38,N_14968,N_14125);
or UO_39 (O_39,N_13802,N_13636);
or UO_40 (O_40,N_14838,N_13702);
xor UO_41 (O_41,N_14154,N_13849);
nor UO_42 (O_42,N_13952,N_13573);
and UO_43 (O_43,N_14992,N_14907);
nor UO_44 (O_44,N_13860,N_14071);
xor UO_45 (O_45,N_13567,N_13533);
and UO_46 (O_46,N_13750,N_14187);
nand UO_47 (O_47,N_14628,N_14753);
or UO_48 (O_48,N_14297,N_14474);
and UO_49 (O_49,N_13867,N_14800);
and UO_50 (O_50,N_14117,N_14141);
and UO_51 (O_51,N_14960,N_13795);
and UO_52 (O_52,N_14211,N_14327);
nor UO_53 (O_53,N_14788,N_14210);
or UO_54 (O_54,N_14483,N_14526);
or UO_55 (O_55,N_13539,N_13887);
nand UO_56 (O_56,N_13900,N_14381);
nor UO_57 (O_57,N_13701,N_14650);
nor UO_58 (O_58,N_14076,N_14138);
and UO_59 (O_59,N_14904,N_14684);
nand UO_60 (O_60,N_13699,N_14202);
nand UO_61 (O_61,N_14576,N_14671);
and UO_62 (O_62,N_14269,N_14631);
nor UO_63 (O_63,N_14497,N_14449);
nor UO_64 (O_64,N_13956,N_14803);
and UO_65 (O_65,N_14597,N_14761);
nor UO_66 (O_66,N_13871,N_14936);
nor UO_67 (O_67,N_13650,N_14926);
or UO_68 (O_68,N_13667,N_14359);
nand UO_69 (O_69,N_13678,N_14815);
nand UO_70 (O_70,N_13960,N_13938);
or UO_71 (O_71,N_14280,N_13883);
nand UO_72 (O_72,N_13626,N_13955);
and UO_73 (O_73,N_14683,N_14689);
or UO_74 (O_74,N_13904,N_14847);
nor UO_75 (O_75,N_13719,N_13912);
nor UO_76 (O_76,N_14927,N_14466);
nor UO_77 (O_77,N_14307,N_14468);
nor UO_78 (O_78,N_13930,N_13821);
nand UO_79 (O_79,N_13859,N_14962);
xnor UO_80 (O_80,N_14718,N_14073);
xor UO_81 (O_81,N_13727,N_13959);
nor UO_82 (O_82,N_14638,N_14190);
xor UO_83 (O_83,N_13595,N_13672);
or UO_84 (O_84,N_14313,N_13580);
or UO_85 (O_85,N_13680,N_14422);
nor UO_86 (O_86,N_14743,N_14682);
nand UO_87 (O_87,N_13758,N_14932);
nor UO_88 (O_88,N_14382,N_14456);
nand UO_89 (O_89,N_13906,N_13850);
nor UO_90 (O_90,N_14952,N_14048);
nor UO_91 (O_91,N_14388,N_14373);
and UO_92 (O_92,N_14467,N_13820);
nor UO_93 (O_93,N_14981,N_13826);
or UO_94 (O_94,N_14731,N_14206);
and UO_95 (O_95,N_13577,N_14471);
and UO_96 (O_96,N_14661,N_14400);
and UO_97 (O_97,N_13766,N_14599);
nand UO_98 (O_98,N_13894,N_14762);
nor UO_99 (O_99,N_13877,N_14620);
and UO_100 (O_100,N_14173,N_14544);
xor UO_101 (O_101,N_14558,N_14700);
and UO_102 (O_102,N_13570,N_14880);
or UO_103 (O_103,N_14160,N_13676);
nor UO_104 (O_104,N_14476,N_14737);
and UO_105 (O_105,N_14458,N_14389);
or UO_106 (O_106,N_14836,N_13962);
and UO_107 (O_107,N_14984,N_13888);
and UO_108 (O_108,N_14287,N_14873);
nand UO_109 (O_109,N_14464,N_13884);
and UO_110 (O_110,N_14993,N_13926);
and UO_111 (O_111,N_14922,N_14510);
nand UO_112 (O_112,N_13568,N_13585);
nand UO_113 (O_113,N_13932,N_14738);
nand UO_114 (O_114,N_14266,N_13958);
nor UO_115 (O_115,N_14401,N_14222);
or UO_116 (O_116,N_13527,N_14943);
nand UO_117 (O_117,N_14088,N_14424);
and UO_118 (O_118,N_14176,N_14941);
nor UO_119 (O_119,N_14583,N_14227);
and UO_120 (O_120,N_14491,N_13770);
and UO_121 (O_121,N_14888,N_13939);
or UO_122 (O_122,N_14033,N_14957);
or UO_123 (O_123,N_14161,N_14890);
or UO_124 (O_124,N_14040,N_14714);
or UO_125 (O_125,N_13554,N_13753);
nor UO_126 (O_126,N_14075,N_14336);
and UO_127 (O_127,N_14812,N_14241);
nand UO_128 (O_128,N_13870,N_14180);
or UO_129 (O_129,N_13518,N_14035);
or UO_130 (O_130,N_14963,N_13616);
nand UO_131 (O_131,N_14523,N_13658);
xor UO_132 (O_132,N_14273,N_14600);
nor UO_133 (O_133,N_13604,N_14525);
xor UO_134 (O_134,N_14658,N_14403);
nand UO_135 (O_135,N_14126,N_14421);
nand UO_136 (O_136,N_13519,N_14964);
or UO_137 (O_137,N_13671,N_13981);
nor UO_138 (O_138,N_13982,N_14263);
nand UO_139 (O_139,N_14262,N_13504);
nor UO_140 (O_140,N_14619,N_13510);
and UO_141 (O_141,N_13892,N_14027);
and UO_142 (O_142,N_14770,N_14635);
nor UO_143 (O_143,N_14844,N_14802);
xnor UO_144 (O_144,N_14586,N_14061);
and UO_145 (O_145,N_14675,N_13713);
and UO_146 (O_146,N_14825,N_14240);
or UO_147 (O_147,N_14605,N_14512);
or UO_148 (O_148,N_13738,N_13907);
nand UO_149 (O_149,N_13865,N_14997);
nand UO_150 (O_150,N_14787,N_13530);
nand UO_151 (O_151,N_13863,N_13605);
nor UO_152 (O_152,N_14191,N_13593);
and UO_153 (O_153,N_14648,N_14704);
nor UO_154 (O_154,N_14751,N_13505);
nand UO_155 (O_155,N_14411,N_13876);
and UO_156 (O_156,N_14056,N_13839);
nor UO_157 (O_157,N_14477,N_14022);
or UO_158 (O_158,N_14224,N_14514);
and UO_159 (O_159,N_14877,N_14221);
and UO_160 (O_160,N_14238,N_14332);
nand UO_161 (O_161,N_14829,N_14301);
or UO_162 (O_162,N_13603,N_14338);
xor UO_163 (O_163,N_13698,N_14921);
xor UO_164 (O_164,N_13746,N_14213);
nor UO_165 (O_165,N_14032,N_13972);
nand UO_166 (O_166,N_14604,N_14255);
or UO_167 (O_167,N_14613,N_13726);
nor UO_168 (O_168,N_13662,N_13708);
nor UO_169 (O_169,N_14341,N_13964);
nor UO_170 (O_170,N_13936,N_14598);
nand UO_171 (O_171,N_14113,N_13542);
nand UO_172 (O_172,N_14184,N_13633);
xor UO_173 (O_173,N_13660,N_13809);
or UO_174 (O_174,N_13824,N_13692);
nand UO_175 (O_175,N_14366,N_13575);
or UO_176 (O_176,N_13797,N_14031);
or UO_177 (O_177,N_14444,N_13862);
or UO_178 (O_178,N_13583,N_14895);
or UO_179 (O_179,N_14104,N_13923);
nand UO_180 (O_180,N_14734,N_14839);
and UO_181 (O_181,N_14492,N_14320);
nor UO_182 (O_182,N_13927,N_14150);
and UO_183 (O_183,N_14530,N_13931);
nor UO_184 (O_184,N_13754,N_13975);
or UO_185 (O_185,N_14264,N_13563);
and UO_186 (O_186,N_13748,N_13646);
or UO_187 (O_187,N_14773,N_14132);
and UO_188 (O_188,N_14654,N_14950);
or UO_189 (O_189,N_13917,N_14845);
nand UO_190 (O_190,N_13811,N_13584);
nand UO_191 (O_191,N_14995,N_13559);
nand UO_192 (O_192,N_14472,N_13810);
nor UO_193 (O_193,N_13875,N_14175);
and UO_194 (O_194,N_14517,N_14766);
nor UO_195 (O_195,N_14869,N_13711);
or UO_196 (O_196,N_14493,N_14858);
nor UO_197 (O_197,N_14391,N_14884);
nand UO_198 (O_198,N_13998,N_14854);
and UO_199 (O_199,N_13744,N_14402);
nand UO_200 (O_200,N_13558,N_14397);
nor UO_201 (O_201,N_13665,N_14096);
or UO_202 (O_202,N_14798,N_13789);
nand UO_203 (O_203,N_13745,N_14588);
xor UO_204 (O_204,N_14701,N_14833);
nand UO_205 (O_205,N_14271,N_14988);
and UO_206 (O_206,N_14171,N_13521);
nand UO_207 (O_207,N_14272,N_14900);
nor UO_208 (O_208,N_14496,N_14819);
nand UO_209 (O_209,N_14719,N_14298);
and UO_210 (O_210,N_14668,N_14087);
or UO_211 (O_211,N_14199,N_13919);
nor UO_212 (O_212,N_13589,N_13694);
nor UO_213 (O_213,N_14356,N_14246);
nand UO_214 (O_214,N_14404,N_14129);
xor UO_215 (O_215,N_14908,N_14503);
or UO_216 (O_216,N_13893,N_14824);
and UO_217 (O_217,N_13918,N_14674);
or UO_218 (O_218,N_13796,N_14678);
nand UO_219 (O_219,N_14127,N_14267);
and UO_220 (O_220,N_13957,N_13967);
xnor UO_221 (O_221,N_14808,N_14946);
and UO_222 (O_222,N_14178,N_14121);
or UO_223 (O_223,N_13823,N_14861);
nand UO_224 (O_224,N_14285,N_14352);
nand UO_225 (O_225,N_13514,N_13831);
nand UO_226 (O_226,N_14479,N_14923);
nand UO_227 (O_227,N_13793,N_13985);
or UO_228 (O_228,N_14256,N_14550);
or UO_229 (O_229,N_14316,N_14251);
nor UO_230 (O_230,N_14000,N_14448);
and UO_231 (O_231,N_14165,N_14367);
and UO_232 (O_232,N_14303,N_14876);
and UO_233 (O_233,N_14469,N_14655);
nand UO_234 (O_234,N_14857,N_13690);
nor UO_235 (O_235,N_13594,N_13717);
nand UO_236 (O_236,N_13649,N_14965);
or UO_237 (O_237,N_14693,N_14551);
nand UO_238 (O_238,N_14198,N_14547);
nand UO_239 (O_239,N_13661,N_14818);
nor UO_240 (O_240,N_14459,N_14556);
xnor UO_241 (O_241,N_13788,N_14691);
xor UO_242 (O_242,N_14567,N_13891);
or UO_243 (O_243,N_14694,N_13525);
or UO_244 (O_244,N_14982,N_14630);
and UO_245 (O_245,N_14771,N_13742);
or UO_246 (O_246,N_13597,N_13762);
nand UO_247 (O_247,N_13734,N_14928);
nor UO_248 (O_248,N_14615,N_14782);
nor UO_249 (O_249,N_14897,N_14883);
nand UO_250 (O_250,N_14610,N_14326);
nor UO_251 (O_251,N_14083,N_14723);
or UO_252 (O_252,N_14004,N_14485);
or UO_253 (O_253,N_14821,N_14398);
nand UO_254 (O_254,N_14754,N_14632);
or UO_255 (O_255,N_14177,N_14915);
and UO_256 (O_256,N_13733,N_14405);
nor UO_257 (O_257,N_13925,N_13610);
nor UO_258 (O_258,N_14841,N_14979);
and UO_259 (O_259,N_14989,N_13945);
or UO_260 (O_260,N_13703,N_14640);
or UO_261 (O_261,N_14616,N_14757);
or UO_262 (O_262,N_14235,N_14112);
and UO_263 (O_263,N_13949,N_14623);
nor UO_264 (O_264,N_13579,N_14079);
nand UO_265 (O_265,N_14482,N_14406);
nand UO_266 (O_266,N_13785,N_14959);
xnor UO_267 (O_267,N_13965,N_14188);
or UO_268 (O_268,N_14109,N_13774);
nand UO_269 (O_269,N_14057,N_14186);
nor UO_270 (O_270,N_13805,N_14670);
and UO_271 (O_271,N_14807,N_13869);
or UO_272 (O_272,N_13971,N_14454);
or UO_273 (O_273,N_14064,N_13848);
nor UO_274 (O_274,N_13562,N_13757);
or UO_275 (O_275,N_13922,N_14453);
nand UO_276 (O_276,N_14536,N_14553);
and UO_277 (O_277,N_13872,N_14930);
or UO_278 (O_278,N_14561,N_13652);
nor UO_279 (O_279,N_14542,N_13761);
or UO_280 (O_280,N_14124,N_14058);
nand UO_281 (O_281,N_14101,N_14130);
and UO_282 (O_282,N_14144,N_13536);
nor UO_283 (O_283,N_13778,N_14985);
or UO_284 (O_284,N_14651,N_14348);
nand UO_285 (O_285,N_14419,N_13670);
or UO_286 (O_286,N_14261,N_14013);
xnor UO_287 (O_287,N_13628,N_14009);
xnor UO_288 (O_288,N_14806,N_14026);
and UO_289 (O_289,N_13970,N_14592);
or UO_290 (O_290,N_13674,N_13974);
nor UO_291 (O_291,N_13764,N_14662);
and UO_292 (O_292,N_14882,N_14748);
or UO_293 (O_293,N_14775,N_13599);
nand UO_294 (O_294,N_13647,N_14887);
nor UO_295 (O_295,N_14428,N_13878);
and UO_296 (O_296,N_14945,N_13644);
or UO_297 (O_297,N_14817,N_14832);
nor UO_298 (O_298,N_14805,N_14527);
or UO_299 (O_299,N_13969,N_14868);
or UO_300 (O_300,N_13532,N_14295);
nand UO_301 (O_301,N_14502,N_13684);
and UO_302 (O_302,N_13771,N_14480);
and UO_303 (O_303,N_13560,N_14374);
and UO_304 (O_304,N_14560,N_14874);
nand UO_305 (O_305,N_14209,N_14543);
nor UO_306 (O_306,N_14218,N_14772);
and UO_307 (O_307,N_13913,N_13873);
nand UO_308 (O_308,N_14478,N_14695);
nor UO_309 (O_309,N_14168,N_14500);
nand UO_310 (O_310,N_14690,N_14573);
or UO_311 (O_311,N_14840,N_14511);
nor UO_312 (O_312,N_14335,N_14357);
xnor UO_313 (O_313,N_14302,N_14450);
nand UO_314 (O_314,N_13845,N_13966);
nor UO_315 (O_315,N_14565,N_14499);
nand UO_316 (O_316,N_14439,N_14629);
and UO_317 (O_317,N_14201,N_14413);
nor UO_318 (O_318,N_14886,N_14164);
nor UO_319 (O_319,N_14166,N_14855);
nor UO_320 (O_320,N_14860,N_14970);
nand UO_321 (O_321,N_14739,N_13706);
and UO_322 (O_322,N_14460,N_13908);
or UO_323 (O_323,N_14777,N_14826);
and UO_324 (O_324,N_14385,N_13895);
nand UO_325 (O_325,N_14259,N_14437);
nand UO_326 (O_326,N_14776,N_14768);
nor UO_327 (O_327,N_14115,N_14275);
nand UO_328 (O_328,N_14584,N_13992);
or UO_329 (O_329,N_14612,N_14089);
and UO_330 (O_330,N_14368,N_13818);
nand UO_331 (O_331,N_13516,N_14917);
or UO_332 (O_332,N_14781,N_13507);
and UO_333 (O_333,N_14937,N_14919);
nand UO_334 (O_334,N_13800,N_14879);
or UO_335 (O_335,N_14916,N_14896);
and UO_336 (O_336,N_14068,N_14994);
and UO_337 (O_337,N_14149,N_14370);
or UO_338 (O_338,N_13557,N_13576);
nor UO_339 (O_339,N_14680,N_14980);
or UO_340 (O_340,N_14579,N_13747);
xnor UO_341 (O_341,N_14025,N_13654);
or UO_342 (O_342,N_13833,N_14473);
and UO_343 (O_343,N_14733,N_14785);
nand UO_344 (O_344,N_14183,N_14169);
or UO_345 (O_345,N_14053,N_14220);
and UO_346 (O_346,N_14999,N_14044);
and UO_347 (O_347,N_14060,N_13765);
and UO_348 (O_348,N_13808,N_13751);
nand UO_349 (O_349,N_14804,N_14595);
and UO_350 (O_350,N_13787,N_14189);
nor UO_351 (O_351,N_14430,N_13729);
nand UO_352 (O_352,N_14568,N_13600);
and UO_353 (O_353,N_14533,N_14535);
and UO_354 (O_354,N_14069,N_13639);
nor UO_355 (O_355,N_14848,N_14355);
or UO_356 (O_356,N_13720,N_14559);
nand UO_357 (O_357,N_14717,N_14607);
or UO_358 (O_358,N_13780,N_14010);
or UO_359 (O_359,N_14752,N_13947);
nor UO_360 (O_360,N_13954,N_14742);
nor UO_361 (O_361,N_14151,N_14685);
or UO_362 (O_362,N_14353,N_14956);
nor UO_363 (O_363,N_14955,N_14170);
or UO_364 (O_364,N_14663,N_14153);
nor UO_365 (O_365,N_14669,N_14786);
xnor UO_366 (O_366,N_13598,N_14828);
or UO_367 (O_367,N_14300,N_14866);
or UO_368 (O_368,N_14822,N_14137);
and UO_369 (O_369,N_14344,N_14637);
nor UO_370 (O_370,N_13866,N_14747);
and UO_371 (O_371,N_13739,N_14667);
and UO_372 (O_372,N_14376,N_14243);
nor UO_373 (O_373,N_13921,N_14870);
or UO_374 (O_374,N_13986,N_14931);
nor UO_375 (O_375,N_13624,N_13933);
and UO_376 (O_376,N_13641,N_13704);
xor UO_377 (O_377,N_14614,N_14148);
and UO_378 (O_378,N_14712,N_14849);
nor UO_379 (O_379,N_13812,N_13623);
nand UO_380 (O_380,N_14652,N_14940);
or UO_381 (O_381,N_14265,N_13806);
nor UO_382 (O_382,N_14349,N_14343);
nor UO_383 (O_383,N_14954,N_13775);
and UO_384 (O_384,N_13503,N_14107);
xor UO_385 (O_385,N_14342,N_14634);
nand UO_386 (O_386,N_14394,N_13803);
nor UO_387 (O_387,N_14672,N_13944);
nor UO_388 (O_388,N_13642,N_14230);
or UO_389 (O_389,N_13991,N_14461);
or UO_390 (O_390,N_14253,N_14769);
or UO_391 (O_391,N_14572,N_14587);
and UO_392 (O_392,N_13586,N_13687);
or UO_393 (O_393,N_13535,N_13842);
nand UO_394 (O_394,N_13827,N_14534);
nand UO_395 (O_395,N_14283,N_13976);
and UO_396 (O_396,N_13668,N_13512);
and UO_397 (O_397,N_13799,N_14318);
nor UO_398 (O_398,N_14519,N_14395);
nand UO_399 (O_399,N_14347,N_14646);
nand UO_400 (O_400,N_13696,N_14028);
and UO_401 (O_401,N_14557,N_14249);
or UO_402 (O_402,N_13963,N_14046);
and UO_403 (O_403,N_13553,N_13953);
nand UO_404 (O_404,N_14912,N_14323);
and UO_405 (O_405,N_14445,N_14438);
or UO_406 (O_406,N_13882,N_14293);
and UO_407 (O_407,N_13685,N_13940);
or UO_408 (O_408,N_14580,N_14918);
nand UO_409 (O_409,N_14155,N_14350);
or UO_410 (O_410,N_13943,N_14756);
nor UO_411 (O_411,N_14602,N_14909);
and UO_412 (O_412,N_13637,N_14012);
nor UO_413 (O_413,N_13659,N_14707);
or UO_414 (O_414,N_14594,N_13950);
nand UO_415 (O_415,N_13890,N_14092);
nor UO_416 (O_416,N_14961,N_14563);
and UO_417 (O_417,N_13522,N_13691);
nand UO_418 (O_418,N_14721,N_14258);
nor UO_419 (O_419,N_14767,N_14384);
xnor UO_420 (O_420,N_14363,N_13858);
nand UO_421 (O_421,N_14760,N_13951);
or UO_422 (O_422,N_14834,N_14062);
nor UO_423 (O_423,N_13693,N_14910);
or UO_424 (O_424,N_13688,N_13621);
nand UO_425 (O_425,N_13537,N_14337);
and UO_426 (O_426,N_13643,N_13564);
nand UO_427 (O_427,N_13531,N_14319);
nand UO_428 (O_428,N_13715,N_14509);
nor UO_429 (O_429,N_14005,N_14072);
nor UO_430 (O_430,N_14564,N_14328);
nand UO_431 (O_431,N_14159,N_13879);
and UO_432 (O_432,N_14346,N_14393);
xnor UO_433 (O_433,N_13830,N_14974);
and UO_434 (O_434,N_14440,N_14475);
nand UO_435 (O_435,N_13889,N_13655);
or UO_436 (O_436,N_13617,N_14516);
nand UO_437 (O_437,N_14094,N_14038);
or UO_438 (O_438,N_14765,N_14881);
nand UO_439 (O_439,N_14233,N_14716);
nand UO_440 (O_440,N_14653,N_14749);
or UO_441 (O_441,N_14090,N_13500);
or UO_442 (O_442,N_14494,N_14609);
or UO_443 (O_443,N_13509,N_14055);
or UO_444 (O_444,N_14452,N_14065);
and UO_445 (O_445,N_13545,N_13571);
nor UO_446 (O_446,N_14324,N_14490);
and UO_447 (O_447,N_14641,N_13705);
nor UO_448 (O_448,N_14034,N_13517);
nor UO_449 (O_449,N_13732,N_14835);
or UO_450 (O_450,N_14023,N_14093);
and UO_451 (O_451,N_13737,N_14986);
nor UO_452 (O_452,N_14383,N_14853);
nand UO_453 (O_453,N_14816,N_14814);
and UO_454 (O_454,N_14434,N_14278);
nor UO_455 (O_455,N_14436,N_14862);
xnor UO_456 (O_456,N_14843,N_14174);
xnor UO_457 (O_457,N_14024,N_14486);
nor UO_458 (O_458,N_14528,N_14575);
nor UO_459 (O_459,N_14045,N_14618);
nand UO_460 (O_460,N_14279,N_13524);
xor UO_461 (O_461,N_14260,N_13716);
nand UO_462 (O_462,N_13635,N_14416);
or UO_463 (O_463,N_13638,N_14501);
nand UO_464 (O_464,N_13613,N_14409);
nand UO_465 (O_465,N_14958,N_14913);
xor UO_466 (O_466,N_14990,N_13648);
nand UO_467 (O_467,N_14292,N_14116);
nand UO_468 (O_468,N_13838,N_13861);
and UO_469 (O_469,N_13634,N_13700);
nand UO_470 (O_470,N_14192,N_14006);
xor UO_471 (O_471,N_14311,N_14105);
nand UO_472 (O_472,N_13682,N_14225);
or UO_473 (O_473,N_13928,N_14949);
and UO_474 (O_474,N_14304,N_13844);
nand UO_475 (O_475,N_13999,N_14158);
or UO_476 (O_476,N_14626,N_14537);
nand UO_477 (O_477,N_14237,N_14420);
nand UO_478 (O_478,N_14778,N_13669);
or UO_479 (O_479,N_14215,N_14289);
or UO_480 (O_480,N_14784,N_14539);
or UO_481 (O_481,N_14415,N_14294);
nor UO_482 (O_482,N_13618,N_13790);
xor UO_483 (O_483,N_13578,N_14410);
nor UO_484 (O_484,N_13569,N_14933);
or UO_485 (O_485,N_14601,N_13898);
and UO_486 (O_486,N_13677,N_13590);
and UO_487 (O_487,N_14172,N_13606);
or UO_488 (O_488,N_14228,N_13763);
or UO_489 (O_489,N_14208,N_13611);
nand UO_490 (O_490,N_13506,N_14677);
and UO_491 (O_491,N_14016,N_14795);
xor UO_492 (O_492,N_14226,N_13836);
nor UO_493 (O_493,N_14231,N_14085);
nand UO_494 (O_494,N_14426,N_14443);
and UO_495 (O_495,N_14157,N_14589);
and UO_496 (O_496,N_14859,N_14442);
or UO_497 (O_497,N_14715,N_14811);
nor UO_498 (O_498,N_14134,N_13743);
nand UO_499 (O_499,N_13741,N_14078);
nor UO_500 (O_500,N_14203,N_13977);
or UO_501 (O_501,N_14001,N_14703);
and UO_502 (O_502,N_14972,N_14207);
nand UO_503 (O_503,N_14002,N_14441);
nor UO_504 (O_504,N_14330,N_14978);
or UO_505 (O_505,N_13581,N_14934);
or UO_506 (O_506,N_14549,N_14020);
nand UO_507 (O_507,N_14362,N_14360);
nand UO_508 (O_508,N_14070,N_13526);
nand UO_509 (O_509,N_14457,N_14763);
nor UO_510 (O_510,N_13714,N_13807);
nand UO_511 (O_511,N_14697,N_14100);
nand UO_512 (O_512,N_14133,N_14179);
or UO_513 (O_513,N_14656,N_14673);
and UO_514 (O_514,N_14699,N_14182);
nand UO_515 (O_515,N_14074,N_13629);
and UO_516 (O_516,N_14372,N_13679);
nor UO_517 (O_517,N_13804,N_14746);
or UO_518 (O_518,N_13915,N_14507);
or UO_519 (O_519,N_13857,N_13995);
xnor UO_520 (O_520,N_14244,N_14593);
xnor UO_521 (O_521,N_14531,N_13825);
or UO_522 (O_522,N_14948,N_14894);
and UO_523 (O_523,N_13760,N_13768);
xor UO_524 (O_524,N_14135,N_14152);
nand UO_525 (O_525,N_13749,N_14007);
or UO_526 (O_526,N_14103,N_14392);
nand UO_527 (O_527,N_14729,N_13941);
or UO_528 (O_528,N_13686,N_14736);
nor UO_529 (O_529,N_14080,N_14377);
nand UO_530 (O_530,N_13934,N_13905);
or UO_531 (O_531,N_14713,N_14666);
nor UO_532 (O_532,N_14705,N_14050);
and UO_533 (O_533,N_13868,N_14063);
nand UO_534 (O_534,N_14334,N_14809);
xor UO_535 (O_535,N_14451,N_13856);
nand UO_536 (O_536,N_14590,N_14147);
or UO_537 (O_537,N_13538,N_13651);
nor UO_538 (O_538,N_14555,N_14545);
and UO_539 (O_539,N_14566,N_14649);
nand UO_540 (O_540,N_14939,N_13731);
nand UO_541 (O_541,N_13712,N_14973);
or UO_542 (O_542,N_14242,N_14591);
and UO_543 (O_543,N_14250,N_13973);
and UO_544 (O_544,N_14899,N_14929);
or UO_545 (O_545,N_14315,N_14942);
nand UO_546 (O_546,N_13776,N_14037);
nand UO_547 (O_547,N_14387,N_14212);
and UO_548 (O_548,N_14920,N_13772);
nand UO_549 (O_549,N_14864,N_14518);
or UO_550 (O_550,N_14412,N_13847);
or UO_551 (O_551,N_14730,N_14789);
xnor UO_552 (O_552,N_14396,N_14708);
and UO_553 (O_553,N_14975,N_14122);
nand UO_554 (O_554,N_14003,N_14433);
nor UO_555 (O_555,N_13615,N_13523);
or UO_556 (O_556,N_13515,N_14783);
nand UO_557 (O_557,N_13502,N_13666);
or UO_558 (O_558,N_14167,N_14850);
and UO_559 (O_559,N_13730,N_13556);
nor UO_560 (O_560,N_14790,N_13814);
nor UO_561 (O_561,N_14059,N_14317);
nand UO_562 (O_562,N_14194,N_14820);
or UO_563 (O_563,N_14938,N_14902);
nor UO_564 (O_564,N_14162,N_14252);
or UO_565 (O_565,N_13718,N_13612);
and UO_566 (O_566,N_13543,N_14585);
and UO_567 (O_567,N_14546,N_13815);
or UO_568 (O_568,N_13864,N_13572);
or UO_569 (O_569,N_14099,N_14333);
or UO_570 (O_570,N_13592,N_13620);
and UO_571 (O_571,N_13528,N_14306);
or UO_572 (O_572,N_13657,N_14017);
nand UO_573 (O_573,N_14143,N_13631);
nand UO_574 (O_574,N_13596,N_14644);
or UO_575 (O_575,N_13552,N_14432);
and UO_576 (O_576,N_14128,N_13695);
and UO_577 (O_577,N_13547,N_14741);
nand UO_578 (O_578,N_13946,N_14810);
nand UO_579 (O_579,N_14049,N_13798);
nor UO_580 (O_580,N_14627,N_14369);
and UO_581 (O_581,N_14131,N_13574);
and UO_582 (O_582,N_14744,N_13980);
and UO_583 (O_583,N_14903,N_14722);
nand UO_584 (O_584,N_13607,N_14779);
or UO_585 (O_585,N_14030,N_14312);
nor UO_586 (O_586,N_13779,N_14504);
nand UO_587 (O_587,N_14645,N_13885);
or UO_588 (O_588,N_13736,N_14633);
and UO_589 (O_589,N_14217,N_14797);
or UO_590 (O_590,N_14686,N_14755);
nand UO_591 (O_591,N_14831,N_14291);
nor UO_592 (O_592,N_14540,N_14953);
or UO_593 (O_593,N_14532,N_14358);
or UO_594 (O_594,N_13948,N_14725);
nand UO_595 (O_595,N_13961,N_14288);
nor UO_596 (O_596,N_14462,N_14282);
nor UO_597 (O_597,N_14554,N_14758);
nor UO_598 (O_598,N_14270,N_13735);
nor UO_599 (O_599,N_14522,N_14570);
nand UO_600 (O_600,N_14310,N_13619);
or UO_601 (O_601,N_14659,N_14463);
nand UO_602 (O_602,N_14976,N_13608);
nand UO_603 (O_603,N_14205,N_14998);
or UO_604 (O_604,N_13841,N_13759);
nand UO_605 (O_605,N_14720,N_14139);
nand UO_606 (O_606,N_14538,N_14054);
xnor UO_607 (O_607,N_13840,N_13855);
and UO_608 (O_608,N_14603,N_14687);
and UO_609 (O_609,N_14234,N_14196);
and UO_610 (O_610,N_14284,N_13640);
or UO_611 (O_611,N_14248,N_13837);
nor UO_612 (O_612,N_13784,N_14418);
xor UO_613 (O_613,N_13929,N_13681);
and UO_614 (O_614,N_14321,N_14290);
or UO_615 (O_615,N_14608,N_14245);
and UO_616 (O_616,N_14123,N_13555);
or UO_617 (O_617,N_13874,N_13663);
nor UO_618 (O_618,N_14911,N_13508);
or UO_619 (O_619,N_13756,N_14429);
nor UO_620 (O_620,N_13709,N_14386);
nand UO_621 (O_621,N_13550,N_13968);
and UO_622 (O_622,N_14987,N_13534);
and UO_623 (O_623,N_13801,N_13937);
or UO_624 (O_624,N_14966,N_13902);
or UO_625 (O_625,N_14571,N_14520);
nor UO_626 (O_626,N_14947,N_13632);
or UO_627 (O_627,N_13978,N_13916);
nor UO_628 (O_628,N_14481,N_13832);
nand UO_629 (O_629,N_14276,N_14489);
or UO_630 (O_630,N_14219,N_13529);
nor UO_631 (O_631,N_14871,N_14029);
and UO_632 (O_632,N_14643,N_14111);
or UO_633 (O_633,N_14951,N_14905);
and UO_634 (O_634,N_14837,N_14091);
nand UO_635 (O_635,N_14764,N_14257);
or UO_636 (O_636,N_13896,N_14120);
xnor UO_637 (O_637,N_13609,N_13513);
xnor UO_638 (O_638,N_14431,N_14801);
and UO_639 (O_639,N_14380,N_13587);
nand UO_640 (O_640,N_14077,N_14039);
nand UO_641 (O_641,N_14505,N_14706);
xor UO_642 (O_642,N_13834,N_14698);
xor UO_643 (O_643,N_14340,N_14145);
or UO_644 (O_644,N_13777,N_14247);
nor UO_645 (O_645,N_13910,N_14067);
nor UO_646 (O_646,N_14679,N_14399);
or UO_647 (O_647,N_13816,N_13843);
or UO_648 (O_648,N_14696,N_14136);
nor UO_649 (O_649,N_14827,N_13675);
or UO_650 (O_650,N_14142,N_14813);
and UO_651 (O_651,N_13673,N_14688);
and UO_652 (O_652,N_14799,N_13942);
xnor UO_653 (O_653,N_14239,N_14582);
and UO_654 (O_654,N_13520,N_13783);
nand UO_655 (O_655,N_14711,N_14846);
or UO_656 (O_656,N_14236,N_14322);
or UO_657 (O_657,N_14286,N_14015);
or UO_658 (O_658,N_14581,N_14447);
or UO_659 (O_659,N_13822,N_14924);
nand UO_660 (O_660,N_14102,N_13786);
or UO_661 (O_661,N_14750,N_14647);
nand UO_662 (O_662,N_13540,N_13935);
and UO_663 (O_663,N_14548,N_14223);
nand UO_664 (O_664,N_14792,N_14796);
and UO_665 (O_665,N_14944,N_13755);
or UO_666 (O_666,N_13728,N_14856);
and UO_667 (O_667,N_14971,N_14495);
and UO_668 (O_668,N_14229,N_14193);
and UO_669 (O_669,N_14487,N_13984);
and UO_670 (O_670,N_14625,N_13721);
nor UO_671 (O_671,N_14214,N_14878);
nor UO_672 (O_672,N_13546,N_14893);
nand UO_673 (O_673,N_13993,N_13990);
xnor UO_674 (O_674,N_13723,N_13653);
nor UO_675 (O_675,N_14407,N_13725);
and UO_676 (O_676,N_13854,N_14506);
and UO_677 (O_677,N_14578,N_13924);
or UO_678 (O_678,N_14119,N_14709);
xor UO_679 (O_679,N_13544,N_14889);
or UO_680 (O_680,N_14606,N_14577);
xnor UO_681 (O_681,N_14082,N_13987);
xnor UO_682 (O_682,N_14665,N_14066);
xor UO_683 (O_683,N_14574,N_14983);
nor UO_684 (O_684,N_13549,N_13683);
or UO_685 (O_685,N_14622,N_14296);
or UO_686 (O_686,N_14508,N_14977);
and UO_687 (O_687,N_14842,N_14197);
nor UO_688 (O_688,N_14794,N_13707);
nor UO_689 (O_689,N_14515,N_14305);
or UO_690 (O_690,N_13689,N_14906);
and UO_691 (O_691,N_13817,N_14642);
nand UO_692 (O_692,N_14042,N_14914);
and UO_693 (O_693,N_14569,N_14371);
nor UO_694 (O_694,N_14967,N_14621);
or UO_695 (O_695,N_14793,N_13880);
nand UO_696 (O_696,N_14935,N_14423);
nand UO_697 (O_697,N_13656,N_13710);
nor UO_698 (O_698,N_13769,N_13983);
or UO_699 (O_699,N_14676,N_14852);
nand UO_700 (O_700,N_14774,N_14331);
nor UO_701 (O_701,N_13511,N_14484);
and UO_702 (O_702,N_13773,N_14378);
and UO_703 (O_703,N_14867,N_13582);
or UO_704 (O_704,N_14097,N_14216);
or UO_705 (O_705,N_14901,N_13994);
nor UO_706 (O_706,N_14740,N_13697);
or UO_707 (O_707,N_14052,N_13819);
nor UO_708 (O_708,N_14008,N_14018);
or UO_709 (O_709,N_14021,N_14019);
or UO_710 (O_710,N_14308,N_14681);
and UO_711 (O_711,N_14011,N_13724);
nor UO_712 (O_712,N_13588,N_14364);
nor UO_713 (O_713,N_13630,N_13541);
xor UO_714 (O_714,N_13782,N_13622);
and UO_715 (O_715,N_14106,N_13853);
nor UO_716 (O_716,N_14724,N_14351);
xor UO_717 (O_717,N_14435,N_14892);
or UO_718 (O_718,N_14086,N_13565);
xor UO_719 (O_719,N_14851,N_14891);
nor UO_720 (O_720,N_14513,N_14664);
nor UO_721 (O_721,N_13767,N_14875);
or UO_722 (O_722,N_14051,N_14991);
nand UO_723 (O_723,N_14624,N_13781);
nor UO_724 (O_724,N_14098,N_14361);
nand UO_725 (O_725,N_14759,N_13813);
nand UO_726 (O_726,N_14084,N_14047);
or UO_727 (O_727,N_14552,N_13792);
or UO_728 (O_728,N_14339,N_14200);
nand UO_729 (O_729,N_14660,N_14277);
nor UO_730 (O_730,N_14529,N_14611);
or UO_731 (O_731,N_14354,N_13914);
nand UO_732 (O_732,N_14329,N_13645);
nand UO_733 (O_733,N_14425,N_13997);
and UO_734 (O_734,N_14110,N_14414);
and UO_735 (O_735,N_14140,N_13602);
and UO_736 (O_736,N_14314,N_14521);
and UO_737 (O_737,N_14727,N_13846);
nor UO_738 (O_738,N_13989,N_14498);
or UO_739 (O_739,N_13551,N_14732);
nor UO_740 (O_740,N_14156,N_14692);
or UO_741 (O_741,N_13664,N_14325);
nand UO_742 (O_742,N_13920,N_14232);
and UO_743 (O_743,N_14830,N_14146);
or UO_744 (O_744,N_14365,N_14823);
or UO_745 (O_745,N_14465,N_14036);
or UO_746 (O_746,N_13881,N_14726);
and UO_747 (O_747,N_13828,N_14195);
nor UO_748 (O_748,N_13566,N_14702);
or UO_749 (O_749,N_13909,N_13625);
nor UO_750 (O_750,N_13564,N_14279);
nand UO_751 (O_751,N_14432,N_14327);
nor UO_752 (O_752,N_14880,N_14986);
nand UO_753 (O_753,N_14282,N_14655);
nand UO_754 (O_754,N_14745,N_13549);
nand UO_755 (O_755,N_14205,N_13604);
nor UO_756 (O_756,N_14187,N_14577);
nor UO_757 (O_757,N_14306,N_14445);
and UO_758 (O_758,N_14391,N_14628);
and UO_759 (O_759,N_14531,N_13789);
xor UO_760 (O_760,N_14573,N_13742);
nor UO_761 (O_761,N_14986,N_13775);
or UO_762 (O_762,N_14286,N_14571);
or UO_763 (O_763,N_14156,N_14449);
or UO_764 (O_764,N_14028,N_14977);
nor UO_765 (O_765,N_14712,N_14352);
xnor UO_766 (O_766,N_14257,N_14775);
nand UO_767 (O_767,N_14172,N_14597);
nand UO_768 (O_768,N_13937,N_14872);
nor UO_769 (O_769,N_14837,N_14671);
or UO_770 (O_770,N_14480,N_14413);
and UO_771 (O_771,N_14629,N_14080);
xor UO_772 (O_772,N_14076,N_14119);
nor UO_773 (O_773,N_14054,N_14823);
or UO_774 (O_774,N_14436,N_14533);
and UO_775 (O_775,N_14448,N_14729);
nor UO_776 (O_776,N_14474,N_14718);
or UO_777 (O_777,N_13569,N_14658);
or UO_778 (O_778,N_13527,N_14105);
or UO_779 (O_779,N_14971,N_13579);
or UO_780 (O_780,N_13914,N_14233);
nand UO_781 (O_781,N_14569,N_14654);
xor UO_782 (O_782,N_14055,N_14542);
nand UO_783 (O_783,N_13981,N_13907);
xor UO_784 (O_784,N_13770,N_14342);
or UO_785 (O_785,N_14097,N_14368);
and UO_786 (O_786,N_14312,N_14561);
nand UO_787 (O_787,N_14220,N_13747);
nor UO_788 (O_788,N_13989,N_13737);
or UO_789 (O_789,N_13544,N_14579);
and UO_790 (O_790,N_14778,N_14097);
or UO_791 (O_791,N_14767,N_14583);
or UO_792 (O_792,N_13600,N_13759);
nor UO_793 (O_793,N_14208,N_14100);
nor UO_794 (O_794,N_14548,N_13991);
and UO_795 (O_795,N_14375,N_13555);
or UO_796 (O_796,N_13516,N_13649);
nand UO_797 (O_797,N_14857,N_14476);
xnor UO_798 (O_798,N_14957,N_14322);
or UO_799 (O_799,N_14271,N_14600);
nand UO_800 (O_800,N_14273,N_14550);
nor UO_801 (O_801,N_14891,N_13842);
nor UO_802 (O_802,N_14561,N_13848);
nand UO_803 (O_803,N_14594,N_14438);
or UO_804 (O_804,N_14013,N_13656);
or UO_805 (O_805,N_14423,N_14429);
nor UO_806 (O_806,N_14633,N_13541);
nor UO_807 (O_807,N_14146,N_14900);
xnor UO_808 (O_808,N_13594,N_14256);
or UO_809 (O_809,N_14643,N_13914);
nand UO_810 (O_810,N_14328,N_13595);
and UO_811 (O_811,N_14511,N_14367);
and UO_812 (O_812,N_13607,N_14632);
nor UO_813 (O_813,N_14571,N_14502);
or UO_814 (O_814,N_14905,N_13877);
or UO_815 (O_815,N_14593,N_14501);
nor UO_816 (O_816,N_14350,N_14137);
or UO_817 (O_817,N_14512,N_13765);
or UO_818 (O_818,N_14446,N_14397);
and UO_819 (O_819,N_14046,N_14887);
nor UO_820 (O_820,N_14762,N_14026);
nor UO_821 (O_821,N_14930,N_14228);
or UO_822 (O_822,N_14432,N_14653);
or UO_823 (O_823,N_14434,N_14899);
nand UO_824 (O_824,N_13639,N_13851);
nor UO_825 (O_825,N_14816,N_14144);
nand UO_826 (O_826,N_14207,N_13961);
nand UO_827 (O_827,N_14368,N_14197);
xnor UO_828 (O_828,N_14176,N_14690);
and UO_829 (O_829,N_13887,N_13541);
or UO_830 (O_830,N_13704,N_14209);
nor UO_831 (O_831,N_14137,N_14767);
or UO_832 (O_832,N_14469,N_14658);
nor UO_833 (O_833,N_13565,N_14432);
nand UO_834 (O_834,N_14074,N_13860);
and UO_835 (O_835,N_13849,N_14000);
or UO_836 (O_836,N_13785,N_14329);
and UO_837 (O_837,N_13685,N_14470);
nand UO_838 (O_838,N_14337,N_13875);
nand UO_839 (O_839,N_14298,N_14822);
nand UO_840 (O_840,N_13998,N_14697);
xnor UO_841 (O_841,N_14409,N_14591);
nand UO_842 (O_842,N_13996,N_13791);
nand UO_843 (O_843,N_14102,N_14113);
or UO_844 (O_844,N_14229,N_13792);
and UO_845 (O_845,N_14947,N_14089);
or UO_846 (O_846,N_14299,N_14104);
or UO_847 (O_847,N_14685,N_13794);
nand UO_848 (O_848,N_14194,N_14515);
nand UO_849 (O_849,N_14720,N_14540);
or UO_850 (O_850,N_13888,N_14463);
nor UO_851 (O_851,N_14959,N_14697);
and UO_852 (O_852,N_14722,N_13877);
nor UO_853 (O_853,N_14891,N_14513);
and UO_854 (O_854,N_14368,N_14786);
or UO_855 (O_855,N_14266,N_14647);
nor UO_856 (O_856,N_14796,N_14013);
and UO_857 (O_857,N_14023,N_13944);
nand UO_858 (O_858,N_14174,N_13675);
nand UO_859 (O_859,N_14105,N_14931);
or UO_860 (O_860,N_14430,N_14566);
or UO_861 (O_861,N_14794,N_14538);
nand UO_862 (O_862,N_13772,N_14451);
or UO_863 (O_863,N_14134,N_14214);
xnor UO_864 (O_864,N_13504,N_14356);
and UO_865 (O_865,N_14345,N_14358);
nor UO_866 (O_866,N_14004,N_14864);
nor UO_867 (O_867,N_13579,N_13517);
nor UO_868 (O_868,N_13547,N_14144);
and UO_869 (O_869,N_14958,N_14886);
nor UO_870 (O_870,N_14784,N_14338);
or UO_871 (O_871,N_13602,N_13844);
nand UO_872 (O_872,N_14799,N_14679);
nor UO_873 (O_873,N_13716,N_14020);
and UO_874 (O_874,N_13702,N_13690);
or UO_875 (O_875,N_14894,N_14579);
nor UO_876 (O_876,N_13971,N_13626);
nor UO_877 (O_877,N_14019,N_13981);
nor UO_878 (O_878,N_14457,N_14268);
xnor UO_879 (O_879,N_14144,N_13816);
or UO_880 (O_880,N_14565,N_14177);
nand UO_881 (O_881,N_14829,N_14412);
nor UO_882 (O_882,N_14872,N_13961);
xnor UO_883 (O_883,N_13773,N_14828);
and UO_884 (O_884,N_14532,N_14555);
nand UO_885 (O_885,N_14773,N_14989);
nor UO_886 (O_886,N_14932,N_14595);
nor UO_887 (O_887,N_13965,N_14121);
or UO_888 (O_888,N_14424,N_14206);
and UO_889 (O_889,N_14269,N_14575);
nor UO_890 (O_890,N_14869,N_14683);
and UO_891 (O_891,N_14241,N_13850);
nor UO_892 (O_892,N_13701,N_14835);
nor UO_893 (O_893,N_14013,N_13674);
nor UO_894 (O_894,N_13647,N_13512);
nor UO_895 (O_895,N_14247,N_14294);
and UO_896 (O_896,N_13960,N_14911);
nor UO_897 (O_897,N_14877,N_14296);
nor UO_898 (O_898,N_14329,N_14855);
nor UO_899 (O_899,N_14355,N_13561);
or UO_900 (O_900,N_13522,N_14620);
xnor UO_901 (O_901,N_14805,N_14432);
and UO_902 (O_902,N_13582,N_13831);
and UO_903 (O_903,N_14320,N_13854);
nand UO_904 (O_904,N_14617,N_14289);
and UO_905 (O_905,N_14251,N_13657);
and UO_906 (O_906,N_14511,N_13632);
or UO_907 (O_907,N_14475,N_14915);
or UO_908 (O_908,N_14436,N_14800);
and UO_909 (O_909,N_14325,N_13507);
xnor UO_910 (O_910,N_13845,N_14236);
or UO_911 (O_911,N_14203,N_13539);
or UO_912 (O_912,N_13510,N_13810);
or UO_913 (O_913,N_14747,N_14542);
nand UO_914 (O_914,N_14141,N_14436);
nor UO_915 (O_915,N_13527,N_14230);
and UO_916 (O_916,N_13545,N_14163);
and UO_917 (O_917,N_13905,N_13818);
and UO_918 (O_918,N_13917,N_13500);
nand UO_919 (O_919,N_14822,N_14926);
nor UO_920 (O_920,N_14708,N_14266);
nor UO_921 (O_921,N_14491,N_14798);
nand UO_922 (O_922,N_13807,N_14458);
and UO_923 (O_923,N_14540,N_14821);
and UO_924 (O_924,N_13616,N_14349);
or UO_925 (O_925,N_13969,N_14918);
nand UO_926 (O_926,N_14518,N_14011);
or UO_927 (O_927,N_14527,N_14815);
nor UO_928 (O_928,N_13980,N_13765);
or UO_929 (O_929,N_13635,N_13873);
nand UO_930 (O_930,N_14766,N_14434);
and UO_931 (O_931,N_14032,N_14013);
or UO_932 (O_932,N_14622,N_14060);
or UO_933 (O_933,N_14972,N_13691);
or UO_934 (O_934,N_14106,N_13542);
and UO_935 (O_935,N_14482,N_14584);
nor UO_936 (O_936,N_13842,N_14921);
or UO_937 (O_937,N_13799,N_14791);
and UO_938 (O_938,N_14867,N_14125);
nor UO_939 (O_939,N_13830,N_14778);
nand UO_940 (O_940,N_14603,N_13933);
xnor UO_941 (O_941,N_14230,N_14636);
nand UO_942 (O_942,N_14341,N_14957);
xor UO_943 (O_943,N_13765,N_13532);
xor UO_944 (O_944,N_13788,N_14501);
nand UO_945 (O_945,N_14236,N_13859);
or UO_946 (O_946,N_14139,N_14548);
nand UO_947 (O_947,N_14420,N_14188);
nand UO_948 (O_948,N_14416,N_13816);
or UO_949 (O_949,N_14232,N_14838);
or UO_950 (O_950,N_14921,N_14257);
or UO_951 (O_951,N_13691,N_14136);
xnor UO_952 (O_952,N_14346,N_14818);
and UO_953 (O_953,N_14762,N_13692);
nor UO_954 (O_954,N_13512,N_13640);
nand UO_955 (O_955,N_14706,N_13700);
or UO_956 (O_956,N_14289,N_13796);
nor UO_957 (O_957,N_14625,N_14493);
or UO_958 (O_958,N_14211,N_14592);
nand UO_959 (O_959,N_13654,N_14853);
and UO_960 (O_960,N_14448,N_14548);
nand UO_961 (O_961,N_13850,N_13951);
and UO_962 (O_962,N_14987,N_14393);
nor UO_963 (O_963,N_13916,N_14987);
xnor UO_964 (O_964,N_14435,N_13793);
nand UO_965 (O_965,N_14397,N_14023);
or UO_966 (O_966,N_14229,N_14719);
nand UO_967 (O_967,N_13618,N_14917);
and UO_968 (O_968,N_14640,N_13836);
or UO_969 (O_969,N_14031,N_14042);
or UO_970 (O_970,N_13744,N_14339);
nor UO_971 (O_971,N_14053,N_14575);
nand UO_972 (O_972,N_14029,N_14016);
nand UO_973 (O_973,N_13557,N_14358);
or UO_974 (O_974,N_14659,N_14004);
and UO_975 (O_975,N_14042,N_14110);
nor UO_976 (O_976,N_14840,N_14739);
nor UO_977 (O_977,N_14898,N_13727);
xnor UO_978 (O_978,N_13737,N_13869);
nor UO_979 (O_979,N_14462,N_13674);
or UO_980 (O_980,N_14698,N_13721);
or UO_981 (O_981,N_14882,N_14870);
xor UO_982 (O_982,N_14785,N_14984);
xor UO_983 (O_983,N_14795,N_14631);
and UO_984 (O_984,N_14493,N_13535);
nand UO_985 (O_985,N_13937,N_13685);
or UO_986 (O_986,N_14038,N_14410);
nand UO_987 (O_987,N_14287,N_13943);
xor UO_988 (O_988,N_14095,N_14591);
xor UO_989 (O_989,N_14991,N_14596);
or UO_990 (O_990,N_14899,N_14970);
nor UO_991 (O_991,N_14608,N_14558);
nor UO_992 (O_992,N_14915,N_14749);
and UO_993 (O_993,N_14528,N_13693);
or UO_994 (O_994,N_14985,N_14632);
nand UO_995 (O_995,N_14967,N_14553);
nand UO_996 (O_996,N_13854,N_13989);
and UO_997 (O_997,N_14968,N_14134);
nor UO_998 (O_998,N_14621,N_14578);
and UO_999 (O_999,N_14351,N_14278);
nor UO_1000 (O_1000,N_13916,N_14873);
nand UO_1001 (O_1001,N_14603,N_13777);
or UO_1002 (O_1002,N_14678,N_13955);
nand UO_1003 (O_1003,N_13696,N_13624);
or UO_1004 (O_1004,N_13814,N_14884);
nor UO_1005 (O_1005,N_14305,N_13846);
or UO_1006 (O_1006,N_14605,N_14040);
or UO_1007 (O_1007,N_13796,N_14986);
xnor UO_1008 (O_1008,N_14630,N_14489);
nand UO_1009 (O_1009,N_14193,N_13645);
nand UO_1010 (O_1010,N_13802,N_13546);
or UO_1011 (O_1011,N_14872,N_13532);
or UO_1012 (O_1012,N_13733,N_13930);
nor UO_1013 (O_1013,N_14519,N_13984);
nor UO_1014 (O_1014,N_13829,N_14829);
and UO_1015 (O_1015,N_14195,N_14118);
nor UO_1016 (O_1016,N_14229,N_13651);
and UO_1017 (O_1017,N_14370,N_14331);
or UO_1018 (O_1018,N_14325,N_14403);
or UO_1019 (O_1019,N_14846,N_14320);
nand UO_1020 (O_1020,N_14724,N_13693);
and UO_1021 (O_1021,N_14005,N_13925);
nand UO_1022 (O_1022,N_14050,N_14640);
xnor UO_1023 (O_1023,N_14432,N_14910);
xnor UO_1024 (O_1024,N_13887,N_14021);
nor UO_1025 (O_1025,N_14036,N_14959);
and UO_1026 (O_1026,N_14121,N_14557);
and UO_1027 (O_1027,N_14829,N_13560);
nand UO_1028 (O_1028,N_14591,N_14325);
and UO_1029 (O_1029,N_14020,N_14171);
and UO_1030 (O_1030,N_14696,N_14486);
or UO_1031 (O_1031,N_14207,N_13981);
xor UO_1032 (O_1032,N_14750,N_14517);
xnor UO_1033 (O_1033,N_13878,N_13911);
nand UO_1034 (O_1034,N_14508,N_13933);
nand UO_1035 (O_1035,N_14419,N_14088);
nor UO_1036 (O_1036,N_14902,N_14211);
and UO_1037 (O_1037,N_13534,N_14069);
nor UO_1038 (O_1038,N_14440,N_14719);
xor UO_1039 (O_1039,N_14065,N_13580);
nor UO_1040 (O_1040,N_14981,N_14709);
nor UO_1041 (O_1041,N_14338,N_14262);
nand UO_1042 (O_1042,N_14198,N_13542);
xor UO_1043 (O_1043,N_14042,N_13826);
nor UO_1044 (O_1044,N_14798,N_13568);
nand UO_1045 (O_1045,N_13899,N_13615);
xnor UO_1046 (O_1046,N_14620,N_14655);
or UO_1047 (O_1047,N_14748,N_14886);
nand UO_1048 (O_1048,N_14643,N_14871);
xnor UO_1049 (O_1049,N_14080,N_14405);
and UO_1050 (O_1050,N_14796,N_13572);
nand UO_1051 (O_1051,N_14989,N_14907);
and UO_1052 (O_1052,N_14385,N_14709);
nand UO_1053 (O_1053,N_13572,N_14370);
and UO_1054 (O_1054,N_13665,N_13972);
and UO_1055 (O_1055,N_14961,N_13966);
and UO_1056 (O_1056,N_14076,N_13649);
and UO_1057 (O_1057,N_14943,N_13991);
or UO_1058 (O_1058,N_14902,N_14426);
and UO_1059 (O_1059,N_14704,N_14328);
nand UO_1060 (O_1060,N_13814,N_14725);
or UO_1061 (O_1061,N_13639,N_13722);
nand UO_1062 (O_1062,N_13683,N_14702);
or UO_1063 (O_1063,N_13801,N_14566);
and UO_1064 (O_1064,N_14469,N_14173);
nand UO_1065 (O_1065,N_13572,N_13727);
nor UO_1066 (O_1066,N_13814,N_14651);
nor UO_1067 (O_1067,N_14603,N_14231);
nor UO_1068 (O_1068,N_13827,N_14110);
and UO_1069 (O_1069,N_13858,N_14342);
and UO_1070 (O_1070,N_14045,N_14641);
or UO_1071 (O_1071,N_13958,N_14429);
nand UO_1072 (O_1072,N_14628,N_14704);
and UO_1073 (O_1073,N_14872,N_14762);
or UO_1074 (O_1074,N_14687,N_13670);
and UO_1075 (O_1075,N_14996,N_14642);
or UO_1076 (O_1076,N_14830,N_14870);
nand UO_1077 (O_1077,N_14060,N_14504);
or UO_1078 (O_1078,N_14654,N_14647);
nand UO_1079 (O_1079,N_14371,N_14276);
nand UO_1080 (O_1080,N_14695,N_14562);
nand UO_1081 (O_1081,N_14655,N_14201);
or UO_1082 (O_1082,N_13559,N_13949);
and UO_1083 (O_1083,N_14856,N_13578);
nor UO_1084 (O_1084,N_14389,N_13804);
xnor UO_1085 (O_1085,N_14535,N_14390);
and UO_1086 (O_1086,N_14015,N_13559);
or UO_1087 (O_1087,N_13760,N_13981);
and UO_1088 (O_1088,N_14395,N_13856);
and UO_1089 (O_1089,N_14049,N_14404);
or UO_1090 (O_1090,N_13556,N_14208);
or UO_1091 (O_1091,N_14144,N_14708);
nor UO_1092 (O_1092,N_14366,N_14671);
or UO_1093 (O_1093,N_13714,N_14628);
or UO_1094 (O_1094,N_13792,N_14674);
or UO_1095 (O_1095,N_14139,N_14688);
or UO_1096 (O_1096,N_14748,N_13609);
and UO_1097 (O_1097,N_13505,N_14572);
nor UO_1098 (O_1098,N_14762,N_14686);
and UO_1099 (O_1099,N_14517,N_14010);
and UO_1100 (O_1100,N_14779,N_14381);
xor UO_1101 (O_1101,N_14608,N_13820);
xnor UO_1102 (O_1102,N_13558,N_13798);
nand UO_1103 (O_1103,N_14543,N_14568);
nand UO_1104 (O_1104,N_14012,N_14799);
xor UO_1105 (O_1105,N_14365,N_14133);
or UO_1106 (O_1106,N_14648,N_14101);
and UO_1107 (O_1107,N_14012,N_14789);
nor UO_1108 (O_1108,N_14497,N_13958);
nand UO_1109 (O_1109,N_13630,N_13884);
nor UO_1110 (O_1110,N_13808,N_14999);
nor UO_1111 (O_1111,N_14052,N_14014);
nand UO_1112 (O_1112,N_14927,N_13571);
xnor UO_1113 (O_1113,N_14533,N_13909);
and UO_1114 (O_1114,N_14118,N_14965);
nor UO_1115 (O_1115,N_14172,N_14970);
and UO_1116 (O_1116,N_14375,N_13900);
or UO_1117 (O_1117,N_14917,N_14373);
and UO_1118 (O_1118,N_14492,N_13780);
or UO_1119 (O_1119,N_14453,N_14440);
or UO_1120 (O_1120,N_14714,N_13674);
nor UO_1121 (O_1121,N_14204,N_14474);
xnor UO_1122 (O_1122,N_13981,N_13589);
nor UO_1123 (O_1123,N_14976,N_14478);
nand UO_1124 (O_1124,N_14427,N_14744);
nand UO_1125 (O_1125,N_13761,N_13915);
and UO_1126 (O_1126,N_14595,N_14446);
xnor UO_1127 (O_1127,N_14023,N_13768);
nand UO_1128 (O_1128,N_14483,N_14503);
and UO_1129 (O_1129,N_14150,N_13594);
and UO_1130 (O_1130,N_14035,N_13550);
nor UO_1131 (O_1131,N_13682,N_14078);
nor UO_1132 (O_1132,N_14533,N_14995);
and UO_1133 (O_1133,N_14337,N_14738);
nor UO_1134 (O_1134,N_13701,N_14087);
nand UO_1135 (O_1135,N_14232,N_14640);
nor UO_1136 (O_1136,N_13971,N_13682);
xor UO_1137 (O_1137,N_14757,N_14024);
or UO_1138 (O_1138,N_14075,N_14326);
xor UO_1139 (O_1139,N_13809,N_14688);
and UO_1140 (O_1140,N_13799,N_14676);
or UO_1141 (O_1141,N_13683,N_14126);
nor UO_1142 (O_1142,N_14982,N_14656);
or UO_1143 (O_1143,N_13826,N_13656);
nor UO_1144 (O_1144,N_13932,N_14722);
nand UO_1145 (O_1145,N_13501,N_14128);
nand UO_1146 (O_1146,N_14412,N_14825);
nand UO_1147 (O_1147,N_14445,N_14700);
or UO_1148 (O_1148,N_14129,N_14684);
or UO_1149 (O_1149,N_13778,N_14980);
nand UO_1150 (O_1150,N_14921,N_14704);
nand UO_1151 (O_1151,N_14092,N_14094);
and UO_1152 (O_1152,N_14910,N_14638);
nor UO_1153 (O_1153,N_13793,N_14176);
or UO_1154 (O_1154,N_13852,N_14994);
nor UO_1155 (O_1155,N_14262,N_13848);
nor UO_1156 (O_1156,N_13723,N_14492);
nor UO_1157 (O_1157,N_14850,N_13840);
xor UO_1158 (O_1158,N_13517,N_14274);
nand UO_1159 (O_1159,N_14429,N_14572);
or UO_1160 (O_1160,N_14947,N_14268);
nand UO_1161 (O_1161,N_14214,N_14342);
or UO_1162 (O_1162,N_13884,N_13638);
xor UO_1163 (O_1163,N_13964,N_14264);
and UO_1164 (O_1164,N_13672,N_14045);
nand UO_1165 (O_1165,N_13501,N_14407);
or UO_1166 (O_1166,N_14089,N_13623);
or UO_1167 (O_1167,N_14041,N_14884);
and UO_1168 (O_1168,N_14035,N_13696);
nor UO_1169 (O_1169,N_14366,N_13579);
and UO_1170 (O_1170,N_14688,N_14727);
or UO_1171 (O_1171,N_13617,N_14874);
nand UO_1172 (O_1172,N_14719,N_14883);
and UO_1173 (O_1173,N_13794,N_13545);
or UO_1174 (O_1174,N_14301,N_14351);
or UO_1175 (O_1175,N_14817,N_14098);
nand UO_1176 (O_1176,N_13732,N_14648);
or UO_1177 (O_1177,N_13670,N_14821);
and UO_1178 (O_1178,N_14832,N_14236);
nor UO_1179 (O_1179,N_14006,N_13862);
nand UO_1180 (O_1180,N_13775,N_14544);
nand UO_1181 (O_1181,N_14204,N_13729);
nand UO_1182 (O_1182,N_14224,N_14434);
nor UO_1183 (O_1183,N_14811,N_13527);
or UO_1184 (O_1184,N_14415,N_14620);
and UO_1185 (O_1185,N_14442,N_13970);
and UO_1186 (O_1186,N_14126,N_14772);
nand UO_1187 (O_1187,N_14673,N_13658);
nand UO_1188 (O_1188,N_14919,N_14794);
xor UO_1189 (O_1189,N_14401,N_13970);
nor UO_1190 (O_1190,N_13688,N_14222);
or UO_1191 (O_1191,N_14942,N_14588);
nand UO_1192 (O_1192,N_14405,N_13806);
or UO_1193 (O_1193,N_13832,N_14863);
or UO_1194 (O_1194,N_13902,N_14001);
or UO_1195 (O_1195,N_14889,N_14758);
and UO_1196 (O_1196,N_14003,N_14629);
nand UO_1197 (O_1197,N_13977,N_14429);
and UO_1198 (O_1198,N_14806,N_14085);
or UO_1199 (O_1199,N_13636,N_13509);
nor UO_1200 (O_1200,N_14947,N_14229);
nor UO_1201 (O_1201,N_14497,N_13568);
or UO_1202 (O_1202,N_14669,N_14133);
nand UO_1203 (O_1203,N_14197,N_13871);
nor UO_1204 (O_1204,N_14120,N_13931);
or UO_1205 (O_1205,N_14646,N_14238);
nand UO_1206 (O_1206,N_13988,N_13994);
or UO_1207 (O_1207,N_14871,N_14053);
nand UO_1208 (O_1208,N_14987,N_14824);
and UO_1209 (O_1209,N_13613,N_13691);
or UO_1210 (O_1210,N_13699,N_13802);
or UO_1211 (O_1211,N_14967,N_14966);
or UO_1212 (O_1212,N_14778,N_14574);
nand UO_1213 (O_1213,N_13806,N_14899);
nand UO_1214 (O_1214,N_14749,N_14545);
and UO_1215 (O_1215,N_14880,N_14185);
or UO_1216 (O_1216,N_14385,N_13992);
and UO_1217 (O_1217,N_13687,N_14547);
and UO_1218 (O_1218,N_14935,N_14963);
and UO_1219 (O_1219,N_14996,N_14244);
nor UO_1220 (O_1220,N_13921,N_13570);
and UO_1221 (O_1221,N_14250,N_13500);
nand UO_1222 (O_1222,N_14092,N_13646);
nand UO_1223 (O_1223,N_13922,N_14423);
or UO_1224 (O_1224,N_13924,N_14537);
nor UO_1225 (O_1225,N_14520,N_13692);
and UO_1226 (O_1226,N_14123,N_14399);
nand UO_1227 (O_1227,N_13655,N_14025);
and UO_1228 (O_1228,N_13565,N_13929);
and UO_1229 (O_1229,N_14202,N_13963);
nand UO_1230 (O_1230,N_13663,N_13579);
nor UO_1231 (O_1231,N_14781,N_14337);
nand UO_1232 (O_1232,N_13574,N_14423);
nand UO_1233 (O_1233,N_13588,N_13626);
and UO_1234 (O_1234,N_14539,N_13564);
and UO_1235 (O_1235,N_14916,N_13547);
or UO_1236 (O_1236,N_13886,N_13743);
or UO_1237 (O_1237,N_14377,N_14761);
xnor UO_1238 (O_1238,N_14243,N_13789);
nor UO_1239 (O_1239,N_14899,N_13876);
or UO_1240 (O_1240,N_13731,N_14871);
nand UO_1241 (O_1241,N_13769,N_14331);
and UO_1242 (O_1242,N_14549,N_14292);
nand UO_1243 (O_1243,N_14708,N_14883);
and UO_1244 (O_1244,N_13957,N_13744);
or UO_1245 (O_1245,N_14823,N_14282);
or UO_1246 (O_1246,N_14086,N_13869);
and UO_1247 (O_1247,N_14438,N_14526);
nor UO_1248 (O_1248,N_14547,N_14271);
or UO_1249 (O_1249,N_14313,N_14856);
nor UO_1250 (O_1250,N_14303,N_14338);
xor UO_1251 (O_1251,N_14472,N_13553);
or UO_1252 (O_1252,N_14571,N_14063);
xor UO_1253 (O_1253,N_14470,N_14226);
and UO_1254 (O_1254,N_14475,N_14369);
or UO_1255 (O_1255,N_13563,N_14135);
or UO_1256 (O_1256,N_13934,N_14263);
or UO_1257 (O_1257,N_13915,N_14777);
nand UO_1258 (O_1258,N_14713,N_13671);
nor UO_1259 (O_1259,N_14656,N_14310);
and UO_1260 (O_1260,N_14059,N_14192);
or UO_1261 (O_1261,N_13797,N_14886);
nand UO_1262 (O_1262,N_14619,N_13656);
or UO_1263 (O_1263,N_13879,N_13997);
nand UO_1264 (O_1264,N_14737,N_13927);
or UO_1265 (O_1265,N_13664,N_14813);
nor UO_1266 (O_1266,N_13724,N_14439);
and UO_1267 (O_1267,N_13621,N_14498);
nor UO_1268 (O_1268,N_14158,N_13803);
nand UO_1269 (O_1269,N_14992,N_13972);
or UO_1270 (O_1270,N_14470,N_14300);
or UO_1271 (O_1271,N_14226,N_14436);
or UO_1272 (O_1272,N_14301,N_14438);
nand UO_1273 (O_1273,N_14060,N_14597);
xnor UO_1274 (O_1274,N_13731,N_14334);
nor UO_1275 (O_1275,N_14141,N_14903);
nor UO_1276 (O_1276,N_13907,N_13535);
nor UO_1277 (O_1277,N_13525,N_14869);
and UO_1278 (O_1278,N_13767,N_14352);
nand UO_1279 (O_1279,N_13648,N_13764);
xor UO_1280 (O_1280,N_14018,N_14471);
nor UO_1281 (O_1281,N_14909,N_13879);
or UO_1282 (O_1282,N_13606,N_14169);
nand UO_1283 (O_1283,N_14911,N_13873);
or UO_1284 (O_1284,N_14023,N_13760);
or UO_1285 (O_1285,N_14676,N_14233);
or UO_1286 (O_1286,N_14965,N_13919);
or UO_1287 (O_1287,N_14033,N_13524);
and UO_1288 (O_1288,N_13898,N_14900);
nand UO_1289 (O_1289,N_13601,N_13610);
nand UO_1290 (O_1290,N_14609,N_13876);
nand UO_1291 (O_1291,N_13965,N_13737);
xor UO_1292 (O_1292,N_13989,N_13902);
and UO_1293 (O_1293,N_14454,N_14611);
nor UO_1294 (O_1294,N_13896,N_13686);
nor UO_1295 (O_1295,N_14127,N_13899);
nor UO_1296 (O_1296,N_14190,N_13716);
nand UO_1297 (O_1297,N_13825,N_14326);
nand UO_1298 (O_1298,N_13871,N_14509);
nor UO_1299 (O_1299,N_14753,N_13834);
or UO_1300 (O_1300,N_13859,N_14355);
and UO_1301 (O_1301,N_13656,N_14825);
xor UO_1302 (O_1302,N_14490,N_13564);
nand UO_1303 (O_1303,N_14244,N_13830);
nand UO_1304 (O_1304,N_14022,N_14998);
nand UO_1305 (O_1305,N_14300,N_14976);
or UO_1306 (O_1306,N_14208,N_14528);
and UO_1307 (O_1307,N_14451,N_13602);
xnor UO_1308 (O_1308,N_14587,N_14963);
nor UO_1309 (O_1309,N_14922,N_14913);
nor UO_1310 (O_1310,N_13531,N_14486);
nand UO_1311 (O_1311,N_14819,N_13934);
nand UO_1312 (O_1312,N_13780,N_13867);
or UO_1313 (O_1313,N_14823,N_14338);
or UO_1314 (O_1314,N_14359,N_14322);
or UO_1315 (O_1315,N_14009,N_13934);
and UO_1316 (O_1316,N_14432,N_14590);
and UO_1317 (O_1317,N_13544,N_14789);
or UO_1318 (O_1318,N_14012,N_13603);
nor UO_1319 (O_1319,N_14677,N_14599);
and UO_1320 (O_1320,N_14012,N_13690);
and UO_1321 (O_1321,N_14353,N_14677);
and UO_1322 (O_1322,N_13626,N_13540);
nor UO_1323 (O_1323,N_14560,N_14047);
or UO_1324 (O_1324,N_14787,N_14945);
or UO_1325 (O_1325,N_14705,N_14998);
nand UO_1326 (O_1326,N_13982,N_14932);
nor UO_1327 (O_1327,N_14101,N_14974);
nand UO_1328 (O_1328,N_14002,N_14088);
and UO_1329 (O_1329,N_14149,N_14107);
nand UO_1330 (O_1330,N_14296,N_14589);
or UO_1331 (O_1331,N_14813,N_13586);
or UO_1332 (O_1332,N_14637,N_14591);
xor UO_1333 (O_1333,N_14873,N_14392);
or UO_1334 (O_1334,N_14710,N_14217);
or UO_1335 (O_1335,N_14223,N_14282);
nand UO_1336 (O_1336,N_14431,N_14926);
and UO_1337 (O_1337,N_13667,N_14151);
and UO_1338 (O_1338,N_14978,N_14756);
nand UO_1339 (O_1339,N_14236,N_14184);
xor UO_1340 (O_1340,N_14704,N_14427);
and UO_1341 (O_1341,N_13840,N_14639);
or UO_1342 (O_1342,N_14924,N_13726);
nor UO_1343 (O_1343,N_14768,N_13872);
and UO_1344 (O_1344,N_14829,N_13994);
nand UO_1345 (O_1345,N_13886,N_13504);
nor UO_1346 (O_1346,N_14805,N_14458);
or UO_1347 (O_1347,N_14577,N_14902);
nand UO_1348 (O_1348,N_14514,N_13560);
nor UO_1349 (O_1349,N_13908,N_13709);
and UO_1350 (O_1350,N_13875,N_14873);
or UO_1351 (O_1351,N_14580,N_13678);
xnor UO_1352 (O_1352,N_13953,N_13535);
nand UO_1353 (O_1353,N_13988,N_13974);
nand UO_1354 (O_1354,N_13716,N_14951);
nor UO_1355 (O_1355,N_14276,N_14046);
nor UO_1356 (O_1356,N_13978,N_14487);
nand UO_1357 (O_1357,N_13687,N_14640);
nor UO_1358 (O_1358,N_14277,N_13877);
nor UO_1359 (O_1359,N_14079,N_14017);
nand UO_1360 (O_1360,N_13687,N_14226);
nand UO_1361 (O_1361,N_14444,N_14603);
nand UO_1362 (O_1362,N_14557,N_13803);
or UO_1363 (O_1363,N_14312,N_14000);
or UO_1364 (O_1364,N_13979,N_14176);
nand UO_1365 (O_1365,N_14437,N_14507);
and UO_1366 (O_1366,N_13523,N_14118);
nand UO_1367 (O_1367,N_13551,N_13843);
nand UO_1368 (O_1368,N_13834,N_13619);
nand UO_1369 (O_1369,N_13928,N_14749);
and UO_1370 (O_1370,N_14112,N_13666);
nand UO_1371 (O_1371,N_14421,N_14287);
and UO_1372 (O_1372,N_14412,N_14665);
nor UO_1373 (O_1373,N_14833,N_14775);
and UO_1374 (O_1374,N_14724,N_14827);
or UO_1375 (O_1375,N_14853,N_14400);
and UO_1376 (O_1376,N_13559,N_13931);
and UO_1377 (O_1377,N_13996,N_14715);
nor UO_1378 (O_1378,N_13562,N_13582);
nand UO_1379 (O_1379,N_14500,N_13751);
and UO_1380 (O_1380,N_14311,N_13587);
or UO_1381 (O_1381,N_13830,N_14649);
nor UO_1382 (O_1382,N_14841,N_14831);
nor UO_1383 (O_1383,N_14794,N_13664);
or UO_1384 (O_1384,N_14144,N_13988);
and UO_1385 (O_1385,N_13736,N_13920);
and UO_1386 (O_1386,N_13927,N_14122);
nor UO_1387 (O_1387,N_14758,N_14365);
and UO_1388 (O_1388,N_13505,N_14687);
or UO_1389 (O_1389,N_14622,N_14951);
or UO_1390 (O_1390,N_14649,N_14739);
nand UO_1391 (O_1391,N_13677,N_14409);
nor UO_1392 (O_1392,N_14208,N_14355);
nor UO_1393 (O_1393,N_14808,N_14587);
xor UO_1394 (O_1394,N_14791,N_13781);
xnor UO_1395 (O_1395,N_14542,N_14720);
nand UO_1396 (O_1396,N_14820,N_14772);
nor UO_1397 (O_1397,N_14614,N_13931);
nor UO_1398 (O_1398,N_13859,N_14376);
and UO_1399 (O_1399,N_14779,N_14925);
nand UO_1400 (O_1400,N_14583,N_14077);
and UO_1401 (O_1401,N_14472,N_14927);
nand UO_1402 (O_1402,N_14431,N_14406);
nor UO_1403 (O_1403,N_14757,N_14708);
or UO_1404 (O_1404,N_14726,N_14157);
and UO_1405 (O_1405,N_14359,N_14083);
nor UO_1406 (O_1406,N_14038,N_14481);
nor UO_1407 (O_1407,N_13592,N_14569);
nor UO_1408 (O_1408,N_13917,N_13956);
and UO_1409 (O_1409,N_13882,N_14382);
nor UO_1410 (O_1410,N_14211,N_14479);
nand UO_1411 (O_1411,N_14209,N_14933);
nand UO_1412 (O_1412,N_14097,N_13704);
xnor UO_1413 (O_1413,N_13947,N_14912);
and UO_1414 (O_1414,N_14065,N_13761);
xor UO_1415 (O_1415,N_14757,N_13624);
nor UO_1416 (O_1416,N_14071,N_13788);
xor UO_1417 (O_1417,N_14451,N_13741);
xor UO_1418 (O_1418,N_13602,N_13833);
or UO_1419 (O_1419,N_14446,N_14923);
or UO_1420 (O_1420,N_14396,N_14752);
nand UO_1421 (O_1421,N_14200,N_14264);
nor UO_1422 (O_1422,N_14405,N_14984);
nor UO_1423 (O_1423,N_14231,N_13658);
or UO_1424 (O_1424,N_13556,N_14588);
and UO_1425 (O_1425,N_14821,N_14367);
or UO_1426 (O_1426,N_14955,N_14716);
or UO_1427 (O_1427,N_14842,N_14232);
nand UO_1428 (O_1428,N_13642,N_14214);
nand UO_1429 (O_1429,N_14774,N_14209);
or UO_1430 (O_1430,N_14157,N_14775);
or UO_1431 (O_1431,N_14419,N_14717);
or UO_1432 (O_1432,N_14122,N_14523);
or UO_1433 (O_1433,N_13742,N_14007);
or UO_1434 (O_1434,N_14840,N_14482);
and UO_1435 (O_1435,N_14180,N_13791);
or UO_1436 (O_1436,N_13552,N_13889);
and UO_1437 (O_1437,N_13948,N_13599);
and UO_1438 (O_1438,N_13548,N_14810);
nor UO_1439 (O_1439,N_13620,N_13956);
nand UO_1440 (O_1440,N_13783,N_13750);
xor UO_1441 (O_1441,N_14975,N_14529);
nor UO_1442 (O_1442,N_13682,N_14917);
and UO_1443 (O_1443,N_14890,N_14594);
nor UO_1444 (O_1444,N_14758,N_14337);
nand UO_1445 (O_1445,N_14120,N_14431);
nand UO_1446 (O_1446,N_14550,N_13665);
or UO_1447 (O_1447,N_14766,N_14683);
or UO_1448 (O_1448,N_14370,N_14539);
nor UO_1449 (O_1449,N_14255,N_13685);
nor UO_1450 (O_1450,N_13885,N_14268);
and UO_1451 (O_1451,N_13888,N_14447);
nor UO_1452 (O_1452,N_14748,N_13831);
nand UO_1453 (O_1453,N_13828,N_14687);
xnor UO_1454 (O_1454,N_14216,N_13783);
nor UO_1455 (O_1455,N_14214,N_14629);
nor UO_1456 (O_1456,N_13595,N_14515);
nand UO_1457 (O_1457,N_13813,N_14595);
nand UO_1458 (O_1458,N_14782,N_14581);
and UO_1459 (O_1459,N_14238,N_13931);
nand UO_1460 (O_1460,N_14184,N_14609);
nor UO_1461 (O_1461,N_14227,N_13758);
nand UO_1462 (O_1462,N_14859,N_13556);
nand UO_1463 (O_1463,N_13854,N_13971);
nor UO_1464 (O_1464,N_14664,N_13972);
and UO_1465 (O_1465,N_13977,N_14910);
nor UO_1466 (O_1466,N_13745,N_13765);
nand UO_1467 (O_1467,N_14492,N_14478);
or UO_1468 (O_1468,N_13920,N_14113);
xor UO_1469 (O_1469,N_13574,N_13953);
nand UO_1470 (O_1470,N_13742,N_14176);
nor UO_1471 (O_1471,N_14091,N_13818);
or UO_1472 (O_1472,N_14737,N_13671);
and UO_1473 (O_1473,N_14315,N_14280);
nand UO_1474 (O_1474,N_14371,N_14090);
nand UO_1475 (O_1475,N_14048,N_14285);
nor UO_1476 (O_1476,N_14952,N_14274);
or UO_1477 (O_1477,N_14067,N_14418);
or UO_1478 (O_1478,N_13649,N_14416);
nand UO_1479 (O_1479,N_14023,N_14103);
nand UO_1480 (O_1480,N_14384,N_14213);
and UO_1481 (O_1481,N_13537,N_13723);
and UO_1482 (O_1482,N_14671,N_14802);
or UO_1483 (O_1483,N_13573,N_14823);
nor UO_1484 (O_1484,N_14335,N_14171);
xor UO_1485 (O_1485,N_14567,N_14676);
nand UO_1486 (O_1486,N_14843,N_14953);
nor UO_1487 (O_1487,N_13556,N_14872);
nand UO_1488 (O_1488,N_14319,N_14914);
or UO_1489 (O_1489,N_14152,N_14490);
and UO_1490 (O_1490,N_14216,N_13832);
nor UO_1491 (O_1491,N_13744,N_14428);
and UO_1492 (O_1492,N_13892,N_14731);
and UO_1493 (O_1493,N_14947,N_13919);
and UO_1494 (O_1494,N_13505,N_14216);
and UO_1495 (O_1495,N_14779,N_14172);
or UO_1496 (O_1496,N_14223,N_14478);
nand UO_1497 (O_1497,N_14923,N_14615);
nand UO_1498 (O_1498,N_14949,N_14131);
nor UO_1499 (O_1499,N_14246,N_14574);
or UO_1500 (O_1500,N_13593,N_14880);
and UO_1501 (O_1501,N_13541,N_14418);
and UO_1502 (O_1502,N_14836,N_14786);
nand UO_1503 (O_1503,N_14744,N_14410);
nor UO_1504 (O_1504,N_13563,N_13841);
nor UO_1505 (O_1505,N_13681,N_14903);
nand UO_1506 (O_1506,N_13632,N_13727);
nor UO_1507 (O_1507,N_13980,N_14331);
nand UO_1508 (O_1508,N_13768,N_13958);
xnor UO_1509 (O_1509,N_14863,N_14774);
xnor UO_1510 (O_1510,N_14865,N_14544);
nor UO_1511 (O_1511,N_14502,N_13991);
xor UO_1512 (O_1512,N_14084,N_14957);
or UO_1513 (O_1513,N_14144,N_14867);
and UO_1514 (O_1514,N_14184,N_13708);
and UO_1515 (O_1515,N_14730,N_13860);
nor UO_1516 (O_1516,N_14152,N_14038);
nor UO_1517 (O_1517,N_14938,N_14243);
nor UO_1518 (O_1518,N_14867,N_14190);
nor UO_1519 (O_1519,N_14071,N_13508);
and UO_1520 (O_1520,N_14988,N_14970);
xor UO_1521 (O_1521,N_14672,N_14981);
nand UO_1522 (O_1522,N_13523,N_14151);
nor UO_1523 (O_1523,N_14211,N_14968);
or UO_1524 (O_1524,N_14564,N_14796);
nand UO_1525 (O_1525,N_14027,N_13837);
nor UO_1526 (O_1526,N_13700,N_14593);
or UO_1527 (O_1527,N_14979,N_14278);
nor UO_1528 (O_1528,N_13647,N_14863);
and UO_1529 (O_1529,N_14106,N_14907);
nand UO_1530 (O_1530,N_13891,N_13518);
nand UO_1531 (O_1531,N_13721,N_13747);
nor UO_1532 (O_1532,N_14459,N_14401);
and UO_1533 (O_1533,N_13640,N_14276);
or UO_1534 (O_1534,N_14689,N_13861);
or UO_1535 (O_1535,N_14142,N_13693);
nor UO_1536 (O_1536,N_14882,N_13628);
or UO_1537 (O_1537,N_14226,N_14163);
and UO_1538 (O_1538,N_14315,N_14583);
and UO_1539 (O_1539,N_14952,N_14325);
or UO_1540 (O_1540,N_14177,N_13922);
and UO_1541 (O_1541,N_14249,N_14472);
nand UO_1542 (O_1542,N_13831,N_13783);
nand UO_1543 (O_1543,N_14354,N_13652);
nor UO_1544 (O_1544,N_13760,N_13671);
nand UO_1545 (O_1545,N_14799,N_14280);
or UO_1546 (O_1546,N_14314,N_14452);
nor UO_1547 (O_1547,N_14214,N_14761);
nor UO_1548 (O_1548,N_14167,N_13893);
nand UO_1549 (O_1549,N_13786,N_14308);
nand UO_1550 (O_1550,N_14890,N_13625);
nand UO_1551 (O_1551,N_13942,N_13997);
or UO_1552 (O_1552,N_13645,N_14438);
and UO_1553 (O_1553,N_14326,N_14338);
nand UO_1554 (O_1554,N_14371,N_14490);
nand UO_1555 (O_1555,N_14864,N_13608);
nand UO_1556 (O_1556,N_14293,N_13870);
nand UO_1557 (O_1557,N_13541,N_14209);
or UO_1558 (O_1558,N_14934,N_14941);
nor UO_1559 (O_1559,N_13570,N_14086);
xor UO_1560 (O_1560,N_13506,N_14367);
nand UO_1561 (O_1561,N_14187,N_14447);
or UO_1562 (O_1562,N_14947,N_13712);
nor UO_1563 (O_1563,N_14647,N_14164);
nand UO_1564 (O_1564,N_14686,N_13806);
and UO_1565 (O_1565,N_14007,N_14467);
nand UO_1566 (O_1566,N_14876,N_14206);
and UO_1567 (O_1567,N_14150,N_14992);
nand UO_1568 (O_1568,N_13773,N_14196);
nand UO_1569 (O_1569,N_14266,N_13784);
nor UO_1570 (O_1570,N_13515,N_14214);
nor UO_1571 (O_1571,N_14504,N_14482);
nor UO_1572 (O_1572,N_14659,N_14166);
nand UO_1573 (O_1573,N_13560,N_14159);
nor UO_1574 (O_1574,N_14150,N_14380);
nor UO_1575 (O_1575,N_14313,N_14606);
xnor UO_1576 (O_1576,N_14656,N_14360);
or UO_1577 (O_1577,N_14365,N_14063);
nand UO_1578 (O_1578,N_14549,N_14648);
xor UO_1579 (O_1579,N_14596,N_14135);
or UO_1580 (O_1580,N_13710,N_14474);
xor UO_1581 (O_1581,N_14095,N_14164);
nand UO_1582 (O_1582,N_14604,N_14179);
and UO_1583 (O_1583,N_14474,N_14978);
or UO_1584 (O_1584,N_14514,N_14767);
nand UO_1585 (O_1585,N_14730,N_14795);
or UO_1586 (O_1586,N_14741,N_13587);
or UO_1587 (O_1587,N_13708,N_14958);
and UO_1588 (O_1588,N_14548,N_14505);
and UO_1589 (O_1589,N_13681,N_14965);
xnor UO_1590 (O_1590,N_14778,N_14892);
nor UO_1591 (O_1591,N_13823,N_14047);
or UO_1592 (O_1592,N_14885,N_13523);
nand UO_1593 (O_1593,N_14691,N_13820);
nand UO_1594 (O_1594,N_14701,N_14986);
or UO_1595 (O_1595,N_14878,N_14431);
nand UO_1596 (O_1596,N_14177,N_14212);
nor UO_1597 (O_1597,N_14960,N_14729);
xnor UO_1598 (O_1598,N_14192,N_14868);
or UO_1599 (O_1599,N_14293,N_14084);
xor UO_1600 (O_1600,N_14499,N_13716);
or UO_1601 (O_1601,N_13807,N_14138);
nand UO_1602 (O_1602,N_14249,N_14787);
and UO_1603 (O_1603,N_14377,N_14411);
and UO_1604 (O_1604,N_14315,N_14371);
nand UO_1605 (O_1605,N_14575,N_14602);
xnor UO_1606 (O_1606,N_14882,N_13972);
nand UO_1607 (O_1607,N_14166,N_14177);
nand UO_1608 (O_1608,N_14966,N_14483);
and UO_1609 (O_1609,N_13968,N_13979);
and UO_1610 (O_1610,N_14372,N_14494);
and UO_1611 (O_1611,N_13776,N_14815);
or UO_1612 (O_1612,N_14998,N_14291);
or UO_1613 (O_1613,N_14629,N_14539);
xor UO_1614 (O_1614,N_14250,N_13885);
xor UO_1615 (O_1615,N_14807,N_14653);
nor UO_1616 (O_1616,N_14844,N_14034);
and UO_1617 (O_1617,N_14129,N_13936);
or UO_1618 (O_1618,N_14728,N_14496);
or UO_1619 (O_1619,N_13999,N_13879);
nand UO_1620 (O_1620,N_14428,N_14687);
or UO_1621 (O_1621,N_14348,N_13601);
nand UO_1622 (O_1622,N_14443,N_14228);
nor UO_1623 (O_1623,N_14988,N_14501);
or UO_1624 (O_1624,N_14136,N_14598);
nand UO_1625 (O_1625,N_13768,N_14294);
nor UO_1626 (O_1626,N_14725,N_14559);
and UO_1627 (O_1627,N_14060,N_14976);
nor UO_1628 (O_1628,N_14303,N_13797);
or UO_1629 (O_1629,N_14333,N_14469);
and UO_1630 (O_1630,N_14906,N_14919);
and UO_1631 (O_1631,N_14060,N_13950);
and UO_1632 (O_1632,N_14443,N_13962);
xnor UO_1633 (O_1633,N_14635,N_14061);
nand UO_1634 (O_1634,N_14320,N_14019);
or UO_1635 (O_1635,N_13558,N_13954);
nand UO_1636 (O_1636,N_13970,N_14245);
nor UO_1637 (O_1637,N_14326,N_14644);
and UO_1638 (O_1638,N_14633,N_14449);
or UO_1639 (O_1639,N_14561,N_13639);
and UO_1640 (O_1640,N_13529,N_13850);
or UO_1641 (O_1641,N_14728,N_14002);
nand UO_1642 (O_1642,N_14528,N_14722);
and UO_1643 (O_1643,N_14847,N_14552);
or UO_1644 (O_1644,N_14206,N_13918);
nand UO_1645 (O_1645,N_14228,N_14688);
and UO_1646 (O_1646,N_14617,N_14960);
and UO_1647 (O_1647,N_14457,N_13516);
or UO_1648 (O_1648,N_13954,N_14857);
xor UO_1649 (O_1649,N_14386,N_14710);
nor UO_1650 (O_1650,N_13598,N_14947);
xnor UO_1651 (O_1651,N_14439,N_13737);
xnor UO_1652 (O_1652,N_13507,N_14293);
and UO_1653 (O_1653,N_14932,N_14993);
and UO_1654 (O_1654,N_14906,N_13534);
or UO_1655 (O_1655,N_14852,N_14105);
and UO_1656 (O_1656,N_14854,N_13756);
or UO_1657 (O_1657,N_14719,N_13956);
xnor UO_1658 (O_1658,N_14321,N_13712);
nor UO_1659 (O_1659,N_14077,N_13842);
nor UO_1660 (O_1660,N_13713,N_13794);
xnor UO_1661 (O_1661,N_13641,N_13668);
nand UO_1662 (O_1662,N_13764,N_14363);
or UO_1663 (O_1663,N_13633,N_14469);
nand UO_1664 (O_1664,N_14108,N_14772);
and UO_1665 (O_1665,N_14841,N_13614);
or UO_1666 (O_1666,N_13521,N_14220);
nand UO_1667 (O_1667,N_14193,N_13661);
nor UO_1668 (O_1668,N_14129,N_14376);
or UO_1669 (O_1669,N_14481,N_14750);
nor UO_1670 (O_1670,N_14131,N_14016);
and UO_1671 (O_1671,N_13889,N_14914);
or UO_1672 (O_1672,N_14926,N_14851);
nand UO_1673 (O_1673,N_13712,N_13624);
nand UO_1674 (O_1674,N_14767,N_14906);
and UO_1675 (O_1675,N_14471,N_14103);
or UO_1676 (O_1676,N_14685,N_14316);
nor UO_1677 (O_1677,N_13926,N_14964);
nand UO_1678 (O_1678,N_14232,N_14241);
and UO_1679 (O_1679,N_14159,N_13607);
or UO_1680 (O_1680,N_14887,N_14949);
and UO_1681 (O_1681,N_13859,N_14380);
and UO_1682 (O_1682,N_13627,N_14022);
or UO_1683 (O_1683,N_14756,N_13837);
nand UO_1684 (O_1684,N_13945,N_13531);
xnor UO_1685 (O_1685,N_14324,N_13954);
or UO_1686 (O_1686,N_14076,N_13629);
or UO_1687 (O_1687,N_13624,N_14484);
or UO_1688 (O_1688,N_14057,N_13643);
nor UO_1689 (O_1689,N_14962,N_14147);
nand UO_1690 (O_1690,N_14122,N_14756);
xnor UO_1691 (O_1691,N_14137,N_13661);
xnor UO_1692 (O_1692,N_14565,N_13666);
nor UO_1693 (O_1693,N_14257,N_14031);
nand UO_1694 (O_1694,N_14686,N_13526);
nor UO_1695 (O_1695,N_14041,N_14349);
nor UO_1696 (O_1696,N_14272,N_13725);
nand UO_1697 (O_1697,N_14925,N_13626);
xor UO_1698 (O_1698,N_13984,N_14540);
and UO_1699 (O_1699,N_14041,N_13699);
nor UO_1700 (O_1700,N_13735,N_14003);
nand UO_1701 (O_1701,N_14412,N_14599);
nor UO_1702 (O_1702,N_14945,N_14596);
nor UO_1703 (O_1703,N_14764,N_14015);
nand UO_1704 (O_1704,N_13576,N_14843);
or UO_1705 (O_1705,N_14967,N_14120);
nand UO_1706 (O_1706,N_14858,N_14285);
nor UO_1707 (O_1707,N_13950,N_14246);
and UO_1708 (O_1708,N_14390,N_14532);
nand UO_1709 (O_1709,N_14613,N_13533);
and UO_1710 (O_1710,N_14145,N_13606);
nand UO_1711 (O_1711,N_13686,N_14165);
xnor UO_1712 (O_1712,N_13530,N_13614);
nor UO_1713 (O_1713,N_13575,N_13683);
nand UO_1714 (O_1714,N_14515,N_14061);
or UO_1715 (O_1715,N_14434,N_13509);
nand UO_1716 (O_1716,N_13765,N_14300);
xnor UO_1717 (O_1717,N_14015,N_14940);
nor UO_1718 (O_1718,N_14985,N_14654);
xor UO_1719 (O_1719,N_14626,N_13779);
nand UO_1720 (O_1720,N_14926,N_14049);
and UO_1721 (O_1721,N_14743,N_13686);
and UO_1722 (O_1722,N_14116,N_14447);
or UO_1723 (O_1723,N_14248,N_14014);
or UO_1724 (O_1724,N_14102,N_14254);
xnor UO_1725 (O_1725,N_14586,N_13949);
nor UO_1726 (O_1726,N_14561,N_13678);
nand UO_1727 (O_1727,N_14772,N_13801);
and UO_1728 (O_1728,N_13802,N_14022);
or UO_1729 (O_1729,N_13558,N_14547);
xor UO_1730 (O_1730,N_14898,N_14044);
nand UO_1731 (O_1731,N_14168,N_14989);
xnor UO_1732 (O_1732,N_13586,N_13995);
nand UO_1733 (O_1733,N_13986,N_14808);
and UO_1734 (O_1734,N_14102,N_13700);
nand UO_1735 (O_1735,N_13597,N_14930);
nand UO_1736 (O_1736,N_14735,N_13879);
and UO_1737 (O_1737,N_14231,N_13887);
and UO_1738 (O_1738,N_13890,N_14336);
and UO_1739 (O_1739,N_13549,N_13513);
and UO_1740 (O_1740,N_14873,N_14932);
or UO_1741 (O_1741,N_14555,N_13912);
and UO_1742 (O_1742,N_14674,N_14003);
nand UO_1743 (O_1743,N_13924,N_13745);
or UO_1744 (O_1744,N_13913,N_13802);
and UO_1745 (O_1745,N_14529,N_13908);
nand UO_1746 (O_1746,N_13970,N_14439);
or UO_1747 (O_1747,N_14716,N_13994);
or UO_1748 (O_1748,N_14257,N_13636);
or UO_1749 (O_1749,N_14624,N_13687);
and UO_1750 (O_1750,N_14113,N_14027);
or UO_1751 (O_1751,N_13689,N_14096);
or UO_1752 (O_1752,N_14361,N_14436);
or UO_1753 (O_1753,N_14786,N_14420);
nand UO_1754 (O_1754,N_14161,N_13734);
and UO_1755 (O_1755,N_14718,N_13810);
nand UO_1756 (O_1756,N_14202,N_14297);
nand UO_1757 (O_1757,N_14580,N_13859);
or UO_1758 (O_1758,N_14112,N_14174);
and UO_1759 (O_1759,N_13829,N_14260);
or UO_1760 (O_1760,N_13579,N_14602);
xor UO_1761 (O_1761,N_14866,N_13507);
nand UO_1762 (O_1762,N_14535,N_14676);
and UO_1763 (O_1763,N_14229,N_14174);
and UO_1764 (O_1764,N_13983,N_14029);
or UO_1765 (O_1765,N_14957,N_14436);
or UO_1766 (O_1766,N_13549,N_14297);
and UO_1767 (O_1767,N_14152,N_14417);
and UO_1768 (O_1768,N_14107,N_14898);
xor UO_1769 (O_1769,N_14785,N_14819);
nand UO_1770 (O_1770,N_13633,N_14741);
or UO_1771 (O_1771,N_14171,N_14097);
nand UO_1772 (O_1772,N_14637,N_14782);
nor UO_1773 (O_1773,N_14855,N_14730);
xnor UO_1774 (O_1774,N_14756,N_14424);
or UO_1775 (O_1775,N_13863,N_13633);
nor UO_1776 (O_1776,N_14549,N_13743);
nand UO_1777 (O_1777,N_13593,N_14156);
nor UO_1778 (O_1778,N_13602,N_13725);
nand UO_1779 (O_1779,N_14037,N_14520);
nor UO_1780 (O_1780,N_14660,N_13742);
or UO_1781 (O_1781,N_14275,N_14565);
nand UO_1782 (O_1782,N_14278,N_13883);
nand UO_1783 (O_1783,N_14312,N_14414);
nand UO_1784 (O_1784,N_14472,N_14615);
or UO_1785 (O_1785,N_13847,N_13795);
and UO_1786 (O_1786,N_14272,N_14553);
nor UO_1787 (O_1787,N_14160,N_14837);
nor UO_1788 (O_1788,N_14593,N_13826);
and UO_1789 (O_1789,N_14125,N_14838);
or UO_1790 (O_1790,N_14138,N_14445);
or UO_1791 (O_1791,N_14968,N_14831);
xor UO_1792 (O_1792,N_13772,N_14900);
and UO_1793 (O_1793,N_14033,N_14592);
or UO_1794 (O_1794,N_13635,N_14144);
nand UO_1795 (O_1795,N_14150,N_14512);
and UO_1796 (O_1796,N_14518,N_13772);
nand UO_1797 (O_1797,N_13958,N_14078);
xor UO_1798 (O_1798,N_14122,N_13714);
or UO_1799 (O_1799,N_14567,N_14825);
nor UO_1800 (O_1800,N_14078,N_14205);
or UO_1801 (O_1801,N_13576,N_14208);
and UO_1802 (O_1802,N_14465,N_14776);
nand UO_1803 (O_1803,N_14182,N_14324);
nor UO_1804 (O_1804,N_13884,N_14521);
xor UO_1805 (O_1805,N_13713,N_14566);
and UO_1806 (O_1806,N_14440,N_13647);
and UO_1807 (O_1807,N_14984,N_14222);
nor UO_1808 (O_1808,N_14920,N_13728);
and UO_1809 (O_1809,N_14892,N_13650);
or UO_1810 (O_1810,N_13856,N_13857);
nor UO_1811 (O_1811,N_13802,N_13821);
or UO_1812 (O_1812,N_14826,N_13581);
nor UO_1813 (O_1813,N_14641,N_14708);
and UO_1814 (O_1814,N_14459,N_14511);
xnor UO_1815 (O_1815,N_14423,N_13728);
or UO_1816 (O_1816,N_14668,N_14416);
and UO_1817 (O_1817,N_14205,N_14917);
nor UO_1818 (O_1818,N_14258,N_14548);
nand UO_1819 (O_1819,N_14088,N_13738);
and UO_1820 (O_1820,N_14938,N_14462);
nor UO_1821 (O_1821,N_13560,N_14027);
nand UO_1822 (O_1822,N_14758,N_13526);
nor UO_1823 (O_1823,N_13792,N_14793);
or UO_1824 (O_1824,N_13958,N_14247);
nand UO_1825 (O_1825,N_14289,N_13956);
nor UO_1826 (O_1826,N_14858,N_13648);
and UO_1827 (O_1827,N_14099,N_13737);
and UO_1828 (O_1828,N_13716,N_13885);
and UO_1829 (O_1829,N_13672,N_14235);
nor UO_1830 (O_1830,N_14176,N_14389);
nor UO_1831 (O_1831,N_14717,N_14483);
nor UO_1832 (O_1832,N_13652,N_14322);
or UO_1833 (O_1833,N_14798,N_13689);
nand UO_1834 (O_1834,N_14124,N_14771);
and UO_1835 (O_1835,N_14102,N_14192);
and UO_1836 (O_1836,N_13996,N_14522);
or UO_1837 (O_1837,N_13568,N_14482);
or UO_1838 (O_1838,N_14259,N_14528);
nor UO_1839 (O_1839,N_14064,N_14569);
nand UO_1840 (O_1840,N_14421,N_14947);
and UO_1841 (O_1841,N_14585,N_14368);
nand UO_1842 (O_1842,N_13868,N_14826);
nor UO_1843 (O_1843,N_13727,N_14263);
xnor UO_1844 (O_1844,N_14259,N_13575);
or UO_1845 (O_1845,N_13939,N_14316);
and UO_1846 (O_1846,N_13848,N_14176);
nand UO_1847 (O_1847,N_14339,N_14003);
xor UO_1848 (O_1848,N_14209,N_14959);
or UO_1849 (O_1849,N_14482,N_14844);
nor UO_1850 (O_1850,N_13728,N_13956);
nand UO_1851 (O_1851,N_13951,N_14341);
or UO_1852 (O_1852,N_14668,N_14265);
nor UO_1853 (O_1853,N_13599,N_14735);
nor UO_1854 (O_1854,N_13990,N_14597);
or UO_1855 (O_1855,N_14740,N_13783);
or UO_1856 (O_1856,N_13752,N_13941);
and UO_1857 (O_1857,N_14020,N_14526);
or UO_1858 (O_1858,N_13774,N_14576);
and UO_1859 (O_1859,N_14759,N_14829);
or UO_1860 (O_1860,N_13756,N_14544);
or UO_1861 (O_1861,N_13727,N_13680);
or UO_1862 (O_1862,N_14077,N_13527);
and UO_1863 (O_1863,N_14892,N_14166);
or UO_1864 (O_1864,N_13560,N_13792);
or UO_1865 (O_1865,N_14824,N_14135);
or UO_1866 (O_1866,N_13790,N_13739);
xnor UO_1867 (O_1867,N_13873,N_14289);
or UO_1868 (O_1868,N_14957,N_14713);
and UO_1869 (O_1869,N_14133,N_13581);
and UO_1870 (O_1870,N_13961,N_13773);
nand UO_1871 (O_1871,N_13989,N_14985);
and UO_1872 (O_1872,N_14484,N_13914);
xnor UO_1873 (O_1873,N_13595,N_14478);
or UO_1874 (O_1874,N_14302,N_13692);
and UO_1875 (O_1875,N_14982,N_14721);
nand UO_1876 (O_1876,N_14471,N_13921);
xor UO_1877 (O_1877,N_13894,N_14395);
and UO_1878 (O_1878,N_14521,N_14110);
or UO_1879 (O_1879,N_14398,N_14106);
nor UO_1880 (O_1880,N_13590,N_13665);
nor UO_1881 (O_1881,N_14356,N_14211);
or UO_1882 (O_1882,N_13831,N_13621);
or UO_1883 (O_1883,N_14574,N_13727);
and UO_1884 (O_1884,N_13860,N_14090);
and UO_1885 (O_1885,N_14851,N_14677);
xor UO_1886 (O_1886,N_14944,N_14959);
and UO_1887 (O_1887,N_14782,N_14224);
and UO_1888 (O_1888,N_14950,N_14469);
nor UO_1889 (O_1889,N_13551,N_13684);
and UO_1890 (O_1890,N_14326,N_14426);
xnor UO_1891 (O_1891,N_13947,N_13818);
or UO_1892 (O_1892,N_14514,N_14307);
nor UO_1893 (O_1893,N_14558,N_14019);
or UO_1894 (O_1894,N_13905,N_14632);
nand UO_1895 (O_1895,N_14312,N_14880);
or UO_1896 (O_1896,N_14409,N_14320);
xnor UO_1897 (O_1897,N_13975,N_13877);
or UO_1898 (O_1898,N_14070,N_14098);
nand UO_1899 (O_1899,N_13759,N_14508);
nand UO_1900 (O_1900,N_14268,N_14270);
nor UO_1901 (O_1901,N_14718,N_14745);
or UO_1902 (O_1902,N_14025,N_14318);
or UO_1903 (O_1903,N_14811,N_14195);
or UO_1904 (O_1904,N_13632,N_14778);
and UO_1905 (O_1905,N_14404,N_14822);
and UO_1906 (O_1906,N_14529,N_14504);
and UO_1907 (O_1907,N_13837,N_14638);
nor UO_1908 (O_1908,N_13840,N_14217);
nand UO_1909 (O_1909,N_14034,N_13781);
nor UO_1910 (O_1910,N_14782,N_14709);
or UO_1911 (O_1911,N_14325,N_14771);
and UO_1912 (O_1912,N_14979,N_14354);
or UO_1913 (O_1913,N_13580,N_13655);
and UO_1914 (O_1914,N_13867,N_14340);
nor UO_1915 (O_1915,N_14716,N_14292);
or UO_1916 (O_1916,N_13581,N_14889);
nand UO_1917 (O_1917,N_13825,N_14750);
and UO_1918 (O_1918,N_14027,N_13514);
nor UO_1919 (O_1919,N_14748,N_13652);
nor UO_1920 (O_1920,N_13727,N_13502);
or UO_1921 (O_1921,N_14394,N_14069);
nand UO_1922 (O_1922,N_13880,N_13847);
and UO_1923 (O_1923,N_14236,N_13834);
or UO_1924 (O_1924,N_13876,N_14232);
nand UO_1925 (O_1925,N_14063,N_13938);
or UO_1926 (O_1926,N_13507,N_14282);
nor UO_1927 (O_1927,N_14919,N_14345);
nor UO_1928 (O_1928,N_13964,N_14241);
nor UO_1929 (O_1929,N_14634,N_14592);
and UO_1930 (O_1930,N_14171,N_13752);
and UO_1931 (O_1931,N_14061,N_13781);
nand UO_1932 (O_1932,N_14161,N_14304);
nor UO_1933 (O_1933,N_14010,N_14022);
and UO_1934 (O_1934,N_13565,N_14708);
or UO_1935 (O_1935,N_14185,N_14902);
xor UO_1936 (O_1936,N_13967,N_14987);
nand UO_1937 (O_1937,N_14470,N_14075);
nand UO_1938 (O_1938,N_14893,N_13544);
and UO_1939 (O_1939,N_14563,N_14458);
nand UO_1940 (O_1940,N_13751,N_14743);
or UO_1941 (O_1941,N_14116,N_13717);
or UO_1942 (O_1942,N_13966,N_13522);
or UO_1943 (O_1943,N_14521,N_14471);
and UO_1944 (O_1944,N_14983,N_14071);
nand UO_1945 (O_1945,N_14489,N_14885);
and UO_1946 (O_1946,N_14829,N_14821);
or UO_1947 (O_1947,N_13611,N_14438);
nor UO_1948 (O_1948,N_13615,N_14356);
or UO_1949 (O_1949,N_13697,N_14627);
nand UO_1950 (O_1950,N_13976,N_14578);
or UO_1951 (O_1951,N_14112,N_14637);
or UO_1952 (O_1952,N_14770,N_14327);
nand UO_1953 (O_1953,N_13830,N_14887);
xnor UO_1954 (O_1954,N_13535,N_14969);
nor UO_1955 (O_1955,N_14568,N_14002);
nand UO_1956 (O_1956,N_14225,N_14663);
nand UO_1957 (O_1957,N_14627,N_13982);
nand UO_1958 (O_1958,N_14389,N_14162);
and UO_1959 (O_1959,N_14740,N_13807);
or UO_1960 (O_1960,N_13762,N_14126);
and UO_1961 (O_1961,N_14612,N_13970);
and UO_1962 (O_1962,N_14306,N_14450);
nor UO_1963 (O_1963,N_14681,N_13662);
xnor UO_1964 (O_1964,N_14581,N_13826);
or UO_1965 (O_1965,N_13957,N_13717);
nand UO_1966 (O_1966,N_14053,N_13679);
nand UO_1967 (O_1967,N_14817,N_14555);
and UO_1968 (O_1968,N_13566,N_14401);
and UO_1969 (O_1969,N_14563,N_13952);
nand UO_1970 (O_1970,N_14675,N_14559);
or UO_1971 (O_1971,N_14381,N_13632);
nand UO_1972 (O_1972,N_14428,N_13675);
nand UO_1973 (O_1973,N_14300,N_13569);
nor UO_1974 (O_1974,N_14772,N_14739);
nor UO_1975 (O_1975,N_14693,N_14395);
nor UO_1976 (O_1976,N_13561,N_13771);
nor UO_1977 (O_1977,N_14600,N_13507);
nand UO_1978 (O_1978,N_14828,N_13640);
nor UO_1979 (O_1979,N_14630,N_14689);
or UO_1980 (O_1980,N_13658,N_14530);
and UO_1981 (O_1981,N_14063,N_14878);
nand UO_1982 (O_1982,N_14146,N_13665);
and UO_1983 (O_1983,N_13642,N_13883);
nor UO_1984 (O_1984,N_14989,N_13813);
or UO_1985 (O_1985,N_13683,N_13665);
nor UO_1986 (O_1986,N_14058,N_13556);
or UO_1987 (O_1987,N_13928,N_14493);
nor UO_1988 (O_1988,N_14455,N_14763);
and UO_1989 (O_1989,N_14668,N_14625);
and UO_1990 (O_1990,N_14053,N_13609);
and UO_1991 (O_1991,N_14711,N_14374);
xnor UO_1992 (O_1992,N_13886,N_14911);
and UO_1993 (O_1993,N_13696,N_14959);
nand UO_1994 (O_1994,N_14362,N_14966);
or UO_1995 (O_1995,N_14210,N_14500);
and UO_1996 (O_1996,N_14132,N_14971);
or UO_1997 (O_1997,N_14178,N_13764);
nand UO_1998 (O_1998,N_13858,N_14485);
and UO_1999 (O_1999,N_14232,N_14788);
endmodule