module basic_750_5000_1000_2_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2504,N_2505,N_2506,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2516,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2532,N_2533,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2545,N_2547,N_2548,N_2549,N_2550,N_2551,N_2553,N_2554,N_2556,N_2557,N_2559,N_2560,N_2561,N_2563,N_2564,N_2565,N_2567,N_2569,N_2570,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2618,N_2619,N_2620,N_2622,N_2623,N_2625,N_2626,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2662,N_2663,N_2664,N_2665,N_2667,N_2668,N_2669,N_2670,N_2671,N_2673,N_2674,N_2675,N_2677,N_2678,N_2679,N_2681,N_2682,N_2683,N_2685,N_2686,N_2688,N_2689,N_2690,N_2692,N_2693,N_2694,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2705,N_2706,N_2707,N_2708,N_2710,N_2712,N_2713,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2763,N_2765,N_2766,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2780,N_2781,N_2782,N_2783,N_2784,N_2787,N_2788,N_2790,N_2792,N_2793,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2807,N_2809,N_2810,N_2811,N_2812,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2822,N_2823,N_2826,N_2827,N_2828,N_2829,N_2830,N_2832,N_2833,N_2834,N_2835,N_2837,N_2838,N_2839,N_2840,N_2841,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2864,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2913,N_2914,N_2917,N_2919,N_2920,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2931,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2947,N_2949,N_2950,N_2951,N_2952,N_2953,N_2956,N_2959,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2979,N_2980,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3007,N_3008,N_3011,N_3012,N_3013,N_3015,N_3017,N_3018,N_3019,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3073,N_3076,N_3077,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3091,N_3092,N_3093,N_3094,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3111,N_3113,N_3114,N_3115,N_3117,N_3118,N_3119,N_3120,N_3123,N_3124,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3147,N_3148,N_3149,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3160,N_3161,N_3162,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3172,N_3174,N_3175,N_3178,N_3179,N_3182,N_3183,N_3184,N_3185,N_3186,N_3188,N_3189,N_3190,N_3191,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3200,N_3201,N_3202,N_3204,N_3205,N_3207,N_3208,N_3211,N_3212,N_3213,N_3214,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3227,N_3228,N_3229,N_3232,N_3234,N_3235,N_3236,N_3237,N_3238,N_3240,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3259,N_3260,N_3261,N_3264,N_3266,N_3268,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3290,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3308,N_3310,N_3312,N_3313,N_3315,N_3316,N_3317,N_3320,N_3323,N_3324,N_3325,N_3326,N_3327,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3337,N_3338,N_3339,N_3340,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3385,N_3387,N_3388,N_3390,N_3392,N_3394,N_3395,N_3396,N_3397,N_3399,N_3400,N_3401,N_3402,N_3403,N_3405,N_3407,N_3408,N_3410,N_3411,N_3412,N_3413,N_3415,N_3417,N_3418,N_3419,N_3420,N_3422,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3432,N_3433,N_3435,N_3436,N_3438,N_3439,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3450,N_3451,N_3452,N_3454,N_3455,N_3456,N_3457,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3466,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3493,N_3494,N_3496,N_3498,N_3499,N_3502,N_3503,N_3504,N_3505,N_3507,N_3508,N_3511,N_3512,N_3513,N_3514,N_3515,N_3519,N_3520,N_3521,N_3522,N_3524,N_3525,N_3527,N_3528,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3547,N_3548,N_3549,N_3550,N_3552,N_3553,N_3554,N_3555,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3566,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3590,N_3591,N_3592,N_3593,N_3594,N_3596,N_3598,N_3599,N_3602,N_3603,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3613,N_3614,N_3615,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3644,N_3645,N_3646,N_3648,N_3650,N_3651,N_3652,N_3653,N_3654,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3678,N_3679,N_3680,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3689,N_3690,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3713,N_3714,N_3716,N_3717,N_3718,N_3720,N_3722,N_3723,N_3724,N_3726,N_3727,N_3728,N_3733,N_3734,N_3735,N_3736,N_3739,N_3741,N_3742,N_3744,N_3746,N_3747,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3759,N_3760,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3771,N_3772,N_3773,N_3775,N_3776,N_3777,N_3778,N_3780,N_3781,N_3782,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3821,N_3823,N_3824,N_3825,N_3826,N_3827,N_3829,N_3831,N_3832,N_3833,N_3836,N_3837,N_3838,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3862,N_3863,N_3867,N_3869,N_3870,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3885,N_3886,N_3888,N_3889,N_3890,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3930,N_3932,N_3933,N_3936,N_3937,N_3939,N_3940,N_3941,N_3942,N_3943,N_3945,N_3947,N_3948,N_3951,N_3952,N_3953,N_3954,N_3956,N_3957,N_3958,N_3959,N_3960,N_3963,N_3965,N_3967,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3983,N_3985,N_3986,N_3987,N_3989,N_3990,N_3993,N_3994,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4016,N_4017,N_4018,N_4019,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4035,N_4036,N_4037,N_4038,N_4039,N_4041,N_4042,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4057,N_4059,N_4060,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4102,N_4104,N_4105,N_4106,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4159,N_4160,N_4161,N_4162,N_4163,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4173,N_4174,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4185,N_4186,N_4187,N_4189,N_4191,N_4192,N_4193,N_4194,N_4195,N_4198,N_4199,N_4200,N_4202,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4226,N_4227,N_4228,N_4229,N_4230,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4263,N_4265,N_4266,N_4267,N_4268,N_4269,N_4271,N_4272,N_4273,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4292,N_4294,N_4295,N_4296,N_4298,N_4299,N_4300,N_4301,N_4302,N_4304,N_4305,N_4306,N_4307,N_4308,N_4310,N_4311,N_4313,N_4314,N_4316,N_4317,N_4318,N_4320,N_4321,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4355,N_4356,N_4357,N_4360,N_4362,N_4364,N_4365,N_4366,N_4368,N_4369,N_4371,N_4372,N_4373,N_4374,N_4376,N_4377,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4387,N_4388,N_4389,N_4391,N_4392,N_4393,N_4394,N_4396,N_4398,N_4399,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4410,N_4412,N_4413,N_4414,N_4415,N_4417,N_4418,N_4420,N_4421,N_4423,N_4424,N_4426,N_4427,N_4429,N_4431,N_4432,N_4433,N_4436,N_4437,N_4438,N_4440,N_4441,N_4442,N_4444,N_4445,N_4447,N_4448,N_4449,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4462,N_4463,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4482,N_4483,N_4484,N_4485,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4509,N_4510,N_4511,N_4512,N_4513,N_4516,N_4517,N_4519,N_4520,N_4521,N_4522,N_4523,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4534,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4544,N_4545,N_4546,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4556,N_4557,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4569,N_4570,N_4571,N_4572,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4583,N_4584,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4609,N_4610,N_4611,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4625,N_4627,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4639,N_4640,N_4641,N_4642,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4653,N_4654,N_4655,N_4656,N_4657,N_4659,N_4660,N_4661,N_4662,N_4664,N_4665,N_4667,N_4668,N_4669,N_4670,N_4671,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4684,N_4685,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4695,N_4698,N_4699,N_4700,N_4701,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4710,N_4711,N_4712,N_4713,N_4715,N_4716,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4728,N_4729,N_4731,N_4733,N_4734,N_4735,N_4736,N_4737,N_4739,N_4740,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4752,N_4753,N_4754,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4779,N_4780,N_4781,N_4782,N_4783,N_4787,N_4788,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4839,N_4840,N_4841,N_4843,N_4844,N_4845,N_4846,N_4849,N_4850,N_4852,N_4853,N_4855,N_4856,N_4857,N_4858,N_4859,N_4861,N_4862,N_4864,N_4865,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4885,N_4887,N_4888,N_4890,N_4893,N_4895,N_4896,N_4897,N_4898,N_4899,N_4903,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4916,N_4917,N_4918,N_4920,N_4921,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4931,N_4933,N_4934,N_4935,N_4937,N_4939,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4970,N_4971,N_4972,N_4973,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4987,N_4988,N_4989,N_4990,N_4994,N_4995,N_4997,N_4998,N_4999;
or U0 (N_0,In_530,In_115);
and U1 (N_1,In_337,In_414);
or U2 (N_2,In_16,In_598);
nand U3 (N_3,In_244,In_657);
or U4 (N_4,In_617,In_384);
or U5 (N_5,In_445,In_717);
xor U6 (N_6,In_694,In_167);
nand U7 (N_7,In_381,In_301);
and U8 (N_8,In_524,In_538);
nand U9 (N_9,In_300,In_701);
and U10 (N_10,In_472,In_440);
or U11 (N_11,In_361,In_41);
and U12 (N_12,In_336,In_290);
and U13 (N_13,In_747,In_29);
and U14 (N_14,In_486,In_111);
and U15 (N_15,In_628,In_233);
or U16 (N_16,In_514,In_122);
nand U17 (N_17,In_711,In_293);
nand U18 (N_18,In_456,In_629);
or U19 (N_19,In_296,In_263);
nor U20 (N_20,In_407,In_674);
xnor U21 (N_21,In_183,In_699);
nor U22 (N_22,In_412,In_75);
nand U23 (N_23,In_579,In_606);
nor U24 (N_24,In_248,In_366);
nor U25 (N_25,In_600,In_80);
nand U26 (N_26,In_370,In_220);
xnor U27 (N_27,In_282,In_663);
nand U28 (N_28,In_665,In_613);
and U29 (N_29,In_395,In_119);
and U30 (N_30,In_174,In_466);
or U31 (N_31,In_481,In_417);
and U32 (N_32,In_670,In_311);
or U33 (N_33,In_177,In_705);
nor U34 (N_34,In_572,In_398);
and U35 (N_35,In_616,In_159);
or U36 (N_36,In_340,In_360);
or U37 (N_37,In_238,In_592);
nor U38 (N_38,In_17,In_131);
nor U39 (N_39,In_744,In_79);
or U40 (N_40,In_27,In_583);
nand U41 (N_41,In_275,In_318);
nand U42 (N_42,In_170,In_353);
and U43 (N_43,In_324,In_476);
or U44 (N_44,In_518,In_568);
or U45 (N_45,In_327,In_432);
nor U46 (N_46,In_22,In_684);
nand U47 (N_47,In_439,In_457);
or U48 (N_48,In_737,In_304);
nand U49 (N_49,In_430,In_371);
and U50 (N_50,In_543,In_148);
and U51 (N_51,In_206,In_356);
or U52 (N_52,In_165,In_287);
and U53 (N_53,In_349,In_721);
and U54 (N_54,In_100,In_603);
or U55 (N_55,In_639,In_215);
nand U56 (N_56,In_186,In_72);
nand U57 (N_57,In_685,In_709);
and U58 (N_58,In_310,In_470);
nand U59 (N_59,In_557,In_633);
and U60 (N_60,In_124,In_362);
or U61 (N_61,In_139,In_230);
or U62 (N_62,In_658,In_143);
or U63 (N_63,In_601,In_6);
and U64 (N_64,In_36,In_730);
nor U65 (N_65,In_621,In_178);
nor U66 (N_66,In_333,In_660);
nor U67 (N_67,In_331,In_279);
nor U68 (N_68,In_526,In_461);
or U69 (N_69,In_224,In_489);
nand U70 (N_70,In_130,In_295);
nand U71 (N_71,In_96,In_582);
and U72 (N_72,In_490,In_671);
nand U73 (N_73,In_630,In_508);
nand U74 (N_74,In_385,In_452);
and U75 (N_75,In_650,In_483);
nand U76 (N_76,In_229,In_307);
and U77 (N_77,In_597,In_471);
nor U78 (N_78,In_453,In_49);
nor U79 (N_79,In_271,In_382);
and U80 (N_80,In_302,In_442);
and U81 (N_81,In_716,In_259);
nand U82 (N_82,In_506,In_61);
nor U83 (N_83,In_67,In_492);
or U84 (N_84,In_463,In_644);
nand U85 (N_85,In_460,In_351);
or U86 (N_86,In_163,In_535);
nand U87 (N_87,In_200,In_609);
and U88 (N_88,In_677,In_433);
nor U89 (N_89,In_522,In_221);
nor U90 (N_90,In_156,In_107);
and U91 (N_91,In_653,In_517);
nand U92 (N_92,In_624,In_493);
nor U93 (N_93,In_113,In_208);
or U94 (N_94,In_212,In_98);
nand U95 (N_95,In_54,In_559);
or U96 (N_96,In_140,In_235);
nand U97 (N_97,In_288,In_724);
and U98 (N_98,In_249,In_531);
nand U99 (N_99,In_74,In_306);
nor U100 (N_100,In_93,In_438);
or U101 (N_101,In_210,In_561);
nand U102 (N_102,In_689,In_283);
nand U103 (N_103,In_323,In_291);
and U104 (N_104,In_733,In_478);
or U105 (N_105,In_241,In_652);
nor U106 (N_106,In_24,In_71);
and U107 (N_107,In_268,In_151);
nand U108 (N_108,In_570,In_297);
nand U109 (N_109,In_4,In_133);
nand U110 (N_110,In_242,In_343);
and U111 (N_111,In_569,In_15);
nor U112 (N_112,In_722,In_181);
nand U113 (N_113,In_97,In_128);
nor U114 (N_114,In_649,In_120);
and U115 (N_115,In_399,In_626);
nand U116 (N_116,In_718,In_147);
and U117 (N_117,In_618,In_607);
nand U118 (N_118,In_545,In_428);
nand U119 (N_119,In_541,In_467);
nand U120 (N_120,In_222,In_686);
nand U121 (N_121,In_392,In_389);
and U122 (N_122,In_298,In_155);
nor U123 (N_123,In_552,In_416);
nor U124 (N_124,In_421,In_105);
nand U125 (N_125,In_313,In_95);
nand U126 (N_126,In_741,In_116);
or U127 (N_127,In_203,In_668);
and U128 (N_128,In_134,In_51);
nor U129 (N_129,In_710,In_114);
or U130 (N_130,In_34,In_89);
or U131 (N_131,In_218,In_525);
or U132 (N_132,In_145,In_544);
or U133 (N_133,In_553,In_488);
nor U134 (N_134,In_123,In_317);
or U135 (N_135,In_566,In_136);
or U136 (N_136,In_329,In_448);
nor U137 (N_137,In_158,In_546);
nand U138 (N_138,In_459,In_322);
nor U139 (N_139,In_620,In_697);
and U140 (N_140,In_47,In_443);
nand U141 (N_141,In_176,In_519);
nor U142 (N_142,In_247,In_664);
and U143 (N_143,In_109,In_556);
nor U144 (N_144,In_18,In_70);
nor U145 (N_145,In_272,In_405);
nor U146 (N_146,In_437,In_104);
nand U147 (N_147,In_704,In_394);
nand U148 (N_148,In_496,In_435);
or U149 (N_149,In_189,In_184);
nand U150 (N_150,In_396,In_73);
and U151 (N_151,In_129,In_286);
nand U152 (N_152,In_328,In_19);
and U153 (N_153,In_213,In_53);
and U154 (N_154,In_719,In_610);
xor U155 (N_155,In_692,In_415);
and U156 (N_156,In_202,In_266);
and U157 (N_157,In_125,In_11);
or U158 (N_158,In_108,In_444);
nor U159 (N_159,In_270,In_35);
or U160 (N_160,In_182,In_599);
nand U161 (N_161,In_565,In_258);
nand U162 (N_162,In_154,In_118);
nand U163 (N_163,In_708,In_539);
nand U164 (N_164,In_547,In_192);
xnor U165 (N_165,In_162,In_110);
nand U166 (N_166,In_216,In_254);
nand U167 (N_167,In_339,In_742);
or U168 (N_168,In_634,In_500);
nor U169 (N_169,In_408,In_294);
and U170 (N_170,In_198,In_369);
or U171 (N_171,In_669,In_625);
and U172 (N_172,In_427,In_277);
and U173 (N_173,In_646,In_431);
nor U174 (N_174,In_739,In_46);
nor U175 (N_175,In_92,In_37);
nand U176 (N_176,In_595,In_83);
xor U177 (N_177,In_316,In_12);
nand U178 (N_178,In_341,In_503);
or U179 (N_179,In_269,In_121);
nand U180 (N_180,In_373,In_693);
nand U181 (N_181,In_315,In_391);
nor U182 (N_182,In_179,In_214);
nand U183 (N_183,In_289,In_454);
and U184 (N_184,In_7,In_587);
nor U185 (N_185,In_175,In_554);
and U186 (N_186,In_409,In_64);
or U187 (N_187,In_205,In_90);
nand U188 (N_188,In_255,In_661);
nand U189 (N_189,In_511,In_707);
or U190 (N_190,In_169,In_513);
nor U191 (N_191,In_484,In_720);
nor U192 (N_192,In_462,In_387);
nor U193 (N_193,In_573,In_374);
nor U194 (N_194,In_560,In_659);
nand U195 (N_195,In_403,In_577);
nor U196 (N_196,In_355,In_586);
or U197 (N_197,In_1,In_564);
xor U198 (N_198,In_66,In_365);
or U199 (N_199,In_691,In_728);
nand U200 (N_200,In_228,In_173);
or U201 (N_201,In_429,In_250);
or U202 (N_202,In_528,In_91);
or U203 (N_203,In_731,In_326);
and U204 (N_204,In_201,In_729);
and U205 (N_205,In_33,In_354);
or U206 (N_206,In_135,In_44);
nand U207 (N_207,In_527,In_636);
and U208 (N_208,In_112,In_594);
or U209 (N_209,In_474,In_14);
nor U210 (N_210,In_563,In_171);
nand U211 (N_211,In_5,In_725);
or U212 (N_212,In_498,In_501);
nor U213 (N_213,In_672,In_204);
nand U214 (N_214,In_550,In_132);
or U215 (N_215,In_520,In_191);
nand U216 (N_216,In_190,In_161);
nand U217 (N_217,In_487,In_342);
nand U218 (N_218,In_166,In_319);
nand U219 (N_219,In_168,In_284);
and U220 (N_220,In_357,In_655);
nor U221 (N_221,In_676,In_332);
nand U222 (N_222,In_548,In_376);
or U223 (N_223,In_464,In_714);
and U224 (N_224,In_736,In_312);
nor U225 (N_225,In_211,In_651);
nand U226 (N_226,In_584,In_345);
and U227 (N_227,In_540,In_23);
and U228 (N_228,In_509,In_611);
nand U229 (N_229,In_101,In_62);
nand U230 (N_230,In_185,In_436);
or U231 (N_231,In_127,In_292);
and U232 (N_232,In_262,In_473);
nor U233 (N_233,In_627,In_378);
nand U234 (N_234,In_605,In_726);
nor U235 (N_235,In_450,In_58);
or U236 (N_236,In_642,In_278);
nand U237 (N_237,In_732,In_38);
nor U238 (N_238,In_223,In_648);
nand U239 (N_239,In_193,In_334);
and U240 (N_240,In_146,In_142);
or U241 (N_241,In_225,In_13);
nor U242 (N_242,In_314,In_590);
nand U243 (N_243,In_604,In_172);
nand U244 (N_244,In_375,In_358);
or U245 (N_245,In_48,In_465);
and U246 (N_246,In_533,In_25);
xnor U247 (N_247,In_364,In_441);
or U248 (N_248,In_700,In_153);
nor U249 (N_249,In_688,In_702);
and U250 (N_250,In_523,In_749);
and U251 (N_251,In_31,In_542);
or U252 (N_252,In_390,In_256);
nor U253 (N_253,In_643,In_401);
nand U254 (N_254,In_305,In_551);
and U255 (N_255,In_232,In_424);
nand U256 (N_256,In_614,In_638);
or U257 (N_257,In_695,In_320);
nand U258 (N_258,In_683,In_469);
and U259 (N_259,In_529,In_240);
or U260 (N_260,In_422,In_141);
and U261 (N_261,In_502,In_50);
and U262 (N_262,In_510,In_562);
and U263 (N_263,In_102,In_348);
and U264 (N_264,In_45,In_420);
and U265 (N_265,In_68,In_9);
and U266 (N_266,In_404,In_706);
and U267 (N_267,In_94,In_372);
nand U268 (N_268,In_679,In_30);
nor U269 (N_269,In_678,In_580);
or U270 (N_270,In_207,In_265);
nand U271 (N_271,In_26,In_377);
nand U272 (N_272,In_69,In_589);
or U273 (N_273,In_734,In_63);
or U274 (N_274,In_219,In_76);
and U275 (N_275,In_137,In_451);
xor U276 (N_276,In_507,In_713);
and U277 (N_277,In_619,In_363);
or U278 (N_278,In_723,In_126);
and U279 (N_279,In_65,In_257);
nand U280 (N_280,In_379,In_88);
nand U281 (N_281,In_60,In_195);
nand U282 (N_282,In_346,In_197);
and U283 (N_283,In_81,In_252);
or U284 (N_284,In_187,In_696);
and U285 (N_285,In_637,In_578);
and U286 (N_286,In_393,In_144);
or U287 (N_287,In_675,In_55);
and U288 (N_288,In_475,In_234);
or U289 (N_289,In_84,In_571);
and U290 (N_290,In_309,In_209);
or U291 (N_291,In_491,In_138);
or U292 (N_292,In_662,In_641);
nor U293 (N_293,In_534,In_164);
or U294 (N_294,In_574,In_690);
and U295 (N_295,In_419,In_82);
and U296 (N_296,In_152,In_632);
nor U297 (N_297,In_581,In_681);
and U298 (N_298,In_727,In_330);
or U299 (N_299,In_85,In_386);
and U300 (N_300,In_576,In_87);
or U301 (N_301,In_400,In_423);
nand U302 (N_302,In_180,In_426);
or U303 (N_303,In_347,In_264);
nand U304 (N_304,In_231,In_103);
and U305 (N_305,In_199,In_56);
xor U306 (N_306,In_499,In_359);
nor U307 (N_307,In_458,In_52);
nand U308 (N_308,In_494,In_246);
and U309 (N_309,In_588,In_504);
nor U310 (N_310,In_656,In_239);
nand U311 (N_311,In_703,In_715);
nand U312 (N_312,In_285,In_43);
nand U313 (N_313,In_698,In_615);
nand U314 (N_314,In_253,In_157);
nand U315 (N_315,In_303,In_558);
nand U316 (N_316,In_645,In_194);
nand U317 (N_317,In_40,In_555);
and U318 (N_318,In_712,In_575);
and U319 (N_319,In_468,In_299);
or U320 (N_320,In_667,In_383);
nor U321 (N_321,In_281,In_682);
nor U322 (N_322,In_308,In_77);
or U323 (N_323,In_406,In_78);
nor U324 (N_324,In_748,In_647);
and U325 (N_325,In_196,In_521);
and U326 (N_326,In_505,In_352);
nor U327 (N_327,In_434,In_267);
and U328 (N_328,In_367,In_160);
and U329 (N_329,In_479,In_261);
nor U330 (N_330,In_86,In_640);
or U331 (N_331,In_485,In_99);
and U332 (N_332,In_673,In_593);
or U333 (N_333,In_532,In_623);
nand U334 (N_334,In_251,In_495);
or U335 (N_335,In_188,In_260);
nor U336 (N_336,In_743,In_515);
and U337 (N_337,In_39,In_150);
nor U338 (N_338,In_635,In_622);
and U339 (N_339,In_280,In_536);
or U340 (N_340,In_516,In_745);
nand U341 (N_341,In_20,In_447);
nand U342 (N_342,In_338,In_106);
and U343 (N_343,In_735,In_549);
nor U344 (N_344,In_631,In_608);
nor U345 (N_345,In_449,In_325);
nor U346 (N_346,In_117,In_680);
and U347 (N_347,In_537,In_32);
and U348 (N_348,In_149,In_687);
nor U349 (N_349,In_217,In_413);
and U350 (N_350,In_425,In_567);
nor U351 (N_351,In_57,In_2);
and U352 (N_352,In_738,In_226);
nor U353 (N_353,In_446,In_59);
nand U354 (N_354,In_477,In_482);
nor U355 (N_355,In_321,In_480);
or U356 (N_356,In_418,In_227);
and U357 (N_357,In_350,In_612);
nor U358 (N_358,In_28,In_276);
nand U359 (N_359,In_274,In_591);
nor U360 (N_360,In_236,In_746);
nand U361 (N_361,In_243,In_368);
nand U362 (N_362,In_410,In_455);
nand U363 (N_363,In_654,In_388);
nand U364 (N_364,In_42,In_497);
xnor U365 (N_365,In_21,In_245);
or U366 (N_366,In_411,In_3);
or U367 (N_367,In_512,In_397);
and U368 (N_368,In_8,In_273);
nand U369 (N_369,In_596,In_402);
nand U370 (N_370,In_10,In_380);
or U371 (N_371,In_237,In_740);
and U372 (N_372,In_344,In_585);
nand U373 (N_373,In_0,In_666);
or U374 (N_374,In_602,In_335);
nor U375 (N_375,In_682,In_526);
nand U376 (N_376,In_5,In_608);
and U377 (N_377,In_393,In_78);
nand U378 (N_378,In_450,In_300);
or U379 (N_379,In_55,In_661);
nor U380 (N_380,In_85,In_671);
and U381 (N_381,In_481,In_350);
nand U382 (N_382,In_579,In_392);
xnor U383 (N_383,In_382,In_113);
or U384 (N_384,In_11,In_328);
nor U385 (N_385,In_41,In_690);
nand U386 (N_386,In_239,In_277);
nor U387 (N_387,In_675,In_142);
and U388 (N_388,In_660,In_271);
and U389 (N_389,In_448,In_668);
and U390 (N_390,In_74,In_93);
xnor U391 (N_391,In_516,In_224);
nor U392 (N_392,In_196,In_640);
and U393 (N_393,In_197,In_344);
and U394 (N_394,In_102,In_178);
nand U395 (N_395,In_591,In_560);
nand U396 (N_396,In_450,In_725);
xnor U397 (N_397,In_680,In_335);
or U398 (N_398,In_248,In_333);
nand U399 (N_399,In_478,In_718);
or U400 (N_400,In_728,In_610);
nand U401 (N_401,In_44,In_589);
nor U402 (N_402,In_123,In_235);
nand U403 (N_403,In_325,In_45);
nor U404 (N_404,In_189,In_182);
and U405 (N_405,In_562,In_154);
nor U406 (N_406,In_123,In_102);
and U407 (N_407,In_3,In_451);
nor U408 (N_408,In_740,In_138);
nand U409 (N_409,In_149,In_366);
or U410 (N_410,In_76,In_335);
nor U411 (N_411,In_510,In_374);
nor U412 (N_412,In_30,In_608);
and U413 (N_413,In_195,In_459);
nor U414 (N_414,In_387,In_147);
nand U415 (N_415,In_180,In_96);
nor U416 (N_416,In_591,In_497);
or U417 (N_417,In_364,In_12);
or U418 (N_418,In_741,In_140);
nor U419 (N_419,In_731,In_390);
nand U420 (N_420,In_250,In_246);
nor U421 (N_421,In_396,In_229);
nor U422 (N_422,In_718,In_619);
and U423 (N_423,In_291,In_452);
nor U424 (N_424,In_186,In_467);
and U425 (N_425,In_564,In_280);
nor U426 (N_426,In_556,In_175);
and U427 (N_427,In_101,In_495);
nor U428 (N_428,In_60,In_576);
xnor U429 (N_429,In_399,In_181);
and U430 (N_430,In_45,In_66);
and U431 (N_431,In_692,In_399);
and U432 (N_432,In_651,In_610);
nand U433 (N_433,In_340,In_253);
nand U434 (N_434,In_271,In_128);
nor U435 (N_435,In_521,In_113);
or U436 (N_436,In_439,In_294);
and U437 (N_437,In_2,In_568);
nor U438 (N_438,In_293,In_404);
nand U439 (N_439,In_694,In_674);
nand U440 (N_440,In_172,In_434);
nand U441 (N_441,In_615,In_128);
nand U442 (N_442,In_165,In_206);
nand U443 (N_443,In_546,In_473);
nand U444 (N_444,In_352,In_615);
or U445 (N_445,In_504,In_200);
and U446 (N_446,In_716,In_290);
or U447 (N_447,In_504,In_660);
or U448 (N_448,In_459,In_258);
and U449 (N_449,In_440,In_649);
nand U450 (N_450,In_499,In_5);
xor U451 (N_451,In_518,In_495);
and U452 (N_452,In_260,In_561);
nor U453 (N_453,In_592,In_388);
or U454 (N_454,In_633,In_61);
or U455 (N_455,In_150,In_102);
nand U456 (N_456,In_675,In_66);
xnor U457 (N_457,In_490,In_281);
nor U458 (N_458,In_639,In_139);
nor U459 (N_459,In_559,In_38);
or U460 (N_460,In_108,In_127);
and U461 (N_461,In_604,In_250);
and U462 (N_462,In_599,In_139);
and U463 (N_463,In_606,In_170);
nand U464 (N_464,In_731,In_553);
and U465 (N_465,In_13,In_331);
nand U466 (N_466,In_504,In_378);
or U467 (N_467,In_250,In_2);
or U468 (N_468,In_418,In_304);
xor U469 (N_469,In_433,In_168);
nor U470 (N_470,In_76,In_401);
nor U471 (N_471,In_575,In_273);
nand U472 (N_472,In_343,In_366);
nand U473 (N_473,In_38,In_675);
nand U474 (N_474,In_746,In_125);
xnor U475 (N_475,In_662,In_117);
and U476 (N_476,In_79,In_630);
nand U477 (N_477,In_238,In_58);
or U478 (N_478,In_599,In_651);
nor U479 (N_479,In_622,In_351);
or U480 (N_480,In_62,In_438);
nor U481 (N_481,In_609,In_284);
or U482 (N_482,In_280,In_181);
nand U483 (N_483,In_139,In_68);
nand U484 (N_484,In_741,In_196);
and U485 (N_485,In_181,In_651);
nand U486 (N_486,In_176,In_682);
or U487 (N_487,In_305,In_89);
nor U488 (N_488,In_45,In_599);
nor U489 (N_489,In_247,In_261);
nand U490 (N_490,In_270,In_611);
and U491 (N_491,In_586,In_192);
nand U492 (N_492,In_439,In_655);
nor U493 (N_493,In_616,In_651);
nand U494 (N_494,In_562,In_613);
nor U495 (N_495,In_212,In_684);
and U496 (N_496,In_557,In_380);
and U497 (N_497,In_0,In_585);
nand U498 (N_498,In_652,In_263);
or U499 (N_499,In_621,In_734);
nor U500 (N_500,In_113,In_24);
nand U501 (N_501,In_22,In_242);
nand U502 (N_502,In_75,In_558);
nand U503 (N_503,In_288,In_440);
nand U504 (N_504,In_573,In_497);
and U505 (N_505,In_89,In_516);
xnor U506 (N_506,In_314,In_591);
and U507 (N_507,In_189,In_617);
or U508 (N_508,In_658,In_328);
or U509 (N_509,In_507,In_526);
or U510 (N_510,In_362,In_681);
nor U511 (N_511,In_351,In_424);
and U512 (N_512,In_557,In_673);
nor U513 (N_513,In_403,In_547);
nand U514 (N_514,In_145,In_703);
or U515 (N_515,In_639,In_54);
nand U516 (N_516,In_651,In_104);
nand U517 (N_517,In_220,In_480);
nand U518 (N_518,In_217,In_105);
and U519 (N_519,In_472,In_689);
or U520 (N_520,In_234,In_381);
nand U521 (N_521,In_272,In_522);
or U522 (N_522,In_591,In_96);
nor U523 (N_523,In_571,In_441);
xor U524 (N_524,In_395,In_602);
and U525 (N_525,In_532,In_516);
or U526 (N_526,In_711,In_670);
xor U527 (N_527,In_254,In_525);
xor U528 (N_528,In_391,In_168);
or U529 (N_529,In_388,In_107);
nand U530 (N_530,In_575,In_518);
and U531 (N_531,In_254,In_670);
nand U532 (N_532,In_145,In_275);
nand U533 (N_533,In_677,In_438);
or U534 (N_534,In_749,In_282);
xnor U535 (N_535,In_748,In_325);
nor U536 (N_536,In_149,In_609);
nor U537 (N_537,In_541,In_141);
and U538 (N_538,In_353,In_321);
nand U539 (N_539,In_246,In_713);
nand U540 (N_540,In_453,In_532);
nor U541 (N_541,In_393,In_245);
and U542 (N_542,In_132,In_334);
and U543 (N_543,In_428,In_221);
nor U544 (N_544,In_416,In_28);
nor U545 (N_545,In_585,In_442);
nor U546 (N_546,In_33,In_518);
or U547 (N_547,In_392,In_321);
nor U548 (N_548,In_447,In_706);
or U549 (N_549,In_513,In_2);
or U550 (N_550,In_27,In_110);
or U551 (N_551,In_269,In_124);
and U552 (N_552,In_219,In_93);
nor U553 (N_553,In_193,In_384);
nor U554 (N_554,In_664,In_217);
and U555 (N_555,In_527,In_612);
and U556 (N_556,In_168,In_393);
nand U557 (N_557,In_551,In_18);
nand U558 (N_558,In_525,In_23);
or U559 (N_559,In_540,In_654);
or U560 (N_560,In_681,In_31);
nor U561 (N_561,In_570,In_174);
and U562 (N_562,In_710,In_466);
and U563 (N_563,In_719,In_214);
nor U564 (N_564,In_598,In_328);
xnor U565 (N_565,In_545,In_226);
or U566 (N_566,In_591,In_510);
and U567 (N_567,In_476,In_381);
and U568 (N_568,In_535,In_628);
or U569 (N_569,In_34,In_676);
or U570 (N_570,In_242,In_540);
nor U571 (N_571,In_241,In_669);
xor U572 (N_572,In_8,In_369);
nor U573 (N_573,In_342,In_22);
or U574 (N_574,In_121,In_201);
nor U575 (N_575,In_301,In_113);
and U576 (N_576,In_49,In_261);
nand U577 (N_577,In_100,In_283);
xor U578 (N_578,In_623,In_258);
nor U579 (N_579,In_245,In_47);
and U580 (N_580,In_417,In_180);
or U581 (N_581,In_97,In_669);
or U582 (N_582,In_564,In_162);
nor U583 (N_583,In_68,In_338);
nand U584 (N_584,In_223,In_120);
or U585 (N_585,In_379,In_242);
xor U586 (N_586,In_322,In_76);
or U587 (N_587,In_739,In_523);
and U588 (N_588,In_195,In_279);
or U589 (N_589,In_643,In_448);
nand U590 (N_590,In_591,In_513);
and U591 (N_591,In_549,In_477);
and U592 (N_592,In_549,In_171);
or U593 (N_593,In_165,In_431);
nor U594 (N_594,In_81,In_387);
nand U595 (N_595,In_67,In_387);
or U596 (N_596,In_492,In_535);
nor U597 (N_597,In_36,In_677);
and U598 (N_598,In_345,In_187);
or U599 (N_599,In_188,In_65);
and U600 (N_600,In_78,In_622);
nand U601 (N_601,In_509,In_269);
and U602 (N_602,In_336,In_562);
nand U603 (N_603,In_284,In_105);
or U604 (N_604,In_736,In_234);
nor U605 (N_605,In_390,In_690);
nand U606 (N_606,In_673,In_220);
nand U607 (N_607,In_441,In_53);
and U608 (N_608,In_66,In_99);
and U609 (N_609,In_231,In_270);
nor U610 (N_610,In_480,In_688);
nor U611 (N_611,In_212,In_123);
or U612 (N_612,In_623,In_167);
and U613 (N_613,In_633,In_126);
nand U614 (N_614,In_205,In_207);
or U615 (N_615,In_199,In_380);
nand U616 (N_616,In_676,In_749);
and U617 (N_617,In_132,In_297);
and U618 (N_618,In_32,In_405);
nor U619 (N_619,In_209,In_490);
and U620 (N_620,In_301,In_511);
and U621 (N_621,In_545,In_232);
xnor U622 (N_622,In_99,In_116);
nand U623 (N_623,In_1,In_446);
and U624 (N_624,In_373,In_68);
and U625 (N_625,In_20,In_730);
or U626 (N_626,In_562,In_520);
nor U627 (N_627,In_236,In_537);
or U628 (N_628,In_289,In_417);
and U629 (N_629,In_436,In_666);
xnor U630 (N_630,In_384,In_608);
and U631 (N_631,In_362,In_551);
nand U632 (N_632,In_15,In_169);
nor U633 (N_633,In_240,In_291);
nand U634 (N_634,In_746,In_216);
and U635 (N_635,In_24,In_511);
or U636 (N_636,In_463,In_92);
nor U637 (N_637,In_164,In_268);
or U638 (N_638,In_723,In_40);
or U639 (N_639,In_331,In_265);
nor U640 (N_640,In_279,In_611);
and U641 (N_641,In_342,In_78);
nand U642 (N_642,In_560,In_615);
nand U643 (N_643,In_658,In_154);
nor U644 (N_644,In_215,In_349);
and U645 (N_645,In_684,In_679);
and U646 (N_646,In_197,In_587);
or U647 (N_647,In_736,In_168);
or U648 (N_648,In_537,In_659);
nand U649 (N_649,In_155,In_630);
or U650 (N_650,In_199,In_357);
nor U651 (N_651,In_353,In_625);
or U652 (N_652,In_207,In_638);
nand U653 (N_653,In_235,In_201);
nand U654 (N_654,In_78,In_662);
nor U655 (N_655,In_409,In_258);
nand U656 (N_656,In_359,In_391);
or U657 (N_657,In_655,In_600);
xnor U658 (N_658,In_481,In_60);
nand U659 (N_659,In_623,In_443);
or U660 (N_660,In_632,In_116);
nand U661 (N_661,In_359,In_612);
and U662 (N_662,In_384,In_80);
nor U663 (N_663,In_170,In_238);
xnor U664 (N_664,In_411,In_542);
nand U665 (N_665,In_518,In_148);
and U666 (N_666,In_675,In_687);
or U667 (N_667,In_186,In_529);
or U668 (N_668,In_543,In_622);
nor U669 (N_669,In_103,In_228);
nor U670 (N_670,In_701,In_128);
and U671 (N_671,In_584,In_162);
or U672 (N_672,In_0,In_8);
nand U673 (N_673,In_504,In_421);
and U674 (N_674,In_76,In_278);
and U675 (N_675,In_187,In_566);
nand U676 (N_676,In_341,In_486);
nor U677 (N_677,In_355,In_693);
nor U678 (N_678,In_432,In_514);
nor U679 (N_679,In_209,In_593);
and U680 (N_680,In_203,In_396);
and U681 (N_681,In_238,In_603);
or U682 (N_682,In_272,In_479);
nor U683 (N_683,In_695,In_660);
and U684 (N_684,In_364,In_409);
or U685 (N_685,In_725,In_142);
nor U686 (N_686,In_245,In_655);
nor U687 (N_687,In_534,In_389);
or U688 (N_688,In_594,In_749);
or U689 (N_689,In_212,In_143);
nand U690 (N_690,In_444,In_150);
nand U691 (N_691,In_197,In_643);
and U692 (N_692,In_307,In_265);
nand U693 (N_693,In_1,In_58);
and U694 (N_694,In_585,In_509);
or U695 (N_695,In_562,In_181);
nand U696 (N_696,In_73,In_506);
nand U697 (N_697,In_277,In_100);
xnor U698 (N_698,In_137,In_241);
nor U699 (N_699,In_691,In_1);
and U700 (N_700,In_547,In_359);
and U701 (N_701,In_409,In_740);
nand U702 (N_702,In_634,In_656);
nor U703 (N_703,In_18,In_616);
nand U704 (N_704,In_397,In_504);
and U705 (N_705,In_662,In_727);
and U706 (N_706,In_338,In_198);
nor U707 (N_707,In_11,In_482);
nand U708 (N_708,In_684,In_340);
nand U709 (N_709,In_364,In_192);
nor U710 (N_710,In_90,In_466);
nand U711 (N_711,In_667,In_256);
or U712 (N_712,In_308,In_438);
and U713 (N_713,In_628,In_569);
nor U714 (N_714,In_291,In_230);
nor U715 (N_715,In_138,In_524);
nor U716 (N_716,In_272,In_359);
nor U717 (N_717,In_634,In_425);
nor U718 (N_718,In_380,In_410);
xor U719 (N_719,In_358,In_473);
nand U720 (N_720,In_7,In_108);
nor U721 (N_721,In_709,In_559);
and U722 (N_722,In_686,In_62);
nand U723 (N_723,In_668,In_351);
or U724 (N_724,In_632,In_159);
nand U725 (N_725,In_286,In_127);
nand U726 (N_726,In_337,In_356);
and U727 (N_727,In_209,In_535);
or U728 (N_728,In_605,In_469);
or U729 (N_729,In_698,In_538);
or U730 (N_730,In_163,In_412);
and U731 (N_731,In_680,In_549);
xor U732 (N_732,In_631,In_633);
and U733 (N_733,In_498,In_382);
and U734 (N_734,In_237,In_600);
nand U735 (N_735,In_551,In_69);
and U736 (N_736,In_222,In_457);
nor U737 (N_737,In_282,In_374);
nor U738 (N_738,In_533,In_70);
nand U739 (N_739,In_163,In_719);
and U740 (N_740,In_135,In_508);
and U741 (N_741,In_250,In_218);
and U742 (N_742,In_119,In_364);
nor U743 (N_743,In_728,In_336);
nor U744 (N_744,In_722,In_735);
or U745 (N_745,In_551,In_709);
or U746 (N_746,In_501,In_322);
nand U747 (N_747,In_686,In_611);
nor U748 (N_748,In_393,In_420);
or U749 (N_749,In_597,In_506);
or U750 (N_750,In_449,In_679);
nor U751 (N_751,In_329,In_450);
nor U752 (N_752,In_406,In_91);
or U753 (N_753,In_41,In_465);
nand U754 (N_754,In_145,In_111);
or U755 (N_755,In_332,In_661);
nor U756 (N_756,In_76,In_339);
or U757 (N_757,In_187,In_447);
nor U758 (N_758,In_501,In_599);
and U759 (N_759,In_140,In_745);
nor U760 (N_760,In_129,In_747);
or U761 (N_761,In_616,In_41);
nand U762 (N_762,In_164,In_128);
and U763 (N_763,In_195,In_524);
or U764 (N_764,In_474,In_716);
or U765 (N_765,In_428,In_573);
nand U766 (N_766,In_99,In_189);
or U767 (N_767,In_60,In_681);
nor U768 (N_768,In_130,In_106);
or U769 (N_769,In_366,In_74);
or U770 (N_770,In_28,In_159);
or U771 (N_771,In_233,In_83);
nor U772 (N_772,In_458,In_720);
and U773 (N_773,In_679,In_109);
and U774 (N_774,In_682,In_255);
nand U775 (N_775,In_158,In_677);
nor U776 (N_776,In_625,In_712);
and U777 (N_777,In_396,In_662);
nand U778 (N_778,In_152,In_174);
nor U779 (N_779,In_603,In_132);
nand U780 (N_780,In_268,In_696);
or U781 (N_781,In_581,In_29);
and U782 (N_782,In_731,In_192);
or U783 (N_783,In_297,In_261);
nand U784 (N_784,In_285,In_228);
or U785 (N_785,In_377,In_670);
nand U786 (N_786,In_57,In_512);
nand U787 (N_787,In_376,In_487);
nor U788 (N_788,In_525,In_713);
and U789 (N_789,In_569,In_369);
nand U790 (N_790,In_90,In_53);
and U791 (N_791,In_294,In_145);
nand U792 (N_792,In_38,In_455);
nor U793 (N_793,In_94,In_239);
nand U794 (N_794,In_671,In_527);
or U795 (N_795,In_440,In_123);
xor U796 (N_796,In_126,In_281);
nand U797 (N_797,In_355,In_430);
or U798 (N_798,In_186,In_343);
and U799 (N_799,In_379,In_61);
and U800 (N_800,In_101,In_627);
or U801 (N_801,In_477,In_638);
nand U802 (N_802,In_289,In_263);
or U803 (N_803,In_492,In_730);
or U804 (N_804,In_312,In_437);
nor U805 (N_805,In_135,In_271);
nand U806 (N_806,In_459,In_682);
and U807 (N_807,In_43,In_413);
nand U808 (N_808,In_286,In_382);
xnor U809 (N_809,In_62,In_173);
nand U810 (N_810,In_589,In_169);
nand U811 (N_811,In_10,In_287);
nor U812 (N_812,In_267,In_722);
nand U813 (N_813,In_634,In_394);
nor U814 (N_814,In_238,In_50);
nand U815 (N_815,In_479,In_438);
xor U816 (N_816,In_706,In_510);
and U817 (N_817,In_264,In_247);
or U818 (N_818,In_15,In_355);
or U819 (N_819,In_310,In_486);
nor U820 (N_820,In_124,In_635);
and U821 (N_821,In_346,In_363);
or U822 (N_822,In_195,In_586);
nand U823 (N_823,In_368,In_341);
or U824 (N_824,In_605,In_82);
and U825 (N_825,In_490,In_213);
nand U826 (N_826,In_392,In_279);
xnor U827 (N_827,In_310,In_165);
nand U828 (N_828,In_300,In_707);
or U829 (N_829,In_633,In_636);
nor U830 (N_830,In_190,In_328);
and U831 (N_831,In_648,In_704);
nor U832 (N_832,In_580,In_596);
nor U833 (N_833,In_49,In_416);
nor U834 (N_834,In_262,In_218);
nand U835 (N_835,In_474,In_153);
nand U836 (N_836,In_701,In_583);
or U837 (N_837,In_288,In_301);
nor U838 (N_838,In_691,In_24);
nand U839 (N_839,In_719,In_347);
xor U840 (N_840,In_486,In_386);
nand U841 (N_841,In_606,In_174);
nand U842 (N_842,In_256,In_428);
and U843 (N_843,In_469,In_673);
and U844 (N_844,In_722,In_719);
nor U845 (N_845,In_423,In_31);
nand U846 (N_846,In_288,In_281);
or U847 (N_847,In_327,In_675);
nand U848 (N_848,In_80,In_58);
nand U849 (N_849,In_339,In_61);
nand U850 (N_850,In_313,In_399);
and U851 (N_851,In_284,In_382);
xor U852 (N_852,In_718,In_264);
and U853 (N_853,In_499,In_246);
nand U854 (N_854,In_678,In_379);
and U855 (N_855,In_484,In_338);
nand U856 (N_856,In_88,In_608);
and U857 (N_857,In_223,In_533);
nand U858 (N_858,In_74,In_440);
and U859 (N_859,In_498,In_270);
nor U860 (N_860,In_19,In_477);
nor U861 (N_861,In_646,In_19);
nor U862 (N_862,In_446,In_184);
nor U863 (N_863,In_154,In_249);
nor U864 (N_864,In_238,In_179);
nand U865 (N_865,In_319,In_508);
nand U866 (N_866,In_321,In_83);
and U867 (N_867,In_221,In_679);
xnor U868 (N_868,In_57,In_399);
or U869 (N_869,In_566,In_307);
nand U870 (N_870,In_163,In_132);
nand U871 (N_871,In_343,In_64);
nand U872 (N_872,In_305,In_278);
or U873 (N_873,In_193,In_17);
nor U874 (N_874,In_61,In_167);
nand U875 (N_875,In_589,In_70);
or U876 (N_876,In_596,In_653);
xor U877 (N_877,In_703,In_175);
nand U878 (N_878,In_694,In_264);
nor U879 (N_879,In_128,In_202);
nand U880 (N_880,In_229,In_299);
or U881 (N_881,In_632,In_521);
and U882 (N_882,In_124,In_14);
nand U883 (N_883,In_402,In_685);
nor U884 (N_884,In_591,In_114);
or U885 (N_885,In_49,In_100);
nor U886 (N_886,In_293,In_426);
or U887 (N_887,In_647,In_284);
or U888 (N_888,In_270,In_545);
and U889 (N_889,In_213,In_269);
or U890 (N_890,In_605,In_87);
or U891 (N_891,In_67,In_745);
nor U892 (N_892,In_96,In_690);
nor U893 (N_893,In_206,In_90);
nand U894 (N_894,In_182,In_694);
nor U895 (N_895,In_20,In_207);
nand U896 (N_896,In_288,In_602);
nor U897 (N_897,In_270,In_650);
or U898 (N_898,In_57,In_243);
nand U899 (N_899,In_746,In_540);
or U900 (N_900,In_502,In_501);
or U901 (N_901,In_146,In_628);
and U902 (N_902,In_555,In_234);
nor U903 (N_903,In_497,In_322);
nand U904 (N_904,In_471,In_370);
and U905 (N_905,In_127,In_575);
nor U906 (N_906,In_338,In_360);
and U907 (N_907,In_104,In_89);
nand U908 (N_908,In_637,In_138);
or U909 (N_909,In_625,In_500);
nor U910 (N_910,In_246,In_690);
nand U911 (N_911,In_435,In_201);
or U912 (N_912,In_534,In_508);
or U913 (N_913,In_142,In_604);
or U914 (N_914,In_414,In_671);
nand U915 (N_915,In_177,In_280);
and U916 (N_916,In_430,In_353);
or U917 (N_917,In_288,In_580);
nor U918 (N_918,In_610,In_92);
nand U919 (N_919,In_136,In_505);
nor U920 (N_920,In_400,In_599);
nand U921 (N_921,In_736,In_684);
xor U922 (N_922,In_578,In_109);
or U923 (N_923,In_458,In_58);
nand U924 (N_924,In_711,In_61);
and U925 (N_925,In_199,In_100);
nor U926 (N_926,In_738,In_512);
nor U927 (N_927,In_27,In_627);
and U928 (N_928,In_527,In_167);
and U929 (N_929,In_416,In_351);
and U930 (N_930,In_460,In_461);
or U931 (N_931,In_473,In_525);
and U932 (N_932,In_661,In_705);
nor U933 (N_933,In_625,In_314);
nand U934 (N_934,In_128,In_451);
and U935 (N_935,In_491,In_586);
and U936 (N_936,In_466,In_220);
nand U937 (N_937,In_241,In_417);
xor U938 (N_938,In_597,In_141);
or U939 (N_939,In_557,In_169);
nand U940 (N_940,In_709,In_239);
and U941 (N_941,In_568,In_536);
and U942 (N_942,In_635,In_659);
and U943 (N_943,In_697,In_122);
nand U944 (N_944,In_472,In_468);
nand U945 (N_945,In_194,In_643);
or U946 (N_946,In_70,In_146);
or U947 (N_947,In_397,In_499);
nand U948 (N_948,In_577,In_533);
nand U949 (N_949,In_418,In_666);
nand U950 (N_950,In_587,In_688);
nor U951 (N_951,In_154,In_17);
nor U952 (N_952,In_440,In_701);
and U953 (N_953,In_470,In_10);
and U954 (N_954,In_242,In_370);
nand U955 (N_955,In_601,In_578);
nor U956 (N_956,In_180,In_510);
nor U957 (N_957,In_250,In_728);
and U958 (N_958,In_383,In_407);
nand U959 (N_959,In_544,In_15);
nand U960 (N_960,In_1,In_270);
or U961 (N_961,In_339,In_605);
nor U962 (N_962,In_9,In_652);
and U963 (N_963,In_121,In_290);
or U964 (N_964,In_385,In_481);
nand U965 (N_965,In_458,In_672);
or U966 (N_966,In_196,In_181);
and U967 (N_967,In_680,In_124);
or U968 (N_968,In_675,In_354);
nor U969 (N_969,In_191,In_627);
or U970 (N_970,In_180,In_452);
or U971 (N_971,In_478,In_528);
nand U972 (N_972,In_490,In_249);
nor U973 (N_973,In_404,In_444);
nor U974 (N_974,In_481,In_148);
or U975 (N_975,In_545,In_244);
nor U976 (N_976,In_361,In_590);
and U977 (N_977,In_223,In_183);
nor U978 (N_978,In_487,In_90);
or U979 (N_979,In_367,In_148);
nand U980 (N_980,In_417,In_35);
nand U981 (N_981,In_365,In_697);
nor U982 (N_982,In_159,In_705);
nor U983 (N_983,In_279,In_312);
nand U984 (N_984,In_671,In_469);
and U985 (N_985,In_504,In_627);
and U986 (N_986,In_224,In_168);
or U987 (N_987,In_444,In_684);
nand U988 (N_988,In_549,In_117);
or U989 (N_989,In_102,In_582);
and U990 (N_990,In_299,In_616);
nand U991 (N_991,In_701,In_392);
or U992 (N_992,In_648,In_583);
or U993 (N_993,In_26,In_323);
nor U994 (N_994,In_555,In_123);
and U995 (N_995,In_135,In_570);
nand U996 (N_996,In_599,In_243);
or U997 (N_997,In_142,In_42);
and U998 (N_998,In_571,In_124);
nor U999 (N_999,In_246,In_39);
and U1000 (N_1000,In_494,In_625);
xnor U1001 (N_1001,In_733,In_578);
nor U1002 (N_1002,In_386,In_490);
nor U1003 (N_1003,In_468,In_21);
nor U1004 (N_1004,In_715,In_633);
and U1005 (N_1005,In_13,In_451);
and U1006 (N_1006,In_701,In_560);
or U1007 (N_1007,In_148,In_215);
or U1008 (N_1008,In_194,In_209);
nand U1009 (N_1009,In_195,In_694);
and U1010 (N_1010,In_682,In_688);
nor U1011 (N_1011,In_438,In_329);
or U1012 (N_1012,In_375,In_270);
nor U1013 (N_1013,In_356,In_449);
nand U1014 (N_1014,In_147,In_485);
nor U1015 (N_1015,In_603,In_280);
nor U1016 (N_1016,In_725,In_634);
or U1017 (N_1017,In_329,In_84);
and U1018 (N_1018,In_165,In_619);
nand U1019 (N_1019,In_130,In_664);
or U1020 (N_1020,In_250,In_454);
nor U1021 (N_1021,In_198,In_371);
or U1022 (N_1022,In_121,In_114);
nor U1023 (N_1023,In_486,In_402);
nor U1024 (N_1024,In_103,In_396);
and U1025 (N_1025,In_720,In_519);
nand U1026 (N_1026,In_219,In_113);
and U1027 (N_1027,In_552,In_623);
or U1028 (N_1028,In_331,In_529);
nand U1029 (N_1029,In_58,In_467);
or U1030 (N_1030,In_602,In_306);
and U1031 (N_1031,In_39,In_158);
or U1032 (N_1032,In_725,In_486);
and U1033 (N_1033,In_29,In_553);
nor U1034 (N_1034,In_15,In_417);
and U1035 (N_1035,In_556,In_86);
and U1036 (N_1036,In_316,In_216);
or U1037 (N_1037,In_107,In_701);
and U1038 (N_1038,In_682,In_421);
nand U1039 (N_1039,In_390,In_718);
nor U1040 (N_1040,In_583,In_542);
and U1041 (N_1041,In_463,In_578);
nor U1042 (N_1042,In_668,In_148);
or U1043 (N_1043,In_555,In_382);
or U1044 (N_1044,In_331,In_24);
xor U1045 (N_1045,In_224,In_563);
nand U1046 (N_1046,In_634,In_76);
nor U1047 (N_1047,In_324,In_708);
or U1048 (N_1048,In_376,In_240);
or U1049 (N_1049,In_107,In_253);
or U1050 (N_1050,In_574,In_546);
and U1051 (N_1051,In_158,In_291);
and U1052 (N_1052,In_642,In_82);
and U1053 (N_1053,In_290,In_601);
nand U1054 (N_1054,In_705,In_199);
or U1055 (N_1055,In_148,In_76);
nor U1056 (N_1056,In_655,In_115);
or U1057 (N_1057,In_601,In_488);
nor U1058 (N_1058,In_408,In_432);
nor U1059 (N_1059,In_22,In_30);
or U1060 (N_1060,In_424,In_94);
or U1061 (N_1061,In_447,In_29);
or U1062 (N_1062,In_146,In_481);
nor U1063 (N_1063,In_281,In_451);
xor U1064 (N_1064,In_492,In_209);
or U1065 (N_1065,In_527,In_488);
and U1066 (N_1066,In_312,In_529);
nor U1067 (N_1067,In_445,In_114);
and U1068 (N_1068,In_254,In_34);
or U1069 (N_1069,In_45,In_587);
nand U1070 (N_1070,In_630,In_377);
or U1071 (N_1071,In_140,In_629);
or U1072 (N_1072,In_676,In_597);
nand U1073 (N_1073,In_120,In_208);
or U1074 (N_1074,In_218,In_556);
xor U1075 (N_1075,In_306,In_359);
and U1076 (N_1076,In_240,In_248);
nand U1077 (N_1077,In_280,In_168);
nand U1078 (N_1078,In_329,In_270);
xor U1079 (N_1079,In_663,In_187);
and U1080 (N_1080,In_470,In_614);
nor U1081 (N_1081,In_472,In_542);
nor U1082 (N_1082,In_3,In_444);
or U1083 (N_1083,In_518,In_499);
nand U1084 (N_1084,In_119,In_621);
xor U1085 (N_1085,In_177,In_667);
nand U1086 (N_1086,In_38,In_49);
and U1087 (N_1087,In_98,In_625);
xnor U1088 (N_1088,In_86,In_14);
or U1089 (N_1089,In_449,In_287);
and U1090 (N_1090,In_589,In_722);
and U1091 (N_1091,In_534,In_136);
nor U1092 (N_1092,In_359,In_55);
and U1093 (N_1093,In_424,In_605);
or U1094 (N_1094,In_466,In_508);
or U1095 (N_1095,In_90,In_428);
nor U1096 (N_1096,In_61,In_578);
nand U1097 (N_1097,In_687,In_396);
nand U1098 (N_1098,In_157,In_256);
nand U1099 (N_1099,In_277,In_139);
and U1100 (N_1100,In_386,In_563);
nor U1101 (N_1101,In_100,In_391);
nor U1102 (N_1102,In_535,In_173);
nand U1103 (N_1103,In_243,In_658);
nand U1104 (N_1104,In_522,In_404);
nand U1105 (N_1105,In_607,In_577);
and U1106 (N_1106,In_737,In_699);
nand U1107 (N_1107,In_117,In_214);
nand U1108 (N_1108,In_20,In_298);
nor U1109 (N_1109,In_161,In_687);
or U1110 (N_1110,In_141,In_661);
nor U1111 (N_1111,In_437,In_6);
or U1112 (N_1112,In_382,In_19);
nand U1113 (N_1113,In_674,In_163);
nand U1114 (N_1114,In_273,In_674);
or U1115 (N_1115,In_638,In_400);
nor U1116 (N_1116,In_407,In_419);
and U1117 (N_1117,In_544,In_210);
nand U1118 (N_1118,In_404,In_40);
or U1119 (N_1119,In_51,In_163);
xor U1120 (N_1120,In_105,In_285);
or U1121 (N_1121,In_307,In_181);
and U1122 (N_1122,In_566,In_502);
and U1123 (N_1123,In_510,In_661);
and U1124 (N_1124,In_595,In_328);
nand U1125 (N_1125,In_452,In_517);
nand U1126 (N_1126,In_419,In_715);
nor U1127 (N_1127,In_44,In_372);
nor U1128 (N_1128,In_595,In_707);
nand U1129 (N_1129,In_59,In_374);
nand U1130 (N_1130,In_626,In_13);
and U1131 (N_1131,In_478,In_349);
nor U1132 (N_1132,In_491,In_740);
or U1133 (N_1133,In_638,In_518);
and U1134 (N_1134,In_625,In_337);
or U1135 (N_1135,In_272,In_656);
and U1136 (N_1136,In_164,In_34);
and U1137 (N_1137,In_322,In_351);
nor U1138 (N_1138,In_19,In_593);
nand U1139 (N_1139,In_159,In_732);
and U1140 (N_1140,In_530,In_143);
nand U1141 (N_1141,In_514,In_301);
and U1142 (N_1142,In_587,In_222);
nor U1143 (N_1143,In_207,In_156);
nor U1144 (N_1144,In_169,In_168);
xor U1145 (N_1145,In_196,In_264);
and U1146 (N_1146,In_521,In_452);
or U1147 (N_1147,In_346,In_679);
nor U1148 (N_1148,In_82,In_217);
or U1149 (N_1149,In_380,In_286);
or U1150 (N_1150,In_372,In_97);
nand U1151 (N_1151,In_707,In_463);
nand U1152 (N_1152,In_535,In_4);
or U1153 (N_1153,In_160,In_525);
nand U1154 (N_1154,In_221,In_246);
or U1155 (N_1155,In_420,In_709);
or U1156 (N_1156,In_307,In_422);
nor U1157 (N_1157,In_620,In_208);
nor U1158 (N_1158,In_728,In_465);
and U1159 (N_1159,In_280,In_486);
and U1160 (N_1160,In_295,In_621);
or U1161 (N_1161,In_280,In_236);
nand U1162 (N_1162,In_16,In_563);
xnor U1163 (N_1163,In_682,In_661);
nand U1164 (N_1164,In_101,In_329);
or U1165 (N_1165,In_168,In_240);
or U1166 (N_1166,In_80,In_561);
nand U1167 (N_1167,In_643,In_409);
and U1168 (N_1168,In_718,In_460);
nor U1169 (N_1169,In_330,In_729);
or U1170 (N_1170,In_657,In_438);
or U1171 (N_1171,In_622,In_359);
or U1172 (N_1172,In_221,In_197);
nand U1173 (N_1173,In_655,In_157);
or U1174 (N_1174,In_695,In_595);
nand U1175 (N_1175,In_593,In_21);
or U1176 (N_1176,In_389,In_591);
and U1177 (N_1177,In_274,In_395);
nand U1178 (N_1178,In_652,In_545);
nand U1179 (N_1179,In_715,In_46);
or U1180 (N_1180,In_107,In_715);
or U1181 (N_1181,In_73,In_134);
or U1182 (N_1182,In_213,In_105);
nor U1183 (N_1183,In_627,In_50);
and U1184 (N_1184,In_660,In_490);
nand U1185 (N_1185,In_290,In_732);
nand U1186 (N_1186,In_418,In_22);
nor U1187 (N_1187,In_591,In_649);
nor U1188 (N_1188,In_742,In_402);
nor U1189 (N_1189,In_65,In_374);
or U1190 (N_1190,In_555,In_453);
nand U1191 (N_1191,In_221,In_721);
or U1192 (N_1192,In_720,In_11);
nand U1193 (N_1193,In_71,In_600);
nand U1194 (N_1194,In_594,In_29);
nor U1195 (N_1195,In_703,In_735);
nor U1196 (N_1196,In_748,In_71);
and U1197 (N_1197,In_578,In_683);
and U1198 (N_1198,In_181,In_259);
nor U1199 (N_1199,In_156,In_724);
nor U1200 (N_1200,In_130,In_412);
and U1201 (N_1201,In_410,In_337);
and U1202 (N_1202,In_45,In_547);
and U1203 (N_1203,In_700,In_63);
nor U1204 (N_1204,In_50,In_562);
and U1205 (N_1205,In_724,In_297);
nor U1206 (N_1206,In_237,In_479);
xnor U1207 (N_1207,In_657,In_298);
and U1208 (N_1208,In_488,In_83);
and U1209 (N_1209,In_245,In_460);
nor U1210 (N_1210,In_721,In_102);
nor U1211 (N_1211,In_216,In_380);
or U1212 (N_1212,In_377,In_306);
or U1213 (N_1213,In_151,In_515);
and U1214 (N_1214,In_515,In_153);
and U1215 (N_1215,In_303,In_236);
and U1216 (N_1216,In_0,In_160);
nand U1217 (N_1217,In_691,In_683);
xnor U1218 (N_1218,In_491,In_652);
nand U1219 (N_1219,In_42,In_298);
nand U1220 (N_1220,In_162,In_264);
nor U1221 (N_1221,In_258,In_692);
nand U1222 (N_1222,In_156,In_496);
nand U1223 (N_1223,In_497,In_728);
nor U1224 (N_1224,In_580,In_34);
or U1225 (N_1225,In_602,In_385);
nand U1226 (N_1226,In_29,In_175);
nor U1227 (N_1227,In_317,In_275);
nor U1228 (N_1228,In_491,In_617);
and U1229 (N_1229,In_738,In_652);
nor U1230 (N_1230,In_498,In_684);
nor U1231 (N_1231,In_209,In_436);
or U1232 (N_1232,In_588,In_262);
nand U1233 (N_1233,In_500,In_394);
and U1234 (N_1234,In_600,In_472);
or U1235 (N_1235,In_570,In_484);
or U1236 (N_1236,In_324,In_116);
nand U1237 (N_1237,In_539,In_410);
and U1238 (N_1238,In_434,In_662);
and U1239 (N_1239,In_230,In_170);
nand U1240 (N_1240,In_663,In_407);
and U1241 (N_1241,In_655,In_152);
or U1242 (N_1242,In_368,In_749);
or U1243 (N_1243,In_179,In_360);
nor U1244 (N_1244,In_83,In_574);
and U1245 (N_1245,In_368,In_57);
or U1246 (N_1246,In_18,In_441);
or U1247 (N_1247,In_2,In_291);
nand U1248 (N_1248,In_549,In_419);
or U1249 (N_1249,In_521,In_343);
nor U1250 (N_1250,In_470,In_661);
or U1251 (N_1251,In_330,In_499);
or U1252 (N_1252,In_490,In_190);
nor U1253 (N_1253,In_723,In_508);
and U1254 (N_1254,In_516,In_219);
and U1255 (N_1255,In_337,In_307);
nor U1256 (N_1256,In_538,In_581);
nor U1257 (N_1257,In_492,In_183);
and U1258 (N_1258,In_654,In_342);
and U1259 (N_1259,In_745,In_452);
nor U1260 (N_1260,In_358,In_148);
or U1261 (N_1261,In_339,In_355);
nand U1262 (N_1262,In_112,In_385);
or U1263 (N_1263,In_359,In_423);
or U1264 (N_1264,In_706,In_164);
and U1265 (N_1265,In_243,In_391);
nor U1266 (N_1266,In_543,In_736);
or U1267 (N_1267,In_57,In_304);
nand U1268 (N_1268,In_243,In_367);
or U1269 (N_1269,In_280,In_241);
nor U1270 (N_1270,In_260,In_607);
nand U1271 (N_1271,In_92,In_36);
nor U1272 (N_1272,In_539,In_218);
nor U1273 (N_1273,In_155,In_281);
nand U1274 (N_1274,In_470,In_300);
xnor U1275 (N_1275,In_282,In_410);
xnor U1276 (N_1276,In_732,In_584);
nand U1277 (N_1277,In_677,In_514);
and U1278 (N_1278,In_460,In_478);
or U1279 (N_1279,In_451,In_532);
and U1280 (N_1280,In_653,In_642);
and U1281 (N_1281,In_154,In_204);
and U1282 (N_1282,In_292,In_520);
nor U1283 (N_1283,In_325,In_307);
or U1284 (N_1284,In_386,In_37);
nand U1285 (N_1285,In_437,In_601);
and U1286 (N_1286,In_156,In_202);
and U1287 (N_1287,In_535,In_186);
nand U1288 (N_1288,In_211,In_524);
nor U1289 (N_1289,In_204,In_622);
and U1290 (N_1290,In_522,In_733);
nor U1291 (N_1291,In_639,In_285);
and U1292 (N_1292,In_645,In_488);
or U1293 (N_1293,In_617,In_22);
and U1294 (N_1294,In_112,In_100);
nand U1295 (N_1295,In_525,In_203);
or U1296 (N_1296,In_685,In_457);
nor U1297 (N_1297,In_352,In_160);
nor U1298 (N_1298,In_304,In_464);
nand U1299 (N_1299,In_219,In_507);
or U1300 (N_1300,In_54,In_33);
xor U1301 (N_1301,In_254,In_577);
nand U1302 (N_1302,In_170,In_406);
or U1303 (N_1303,In_719,In_90);
or U1304 (N_1304,In_389,In_338);
or U1305 (N_1305,In_226,In_633);
nor U1306 (N_1306,In_273,In_743);
and U1307 (N_1307,In_191,In_582);
nand U1308 (N_1308,In_356,In_640);
nand U1309 (N_1309,In_469,In_672);
nor U1310 (N_1310,In_332,In_455);
nor U1311 (N_1311,In_683,In_556);
nor U1312 (N_1312,In_232,In_214);
nand U1313 (N_1313,In_667,In_713);
nand U1314 (N_1314,In_222,In_679);
or U1315 (N_1315,In_450,In_260);
or U1316 (N_1316,In_654,In_534);
nand U1317 (N_1317,In_212,In_691);
xor U1318 (N_1318,In_293,In_348);
or U1319 (N_1319,In_548,In_213);
xor U1320 (N_1320,In_82,In_644);
or U1321 (N_1321,In_243,In_504);
and U1322 (N_1322,In_539,In_21);
or U1323 (N_1323,In_272,In_185);
or U1324 (N_1324,In_200,In_25);
nor U1325 (N_1325,In_749,In_331);
or U1326 (N_1326,In_319,In_192);
or U1327 (N_1327,In_169,In_66);
and U1328 (N_1328,In_524,In_264);
and U1329 (N_1329,In_718,In_652);
nor U1330 (N_1330,In_33,In_728);
nor U1331 (N_1331,In_518,In_390);
nand U1332 (N_1332,In_80,In_601);
or U1333 (N_1333,In_154,In_524);
nand U1334 (N_1334,In_130,In_44);
and U1335 (N_1335,In_658,In_261);
nor U1336 (N_1336,In_407,In_707);
xor U1337 (N_1337,In_502,In_497);
nand U1338 (N_1338,In_451,In_261);
and U1339 (N_1339,In_127,In_167);
or U1340 (N_1340,In_741,In_637);
or U1341 (N_1341,In_558,In_291);
nor U1342 (N_1342,In_190,In_411);
nand U1343 (N_1343,In_179,In_553);
nor U1344 (N_1344,In_446,In_241);
nand U1345 (N_1345,In_740,In_33);
and U1346 (N_1346,In_105,In_243);
or U1347 (N_1347,In_506,In_346);
or U1348 (N_1348,In_608,In_718);
nor U1349 (N_1349,In_482,In_32);
or U1350 (N_1350,In_438,In_609);
nor U1351 (N_1351,In_638,In_267);
nand U1352 (N_1352,In_125,In_436);
and U1353 (N_1353,In_442,In_397);
and U1354 (N_1354,In_453,In_23);
nand U1355 (N_1355,In_128,In_74);
nand U1356 (N_1356,In_147,In_675);
nand U1357 (N_1357,In_17,In_507);
nand U1358 (N_1358,In_537,In_610);
and U1359 (N_1359,In_17,In_713);
and U1360 (N_1360,In_593,In_566);
nand U1361 (N_1361,In_611,In_455);
and U1362 (N_1362,In_508,In_82);
and U1363 (N_1363,In_20,In_457);
nand U1364 (N_1364,In_415,In_727);
or U1365 (N_1365,In_719,In_378);
or U1366 (N_1366,In_666,In_294);
or U1367 (N_1367,In_321,In_513);
or U1368 (N_1368,In_704,In_100);
nor U1369 (N_1369,In_689,In_322);
or U1370 (N_1370,In_735,In_199);
or U1371 (N_1371,In_321,In_490);
and U1372 (N_1372,In_422,In_181);
or U1373 (N_1373,In_201,In_490);
nand U1374 (N_1374,In_456,In_143);
nand U1375 (N_1375,In_605,In_237);
nor U1376 (N_1376,In_479,In_209);
nand U1377 (N_1377,In_265,In_346);
and U1378 (N_1378,In_512,In_722);
nor U1379 (N_1379,In_629,In_589);
nor U1380 (N_1380,In_191,In_90);
nor U1381 (N_1381,In_165,In_410);
or U1382 (N_1382,In_310,In_454);
nor U1383 (N_1383,In_189,In_298);
and U1384 (N_1384,In_478,In_601);
and U1385 (N_1385,In_543,In_10);
and U1386 (N_1386,In_164,In_721);
and U1387 (N_1387,In_511,In_362);
nor U1388 (N_1388,In_577,In_743);
nor U1389 (N_1389,In_372,In_320);
nand U1390 (N_1390,In_520,In_318);
nor U1391 (N_1391,In_482,In_88);
and U1392 (N_1392,In_579,In_28);
and U1393 (N_1393,In_283,In_535);
nand U1394 (N_1394,In_372,In_587);
or U1395 (N_1395,In_374,In_229);
nand U1396 (N_1396,In_125,In_241);
and U1397 (N_1397,In_427,In_526);
or U1398 (N_1398,In_534,In_707);
and U1399 (N_1399,In_58,In_620);
and U1400 (N_1400,In_152,In_85);
nor U1401 (N_1401,In_557,In_331);
or U1402 (N_1402,In_272,In_630);
nand U1403 (N_1403,In_551,In_434);
and U1404 (N_1404,In_748,In_190);
nand U1405 (N_1405,In_712,In_161);
nor U1406 (N_1406,In_709,In_166);
or U1407 (N_1407,In_557,In_58);
and U1408 (N_1408,In_440,In_432);
nor U1409 (N_1409,In_411,In_361);
or U1410 (N_1410,In_27,In_305);
nor U1411 (N_1411,In_312,In_168);
nand U1412 (N_1412,In_213,In_22);
xor U1413 (N_1413,In_538,In_494);
nand U1414 (N_1414,In_492,In_605);
or U1415 (N_1415,In_125,In_130);
nor U1416 (N_1416,In_735,In_55);
or U1417 (N_1417,In_98,In_307);
and U1418 (N_1418,In_122,In_263);
or U1419 (N_1419,In_445,In_730);
or U1420 (N_1420,In_617,In_65);
nand U1421 (N_1421,In_513,In_383);
nand U1422 (N_1422,In_110,In_233);
nor U1423 (N_1423,In_133,In_492);
and U1424 (N_1424,In_548,In_449);
nand U1425 (N_1425,In_248,In_662);
nor U1426 (N_1426,In_72,In_274);
nor U1427 (N_1427,In_148,In_618);
nor U1428 (N_1428,In_399,In_701);
or U1429 (N_1429,In_599,In_396);
and U1430 (N_1430,In_472,In_438);
nor U1431 (N_1431,In_28,In_336);
nand U1432 (N_1432,In_573,In_76);
and U1433 (N_1433,In_621,In_692);
nor U1434 (N_1434,In_91,In_493);
nand U1435 (N_1435,In_256,In_303);
nor U1436 (N_1436,In_369,In_10);
or U1437 (N_1437,In_508,In_539);
nand U1438 (N_1438,In_442,In_363);
nand U1439 (N_1439,In_78,In_7);
nand U1440 (N_1440,In_405,In_489);
and U1441 (N_1441,In_667,In_106);
or U1442 (N_1442,In_322,In_668);
or U1443 (N_1443,In_491,In_686);
or U1444 (N_1444,In_246,In_132);
nor U1445 (N_1445,In_433,In_78);
nor U1446 (N_1446,In_7,In_576);
and U1447 (N_1447,In_728,In_242);
and U1448 (N_1448,In_567,In_591);
xnor U1449 (N_1449,In_82,In_431);
nor U1450 (N_1450,In_529,In_670);
or U1451 (N_1451,In_112,In_143);
xor U1452 (N_1452,In_516,In_281);
or U1453 (N_1453,In_249,In_707);
and U1454 (N_1454,In_740,In_28);
nor U1455 (N_1455,In_741,In_737);
nor U1456 (N_1456,In_335,In_457);
nand U1457 (N_1457,In_195,In_364);
nand U1458 (N_1458,In_744,In_67);
and U1459 (N_1459,In_58,In_51);
or U1460 (N_1460,In_596,In_528);
nor U1461 (N_1461,In_301,In_691);
nor U1462 (N_1462,In_430,In_662);
nand U1463 (N_1463,In_92,In_484);
nand U1464 (N_1464,In_443,In_694);
or U1465 (N_1465,In_271,In_176);
nor U1466 (N_1466,In_475,In_16);
nor U1467 (N_1467,In_722,In_108);
nor U1468 (N_1468,In_570,In_743);
and U1469 (N_1469,In_242,In_619);
nor U1470 (N_1470,In_218,In_37);
and U1471 (N_1471,In_663,In_506);
and U1472 (N_1472,In_201,In_58);
and U1473 (N_1473,In_178,In_214);
or U1474 (N_1474,In_380,In_212);
nand U1475 (N_1475,In_169,In_318);
or U1476 (N_1476,In_186,In_459);
nor U1477 (N_1477,In_644,In_359);
or U1478 (N_1478,In_366,In_642);
nor U1479 (N_1479,In_233,In_668);
or U1480 (N_1480,In_106,In_659);
nand U1481 (N_1481,In_412,In_328);
and U1482 (N_1482,In_363,In_661);
nand U1483 (N_1483,In_546,In_570);
nor U1484 (N_1484,In_169,In_120);
nor U1485 (N_1485,In_714,In_24);
nor U1486 (N_1486,In_419,In_184);
xor U1487 (N_1487,In_343,In_73);
nor U1488 (N_1488,In_317,In_383);
or U1489 (N_1489,In_256,In_228);
and U1490 (N_1490,In_284,In_338);
nand U1491 (N_1491,In_46,In_31);
and U1492 (N_1492,In_21,In_748);
or U1493 (N_1493,In_740,In_528);
nand U1494 (N_1494,In_612,In_315);
or U1495 (N_1495,In_699,In_431);
or U1496 (N_1496,In_427,In_159);
and U1497 (N_1497,In_726,In_342);
nor U1498 (N_1498,In_556,In_504);
and U1499 (N_1499,In_151,In_198);
nor U1500 (N_1500,In_408,In_51);
nand U1501 (N_1501,In_299,In_724);
and U1502 (N_1502,In_135,In_273);
nor U1503 (N_1503,In_677,In_529);
nor U1504 (N_1504,In_281,In_661);
nor U1505 (N_1505,In_509,In_383);
or U1506 (N_1506,In_410,In_184);
nor U1507 (N_1507,In_307,In_732);
and U1508 (N_1508,In_443,In_212);
and U1509 (N_1509,In_653,In_314);
nand U1510 (N_1510,In_362,In_606);
or U1511 (N_1511,In_745,In_73);
nand U1512 (N_1512,In_688,In_398);
nor U1513 (N_1513,In_483,In_643);
nor U1514 (N_1514,In_692,In_667);
nand U1515 (N_1515,In_680,In_17);
and U1516 (N_1516,In_165,In_338);
nand U1517 (N_1517,In_667,In_508);
or U1518 (N_1518,In_274,In_529);
or U1519 (N_1519,In_443,In_571);
nand U1520 (N_1520,In_377,In_528);
nand U1521 (N_1521,In_252,In_152);
nor U1522 (N_1522,In_59,In_473);
nor U1523 (N_1523,In_204,In_225);
or U1524 (N_1524,In_214,In_380);
nand U1525 (N_1525,In_365,In_323);
nand U1526 (N_1526,In_698,In_192);
nor U1527 (N_1527,In_593,In_637);
or U1528 (N_1528,In_645,In_538);
nor U1529 (N_1529,In_333,In_133);
or U1530 (N_1530,In_183,In_167);
nand U1531 (N_1531,In_687,In_53);
or U1532 (N_1532,In_436,In_165);
and U1533 (N_1533,In_476,In_646);
or U1534 (N_1534,In_161,In_617);
nand U1535 (N_1535,In_311,In_691);
or U1536 (N_1536,In_556,In_376);
nor U1537 (N_1537,In_350,In_381);
nor U1538 (N_1538,In_294,In_516);
and U1539 (N_1539,In_76,In_341);
or U1540 (N_1540,In_227,In_607);
nor U1541 (N_1541,In_427,In_361);
and U1542 (N_1542,In_186,In_275);
or U1543 (N_1543,In_99,In_22);
nand U1544 (N_1544,In_338,In_58);
and U1545 (N_1545,In_634,In_166);
nand U1546 (N_1546,In_383,In_659);
and U1547 (N_1547,In_189,In_297);
and U1548 (N_1548,In_10,In_283);
xor U1549 (N_1549,In_48,In_560);
or U1550 (N_1550,In_142,In_6);
nand U1551 (N_1551,In_362,In_343);
or U1552 (N_1552,In_640,In_471);
nand U1553 (N_1553,In_455,In_17);
and U1554 (N_1554,In_301,In_148);
nor U1555 (N_1555,In_237,In_258);
and U1556 (N_1556,In_180,In_537);
nand U1557 (N_1557,In_339,In_678);
and U1558 (N_1558,In_469,In_434);
nand U1559 (N_1559,In_240,In_548);
nor U1560 (N_1560,In_506,In_305);
and U1561 (N_1561,In_565,In_744);
nand U1562 (N_1562,In_379,In_339);
nor U1563 (N_1563,In_230,In_437);
nand U1564 (N_1564,In_58,In_696);
nor U1565 (N_1565,In_101,In_662);
or U1566 (N_1566,In_198,In_300);
or U1567 (N_1567,In_42,In_185);
and U1568 (N_1568,In_360,In_43);
nor U1569 (N_1569,In_541,In_104);
and U1570 (N_1570,In_220,In_12);
nand U1571 (N_1571,In_471,In_716);
and U1572 (N_1572,In_252,In_312);
nor U1573 (N_1573,In_257,In_374);
nor U1574 (N_1574,In_544,In_674);
and U1575 (N_1575,In_642,In_507);
or U1576 (N_1576,In_118,In_600);
nor U1577 (N_1577,In_722,In_12);
and U1578 (N_1578,In_660,In_457);
xor U1579 (N_1579,In_675,In_497);
nor U1580 (N_1580,In_518,In_505);
nor U1581 (N_1581,In_86,In_213);
or U1582 (N_1582,In_747,In_686);
nor U1583 (N_1583,In_742,In_39);
or U1584 (N_1584,In_267,In_742);
and U1585 (N_1585,In_417,In_434);
and U1586 (N_1586,In_145,In_136);
or U1587 (N_1587,In_110,In_435);
nand U1588 (N_1588,In_167,In_364);
nand U1589 (N_1589,In_117,In_554);
or U1590 (N_1590,In_574,In_462);
and U1591 (N_1591,In_270,In_653);
or U1592 (N_1592,In_263,In_667);
nand U1593 (N_1593,In_439,In_729);
nand U1594 (N_1594,In_134,In_684);
nor U1595 (N_1595,In_670,In_150);
or U1596 (N_1596,In_118,In_407);
and U1597 (N_1597,In_132,In_265);
and U1598 (N_1598,In_333,In_631);
or U1599 (N_1599,In_545,In_495);
nand U1600 (N_1600,In_449,In_354);
xnor U1601 (N_1601,In_555,In_634);
nand U1602 (N_1602,In_517,In_554);
nand U1603 (N_1603,In_445,In_671);
and U1604 (N_1604,In_731,In_380);
nor U1605 (N_1605,In_349,In_169);
nand U1606 (N_1606,In_381,In_351);
nand U1607 (N_1607,In_119,In_366);
nand U1608 (N_1608,In_553,In_721);
nand U1609 (N_1609,In_355,In_686);
nor U1610 (N_1610,In_744,In_688);
nand U1611 (N_1611,In_680,In_358);
nor U1612 (N_1612,In_255,In_651);
and U1613 (N_1613,In_167,In_501);
and U1614 (N_1614,In_533,In_297);
and U1615 (N_1615,In_132,In_565);
or U1616 (N_1616,In_202,In_271);
nor U1617 (N_1617,In_221,In_311);
and U1618 (N_1618,In_373,In_344);
nand U1619 (N_1619,In_123,In_486);
nand U1620 (N_1620,In_29,In_710);
and U1621 (N_1621,In_168,In_611);
or U1622 (N_1622,In_270,In_610);
nand U1623 (N_1623,In_290,In_729);
or U1624 (N_1624,In_539,In_747);
nand U1625 (N_1625,In_488,In_267);
nand U1626 (N_1626,In_491,In_470);
or U1627 (N_1627,In_18,In_688);
nand U1628 (N_1628,In_543,In_353);
nor U1629 (N_1629,In_561,In_711);
xnor U1630 (N_1630,In_100,In_388);
nand U1631 (N_1631,In_477,In_465);
nand U1632 (N_1632,In_563,In_304);
nand U1633 (N_1633,In_721,In_78);
and U1634 (N_1634,In_613,In_4);
and U1635 (N_1635,In_156,In_433);
nor U1636 (N_1636,In_185,In_293);
nor U1637 (N_1637,In_621,In_402);
nor U1638 (N_1638,In_215,In_168);
nor U1639 (N_1639,In_749,In_91);
and U1640 (N_1640,In_481,In_41);
or U1641 (N_1641,In_261,In_120);
nor U1642 (N_1642,In_687,In_415);
and U1643 (N_1643,In_11,In_55);
nand U1644 (N_1644,In_520,In_468);
or U1645 (N_1645,In_607,In_197);
nor U1646 (N_1646,In_286,In_533);
or U1647 (N_1647,In_151,In_614);
and U1648 (N_1648,In_78,In_456);
nor U1649 (N_1649,In_686,In_135);
or U1650 (N_1650,In_238,In_159);
and U1651 (N_1651,In_379,In_78);
nor U1652 (N_1652,In_718,In_32);
and U1653 (N_1653,In_666,In_466);
and U1654 (N_1654,In_703,In_378);
nor U1655 (N_1655,In_35,In_693);
or U1656 (N_1656,In_742,In_141);
nand U1657 (N_1657,In_711,In_333);
nor U1658 (N_1658,In_352,In_521);
nand U1659 (N_1659,In_607,In_699);
and U1660 (N_1660,In_112,In_481);
nor U1661 (N_1661,In_192,In_720);
and U1662 (N_1662,In_378,In_581);
nand U1663 (N_1663,In_511,In_198);
or U1664 (N_1664,In_274,In_237);
nor U1665 (N_1665,In_365,In_216);
or U1666 (N_1666,In_355,In_538);
nor U1667 (N_1667,In_121,In_242);
and U1668 (N_1668,In_66,In_688);
nor U1669 (N_1669,In_174,In_445);
and U1670 (N_1670,In_492,In_4);
xnor U1671 (N_1671,In_477,In_7);
nand U1672 (N_1672,In_464,In_361);
nor U1673 (N_1673,In_707,In_694);
or U1674 (N_1674,In_338,In_102);
nand U1675 (N_1675,In_21,In_583);
or U1676 (N_1676,In_650,In_533);
or U1677 (N_1677,In_703,In_400);
or U1678 (N_1678,In_722,In_294);
and U1679 (N_1679,In_106,In_195);
and U1680 (N_1680,In_22,In_338);
nor U1681 (N_1681,In_623,In_297);
nor U1682 (N_1682,In_308,In_78);
nand U1683 (N_1683,In_556,In_627);
nor U1684 (N_1684,In_310,In_274);
nand U1685 (N_1685,In_301,In_86);
or U1686 (N_1686,In_60,In_86);
nor U1687 (N_1687,In_118,In_235);
and U1688 (N_1688,In_196,In_641);
nand U1689 (N_1689,In_69,In_87);
and U1690 (N_1690,In_279,In_712);
nor U1691 (N_1691,In_45,In_465);
or U1692 (N_1692,In_358,In_273);
and U1693 (N_1693,In_664,In_433);
nor U1694 (N_1694,In_668,In_412);
or U1695 (N_1695,In_328,In_554);
xnor U1696 (N_1696,In_424,In_113);
and U1697 (N_1697,In_310,In_150);
nor U1698 (N_1698,In_600,In_660);
nor U1699 (N_1699,In_505,In_299);
nand U1700 (N_1700,In_59,In_157);
and U1701 (N_1701,In_86,In_345);
nand U1702 (N_1702,In_274,In_179);
nand U1703 (N_1703,In_685,In_628);
nand U1704 (N_1704,In_68,In_171);
nand U1705 (N_1705,In_255,In_301);
or U1706 (N_1706,In_377,In_204);
nand U1707 (N_1707,In_81,In_631);
xor U1708 (N_1708,In_174,In_191);
or U1709 (N_1709,In_387,In_528);
and U1710 (N_1710,In_295,In_408);
xor U1711 (N_1711,In_18,In_55);
and U1712 (N_1712,In_672,In_272);
nand U1713 (N_1713,In_208,In_54);
nor U1714 (N_1714,In_700,In_584);
or U1715 (N_1715,In_419,In_412);
or U1716 (N_1716,In_242,In_518);
nor U1717 (N_1717,In_306,In_18);
and U1718 (N_1718,In_669,In_106);
xor U1719 (N_1719,In_27,In_184);
or U1720 (N_1720,In_10,In_365);
or U1721 (N_1721,In_412,In_36);
or U1722 (N_1722,In_425,In_721);
nand U1723 (N_1723,In_84,In_728);
nor U1724 (N_1724,In_543,In_416);
and U1725 (N_1725,In_225,In_131);
nor U1726 (N_1726,In_657,In_515);
or U1727 (N_1727,In_94,In_190);
or U1728 (N_1728,In_463,In_62);
nor U1729 (N_1729,In_117,In_539);
nand U1730 (N_1730,In_341,In_202);
nor U1731 (N_1731,In_57,In_114);
nand U1732 (N_1732,In_405,In_391);
nand U1733 (N_1733,In_649,In_232);
nor U1734 (N_1734,In_715,In_432);
or U1735 (N_1735,In_230,In_237);
nand U1736 (N_1736,In_106,In_518);
nand U1737 (N_1737,In_217,In_111);
nand U1738 (N_1738,In_62,In_536);
nor U1739 (N_1739,In_664,In_191);
nor U1740 (N_1740,In_3,In_153);
or U1741 (N_1741,In_465,In_307);
nor U1742 (N_1742,In_620,In_223);
or U1743 (N_1743,In_561,In_105);
nand U1744 (N_1744,In_212,In_686);
and U1745 (N_1745,In_249,In_118);
and U1746 (N_1746,In_57,In_447);
and U1747 (N_1747,In_610,In_721);
and U1748 (N_1748,In_478,In_512);
and U1749 (N_1749,In_457,In_10);
and U1750 (N_1750,In_641,In_347);
nand U1751 (N_1751,In_420,In_576);
nor U1752 (N_1752,In_595,In_379);
and U1753 (N_1753,In_257,In_462);
and U1754 (N_1754,In_121,In_214);
or U1755 (N_1755,In_491,In_270);
and U1756 (N_1756,In_555,In_308);
and U1757 (N_1757,In_715,In_144);
and U1758 (N_1758,In_113,In_659);
and U1759 (N_1759,In_63,In_119);
and U1760 (N_1760,In_302,In_168);
or U1761 (N_1761,In_438,In_523);
nor U1762 (N_1762,In_195,In_601);
and U1763 (N_1763,In_488,In_367);
nor U1764 (N_1764,In_229,In_669);
nor U1765 (N_1765,In_503,In_558);
and U1766 (N_1766,In_268,In_383);
and U1767 (N_1767,In_25,In_513);
nand U1768 (N_1768,In_626,In_173);
or U1769 (N_1769,In_23,In_446);
and U1770 (N_1770,In_650,In_731);
xor U1771 (N_1771,In_521,In_68);
nor U1772 (N_1772,In_156,In_364);
or U1773 (N_1773,In_586,In_408);
or U1774 (N_1774,In_507,In_42);
or U1775 (N_1775,In_537,In_197);
and U1776 (N_1776,In_344,In_671);
nor U1777 (N_1777,In_395,In_479);
or U1778 (N_1778,In_730,In_55);
nand U1779 (N_1779,In_454,In_242);
or U1780 (N_1780,In_347,In_656);
and U1781 (N_1781,In_693,In_492);
or U1782 (N_1782,In_742,In_309);
nand U1783 (N_1783,In_384,In_66);
or U1784 (N_1784,In_30,In_660);
and U1785 (N_1785,In_251,In_95);
nor U1786 (N_1786,In_316,In_495);
xor U1787 (N_1787,In_683,In_172);
and U1788 (N_1788,In_533,In_291);
or U1789 (N_1789,In_588,In_670);
nor U1790 (N_1790,In_9,In_641);
or U1791 (N_1791,In_79,In_487);
nand U1792 (N_1792,In_41,In_379);
and U1793 (N_1793,In_507,In_704);
and U1794 (N_1794,In_638,In_134);
or U1795 (N_1795,In_66,In_372);
nor U1796 (N_1796,In_631,In_671);
or U1797 (N_1797,In_220,In_84);
nor U1798 (N_1798,In_173,In_472);
and U1799 (N_1799,In_162,In_600);
nand U1800 (N_1800,In_188,In_732);
and U1801 (N_1801,In_101,In_403);
nor U1802 (N_1802,In_385,In_105);
nand U1803 (N_1803,In_43,In_498);
or U1804 (N_1804,In_93,In_693);
nand U1805 (N_1805,In_84,In_113);
nand U1806 (N_1806,In_195,In_650);
and U1807 (N_1807,In_326,In_665);
nor U1808 (N_1808,In_386,In_701);
nand U1809 (N_1809,In_360,In_503);
nor U1810 (N_1810,In_183,In_474);
and U1811 (N_1811,In_466,In_176);
nor U1812 (N_1812,In_224,In_104);
nand U1813 (N_1813,In_359,In_127);
nand U1814 (N_1814,In_73,In_2);
and U1815 (N_1815,In_241,In_680);
nand U1816 (N_1816,In_55,In_635);
and U1817 (N_1817,In_180,In_657);
nand U1818 (N_1818,In_664,In_134);
nand U1819 (N_1819,In_362,In_12);
or U1820 (N_1820,In_574,In_382);
nand U1821 (N_1821,In_37,In_449);
xnor U1822 (N_1822,In_608,In_333);
or U1823 (N_1823,In_237,In_110);
nand U1824 (N_1824,In_174,In_524);
nand U1825 (N_1825,In_20,In_727);
nor U1826 (N_1826,In_508,In_179);
nand U1827 (N_1827,In_593,In_552);
or U1828 (N_1828,In_294,In_132);
nor U1829 (N_1829,In_233,In_373);
nor U1830 (N_1830,In_158,In_619);
xnor U1831 (N_1831,In_575,In_388);
or U1832 (N_1832,In_180,In_618);
nand U1833 (N_1833,In_402,In_27);
or U1834 (N_1834,In_198,In_25);
and U1835 (N_1835,In_516,In_531);
and U1836 (N_1836,In_288,In_32);
nor U1837 (N_1837,In_310,In_23);
nand U1838 (N_1838,In_62,In_246);
or U1839 (N_1839,In_521,In_711);
nand U1840 (N_1840,In_121,In_297);
nor U1841 (N_1841,In_619,In_149);
nand U1842 (N_1842,In_217,In_114);
or U1843 (N_1843,In_666,In_423);
or U1844 (N_1844,In_444,In_714);
nand U1845 (N_1845,In_368,In_526);
nor U1846 (N_1846,In_182,In_645);
or U1847 (N_1847,In_566,In_703);
or U1848 (N_1848,In_186,In_530);
nand U1849 (N_1849,In_268,In_184);
nand U1850 (N_1850,In_334,In_724);
nand U1851 (N_1851,In_340,In_294);
nor U1852 (N_1852,In_555,In_627);
or U1853 (N_1853,In_262,In_179);
and U1854 (N_1854,In_555,In_482);
nand U1855 (N_1855,In_717,In_379);
nor U1856 (N_1856,In_740,In_357);
or U1857 (N_1857,In_364,In_266);
and U1858 (N_1858,In_719,In_534);
nor U1859 (N_1859,In_608,In_580);
and U1860 (N_1860,In_133,In_608);
or U1861 (N_1861,In_110,In_596);
nand U1862 (N_1862,In_607,In_589);
nor U1863 (N_1863,In_41,In_415);
or U1864 (N_1864,In_82,In_13);
and U1865 (N_1865,In_686,In_0);
and U1866 (N_1866,In_290,In_389);
or U1867 (N_1867,In_105,In_80);
or U1868 (N_1868,In_607,In_471);
and U1869 (N_1869,In_295,In_445);
and U1870 (N_1870,In_734,In_455);
and U1871 (N_1871,In_547,In_630);
nand U1872 (N_1872,In_113,In_401);
or U1873 (N_1873,In_227,In_249);
nor U1874 (N_1874,In_135,In_575);
nor U1875 (N_1875,In_197,In_659);
or U1876 (N_1876,In_728,In_177);
nor U1877 (N_1877,In_207,In_360);
or U1878 (N_1878,In_314,In_184);
nand U1879 (N_1879,In_318,In_79);
nor U1880 (N_1880,In_361,In_11);
or U1881 (N_1881,In_489,In_389);
and U1882 (N_1882,In_632,In_593);
or U1883 (N_1883,In_688,In_617);
xor U1884 (N_1884,In_532,In_568);
nand U1885 (N_1885,In_147,In_526);
nor U1886 (N_1886,In_202,In_452);
and U1887 (N_1887,In_722,In_44);
and U1888 (N_1888,In_583,In_111);
or U1889 (N_1889,In_624,In_479);
xor U1890 (N_1890,In_567,In_271);
nor U1891 (N_1891,In_470,In_108);
and U1892 (N_1892,In_19,In_252);
nor U1893 (N_1893,In_309,In_598);
or U1894 (N_1894,In_730,In_584);
and U1895 (N_1895,In_321,In_627);
nor U1896 (N_1896,In_733,In_621);
or U1897 (N_1897,In_489,In_275);
and U1898 (N_1898,In_206,In_441);
and U1899 (N_1899,In_232,In_22);
nor U1900 (N_1900,In_118,In_630);
nand U1901 (N_1901,In_592,In_353);
and U1902 (N_1902,In_200,In_322);
nor U1903 (N_1903,In_98,In_695);
nor U1904 (N_1904,In_641,In_509);
nand U1905 (N_1905,In_702,In_37);
and U1906 (N_1906,In_284,In_719);
and U1907 (N_1907,In_462,In_209);
nand U1908 (N_1908,In_344,In_183);
or U1909 (N_1909,In_655,In_295);
nor U1910 (N_1910,In_268,In_466);
or U1911 (N_1911,In_288,In_310);
nand U1912 (N_1912,In_181,In_538);
and U1913 (N_1913,In_585,In_505);
or U1914 (N_1914,In_294,In_406);
and U1915 (N_1915,In_14,In_407);
nor U1916 (N_1916,In_193,In_478);
nor U1917 (N_1917,In_323,In_25);
nor U1918 (N_1918,In_103,In_257);
and U1919 (N_1919,In_483,In_505);
or U1920 (N_1920,In_471,In_455);
and U1921 (N_1921,In_703,In_479);
nand U1922 (N_1922,In_621,In_716);
nor U1923 (N_1923,In_600,In_58);
and U1924 (N_1924,In_271,In_469);
nor U1925 (N_1925,In_66,In_442);
and U1926 (N_1926,In_234,In_367);
and U1927 (N_1927,In_312,In_387);
and U1928 (N_1928,In_448,In_748);
and U1929 (N_1929,In_370,In_386);
and U1930 (N_1930,In_464,In_317);
nor U1931 (N_1931,In_463,In_177);
nand U1932 (N_1932,In_624,In_103);
and U1933 (N_1933,In_160,In_643);
nand U1934 (N_1934,In_228,In_453);
and U1935 (N_1935,In_79,In_653);
nand U1936 (N_1936,In_155,In_109);
and U1937 (N_1937,In_680,In_570);
or U1938 (N_1938,In_256,In_321);
nand U1939 (N_1939,In_387,In_684);
nand U1940 (N_1940,In_653,In_364);
nor U1941 (N_1941,In_525,In_169);
and U1942 (N_1942,In_334,In_232);
nand U1943 (N_1943,In_304,In_452);
and U1944 (N_1944,In_432,In_309);
or U1945 (N_1945,In_473,In_78);
nor U1946 (N_1946,In_108,In_300);
and U1947 (N_1947,In_744,In_728);
nor U1948 (N_1948,In_497,In_734);
or U1949 (N_1949,In_658,In_731);
nand U1950 (N_1950,In_429,In_399);
nor U1951 (N_1951,In_447,In_633);
nand U1952 (N_1952,In_406,In_409);
or U1953 (N_1953,In_32,In_107);
nor U1954 (N_1954,In_733,In_470);
or U1955 (N_1955,In_530,In_712);
or U1956 (N_1956,In_349,In_426);
nor U1957 (N_1957,In_295,In_357);
nand U1958 (N_1958,In_604,In_90);
nor U1959 (N_1959,In_15,In_729);
xor U1960 (N_1960,In_660,In_467);
nand U1961 (N_1961,In_736,In_310);
and U1962 (N_1962,In_320,In_283);
or U1963 (N_1963,In_13,In_97);
or U1964 (N_1964,In_613,In_736);
nor U1965 (N_1965,In_531,In_28);
nor U1966 (N_1966,In_691,In_52);
nor U1967 (N_1967,In_573,In_412);
nand U1968 (N_1968,In_302,In_252);
and U1969 (N_1969,In_394,In_53);
or U1970 (N_1970,In_453,In_443);
xor U1971 (N_1971,In_197,In_74);
and U1972 (N_1972,In_702,In_109);
and U1973 (N_1973,In_428,In_691);
and U1974 (N_1974,In_396,In_616);
nor U1975 (N_1975,In_155,In_294);
or U1976 (N_1976,In_537,In_635);
and U1977 (N_1977,In_324,In_249);
and U1978 (N_1978,In_367,In_611);
or U1979 (N_1979,In_82,In_152);
nand U1980 (N_1980,In_83,In_388);
and U1981 (N_1981,In_406,In_513);
nand U1982 (N_1982,In_703,In_417);
nand U1983 (N_1983,In_572,In_258);
and U1984 (N_1984,In_369,In_107);
nand U1985 (N_1985,In_338,In_105);
or U1986 (N_1986,In_275,In_555);
nor U1987 (N_1987,In_172,In_404);
nand U1988 (N_1988,In_304,In_25);
nor U1989 (N_1989,In_435,In_607);
or U1990 (N_1990,In_749,In_408);
nor U1991 (N_1991,In_513,In_251);
nand U1992 (N_1992,In_686,In_683);
and U1993 (N_1993,In_326,In_709);
or U1994 (N_1994,In_451,In_283);
or U1995 (N_1995,In_280,In_590);
nand U1996 (N_1996,In_56,In_641);
nand U1997 (N_1997,In_597,In_288);
and U1998 (N_1998,In_220,In_411);
nand U1999 (N_1999,In_10,In_81);
nand U2000 (N_2000,In_47,In_439);
nand U2001 (N_2001,In_5,In_293);
and U2002 (N_2002,In_288,In_411);
nor U2003 (N_2003,In_5,In_131);
and U2004 (N_2004,In_632,In_749);
and U2005 (N_2005,In_259,In_89);
nand U2006 (N_2006,In_651,In_678);
nand U2007 (N_2007,In_454,In_732);
nand U2008 (N_2008,In_232,In_299);
or U2009 (N_2009,In_255,In_149);
or U2010 (N_2010,In_226,In_353);
xnor U2011 (N_2011,In_716,In_357);
nor U2012 (N_2012,In_494,In_430);
or U2013 (N_2013,In_87,In_221);
nor U2014 (N_2014,In_159,In_21);
nor U2015 (N_2015,In_662,In_123);
nor U2016 (N_2016,In_419,In_576);
nand U2017 (N_2017,In_597,In_589);
or U2018 (N_2018,In_147,In_716);
nand U2019 (N_2019,In_264,In_588);
nor U2020 (N_2020,In_564,In_441);
and U2021 (N_2021,In_282,In_91);
or U2022 (N_2022,In_202,In_184);
nor U2023 (N_2023,In_24,In_312);
nand U2024 (N_2024,In_156,In_481);
nand U2025 (N_2025,In_702,In_129);
or U2026 (N_2026,In_608,In_229);
and U2027 (N_2027,In_396,In_227);
nor U2028 (N_2028,In_500,In_406);
or U2029 (N_2029,In_136,In_703);
nand U2030 (N_2030,In_533,In_711);
nand U2031 (N_2031,In_86,In_140);
and U2032 (N_2032,In_348,In_14);
and U2033 (N_2033,In_741,In_490);
and U2034 (N_2034,In_372,In_93);
nand U2035 (N_2035,In_174,In_483);
and U2036 (N_2036,In_88,In_176);
and U2037 (N_2037,In_315,In_151);
or U2038 (N_2038,In_182,In_557);
or U2039 (N_2039,In_146,In_103);
nand U2040 (N_2040,In_195,In_689);
or U2041 (N_2041,In_735,In_522);
or U2042 (N_2042,In_627,In_20);
or U2043 (N_2043,In_378,In_312);
and U2044 (N_2044,In_612,In_452);
or U2045 (N_2045,In_605,In_190);
or U2046 (N_2046,In_43,In_417);
and U2047 (N_2047,In_139,In_56);
nand U2048 (N_2048,In_126,In_374);
or U2049 (N_2049,In_623,In_272);
or U2050 (N_2050,In_149,In_137);
nand U2051 (N_2051,In_146,In_596);
and U2052 (N_2052,In_598,In_223);
and U2053 (N_2053,In_749,In_428);
and U2054 (N_2054,In_732,In_384);
nand U2055 (N_2055,In_568,In_655);
or U2056 (N_2056,In_379,In_705);
and U2057 (N_2057,In_477,In_669);
or U2058 (N_2058,In_493,In_193);
nand U2059 (N_2059,In_677,In_702);
and U2060 (N_2060,In_286,In_86);
and U2061 (N_2061,In_182,In_554);
and U2062 (N_2062,In_383,In_79);
or U2063 (N_2063,In_131,In_275);
nor U2064 (N_2064,In_519,In_681);
and U2065 (N_2065,In_412,In_52);
nand U2066 (N_2066,In_265,In_679);
nor U2067 (N_2067,In_310,In_726);
nor U2068 (N_2068,In_194,In_545);
and U2069 (N_2069,In_375,In_248);
nor U2070 (N_2070,In_643,In_418);
or U2071 (N_2071,In_473,In_330);
nand U2072 (N_2072,In_308,In_39);
and U2073 (N_2073,In_214,In_249);
nand U2074 (N_2074,In_722,In_9);
nor U2075 (N_2075,In_431,In_248);
and U2076 (N_2076,In_590,In_414);
nand U2077 (N_2077,In_665,In_446);
nor U2078 (N_2078,In_653,In_136);
or U2079 (N_2079,In_103,In_444);
nor U2080 (N_2080,In_119,In_543);
and U2081 (N_2081,In_577,In_415);
nand U2082 (N_2082,In_379,In_435);
or U2083 (N_2083,In_187,In_508);
or U2084 (N_2084,In_699,In_330);
nor U2085 (N_2085,In_135,In_31);
or U2086 (N_2086,In_304,In_99);
or U2087 (N_2087,In_540,In_176);
and U2088 (N_2088,In_363,In_182);
and U2089 (N_2089,In_680,In_648);
nor U2090 (N_2090,In_335,In_177);
or U2091 (N_2091,In_682,In_44);
and U2092 (N_2092,In_701,In_206);
nand U2093 (N_2093,In_438,In_242);
and U2094 (N_2094,In_390,In_159);
nor U2095 (N_2095,In_518,In_342);
xnor U2096 (N_2096,In_639,In_307);
and U2097 (N_2097,In_724,In_125);
nand U2098 (N_2098,In_120,In_236);
or U2099 (N_2099,In_548,In_483);
nor U2100 (N_2100,In_213,In_566);
and U2101 (N_2101,In_7,In_324);
nand U2102 (N_2102,In_275,In_35);
nor U2103 (N_2103,In_637,In_675);
nor U2104 (N_2104,In_201,In_319);
nand U2105 (N_2105,In_221,In_509);
and U2106 (N_2106,In_388,In_555);
xnor U2107 (N_2107,In_700,In_116);
or U2108 (N_2108,In_184,In_602);
and U2109 (N_2109,In_469,In_183);
and U2110 (N_2110,In_620,In_484);
nor U2111 (N_2111,In_329,In_343);
nor U2112 (N_2112,In_706,In_241);
or U2113 (N_2113,In_534,In_509);
xnor U2114 (N_2114,In_444,In_539);
and U2115 (N_2115,In_52,In_403);
nor U2116 (N_2116,In_535,In_269);
nor U2117 (N_2117,In_507,In_330);
nor U2118 (N_2118,In_273,In_306);
or U2119 (N_2119,In_57,In_458);
or U2120 (N_2120,In_676,In_447);
and U2121 (N_2121,In_76,In_88);
or U2122 (N_2122,In_454,In_370);
and U2123 (N_2123,In_581,In_412);
or U2124 (N_2124,In_48,In_126);
and U2125 (N_2125,In_57,In_297);
or U2126 (N_2126,In_81,In_196);
nor U2127 (N_2127,In_731,In_58);
or U2128 (N_2128,In_242,In_431);
and U2129 (N_2129,In_137,In_348);
nor U2130 (N_2130,In_465,In_490);
nor U2131 (N_2131,In_37,In_222);
nor U2132 (N_2132,In_665,In_547);
nand U2133 (N_2133,In_75,In_382);
and U2134 (N_2134,In_74,In_15);
nor U2135 (N_2135,In_699,In_627);
or U2136 (N_2136,In_45,In_141);
nand U2137 (N_2137,In_84,In_144);
and U2138 (N_2138,In_649,In_334);
nand U2139 (N_2139,In_723,In_69);
and U2140 (N_2140,In_330,In_171);
nand U2141 (N_2141,In_673,In_103);
nor U2142 (N_2142,In_575,In_693);
and U2143 (N_2143,In_135,In_199);
xor U2144 (N_2144,In_489,In_313);
or U2145 (N_2145,In_550,In_476);
or U2146 (N_2146,In_242,In_246);
nand U2147 (N_2147,In_694,In_214);
nand U2148 (N_2148,In_365,In_561);
or U2149 (N_2149,In_100,In_219);
nor U2150 (N_2150,In_429,In_610);
nor U2151 (N_2151,In_702,In_326);
or U2152 (N_2152,In_612,In_483);
nor U2153 (N_2153,In_440,In_558);
or U2154 (N_2154,In_10,In_214);
xnor U2155 (N_2155,In_238,In_310);
nor U2156 (N_2156,In_461,In_688);
nor U2157 (N_2157,In_397,In_611);
nor U2158 (N_2158,In_422,In_116);
nor U2159 (N_2159,In_701,In_387);
nor U2160 (N_2160,In_429,In_37);
nand U2161 (N_2161,In_218,In_45);
nand U2162 (N_2162,In_11,In_692);
or U2163 (N_2163,In_147,In_21);
or U2164 (N_2164,In_276,In_449);
nor U2165 (N_2165,In_103,In_287);
or U2166 (N_2166,In_321,In_29);
nor U2167 (N_2167,In_677,In_453);
nand U2168 (N_2168,In_625,In_100);
nor U2169 (N_2169,In_306,In_338);
or U2170 (N_2170,In_219,In_400);
or U2171 (N_2171,In_437,In_118);
or U2172 (N_2172,In_78,In_522);
nand U2173 (N_2173,In_144,In_490);
nand U2174 (N_2174,In_514,In_151);
or U2175 (N_2175,In_195,In_213);
and U2176 (N_2176,In_289,In_663);
nor U2177 (N_2177,In_278,In_315);
nand U2178 (N_2178,In_446,In_381);
nand U2179 (N_2179,In_180,In_32);
nand U2180 (N_2180,In_410,In_293);
nor U2181 (N_2181,In_102,In_110);
or U2182 (N_2182,In_670,In_74);
nand U2183 (N_2183,In_465,In_310);
xor U2184 (N_2184,In_613,In_634);
xnor U2185 (N_2185,In_132,In_207);
and U2186 (N_2186,In_649,In_508);
nor U2187 (N_2187,In_145,In_459);
and U2188 (N_2188,In_482,In_389);
or U2189 (N_2189,In_661,In_519);
or U2190 (N_2190,In_425,In_152);
nand U2191 (N_2191,In_549,In_486);
and U2192 (N_2192,In_75,In_335);
nand U2193 (N_2193,In_726,In_447);
nor U2194 (N_2194,In_227,In_330);
nand U2195 (N_2195,In_721,In_205);
nand U2196 (N_2196,In_299,In_95);
nor U2197 (N_2197,In_173,In_598);
and U2198 (N_2198,In_75,In_147);
nand U2199 (N_2199,In_427,In_132);
and U2200 (N_2200,In_471,In_618);
nor U2201 (N_2201,In_423,In_417);
and U2202 (N_2202,In_337,In_281);
or U2203 (N_2203,In_84,In_597);
or U2204 (N_2204,In_182,In_510);
nand U2205 (N_2205,In_428,In_659);
or U2206 (N_2206,In_529,In_97);
nor U2207 (N_2207,In_643,In_128);
or U2208 (N_2208,In_494,In_166);
nor U2209 (N_2209,In_133,In_491);
or U2210 (N_2210,In_391,In_345);
and U2211 (N_2211,In_570,In_216);
and U2212 (N_2212,In_353,In_286);
nand U2213 (N_2213,In_124,In_401);
nand U2214 (N_2214,In_128,In_479);
and U2215 (N_2215,In_283,In_392);
or U2216 (N_2216,In_575,In_10);
nor U2217 (N_2217,In_423,In_687);
nor U2218 (N_2218,In_314,In_149);
or U2219 (N_2219,In_11,In_199);
or U2220 (N_2220,In_207,In_706);
nand U2221 (N_2221,In_102,In_412);
nor U2222 (N_2222,In_719,In_75);
and U2223 (N_2223,In_421,In_59);
nand U2224 (N_2224,In_90,In_531);
or U2225 (N_2225,In_205,In_398);
xnor U2226 (N_2226,In_463,In_74);
xor U2227 (N_2227,In_345,In_157);
and U2228 (N_2228,In_12,In_118);
and U2229 (N_2229,In_646,In_390);
nor U2230 (N_2230,In_296,In_706);
nor U2231 (N_2231,In_382,In_590);
nand U2232 (N_2232,In_333,In_435);
and U2233 (N_2233,In_457,In_184);
or U2234 (N_2234,In_287,In_625);
nor U2235 (N_2235,In_708,In_565);
and U2236 (N_2236,In_600,In_127);
nor U2237 (N_2237,In_139,In_535);
nand U2238 (N_2238,In_671,In_255);
and U2239 (N_2239,In_279,In_207);
xnor U2240 (N_2240,In_714,In_690);
or U2241 (N_2241,In_472,In_373);
nor U2242 (N_2242,In_257,In_270);
or U2243 (N_2243,In_245,In_552);
xnor U2244 (N_2244,In_371,In_674);
or U2245 (N_2245,In_660,In_103);
nand U2246 (N_2246,In_384,In_33);
or U2247 (N_2247,In_228,In_648);
and U2248 (N_2248,In_5,In_671);
nor U2249 (N_2249,In_719,In_660);
or U2250 (N_2250,In_485,In_186);
nand U2251 (N_2251,In_389,In_196);
or U2252 (N_2252,In_404,In_615);
xor U2253 (N_2253,In_262,In_314);
nand U2254 (N_2254,In_676,In_564);
and U2255 (N_2255,In_472,In_486);
or U2256 (N_2256,In_57,In_485);
nand U2257 (N_2257,In_141,In_712);
or U2258 (N_2258,In_42,In_482);
nor U2259 (N_2259,In_368,In_62);
or U2260 (N_2260,In_103,In_182);
xor U2261 (N_2261,In_616,In_353);
nor U2262 (N_2262,In_367,In_533);
or U2263 (N_2263,In_34,In_521);
or U2264 (N_2264,In_376,In_160);
nor U2265 (N_2265,In_659,In_688);
or U2266 (N_2266,In_232,In_528);
nor U2267 (N_2267,In_298,In_328);
nand U2268 (N_2268,In_253,In_453);
xnor U2269 (N_2269,In_408,In_85);
and U2270 (N_2270,In_121,In_101);
and U2271 (N_2271,In_296,In_503);
nor U2272 (N_2272,In_63,In_376);
and U2273 (N_2273,In_629,In_43);
or U2274 (N_2274,In_250,In_439);
nand U2275 (N_2275,In_40,In_38);
or U2276 (N_2276,In_731,In_403);
nand U2277 (N_2277,In_637,In_620);
and U2278 (N_2278,In_49,In_727);
or U2279 (N_2279,In_556,In_666);
or U2280 (N_2280,In_103,In_677);
nand U2281 (N_2281,In_273,In_317);
and U2282 (N_2282,In_61,In_27);
nor U2283 (N_2283,In_157,In_416);
or U2284 (N_2284,In_97,In_346);
nor U2285 (N_2285,In_64,In_385);
or U2286 (N_2286,In_92,In_124);
nand U2287 (N_2287,In_28,In_207);
nor U2288 (N_2288,In_243,In_183);
and U2289 (N_2289,In_600,In_656);
or U2290 (N_2290,In_580,In_637);
or U2291 (N_2291,In_381,In_461);
or U2292 (N_2292,In_230,In_52);
or U2293 (N_2293,In_32,In_652);
and U2294 (N_2294,In_708,In_108);
nor U2295 (N_2295,In_722,In_501);
nand U2296 (N_2296,In_206,In_442);
nand U2297 (N_2297,In_492,In_571);
nand U2298 (N_2298,In_35,In_473);
nor U2299 (N_2299,In_482,In_532);
xnor U2300 (N_2300,In_662,In_613);
or U2301 (N_2301,In_332,In_85);
nor U2302 (N_2302,In_198,In_570);
nand U2303 (N_2303,In_704,In_352);
nor U2304 (N_2304,In_175,In_317);
nor U2305 (N_2305,In_127,In_227);
and U2306 (N_2306,In_49,In_565);
nor U2307 (N_2307,In_457,In_441);
or U2308 (N_2308,In_382,In_160);
and U2309 (N_2309,In_421,In_427);
and U2310 (N_2310,In_144,In_115);
or U2311 (N_2311,In_626,In_302);
and U2312 (N_2312,In_551,In_518);
nand U2313 (N_2313,In_281,In_345);
and U2314 (N_2314,In_331,In_310);
and U2315 (N_2315,In_254,In_680);
or U2316 (N_2316,In_680,In_123);
or U2317 (N_2317,In_75,In_205);
nor U2318 (N_2318,In_631,In_93);
or U2319 (N_2319,In_682,In_626);
and U2320 (N_2320,In_629,In_405);
nand U2321 (N_2321,In_222,In_474);
or U2322 (N_2322,In_673,In_6);
or U2323 (N_2323,In_168,In_304);
nand U2324 (N_2324,In_616,In_411);
or U2325 (N_2325,In_584,In_373);
nand U2326 (N_2326,In_235,In_43);
nand U2327 (N_2327,In_578,In_457);
or U2328 (N_2328,In_740,In_712);
nand U2329 (N_2329,In_519,In_273);
nor U2330 (N_2330,In_118,In_465);
or U2331 (N_2331,In_613,In_463);
nor U2332 (N_2332,In_65,In_461);
nand U2333 (N_2333,In_393,In_553);
nand U2334 (N_2334,In_551,In_297);
nand U2335 (N_2335,In_443,In_591);
nand U2336 (N_2336,In_519,In_43);
or U2337 (N_2337,In_237,In_3);
nand U2338 (N_2338,In_434,In_367);
nand U2339 (N_2339,In_697,In_682);
nand U2340 (N_2340,In_559,In_735);
and U2341 (N_2341,In_113,In_732);
or U2342 (N_2342,In_651,In_694);
and U2343 (N_2343,In_521,In_386);
nand U2344 (N_2344,In_406,In_374);
or U2345 (N_2345,In_242,In_311);
and U2346 (N_2346,In_97,In_707);
nor U2347 (N_2347,In_325,In_589);
nor U2348 (N_2348,In_407,In_349);
and U2349 (N_2349,In_421,In_170);
or U2350 (N_2350,In_687,In_302);
nor U2351 (N_2351,In_574,In_104);
and U2352 (N_2352,In_73,In_669);
and U2353 (N_2353,In_523,In_493);
or U2354 (N_2354,In_94,In_737);
nor U2355 (N_2355,In_175,In_465);
nand U2356 (N_2356,In_693,In_371);
or U2357 (N_2357,In_26,In_480);
nor U2358 (N_2358,In_591,In_179);
nand U2359 (N_2359,In_41,In_459);
nor U2360 (N_2360,In_677,In_21);
or U2361 (N_2361,In_682,In_182);
and U2362 (N_2362,In_313,In_720);
nor U2363 (N_2363,In_651,In_22);
nand U2364 (N_2364,In_454,In_12);
or U2365 (N_2365,In_98,In_590);
and U2366 (N_2366,In_532,In_604);
and U2367 (N_2367,In_500,In_198);
nor U2368 (N_2368,In_66,In_292);
xor U2369 (N_2369,In_650,In_144);
and U2370 (N_2370,In_614,In_461);
nor U2371 (N_2371,In_502,In_714);
nand U2372 (N_2372,In_436,In_89);
nor U2373 (N_2373,In_389,In_438);
nand U2374 (N_2374,In_34,In_5);
and U2375 (N_2375,In_662,In_308);
nor U2376 (N_2376,In_456,In_583);
nor U2377 (N_2377,In_56,In_550);
or U2378 (N_2378,In_49,In_13);
or U2379 (N_2379,In_235,In_145);
or U2380 (N_2380,In_351,In_141);
nand U2381 (N_2381,In_72,In_616);
nor U2382 (N_2382,In_648,In_135);
and U2383 (N_2383,In_82,In_570);
nand U2384 (N_2384,In_124,In_89);
or U2385 (N_2385,In_468,In_107);
nor U2386 (N_2386,In_739,In_735);
and U2387 (N_2387,In_95,In_612);
and U2388 (N_2388,In_303,In_202);
nand U2389 (N_2389,In_270,In_322);
nand U2390 (N_2390,In_612,In_65);
and U2391 (N_2391,In_0,In_747);
nor U2392 (N_2392,In_352,In_178);
and U2393 (N_2393,In_531,In_571);
or U2394 (N_2394,In_605,In_7);
or U2395 (N_2395,In_132,In_639);
nor U2396 (N_2396,In_437,In_695);
and U2397 (N_2397,In_640,In_578);
nor U2398 (N_2398,In_125,In_602);
nand U2399 (N_2399,In_554,In_294);
and U2400 (N_2400,In_189,In_281);
or U2401 (N_2401,In_700,In_554);
nor U2402 (N_2402,In_560,In_661);
xor U2403 (N_2403,In_621,In_730);
nor U2404 (N_2404,In_682,In_643);
or U2405 (N_2405,In_660,In_64);
or U2406 (N_2406,In_386,In_451);
nor U2407 (N_2407,In_451,In_24);
or U2408 (N_2408,In_645,In_451);
xor U2409 (N_2409,In_613,In_593);
nand U2410 (N_2410,In_697,In_742);
and U2411 (N_2411,In_683,In_50);
xor U2412 (N_2412,In_590,In_512);
nand U2413 (N_2413,In_560,In_712);
nor U2414 (N_2414,In_258,In_139);
nand U2415 (N_2415,In_39,In_74);
and U2416 (N_2416,In_195,In_246);
nor U2417 (N_2417,In_215,In_532);
nand U2418 (N_2418,In_509,In_348);
nor U2419 (N_2419,In_462,In_715);
and U2420 (N_2420,In_71,In_532);
or U2421 (N_2421,In_571,In_679);
and U2422 (N_2422,In_283,In_476);
nand U2423 (N_2423,In_318,In_32);
or U2424 (N_2424,In_393,In_258);
nand U2425 (N_2425,In_153,In_435);
nand U2426 (N_2426,In_454,In_346);
nand U2427 (N_2427,In_362,In_408);
or U2428 (N_2428,In_250,In_517);
nand U2429 (N_2429,In_374,In_329);
nand U2430 (N_2430,In_52,In_440);
or U2431 (N_2431,In_435,In_722);
or U2432 (N_2432,In_122,In_102);
nor U2433 (N_2433,In_342,In_411);
nand U2434 (N_2434,In_117,In_698);
nor U2435 (N_2435,In_144,In_704);
or U2436 (N_2436,In_216,In_151);
nand U2437 (N_2437,In_557,In_154);
or U2438 (N_2438,In_258,In_326);
nor U2439 (N_2439,In_201,In_646);
and U2440 (N_2440,In_653,In_10);
nor U2441 (N_2441,In_112,In_534);
or U2442 (N_2442,In_556,In_611);
nor U2443 (N_2443,In_611,In_449);
or U2444 (N_2444,In_167,In_296);
and U2445 (N_2445,In_620,In_677);
nor U2446 (N_2446,In_622,In_264);
nand U2447 (N_2447,In_349,In_61);
nor U2448 (N_2448,In_329,In_139);
nor U2449 (N_2449,In_328,In_326);
and U2450 (N_2450,In_450,In_267);
and U2451 (N_2451,In_91,In_318);
or U2452 (N_2452,In_657,In_349);
nor U2453 (N_2453,In_515,In_514);
nand U2454 (N_2454,In_262,In_228);
or U2455 (N_2455,In_693,In_64);
nor U2456 (N_2456,In_212,In_346);
or U2457 (N_2457,In_308,In_403);
or U2458 (N_2458,In_41,In_565);
nand U2459 (N_2459,In_180,In_182);
and U2460 (N_2460,In_283,In_524);
or U2461 (N_2461,In_196,In_222);
nand U2462 (N_2462,In_101,In_180);
or U2463 (N_2463,In_570,In_134);
nand U2464 (N_2464,In_119,In_97);
and U2465 (N_2465,In_506,In_358);
nor U2466 (N_2466,In_541,In_632);
nand U2467 (N_2467,In_1,In_241);
nor U2468 (N_2468,In_531,In_520);
and U2469 (N_2469,In_404,In_143);
nor U2470 (N_2470,In_578,In_486);
or U2471 (N_2471,In_317,In_468);
and U2472 (N_2472,In_147,In_184);
nor U2473 (N_2473,In_450,In_279);
nand U2474 (N_2474,In_600,In_379);
or U2475 (N_2475,In_185,In_80);
nand U2476 (N_2476,In_309,In_644);
and U2477 (N_2477,In_36,In_274);
or U2478 (N_2478,In_327,In_116);
or U2479 (N_2479,In_141,In_507);
nor U2480 (N_2480,In_306,In_672);
and U2481 (N_2481,In_604,In_219);
or U2482 (N_2482,In_504,In_574);
or U2483 (N_2483,In_49,In_108);
and U2484 (N_2484,In_289,In_712);
and U2485 (N_2485,In_203,In_432);
and U2486 (N_2486,In_171,In_593);
nand U2487 (N_2487,In_495,In_626);
xor U2488 (N_2488,In_413,In_511);
nor U2489 (N_2489,In_467,In_645);
nand U2490 (N_2490,In_65,In_683);
and U2491 (N_2491,In_190,In_299);
nand U2492 (N_2492,In_621,In_690);
nor U2493 (N_2493,In_607,In_293);
and U2494 (N_2494,In_394,In_367);
nor U2495 (N_2495,In_204,In_90);
nor U2496 (N_2496,In_56,In_273);
or U2497 (N_2497,In_211,In_407);
nor U2498 (N_2498,In_186,In_83);
nor U2499 (N_2499,In_26,In_659);
or U2500 (N_2500,N_1331,N_1444);
and U2501 (N_2501,N_30,N_2165);
nor U2502 (N_2502,N_1280,N_1653);
nor U2503 (N_2503,N_1177,N_37);
nor U2504 (N_2504,N_2163,N_2051);
nand U2505 (N_2505,N_2082,N_1725);
nand U2506 (N_2506,N_1135,N_1461);
nor U2507 (N_2507,N_1965,N_2212);
and U2508 (N_2508,N_236,N_1946);
and U2509 (N_2509,N_632,N_1832);
nor U2510 (N_2510,N_2264,N_2132);
nand U2511 (N_2511,N_1109,N_1776);
nor U2512 (N_2512,N_2145,N_344);
nand U2513 (N_2513,N_1187,N_1614);
and U2514 (N_2514,N_2384,N_1622);
and U2515 (N_2515,N_2293,N_42);
and U2516 (N_2516,N_1524,N_1637);
or U2517 (N_2517,N_1968,N_1894);
nor U2518 (N_2518,N_1247,N_1134);
nor U2519 (N_2519,N_868,N_681);
and U2520 (N_2520,N_63,N_2441);
nand U2521 (N_2521,N_1991,N_2406);
nor U2522 (N_2522,N_2007,N_583);
nand U2523 (N_2523,N_1083,N_2477);
nand U2524 (N_2524,N_43,N_2416);
nor U2525 (N_2525,N_1272,N_1287);
and U2526 (N_2526,N_1679,N_1162);
nor U2527 (N_2527,N_93,N_1147);
nand U2528 (N_2528,N_882,N_2197);
nor U2529 (N_2529,N_836,N_644);
nand U2530 (N_2530,N_452,N_606);
and U2531 (N_2531,N_809,N_148);
and U2532 (N_2532,N_1230,N_1962);
nor U2533 (N_2533,N_4,N_352);
or U2534 (N_2534,N_2249,N_1730);
or U2535 (N_2535,N_394,N_2292);
nand U2536 (N_2536,N_1315,N_2469);
nand U2537 (N_2537,N_663,N_1263);
nor U2538 (N_2538,N_2036,N_370);
or U2539 (N_2539,N_947,N_2490);
or U2540 (N_2540,N_1802,N_1577);
and U2541 (N_2541,N_793,N_1032);
nor U2542 (N_2542,N_1555,N_1954);
and U2543 (N_2543,N_1449,N_2077);
nand U2544 (N_2544,N_319,N_243);
or U2545 (N_2545,N_197,N_639);
or U2546 (N_2546,N_2083,N_1626);
nand U2547 (N_2547,N_780,N_802);
or U2548 (N_2548,N_1342,N_1689);
nor U2549 (N_2549,N_589,N_1706);
nand U2550 (N_2550,N_118,N_465);
and U2551 (N_2551,N_1124,N_1768);
or U2552 (N_2552,N_17,N_1545);
and U2553 (N_2553,N_1349,N_204);
or U2554 (N_2554,N_396,N_1045);
nand U2555 (N_2555,N_1676,N_1085);
nor U2556 (N_2556,N_737,N_634);
and U2557 (N_2557,N_2414,N_2284);
nor U2558 (N_2558,N_1217,N_374);
nand U2559 (N_2559,N_254,N_1463);
nand U2560 (N_2560,N_469,N_2348);
nor U2561 (N_2561,N_1101,N_2426);
and U2562 (N_2562,N_1019,N_419);
nand U2563 (N_2563,N_1932,N_1501);
or U2564 (N_2564,N_298,N_1148);
nand U2565 (N_2565,N_779,N_619);
nor U2566 (N_2566,N_1511,N_1834);
nand U2567 (N_2567,N_772,N_796);
nor U2568 (N_2568,N_1967,N_1738);
nand U2569 (N_2569,N_862,N_1274);
or U2570 (N_2570,N_574,N_1371);
or U2571 (N_2571,N_1901,N_482);
nand U2572 (N_2572,N_925,N_1432);
or U2573 (N_2573,N_937,N_2311);
and U2574 (N_2574,N_2114,N_797);
nor U2575 (N_2575,N_2043,N_1029);
or U2576 (N_2576,N_1119,N_2067);
nand U2577 (N_2577,N_305,N_2494);
nor U2578 (N_2578,N_34,N_2009);
or U2579 (N_2579,N_1726,N_211);
nor U2580 (N_2580,N_1356,N_2300);
and U2581 (N_2581,N_1269,N_2245);
nor U2582 (N_2582,N_1251,N_2241);
nor U2583 (N_2583,N_1510,N_861);
nor U2584 (N_2584,N_1339,N_2252);
and U2585 (N_2585,N_304,N_1030);
xor U2586 (N_2586,N_1757,N_1990);
nand U2587 (N_2587,N_0,N_833);
or U2588 (N_2588,N_1774,N_624);
nand U2589 (N_2589,N_974,N_2331);
and U2590 (N_2590,N_1044,N_637);
or U2591 (N_2591,N_27,N_52);
or U2592 (N_2592,N_1546,N_1733);
or U2593 (N_2593,N_2035,N_1308);
nand U2594 (N_2594,N_1769,N_2094);
nor U2595 (N_2595,N_969,N_2373);
or U2596 (N_2596,N_1721,N_934);
nand U2597 (N_2597,N_1457,N_1139);
or U2598 (N_2598,N_1469,N_1857);
or U2599 (N_2599,N_19,N_159);
or U2600 (N_2600,N_1022,N_1271);
nand U2601 (N_2601,N_1224,N_1068);
xor U2602 (N_2602,N_1131,N_1710);
nor U2603 (N_2603,N_2461,N_203);
and U2604 (N_2604,N_573,N_1541);
nor U2605 (N_2605,N_545,N_2111);
nor U2606 (N_2606,N_2462,N_2156);
or U2607 (N_2607,N_2370,N_1788);
nand U2608 (N_2608,N_2480,N_1050);
and U2609 (N_2609,N_983,N_738);
and U2610 (N_2610,N_1113,N_257);
nor U2611 (N_2611,N_1021,N_1599);
or U2612 (N_2612,N_647,N_744);
nand U2613 (N_2613,N_2183,N_1665);
and U2614 (N_2614,N_15,N_373);
nor U2615 (N_2615,N_1695,N_1326);
or U2616 (N_2616,N_853,N_2261);
nor U2617 (N_2617,N_963,N_669);
nor U2618 (N_2618,N_47,N_985);
or U2619 (N_2619,N_1057,N_2062);
nand U2620 (N_2620,N_713,N_2275);
nor U2621 (N_2621,N_1236,N_390);
nand U2622 (N_2622,N_160,N_1016);
and U2623 (N_2623,N_1896,N_603);
nand U2624 (N_2624,N_912,N_801);
and U2625 (N_2625,N_2305,N_1839);
nand U2626 (N_2626,N_962,N_742);
and U2627 (N_2627,N_308,N_1242);
or U2628 (N_2628,N_363,N_1907);
or U2629 (N_2629,N_1114,N_1570);
or U2630 (N_2630,N_1681,N_847);
or U2631 (N_2631,N_725,N_2115);
nor U2632 (N_2632,N_1041,N_2027);
nand U2633 (N_2633,N_1392,N_917);
nor U2634 (N_2634,N_1741,N_2421);
nand U2635 (N_2635,N_310,N_169);
nor U2636 (N_2636,N_1970,N_894);
nand U2637 (N_2637,N_709,N_1685);
and U2638 (N_2638,N_1631,N_288);
xnor U2639 (N_2639,N_629,N_2060);
or U2640 (N_2640,N_184,N_2203);
or U2641 (N_2641,N_2453,N_2313);
or U2642 (N_2642,N_450,N_2238);
nor U2643 (N_2643,N_913,N_1241);
or U2644 (N_2644,N_2182,N_411);
nand U2645 (N_2645,N_733,N_1402);
or U2646 (N_2646,N_295,N_1426);
or U2647 (N_2647,N_2354,N_763);
nor U2648 (N_2648,N_1483,N_154);
xnor U2649 (N_2649,N_1380,N_783);
or U2650 (N_2650,N_1824,N_817);
and U2651 (N_2651,N_60,N_2129);
or U2652 (N_2652,N_2136,N_1943);
or U2653 (N_2653,N_490,N_1398);
and U2654 (N_2654,N_475,N_1795);
or U2655 (N_2655,N_2096,N_1306);
nor U2656 (N_2656,N_410,N_578);
and U2657 (N_2657,N_1589,N_1488);
nand U2658 (N_2658,N_426,N_514);
nor U2659 (N_2659,N_1898,N_2176);
and U2660 (N_2660,N_189,N_1408);
nor U2661 (N_2661,N_2170,N_198);
nand U2662 (N_2662,N_795,N_501);
nand U2663 (N_2663,N_671,N_989);
or U2664 (N_2664,N_527,N_977);
or U2665 (N_2665,N_628,N_2201);
nand U2666 (N_2666,N_1838,N_479);
or U2667 (N_2667,N_186,N_1663);
or U2668 (N_2668,N_1644,N_289);
and U2669 (N_2669,N_1835,N_904);
nor U2670 (N_2670,N_1034,N_2104);
nor U2671 (N_2671,N_339,N_78);
nor U2672 (N_2672,N_35,N_1979);
nand U2673 (N_2673,N_326,N_851);
nand U2674 (N_2674,N_1982,N_519);
or U2675 (N_2675,N_1530,N_79);
nand U2676 (N_2676,N_1081,N_1645);
or U2677 (N_2677,N_264,N_515);
or U2678 (N_2678,N_1715,N_290);
and U2679 (N_2679,N_2380,N_1110);
and U2680 (N_2680,N_45,N_1406);
nor U2681 (N_2681,N_2338,N_1314);
nor U2682 (N_2682,N_1722,N_2302);
nor U2683 (N_2683,N_621,N_2020);
and U2684 (N_2684,N_991,N_745);
nand U2685 (N_2685,N_706,N_1617);
or U2686 (N_2686,N_1058,N_996);
nor U2687 (N_2687,N_365,N_2396);
and U2688 (N_2688,N_1399,N_2350);
nand U2689 (N_2689,N_2378,N_1949);
nand U2690 (N_2690,N_1132,N_2070);
or U2691 (N_2691,N_380,N_976);
and U2692 (N_2692,N_958,N_966);
nand U2693 (N_2693,N_954,N_22);
nand U2694 (N_2694,N_1522,N_1341);
or U2695 (N_2695,N_129,N_726);
or U2696 (N_2696,N_887,N_1353);
or U2697 (N_2697,N_2117,N_1288);
nor U2698 (N_2698,N_2366,N_1548);
nand U2699 (N_2699,N_1846,N_1092);
or U2700 (N_2700,N_1479,N_366);
or U2701 (N_2701,N_163,N_2003);
nor U2702 (N_2702,N_2088,N_1820);
nand U2703 (N_2703,N_1924,N_1895);
nor U2704 (N_2704,N_275,N_1512);
or U2705 (N_2705,N_769,N_1413);
and U2706 (N_2706,N_1799,N_1194);
nand U2707 (N_2707,N_1075,N_2360);
or U2708 (N_2708,N_1578,N_146);
or U2709 (N_2709,N_1861,N_1520);
and U2710 (N_2710,N_1872,N_1369);
nor U2711 (N_2711,N_2140,N_1378);
and U2712 (N_2712,N_883,N_1870);
or U2713 (N_2713,N_2081,N_1276);
and U2714 (N_2714,N_219,N_2417);
nor U2715 (N_2715,N_1985,N_72);
nor U2716 (N_2716,N_2353,N_2243);
nor U2717 (N_2717,N_1951,N_1993);
nand U2718 (N_2718,N_1616,N_263);
and U2719 (N_2719,N_1875,N_2013);
nand U2720 (N_2720,N_2109,N_432);
nor U2721 (N_2721,N_616,N_1319);
nand U2722 (N_2722,N_1984,N_233);
or U2723 (N_2723,N_655,N_1144);
nor U2724 (N_2724,N_689,N_13);
nor U2725 (N_2725,N_312,N_720);
and U2726 (N_2726,N_2489,N_674);
and U2727 (N_2727,N_1202,N_1580);
nand U2728 (N_2728,N_1865,N_1673);
nand U2729 (N_2729,N_2102,N_2254);
nor U2730 (N_2730,N_447,N_556);
xor U2731 (N_2731,N_1054,N_1905);
nor U2732 (N_2732,N_1783,N_1779);
or U2733 (N_2733,N_549,N_99);
and U2734 (N_2734,N_2475,N_438);
nor U2735 (N_2735,N_1254,N_1833);
or U2736 (N_2736,N_1751,N_784);
nand U2737 (N_2737,N_2403,N_1153);
and U2738 (N_2738,N_617,N_2409);
and U2739 (N_2739,N_10,N_2113);
xor U2740 (N_2740,N_1176,N_250);
xor U2741 (N_2741,N_1261,N_710);
nor U2742 (N_2742,N_1844,N_315);
and U2743 (N_2743,N_2253,N_1975);
or U2744 (N_2744,N_464,N_1091);
nand U2745 (N_2745,N_1037,N_2240);
or U2746 (N_2746,N_586,N_2039);
nor U2747 (N_2747,N_1995,N_1297);
and U2748 (N_2748,N_1055,N_1583);
nand U2749 (N_2749,N_1744,N_865);
nand U2750 (N_2750,N_656,N_2446);
nand U2751 (N_2751,N_1786,N_1734);
or U2752 (N_2752,N_2159,N_2000);
nand U2753 (N_2753,N_1372,N_2231);
nand U2754 (N_2754,N_1585,N_2457);
or U2755 (N_2755,N_1450,N_945);
nand U2756 (N_2756,N_646,N_1493);
or U2757 (N_2757,N_255,N_414);
or U2758 (N_2758,N_1445,N_113);
xnor U2759 (N_2759,N_162,N_1281);
nor U2760 (N_2760,N_2150,N_348);
and U2761 (N_2761,N_2084,N_337);
nand U2762 (N_2762,N_2189,N_256);
or U2763 (N_2763,N_1762,N_1518);
nor U2764 (N_2764,N_1477,N_665);
nor U2765 (N_2765,N_633,N_2087);
or U2766 (N_2766,N_1435,N_1736);
nor U2767 (N_2767,N_325,N_2429);
nand U2768 (N_2768,N_335,N_1486);
nand U2769 (N_2769,N_877,N_2157);
nand U2770 (N_2770,N_2328,N_2357);
and U2771 (N_2771,N_2064,N_201);
and U2772 (N_2772,N_1639,N_2250);
nand U2773 (N_2773,N_3,N_2278);
and U2774 (N_2774,N_615,N_2093);
nand U2775 (N_2775,N_1910,N_2288);
nand U2776 (N_2776,N_415,N_1971);
nand U2777 (N_2777,N_1523,N_433);
or U2778 (N_2778,N_1196,N_224);
or U2779 (N_2779,N_667,N_1652);
nor U2780 (N_2780,N_685,N_200);
nor U2781 (N_2781,N_618,N_378);
nand U2782 (N_2782,N_1816,N_102);
or U2783 (N_2783,N_1879,N_165);
nor U2784 (N_2784,N_1231,N_716);
nor U2785 (N_2785,N_1487,N_2026);
nand U2786 (N_2786,N_392,N_781);
or U2787 (N_2787,N_2308,N_1945);
nand U2788 (N_2788,N_248,N_1340);
nor U2789 (N_2789,N_338,N_1412);
and U2790 (N_2790,N_2079,N_1678);
nand U2791 (N_2791,N_2193,N_543);
and U2792 (N_2792,N_547,N_23);
nor U2793 (N_2793,N_2279,N_920);
nand U2794 (N_2794,N_1036,N_489);
nand U2795 (N_2795,N_539,N_481);
nor U2796 (N_2796,N_732,N_2395);
nor U2797 (N_2797,N_1606,N_1675);
xnor U2798 (N_2798,N_28,N_1748);
nand U2799 (N_2799,N_170,N_658);
and U2800 (N_2800,N_2337,N_1367);
and U2801 (N_2801,N_1623,N_2430);
or U2802 (N_2802,N_919,N_507);
or U2803 (N_2803,N_2319,N_175);
nor U2804 (N_2804,N_1347,N_605);
or U2805 (N_2805,N_1072,N_1211);
nor U2806 (N_2806,N_1576,N_158);
nand U2807 (N_2807,N_1253,N_296);
or U2808 (N_2808,N_100,N_770);
nand U2809 (N_2809,N_125,N_1697);
nand U2810 (N_2810,N_828,N_1246);
and U2811 (N_2811,N_1874,N_1465);
or U2812 (N_2812,N_332,N_1575);
and U2813 (N_2813,N_931,N_2325);
or U2814 (N_2814,N_1437,N_2420);
xnor U2815 (N_2815,N_1690,N_970);
xor U2816 (N_2816,N_1039,N_2251);
or U2817 (N_2817,N_1255,N_1655);
or U2818 (N_2818,N_2194,N_1627);
nand U2819 (N_2819,N_841,N_2323);
and U2820 (N_2820,N_2247,N_1760);
nor U2821 (N_2821,N_461,N_1338);
or U2822 (N_2822,N_1853,N_723);
xnor U2823 (N_2823,N_592,N_283);
or U2824 (N_2824,N_2218,N_252);
and U2825 (N_2825,N_1803,N_630);
and U2826 (N_2826,N_1368,N_379);
nand U2827 (N_2827,N_2398,N_1837);
nor U2828 (N_2828,N_1603,N_97);
nand U2829 (N_2829,N_2041,N_1100);
nand U2830 (N_2830,N_75,N_32);
nor U2831 (N_2831,N_2021,N_495);
and U2832 (N_2832,N_1883,N_1882);
nand U2833 (N_2833,N_36,N_2255);
nand U2834 (N_2834,N_87,N_230);
nor U2835 (N_2835,N_491,N_1699);
and U2836 (N_2836,N_1043,N_1703);
nor U2837 (N_2837,N_1152,N_1698);
and U2838 (N_2838,N_1514,N_2413);
nand U2839 (N_2839,N_2188,N_1442);
nor U2840 (N_2840,N_2207,N_1499);
nand U2841 (N_2841,N_1737,N_231);
and U2842 (N_2842,N_59,N_719);
nor U2843 (N_2843,N_1567,N_971);
or U2844 (N_2844,N_661,N_207);
or U2845 (N_2845,N_1088,N_1554);
nand U2846 (N_2846,N_1931,N_1960);
nand U2847 (N_2847,N_1671,N_441);
nand U2848 (N_2848,N_83,N_1063);
nand U2849 (N_2849,N_1299,N_1983);
nor U2850 (N_2850,N_1852,N_1770);
and U2851 (N_2851,N_2018,N_2340);
or U2852 (N_2852,N_2356,N_553);
nor U2853 (N_2853,N_1552,N_2059);
or U2854 (N_2854,N_875,N_451);
nand U2855 (N_2855,N_1784,N_560);
and U2856 (N_2856,N_171,N_843);
xnor U2857 (N_2857,N_1404,N_346);
xnor U2858 (N_2858,N_1103,N_2485);
or U2859 (N_2859,N_1559,N_1260);
nand U2860 (N_2860,N_176,N_550);
nor U2861 (N_2861,N_1197,N_222);
xnor U2862 (N_2862,N_1796,N_730);
nor U2863 (N_2863,N_1963,N_217);
or U2864 (N_2864,N_739,N_328);
nor U2865 (N_2865,N_2287,N_867);
nor U2866 (N_2866,N_2153,N_64);
nand U2867 (N_2867,N_1336,N_1008);
and U2868 (N_2868,N_1206,N_2491);
nand U2869 (N_2869,N_445,N_529);
xor U2870 (N_2870,N_2233,N_9);
nor U2871 (N_2871,N_1947,N_871);
and U2872 (N_2872,N_152,N_597);
xnor U2873 (N_2873,N_110,N_429);
nand U2874 (N_2874,N_1544,N_1009);
nand U2875 (N_2875,N_2346,N_1999);
or U2876 (N_2876,N_684,N_1621);
nor U2877 (N_2877,N_908,N_112);
or U2878 (N_2878,N_2451,N_1175);
nand U2879 (N_2879,N_557,N_1328);
or U2880 (N_2880,N_1531,N_1505);
nand U2881 (N_2881,N_2042,N_33);
and U2882 (N_2882,N_512,N_878);
and U2883 (N_2883,N_1205,N_1565);
and U2884 (N_2884,N_1948,N_2169);
or U2885 (N_2885,N_577,N_499);
nand U2886 (N_2886,N_551,N_700);
nor U2887 (N_2887,N_1785,N_1601);
and U2888 (N_2888,N_660,N_90);
and U2889 (N_2889,N_398,N_282);
or U2890 (N_2890,N_2133,N_1290);
nand U2891 (N_2891,N_2262,N_1302);
nand U2892 (N_2892,N_16,N_1238);
nor U2893 (N_2893,N_2322,N_260);
nor U2894 (N_2894,N_1452,N_1916);
nand U2895 (N_2895,N_1295,N_1222);
nand U2896 (N_2896,N_1012,N_1344);
nand U2897 (N_2897,N_2387,N_2397);
xor U2898 (N_2898,N_1687,N_1613);
nand U2899 (N_2899,N_1973,N_1052);
and U2900 (N_2900,N_2438,N_2479);
xnor U2901 (N_2901,N_1026,N_1539);
nand U2902 (N_2902,N_360,N_1904);
nand U2903 (N_2903,N_659,N_1952);
nor U2904 (N_2904,N_2160,N_1316);
xnor U2905 (N_2905,N_1379,N_405);
nand U2906 (N_2906,N_55,N_1199);
and U2907 (N_2907,N_1958,N_2347);
nor U2908 (N_2908,N_487,N_1941);
or U2909 (N_2909,N_758,N_2381);
and U2910 (N_2910,N_1660,N_369);
and U2911 (N_2911,N_2092,N_876);
and U2912 (N_2912,N_1656,N_2399);
nand U2913 (N_2913,N_1200,N_1475);
or U2914 (N_2914,N_2200,N_1953);
and U2915 (N_2915,N_2071,N_1223);
nor U2916 (N_2916,N_686,N_2239);
nand U2917 (N_2917,N_940,N_1178);
and U2918 (N_2918,N_866,N_174);
nor U2919 (N_2919,N_1889,N_1822);
and U2920 (N_2920,N_541,N_1772);
and U2921 (N_2921,N_2206,N_2342);
or U2922 (N_2922,N_1998,N_1659);
or U2923 (N_2923,N_1553,N_1533);
or U2924 (N_2924,N_1080,N_1618);
or U2925 (N_2925,N_587,N_1763);
and U2926 (N_2926,N_2364,N_1604);
nor U2927 (N_2927,N_2187,N_1277);
nor U2928 (N_2928,N_2471,N_1818);
or U2929 (N_2929,N_1997,N_2411);
nor U2930 (N_2930,N_2472,N_2168);
nor U2931 (N_2931,N_1562,N_2019);
nand U2932 (N_2932,N_1742,N_400);
or U2933 (N_2933,N_66,N_608);
and U2934 (N_2934,N_722,N_1396);
nor U2935 (N_2935,N_138,N_2326);
and U2936 (N_2936,N_1038,N_1573);
nor U2937 (N_2937,N_2495,N_852);
or U2938 (N_2938,N_2301,N_1296);
or U2939 (N_2939,N_2226,N_2023);
nor U2940 (N_2940,N_620,N_740);
nor U2941 (N_2941,N_1000,N_1279);
nand U2942 (N_2942,N_1672,N_611);
or U2943 (N_2943,N_698,N_929);
and U2944 (N_2944,N_1922,N_522);
nor U2945 (N_2945,N_1534,N_2220);
or U2946 (N_2946,N_2237,N_2031);
or U2947 (N_2947,N_388,N_1773);
nand U2948 (N_2948,N_670,N_840);
and U2949 (N_2949,N_679,N_1275);
or U2950 (N_2950,N_1992,N_51);
and U2951 (N_2951,N_1876,N_14);
nand U2952 (N_2952,N_1608,N_2336);
nand U2953 (N_2953,N_623,N_262);
nor U2954 (N_2954,N_1863,N_1258);
or U2955 (N_2955,N_704,N_2427);
nand U2956 (N_2956,N_1179,N_1859);
and U2957 (N_2957,N_436,N_1086);
nor U2958 (N_2958,N_2367,N_1159);
nor U2959 (N_2959,N_2468,N_1836);
or U2960 (N_2960,N_1688,N_1307);
nor U2961 (N_2961,N_1749,N_778);
nand U2962 (N_2962,N_1921,N_2123);
or U2963 (N_2963,N_71,N_155);
nor U2964 (N_2964,N_2418,N_717);
nand U2965 (N_2965,N_999,N_749);
or U2966 (N_2966,N_1677,N_316);
nor U2967 (N_2967,N_576,N_1017);
or U2968 (N_2968,N_2415,N_1237);
nand U2969 (N_2969,N_1716,N_2152);
nor U2970 (N_2970,N_1366,N_2432);
nor U2971 (N_2971,N_1428,N_1847);
or U2972 (N_2972,N_1765,N_1825);
or U2973 (N_2973,N_855,N_2131);
nand U2974 (N_2974,N_1775,N_2038);
or U2975 (N_2975,N_216,N_208);
nor U2976 (N_2976,N_2134,N_1754);
or U2977 (N_2977,N_1128,N_135);
nor U2978 (N_2978,N_77,N_1133);
or U2979 (N_2979,N_1624,N_2267);
nand U2980 (N_2980,N_1106,N_1902);
or U2981 (N_2981,N_2091,N_1858);
and U2982 (N_2982,N_1264,N_1764);
nand U2983 (N_2983,N_2400,N_638);
or U2984 (N_2984,N_820,N_1023);
nor U2985 (N_2985,N_393,N_40);
or U2986 (N_2986,N_1439,N_1930);
nor U2987 (N_2987,N_349,N_1704);
nor U2988 (N_2988,N_1142,N_2010);
or U2989 (N_2989,N_496,N_2496);
or U2990 (N_2990,N_2382,N_1972);
and U2991 (N_2991,N_1313,N_1337);
nor U2992 (N_2992,N_1572,N_844);
and U2993 (N_2993,N_1966,N_2143);
nand U2994 (N_2994,N_96,N_2055);
and U2995 (N_2995,N_381,N_2099);
nand U2996 (N_2996,N_1674,N_677);
nor U2997 (N_2997,N_1923,N_1429);
nand U2998 (N_2998,N_761,N_2173);
or U2999 (N_2999,N_649,N_1431);
nor U3000 (N_3000,N_462,N_1915);
and U3001 (N_3001,N_2412,N_1228);
nor U3002 (N_3002,N_247,N_886);
or U3003 (N_3003,N_682,N_1105);
or U3004 (N_3004,N_736,N_2389);
and U3005 (N_3005,N_2100,N_800);
and U3006 (N_3006,N_1459,N_1550);
nor U3007 (N_3007,N_1629,N_418);
or U3008 (N_3008,N_1416,N_1917);
nand U3009 (N_3009,N_1409,N_106);
or U3010 (N_3010,N_375,N_1181);
nor U3011 (N_3011,N_1259,N_1702);
nand U3012 (N_3012,N_2139,N_997);
and U3013 (N_3013,N_1121,N_2466);
nor U3014 (N_3014,N_1138,N_554);
or U3015 (N_3015,N_641,N_1434);
and U3016 (N_3016,N_377,N_459);
and U3017 (N_3017,N_1938,N_1605);
or U3018 (N_3018,N_2029,N_1934);
nand U3019 (N_3019,N_1735,N_1311);
or U3020 (N_3020,N_2390,N_478);
nor U3021 (N_3021,N_494,N_2221);
nand U3022 (N_3022,N_562,N_1304);
nor U3023 (N_3023,N_1383,N_116);
nand U3024 (N_3024,N_901,N_2434);
and U3025 (N_3025,N_822,N_1136);
nand U3026 (N_3026,N_2377,N_1028);
nand U3027 (N_3027,N_1756,N_1828);
nor U3028 (N_3028,N_1897,N_536);
or U3029 (N_3029,N_1586,N_26);
nand U3030 (N_3030,N_2135,N_785);
nand U3031 (N_3031,N_2470,N_752);
nor U3032 (N_3032,N_708,N_1393);
nand U3033 (N_3033,N_930,N_440);
and U3034 (N_3034,N_2112,N_1890);
or U3035 (N_3035,N_924,N_2391);
and U3036 (N_3036,N_1593,N_2242);
and U3037 (N_3037,N_1001,N_156);
nor U3038 (N_3038,N_237,N_1630);
nand U3039 (N_3039,N_427,N_1292);
nor U3040 (N_3040,N_2260,N_49);
nor U3041 (N_3041,N_329,N_147);
or U3042 (N_3042,N_2459,N_1115);
nand U3043 (N_3043,N_1549,N_1758);
nor U3044 (N_3044,N_229,N_728);
nand U3045 (N_3045,N_1778,N_2303);
or U3046 (N_3046,N_790,N_460);
nor U3047 (N_3047,N_1880,N_1806);
nand U3048 (N_3048,N_1183,N_408);
or U3049 (N_3049,N_190,N_727);
or U3050 (N_3050,N_747,N_2329);
and U3051 (N_3051,N_959,N_1195);
or U3052 (N_3052,N_1503,N_1289);
nor U3053 (N_3053,N_1650,N_1352);
or U3054 (N_3054,N_1240,N_2355);
nor U3055 (N_3055,N_835,N_1829);
xor U3056 (N_3056,N_195,N_1423);
or U3057 (N_3057,N_362,N_303);
or U3058 (N_3058,N_1458,N_1885);
nor U3059 (N_3059,N_1190,N_1911);
nand U3060 (N_3060,N_1168,N_417);
nand U3061 (N_3061,N_180,N_542);
and U3062 (N_3062,N_1112,N_1691);
and U3063 (N_3063,N_2372,N_2258);
nand U3064 (N_3064,N_2339,N_2030);
and U3065 (N_3065,N_1362,N_645);
or U3066 (N_3066,N_1819,N_1940);
nor U3067 (N_3067,N_1743,N_2151);
nand U3068 (N_3068,N_2068,N_123);
nor U3069 (N_3069,N_2358,N_631);
and U3070 (N_3070,N_1638,N_1118);
and U3071 (N_3071,N_1448,N_653);
xnor U3072 (N_3072,N_1654,N_2297);
and U3073 (N_3073,N_2138,N_1403);
nand U3074 (N_3074,N_108,N_191);
nand U3075 (N_3075,N_2435,N_848);
nand U3076 (N_3076,N_2137,N_1407);
nor U3077 (N_3077,N_466,N_401);
and U3078 (N_3078,N_2161,N_89);
and U3079 (N_3079,N_526,N_982);
nor U3080 (N_3080,N_760,N_2191);
nand U3081 (N_3081,N_909,N_2110);
and U3082 (N_3082,N_2345,N_1810);
and U3083 (N_3083,N_537,N_1723);
nand U3084 (N_3084,N_2155,N_799);
nor U3085 (N_3085,N_1517,N_2141);
nand U3086 (N_3086,N_1234,N_1651);
or U3087 (N_3087,N_2204,N_1286);
nor U3088 (N_3088,N_1950,N_1711);
nand U3089 (N_3089,N_1658,N_134);
nor U3090 (N_3090,N_1474,N_2383);
nand U3091 (N_3091,N_2487,N_2265);
and U3092 (N_3092,N_1361,N_729);
nor U3093 (N_3093,N_1789,N_41);
nor U3094 (N_3094,N_816,N_510);
and U3095 (N_3095,N_1268,N_412);
or U3096 (N_3096,N_821,N_1345);
nand U3097 (N_3097,N_94,N_2317);
nand U3098 (N_3098,N_910,N_794);
nor U3099 (N_3099,N_149,N_652);
nand U3100 (N_3100,N_1502,N_1684);
nor U3101 (N_3101,N_358,N_1294);
nand U3102 (N_3102,N_357,N_213);
nor U3103 (N_3103,N_1157,N_2343);
nand U3104 (N_3104,N_1174,N_69);
or U3105 (N_3105,N_1537,N_1169);
nor U3106 (N_3106,N_437,N_687);
and U3107 (N_3107,N_1926,N_1391);
and U3108 (N_3108,N_2089,N_1024);
and U3109 (N_3109,N_1862,N_972);
nor U3110 (N_3110,N_981,N_1964);
and U3111 (N_3111,N_95,N_1123);
or U3112 (N_3112,N_614,N_1117);
nor U3113 (N_3113,N_2270,N_2443);
and U3114 (N_3114,N_1208,N_220);
and U3115 (N_3115,N_642,N_105);
nor U3116 (N_3116,N_1099,N_1250);
nand U3117 (N_3117,N_2002,N_136);
nor U3118 (N_3118,N_1415,N_635);
and U3119 (N_3119,N_2499,N_839);
and U3120 (N_3120,N_1597,N_104);
nand U3121 (N_3121,N_1184,N_888);
nand U3122 (N_3122,N_1628,N_1320);
nor U3123 (N_3123,N_1719,N_1478);
nand U3124 (N_3124,N_2186,N_144);
and U3125 (N_3125,N_584,N_2299);
and U3126 (N_3126,N_705,N_563);
or U3127 (N_3127,N_274,N_1694);
and U3128 (N_3128,N_2078,N_1332);
or U3129 (N_3129,N_2458,N_1670);
nand U3130 (N_3130,N_76,N_306);
and U3131 (N_3131,N_1591,N_788);
nor U3132 (N_3132,N_753,N_1526);
and U3133 (N_3133,N_1823,N_1595);
nor U3134 (N_3134,N_899,N_1705);
or U3135 (N_3135,N_1579,N_804);
and U3136 (N_3136,N_1888,N_995);
nand U3137 (N_3137,N_1724,N_1635);
or U3138 (N_3138,N_1571,N_825);
or U3139 (N_3139,N_1750,N_2309);
or U3140 (N_3140,N_1532,N_1974);
or U3141 (N_3141,N_1171,N_2172);
nand U3142 (N_3142,N_1536,N_280);
nand U3143 (N_3143,N_1661,N_1759);
nand U3144 (N_3144,N_1060,N_1557);
or U3145 (N_3145,N_114,N_776);
and U3146 (N_3146,N_317,N_2097);
nor U3147 (N_3147,N_1619,N_2401);
and U3148 (N_3148,N_2069,N_409);
nand U3149 (N_3149,N_1851,N_818);
nand U3150 (N_3150,N_854,N_850);
and U3151 (N_3151,N_579,N_387);
or U3152 (N_3152,N_57,N_980);
or U3153 (N_3153,N_1800,N_1317);
nor U3154 (N_3154,N_1731,N_2283);
nand U3155 (N_3155,N_261,N_905);
nor U3156 (N_3156,N_768,N_1632);
nor U3157 (N_3157,N_591,N_444);
and U3158 (N_3158,N_756,N_1020);
or U3159 (N_3159,N_973,N_1791);
nand U3160 (N_3160,N_1664,N_651);
nor U3161 (N_3161,N_353,N_1521);
or U3162 (N_3162,N_2442,N_535);
nand U3163 (N_3163,N_2271,N_1140);
and U3164 (N_3164,N_2101,N_1443);
or U3165 (N_3165,N_1994,N_872);
and U3166 (N_3166,N_1602,N_1494);
and U3167 (N_3167,N_320,N_731);
and U3168 (N_3168,N_846,N_183);
xor U3169 (N_3169,N_1400,N_1104);
nand U3170 (N_3170,N_714,N_1248);
nand U3171 (N_3171,N_2392,N_1303);
nor U3172 (N_3172,N_1212,N_518);
and U3173 (N_3173,N_448,N_2190);
nand U3174 (N_3174,N_1472,N_1387);
nor U3175 (N_3175,N_351,N_525);
and U3176 (N_3176,N_368,N_1158);
nor U3177 (N_3177,N_2290,N_2048);
and U3178 (N_3178,N_1137,N_20);
nor U3179 (N_3179,N_1321,N_1385);
and U3180 (N_3180,N_1278,N_2044);
and U3181 (N_3181,N_430,N_340);
xnor U3182 (N_3182,N_2144,N_1584);
or U3183 (N_3183,N_791,N_2407);
and U3184 (N_3184,N_2011,N_2428);
or U3185 (N_3185,N_1787,N_2224);
or U3186 (N_3186,N_223,N_2054);
or U3187 (N_3187,N_1781,N_265);
or U3188 (N_3188,N_2066,N_1692);
and U3189 (N_3189,N_935,N_2404);
nor U3190 (N_3190,N_1936,N_2437);
and U3191 (N_3191,N_1986,N_443);
or U3192 (N_3192,N_1257,N_1489);
or U3193 (N_3193,N_798,N_2005);
nand U3194 (N_3194,N_1419,N_1375);
and U3195 (N_3195,N_2198,N_1323);
nand U3196 (N_3196,N_292,N_968);
nand U3197 (N_3197,N_1484,N_1817);
and U3198 (N_3198,N_1388,N_1421);
and U3199 (N_3199,N_141,N_1809);
or U3200 (N_3200,N_1740,N_1007);
and U3201 (N_3201,N_609,N_1401);
and U3202 (N_3202,N_407,N_911);
and U3203 (N_3203,N_1476,N_1031);
or U3204 (N_3204,N_371,N_1831);
and U3205 (N_3205,N_533,N_914);
nand U3206 (N_3206,N_1180,N_517);
nand U3207 (N_3207,N_1414,N_524);
or U3208 (N_3208,N_898,N_2058);
or U3209 (N_3209,N_1422,N_826);
nand U3210 (N_3210,N_1358,N_1076);
nand U3211 (N_3211,N_1987,N_1035);
and U3212 (N_3212,N_897,N_1826);
and U3213 (N_3213,N_2422,N_1093);
xor U3214 (N_3214,N_602,N_382);
and U3215 (N_3215,N_1047,N_299);
or U3216 (N_3216,N_1364,N_2314);
or U3217 (N_3217,N_1961,N_552);
or U3218 (N_3218,N_933,N_808);
xor U3219 (N_3219,N_1239,N_1267);
and U3220 (N_3220,N_1284,N_1793);
or U3221 (N_3221,N_1351,N_1470);
nand U3222 (N_3222,N_1051,N_1411);
nor U3223 (N_3223,N_892,N_1790);
nor U3224 (N_3224,N_814,N_425);
or U3225 (N_3225,N_1871,N_1069);
or U3226 (N_3226,N_950,N_666);
nor U3227 (N_3227,N_1209,N_902);
nand U3228 (N_3228,N_467,N_498);
nor U3229 (N_3229,N_594,N_748);
or U3230 (N_3230,N_1551,N_1084);
or U3231 (N_3231,N_960,N_140);
nor U3232 (N_3232,N_1797,N_585);
and U3233 (N_3233,N_179,N_521);
and U3234 (N_3234,N_2006,N_1841);
and U3235 (N_3235,N_650,N_1436);
and U3236 (N_3236,N_565,N_259);
nand U3237 (N_3237,N_984,N_856);
or U3238 (N_3238,N_1027,N_2361);
nand U3239 (N_3239,N_927,N_1668);
and U3240 (N_3240,N_177,N_1430);
or U3241 (N_3241,N_857,N_1855);
nand U3242 (N_3242,N_2256,N_206);
or U3243 (N_3243,N_1218,N_391);
nand U3244 (N_3244,N_1167,N_268);
nand U3245 (N_3245,N_115,N_1373);
or U3246 (N_3246,N_2375,N_61);
nor U3247 (N_3247,N_2269,N_531);
nand U3248 (N_3248,N_715,N_376);
and U3249 (N_3249,N_1877,N_805);
nand U3250 (N_3250,N_85,N_1166);
and U3251 (N_3251,N_1718,N_1811);
or U3252 (N_3252,N_622,N_824);
nand U3253 (N_3253,N_907,N_900);
nand U3254 (N_3254,N_889,N_1588);
nor U3255 (N_3255,N_356,N_2049);
and U3256 (N_3256,N_471,N_1955);
nand U3257 (N_3257,N_1600,N_2484);
or U3258 (N_3258,N_569,N_2202);
nand U3259 (N_3259,N_446,N_509);
and U3260 (N_3260,N_1154,N_965);
nand U3261 (N_3261,N_1151,N_1);
nand U3262 (N_3262,N_1219,N_923);
and U3263 (N_3263,N_1079,N_2025);
xnor U3264 (N_3264,N_1046,N_2056);
and U3265 (N_3265,N_1566,N_640);
nor U3266 (N_3266,N_2046,N_1418);
and U3267 (N_3267,N_2333,N_1568);
xor U3268 (N_3268,N_2431,N_755);
nor U3269 (N_3269,N_2047,N_1807);
nor U3270 (N_3270,N_167,N_1929);
and U3271 (N_3271,N_863,N_1210);
nand U3272 (N_3272,N_497,N_1440);
or U3273 (N_3273,N_321,N_2332);
or U3274 (N_3274,N_1939,N_1053);
nor U3275 (N_3275,N_2040,N_948);
nor U3276 (N_3276,N_1013,N_2341);
and U3277 (N_3277,N_192,N_2294);
xnor U3278 (N_3278,N_1657,N_2106);
xor U3279 (N_3279,N_2497,N_1141);
nand U3280 (N_3280,N_506,N_1777);
nor U3281 (N_3281,N_1558,N_572);
nor U3282 (N_3282,N_1881,N_293);
or U3283 (N_3283,N_2063,N_2473);
nor U3284 (N_3284,N_477,N_1845);
and U3285 (N_3285,N_1513,N_743);
and U3286 (N_3286,N_1149,N_975);
nor U3287 (N_3287,N_2122,N_124);
nor U3288 (N_3288,N_2324,N_1125);
or U3289 (N_3289,N_2235,N_194);
nand U3290 (N_3290,N_500,N_2185);
nand U3291 (N_3291,N_48,N_2405);
and U3292 (N_3292,N_2142,N_1497);
nor U3293 (N_3293,N_1988,N_1309);
and U3294 (N_3294,N_39,N_2196);
nor U3295 (N_3295,N_1538,N_2177);
nor U3296 (N_3296,N_1977,N_2433);
nand U3297 (N_3297,N_559,N_1130);
and U3298 (N_3298,N_1334,N_58);
and U3299 (N_3299,N_1061,N_395);
and U3300 (N_3300,N_873,N_595);
or U3301 (N_3301,N_188,N_2320);
or U3302 (N_3302,N_1301,N_2234);
and U3303 (N_3303,N_789,N_829);
nor U3304 (N_3304,N_2274,N_1360);
nor U3305 (N_3305,N_2257,N_1683);
or U3306 (N_3306,N_1049,N_1357);
or U3307 (N_3307,N_127,N_86);
nor U3308 (N_3308,N_285,N_2419);
nand U3309 (N_3309,N_384,N_1893);
or U3310 (N_3310,N_567,N_251);
and U3311 (N_3311,N_1087,N_294);
or U3312 (N_3312,N_1417,N_1160);
nor U3313 (N_3313,N_1729,N_1739);
nand U3314 (N_3314,N_218,N_1410);
nor U3315 (N_3315,N_434,N_8);
or U3316 (N_3316,N_2050,N_610);
and U3317 (N_3317,N_1456,N_648);
nor U3318 (N_3318,N_1610,N_2214);
nand U3319 (N_3319,N_1064,N_815);
and U3320 (N_3320,N_2147,N_1298);
nor U3321 (N_3321,N_485,N_455);
xor U3322 (N_3322,N_1122,N_107);
or U3323 (N_3323,N_672,N_486);
nand U3324 (N_3324,N_1900,N_1891);
nand U3325 (N_3325,N_528,N_1389);
or U3326 (N_3326,N_590,N_1164);
and U3327 (N_3327,N_2004,N_1581);
xor U3328 (N_3328,N_67,N_2057);
or U3329 (N_3329,N_73,N_1395);
and U3330 (N_3330,N_454,N_1438);
or U3331 (N_3331,N_1633,N_2146);
or U3332 (N_3332,N_1172,N_1186);
nand U3333 (N_3333,N_1981,N_636);
nand U3334 (N_3334,N_273,N_1390);
nor U3335 (N_3335,N_1814,N_196);
and U3336 (N_3336,N_1188,N_2232);
nor U3337 (N_3337,N_1330,N_1343);
and U3338 (N_3338,N_119,N_210);
nor U3339 (N_3339,N_420,N_2465);
xnor U3340 (N_3340,N_695,N_823);
and U3341 (N_3341,N_1564,N_2107);
nor U3342 (N_3342,N_240,N_1370);
and U3343 (N_3343,N_355,N_2463);
xor U3344 (N_3344,N_334,N_449);
or U3345 (N_3345,N_1866,N_1596);
nand U3346 (N_3346,N_399,N_890);
nand U3347 (N_3347,N_1018,N_2455);
nor U3348 (N_3348,N_139,N_943);
nor U3349 (N_3349,N_241,N_1094);
nand U3350 (N_3350,N_2277,N_1173);
nor U3351 (N_3351,N_270,N_2128);
and U3352 (N_3352,N_131,N_1192);
or U3353 (N_3353,N_1146,N_1492);
and U3354 (N_3354,N_1096,N_164);
nor U3355 (N_3355,N_2488,N_765);
and U3356 (N_3356,N_249,N_111);
nand U3357 (N_3357,N_859,N_62);
nor U3358 (N_3358,N_2362,N_1519);
and U3359 (N_3359,N_1899,N_936);
or U3360 (N_3360,N_2321,N_1333);
or U3361 (N_3361,N_1235,N_238);
and U3362 (N_3362,N_953,N_327);
nand U3363 (N_3363,N_2273,N_1693);
and U3364 (N_3364,N_2033,N_453);
nor U3365 (N_3365,N_2095,N_718);
and U3366 (N_3366,N_1782,N_1225);
nor U3367 (N_3367,N_2266,N_1937);
and U3368 (N_3368,N_2281,N_922);
or U3369 (N_3369,N_1969,N_1867);
and U3370 (N_3370,N_2181,N_2072);
or U3371 (N_3371,N_1528,N_1496);
and U3372 (N_3372,N_1515,N_2126);
and U3373 (N_3373,N_2285,N_269);
nor U3374 (N_3374,N_2312,N_757);
or U3375 (N_3375,N_2318,N_1156);
nand U3376 (N_3376,N_1634,N_65);
or U3377 (N_3377,N_2195,N_1560);
xnor U3378 (N_3378,N_697,N_944);
nor U3379 (N_3379,N_891,N_2478);
nor U3380 (N_3380,N_1753,N_271);
nand U3381 (N_3381,N_879,N_504);
nor U3382 (N_3382,N_145,N_2306);
or U3383 (N_3383,N_811,N_239);
or U3384 (N_3384,N_1363,N_1381);
or U3385 (N_3385,N_2154,N_1767);
or U3386 (N_3386,N_359,N_693);
or U3387 (N_3387,N_1516,N_2213);
nand U3388 (N_3388,N_2327,N_2244);
nor U3389 (N_3389,N_746,N_46);
nand U3390 (N_3390,N_1005,N_331);
or U3391 (N_3391,N_2118,N_226);
and U3392 (N_3392,N_1059,N_1244);
and U3393 (N_3393,N_5,N_2149);
or U3394 (N_3394,N_1048,N_281);
nand U3395 (N_3395,N_2464,N_2125);
xor U3396 (N_3396,N_2483,N_354);
nor U3397 (N_3397,N_2045,N_2219);
and U3398 (N_3398,N_2263,N_12);
nand U3399 (N_3399,N_2423,N_2120);
nand U3400 (N_3400,N_956,N_168);
nor U3401 (N_3401,N_56,N_2024);
or U3402 (N_3402,N_82,N_978);
or U3403 (N_3403,N_1590,N_607);
nor U3404 (N_3404,N_1095,N_2121);
and U3405 (N_3405,N_1424,N_225);
or U3406 (N_3406,N_2456,N_1609);
nor U3407 (N_3407,N_2037,N_2105);
and U3408 (N_3408,N_1189,N_1120);
or U3409 (N_3409,N_625,N_2119);
nand U3410 (N_3410,N_29,N_372);
or U3411 (N_3411,N_1556,N_1420);
and U3412 (N_3412,N_1906,N_1495);
nor U3413 (N_3413,N_1842,N_2467);
nor U3414 (N_3414,N_699,N_185);
and U3415 (N_3415,N_939,N_1374);
nand U3416 (N_3416,N_1830,N_2171);
nor U3417 (N_3417,N_775,N_1850);
or U3418 (N_3418,N_142,N_885);
and U3419 (N_3419,N_792,N_2076);
nand U3420 (N_3420,N_2248,N_1090);
nand U3421 (N_3421,N_774,N_1620);
and U3422 (N_3422,N_1913,N_511);
or U3423 (N_3423,N_1453,N_2334);
or U3424 (N_3424,N_103,N_2276);
nor U3425 (N_3425,N_1365,N_2492);
nand U3426 (N_3426,N_7,N_74);
nor U3427 (N_3427,N_964,N_1849);
nor U3428 (N_3428,N_2065,N_1491);
nand U3429 (N_3429,N_2368,N_1350);
nand U3430 (N_3430,N_558,N_810);
or U3431 (N_3431,N_601,N_1467);
nor U3432 (N_3432,N_1215,N_1346);
and U3433 (N_3433,N_221,N_245);
nand U3434 (N_3434,N_932,N_150);
or U3435 (N_3435,N_596,N_1569);
xnor U3436 (N_3436,N_397,N_1074);
nor U3437 (N_3437,N_2474,N_157);
nor U3438 (N_3438,N_2209,N_837);
and U3439 (N_3439,N_2482,N_951);
or U3440 (N_3440,N_1701,N_967);
and U3441 (N_3441,N_1615,N_845);
and U3442 (N_3442,N_721,N_2481);
nand U3443 (N_3443,N_881,N_1116);
or U3444 (N_3444,N_284,N_2016);
and U3445 (N_3445,N_673,N_1884);
or U3446 (N_3446,N_992,N_323);
and U3447 (N_3447,N_242,N_2307);
nand U3448 (N_3448,N_513,N_1794);
nor U3449 (N_3449,N_182,N_1682);
or U3450 (N_3450,N_439,N_1801);
nor U3451 (N_3451,N_827,N_662);
or U3452 (N_3452,N_345,N_2424);
or U3453 (N_3453,N_2445,N_2228);
xor U3454 (N_3454,N_1441,N_1067);
and U3455 (N_3455,N_428,N_2074);
or U3456 (N_3456,N_1746,N_994);
or U3457 (N_3457,N_1312,N_480);
or U3458 (N_3458,N_1766,N_1376);
nor U3459 (N_3459,N_297,N_2374);
nand U3460 (N_3460,N_571,N_1498);
nand U3461 (N_3461,N_2436,N_2211);
xnor U3462 (N_3462,N_1354,N_2164);
or U3463 (N_3463,N_1509,N_18);
or U3464 (N_3464,N_151,N_1843);
nor U3465 (N_3465,N_1978,N_314);
nand U3466 (N_3466,N_1214,N_2351);
or U3467 (N_3467,N_690,N_1155);
nor U3468 (N_3468,N_279,N_1033);
and U3469 (N_3469,N_2454,N_1592);
nand U3470 (N_3470,N_456,N_2227);
nand U3471 (N_3471,N_979,N_1481);
or U3472 (N_3472,N_1460,N_1129);
or U3473 (N_3473,N_1335,N_1827);
nor U3474 (N_3474,N_2369,N_1229);
and U3475 (N_3475,N_735,N_1108);
nand U3476 (N_3476,N_130,N_1959);
and U3477 (N_3477,N_287,N_1127);
and U3478 (N_3478,N_2158,N_286);
nand U3479 (N_3479,N_1102,N_468);
and U3480 (N_3480,N_2,N_1886);
and U3481 (N_3481,N_1506,N_435);
nand U3482 (N_3482,N_1649,N_413);
and U3483 (N_3483,N_342,N_1300);
nor U3484 (N_3484,N_555,N_1856);
nand U3485 (N_3485,N_2008,N_581);
or U3486 (N_3486,N_92,N_2410);
nor U3487 (N_3487,N_786,N_2162);
or U3488 (N_3488,N_68,N_215);
nand U3489 (N_3489,N_1324,N_1201);
nand U3490 (N_3490,N_505,N_668);
and U3491 (N_3491,N_880,N_762);
nand U3492 (N_3492,N_2192,N_322);
or U3493 (N_3493,N_1732,N_2127);
nand U3494 (N_3494,N_21,N_2130);
nand U3495 (N_3495,N_2296,N_1928);
nand U3496 (N_3496,N_1641,N_442);
or U3497 (N_3497,N_2388,N_2448);
or U3498 (N_3498,N_173,N_1163);
nor U3499 (N_3499,N_1462,N_181);
nand U3500 (N_3500,N_1077,N_759);
or U3501 (N_3501,N_267,N_2075);
or U3502 (N_3502,N_80,N_1504);
nand U3503 (N_3503,N_1976,N_1798);
xnor U3504 (N_3504,N_484,N_1040);
or U3505 (N_3505,N_1667,N_2365);
or U3506 (N_3506,N_540,N_416);
or U3507 (N_3507,N_1359,N_946);
or U3508 (N_3508,N_266,N_1543);
nand U3509 (N_3509,N_508,N_1454);
or U3510 (N_3510,N_683,N_1612);
and U3511 (N_3511,N_1728,N_2053);
nand U3512 (N_3512,N_1056,N_1468);
or U3513 (N_3513,N_754,N_1755);
nand U3514 (N_3514,N_1220,N_2015);
and U3515 (N_3515,N_2216,N_1025);
or U3516 (N_3516,N_258,N_488);
nor U3517 (N_3517,N_1232,N_1535);
and U3518 (N_3518,N_2179,N_493);
and U3519 (N_3519,N_1098,N_161);
or U3520 (N_3520,N_389,N_2439);
nand U3521 (N_3521,N_386,N_703);
nand U3522 (N_3522,N_383,N_1490);
and U3523 (N_3523,N_701,N_990);
nand U3524 (N_3524,N_2116,N_209);
nor U3525 (N_3525,N_2166,N_830);
and U3526 (N_3526,N_741,N_1996);
nand U3527 (N_3527,N_1686,N_2184);
nand U3528 (N_3528,N_122,N_277);
and U3529 (N_3529,N_1283,N_941);
nand U3530 (N_3530,N_538,N_712);
or U3531 (N_3531,N_570,N_952);
and U3532 (N_3532,N_1919,N_1329);
or U3533 (N_3533,N_643,N_1561);
and U3534 (N_3534,N_2017,N_2210);
nor U3535 (N_3535,N_1868,N_2086);
nor U3536 (N_3536,N_1848,N_986);
or U3537 (N_3537,N_1860,N_276);
and U3538 (N_3538,N_1662,N_385);
or U3539 (N_3539,N_1262,N_333);
and U3540 (N_3540,N_2498,N_2335);
or U3541 (N_3541,N_1318,N_803);
nand U3542 (N_3542,N_1574,N_1170);
or U3543 (N_3543,N_869,N_1507);
and U3544 (N_3544,N_2316,N_406);
nor U3545 (N_3545,N_492,N_81);
nand U3546 (N_3546,N_109,N_2085);
nand U3547 (N_3547,N_1006,N_1293);
nand U3548 (N_3548,N_2282,N_302);
nor U3549 (N_3549,N_212,N_831);
or U3550 (N_3550,N_53,N_1089);
and U3551 (N_3551,N_1887,N_431);
nand U3552 (N_3552,N_1813,N_1944);
nand U3553 (N_3553,N_2229,N_1325);
and U3554 (N_3554,N_1322,N_324);
nand U3555 (N_3555,N_1636,N_2246);
or U3556 (N_3556,N_1216,N_1607);
or U3557 (N_3557,N_473,N_1377);
or U3558 (N_3558,N_750,N_2440);
and U3559 (N_3559,N_657,N_350);
nand U3560 (N_3560,N_1145,N_1185);
or U3561 (N_3561,N_343,N_1525);
nand U3562 (N_3562,N_1305,N_1233);
nand U3563 (N_3563,N_330,N_1256);
nor U3564 (N_3564,N_1792,N_2385);
nand U3565 (N_3565,N_2034,N_819);
nor U3566 (N_3566,N_564,N_724);
nor U3567 (N_3567,N_1542,N_301);
nor U3568 (N_3568,N_1243,N_272);
or U3569 (N_3569,N_874,N_403);
or U3570 (N_3570,N_2295,N_503);
or U3571 (N_3571,N_1249,N_1464);
nand U3572 (N_3572,N_858,N_2180);
nand U3573 (N_3573,N_957,N_1582);
or U3574 (N_3574,N_1004,N_404);
and U3575 (N_3575,N_530,N_2175);
nor U3576 (N_3576,N_2408,N_1598);
or U3577 (N_3577,N_1696,N_2376);
and U3578 (N_3578,N_832,N_311);
xnor U3579 (N_3579,N_474,N_1397);
and U3580 (N_3580,N_1070,N_1348);
nand U3581 (N_3581,N_696,N_787);
and U3582 (N_3582,N_1854,N_44);
nand U3583 (N_3583,N_2402,N_1065);
or U3584 (N_3584,N_1989,N_903);
and U3585 (N_3585,N_1643,N_1394);
and U3586 (N_3586,N_675,N_1680);
nand U3587 (N_3587,N_153,N_1193);
nand U3588 (N_3588,N_2090,N_1980);
nor U3589 (N_3589,N_2486,N_117);
or U3590 (N_3590,N_2073,N_422);
nor U3591 (N_3591,N_2460,N_2174);
nor U3592 (N_3592,N_2386,N_1935);
nand U3593 (N_3593,N_1042,N_199);
and U3594 (N_3594,N_126,N_2298);
nor U3595 (N_3595,N_1165,N_1252);
nand U3596 (N_3596,N_771,N_921);
nor U3597 (N_3597,N_1587,N_1213);
nand U3598 (N_3598,N_1382,N_1150);
nor U3599 (N_3599,N_2449,N_918);
nand U3600 (N_3600,N_1642,N_2124);
and U3601 (N_3601,N_1245,N_568);
or U3602 (N_3602,N_1327,N_421);
nor U3603 (N_3603,N_1204,N_2230);
or U3604 (N_3604,N_1014,N_2061);
nand U3605 (N_3605,N_1291,N_2208);
or U3606 (N_3606,N_2178,N_955);
or U3607 (N_3607,N_534,N_1433);
nor U3608 (N_3608,N_2363,N_364);
nand U3609 (N_3609,N_1563,N_54);
or U3610 (N_3610,N_214,N_336);
nor U3611 (N_3611,N_1918,N_516);
nor U3612 (N_3612,N_88,N_626);
or U3613 (N_3613,N_884,N_813);
nand U3614 (N_3614,N_187,N_680);
nor U3615 (N_3615,N_2447,N_1611);
or U3616 (N_3616,N_1815,N_782);
and U3617 (N_3617,N_764,N_916);
nor U3618 (N_3618,N_604,N_2028);
or U3619 (N_3619,N_291,N_654);
xor U3620 (N_3620,N_1808,N_1405);
xnor U3621 (N_3621,N_2349,N_2259);
xor U3622 (N_3622,N_2217,N_120);
and U3623 (N_3623,N_988,N_1727);
and U3624 (N_3624,N_1126,N_1745);
xor U3625 (N_3625,N_1010,N_777);
and U3626 (N_3626,N_812,N_202);
nand U3627 (N_3627,N_1473,N_1717);
nand U3628 (N_3628,N_166,N_520);
or U3629 (N_3629,N_664,N_2103);
xnor U3630 (N_3630,N_502,N_860);
nor U3631 (N_3631,N_1547,N_1273);
nor U3632 (N_3632,N_227,N_1666);
or U3633 (N_3633,N_1625,N_2148);
nor U3634 (N_3634,N_593,N_1427);
or U3635 (N_3635,N_172,N_458);
nor U3636 (N_3636,N_2371,N_1221);
and U3637 (N_3637,N_2315,N_1471);
and U3638 (N_3638,N_1451,N_341);
nand U3639 (N_3639,N_2280,N_2393);
nor U3640 (N_3640,N_532,N_2098);
or U3641 (N_3641,N_588,N_1107);
and U3642 (N_3642,N_2080,N_309);
xnor U3643 (N_3643,N_1708,N_1925);
or U3644 (N_3644,N_707,N_367);
nor U3645 (N_3645,N_1707,N_178);
nor U3646 (N_3646,N_1485,N_1386);
and U3647 (N_3647,N_1640,N_734);
nand U3648 (N_3648,N_711,N_2223);
nor U3649 (N_3649,N_834,N_1482);
or U3650 (N_3650,N_1909,N_1933);
nor U3651 (N_3651,N_676,N_2052);
or U3652 (N_3652,N_598,N_235);
or U3653 (N_3653,N_691,N_2289);
or U3654 (N_3654,N_613,N_1447);
nor U3655 (N_3655,N_423,N_926);
nor U3656 (N_3656,N_2012,N_1927);
nor U3657 (N_3657,N_1709,N_1878);
and U3658 (N_3658,N_2450,N_2476);
nand U3659 (N_3659,N_1761,N_318);
nor U3660 (N_3660,N_1869,N_1713);
nand U3661 (N_3661,N_1747,N_1780);
nor U3662 (N_3662,N_132,N_1812);
or U3663 (N_3663,N_751,N_678);
or U3664 (N_3664,N_98,N_1903);
nor U3665 (N_3665,N_582,N_938);
and U3666 (N_3666,N_1203,N_1527);
nor U3667 (N_3667,N_546,N_228);
nand U3668 (N_3668,N_1594,N_895);
nand U3669 (N_3669,N_307,N_1073);
nand U3670 (N_3670,N_575,N_70);
or U3671 (N_3671,N_807,N_1355);
and U3672 (N_3672,N_849,N_476);
nor U3673 (N_3673,N_402,N_313);
or U3674 (N_3674,N_1425,N_1191);
nand U3675 (N_3675,N_1480,N_1078);
and U3676 (N_3676,N_773,N_870);
and U3677 (N_3677,N_133,N_2493);
nor U3678 (N_3678,N_1840,N_91);
and U3679 (N_3679,N_1282,N_483);
or U3680 (N_3680,N_2330,N_1714);
and U3681 (N_3681,N_1508,N_2032);
and U3682 (N_3682,N_2344,N_1066);
nand U3683 (N_3683,N_193,N_548);
nor U3684 (N_3684,N_1003,N_1446);
or U3685 (N_3685,N_101,N_2167);
nor U3686 (N_3686,N_1161,N_470);
or U3687 (N_3687,N_1646,N_906);
and U3688 (N_3688,N_1892,N_2310);
or U3689 (N_3689,N_864,N_457);
nand U3690 (N_3690,N_544,N_766);
xnor U3691 (N_3691,N_121,N_1864);
or U3692 (N_3692,N_1529,N_2222);
nand U3693 (N_3693,N_2379,N_1873);
xnor U3694 (N_3694,N_347,N_1226);
and U3695 (N_3695,N_1227,N_137);
nand U3696 (N_3696,N_928,N_128);
nand U3697 (N_3697,N_806,N_1384);
and U3698 (N_3698,N_2225,N_1920);
nor U3699 (N_3699,N_1804,N_1082);
nand U3700 (N_3700,N_896,N_6);
nor U3701 (N_3701,N_1143,N_702);
and U3702 (N_3702,N_1310,N_767);
nor U3703 (N_3703,N_1942,N_1466);
and U3704 (N_3704,N_2286,N_612);
nand U3705 (N_3705,N_2236,N_1270);
and U3706 (N_3706,N_143,N_2352);
or U3707 (N_3707,N_2425,N_2394);
or U3708 (N_3708,N_84,N_1455);
nor U3709 (N_3709,N_1912,N_998);
xor U3710 (N_3710,N_961,N_1111);
or U3711 (N_3711,N_1648,N_424);
and U3712 (N_3712,N_2014,N_1071);
or U3713 (N_3713,N_361,N_580);
or U3714 (N_3714,N_232,N_2444);
nor U3715 (N_3715,N_38,N_2359);
nand U3716 (N_3716,N_893,N_2215);
nor U3717 (N_3717,N_1647,N_278);
or U3718 (N_3718,N_1805,N_627);
nand U3719 (N_3719,N_1097,N_1771);
nand U3720 (N_3720,N_1821,N_1015);
nor U3721 (N_3721,N_523,N_1752);
nand U3722 (N_3722,N_915,N_1207);
and U3723 (N_3723,N_1957,N_2304);
or U3724 (N_3724,N_1540,N_993);
and U3725 (N_3725,N_1002,N_463);
nor U3726 (N_3726,N_1198,N_50);
nor U3727 (N_3727,N_838,N_561);
nand U3728 (N_3728,N_688,N_2452);
nor U3729 (N_3729,N_949,N_2268);
nand U3730 (N_3730,N_253,N_1908);
or U3731 (N_3731,N_2022,N_1500);
nand U3732 (N_3732,N_1956,N_600);
or U3733 (N_3733,N_1712,N_1720);
nand U3734 (N_3734,N_25,N_2108);
or U3735 (N_3735,N_234,N_300);
or U3736 (N_3736,N_2272,N_1700);
nor U3737 (N_3737,N_599,N_694);
or U3738 (N_3738,N_246,N_692);
and U3739 (N_3739,N_2291,N_244);
xor U3740 (N_3740,N_31,N_1182);
nor U3741 (N_3741,N_987,N_11);
or U3742 (N_3742,N_1669,N_842);
nand U3743 (N_3743,N_1266,N_2205);
or U3744 (N_3744,N_1285,N_942);
nand U3745 (N_3745,N_1062,N_566);
nor U3746 (N_3746,N_1265,N_24);
nor U3747 (N_3747,N_2001,N_472);
and U3748 (N_3748,N_1011,N_205);
nor U3749 (N_3749,N_2199,N_1914);
nand U3750 (N_3750,N_1600,N_1531);
nor U3751 (N_3751,N_100,N_143);
and U3752 (N_3752,N_2484,N_2461);
nor U3753 (N_3753,N_1384,N_690);
nand U3754 (N_3754,N_295,N_2426);
or U3755 (N_3755,N_984,N_1544);
nor U3756 (N_3756,N_2445,N_2024);
or U3757 (N_3757,N_1367,N_1810);
nor U3758 (N_3758,N_734,N_220);
nor U3759 (N_3759,N_1750,N_2390);
and U3760 (N_3760,N_1501,N_1739);
nand U3761 (N_3761,N_215,N_1567);
nand U3762 (N_3762,N_2314,N_1615);
and U3763 (N_3763,N_2294,N_1103);
or U3764 (N_3764,N_1181,N_858);
xor U3765 (N_3765,N_845,N_618);
nand U3766 (N_3766,N_271,N_1876);
or U3767 (N_3767,N_418,N_1790);
or U3768 (N_3768,N_840,N_1022);
nand U3769 (N_3769,N_897,N_813);
nor U3770 (N_3770,N_2331,N_1111);
nand U3771 (N_3771,N_492,N_2372);
nor U3772 (N_3772,N_975,N_1394);
nand U3773 (N_3773,N_1728,N_2498);
xnor U3774 (N_3774,N_233,N_2124);
xnor U3775 (N_3775,N_1986,N_1571);
xnor U3776 (N_3776,N_1847,N_975);
or U3777 (N_3777,N_1336,N_1460);
nor U3778 (N_3778,N_2269,N_811);
nor U3779 (N_3779,N_1858,N_2201);
and U3780 (N_3780,N_1473,N_947);
or U3781 (N_3781,N_2044,N_1511);
or U3782 (N_3782,N_412,N_1985);
or U3783 (N_3783,N_200,N_570);
nor U3784 (N_3784,N_2096,N_1396);
xor U3785 (N_3785,N_348,N_1081);
or U3786 (N_3786,N_778,N_1371);
nand U3787 (N_3787,N_246,N_90);
or U3788 (N_3788,N_876,N_162);
nand U3789 (N_3789,N_2370,N_1776);
nor U3790 (N_3790,N_1866,N_2080);
or U3791 (N_3791,N_201,N_1501);
or U3792 (N_3792,N_1606,N_1177);
or U3793 (N_3793,N_815,N_1767);
or U3794 (N_3794,N_46,N_920);
nand U3795 (N_3795,N_2149,N_1520);
nor U3796 (N_3796,N_507,N_2481);
nand U3797 (N_3797,N_852,N_820);
nand U3798 (N_3798,N_2262,N_84);
or U3799 (N_3799,N_1277,N_702);
and U3800 (N_3800,N_946,N_596);
nand U3801 (N_3801,N_1111,N_1579);
or U3802 (N_3802,N_1647,N_2426);
nor U3803 (N_3803,N_898,N_345);
or U3804 (N_3804,N_1080,N_981);
or U3805 (N_3805,N_301,N_2268);
and U3806 (N_3806,N_2468,N_2405);
nor U3807 (N_3807,N_40,N_1928);
nand U3808 (N_3808,N_1223,N_2006);
or U3809 (N_3809,N_1179,N_200);
nand U3810 (N_3810,N_1444,N_884);
or U3811 (N_3811,N_2088,N_247);
or U3812 (N_3812,N_305,N_280);
nor U3813 (N_3813,N_1049,N_1007);
and U3814 (N_3814,N_2155,N_260);
nor U3815 (N_3815,N_2004,N_2046);
and U3816 (N_3816,N_722,N_2140);
and U3817 (N_3817,N_258,N_849);
nor U3818 (N_3818,N_2336,N_1695);
and U3819 (N_3819,N_1007,N_1574);
nand U3820 (N_3820,N_819,N_2142);
xor U3821 (N_3821,N_1320,N_180);
nor U3822 (N_3822,N_1404,N_1253);
nor U3823 (N_3823,N_2204,N_1362);
xor U3824 (N_3824,N_1950,N_2204);
or U3825 (N_3825,N_2304,N_134);
nand U3826 (N_3826,N_947,N_1903);
and U3827 (N_3827,N_2354,N_205);
nand U3828 (N_3828,N_2286,N_1693);
nand U3829 (N_3829,N_427,N_98);
nor U3830 (N_3830,N_735,N_1333);
nor U3831 (N_3831,N_2207,N_1014);
or U3832 (N_3832,N_2453,N_1512);
or U3833 (N_3833,N_947,N_431);
and U3834 (N_3834,N_1438,N_1825);
or U3835 (N_3835,N_2301,N_426);
or U3836 (N_3836,N_1873,N_547);
nor U3837 (N_3837,N_1517,N_1847);
nand U3838 (N_3838,N_502,N_2335);
nor U3839 (N_3839,N_1954,N_728);
nand U3840 (N_3840,N_1005,N_396);
or U3841 (N_3841,N_1531,N_1029);
and U3842 (N_3842,N_255,N_591);
xnor U3843 (N_3843,N_421,N_1749);
nor U3844 (N_3844,N_490,N_1074);
and U3845 (N_3845,N_546,N_1405);
nand U3846 (N_3846,N_1459,N_2471);
and U3847 (N_3847,N_547,N_1942);
and U3848 (N_3848,N_2113,N_1951);
and U3849 (N_3849,N_1010,N_1503);
and U3850 (N_3850,N_779,N_2085);
and U3851 (N_3851,N_515,N_542);
or U3852 (N_3852,N_799,N_425);
nand U3853 (N_3853,N_1377,N_2477);
nor U3854 (N_3854,N_1400,N_518);
or U3855 (N_3855,N_1757,N_255);
or U3856 (N_3856,N_716,N_213);
nand U3857 (N_3857,N_1462,N_2153);
and U3858 (N_3858,N_1398,N_95);
and U3859 (N_3859,N_1773,N_646);
or U3860 (N_3860,N_1364,N_2421);
nor U3861 (N_3861,N_1660,N_1369);
and U3862 (N_3862,N_449,N_1769);
nand U3863 (N_3863,N_2435,N_2168);
nor U3864 (N_3864,N_2406,N_1790);
and U3865 (N_3865,N_1940,N_1217);
or U3866 (N_3866,N_2398,N_1909);
nor U3867 (N_3867,N_2328,N_2300);
and U3868 (N_3868,N_920,N_791);
or U3869 (N_3869,N_661,N_1175);
nand U3870 (N_3870,N_1356,N_1650);
or U3871 (N_3871,N_199,N_618);
and U3872 (N_3872,N_733,N_1362);
or U3873 (N_3873,N_2026,N_150);
and U3874 (N_3874,N_2040,N_608);
or U3875 (N_3875,N_982,N_866);
nor U3876 (N_3876,N_632,N_2082);
or U3877 (N_3877,N_1258,N_277);
xnor U3878 (N_3878,N_365,N_1387);
nand U3879 (N_3879,N_774,N_2441);
nor U3880 (N_3880,N_669,N_476);
nand U3881 (N_3881,N_555,N_936);
nor U3882 (N_3882,N_799,N_1161);
nand U3883 (N_3883,N_282,N_2023);
nand U3884 (N_3884,N_428,N_1208);
nor U3885 (N_3885,N_1474,N_2465);
and U3886 (N_3886,N_944,N_2078);
nand U3887 (N_3887,N_1682,N_292);
and U3888 (N_3888,N_429,N_2022);
nand U3889 (N_3889,N_132,N_2487);
nand U3890 (N_3890,N_2120,N_728);
nand U3891 (N_3891,N_121,N_2140);
nor U3892 (N_3892,N_2030,N_1154);
or U3893 (N_3893,N_1180,N_576);
and U3894 (N_3894,N_311,N_530);
nand U3895 (N_3895,N_584,N_610);
nor U3896 (N_3896,N_1156,N_1852);
and U3897 (N_3897,N_1726,N_1319);
nand U3898 (N_3898,N_302,N_651);
nand U3899 (N_3899,N_1689,N_821);
xnor U3900 (N_3900,N_436,N_2096);
and U3901 (N_3901,N_1066,N_1843);
nand U3902 (N_3902,N_2354,N_2431);
or U3903 (N_3903,N_1236,N_1604);
and U3904 (N_3904,N_1678,N_1600);
nand U3905 (N_3905,N_1579,N_1480);
nand U3906 (N_3906,N_1429,N_1478);
nand U3907 (N_3907,N_50,N_1967);
nand U3908 (N_3908,N_912,N_53);
xnor U3909 (N_3909,N_1938,N_705);
and U3910 (N_3910,N_1554,N_333);
or U3911 (N_3911,N_1977,N_1627);
and U3912 (N_3912,N_2262,N_1456);
nand U3913 (N_3913,N_825,N_1652);
and U3914 (N_3914,N_1413,N_1833);
and U3915 (N_3915,N_164,N_2034);
nor U3916 (N_3916,N_1247,N_1152);
nor U3917 (N_3917,N_1981,N_793);
nand U3918 (N_3918,N_2175,N_446);
and U3919 (N_3919,N_1985,N_911);
and U3920 (N_3920,N_866,N_417);
xor U3921 (N_3921,N_2229,N_1177);
and U3922 (N_3922,N_2100,N_2494);
or U3923 (N_3923,N_968,N_930);
nor U3924 (N_3924,N_1986,N_2219);
nand U3925 (N_3925,N_2432,N_1125);
nand U3926 (N_3926,N_384,N_1313);
and U3927 (N_3927,N_1056,N_1978);
xnor U3928 (N_3928,N_2262,N_1905);
nor U3929 (N_3929,N_1964,N_80);
and U3930 (N_3930,N_2088,N_1506);
and U3931 (N_3931,N_974,N_532);
nor U3932 (N_3932,N_2284,N_1015);
nor U3933 (N_3933,N_517,N_375);
nand U3934 (N_3934,N_467,N_207);
nor U3935 (N_3935,N_1715,N_1476);
nor U3936 (N_3936,N_329,N_653);
nand U3937 (N_3937,N_2117,N_11);
nor U3938 (N_3938,N_898,N_1556);
and U3939 (N_3939,N_815,N_1649);
or U3940 (N_3940,N_301,N_1752);
nor U3941 (N_3941,N_2133,N_645);
nand U3942 (N_3942,N_2080,N_349);
and U3943 (N_3943,N_649,N_377);
and U3944 (N_3944,N_1551,N_1900);
xnor U3945 (N_3945,N_487,N_128);
nand U3946 (N_3946,N_2499,N_391);
nor U3947 (N_3947,N_1995,N_2073);
nand U3948 (N_3948,N_494,N_168);
or U3949 (N_3949,N_1987,N_1637);
nor U3950 (N_3950,N_1373,N_1507);
nand U3951 (N_3951,N_1845,N_1438);
or U3952 (N_3952,N_864,N_98);
and U3953 (N_3953,N_34,N_398);
or U3954 (N_3954,N_46,N_1166);
nand U3955 (N_3955,N_1580,N_2330);
or U3956 (N_3956,N_981,N_1904);
nand U3957 (N_3957,N_847,N_264);
or U3958 (N_3958,N_712,N_664);
nor U3959 (N_3959,N_5,N_2178);
nand U3960 (N_3960,N_826,N_1178);
and U3961 (N_3961,N_138,N_1606);
or U3962 (N_3962,N_811,N_2451);
xor U3963 (N_3963,N_436,N_1929);
or U3964 (N_3964,N_1574,N_625);
nor U3965 (N_3965,N_1126,N_1517);
or U3966 (N_3966,N_363,N_1741);
or U3967 (N_3967,N_873,N_1311);
nor U3968 (N_3968,N_1085,N_1881);
and U3969 (N_3969,N_1386,N_1116);
nor U3970 (N_3970,N_391,N_212);
or U3971 (N_3971,N_1188,N_1710);
nand U3972 (N_3972,N_412,N_2423);
nand U3973 (N_3973,N_800,N_750);
or U3974 (N_3974,N_1002,N_1001);
or U3975 (N_3975,N_2460,N_2075);
and U3976 (N_3976,N_1074,N_864);
or U3977 (N_3977,N_1040,N_2134);
or U3978 (N_3978,N_787,N_630);
nand U3979 (N_3979,N_2238,N_1329);
or U3980 (N_3980,N_2095,N_1756);
nor U3981 (N_3981,N_1431,N_1621);
and U3982 (N_3982,N_928,N_152);
and U3983 (N_3983,N_686,N_1180);
nor U3984 (N_3984,N_1340,N_2115);
nand U3985 (N_3985,N_1849,N_1422);
and U3986 (N_3986,N_55,N_211);
or U3987 (N_3987,N_322,N_2053);
and U3988 (N_3988,N_28,N_75);
and U3989 (N_3989,N_1839,N_1144);
nor U3990 (N_3990,N_2037,N_164);
nand U3991 (N_3991,N_2058,N_2096);
nor U3992 (N_3992,N_2326,N_769);
nor U3993 (N_3993,N_1653,N_1321);
xor U3994 (N_3994,N_184,N_750);
and U3995 (N_3995,N_1325,N_1249);
or U3996 (N_3996,N_2229,N_1075);
or U3997 (N_3997,N_1019,N_349);
or U3998 (N_3998,N_740,N_1084);
and U3999 (N_3999,N_2305,N_1070);
nand U4000 (N_4000,N_1374,N_99);
nor U4001 (N_4001,N_23,N_1954);
nand U4002 (N_4002,N_1559,N_2001);
or U4003 (N_4003,N_165,N_1199);
nand U4004 (N_4004,N_354,N_34);
nor U4005 (N_4005,N_1348,N_1876);
and U4006 (N_4006,N_1676,N_1666);
or U4007 (N_4007,N_1937,N_1347);
nor U4008 (N_4008,N_2441,N_657);
or U4009 (N_4009,N_2460,N_1166);
nand U4010 (N_4010,N_292,N_404);
nor U4011 (N_4011,N_2301,N_2423);
nor U4012 (N_4012,N_2295,N_1777);
nand U4013 (N_4013,N_753,N_2376);
nand U4014 (N_4014,N_692,N_2457);
or U4015 (N_4015,N_583,N_548);
nor U4016 (N_4016,N_1597,N_1486);
nand U4017 (N_4017,N_138,N_1494);
or U4018 (N_4018,N_604,N_106);
or U4019 (N_4019,N_430,N_675);
or U4020 (N_4020,N_31,N_1850);
and U4021 (N_4021,N_998,N_1060);
or U4022 (N_4022,N_2114,N_1826);
and U4023 (N_4023,N_1152,N_861);
or U4024 (N_4024,N_309,N_312);
or U4025 (N_4025,N_94,N_1043);
xnor U4026 (N_4026,N_1575,N_1089);
or U4027 (N_4027,N_298,N_186);
nor U4028 (N_4028,N_2176,N_2187);
nor U4029 (N_4029,N_714,N_1284);
nor U4030 (N_4030,N_117,N_601);
nand U4031 (N_4031,N_726,N_1);
nor U4032 (N_4032,N_720,N_1376);
nor U4033 (N_4033,N_60,N_1116);
and U4034 (N_4034,N_2054,N_372);
and U4035 (N_4035,N_869,N_326);
and U4036 (N_4036,N_2248,N_2403);
nand U4037 (N_4037,N_577,N_87);
or U4038 (N_4038,N_453,N_472);
nor U4039 (N_4039,N_1071,N_776);
and U4040 (N_4040,N_734,N_2079);
or U4041 (N_4041,N_904,N_2031);
nand U4042 (N_4042,N_1834,N_588);
and U4043 (N_4043,N_2482,N_1377);
nor U4044 (N_4044,N_276,N_2404);
and U4045 (N_4045,N_916,N_734);
nor U4046 (N_4046,N_1864,N_1686);
nor U4047 (N_4047,N_1134,N_2071);
or U4048 (N_4048,N_1382,N_1407);
or U4049 (N_4049,N_2003,N_180);
nand U4050 (N_4050,N_2273,N_2439);
or U4051 (N_4051,N_606,N_904);
nand U4052 (N_4052,N_1717,N_1458);
and U4053 (N_4053,N_2184,N_926);
nand U4054 (N_4054,N_576,N_1048);
nor U4055 (N_4055,N_970,N_483);
or U4056 (N_4056,N_181,N_2010);
nand U4057 (N_4057,N_758,N_2302);
nor U4058 (N_4058,N_1366,N_879);
or U4059 (N_4059,N_689,N_1373);
or U4060 (N_4060,N_965,N_2386);
or U4061 (N_4061,N_34,N_1608);
or U4062 (N_4062,N_1644,N_536);
nor U4063 (N_4063,N_1086,N_141);
and U4064 (N_4064,N_1029,N_16);
xnor U4065 (N_4065,N_2410,N_1883);
or U4066 (N_4066,N_256,N_1029);
xnor U4067 (N_4067,N_820,N_588);
nand U4068 (N_4068,N_198,N_1234);
nand U4069 (N_4069,N_1681,N_1627);
and U4070 (N_4070,N_2282,N_2352);
nor U4071 (N_4071,N_452,N_132);
or U4072 (N_4072,N_2188,N_2029);
nand U4073 (N_4073,N_2318,N_2241);
nand U4074 (N_4074,N_2362,N_861);
nand U4075 (N_4075,N_2082,N_1360);
nand U4076 (N_4076,N_396,N_1524);
and U4077 (N_4077,N_1349,N_1960);
nand U4078 (N_4078,N_376,N_24);
nor U4079 (N_4079,N_19,N_1224);
nand U4080 (N_4080,N_968,N_1662);
nand U4081 (N_4081,N_1661,N_2030);
and U4082 (N_4082,N_1203,N_2343);
and U4083 (N_4083,N_252,N_2034);
or U4084 (N_4084,N_610,N_1174);
or U4085 (N_4085,N_111,N_1582);
nand U4086 (N_4086,N_1998,N_238);
nor U4087 (N_4087,N_187,N_1003);
nor U4088 (N_4088,N_371,N_1979);
nand U4089 (N_4089,N_1056,N_1725);
nor U4090 (N_4090,N_2286,N_653);
or U4091 (N_4091,N_446,N_1718);
nand U4092 (N_4092,N_383,N_2436);
nor U4093 (N_4093,N_1390,N_2355);
nor U4094 (N_4094,N_2456,N_505);
and U4095 (N_4095,N_1649,N_535);
nor U4096 (N_4096,N_1772,N_2236);
nor U4097 (N_4097,N_2178,N_370);
nor U4098 (N_4098,N_2388,N_2421);
nand U4099 (N_4099,N_2336,N_735);
and U4100 (N_4100,N_1329,N_1814);
nor U4101 (N_4101,N_757,N_863);
and U4102 (N_4102,N_1214,N_1420);
or U4103 (N_4103,N_1094,N_1256);
or U4104 (N_4104,N_1173,N_834);
and U4105 (N_4105,N_649,N_2428);
nand U4106 (N_4106,N_270,N_1886);
and U4107 (N_4107,N_1265,N_1184);
nor U4108 (N_4108,N_92,N_1521);
or U4109 (N_4109,N_462,N_276);
or U4110 (N_4110,N_1411,N_1872);
and U4111 (N_4111,N_639,N_911);
xor U4112 (N_4112,N_2342,N_581);
or U4113 (N_4113,N_2327,N_716);
or U4114 (N_4114,N_552,N_2311);
nand U4115 (N_4115,N_1736,N_1197);
nor U4116 (N_4116,N_1450,N_1029);
nand U4117 (N_4117,N_600,N_1579);
and U4118 (N_4118,N_1429,N_19);
or U4119 (N_4119,N_1680,N_1597);
or U4120 (N_4120,N_730,N_339);
and U4121 (N_4121,N_729,N_520);
or U4122 (N_4122,N_1153,N_1364);
or U4123 (N_4123,N_709,N_1617);
nand U4124 (N_4124,N_1250,N_2304);
and U4125 (N_4125,N_1668,N_1228);
and U4126 (N_4126,N_868,N_257);
nor U4127 (N_4127,N_1361,N_2436);
and U4128 (N_4128,N_840,N_1027);
or U4129 (N_4129,N_839,N_722);
and U4130 (N_4130,N_217,N_746);
nor U4131 (N_4131,N_1128,N_2305);
or U4132 (N_4132,N_1416,N_2075);
or U4133 (N_4133,N_1023,N_1794);
and U4134 (N_4134,N_2020,N_82);
xnor U4135 (N_4135,N_315,N_2382);
and U4136 (N_4136,N_1557,N_1284);
and U4137 (N_4137,N_622,N_2024);
nor U4138 (N_4138,N_980,N_160);
or U4139 (N_4139,N_89,N_909);
or U4140 (N_4140,N_49,N_2073);
or U4141 (N_4141,N_351,N_2182);
nor U4142 (N_4142,N_1816,N_1683);
nand U4143 (N_4143,N_1786,N_1832);
or U4144 (N_4144,N_221,N_303);
and U4145 (N_4145,N_519,N_1018);
nand U4146 (N_4146,N_1094,N_1160);
nor U4147 (N_4147,N_2454,N_1771);
or U4148 (N_4148,N_1188,N_2188);
nor U4149 (N_4149,N_1121,N_1789);
and U4150 (N_4150,N_1766,N_1267);
nand U4151 (N_4151,N_881,N_887);
nor U4152 (N_4152,N_580,N_2117);
or U4153 (N_4153,N_1862,N_1659);
nor U4154 (N_4154,N_422,N_1429);
nand U4155 (N_4155,N_325,N_1185);
nor U4156 (N_4156,N_606,N_2164);
and U4157 (N_4157,N_542,N_866);
nor U4158 (N_4158,N_1318,N_532);
nand U4159 (N_4159,N_2152,N_2438);
nor U4160 (N_4160,N_878,N_1569);
nor U4161 (N_4161,N_2335,N_421);
and U4162 (N_4162,N_599,N_812);
or U4163 (N_4163,N_2396,N_1981);
or U4164 (N_4164,N_2100,N_2160);
or U4165 (N_4165,N_923,N_403);
and U4166 (N_4166,N_1709,N_1841);
nor U4167 (N_4167,N_1349,N_823);
nand U4168 (N_4168,N_2303,N_2318);
and U4169 (N_4169,N_1148,N_968);
or U4170 (N_4170,N_2080,N_980);
and U4171 (N_4171,N_2152,N_358);
and U4172 (N_4172,N_1064,N_1757);
nand U4173 (N_4173,N_1598,N_1685);
or U4174 (N_4174,N_992,N_1391);
or U4175 (N_4175,N_570,N_918);
nor U4176 (N_4176,N_1279,N_2333);
or U4177 (N_4177,N_2440,N_1965);
nor U4178 (N_4178,N_1958,N_2192);
and U4179 (N_4179,N_2131,N_1227);
or U4180 (N_4180,N_460,N_1097);
or U4181 (N_4181,N_1951,N_470);
and U4182 (N_4182,N_1106,N_1799);
and U4183 (N_4183,N_1386,N_1623);
and U4184 (N_4184,N_2389,N_2237);
nand U4185 (N_4185,N_334,N_591);
and U4186 (N_4186,N_2348,N_1107);
or U4187 (N_4187,N_1032,N_1175);
nor U4188 (N_4188,N_1014,N_1684);
and U4189 (N_4189,N_2118,N_9);
or U4190 (N_4190,N_2188,N_1393);
nor U4191 (N_4191,N_1734,N_614);
and U4192 (N_4192,N_751,N_405);
nor U4193 (N_4193,N_1194,N_1516);
and U4194 (N_4194,N_2181,N_601);
and U4195 (N_4195,N_1219,N_829);
nand U4196 (N_4196,N_2150,N_755);
and U4197 (N_4197,N_2035,N_250);
and U4198 (N_4198,N_938,N_594);
and U4199 (N_4199,N_2423,N_1327);
or U4200 (N_4200,N_24,N_2096);
and U4201 (N_4201,N_626,N_798);
or U4202 (N_4202,N_347,N_302);
xnor U4203 (N_4203,N_379,N_1529);
nor U4204 (N_4204,N_1331,N_1594);
nand U4205 (N_4205,N_1861,N_1166);
or U4206 (N_4206,N_411,N_1218);
nand U4207 (N_4207,N_1377,N_1529);
nand U4208 (N_4208,N_2267,N_467);
or U4209 (N_4209,N_1556,N_2175);
nor U4210 (N_4210,N_2261,N_1112);
and U4211 (N_4211,N_417,N_203);
nand U4212 (N_4212,N_802,N_2004);
and U4213 (N_4213,N_707,N_2171);
and U4214 (N_4214,N_121,N_2489);
or U4215 (N_4215,N_369,N_457);
nor U4216 (N_4216,N_2226,N_1179);
or U4217 (N_4217,N_1340,N_2156);
and U4218 (N_4218,N_516,N_1372);
or U4219 (N_4219,N_1954,N_1228);
and U4220 (N_4220,N_2049,N_1112);
nand U4221 (N_4221,N_1416,N_1355);
nand U4222 (N_4222,N_1327,N_211);
nor U4223 (N_4223,N_2196,N_2017);
nor U4224 (N_4224,N_841,N_1676);
xnor U4225 (N_4225,N_1956,N_553);
or U4226 (N_4226,N_1330,N_1622);
nand U4227 (N_4227,N_1818,N_1944);
and U4228 (N_4228,N_567,N_1973);
and U4229 (N_4229,N_1936,N_2490);
nand U4230 (N_4230,N_2407,N_342);
and U4231 (N_4231,N_278,N_583);
and U4232 (N_4232,N_2368,N_545);
nor U4233 (N_4233,N_2386,N_1495);
nor U4234 (N_4234,N_1280,N_1405);
nand U4235 (N_4235,N_23,N_1076);
nand U4236 (N_4236,N_363,N_387);
nand U4237 (N_4237,N_1057,N_1946);
nor U4238 (N_4238,N_1350,N_1248);
nand U4239 (N_4239,N_1291,N_569);
or U4240 (N_4240,N_2092,N_66);
nor U4241 (N_4241,N_1386,N_1023);
or U4242 (N_4242,N_1439,N_1689);
nor U4243 (N_4243,N_704,N_792);
or U4244 (N_4244,N_1341,N_1820);
or U4245 (N_4245,N_2031,N_589);
and U4246 (N_4246,N_1706,N_1970);
nand U4247 (N_4247,N_1294,N_2440);
or U4248 (N_4248,N_692,N_56);
and U4249 (N_4249,N_2017,N_1608);
or U4250 (N_4250,N_1901,N_2263);
and U4251 (N_4251,N_1107,N_896);
nor U4252 (N_4252,N_1586,N_433);
xor U4253 (N_4253,N_596,N_789);
or U4254 (N_4254,N_513,N_1412);
and U4255 (N_4255,N_2082,N_675);
nor U4256 (N_4256,N_2155,N_1072);
and U4257 (N_4257,N_355,N_764);
and U4258 (N_4258,N_2082,N_613);
nor U4259 (N_4259,N_1101,N_2240);
and U4260 (N_4260,N_167,N_2376);
or U4261 (N_4261,N_1358,N_2172);
or U4262 (N_4262,N_888,N_2360);
and U4263 (N_4263,N_404,N_1454);
or U4264 (N_4264,N_763,N_2316);
nor U4265 (N_4265,N_196,N_373);
and U4266 (N_4266,N_1316,N_1284);
and U4267 (N_4267,N_2302,N_1530);
or U4268 (N_4268,N_78,N_1929);
and U4269 (N_4269,N_2169,N_2259);
nand U4270 (N_4270,N_2269,N_1218);
nand U4271 (N_4271,N_373,N_1998);
nand U4272 (N_4272,N_1680,N_556);
nand U4273 (N_4273,N_1880,N_2320);
nor U4274 (N_4274,N_602,N_1101);
or U4275 (N_4275,N_208,N_443);
and U4276 (N_4276,N_58,N_143);
and U4277 (N_4277,N_328,N_646);
and U4278 (N_4278,N_231,N_631);
nor U4279 (N_4279,N_1435,N_1252);
nand U4280 (N_4280,N_746,N_686);
and U4281 (N_4281,N_1539,N_972);
nor U4282 (N_4282,N_537,N_2029);
and U4283 (N_4283,N_1485,N_2049);
or U4284 (N_4284,N_622,N_2197);
nand U4285 (N_4285,N_1774,N_1284);
or U4286 (N_4286,N_796,N_442);
nand U4287 (N_4287,N_2177,N_2196);
or U4288 (N_4288,N_799,N_641);
or U4289 (N_4289,N_1069,N_1797);
or U4290 (N_4290,N_620,N_1824);
or U4291 (N_4291,N_847,N_1686);
nor U4292 (N_4292,N_339,N_162);
and U4293 (N_4293,N_316,N_123);
nand U4294 (N_4294,N_10,N_2055);
nand U4295 (N_4295,N_1661,N_1358);
nor U4296 (N_4296,N_462,N_562);
nand U4297 (N_4297,N_1810,N_2230);
nand U4298 (N_4298,N_2419,N_24);
nand U4299 (N_4299,N_2209,N_1446);
and U4300 (N_4300,N_1910,N_1992);
nand U4301 (N_4301,N_1102,N_970);
or U4302 (N_4302,N_1209,N_2459);
or U4303 (N_4303,N_2151,N_353);
nand U4304 (N_4304,N_1665,N_2444);
and U4305 (N_4305,N_2021,N_50);
nand U4306 (N_4306,N_1126,N_1442);
nand U4307 (N_4307,N_425,N_50);
or U4308 (N_4308,N_1678,N_571);
and U4309 (N_4309,N_984,N_723);
nor U4310 (N_4310,N_1683,N_470);
or U4311 (N_4311,N_460,N_664);
nand U4312 (N_4312,N_1735,N_1291);
nor U4313 (N_4313,N_1280,N_68);
nor U4314 (N_4314,N_2154,N_47);
nor U4315 (N_4315,N_1046,N_2219);
nor U4316 (N_4316,N_2484,N_2011);
or U4317 (N_4317,N_227,N_967);
and U4318 (N_4318,N_290,N_1603);
nor U4319 (N_4319,N_527,N_705);
nor U4320 (N_4320,N_654,N_1684);
or U4321 (N_4321,N_2451,N_2416);
or U4322 (N_4322,N_1210,N_2166);
xor U4323 (N_4323,N_807,N_2326);
and U4324 (N_4324,N_1064,N_1218);
or U4325 (N_4325,N_1215,N_2245);
and U4326 (N_4326,N_1041,N_2403);
or U4327 (N_4327,N_2376,N_239);
nand U4328 (N_4328,N_1223,N_1278);
nand U4329 (N_4329,N_2440,N_1826);
or U4330 (N_4330,N_1533,N_562);
and U4331 (N_4331,N_151,N_1612);
and U4332 (N_4332,N_2067,N_1825);
nand U4333 (N_4333,N_1462,N_587);
nor U4334 (N_4334,N_468,N_274);
or U4335 (N_4335,N_2302,N_1823);
or U4336 (N_4336,N_795,N_1094);
and U4337 (N_4337,N_1870,N_1097);
or U4338 (N_4338,N_1555,N_140);
nand U4339 (N_4339,N_2325,N_1053);
or U4340 (N_4340,N_1142,N_502);
nand U4341 (N_4341,N_1246,N_1336);
or U4342 (N_4342,N_2360,N_2270);
nand U4343 (N_4343,N_1567,N_799);
nor U4344 (N_4344,N_549,N_2258);
nor U4345 (N_4345,N_1371,N_2281);
and U4346 (N_4346,N_2246,N_1368);
and U4347 (N_4347,N_1717,N_2328);
or U4348 (N_4348,N_1728,N_1227);
nand U4349 (N_4349,N_1780,N_1759);
nand U4350 (N_4350,N_565,N_2410);
and U4351 (N_4351,N_769,N_739);
nor U4352 (N_4352,N_111,N_572);
or U4353 (N_4353,N_161,N_843);
and U4354 (N_4354,N_36,N_2287);
or U4355 (N_4355,N_1319,N_1636);
nand U4356 (N_4356,N_785,N_1650);
nand U4357 (N_4357,N_1668,N_2150);
or U4358 (N_4358,N_1936,N_1201);
and U4359 (N_4359,N_1047,N_1734);
nor U4360 (N_4360,N_889,N_1261);
and U4361 (N_4361,N_2233,N_1482);
or U4362 (N_4362,N_498,N_678);
xnor U4363 (N_4363,N_1250,N_123);
or U4364 (N_4364,N_325,N_2125);
and U4365 (N_4365,N_1565,N_621);
nor U4366 (N_4366,N_1328,N_2071);
nor U4367 (N_4367,N_2301,N_153);
and U4368 (N_4368,N_943,N_34);
or U4369 (N_4369,N_1403,N_1412);
and U4370 (N_4370,N_223,N_384);
nor U4371 (N_4371,N_127,N_1875);
or U4372 (N_4372,N_1957,N_2478);
xor U4373 (N_4373,N_2114,N_1740);
or U4374 (N_4374,N_1687,N_1285);
or U4375 (N_4375,N_95,N_679);
nor U4376 (N_4376,N_1899,N_1336);
nor U4377 (N_4377,N_1980,N_1323);
nor U4378 (N_4378,N_510,N_1581);
nand U4379 (N_4379,N_967,N_1947);
nand U4380 (N_4380,N_908,N_2010);
nor U4381 (N_4381,N_1878,N_1932);
nor U4382 (N_4382,N_1465,N_751);
nor U4383 (N_4383,N_814,N_1362);
and U4384 (N_4384,N_449,N_329);
nor U4385 (N_4385,N_750,N_1217);
and U4386 (N_4386,N_798,N_2334);
or U4387 (N_4387,N_425,N_924);
xnor U4388 (N_4388,N_551,N_2153);
and U4389 (N_4389,N_1795,N_2214);
and U4390 (N_4390,N_566,N_1910);
nor U4391 (N_4391,N_1533,N_1540);
and U4392 (N_4392,N_329,N_1992);
and U4393 (N_4393,N_1555,N_1261);
nor U4394 (N_4394,N_1815,N_448);
or U4395 (N_4395,N_1223,N_318);
or U4396 (N_4396,N_1769,N_1345);
nor U4397 (N_4397,N_1030,N_485);
and U4398 (N_4398,N_667,N_1202);
and U4399 (N_4399,N_240,N_2040);
nand U4400 (N_4400,N_2072,N_1288);
or U4401 (N_4401,N_30,N_911);
nand U4402 (N_4402,N_326,N_1);
or U4403 (N_4403,N_1917,N_164);
or U4404 (N_4404,N_232,N_1813);
and U4405 (N_4405,N_871,N_1553);
or U4406 (N_4406,N_512,N_1996);
nor U4407 (N_4407,N_656,N_2142);
nand U4408 (N_4408,N_2409,N_2013);
nand U4409 (N_4409,N_553,N_299);
and U4410 (N_4410,N_1551,N_2463);
xor U4411 (N_4411,N_2429,N_1648);
nor U4412 (N_4412,N_1903,N_1694);
nand U4413 (N_4413,N_1804,N_6);
or U4414 (N_4414,N_473,N_966);
and U4415 (N_4415,N_1100,N_1515);
and U4416 (N_4416,N_2114,N_1831);
nand U4417 (N_4417,N_1564,N_2285);
or U4418 (N_4418,N_1175,N_227);
or U4419 (N_4419,N_1270,N_110);
and U4420 (N_4420,N_174,N_1894);
nand U4421 (N_4421,N_674,N_2218);
nand U4422 (N_4422,N_1181,N_1532);
or U4423 (N_4423,N_1173,N_1910);
or U4424 (N_4424,N_1460,N_1251);
or U4425 (N_4425,N_1976,N_2383);
and U4426 (N_4426,N_1153,N_1048);
or U4427 (N_4427,N_1409,N_961);
nor U4428 (N_4428,N_2253,N_462);
or U4429 (N_4429,N_1410,N_2055);
or U4430 (N_4430,N_1035,N_2359);
or U4431 (N_4431,N_974,N_2272);
nor U4432 (N_4432,N_1365,N_1294);
or U4433 (N_4433,N_131,N_657);
nor U4434 (N_4434,N_2461,N_1550);
and U4435 (N_4435,N_31,N_484);
nor U4436 (N_4436,N_2062,N_1033);
and U4437 (N_4437,N_1070,N_1581);
and U4438 (N_4438,N_1725,N_799);
nand U4439 (N_4439,N_1001,N_252);
nor U4440 (N_4440,N_447,N_1317);
or U4441 (N_4441,N_2063,N_203);
nor U4442 (N_4442,N_946,N_2137);
nor U4443 (N_4443,N_215,N_2318);
and U4444 (N_4444,N_163,N_1725);
nand U4445 (N_4445,N_1659,N_906);
nand U4446 (N_4446,N_1272,N_1452);
nor U4447 (N_4447,N_2061,N_2046);
or U4448 (N_4448,N_1794,N_1521);
nor U4449 (N_4449,N_2490,N_28);
nor U4450 (N_4450,N_663,N_2062);
nor U4451 (N_4451,N_555,N_44);
nand U4452 (N_4452,N_1612,N_427);
or U4453 (N_4453,N_904,N_517);
nor U4454 (N_4454,N_571,N_2314);
or U4455 (N_4455,N_1010,N_1355);
and U4456 (N_4456,N_713,N_884);
nor U4457 (N_4457,N_1967,N_1585);
nand U4458 (N_4458,N_1260,N_414);
nand U4459 (N_4459,N_1485,N_308);
nand U4460 (N_4460,N_1567,N_873);
or U4461 (N_4461,N_1492,N_2415);
nor U4462 (N_4462,N_1649,N_393);
nor U4463 (N_4463,N_1149,N_984);
or U4464 (N_4464,N_717,N_623);
nand U4465 (N_4465,N_1927,N_1170);
nand U4466 (N_4466,N_831,N_845);
or U4467 (N_4467,N_1827,N_2066);
or U4468 (N_4468,N_2421,N_1996);
or U4469 (N_4469,N_1980,N_333);
nand U4470 (N_4470,N_2130,N_2125);
nor U4471 (N_4471,N_1891,N_1341);
and U4472 (N_4472,N_2323,N_1063);
nand U4473 (N_4473,N_2367,N_2251);
nand U4474 (N_4474,N_998,N_828);
and U4475 (N_4475,N_2462,N_2396);
or U4476 (N_4476,N_1678,N_464);
or U4477 (N_4477,N_2110,N_2152);
or U4478 (N_4478,N_1477,N_1886);
nand U4479 (N_4479,N_82,N_2359);
and U4480 (N_4480,N_1784,N_1933);
and U4481 (N_4481,N_534,N_2073);
or U4482 (N_4482,N_307,N_2126);
nor U4483 (N_4483,N_2498,N_373);
nor U4484 (N_4484,N_1022,N_962);
nand U4485 (N_4485,N_1609,N_1344);
nand U4486 (N_4486,N_1769,N_2102);
or U4487 (N_4487,N_1384,N_188);
and U4488 (N_4488,N_1327,N_2363);
xor U4489 (N_4489,N_1934,N_2499);
and U4490 (N_4490,N_352,N_423);
or U4491 (N_4491,N_280,N_2113);
and U4492 (N_4492,N_1974,N_1021);
or U4493 (N_4493,N_308,N_204);
nor U4494 (N_4494,N_988,N_2169);
nor U4495 (N_4495,N_1726,N_1235);
xor U4496 (N_4496,N_1026,N_547);
nor U4497 (N_4497,N_828,N_2087);
nor U4498 (N_4498,N_1197,N_817);
xor U4499 (N_4499,N_1008,N_108);
and U4500 (N_4500,N_1370,N_1435);
and U4501 (N_4501,N_1283,N_46);
or U4502 (N_4502,N_401,N_975);
nand U4503 (N_4503,N_638,N_599);
xor U4504 (N_4504,N_693,N_657);
or U4505 (N_4505,N_71,N_938);
or U4506 (N_4506,N_1273,N_202);
nand U4507 (N_4507,N_1304,N_690);
and U4508 (N_4508,N_2082,N_1408);
nor U4509 (N_4509,N_458,N_1971);
or U4510 (N_4510,N_430,N_2088);
nand U4511 (N_4511,N_48,N_16);
or U4512 (N_4512,N_2460,N_2189);
and U4513 (N_4513,N_2254,N_1012);
nand U4514 (N_4514,N_1129,N_1963);
nor U4515 (N_4515,N_190,N_1126);
or U4516 (N_4516,N_2386,N_1475);
or U4517 (N_4517,N_1583,N_1946);
nor U4518 (N_4518,N_1487,N_801);
or U4519 (N_4519,N_2210,N_1569);
nor U4520 (N_4520,N_1997,N_1573);
or U4521 (N_4521,N_1206,N_505);
or U4522 (N_4522,N_2041,N_1698);
nor U4523 (N_4523,N_142,N_2045);
nor U4524 (N_4524,N_88,N_1606);
nand U4525 (N_4525,N_1787,N_2238);
or U4526 (N_4526,N_827,N_210);
nor U4527 (N_4527,N_650,N_2337);
nor U4528 (N_4528,N_1885,N_1790);
or U4529 (N_4529,N_454,N_503);
and U4530 (N_4530,N_1580,N_1357);
nand U4531 (N_4531,N_62,N_2223);
nand U4532 (N_4532,N_1229,N_948);
nor U4533 (N_4533,N_218,N_2008);
nand U4534 (N_4534,N_342,N_1743);
or U4535 (N_4535,N_1766,N_619);
or U4536 (N_4536,N_1626,N_311);
nor U4537 (N_4537,N_1717,N_1581);
or U4538 (N_4538,N_711,N_1248);
and U4539 (N_4539,N_927,N_383);
nand U4540 (N_4540,N_276,N_1056);
nor U4541 (N_4541,N_2183,N_1445);
and U4542 (N_4542,N_2275,N_1589);
or U4543 (N_4543,N_1256,N_1832);
nor U4544 (N_4544,N_1150,N_1381);
nand U4545 (N_4545,N_116,N_1959);
nand U4546 (N_4546,N_1334,N_2333);
nand U4547 (N_4547,N_2426,N_245);
nand U4548 (N_4548,N_2444,N_885);
nand U4549 (N_4549,N_860,N_126);
xor U4550 (N_4550,N_2342,N_1313);
nand U4551 (N_4551,N_1101,N_1929);
nand U4552 (N_4552,N_1660,N_408);
nor U4553 (N_4553,N_1228,N_934);
and U4554 (N_4554,N_933,N_1643);
or U4555 (N_4555,N_1672,N_1560);
and U4556 (N_4556,N_1059,N_1372);
nand U4557 (N_4557,N_1266,N_1432);
nor U4558 (N_4558,N_2110,N_737);
and U4559 (N_4559,N_1609,N_2458);
or U4560 (N_4560,N_1688,N_2482);
nand U4561 (N_4561,N_1803,N_1358);
nor U4562 (N_4562,N_1418,N_1281);
or U4563 (N_4563,N_882,N_376);
nand U4564 (N_4564,N_1981,N_1820);
nor U4565 (N_4565,N_1665,N_1900);
nand U4566 (N_4566,N_2370,N_834);
nand U4567 (N_4567,N_605,N_824);
nor U4568 (N_4568,N_798,N_1998);
nor U4569 (N_4569,N_1487,N_155);
and U4570 (N_4570,N_801,N_945);
and U4571 (N_4571,N_2182,N_137);
and U4572 (N_4572,N_2049,N_1330);
and U4573 (N_4573,N_2059,N_749);
nand U4574 (N_4574,N_2423,N_1156);
and U4575 (N_4575,N_1121,N_862);
xnor U4576 (N_4576,N_1731,N_1182);
or U4577 (N_4577,N_2074,N_2351);
or U4578 (N_4578,N_1162,N_1069);
nand U4579 (N_4579,N_312,N_1105);
and U4580 (N_4580,N_1053,N_1594);
nand U4581 (N_4581,N_1853,N_2406);
or U4582 (N_4582,N_1237,N_1606);
and U4583 (N_4583,N_1620,N_1661);
nand U4584 (N_4584,N_50,N_55);
nor U4585 (N_4585,N_2124,N_2325);
nand U4586 (N_4586,N_1030,N_130);
and U4587 (N_4587,N_134,N_1159);
or U4588 (N_4588,N_565,N_903);
nand U4589 (N_4589,N_258,N_1092);
nor U4590 (N_4590,N_428,N_2481);
or U4591 (N_4591,N_2015,N_139);
or U4592 (N_4592,N_467,N_2073);
or U4593 (N_4593,N_1519,N_449);
nand U4594 (N_4594,N_1441,N_1105);
and U4595 (N_4595,N_1800,N_927);
nor U4596 (N_4596,N_411,N_1433);
nand U4597 (N_4597,N_535,N_850);
nand U4598 (N_4598,N_154,N_948);
and U4599 (N_4599,N_2270,N_1036);
nor U4600 (N_4600,N_1169,N_2332);
and U4601 (N_4601,N_904,N_2057);
nor U4602 (N_4602,N_769,N_1001);
and U4603 (N_4603,N_739,N_1763);
and U4604 (N_4604,N_1168,N_854);
and U4605 (N_4605,N_1924,N_687);
nand U4606 (N_4606,N_2275,N_1923);
nor U4607 (N_4607,N_1191,N_2008);
or U4608 (N_4608,N_1810,N_93);
or U4609 (N_4609,N_857,N_527);
and U4610 (N_4610,N_475,N_1673);
and U4611 (N_4611,N_494,N_2279);
and U4612 (N_4612,N_1929,N_2432);
or U4613 (N_4613,N_1887,N_1136);
nand U4614 (N_4614,N_1011,N_102);
or U4615 (N_4615,N_841,N_1917);
nor U4616 (N_4616,N_692,N_1700);
nand U4617 (N_4617,N_1609,N_950);
nor U4618 (N_4618,N_1606,N_1105);
and U4619 (N_4619,N_2172,N_2004);
and U4620 (N_4620,N_818,N_1766);
xnor U4621 (N_4621,N_1975,N_225);
and U4622 (N_4622,N_866,N_1790);
nor U4623 (N_4623,N_1535,N_2359);
or U4624 (N_4624,N_1413,N_1084);
nor U4625 (N_4625,N_2260,N_2360);
xnor U4626 (N_4626,N_1152,N_1600);
or U4627 (N_4627,N_811,N_549);
and U4628 (N_4628,N_986,N_145);
nor U4629 (N_4629,N_2244,N_2265);
nand U4630 (N_4630,N_313,N_869);
and U4631 (N_4631,N_467,N_517);
nand U4632 (N_4632,N_463,N_997);
or U4633 (N_4633,N_2457,N_330);
nor U4634 (N_4634,N_965,N_567);
nand U4635 (N_4635,N_2200,N_737);
or U4636 (N_4636,N_1533,N_2013);
or U4637 (N_4637,N_1070,N_1881);
nor U4638 (N_4638,N_1587,N_511);
nor U4639 (N_4639,N_932,N_656);
nand U4640 (N_4640,N_981,N_2369);
or U4641 (N_4641,N_1985,N_82);
nor U4642 (N_4642,N_532,N_2236);
nand U4643 (N_4643,N_1973,N_468);
or U4644 (N_4644,N_1140,N_1949);
nand U4645 (N_4645,N_1879,N_203);
nor U4646 (N_4646,N_1007,N_143);
and U4647 (N_4647,N_700,N_2350);
or U4648 (N_4648,N_1522,N_962);
nand U4649 (N_4649,N_761,N_1748);
nand U4650 (N_4650,N_1790,N_380);
or U4651 (N_4651,N_861,N_2175);
or U4652 (N_4652,N_1984,N_1368);
nand U4653 (N_4653,N_832,N_2498);
xor U4654 (N_4654,N_1464,N_1784);
and U4655 (N_4655,N_2240,N_2306);
nor U4656 (N_4656,N_1978,N_1109);
xnor U4657 (N_4657,N_1459,N_1872);
nor U4658 (N_4658,N_1440,N_2214);
or U4659 (N_4659,N_1141,N_2016);
nand U4660 (N_4660,N_362,N_1121);
nand U4661 (N_4661,N_167,N_1250);
nor U4662 (N_4662,N_2354,N_564);
nor U4663 (N_4663,N_819,N_1959);
nor U4664 (N_4664,N_935,N_1477);
nor U4665 (N_4665,N_1919,N_2422);
and U4666 (N_4666,N_393,N_1693);
or U4667 (N_4667,N_2312,N_2495);
or U4668 (N_4668,N_557,N_1935);
nand U4669 (N_4669,N_1056,N_2048);
and U4670 (N_4670,N_826,N_417);
nor U4671 (N_4671,N_344,N_861);
nor U4672 (N_4672,N_1202,N_119);
and U4673 (N_4673,N_425,N_1021);
nor U4674 (N_4674,N_1390,N_1460);
or U4675 (N_4675,N_853,N_969);
or U4676 (N_4676,N_10,N_1721);
nand U4677 (N_4677,N_1280,N_2380);
nor U4678 (N_4678,N_709,N_106);
nand U4679 (N_4679,N_1496,N_2333);
or U4680 (N_4680,N_2272,N_1891);
nor U4681 (N_4681,N_1405,N_2377);
nor U4682 (N_4682,N_1948,N_1805);
nor U4683 (N_4683,N_5,N_1767);
and U4684 (N_4684,N_613,N_2101);
nand U4685 (N_4685,N_1793,N_1232);
or U4686 (N_4686,N_763,N_554);
nand U4687 (N_4687,N_1250,N_417);
or U4688 (N_4688,N_132,N_457);
and U4689 (N_4689,N_212,N_25);
or U4690 (N_4690,N_541,N_395);
nor U4691 (N_4691,N_1717,N_1497);
nand U4692 (N_4692,N_141,N_1774);
or U4693 (N_4693,N_1604,N_264);
and U4694 (N_4694,N_1315,N_2002);
or U4695 (N_4695,N_2066,N_676);
or U4696 (N_4696,N_2392,N_1956);
nor U4697 (N_4697,N_105,N_1758);
and U4698 (N_4698,N_1422,N_1465);
and U4699 (N_4699,N_1100,N_1433);
and U4700 (N_4700,N_555,N_1357);
and U4701 (N_4701,N_1122,N_1559);
and U4702 (N_4702,N_1283,N_1567);
nand U4703 (N_4703,N_1103,N_2403);
and U4704 (N_4704,N_193,N_1368);
or U4705 (N_4705,N_1679,N_1454);
nand U4706 (N_4706,N_1645,N_1093);
and U4707 (N_4707,N_527,N_447);
nor U4708 (N_4708,N_341,N_697);
and U4709 (N_4709,N_2414,N_1246);
or U4710 (N_4710,N_850,N_83);
nor U4711 (N_4711,N_1329,N_1290);
or U4712 (N_4712,N_210,N_1626);
and U4713 (N_4713,N_1067,N_2156);
and U4714 (N_4714,N_200,N_2070);
and U4715 (N_4715,N_1441,N_1648);
or U4716 (N_4716,N_2315,N_1827);
or U4717 (N_4717,N_1431,N_2408);
nor U4718 (N_4718,N_1095,N_2267);
nand U4719 (N_4719,N_214,N_2369);
nor U4720 (N_4720,N_2376,N_1826);
and U4721 (N_4721,N_1771,N_835);
nor U4722 (N_4722,N_313,N_1725);
or U4723 (N_4723,N_456,N_1551);
xnor U4724 (N_4724,N_454,N_2357);
nor U4725 (N_4725,N_33,N_851);
nor U4726 (N_4726,N_1548,N_1117);
nand U4727 (N_4727,N_80,N_160);
nor U4728 (N_4728,N_249,N_16);
nand U4729 (N_4729,N_1954,N_962);
nand U4730 (N_4730,N_2180,N_1511);
or U4731 (N_4731,N_1936,N_1918);
nand U4732 (N_4732,N_2102,N_2232);
or U4733 (N_4733,N_675,N_1253);
nand U4734 (N_4734,N_342,N_141);
nor U4735 (N_4735,N_1606,N_1847);
or U4736 (N_4736,N_2273,N_2250);
and U4737 (N_4737,N_83,N_2466);
and U4738 (N_4738,N_1843,N_2289);
nor U4739 (N_4739,N_1930,N_675);
or U4740 (N_4740,N_1512,N_429);
nand U4741 (N_4741,N_1734,N_906);
nand U4742 (N_4742,N_996,N_1854);
nand U4743 (N_4743,N_1651,N_12);
and U4744 (N_4744,N_1978,N_1252);
nor U4745 (N_4745,N_1088,N_1290);
and U4746 (N_4746,N_402,N_2215);
and U4747 (N_4747,N_487,N_1145);
or U4748 (N_4748,N_1969,N_1722);
nor U4749 (N_4749,N_146,N_2346);
and U4750 (N_4750,N_1904,N_1847);
and U4751 (N_4751,N_1517,N_1998);
nand U4752 (N_4752,N_162,N_787);
and U4753 (N_4753,N_1492,N_646);
xnor U4754 (N_4754,N_511,N_2478);
xor U4755 (N_4755,N_1634,N_81);
xor U4756 (N_4756,N_928,N_2221);
nor U4757 (N_4757,N_119,N_155);
nor U4758 (N_4758,N_1735,N_1772);
and U4759 (N_4759,N_1917,N_1670);
or U4760 (N_4760,N_2139,N_1374);
nand U4761 (N_4761,N_47,N_1588);
nor U4762 (N_4762,N_1234,N_577);
nand U4763 (N_4763,N_2457,N_1407);
nor U4764 (N_4764,N_1542,N_863);
nor U4765 (N_4765,N_875,N_1995);
or U4766 (N_4766,N_1962,N_1511);
or U4767 (N_4767,N_1478,N_130);
and U4768 (N_4768,N_1038,N_1973);
or U4769 (N_4769,N_510,N_1351);
nor U4770 (N_4770,N_2402,N_1671);
and U4771 (N_4771,N_2136,N_1121);
or U4772 (N_4772,N_1315,N_1902);
nor U4773 (N_4773,N_1480,N_654);
nor U4774 (N_4774,N_2440,N_1674);
or U4775 (N_4775,N_53,N_2187);
and U4776 (N_4776,N_1469,N_738);
and U4777 (N_4777,N_1515,N_1097);
and U4778 (N_4778,N_986,N_1065);
and U4779 (N_4779,N_1442,N_339);
nand U4780 (N_4780,N_2096,N_1250);
or U4781 (N_4781,N_2469,N_2228);
nand U4782 (N_4782,N_621,N_2211);
or U4783 (N_4783,N_220,N_2016);
or U4784 (N_4784,N_0,N_1874);
or U4785 (N_4785,N_382,N_2251);
nand U4786 (N_4786,N_502,N_820);
nor U4787 (N_4787,N_1190,N_2373);
nand U4788 (N_4788,N_612,N_1614);
and U4789 (N_4789,N_1480,N_1687);
nor U4790 (N_4790,N_693,N_1501);
nand U4791 (N_4791,N_1626,N_2256);
and U4792 (N_4792,N_1152,N_1444);
nor U4793 (N_4793,N_1131,N_1676);
nand U4794 (N_4794,N_603,N_1521);
nor U4795 (N_4795,N_53,N_168);
and U4796 (N_4796,N_235,N_1185);
or U4797 (N_4797,N_2333,N_2440);
or U4798 (N_4798,N_81,N_2478);
nand U4799 (N_4799,N_1815,N_1427);
nand U4800 (N_4800,N_6,N_1988);
nor U4801 (N_4801,N_371,N_429);
nor U4802 (N_4802,N_1613,N_2242);
nand U4803 (N_4803,N_474,N_517);
nor U4804 (N_4804,N_1870,N_1936);
nand U4805 (N_4805,N_156,N_538);
nand U4806 (N_4806,N_1109,N_1282);
or U4807 (N_4807,N_2476,N_2275);
nor U4808 (N_4808,N_1428,N_1277);
and U4809 (N_4809,N_1215,N_1713);
nor U4810 (N_4810,N_2304,N_117);
or U4811 (N_4811,N_613,N_2194);
nor U4812 (N_4812,N_589,N_2020);
and U4813 (N_4813,N_869,N_818);
nand U4814 (N_4814,N_71,N_1370);
nor U4815 (N_4815,N_1630,N_2468);
and U4816 (N_4816,N_1949,N_802);
or U4817 (N_4817,N_998,N_1527);
nor U4818 (N_4818,N_1960,N_272);
nand U4819 (N_4819,N_336,N_525);
or U4820 (N_4820,N_1894,N_1911);
nor U4821 (N_4821,N_873,N_2361);
or U4822 (N_4822,N_769,N_1875);
and U4823 (N_4823,N_1420,N_1577);
and U4824 (N_4824,N_528,N_649);
and U4825 (N_4825,N_586,N_354);
nor U4826 (N_4826,N_1329,N_4);
nand U4827 (N_4827,N_2023,N_165);
and U4828 (N_4828,N_2110,N_631);
nor U4829 (N_4829,N_1335,N_2099);
nand U4830 (N_4830,N_2111,N_2207);
and U4831 (N_4831,N_2476,N_2206);
nor U4832 (N_4832,N_2104,N_1526);
or U4833 (N_4833,N_2223,N_360);
or U4834 (N_4834,N_2226,N_1863);
and U4835 (N_4835,N_2246,N_892);
nor U4836 (N_4836,N_274,N_96);
and U4837 (N_4837,N_921,N_647);
or U4838 (N_4838,N_2007,N_632);
and U4839 (N_4839,N_1777,N_1925);
nand U4840 (N_4840,N_488,N_901);
nand U4841 (N_4841,N_2451,N_628);
and U4842 (N_4842,N_1706,N_840);
nor U4843 (N_4843,N_2308,N_2432);
nor U4844 (N_4844,N_121,N_2008);
or U4845 (N_4845,N_804,N_1225);
nor U4846 (N_4846,N_1055,N_2036);
or U4847 (N_4847,N_1444,N_1638);
or U4848 (N_4848,N_1468,N_1150);
and U4849 (N_4849,N_2249,N_1324);
and U4850 (N_4850,N_2363,N_2083);
and U4851 (N_4851,N_1373,N_2179);
nand U4852 (N_4852,N_2047,N_349);
or U4853 (N_4853,N_2312,N_2022);
and U4854 (N_4854,N_1261,N_794);
nand U4855 (N_4855,N_265,N_573);
nor U4856 (N_4856,N_1237,N_1457);
nor U4857 (N_4857,N_613,N_531);
nand U4858 (N_4858,N_2010,N_1571);
and U4859 (N_4859,N_1701,N_911);
or U4860 (N_4860,N_754,N_2262);
nand U4861 (N_4861,N_1834,N_851);
or U4862 (N_4862,N_2182,N_508);
and U4863 (N_4863,N_189,N_401);
nand U4864 (N_4864,N_276,N_1437);
nand U4865 (N_4865,N_1774,N_1857);
and U4866 (N_4866,N_2015,N_1094);
nor U4867 (N_4867,N_2305,N_764);
nor U4868 (N_4868,N_2460,N_1306);
or U4869 (N_4869,N_1728,N_1867);
and U4870 (N_4870,N_1298,N_708);
or U4871 (N_4871,N_1749,N_2403);
or U4872 (N_4872,N_893,N_1798);
or U4873 (N_4873,N_418,N_166);
nor U4874 (N_4874,N_955,N_1956);
nor U4875 (N_4875,N_555,N_736);
and U4876 (N_4876,N_1754,N_272);
nand U4877 (N_4877,N_385,N_2140);
nand U4878 (N_4878,N_1649,N_721);
or U4879 (N_4879,N_1237,N_1652);
nor U4880 (N_4880,N_2211,N_651);
and U4881 (N_4881,N_1329,N_1508);
or U4882 (N_4882,N_453,N_1163);
and U4883 (N_4883,N_291,N_974);
and U4884 (N_4884,N_953,N_1);
and U4885 (N_4885,N_1338,N_1621);
or U4886 (N_4886,N_197,N_2178);
and U4887 (N_4887,N_2284,N_949);
and U4888 (N_4888,N_630,N_149);
nor U4889 (N_4889,N_952,N_284);
nand U4890 (N_4890,N_1152,N_230);
nor U4891 (N_4891,N_1005,N_2186);
nor U4892 (N_4892,N_1081,N_2263);
nand U4893 (N_4893,N_1623,N_2024);
or U4894 (N_4894,N_2223,N_1182);
nor U4895 (N_4895,N_2121,N_1149);
and U4896 (N_4896,N_2053,N_1578);
or U4897 (N_4897,N_1286,N_2341);
nand U4898 (N_4898,N_283,N_440);
or U4899 (N_4899,N_44,N_1837);
nor U4900 (N_4900,N_577,N_203);
and U4901 (N_4901,N_474,N_1125);
and U4902 (N_4902,N_2089,N_692);
and U4903 (N_4903,N_2129,N_329);
and U4904 (N_4904,N_1317,N_125);
nor U4905 (N_4905,N_892,N_1798);
xor U4906 (N_4906,N_1909,N_2207);
nand U4907 (N_4907,N_2469,N_2492);
or U4908 (N_4908,N_1513,N_485);
or U4909 (N_4909,N_806,N_848);
or U4910 (N_4910,N_2294,N_1435);
or U4911 (N_4911,N_2283,N_1129);
and U4912 (N_4912,N_800,N_663);
and U4913 (N_4913,N_1702,N_1558);
xnor U4914 (N_4914,N_2018,N_376);
nand U4915 (N_4915,N_1157,N_1489);
xor U4916 (N_4916,N_1699,N_2095);
nand U4917 (N_4917,N_1368,N_1850);
nor U4918 (N_4918,N_2170,N_317);
nand U4919 (N_4919,N_1744,N_487);
xnor U4920 (N_4920,N_1583,N_1122);
or U4921 (N_4921,N_1940,N_709);
nand U4922 (N_4922,N_1411,N_2153);
nor U4923 (N_4923,N_1981,N_103);
or U4924 (N_4924,N_349,N_238);
nand U4925 (N_4925,N_1102,N_999);
nand U4926 (N_4926,N_1762,N_501);
nor U4927 (N_4927,N_138,N_1948);
nor U4928 (N_4928,N_2042,N_1399);
or U4929 (N_4929,N_2455,N_1170);
or U4930 (N_4930,N_506,N_190);
nand U4931 (N_4931,N_1160,N_229);
nor U4932 (N_4932,N_1943,N_559);
and U4933 (N_4933,N_549,N_2441);
and U4934 (N_4934,N_1236,N_2442);
nand U4935 (N_4935,N_2256,N_501);
and U4936 (N_4936,N_1661,N_2132);
or U4937 (N_4937,N_244,N_415);
or U4938 (N_4938,N_2299,N_1805);
xnor U4939 (N_4939,N_1106,N_850);
and U4940 (N_4940,N_534,N_887);
xnor U4941 (N_4941,N_850,N_960);
or U4942 (N_4942,N_2281,N_1963);
nand U4943 (N_4943,N_1706,N_1216);
nand U4944 (N_4944,N_2223,N_1505);
or U4945 (N_4945,N_2354,N_295);
nand U4946 (N_4946,N_2126,N_1698);
nand U4947 (N_4947,N_1138,N_51);
and U4948 (N_4948,N_28,N_713);
or U4949 (N_4949,N_2165,N_1145);
nand U4950 (N_4950,N_1855,N_1199);
nor U4951 (N_4951,N_2381,N_289);
and U4952 (N_4952,N_2031,N_1129);
or U4953 (N_4953,N_383,N_1257);
or U4954 (N_4954,N_1815,N_718);
and U4955 (N_4955,N_1199,N_1090);
nand U4956 (N_4956,N_1557,N_665);
nand U4957 (N_4957,N_80,N_666);
or U4958 (N_4958,N_251,N_761);
or U4959 (N_4959,N_273,N_2316);
or U4960 (N_4960,N_600,N_149);
and U4961 (N_4961,N_706,N_1417);
and U4962 (N_4962,N_2055,N_758);
and U4963 (N_4963,N_1262,N_2248);
nand U4964 (N_4964,N_1321,N_2338);
nand U4965 (N_4965,N_345,N_1292);
nor U4966 (N_4966,N_2151,N_457);
nor U4967 (N_4967,N_229,N_1722);
nand U4968 (N_4968,N_2222,N_1285);
or U4969 (N_4969,N_2072,N_2245);
nor U4970 (N_4970,N_1293,N_86);
nand U4971 (N_4971,N_1450,N_791);
nor U4972 (N_4972,N_2299,N_2287);
or U4973 (N_4973,N_1855,N_2141);
or U4974 (N_4974,N_540,N_1475);
and U4975 (N_4975,N_2080,N_288);
or U4976 (N_4976,N_1175,N_130);
or U4977 (N_4977,N_1474,N_2329);
nand U4978 (N_4978,N_2475,N_1146);
nand U4979 (N_4979,N_1113,N_1330);
xnor U4980 (N_4980,N_1450,N_2339);
and U4981 (N_4981,N_1010,N_2228);
or U4982 (N_4982,N_1086,N_187);
and U4983 (N_4983,N_874,N_1971);
and U4984 (N_4984,N_1857,N_110);
nand U4985 (N_4985,N_1571,N_832);
or U4986 (N_4986,N_1597,N_1611);
and U4987 (N_4987,N_1881,N_400);
or U4988 (N_4988,N_1742,N_1197);
and U4989 (N_4989,N_1152,N_1720);
nand U4990 (N_4990,N_2440,N_2005);
and U4991 (N_4991,N_1866,N_225);
and U4992 (N_4992,N_279,N_2192);
nor U4993 (N_4993,N_948,N_400);
nand U4994 (N_4994,N_943,N_1343);
and U4995 (N_4995,N_1028,N_2276);
or U4996 (N_4996,N_2083,N_826);
and U4997 (N_4997,N_880,N_1353);
or U4998 (N_4998,N_243,N_2142);
and U4999 (N_4999,N_2176,N_1625);
and UO_0 (O_0,N_4069,N_2580);
or UO_1 (O_1,N_2577,N_4594);
or UO_2 (O_2,N_3481,N_4662);
nor UO_3 (O_3,N_4448,N_2894);
and UO_4 (O_4,N_4092,N_4579);
nor UO_5 (O_5,N_3457,N_4458);
and UO_6 (O_6,N_3401,N_4454);
or UO_7 (O_7,N_3870,N_3300);
nor UO_8 (O_8,N_4207,N_3367);
and UO_9 (O_9,N_3965,N_2504);
nand UO_10 (O_10,N_3848,N_3049);
nand UO_11 (O_11,N_2694,N_4129);
and UO_12 (O_12,N_2807,N_4223);
nor UO_13 (O_13,N_4191,N_2605);
nor UO_14 (O_14,N_4452,N_3179);
nor UO_15 (O_15,N_4910,N_3275);
nor UO_16 (O_16,N_2736,N_4338);
nor UO_17 (O_17,N_4830,N_4668);
nand UO_18 (O_18,N_3140,N_3137);
nand UO_19 (O_19,N_3369,N_4731);
or UO_20 (O_20,N_4349,N_3387);
and UO_21 (O_21,N_3424,N_3584);
xor UO_22 (O_22,N_4553,N_3734);
or UO_23 (O_23,N_3573,N_2937);
nor UO_24 (O_24,N_4610,N_3947);
nor UO_25 (O_25,N_2941,N_2978);
nor UO_26 (O_26,N_2600,N_3686);
nand UO_27 (O_27,N_2615,N_4147);
nor UO_28 (O_28,N_4235,N_2977);
xnor UO_29 (O_29,N_3507,N_4382);
nand UO_30 (O_30,N_4016,N_4257);
and UO_31 (O_31,N_3143,N_4456);
or UO_32 (O_32,N_4365,N_2723);
and UO_33 (O_33,N_3914,N_4154);
or UO_34 (O_34,N_4916,N_3277);
nand UO_35 (O_35,N_3471,N_4360);
and UO_36 (O_36,N_4204,N_4011);
nand UO_37 (O_37,N_3813,N_3607);
or UO_38 (O_38,N_4877,N_4739);
and UO_39 (O_39,N_2857,N_3370);
and UO_40 (O_40,N_2656,N_2728);
and UO_41 (O_41,N_4937,N_4394);
nor UO_42 (O_42,N_4339,N_4078);
or UO_43 (O_43,N_4388,N_3858);
nor UO_44 (O_44,N_4391,N_3543);
and UO_45 (O_45,N_3174,N_3034);
or UO_46 (O_46,N_4636,N_3633);
or UO_47 (O_47,N_4987,N_4463);
nand UO_48 (O_48,N_4209,N_3355);
and UO_49 (O_49,N_4522,N_3827);
nor UO_50 (O_50,N_4549,N_4478);
xnor UO_51 (O_51,N_3232,N_3772);
or UO_52 (O_52,N_3583,N_3504);
nand UO_53 (O_53,N_4997,N_3644);
nand UO_54 (O_54,N_3107,N_4761);
nor UO_55 (O_55,N_4145,N_3043);
or UO_56 (O_56,N_4659,N_3156);
nor UO_57 (O_57,N_4237,N_2856);
nor UO_58 (O_58,N_3499,N_3243);
xor UO_59 (O_59,N_4459,N_4157);
or UO_60 (O_60,N_2682,N_3922);
nand UO_61 (O_61,N_3605,N_3245);
nor UO_62 (O_62,N_4898,N_2885);
nor UO_63 (O_63,N_4065,N_2926);
and UO_64 (O_64,N_3552,N_4967);
or UO_65 (O_65,N_2538,N_3376);
and UO_66 (O_66,N_3956,N_4642);
nand UO_67 (O_67,N_4759,N_4979);
or UO_68 (O_68,N_3781,N_4494);
or UO_69 (O_69,N_4352,N_2510);
or UO_70 (O_70,N_3170,N_3845);
nor UO_71 (O_71,N_2843,N_3364);
nand UO_72 (O_72,N_3184,N_4990);
nand UO_73 (O_73,N_3654,N_4824);
and UO_74 (O_74,N_4377,N_2693);
or UO_75 (O_75,N_3771,N_4429);
or UO_76 (O_76,N_4801,N_4942);
nor UO_77 (O_77,N_3475,N_4032);
nor UO_78 (O_78,N_4012,N_4404);
or UO_79 (O_79,N_3057,N_3058);
and UO_80 (O_80,N_2909,N_4473);
nand UO_81 (O_81,N_2610,N_2502);
nor UO_82 (O_82,N_4149,N_2752);
and UO_83 (O_83,N_4657,N_4407);
nor UO_84 (O_84,N_4983,N_3812);
nand UO_85 (O_85,N_2601,N_4146);
and UO_86 (O_86,N_3941,N_3375);
nand UO_87 (O_87,N_4837,N_4169);
and UO_88 (O_88,N_4006,N_4326);
nor UO_89 (O_89,N_3306,N_4595);
nand UO_90 (O_90,N_3070,N_3167);
or UO_91 (O_91,N_2583,N_3670);
or UO_92 (O_92,N_4405,N_2936);
or UO_93 (O_93,N_4173,N_2663);
nand UO_94 (O_94,N_4418,N_3697);
nor UO_95 (O_95,N_3849,N_4998);
nor UO_96 (O_96,N_4320,N_4165);
nand UO_97 (O_97,N_2835,N_4482);
or UO_98 (O_98,N_4711,N_3695);
nor UO_99 (O_99,N_2674,N_4834);
nor UO_100 (O_100,N_2581,N_3632);
or UO_101 (O_101,N_3558,N_2773);
nor UO_102 (O_102,N_4229,N_3018);
or UO_103 (O_103,N_3196,N_3619);
or UO_104 (O_104,N_2922,N_3470);
nor UO_105 (O_105,N_4890,N_3193);
nand UO_106 (O_106,N_2588,N_4712);
nand UO_107 (O_107,N_3227,N_4767);
nor UO_108 (O_108,N_3694,N_4563);
nor UO_109 (O_109,N_3727,N_4144);
nor UO_110 (O_110,N_4426,N_3357);
and UO_111 (O_111,N_3720,N_4019);
and UO_112 (O_112,N_3566,N_3880);
or UO_113 (O_113,N_2819,N_4323);
and UO_114 (O_114,N_4284,N_4740);
or UO_115 (O_115,N_3877,N_4218);
nand UO_116 (O_116,N_3790,N_3303);
nor UO_117 (O_117,N_3902,N_3796);
and UO_118 (O_118,N_4756,N_4649);
or UO_119 (O_119,N_4384,N_2590);
xor UO_120 (O_120,N_2612,N_3222);
or UO_121 (O_121,N_4021,N_3450);
nand UO_122 (O_122,N_2893,N_4166);
and UO_123 (O_123,N_2543,N_3012);
or UO_124 (O_124,N_2940,N_4495);
nand UO_125 (O_125,N_3478,N_4918);
nor UO_126 (O_126,N_3320,N_4420);
nand UO_127 (O_127,N_3060,N_3359);
nor UO_128 (O_128,N_2742,N_2943);
and UO_129 (O_129,N_3911,N_3065);
and UO_130 (O_130,N_4564,N_2633);
and UO_131 (O_131,N_3373,N_4670);
nand UO_132 (O_132,N_3489,N_4633);
nand UO_133 (O_133,N_4051,N_3462);
nor UO_134 (O_134,N_3970,N_3305);
or UO_135 (O_135,N_2602,N_4823);
or UO_136 (O_136,N_3051,N_2659);
and UO_137 (O_137,N_4699,N_2686);
nor UO_138 (O_138,N_2560,N_3212);
or UO_139 (O_139,N_3520,N_2877);
nand UO_140 (O_140,N_4764,N_3186);
nand UO_141 (O_141,N_3208,N_3608);
nand UO_142 (O_142,N_4913,N_4954);
nand UO_143 (O_143,N_4340,N_4307);
and UO_144 (O_144,N_4200,N_3229);
or UO_145 (O_145,N_2520,N_4952);
xor UO_146 (O_146,N_4726,N_3621);
nand UO_147 (O_147,N_4735,N_2673);
and UO_148 (O_148,N_3872,N_4311);
nand UO_149 (O_149,N_3444,N_2867);
nand UO_150 (O_150,N_4462,N_2529);
nand UO_151 (O_151,N_3221,N_4308);
nand UO_152 (O_152,N_4253,N_3936);
nand UO_153 (O_153,N_2541,N_4118);
nand UO_154 (O_154,N_2814,N_3078);
nor UO_155 (O_155,N_3587,N_3415);
or UO_156 (O_156,N_4160,N_3120);
or UO_157 (O_157,N_2995,N_3333);
nand UO_158 (O_158,N_4556,N_3515);
nor UO_159 (O_159,N_4698,N_4471);
or UO_160 (O_160,N_2658,N_3850);
or UO_161 (O_161,N_4423,N_4085);
or UO_162 (O_162,N_3076,N_4846);
nor UO_163 (O_163,N_4677,N_4373);
nand UO_164 (O_164,N_2678,N_4647);
or UO_165 (O_165,N_4899,N_4356);
or UO_166 (O_166,N_2864,N_3765);
nand UO_167 (O_167,N_2774,N_3650);
nor UO_168 (O_168,N_3793,N_4869);
xor UO_169 (O_169,N_4222,N_3591);
and UO_170 (O_170,N_3477,N_3464);
xnor UO_171 (O_171,N_3602,N_3726);
and UO_172 (O_172,N_3066,N_4521);
nand UO_173 (O_173,N_2688,N_3716);
nand UO_174 (O_174,N_3755,N_4119);
nand UO_175 (O_175,N_3576,N_2669);
or UO_176 (O_176,N_2838,N_2696);
nand UO_177 (O_177,N_4206,N_2690);
nor UO_178 (O_178,N_2907,N_3220);
nand UO_179 (O_179,N_4685,N_3618);
or UO_180 (O_180,N_4907,N_3425);
nand UO_181 (O_181,N_4867,N_4684);
nand UO_182 (O_182,N_3568,N_3334);
nor UO_183 (O_183,N_4334,N_4108);
nor UO_184 (O_184,N_3085,N_2769);
xor UO_185 (O_185,N_3004,N_3996);
nor UO_186 (O_186,N_4470,N_3438);
nand UO_187 (O_187,N_2892,N_3948);
or UO_188 (O_188,N_4661,N_3326);
nand UO_189 (O_189,N_2879,N_3068);
xnor UO_190 (O_190,N_2859,N_2965);
nand UO_191 (O_191,N_2961,N_4908);
or UO_192 (O_192,N_4639,N_2671);
and UO_193 (O_193,N_3603,N_3412);
nand UO_194 (O_194,N_3487,N_2553);
nor UO_195 (O_195,N_4542,N_4883);
and UO_196 (O_196,N_4591,N_3157);
or UO_197 (O_197,N_4971,N_3545);
nor UO_198 (O_198,N_3652,N_4194);
and UO_199 (O_199,N_4389,N_3131);
nor UO_200 (O_200,N_3149,N_3801);
and UO_201 (O_201,N_4982,N_2614);
or UO_202 (O_202,N_4619,N_4743);
nor UO_203 (O_203,N_4729,N_4826);
nor UO_204 (O_204,N_4026,N_3189);
and UO_205 (O_205,N_4810,N_2500);
nor UO_206 (O_206,N_4057,N_4999);
and UO_207 (O_207,N_2536,N_3083);
nor UO_208 (O_208,N_2972,N_3540);
and UO_209 (O_209,N_2547,N_3867);
and UO_210 (O_210,N_3238,N_4054);
nor UO_211 (O_211,N_3073,N_2828);
and UO_212 (O_212,N_3183,N_3722);
nand UO_213 (O_213,N_4479,N_4502);
nor UO_214 (O_214,N_4605,N_3324);
and UO_215 (O_215,N_2797,N_3869);
nor UO_216 (O_216,N_2993,N_3017);
or UO_217 (O_217,N_4947,N_4246);
nor UO_218 (O_218,N_4300,N_3466);
or UO_219 (O_219,N_3339,N_4059);
nand UO_220 (O_220,N_4955,N_4500);
or UO_221 (O_221,N_3749,N_3767);
or UO_222 (O_222,N_3714,N_4551);
nor UO_223 (O_223,N_3980,N_2732);
nor UO_224 (O_224,N_4607,N_2639);
or UO_225 (O_225,N_3028,N_3917);
nand UO_226 (O_226,N_4621,N_3901);
or UO_227 (O_227,N_4745,N_2914);
nor UO_228 (O_228,N_3294,N_3704);
and UO_229 (O_229,N_3103,N_3461);
or UO_230 (O_230,N_3211,N_3032);
nand UO_231 (O_231,N_3728,N_2569);
or UO_232 (O_232,N_4734,N_2853);
and UO_233 (O_233,N_4989,N_2757);
and UO_234 (O_234,N_3029,N_4055);
or UO_235 (O_235,N_4920,N_2829);
nand UO_236 (O_236,N_4236,N_3077);
nand UO_237 (O_237,N_4211,N_3488);
or UO_238 (O_238,N_2516,N_2662);
nor UO_239 (O_239,N_3628,N_4557);
and UO_240 (O_240,N_4921,N_3316);
and UO_241 (O_241,N_2613,N_4023);
or UO_242 (O_242,N_4787,N_3895);
and UO_243 (O_243,N_3890,N_4477);
or UO_244 (O_244,N_2683,N_2532);
nand UO_245 (O_245,N_4513,N_4849);
or UO_246 (O_246,N_3349,N_4139);
or UO_247 (O_247,N_4782,N_2905);
or UO_248 (O_248,N_2623,N_4815);
nor UO_249 (O_249,N_3811,N_4758);
and UO_250 (O_250,N_3557,N_3379);
or UO_251 (O_251,N_2755,N_3247);
nor UO_252 (O_252,N_4576,N_4140);
or UO_253 (O_253,N_4168,N_4574);
nor UO_254 (O_254,N_4985,N_4737);
and UO_255 (O_255,N_4344,N_3685);
nand UO_256 (O_256,N_3799,N_4577);
nand UO_257 (O_257,N_4765,N_3883);
nand UO_258 (O_258,N_4820,N_4052);
nand UO_259 (O_259,N_3235,N_3114);
nor UO_260 (O_260,N_3141,N_2524);
nor UO_261 (O_261,N_2597,N_4766);
nand UO_262 (O_262,N_4313,N_4440);
and UO_263 (O_263,N_3023,N_2608);
nor UO_264 (O_264,N_3445,N_4199);
nor UO_265 (O_265,N_4879,N_4704);
or UO_266 (O_266,N_2872,N_3741);
nand UO_267 (O_267,N_3861,N_3224);
nor UO_268 (O_268,N_2729,N_3862);
nor UO_269 (O_269,N_4852,N_2776);
or UO_270 (O_270,N_4695,N_3002);
nand UO_271 (O_271,N_3977,N_3182);
xnor UO_272 (O_272,N_3109,N_4507);
and UO_273 (O_273,N_4733,N_4335);
nor UO_274 (O_274,N_4530,N_3896);
nand UO_275 (O_275,N_3614,N_3606);
xor UO_276 (O_276,N_2622,N_4421);
nor UO_277 (O_277,N_4089,N_3855);
nor UO_278 (O_278,N_3037,N_4893);
and UO_279 (O_279,N_4106,N_4183);
nor UO_280 (O_280,N_4105,N_4926);
nand UO_281 (O_281,N_3846,N_3888);
or UO_282 (O_282,N_3553,N_3842);
or UO_283 (O_283,N_4968,N_4537);
nand UO_284 (O_284,N_2979,N_3069);
nand UO_285 (O_285,N_4254,N_2548);
nand UO_286 (O_286,N_4221,N_3194);
or UO_287 (O_287,N_3297,N_2949);
or UO_288 (O_288,N_2966,N_4009);
nor UO_289 (O_289,N_3671,N_3352);
or UO_290 (O_290,N_3903,N_3806);
or UO_291 (O_291,N_3809,N_4671);
xnor UO_292 (O_292,N_3164,N_3544);
and UO_293 (O_293,N_2572,N_3332);
xor UO_294 (O_294,N_2619,N_3505);
nand UO_295 (O_295,N_4874,N_3763);
nor UO_296 (O_296,N_3292,N_4301);
or UO_297 (O_297,N_3127,N_3974);
and UO_298 (O_298,N_3059,N_4451);
or UO_299 (O_299,N_4857,N_4931);
nor UO_300 (O_300,N_3777,N_4318);
and UO_301 (O_301,N_4682,N_4214);
xor UO_302 (O_302,N_3175,N_4850);
or UO_303 (O_303,N_4757,N_3512);
nand UO_304 (O_304,N_4098,N_3593);
or UO_305 (O_305,N_4004,N_3213);
and UO_306 (O_306,N_3011,N_3629);
nor UO_307 (O_307,N_4793,N_4602);
nand UO_308 (O_308,N_3240,N_3223);
and UO_309 (O_309,N_2650,N_4569);
or UO_310 (O_310,N_2855,N_3105);
or UO_311 (O_311,N_3841,N_4707);
xnor UO_312 (O_312,N_3912,N_4529);
nand UO_313 (O_313,N_3875,N_3108);
nor UO_314 (O_314,N_4374,N_3718);
and UO_315 (O_315,N_2869,N_4821);
and UO_316 (O_316,N_3144,N_4656);
or UO_317 (O_317,N_3272,N_2717);
nand UO_318 (O_318,N_3350,N_2689);
nand UO_319 (O_319,N_4748,N_3791);
nand UO_320 (O_320,N_4870,N_3256);
or UO_321 (O_321,N_3392,N_3945);
nand UO_322 (O_322,N_3524,N_3535);
nor UO_323 (O_323,N_3531,N_3119);
nor UO_324 (O_324,N_4791,N_3061);
and UO_325 (O_325,N_4252,N_3572);
and UO_326 (O_326,N_4369,N_4878);
and UO_327 (O_327,N_2987,N_4104);
nand UO_328 (O_328,N_4832,N_4449);
or UO_329 (O_329,N_3537,N_2595);
or UO_330 (O_330,N_2854,N_2668);
or UO_331 (O_331,N_3853,N_4036);
and UO_332 (O_332,N_3407,N_2737);
or UO_333 (O_333,N_4273,N_3511);
nor UO_334 (O_334,N_2620,N_4136);
and UO_335 (O_335,N_4804,N_3634);
nand UO_336 (O_336,N_3851,N_3093);
and UO_337 (O_337,N_2706,N_2539);
nor UO_338 (O_338,N_2604,N_3863);
and UO_339 (O_339,N_2596,N_2570);
nand UO_340 (O_340,N_4038,N_3635);
nand UO_341 (O_341,N_4841,N_3242);
nand UO_342 (O_342,N_3480,N_3117);
and UO_343 (O_343,N_4615,N_4468);
nand UO_344 (O_344,N_4750,N_2772);
nor UO_345 (O_345,N_4436,N_2822);
or UO_346 (O_346,N_4770,N_4526);
and UO_347 (O_347,N_4445,N_2782);
nand UO_348 (O_348,N_2738,N_4283);
nor UO_349 (O_349,N_3989,N_4792);
nor UO_350 (O_350,N_2803,N_2632);
and UO_351 (O_351,N_3092,N_4289);
and UO_352 (O_352,N_2703,N_4457);
nand UO_353 (O_353,N_3805,N_2889);
or UO_354 (O_354,N_3787,N_3062);
or UO_355 (O_355,N_2733,N_3645);
nand UO_356 (O_356,N_2839,N_3325);
nor UO_357 (O_357,N_4822,N_3651);
nor UO_358 (O_358,N_4381,N_3166);
nand UO_359 (O_359,N_3983,N_4064);
nor UO_360 (O_360,N_4115,N_4512);
nor UO_361 (O_361,N_2519,N_3408);
nor UO_362 (O_362,N_4719,N_4484);
and UO_363 (O_363,N_4799,N_3001);
and UO_364 (O_364,N_4328,N_3709);
nor UO_365 (O_365,N_4066,N_3735);
and UO_366 (O_366,N_2802,N_4143);
nor UO_367 (O_367,N_3155,N_2917);
and UO_368 (O_368,N_4042,N_2935);
and UO_369 (O_369,N_3937,N_2848);
or UO_370 (O_370,N_3399,N_4232);
and UO_371 (O_371,N_2874,N_4071);
nor UO_372 (O_372,N_4306,N_4097);
or UO_373 (O_373,N_4258,N_2777);
or UO_374 (O_374,N_3723,N_4017);
xnor UO_375 (O_375,N_4286,N_3824);
nor UO_376 (O_376,N_2714,N_4072);
and UO_377 (O_377,N_4861,N_3631);
and UO_378 (O_378,N_4583,N_4800);
nand UO_379 (O_379,N_3762,N_3643);
and UO_380 (O_380,N_2518,N_2603);
and UO_381 (O_381,N_4807,N_3669);
nand UO_382 (O_382,N_4035,N_4570);
nor UO_383 (O_383,N_4972,N_2832);
nor UO_384 (O_384,N_3700,N_4567);
and UO_385 (O_385,N_4665,N_2811);
or UO_386 (O_386,N_4944,N_4613);
nand UO_387 (O_387,N_4047,N_3810);
or UO_388 (O_388,N_3807,N_4399);
and UO_389 (O_389,N_3808,N_4465);
and UO_390 (O_390,N_3088,N_4742);
nor UO_391 (O_391,N_4263,N_3889);
nand UO_392 (O_392,N_3234,N_4592);
and UO_393 (O_393,N_3831,N_4620);
nand UO_394 (O_394,N_2908,N_3900);
nand UO_395 (O_395,N_2508,N_3123);
or UO_396 (O_396,N_3750,N_3162);
nor UO_397 (O_397,N_3427,N_4342);
or UO_398 (O_398,N_4278,N_2712);
nand UO_399 (O_399,N_3800,N_2643);
or UO_400 (O_400,N_2760,N_4536);
or UO_401 (O_401,N_3973,N_3266);
and UO_402 (O_402,N_4304,N_3097);
or UO_403 (O_403,N_4132,N_2708);
and UO_404 (O_404,N_2826,N_3832);
or UO_405 (O_405,N_4928,N_3792);
nor UO_406 (O_406,N_4970,N_4584);
or UO_407 (O_407,N_3257,N_3926);
nor UO_408 (O_408,N_2545,N_3997);
nand UO_409 (O_409,N_4614,N_3666);
nor UO_410 (O_410,N_4650,N_3856);
or UO_411 (O_411,N_3857,N_4887);
xnor UO_412 (O_412,N_2745,N_2637);
xnor UO_413 (O_413,N_3636,N_2933);
nor UO_414 (O_414,N_3898,N_2544);
xnor UO_415 (O_415,N_3508,N_4073);
nor UO_416 (O_416,N_2763,N_3460);
or UO_417 (O_417,N_4814,N_4566);
and UO_418 (O_418,N_3639,N_3910);
nand UO_419 (O_419,N_2945,N_2982);
nor UO_420 (O_420,N_2679,N_3676);
or UO_421 (O_421,N_3330,N_4505);
and UO_422 (O_422,N_2713,N_4336);
nor UO_423 (O_423,N_2901,N_2664);
nor UO_424 (O_424,N_4675,N_3773);
nand UO_425 (O_425,N_4267,N_4075);
nand UO_426 (O_426,N_2796,N_4953);
and UO_427 (O_427,N_3041,N_3909);
and UO_428 (O_428,N_3281,N_4599);
and UO_429 (O_429,N_4929,N_4392);
nor UO_430 (O_430,N_4316,N_4385);
nor UO_431 (O_431,N_2593,N_4771);
or UO_432 (O_432,N_3625,N_2734);
and UO_433 (O_433,N_4523,N_4708);
and UO_434 (O_434,N_2512,N_4250);
and UO_435 (O_435,N_3126,N_3930);
and UO_436 (O_436,N_2509,N_3768);
or UO_437 (O_437,N_3456,N_4084);
or UO_438 (O_438,N_4606,N_4213);
nor UO_439 (O_439,N_3397,N_3024);
or UO_440 (O_440,N_3129,N_2751);
nand UO_441 (O_441,N_4635,N_2924);
nand UO_442 (O_442,N_4779,N_4189);
xor UO_443 (O_443,N_3259,N_3469);
nand UO_444 (O_444,N_3285,N_3439);
nor UO_445 (O_445,N_3679,N_3653);
or UO_446 (O_446,N_4131,N_4279);
nor UO_447 (O_447,N_4408,N_3494);
or UO_448 (O_448,N_3736,N_3086);
nand UO_449 (O_449,N_4506,N_4957);
nor UO_450 (O_450,N_3459,N_2640);
and UO_451 (O_451,N_4760,N_2830);
or UO_452 (O_452,N_3252,N_3967);
nor UO_453 (O_453,N_4031,N_3338);
nor UO_454 (O_454,N_4976,N_4722);
or UO_455 (O_455,N_4934,N_3733);
or UO_456 (O_456,N_3582,N_4227);
or UO_457 (O_457,N_4839,N_3172);
nor UO_458 (O_458,N_2533,N_4415);
nor UO_459 (O_459,N_4193,N_2996);
and UO_460 (O_460,N_3682,N_4831);
and UO_461 (O_461,N_4299,N_4074);
nor UO_462 (O_462,N_3894,N_3538);
or UO_463 (O_463,N_4836,N_4387);
or UO_464 (O_464,N_4653,N_3344);
and UO_465 (O_465,N_4355,N_4660);
and UO_466 (O_466,N_4088,N_4504);
nor UO_467 (O_467,N_4678,N_4476);
and UO_468 (O_468,N_3160,N_4281);
nand UO_469 (O_469,N_4362,N_4994);
nor UO_470 (O_470,N_2561,N_3138);
xor UO_471 (O_471,N_4018,N_3153);
nor UO_472 (O_472,N_4240,N_4634);
xnor UO_473 (O_473,N_4109,N_3960);
nor UO_474 (O_474,N_4517,N_3096);
nand UO_475 (O_475,N_4808,N_4376);
nand UO_476 (O_476,N_3045,N_3374);
and UO_477 (O_477,N_3744,N_3396);
nand UO_478 (O_478,N_3672,N_2766);
and UO_479 (O_479,N_3859,N_4087);
nor UO_480 (O_480,N_3785,N_3940);
nor UO_481 (O_481,N_4137,N_3622);
or UO_482 (O_482,N_4219,N_4960);
or UO_483 (O_483,N_4350,N_4432);
nor UO_484 (O_484,N_2675,N_3454);
and UO_485 (O_485,N_3885,N_3347);
or UO_486 (O_486,N_4843,N_4749);
or UO_487 (O_487,N_2812,N_4981);
or UO_488 (O_488,N_4884,N_2980);
or UO_489 (O_489,N_3100,N_4224);
nor UO_490 (O_490,N_3191,N_3429);
nor UO_491 (O_491,N_4781,N_4102);
nor UO_492 (O_492,N_3814,N_3284);
and UO_493 (O_493,N_3204,N_3268);
or UO_494 (O_494,N_4096,N_3276);
and UO_495 (O_495,N_3724,N_4603);
nand UO_496 (O_496,N_4964,N_3951);
nor UO_497 (O_497,N_3452,N_4474);
and UO_498 (O_498,N_2609,N_3541);
or UO_499 (O_499,N_2888,N_4715);
or UO_500 (O_500,N_4803,N_3844);
nor UO_501 (O_501,N_2626,N_4864);
or UO_502 (O_502,N_3053,N_4195);
or UO_503 (O_503,N_3111,N_3084);
or UO_504 (O_504,N_2975,N_3993);
or UO_505 (O_505,N_2715,N_4520);
or UO_506 (O_506,N_2991,N_4427);
nor UO_507 (O_507,N_2522,N_4527);
nand UO_508 (O_508,N_4417,N_3081);
xor UO_509 (O_509,N_4561,N_3482);
nand UO_510 (O_510,N_4001,N_2740);
nand UO_511 (O_511,N_3610,N_4271);
and UO_512 (O_512,N_4720,N_3331);
and UO_513 (O_513,N_2634,N_4924);
or UO_514 (O_514,N_3821,N_4083);
or UO_515 (O_515,N_4817,N_3994);
or UO_516 (O_516,N_3402,N_3754);
nor UO_517 (O_517,N_3939,N_4816);
or UO_518 (O_518,N_4645,N_3742);
or UO_519 (O_519,N_3327,N_2638);
or UO_520 (O_520,N_3395,N_2647);
and UO_521 (O_521,N_3921,N_4724);
nand UO_522 (O_522,N_3417,N_4234);
or UO_523 (O_523,N_3490,N_2897);
and UO_524 (O_524,N_4780,N_3641);
nor UO_525 (O_525,N_4150,N_4501);
or UO_526 (O_526,N_2947,N_3472);
nand UO_527 (O_527,N_4978,N_2513);
nor UO_528 (O_528,N_4265,N_4371);
and UO_529 (O_529,N_4029,N_4490);
xor UO_530 (O_530,N_2891,N_4962);
or UO_531 (O_531,N_4346,N_3400);
or UO_532 (O_532,N_4679,N_3609);
nand UO_533 (O_533,N_2844,N_4777);
nand UO_534 (O_534,N_3640,N_3378);
nand UO_535 (O_535,N_4844,N_4933);
and UO_536 (O_536,N_2882,N_2775);
nor UO_537 (O_537,N_2871,N_2971);
nor UO_538 (O_538,N_4773,N_2787);
and UO_539 (O_539,N_4825,N_4525);
nand UO_540 (O_540,N_4988,N_4251);
or UO_541 (O_541,N_4703,N_4581);
nand UO_542 (O_542,N_3426,N_4939);
or UO_543 (O_543,N_3372,N_4027);
nand UO_544 (O_544,N_4909,N_4746);
nand UO_545 (O_545,N_2636,N_2565);
nand UO_546 (O_546,N_3485,N_2611);
nand UO_547 (O_547,N_3342,N_3562);
nor UO_548 (O_548,N_4896,N_4151);
nand UO_549 (O_549,N_3280,N_3707);
nor UO_550 (O_550,N_4003,N_2730);
nor UO_551 (O_551,N_2649,N_2718);
or UO_552 (O_552,N_2527,N_3496);
nand UO_553 (O_553,N_2594,N_3254);
nand UO_554 (O_554,N_2549,N_4080);
and UO_555 (O_555,N_2506,N_2809);
nor UO_556 (O_556,N_3313,N_3237);
or UO_557 (O_557,N_2556,N_3251);
and UO_558 (O_558,N_2575,N_3190);
nand UO_559 (O_559,N_4447,N_4302);
nor UO_560 (O_560,N_3102,N_2599);
nor UO_561 (O_561,N_4609,N_4676);
or UO_562 (O_562,N_2959,N_4364);
nor UO_563 (O_563,N_4256,N_3789);
nor UO_564 (O_564,N_3843,N_2747);
nand UO_565 (O_565,N_3503,N_4082);
nor UO_566 (O_566,N_3036,N_4277);
and UO_567 (O_567,N_3747,N_2514);
nor UO_568 (O_568,N_4941,N_2870);
nand UO_569 (O_569,N_4865,N_2990);
and UO_570 (O_570,N_2861,N_4805);
and UO_571 (O_571,N_3699,N_2938);
or UO_572 (O_572,N_4202,N_3200);
nand UO_573 (O_573,N_4208,N_2973);
and UO_574 (O_574,N_2985,N_3542);
nand UO_575 (O_575,N_4368,N_2699);
and UO_576 (O_576,N_2923,N_4170);
xor UO_577 (O_577,N_4155,N_3205);
and UO_578 (O_578,N_4689,N_3907);
xnor UO_579 (O_579,N_2585,N_3216);
xor UO_580 (O_580,N_4294,N_3711);
nor UO_581 (O_581,N_3637,N_4623);
nor UO_582 (O_582,N_4324,N_4516);
nand UO_583 (O_583,N_3514,N_2645);
or UO_584 (O_584,N_3405,N_2741);
or UO_585 (O_585,N_3491,N_4048);
nand UO_586 (O_586,N_3683,N_3873);
or UO_587 (O_587,N_4856,N_3923);
and UO_588 (O_588,N_3403,N_4946);
nor UO_589 (O_589,N_3493,N_4680);
nand UO_590 (O_590,N_4260,N_2677);
or UO_591 (O_591,N_4296,N_2858);
or UO_592 (O_592,N_4693,N_4681);
nand UO_593 (O_593,N_4713,N_2902);
or UO_594 (O_594,N_4113,N_4152);
or UO_595 (O_595,N_2847,N_4469);
nand UO_596 (O_596,N_3753,N_3575);
nand UO_597 (O_597,N_2589,N_4333);
nand UO_598 (O_598,N_2641,N_3752);
or UO_599 (O_599,N_3411,N_3380);
nor UO_600 (O_600,N_3371,N_3798);
nor UO_601 (O_601,N_3684,N_2746);
or UO_602 (O_602,N_2665,N_2644);
or UO_603 (O_603,N_4855,N_3555);
and UO_604 (O_604,N_4372,N_3659);
xor UO_605 (O_605,N_3422,N_4244);
nor UO_606 (O_606,N_4276,N_3953);
nand UO_607 (O_607,N_4721,N_3329);
or UO_608 (O_608,N_4488,N_2815);
nor UO_609 (O_609,N_4091,N_3003);
and UO_610 (O_610,N_3340,N_4917);
nor UO_611 (O_611,N_2846,N_3154);
nor UO_612 (O_612,N_3908,N_2725);
or UO_613 (O_613,N_3290,N_4025);
nand UO_614 (O_614,N_4192,N_3273);
nand UO_615 (O_615,N_3563,N_4343);
or UO_616 (O_616,N_4120,N_3354);
or UO_617 (O_617,N_4546,N_4545);
or UO_618 (O_618,N_3188,N_2834);
nand UO_619 (O_619,N_3315,N_2526);
nor UO_620 (O_620,N_3308,N_3698);
and UO_621 (O_621,N_4903,N_4185);
nor UO_622 (O_622,N_2578,N_3757);
and UO_623 (O_623,N_3302,N_2951);
nor UO_624 (O_624,N_4433,N_4587);
xor UO_625 (O_625,N_4725,N_4067);
nand UO_626 (O_626,N_3145,N_4963);
and UO_627 (O_627,N_4077,N_4627);
and UO_628 (O_628,N_4538,N_3443);
and UO_629 (O_629,N_2573,N_3178);
xnor UO_630 (O_630,N_3680,N_3343);
nor UO_631 (O_631,N_2911,N_2781);
and UO_632 (O_632,N_4716,N_3533);
and UO_633 (O_633,N_3775,N_3580);
nand UO_634 (O_634,N_4510,N_3052);
and UO_635 (O_635,N_2817,N_3687);
nand UO_636 (O_636,N_3419,N_3675);
or UO_637 (O_637,N_2739,N_4130);
or UO_638 (O_638,N_3833,N_3739);
nand UO_639 (O_639,N_3648,N_4763);
nand UO_640 (O_640,N_3662,N_4973);
and UO_641 (O_641,N_3432,N_4802);
nand UO_642 (O_642,N_3513,N_3802);
xor UO_643 (O_643,N_4347,N_4897);
or UO_644 (O_644,N_4325,N_2701);
or UO_645 (O_645,N_4692,N_2530);
or UO_646 (O_646,N_3283,N_4961);
nand UO_647 (O_647,N_4540,N_3246);
nor UO_648 (O_648,N_4984,N_4317);
nand UO_649 (O_649,N_4797,N_4845);
nor UO_650 (O_650,N_2887,N_4290);
nand UO_651 (O_651,N_4305,N_2970);
and UO_652 (O_652,N_2895,N_4475);
nand UO_653 (O_653,N_4167,N_3536);
nor UO_654 (O_654,N_2986,N_4028);
and UO_655 (O_655,N_4116,N_3035);
or UO_656 (O_656,N_2537,N_4402);
nand UO_657 (O_657,N_2988,N_4162);
nor UO_658 (O_658,N_4138,N_2720);
and UO_659 (O_659,N_3099,N_4314);
and UO_660 (O_660,N_4245,N_2753);
or UO_661 (O_661,N_4775,N_3282);
nor UO_662 (O_662,N_3050,N_3022);
nor UO_663 (O_663,N_4287,N_4413);
nand UO_664 (O_664,N_2719,N_2592);
nand UO_665 (O_665,N_2584,N_2913);
nand UO_666 (O_666,N_2692,N_4754);
nand UO_667 (O_667,N_3013,N_4868);
and UO_668 (O_668,N_4163,N_2873);
nand UO_669 (O_669,N_4268,N_2567);
or UO_670 (O_670,N_3570,N_3674);
nand UO_671 (O_671,N_3578,N_4437);
nor UO_672 (O_672,N_3087,N_2798);
and UO_673 (O_673,N_3447,N_4292);
nor UO_674 (O_674,N_3197,N_2880);
or UO_675 (O_675,N_3128,N_3975);
and UO_676 (O_676,N_3310,N_2563);
and UO_677 (O_677,N_4927,N_3972);
or UO_678 (O_678,N_4752,N_2919);
and UO_679 (O_679,N_4881,N_4541);
or UO_680 (O_680,N_2554,N_2783);
and UO_681 (O_681,N_3455,N_2681);
or UO_682 (O_682,N_3353,N_2840);
nor UO_683 (O_683,N_3571,N_2962);
xor UO_684 (O_684,N_3217,N_4153);
or UO_685 (O_685,N_4099,N_4248);
nand UO_686 (O_686,N_3385,N_3690);
or UO_687 (O_687,N_4095,N_4275);
nor UO_688 (O_688,N_3532,N_3554);
or UO_689 (O_689,N_4911,N_4117);
or UO_690 (O_690,N_2707,N_3959);
or UO_691 (O_691,N_4617,N_4266);
nor UO_692 (O_692,N_3000,N_3381);
and UO_693 (O_693,N_4885,N_4862);
nor UO_694 (O_694,N_4795,N_3039);
nor UO_695 (O_695,N_4467,N_4285);
or UO_696 (O_696,N_3592,N_4667);
nor UO_697 (O_697,N_2816,N_3560);
or UO_698 (O_698,N_3585,N_3826);
and UO_699 (O_699,N_3927,N_4768);
nor UO_700 (O_700,N_2756,N_3317);
or UO_701 (O_701,N_2788,N_4669);
or UO_702 (O_702,N_2931,N_2852);
or UO_703 (O_703,N_4611,N_3360);
xor UO_704 (O_704,N_4121,N_3042);
nor UO_705 (O_705,N_2765,N_2744);
nand UO_706 (O_706,N_3577,N_2883);
and UO_707 (O_707,N_4269,N_3702);
nor UO_708 (O_708,N_3847,N_3528);
nand UO_709 (O_709,N_2969,N_4041);
nor UO_710 (O_710,N_3638,N_2841);
or UO_711 (O_711,N_4070,N_2927);
nand UO_712 (O_712,N_3534,N_2898);
nand UO_713 (O_713,N_3976,N_4366);
nand UO_714 (O_714,N_4876,N_2654);
or UO_715 (O_715,N_4705,N_4788);
nand UO_716 (O_716,N_2950,N_3031);
and UO_717 (O_717,N_3366,N_4622);
nor UO_718 (O_718,N_4442,N_4076);
or UO_719 (O_719,N_4044,N_3358);
nor UO_720 (O_720,N_4398,N_3301);
nand UO_721 (O_721,N_4604,N_3261);
or UO_722 (O_722,N_2999,N_3928);
nand UO_723 (O_723,N_4135,N_3248);
or UO_724 (O_724,N_2818,N_2700);
and UO_725 (O_725,N_4646,N_4174);
or UO_726 (O_726,N_2535,N_4247);
and UO_727 (O_727,N_3124,N_3337);
and UO_728 (O_728,N_2886,N_3943);
and UO_729 (O_729,N_4010,N_4935);
or UO_730 (O_730,N_4914,N_2521);
and UO_731 (O_731,N_4975,N_3361);
or UO_732 (O_732,N_3476,N_3264);
xnor UO_733 (O_733,N_3236,N_3388);
nor UO_734 (O_734,N_4769,N_4128);
nand UO_735 (O_735,N_3293,N_3304);
nand UO_736 (O_736,N_3346,N_4238);
nand UO_737 (O_737,N_2778,N_3838);
xnor UO_738 (O_738,N_4022,N_3019);
nor UO_739 (O_739,N_3139,N_3782);
or UO_740 (O_740,N_3104,N_3881);
or UO_741 (O_741,N_4178,N_3708);
nor UO_742 (O_742,N_4187,N_4496);
and UO_743 (O_743,N_2564,N_4341);
nor UO_744 (O_744,N_4380,N_4853);
and UO_745 (O_745,N_4701,N_3113);
nand UO_746 (O_746,N_4090,N_2670);
or UO_747 (O_747,N_4840,N_2685);
nand UO_748 (O_748,N_3260,N_3522);
nand UO_749 (O_749,N_2705,N_4310);
nor UO_750 (O_750,N_3451,N_4013);
or UO_751 (O_751,N_4531,N_3368);
nand UO_752 (O_752,N_3147,N_4007);
or UO_753 (O_753,N_3623,N_4046);
nor UO_754 (O_754,N_3703,N_4492);
or UO_755 (O_755,N_4053,N_4827);
and UO_756 (O_756,N_4875,N_4586);
nand UO_757 (O_757,N_3287,N_3906);
or UO_758 (O_758,N_3784,N_3202);
and UO_759 (O_759,N_4210,N_2952);
and UO_760 (O_760,N_2721,N_3999);
or UO_761 (O_761,N_2629,N_4700);
nand UO_762 (O_762,N_3169,N_4133);
nand UO_763 (O_763,N_4156,N_4995);
nor UO_764 (O_764,N_3769,N_3351);
nor UO_765 (O_765,N_2655,N_3530);
nor UO_766 (O_766,N_4772,N_2968);
and UO_767 (O_767,N_2904,N_3474);
and UO_768 (O_768,N_4329,N_3689);
or UO_769 (O_769,N_4233,N_4776);
and UO_770 (O_770,N_4002,N_3987);
nand UO_771 (O_771,N_3920,N_4534);
nor UO_772 (O_772,N_3055,N_3971);
nor UO_773 (O_773,N_3118,N_4487);
and UO_774 (O_774,N_4980,N_2771);
and UO_775 (O_775,N_3954,N_4882);
and UO_776 (O_776,N_2625,N_4588);
nor UO_777 (O_777,N_2862,N_4094);
nand UO_778 (O_778,N_2505,N_2750);
and UO_779 (O_779,N_3932,N_2667);
nand UO_780 (O_780,N_3082,N_3978);
nor UO_781 (O_781,N_4632,N_4736);
nor UO_782 (O_782,N_3098,N_3115);
nand UO_783 (O_783,N_3225,N_4159);
or UO_784 (O_784,N_3519,N_4966);
and UO_785 (O_785,N_3335,N_3759);
or UO_786 (O_786,N_4212,N_4753);
and UO_787 (O_787,N_3296,N_4412);
and UO_788 (O_788,N_3646,N_4596);
nand UO_789 (O_789,N_4228,N_3925);
and UO_790 (O_790,N_3047,N_4282);
and UO_791 (O_791,N_4455,N_4351);
and UO_792 (O_792,N_4008,N_3918);
and UO_793 (O_793,N_2942,N_4142);
and UO_794 (O_794,N_3214,N_4330);
nand UO_795 (O_795,N_4345,N_4664);
nor UO_796 (O_796,N_4393,N_2576);
or UO_797 (O_797,N_3394,N_4063);
nor UO_798 (O_798,N_4794,N_4444);
or UO_799 (O_799,N_4215,N_2761);
or UO_800 (O_800,N_3620,N_3185);
and UO_801 (O_801,N_3897,N_4562);
and UO_802 (O_802,N_4796,N_2630);
nor UO_803 (O_803,N_4489,N_4037);
nand UO_804 (O_804,N_4243,N_4511);
or UO_805 (O_805,N_4161,N_3521);
or UO_806 (O_806,N_3746,N_3030);
xor UO_807 (O_807,N_3594,N_2827);
or UO_808 (O_808,N_2868,N_4706);
or UO_809 (O_809,N_4401,N_4965);
and UO_810 (O_810,N_3253,N_4948);
nand UO_811 (O_811,N_3876,N_4550);
and UO_812 (O_812,N_2845,N_2710);
nor UO_813 (O_813,N_4348,N_3021);
nand UO_814 (O_814,N_3696,N_4005);
xnor UO_815 (O_815,N_2837,N_2928);
nor UO_816 (O_816,N_4357,N_4690);
or UO_817 (O_817,N_3979,N_2875);
and UO_818 (O_818,N_2724,N_4396);
or UO_819 (O_819,N_3630,N_2618);
nand UO_820 (O_820,N_4406,N_3136);
nor UO_821 (O_821,N_4331,N_2906);
nand UO_822 (O_822,N_2768,N_4956);
nand UO_823 (O_823,N_4332,N_3547);
and UO_824 (O_824,N_3101,N_4688);
nor UO_825 (O_825,N_3201,N_2749);
nand UO_826 (O_826,N_2697,N_3751);
nand UO_827 (O_827,N_3776,N_4813);
nand UO_828 (O_828,N_4811,N_3797);
and UO_829 (O_829,N_3586,N_3836);
or UO_830 (O_830,N_3957,N_4589);
and UO_831 (O_831,N_2920,N_3760);
and UO_832 (O_832,N_4050,N_4872);
and UO_833 (O_833,N_3667,N_3786);
nor UO_834 (O_834,N_3271,N_3933);
nor UO_835 (O_835,N_3915,N_3442);
nor UO_836 (O_836,N_4631,N_2702);
or UO_837 (O_837,N_3377,N_4629);
and UO_838 (O_838,N_3498,N_2587);
nor UO_839 (O_839,N_3165,N_3040);
nor UO_840 (O_840,N_4637,N_4045);
or UO_841 (O_841,N_3433,N_4959);
or UO_842 (O_842,N_4895,N_3025);
and UO_843 (O_843,N_4783,N_3067);
and UO_844 (O_844,N_4710,N_4539);
xor UO_845 (O_845,N_3764,N_2896);
nor UO_846 (O_846,N_3435,N_3816);
or UO_847 (O_847,N_2983,N_3706);
or UO_848 (O_848,N_4873,N_3152);
nand UO_849 (O_849,N_3420,N_4641);
nor UO_850 (O_850,N_2994,N_4951);
nor UO_851 (O_851,N_4744,N_4572);
nand UO_852 (O_852,N_4060,N_2964);
and UO_853 (O_853,N_2616,N_3823);
or UO_854 (O_854,N_3678,N_4261);
xor UO_855 (O_855,N_3048,N_3056);
nand UO_856 (O_856,N_4379,N_2540);
xor UO_857 (O_857,N_3701,N_2735);
and UO_858 (O_858,N_4186,N_3080);
or UO_859 (O_859,N_4180,N_2953);
or UO_860 (O_860,N_3295,N_3527);
nand UO_861 (O_861,N_3837,N_4943);
nor UO_862 (O_862,N_4039,N_3473);
nor UO_863 (O_863,N_2657,N_3274);
and UO_864 (O_864,N_2770,N_3054);
nor UO_865 (O_865,N_4337,N_4093);
nor UO_866 (O_866,N_3963,N_3942);
and UO_867 (O_867,N_2944,N_3550);
nand UO_868 (O_868,N_3579,N_2792);
and UO_869 (O_869,N_4255,N_3026);
and UO_870 (O_870,N_3913,N_2934);
or UO_871 (O_871,N_4111,N_4062);
nor UO_872 (O_872,N_4858,N_3161);
nor UO_873 (O_873,N_4198,N_3207);
or UO_874 (O_874,N_4774,N_4249);
nand UO_875 (O_875,N_3219,N_4441);
nor UO_876 (O_876,N_3788,N_4327);
or UO_877 (O_877,N_3130,N_3479);
nand UO_878 (O_878,N_2804,N_4241);
or UO_879 (O_879,N_3780,N_4640);
nor UO_880 (O_880,N_4127,N_3064);
nand UO_881 (O_881,N_3539,N_4945);
nand UO_882 (O_882,N_3094,N_2881);
nor UO_883 (O_883,N_2631,N_4654);
nand UO_884 (O_884,N_3825,N_4747);
nand UO_885 (O_885,N_3756,N_3879);
and UO_886 (O_886,N_3345,N_3410);
nor UO_887 (O_887,N_4601,N_4630);
nor UO_888 (O_888,N_3818,N_4616);
nor UO_889 (O_889,N_4259,N_3428);
or UO_890 (O_890,N_4655,N_2586);
nor UO_891 (O_891,N_4544,N_2525);
and UO_892 (O_892,N_3158,N_3958);
nor UO_893 (O_893,N_3615,N_2793);
xor UO_894 (O_894,N_4431,N_3244);
nor UO_895 (O_895,N_3008,N_3599);
nor UO_896 (O_896,N_2731,N_2557);
or UO_897 (O_897,N_2642,N_4728);
and UO_898 (O_898,N_3559,N_4559);
and UO_899 (O_899,N_3279,N_3899);
nor UO_900 (O_900,N_4491,N_3658);
nand UO_901 (O_901,N_2780,N_3486);
nand UO_902 (O_902,N_3564,N_4226);
or UO_903 (O_903,N_3027,N_2523);
and UO_904 (O_904,N_4519,N_3502);
or UO_905 (O_905,N_3007,N_4950);
nor UO_906 (O_906,N_3135,N_2992);
nand UO_907 (O_907,N_3549,N_4651);
and UO_908 (O_908,N_2653,N_4497);
or UO_909 (O_909,N_3713,N_2963);
nand UO_910 (O_910,N_4977,N_3998);
nor UO_911 (O_911,N_4499,N_4888);
nand UO_912 (O_912,N_2646,N_3581);
xor UO_913 (O_913,N_4580,N_4049);
nor UO_914 (O_914,N_4014,N_4230);
or UO_915 (O_915,N_3692,N_2722);
and UO_916 (O_916,N_3990,N_4833);
or UO_917 (O_917,N_3985,N_4600);
nor UO_918 (O_918,N_2748,N_2759);
or UO_919 (O_919,N_4122,N_2574);
nor UO_920 (O_920,N_4110,N_4509);
or UO_921 (O_921,N_3168,N_3878);
nand UO_922 (O_922,N_4321,N_3795);
and UO_923 (O_923,N_2956,N_3613);
nor UO_924 (O_924,N_4438,N_2800);
or UO_925 (O_925,N_4081,N_4353);
nor UO_926 (O_926,N_2974,N_4000);
nand UO_927 (O_927,N_3660,N_4625);
nand UO_928 (O_928,N_3015,N_2910);
nand UO_929 (O_929,N_4123,N_3148);
nand UO_930 (O_930,N_3916,N_3448);
nor UO_931 (O_931,N_4295,N_4272);
or UO_932 (O_932,N_2925,N_2801);
nand UO_933 (O_933,N_4424,N_3882);
and UO_934 (O_934,N_2582,N_2876);
nor UO_935 (O_935,N_4552,N_4923);
nand UO_936 (O_936,N_4181,N_3413);
and UO_937 (O_937,N_4288,N_3952);
and UO_938 (O_938,N_4182,N_2784);
or UO_939 (O_939,N_2726,N_2550);
nor UO_940 (O_940,N_3874,N_4762);
and UO_941 (O_941,N_4453,N_3365);
nor UO_942 (O_942,N_4578,N_3817);
and UO_943 (O_943,N_3886,N_4410);
and UO_944 (O_944,N_3657,N_3390);
nand UO_945 (O_945,N_3046,N_4205);
and UO_946 (O_946,N_3525,N_4673);
or UO_947 (O_947,N_3436,N_3893);
nand UO_948 (O_948,N_3195,N_2997);
nand UO_949 (O_949,N_3133,N_3693);
nor UO_950 (O_950,N_3905,N_4598);
or UO_951 (O_951,N_4809,N_3463);
or UO_952 (O_952,N_3038,N_3312);
and UO_953 (O_953,N_4648,N_3815);
or UO_954 (O_954,N_4414,N_4030);
and UO_955 (O_955,N_3598,N_3924);
and UO_956 (O_956,N_3986,N_4859);
nand UO_957 (O_957,N_3804,N_4466);
or UO_958 (O_958,N_3483,N_2820);
and UO_959 (O_959,N_2698,N_3668);
or UO_960 (O_960,N_4835,N_4498);
nand UO_961 (O_961,N_4674,N_4124);
nand UO_962 (O_962,N_2860,N_2984);
and UO_963 (O_963,N_2758,N_4220);
nand UO_964 (O_964,N_3286,N_3673);
and UO_965 (O_965,N_2551,N_4242);
or UO_966 (O_966,N_4912,N_4565);
or UO_967 (O_967,N_4298,N_2903);
and UO_968 (O_968,N_3661,N_4280);
nand UO_969 (O_969,N_3778,N_2899);
or UO_970 (O_970,N_4485,N_3255);
or UO_971 (O_971,N_3356,N_3596);
and UO_972 (O_972,N_3132,N_2799);
nor UO_973 (O_973,N_3569,N_2810);
or UO_974 (O_974,N_4723,N_4818);
xor UO_975 (O_975,N_4554,N_3717);
and UO_976 (O_976,N_3561,N_3228);
nand UO_977 (O_977,N_3624,N_3418);
and UO_978 (O_978,N_2648,N_4483);
nor UO_979 (O_979,N_4560,N_3091);
nor UO_980 (O_980,N_4383,N_4806);
nand UO_981 (O_981,N_3323,N_2998);
or UO_982 (O_982,N_3198,N_4597);
nand UO_983 (O_983,N_3382,N_4403);
nand UO_984 (O_984,N_4575,N_2884);
nor UO_985 (O_985,N_3854,N_2559);
nor UO_986 (O_986,N_3548,N_3705);
or UO_987 (O_987,N_4618,N_4179);
nor UO_988 (O_988,N_4503,N_3218);
or UO_989 (O_989,N_4024,N_4590);
and UO_990 (O_990,N_2528,N_4112);
nand UO_991 (O_991,N_2833,N_3803);
and UO_992 (O_992,N_4925,N_4871);
and UO_993 (O_993,N_3348,N_4829);
nor UO_994 (O_994,N_3829,N_3142);
nor UO_995 (O_995,N_4528,N_4126);
and UO_996 (O_996,N_4691,N_3590);
or UO_997 (O_997,N_2790,N_2591);
and UO_998 (O_998,N_2511,N_4571);
or UO_999 (O_999,N_2823,N_3656);
endmodule